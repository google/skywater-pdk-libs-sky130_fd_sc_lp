* File: sky130_fd_sc_lp__einvn_0.spice
* Created: Fri Aug 28 10:32:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvn_0.pex.spice"
.subckt sky130_fd_sc_lp__einvn_0  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_TE_B_M1004_g N_A_28_141#_M1004_s VNB NSHORT L=0.15
+ W=0.42 AD=0.08715 AS=0.1113 PD=0.835 PS=1.37 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 A_224_141# N_A_28_141#_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.08715 PD=0.66 PS=0.835 NRD=18.564 NRS=18.564 M=1 R=2.8
+ SA=75000.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_Z_M1002_d N_A_M1002_g A_224_141# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_TE_B_M1001_g N_A_28_141#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0855057 AS=0.1197 PD=0.80434 PS=1.41 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 A_224_481# N_TE_B_M1003_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.130294 PD=0.88 PS=1.22566 NRD=19.9955 NRS=9.9879 M=1 R=4.26667
+ SA=75000.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_Z_M1000_d N_A_M1000_g A_224_481# VPB PHIGHVT L=0.15 W=0.64 AD=0.1696
+ AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75000.9
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.2895 P=8.33
*
.include "sky130_fd_sc_lp__einvn_0.pxi.spice"
*
.ends
*
*
