* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__einvp_8 A TE VGND VNB VPB VPWR Z
X0 VGND TE a_371_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_371_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 Z A a_365_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_365_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 Z A a_371_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_365_367# a_182_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VPWR a_182_367# a_365_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_365_367# a_182_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_371_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VGND TE a_371_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VGND TE a_371_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VPWR TE a_182_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND TE a_182_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_371_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_365_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_371_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 Z A a_365_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VGND TE a_371_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_371_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_371_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_365_367# a_182_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VPWR a_182_367# a_365_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 Z A a_371_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 VPWR a_182_367# a_365_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_365_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 Z A a_365_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 VPWR a_182_367# a_365_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 a_365_367# a_182_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 a_371_47# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 Z A a_371_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 Z A a_365_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_365_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_371_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 Z A a_371_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
