* File: sky130_fd_sc_lp__einvn_m.spice
* Created: Fri Aug 28 10:33:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvn_m.pex.spice"
.subckt sky130_fd_sc_lp__einvn_m  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_TE_B_M1004_g N_A_47_154#_M1004_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0609 AS=0.1113 PD=0.71 PS=1.37 NRD=2.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 A_218_154# N_A_47_154#_M1000_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0609 PD=0.7 PS=0.71 NRD=24.276 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g A_218_154# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=24.276 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_TE_B_M1002_g N_A_47_154#_M1002_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 A_232_535# N_TE_B_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_Z_M1003_d N_A_M1003_g A_232_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.2895 P=8.33
*
.include "sky130_fd_sc_lp__einvn_m.pxi.spice"
*
.ends
*
*
