* File: sky130_fd_sc_lp__xnor2_m.pex.spice
* Created: Fri Aug 28 11:35:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XNOR2_M%A 3 5 7 11 15 19 23 25 27 36
c46 19 0 1.94133e-19 $X=1.195 $Y=1.28
c47 11 0 7.24622e-20 $X=1.41 $Y=0.66
c48 7 0 1.9934e-19 $X=1.05 $Y=2.32
r49 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.29
+ $Y=1.295 $X2=1.29 $Y2=1.295
r50 27 37 8.63834 $w=5.38e-07 $l=3.9e-07 $layer=LI1_cond $X=1.68 $Y=1.48
+ $X2=1.29 $Y2=1.48
r51 25 37 1.99346 $w=5.38e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.48 $X2=1.29
+ $Y2=1.48
r52 23 25 10.6318 $w=5.38e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.48 $X2=1.2
+ $Y2=1.48
r53 21 36 37.2422 $w=5.1e-07 $l=3.55e-07 $layer=POLY_cond $X=1.23 $Y=1.65
+ $X2=1.23 $Y2=1.295
r54 19 36 1.57362 $w=5.1e-07 $l=1.5e-08 $layer=POLY_cond $X=1.23 $Y=1.28
+ $X2=1.23 $Y2=1.295
r55 5 21 24.7327 $w=5.1e-07 $l=1.5e-07 $layer=POLY_cond $X=1.265 $Y=1.8
+ $X2=1.265 $Y2=1.65
r56 5 15 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.48 $Y=1.8 $X2=1.48
+ $Y2=2.32
r57 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.05 $Y=1.8 $X2=1.05
+ $Y2=2.32
r58 1 19 24.7327 $w=5.1e-07 $l=1.5e-07 $layer=POLY_cond $X=1.195 $Y=1.13
+ $X2=1.195 $Y2=1.28
r59 1 11 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.41 $Y=1.13 $X2=1.41
+ $Y2=0.66
r60 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.98 $Y=1.13 $X2=0.98
+ $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_M%B 3 6 7 8 11 14 15 16 17 22
c51 11 0 3.47049e-20 $X=1.84 $Y=0.66
c52 3 0 3.79214e-19 $X=0.62 $Y=0.66
r53 22 25 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.93 $Y=2.885 $X2=1.93
+ $Y2=2.975
r54 22 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.93 $Y=2.885
+ $X2=1.93 $Y2=2.72
r55 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=2.885 $X2=1.93 $Y2=2.885
r56 16 17 19.7562 $w=2.78e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.83
+ $X2=2.64 $Y2=2.83
r57 16 23 9.4665 $w=2.78e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=2.83 $X2=1.93
+ $Y2=2.83
r58 15 23 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=1.68 $Y=2.83
+ $X2=1.93 $Y2=2.83
r59 14 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.84 $Y=2.32 $X2=1.84
+ $Y2=2.72
r60 11 14 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=1.84 $Y=0.66
+ $X2=1.84 $Y2=2.32
r61 7 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=2.975
+ $X2=1.93 $Y2=2.975
r62 7 8 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.765 $Y=2.975
+ $X2=0.695 $Y2=2.975
r63 3 6 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=0.62 $Y=0.66 $X2=0.62
+ $Y2=2.32
r64 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.62 $Y=2.9
+ $X2=0.695 $Y2=2.975
r65 1 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.62 $Y=2.9 $X2=0.62
+ $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_M%A_56_90# 1 2 7 8 11 15 19 22 23 24 27 29 33
+ 34 39 41
c62 41 0 4.50749e-20 $X=0.835 $Y=2.015
c63 29 0 1.49058e-19 $X=2.205 $Y=2.015
c64 27 0 5.43989e-19 $X=0.835 $Y=2.255
r65 36 39 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=0.325 $Y=0.725
+ $X2=0.405 $Y2=0.725
r66 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.445 $X2=2.29 $Y2=1.445
r67 31 33 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.29 $Y=1.93
+ $X2=2.29 $Y2=1.445
r68 30 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=2.015
+ $X2=0.835 $Y2=2.015
r69 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.205 $Y=2.015
+ $X2=2.29 $Y2=1.93
r70 29 30 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=2.205 $Y=2.015
+ $X2=0.92 $Y2=2.015
r71 25 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=2.1
+ $X2=0.835 $Y2=2.015
r72 25 27 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.835 $Y=2.1
+ $X2=0.835 $Y2=2.255
r73 23 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.015
+ $X2=0.835 $Y2=2.015
r74 23 24 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.75 $Y=2.015
+ $X2=0.41 $Y2=2.015
r75 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.325 $Y=1.93
+ $X2=0.41 $Y2=2.015
r76 21 36 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.325 $Y=0.83
+ $X2=0.325 $Y2=0.725
r77 21 22 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=0.325 $Y=0.83
+ $X2=0.325 $Y2=1.93
r78 18 19 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=2.74 $Y=1.355
+ $X2=2.87 $Y2=1.355
r79 17 34 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.29 $Y=1.43
+ $X2=2.29 $Y2=1.445
r80 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.87 $Y=1.28
+ $X2=2.87 $Y2=1.355
r81 13 15 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.87 $Y=1.28
+ $X2=2.87 $Y2=0.66
r82 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.74 $Y=1.43 $X2=2.74
+ $Y2=1.355
r83 9 11 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2.74 $Y=1.43 $X2=2.74
+ $Y2=2.32
r84 8 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.455 $Y=1.355
+ $X2=2.29 $Y2=1.43
r85 7 18 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.665 $Y=1.355
+ $X2=2.74 $Y2=1.355
r86 7 8 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.665 $Y=1.355
+ $X2=2.455 $Y2=1.355
r87 2 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.695
+ $Y=2.11 $X2=0.835 $Y2=2.255
r88 1 39 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.28
+ $Y=0.45 $X2=0.405 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_M%VPWR 1 2 3 10 12 15 16 18 23 25 27 32 41 45
c37 23 0 1.79874e-19 $X=1.265 $Y=2.385
r38 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 36 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 33 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=1.185 $Y2=3.33
r44 33 35 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 32 44 3.49902 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=3.132 $Y2=3.33
r46 32 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 31 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 28 38 4.51706 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.285 $Y2=3.33
r51 28 30 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.57 $Y=3.33 $X2=0.72
+ $Y2=3.33
r52 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=1.185
+ $Y2=3.33
r53 27 30 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r54 25 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 25 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 20 23 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.185 $Y=2.385
+ $X2=1.265 $Y2=2.385
r57 16 44 3.34488 $w=1.9e-07 $l=1.69245e-07 $layer=LI1_cond $X=3 $Y=3.245
+ $X2=3.132 $Y2=3.33
r58 16 18 52.5359 $w=1.88e-07 $l=9e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.345
r59 15 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=3.33
r60 14 20 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.185 $Y=2.49
+ $X2=1.185 $Y2=2.385
r61 14 15 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.185 $Y=2.49
+ $X2=1.185 $Y2=3.245
r62 10 38 3.24911 $w=3.3e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.405 $Y=3.245
+ $X2=0.285 $Y2=3.33
r63 10 12 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=0.405 $Y=3.245
+ $X2=0.405 $Y2=2.385
r64 3 18 600 $w=1.7e-07 $l=3.10403e-07 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=2.11 $X2=2.99 $Y2=2.345
r65 2 23 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=2.11 $X2=1.265 $Y2=2.385
r66 1 12 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.28
+ $Y=2.11 $X2=0.405 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_M%Y 1 2 9 12 13 14 15 16 23
r25 16 23 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.64 $Y=2.385
+ $X2=2.64 $Y2=2.28
r26 16 34 7.29301 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.555 $Y=2.385
+ $X2=2.39 $Y2=2.385
r27 15 23 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.64 $Y=2.035
+ $X2=2.64 $Y2=2.28
r28 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=2.035
r29 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.665
r30 12 13 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=0.925
+ $X2=2.64 $Y2=1.295
r31 11 12 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.64 $Y=0.83
+ $X2=2.64 $Y2=0.925
r32 9 11 6.36683 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.655 $Y=0.725
+ $X2=2.655 $Y2=0.83
r33 2 34 600 $w=1.7e-07 $l=5.96867e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=2.11 $X2=2.39 $Y2=2.385
r34 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.45 $X2=2.655 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_M%VGND 1 2 10 11 12 14 18 20 27 28 31
c41 28 0 3.47049e-20 $X=3.12 $Y=0
r42 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 25 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.185
+ $Y2=0
r45 25 27 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.28 $Y=0 $X2=3.12
+ $Y2=0
r46 23 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r47 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 20 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.09 $Y=0 $X2=1.185
+ $Y2=0
r49 20 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.72
+ $Y2=0
r50 18 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r51 18 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r52 14 16 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.135 $Y=0.725
+ $X2=2.135 $Y2=0.945
r53 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=0.945
+ $X2=2.135 $Y2=0.945
r54 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.97 $Y=0.945
+ $X2=1.28 $Y2=0.945
r55 8 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.185 $Y=0.86
+ $X2=1.28 $Y2=0.945
r56 8 10 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.185 $Y=0.86
+ $X2=1.185 $Y2=0.725
r57 7 31 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r58 7 10 37.3589 $w=1.88e-07 $l=6.4e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.725
r59 2 14 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=1.915
+ $Y=0.45 $X2=2.135 $Y2=0.725
r60 1 10 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.055
+ $Y=0.45 $X2=1.195 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_M%A_297_90# 1 2 7 11 13
c18 7 0 7.24622e-20 $X=3 $Y=0.355
r19 13 16 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.625 $Y=0.355
+ $X2=1.625 $Y2=0.575
r20 9 11 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=3.095 $Y=0.44
+ $X2=3.095 $Y2=0.595
r21 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=0.355
+ $X2=1.625 $Y2=0.355
r22 7 9 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3 $Y=0.355
+ $X2=3.095 $Y2=0.44
r23 7 8 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3 $Y=0.355 $X2=1.79
+ $Y2=0.355
r24 2 11 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.45 $X2=3.085 $Y2=0.595
r25 1 16 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.45 $X2=1.625 $Y2=0.575
.ends

