* File: sky130_fd_sc_lp__ha_lp.pex.spice
* Created: Wed Sep  2 09:54:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__HA_LP%A_83_153# 1 2 9 12 15 19 21 27 28 32 37 39 41
+ 43
r70 34 37 4.24584 $w=3.78e-07 $l=1.4e-07 $layer=LI1_cond $X=1.415 $Y=0.455
+ $X2=1.555 $Y2=0.455
r71 30 32 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.87 $Y=1.895
+ $X2=1.87 $Y2=2.24
r72 29 39 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.5 $Y=1.81
+ $X2=1.415 $Y2=1.73
r73 28 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.705 $Y=1.81
+ $X2=1.87 $Y2=1.895
r74 28 29 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.705 $Y=1.81
+ $X2=1.5 $Y2=1.81
r75 27 39 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=1.565
+ $X2=1.415 $Y2=1.73
r76 26 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.415 $Y=0.645
+ $X2=1.415 $Y2=0.455
r77 26 27 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.415 $Y=0.645
+ $X2=1.415 $Y2=1.565
r78 24 43 6.32375 $w=3.65e-07 $l=4e-08 $layer=POLY_cond $X=1.035 $Y=1.747
+ $X2=1.075 $Y2=1.747
r79 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.035
+ $Y=1.73 $X2=1.035 $Y2=1.73
r80 21 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=1.73
+ $X2=1.415 $Y2=1.73
r81 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.33 $Y=1.73
+ $X2=1.035 $Y2=1.73
r82 17 43 11.667 $w=2.5e-07 $l=1.83e-07 $layer=POLY_cond $X=1.075 $Y=1.93
+ $X2=1.075 $Y2=1.747
r83 17 19 165.222 $w=2.5e-07 $l=6.65e-07 $layer=POLY_cond $X=1.075 $Y=1.93
+ $X2=1.075 $Y2=2.595
r84 13 24 29.2473 $w=3.65e-07 $l=1.85e-07 $layer=POLY_cond $X=0.85 $Y=1.747
+ $X2=1.035 $Y2=1.747
r85 13 41 32.4387 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.85 $Y=1.747
+ $X2=0.775 $Y2=1.747
r86 13 15 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.85 $Y=1.565
+ $X2=0.85 $Y2=1.105
r87 12 41 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.565 $Y=1.855
+ $X2=0.775 $Y2=1.855
r88 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.49 $Y=1.78
+ $X2=0.565 $Y2=1.855
r89 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.49 $Y=1.78 $X2=0.49
+ $Y2=1.105
r90 2 32 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.73
+ $Y=2.095 $X2=1.87 $Y2=2.24
r91 1 37 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.555 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__HA_LP%A_296_286# 1 2 7 9 13 17 21 25 27 31 33 34 39
+ 43 51 52 53 55 56
c132 33 0 9.89418e-20 $X=3.865 $Y=1.31
c133 9 0 1.20999e-19 $X=1.605 $Y=2.595
r134 56 59 66.9034 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=4.61 $Y=1.39
+ $X2=4.61 $Y2=1.895
r135 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.52
+ $Y=1.39 $X2=4.52 $Y2=1.39
r136 51 52 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.812 $Y=2.475
+ $X2=3.812 $Y2=2.31
r137 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.265 $X2=1.82 $Y2=1.265
r138 43 46 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=1.832 $Y=1.185
+ $X2=1.832 $Y2=1.265
r139 40 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=1.31
+ $X2=3.95 $Y2=1.31
r140 39 55 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=1.31
+ $X2=4.52 $Y2=1.31
r141 39 40 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.355 $Y=1.31
+ $X2=4.035 $Y2=1.31
r142 37 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=1.395
+ $X2=3.95 $Y2=1.31
r143 37 52 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=3.95 $Y=1.395
+ $X2=3.95 $Y2=2.31
r144 33 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=1.31
+ $X2=3.95 $Y2=1.31
r145 33 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.865 $Y=1.31
+ $X2=3.59 $Y2=1.31
r146 29 34 9.53671 $w=2.34e-07 $l=1.93959e-07 $layer=LI1_cond $X=3.425 $Y=1.247
+ $X2=3.59 $Y2=1.31
r147 29 31 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.425 $Y=1.1
+ $X2=3.425 $Y2=0.835
r148 28 43 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.985 $Y=1.185
+ $X2=1.832 $Y2=1.185
r149 27 29 9.53671 $w=2.34e-07 $l=1.93533e-07 $layer=LI1_cond $X=3.26 $Y=1.185
+ $X2=3.425 $Y2=1.247
r150 27 28 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=3.26 $Y=1.185
+ $X2=1.985 $Y2=1.185
r151 23 56 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=4.79 $Y=1.225
+ $X2=4.61 $Y2=1.39
r152 23 25 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.79 $Y=1.225
+ $X2=4.79 $Y2=0.835
r153 21 59 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=4.645 $Y=2.595
+ $X2=4.645 $Y2=1.895
r154 15 56 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=4.43 $Y=1.225
+ $X2=4.61 $Y2=1.39
r155 15 17 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.43 $Y=1.225
+ $X2=4.43 $Y2=0.835
r156 11 47 38.9379 $w=3.62e-07 $l=1.83016e-07 $layer=POLY_cond $X=1.77 $Y=1.1
+ $X2=1.732 $Y2=1.265
r157 11 13 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=1.77 $Y=1.1
+ $X2=1.77 $Y2=0.445
r158 7 47 43.27 $w=3.62e-07 $l=3.4775e-07 $layer=POLY_cond $X=1.605 $Y=1.555
+ $X2=1.732 $Y2=1.265
r159 7 9 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.605 $Y=1.555
+ $X2=1.605 $Y2=2.595
r160 2 51 300 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.615
+ $Y=2.095 $X2=3.755 $Y2=2.475
r161 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.625 $X2=3.425 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__HA_LP%B 3 8 12 18 19 20 21 22 25 26 28 32 33 36 37
+ 38 42 45
c109 36 0 1.20999e-19 $X=2.485 $Y=2.045
c110 33 0 9.89418e-20 $X=3.52 $Y=1.77
c111 32 0 4.077e-19 $X=3.52 $Y=1.77
c112 20 0 8.64737e-20 $X=2.235 $Y=0.88
r113 37 38 8.19535 $w=5.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.485 $Y=2.405
+ $X2=2.485 $Y2=2.775
r114 35 37 6.09114 $w=5.38e-07 $l=2.75e-07 $layer=LI1_cond $X=2.485 $Y=2.13
+ $X2=2.485 $Y2=2.405
r115 35 36 2.23656 $w=4.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=2.13
+ $X2=2.485 $Y2=2.045
r116 33 46 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.77
+ $X2=3.52 $Y2=1.935
r117 33 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.77
+ $X2=3.52 $Y2=1.605
r118 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.52
+ $Y=1.77 $X2=3.52 $Y2=1.77
r119 30 32 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=3.535 $Y=1.96
+ $X2=3.535 $Y2=1.77
r120 29 36 4.86468 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.755 $Y=2.045
+ $X2=2.485 $Y2=2.045
r121 28 30 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.385 $Y=2.045
+ $X2=3.535 $Y2=1.96
r122 28 29 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.385 $Y=2.045
+ $X2=2.755 $Y2=2.045
r123 26 43 31.9995 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.77
+ $X2=2.37 $Y2=1.935
r124 26 42 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.77
+ $X2=2.37 $Y2=1.605
r125 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.77 $X2=2.38 $Y2=1.77
r126 23 36 2.23656 $w=4.35e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.38 $Y=1.96
+ $X2=2.485 $Y2=2.045
r127 23 25 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.38 $Y=1.96
+ $X2=2.38 $Y2=1.77
r128 22 45 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.58 $Y=1.27
+ $X2=3.58 $Y2=1.605
r129 21 22 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=3.61 $Y=1.12
+ $X2=3.61 $Y2=1.27
r130 20 42 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=2.27 $Y=0.88
+ $X2=2.27 $Y2=1.605
r131 19 20 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.235 $Y=0.73
+ $X2=2.235 $Y2=0.88
r132 18 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.64 $Y=0.835
+ $X2=3.64 $Y2=1.12
r133 12 46 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.49 $Y=2.595
+ $X2=3.49 $Y2=1.935
r134 8 43 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.34 $Y=2.595
+ $X2=2.34 $Y2=1.935
r135 3 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.2 $Y=0.445 $X2=2.2
+ $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__HA_LP%A 1 3 8 11 12 13 14 16 21 27 29 31 32 35 37
c97 35 0 1.77619e-19 $X=2.95 $Y=1.615
c98 16 0 7.90742e-20 $X=4.02 $Y=2.595
r99 35 38 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.615
+ $X2=2.95 $Y2=1.78
r100 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.615
+ $X2=2.95 $Y2=1.45
r101 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.615 $X2=2.95 $Y2=1.615
r102 32 36 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.12 $Y=1.615
+ $X2=2.95 $Y2=1.615
r103 30 31 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.035 $Y=1.12
+ $X2=4.035 $Y2=1.27
r104 29 31 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.07 $Y=1.51
+ $X2=4.07 $Y2=1.27
r105 26 27 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=2.86 $Y=0.805
+ $X2=3.135 $Y2=0.805
r106 24 26 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.63 $Y=0.805
+ $X2=2.86 $Y2=0.805
r107 21 30 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4 $Y=0.835 $X2=4
+ $Y2=1.12
r108 18 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4 $Y=0.255 $X2=4
+ $Y2=0.835
r109 14 29 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.02 $Y=1.635
+ $X2=4.02 $Y2=1.51
r110 14 16 238.515 $w=2.5e-07 $l=9.6e-07 $layer=POLY_cond $X=4.02 $Y=1.635
+ $X2=4.02 $Y2=2.595
r111 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.925 $Y=0.18
+ $X2=4 $Y2=0.255
r112 12 13 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=3.925 $Y=0.18
+ $X2=3.21 $Y2=0.18
r113 11 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.135 $Y=0.73
+ $X2=3.135 $Y2=0.805
r114 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.135 $Y=0.255
+ $X2=3.21 $Y2=0.18
r115 10 11 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=3.135 $Y=0.255
+ $X2=3.135 $Y2=0.73
r116 8 38 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.91 $Y=2.595
+ $X2=2.91 $Y2=1.78
r117 4 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.86 $Y=0.88
+ $X2=2.86 $Y2=0.805
r118 4 37 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.86 $Y=0.88
+ $X2=2.86 $Y2=1.45
r119 1 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.63 $Y=0.73
+ $X2=2.63 $Y2=0.805
r120 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.63 $Y=0.73 $X2=2.63
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__HA_LP%SUM 1 2 7 8 9 11 16 17 18 19 20 21 22
r27 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=2.405
+ $X2=0.275 $Y2=2.775
r28 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=2.035
+ $X2=0.275 $Y2=2.405
r29 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=1.665
+ $X2=0.275 $Y2=2.035
r30 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=1.295
+ $X2=0.275 $Y2=1.665
r31 18 36 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.275 $Y=1.295
+ $X2=0.275 $Y2=1.105
r32 17 36 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.275 $Y=0.925
+ $X2=0.275 $Y2=1.105
r33 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=0.555
+ $X2=0.275 $Y2=0.925
r34 13 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.275 $Y=2.865
+ $X2=0.275 $Y2=2.775
r35 9 15 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=2.865 $X2=0.81
+ $Y2=2.95
r36 9 11 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=0.81 $Y=2.865
+ $X2=0.81 $Y2=2.24
r37 8 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.44 $Y=2.95
+ $X2=0.275 $Y2=2.865
r38 7 15 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.645 $Y=2.95
+ $X2=0.81 $Y2=2.95
r39 7 8 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.645 $Y=2.95
+ $X2=0.44 $Y2=2.95
r40 2 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=2.095 $X2=0.81 $Y2=2.95
r41 2 11 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=2.095 $X2=0.81 $Y2=2.24
r42 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.895 $X2=0.275 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__HA_LP%VPWR 1 2 3 12 18 22 27 28 29 31 36 49 50 53 56
r63 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r64 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r65 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r66 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r67 47 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r69 44 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.34 $Y=3.33
+ $X2=3.175 $Y2=3.33
r70 44 46 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.34 $Y=3.33
+ $X2=4.08 $Y2=3.33
r71 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r72 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r73 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 37 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.34 $Y2=3.33
r75 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 36 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.01 $Y=3.33
+ $X2=3.175 $Y2=3.33
r77 36 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.01 $Y=3.33 $X2=2.64
+ $Y2=3.33
r78 34 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r79 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r80 31 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=3.33
+ $X2=1.34 $Y2=3.33
r81 31 33 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=1.175 $Y=3.33 $X2=0.24
+ $Y2=3.33
r82 29 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r83 29 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 29 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r85 27 46 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.38 $Y2=3.33
r87 26 49 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=5.04 $Y2=3.33
r88 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=4.38 $Y2=3.33
r89 22 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.38 $Y=2.24 $X2=4.38
+ $Y2=2.95
r90 20 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=3.245
+ $X2=4.38 $Y2=3.33
r91 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.38 $Y=3.245
+ $X2=4.38 $Y2=2.95
r92 16 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.175 $Y=3.245
+ $X2=3.175 $Y2=3.33
r93 16 18 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.175 $Y=3.245
+ $X2=3.175 $Y2=2.475
r94 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.34 $Y=2.24 $X2=1.34
+ $Y2=2.95
r95 10 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.34 $Y=3.245
+ $X2=1.34 $Y2=3.33
r96 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.34 $Y=3.245
+ $X2=1.34 $Y2=2.95
r97 3 25 400 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=4.145
+ $Y=2.095 $X2=4.38 $Y2=2.95
r98 3 22 400 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=4.145
+ $Y=2.095 $X2=4.38 $Y2=2.24
r99 2 18 300 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=3.035
+ $Y=2.095 $X2=3.175 $Y2=2.475
r100 1 15 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.095 $X2=1.34 $Y2=2.95
r101 1 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.095 $X2=1.34 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__HA_LP%COUT 1 2 7 8 9 10 11 12 13 37 45
r22 38 51 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=4.957 $Y=2.287
+ $X2=4.957 $Y2=2.24
r23 37 49 1.88154 $w=2.43e-07 $l=4e-08 $layer=LI1_cond $X=5.047 $Y=2.035
+ $X2=5.047 $Y2=2.075
r24 23 45 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.005 $Y=0.88
+ $X2=5.005 $Y2=0.925
r25 12 13 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=4.957 $Y=2.405
+ $X2=4.957 $Y2=2.775
r26 12 38 3.19972 $w=4.23e-07 $l=1.18e-07 $layer=LI1_cond $X=4.957 $Y=2.405
+ $X2=4.957 $Y2=2.287
r27 11 51 3.87763 $w=4.23e-07 $l=1.43e-07 $layer=LI1_cond $X=4.957 $Y=2.097
+ $X2=4.957 $Y2=2.24
r28 11 49 2.64642 $w=4.23e-07 $l=2.2e-08 $layer=LI1_cond $X=4.957 $Y=2.097
+ $X2=4.957 $Y2=2.075
r29 11 37 1.08189 $w=2.43e-07 $l=2.3e-08 $layer=LI1_cond $X=5.047 $Y=2.012
+ $X2=5.047 $Y2=2.035
r30 10 11 16.3224 $w=2.43e-07 $l=3.47e-07 $layer=LI1_cond $X=5.047 $Y=1.665
+ $X2=5.047 $Y2=2.012
r31 9 10 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=5.047 $Y=1.295
+ $X2=5.047 $Y2=1.665
r32 9 47 11.7596 $w=2.43e-07 $l=2.5e-07 $layer=LI1_cond $X=5.047 $Y=1.295
+ $X2=5.047 $Y2=1.045
r33 8 47 4.28104 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=5.005 $Y=0.945
+ $X2=5.005 $Y2=1.045
r34 8 45 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=5.005 $Y=0.945
+ $X2=5.005 $Y2=0.925
r35 8 23 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=5.005 $Y=0.825
+ $X2=5.005 $Y2=0.88
r36 7 8 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=5.005 $Y=0.555
+ $X2=5.005 $Y2=0.825
r37 2 51 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.77
+ $Y=2.095 $X2=4.91 $Y2=2.24
r38 1 8 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.625 $X2=5.005 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__HA_LP%VGND 1 2 3 12 16 20 23 24 26 27 28 40 46 47 50
c72 12 0 5.34194e-20 $X=1.065 $Y=1.12
r73 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r74 47 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r75 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r76 44 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.38 $Y=0 $X2=4.215
+ $Y2=0
r77 44 46 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.38 $Y=0 $X2=5.04
+ $Y2=0
r78 40 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=0 $X2=4.215
+ $Y2=0
r79 40 42 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=4.05 $Y=0 $X2=2.64
+ $Y2=0
r80 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r81 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r82 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r83 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r84 32 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r85 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r86 28 51 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r87 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r88 28 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r89 26 38 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.16
+ $Y2=0
r90 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.415
+ $Y2=0
r91 25 42 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.64
+ $Y2=0
r92 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.415
+ $Y2=0
r93 23 31 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=0.72
+ $Y2=0
r94 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=1.025
+ $Y2=0
r95 22 35 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.2
+ $Y2=0
r96 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.025
+ $Y2=0
r97 18 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0
r98 18 20 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0.825
r99 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=0.085
+ $X2=2.415 $Y2=0
r100 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.415 $Y=0.085
+ $X2=2.415 $Y2=0.39
r101 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.025 $Y=0.085
+ $X2=1.025 $Y2=0
r102 10 12 47.7111 $w=2.48e-07 $l=1.035e-06 $layer=LI1_cond $X=1.025 $Y=0.085
+ $X2=1.025 $Y2=1.12
r103 3 20 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.625 $X2=4.215 $Y2=0.825
r104 2 16 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.235 $X2=2.415 $Y2=0.39
r105 1 12 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.925
+ $Y=0.895 $X2=1.065 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LP__HA_LP%A_369_47# 1 2 9 11 12 15
c32 15 0 8.64737e-20 $X=2.845 $Y=0.47
c33 9 0 5.34194e-20 $X=1.985 $Y=0.47
r34 13 15 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=2.885 $Y=0.75
+ $X2=2.885 $Y2=0.47
r35 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.76 $Y=0.835
+ $X2=2.885 $Y2=0.75
r36 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.76 $Y=0.835
+ $X2=2.07 $Y2=0.835
r37 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.945 $Y=0.75
+ $X2=2.07 $Y2=0.835
r38 7 9 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.945 $Y=0.75
+ $X2=1.945 $Y2=0.47
r39 2 15 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.705
+ $Y=0.235 $X2=2.845 $Y2=0.47
r40 1 9 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.235 $X2=1.985 $Y2=0.47
.ends

