* File: sky130_fd_sc_lp__o221a_1.pxi.spice
* Created: Wed Sep  2 10:18:13 2020
* 
x_PM_SKY130_FD_SC_LP__O221A_1%C1 N_C1_M1002_g N_C1_M1003_g N_C1_c_69_n
+ N_C1_c_70_n C1 C1 C1 C1 N_C1_c_72_n C1 PM_SKY130_FD_SC_LP__O221A_1%C1
x_PM_SKY130_FD_SC_LP__O221A_1%B1 N_B1_M1010_g N_B1_M1006_g B1 B1 N_B1_c_111_n
+ N_B1_c_112_n PM_SKY130_FD_SC_LP__O221A_1%B1
x_PM_SKY130_FD_SC_LP__O221A_1%B2 N_B2_M1004_g N_B2_M1000_g B2 N_B2_c_150_n
+ N_B2_c_151_n N_B2_c_152_n PM_SKY130_FD_SC_LP__O221A_1%B2
x_PM_SKY130_FD_SC_LP__O221A_1%A2 N_A2_M1007_g N_A2_M1001_g A2 A2 N_A2_c_188_n
+ N_A2_c_189_n PM_SKY130_FD_SC_LP__O221A_1%A2
x_PM_SKY130_FD_SC_LP__O221A_1%A1 N_A1_M1008_g N_A1_M1011_g A1 N_A1_c_221_n
+ N_A1_c_222_n PM_SKY130_FD_SC_LP__O221A_1%A1
x_PM_SKY130_FD_SC_LP__O221A_1%A_96_49# N_A_96_49#_M1002_s N_A_96_49#_M1003_s
+ N_A_96_49#_M1000_d N_A_96_49#_M1005_g N_A_96_49#_M1009_g N_A_96_49#_c_263_n
+ N_A_96_49#_c_264_n N_A_96_49#_c_252_n N_A_96_49#_c_285_n N_A_96_49#_c_272_n
+ N_A_96_49#_c_294_n N_A_96_49#_c_260_n N_A_96_49#_c_253_n N_A_96_49#_c_254_n
+ N_A_96_49#_c_262_n N_A_96_49#_c_255_n N_A_96_49#_c_256_n N_A_96_49#_c_257_n
+ PM_SKY130_FD_SC_LP__O221A_1%A_96_49#
x_PM_SKY130_FD_SC_LP__O221A_1%VPWR N_VPWR_M1003_d N_VPWR_M1008_d N_VPWR_c_350_n
+ N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n VPWR N_VPWR_c_354_n
+ N_VPWR_c_355_n N_VPWR_c_349_n N_VPWR_c_357_n PM_SKY130_FD_SC_LP__O221A_1%VPWR
x_PM_SKY130_FD_SC_LP__O221A_1%X N_X_M1005_d N_X_M1009_d X X X X X X X X
+ N_X_c_401_n N_X_c_398_n PM_SKY130_FD_SC_LP__O221A_1%X
x_PM_SKY130_FD_SC_LP__O221A_1%A_179_49# N_A_179_49#_M1002_d N_A_179_49#_M1004_d
+ N_A_179_49#_c_423_n N_A_179_49#_c_424_n N_A_179_49#_c_422_n
+ PM_SKY130_FD_SC_LP__O221A_1%A_179_49#
x_PM_SKY130_FD_SC_LP__O221A_1%A_273_49# N_A_273_49#_M1010_d N_A_273_49#_M1007_d
+ N_A_273_49#_c_446_n N_A_273_49#_c_463_p N_A_273_49#_c_447_n
+ PM_SKY130_FD_SC_LP__O221A_1%A_273_49#
x_PM_SKY130_FD_SC_LP__O221A_1%VGND N_VGND_M1007_s N_VGND_M1011_d N_VGND_c_468_n
+ N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n N_VGND_c_473_n
+ VGND N_VGND_c_474_n N_VGND_c_475_n PM_SKY130_FD_SC_LP__O221A_1%VGND
cc_1 VNB N_C1_M1002_g 0.0279212f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=0.665
cc_2 VNB N_C1_c_69_n 0.0416022f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.51
cc_3 VNB N_C1_c_70_n 0.00889595f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.51
cc_4 VNB C1 0.0334075f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_C1_c_72_n 0.0125449f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.51
cc_6 VNB N_B1_M1006_g 0.00579169f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.465
cc_7 VNB B1 0.00286722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_111_n 0.0331104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_112_n 0.0178295f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_10 VNB N_B2_M1000_g 0.0103833f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.465
cc_11 VNB N_B2_c_150_n 0.0316714f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_12 VNB N_B2_c_151_n 0.00385539f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_13 VNB N_B2_c_152_n 0.022105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_M1001_g 0.0108423f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.465
cc_15 VNB A2 0.00942581f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.51
cc_16 VNB N_A2_c_188_n 0.0377127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_189_n 0.0214535f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_18 VNB N_A1_M1008_g 0.00779837f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=0.665
cc_19 VNB A1 0.00347946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_221_n 0.0321476f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_21 VNB N_A1_c_222_n 0.0168033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_96_49#_M1009_g 0.00824724f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_23 VNB N_A_96_49#_c_252_n 0.00321865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_96_49#_c_253_n 0.00176221f $X=-0.19 $Y=-0.245 $X2=0.205 $Y2=1.75
cc_25 VNB N_A_96_49#_c_254_n 0.00433425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_96_49#_c_255_n 0.0036042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_96_49#_c_256_n 0.0375128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_96_49#_c_257_n 0.0201641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_349_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.295
cc_30 VNB X 0.0352475f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.51
cc_31 VNB N_X_c_398_n 0.042066f $X=-0.19 $Y=-0.245 $X2=0.205 $Y2=2.405
cc_32 VNB N_A_179_49#_c_422_n 0.0043955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_273_49#_c_446_n 0.00839969f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.465
cc_34 VNB N_VGND_c_468_n 0.00711065f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.51
cc_35 VNB N_VGND_c_469_n 0.00274151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_470_n 0.0604107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_471_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_472_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_473_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_474_n 0.0233891f $X=-0.19 $Y=-0.245 $X2=0.205 $Y2=1.75
cc_41 VNB N_VGND_c_475_n 0.242449f $X=-0.19 $Y=-0.245 $X2=0.205 $Y2=2.035
cc_42 VPB N_C1_M1003_g 0.0230258f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.465
cc_43 VPB N_C1_c_69_n 0.0150136f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.51
cc_44 VPB N_C1_c_70_n 6.62869e-19 $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.51
cc_45 VPB C1 0.0463462f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_46 VPB N_C1_c_72_n 0.0120169f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.51
cc_47 VPB N_B1_M1006_g 0.0206727f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.465
cc_48 VPB B1 0.00228787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B2_M1000_g 0.0250309f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.465
cc_50 VPB N_A2_M1001_g 0.0237493f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.465
cc_51 VPB N_A1_M1008_g 0.0194425f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=0.665
cc_52 VPB N_A_96_49#_M1009_g 0.025001f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_53 VPB N_A_96_49#_c_252_n 0.00156622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_96_49#_c_260_n 0.0118622f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.295
cc_55 VPB N_A_96_49#_c_253_n 4.12161e-19 $X=-0.19 $Y=1.655 $X2=0.205 $Y2=1.75
cc_56 VPB N_A_96_49#_c_262_n 0.0111851f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.547
cc_57 VPB N_VPWR_c_350_n 0.0055721f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.51
cc_58 VPB N_VPWR_c_351_n 0.00562991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_352_n 0.051873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_353_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_354_n 0.0281856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_355_n 0.0236269f $X=-0.19 $Y=1.655 $X2=0.205 $Y2=1.295
cc_63 VPB N_VPWR_c_349_n 0.0558417f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.295
cc_64 VPB N_VPWR_c_357_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0.205 $Y2=1.75
cc_65 VPB X 0.00201967f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.51
cc_66 VPB X 0.0398164f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_67 VPB N_X_c_401_n 0.0345566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 N_C1_c_70_n N_B1_M1006_g 0.0267714f $X=0.82 $Y=1.51 $X2=0 $Y2=0
cc_69 N_C1_M1002_g B1 3.8043e-19 $X=0.82 $Y=0.665 $X2=0 $Y2=0
cc_70 N_C1_c_70_n B1 7.05823e-19 $X=0.82 $Y=1.51 $X2=0 $Y2=0
cc_71 N_C1_M1002_g N_B1_c_111_n 0.0206051f $X=0.82 $Y=0.665 $X2=0 $Y2=0
cc_72 N_C1_M1002_g N_B1_c_112_n 0.0148812f $X=0.82 $Y=0.665 $X2=0 $Y2=0
cc_73 C1 N_A_96_49#_c_263_n 0.0194487f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_74 N_C1_M1003_g N_A_96_49#_c_264_n 0.0113245f $X=0.82 $Y=2.465 $X2=0 $Y2=0
cc_75 C1 N_A_96_49#_c_264_n 0.0372284f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_76 N_C1_M1002_g N_A_96_49#_c_252_n 0.00505411f $X=0.82 $Y=0.665 $X2=0 $Y2=0
cc_77 N_C1_M1003_g N_A_96_49#_c_252_n 0.00782041f $X=0.82 $Y=2.465 $X2=0 $Y2=0
cc_78 N_C1_c_70_n N_A_96_49#_c_252_n 0.0102553f $X=0.82 $Y=1.51 $X2=0 $Y2=0
cc_79 C1 N_A_96_49#_c_252_n 0.00614565f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 C1 N_A_96_49#_c_252_n 0.00652378f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_81 N_C1_c_72_n N_A_96_49#_c_252_n 0.0264609f $X=0.42 $Y=1.51 $X2=0 $Y2=0
cc_82 N_C1_M1003_g N_A_96_49#_c_272_n 0.0124366f $X=0.82 $Y=2.465 $X2=0 $Y2=0
cc_83 N_C1_c_69_n N_A_96_49#_c_272_n 0.00565431f $X=0.745 $Y=1.51 $X2=0 $Y2=0
cc_84 C1 N_A_96_49#_c_272_n 0.0142331f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_85 N_C1_c_72_n N_A_96_49#_c_272_n 0.00532375f $X=0.42 $Y=1.51 $X2=0 $Y2=0
cc_86 N_C1_M1002_g N_A_96_49#_c_254_n 0.0128526f $X=0.82 $Y=0.665 $X2=0 $Y2=0
cc_87 N_C1_c_69_n N_A_96_49#_c_254_n 0.00831114f $X=0.745 $Y=1.51 $X2=0 $Y2=0
cc_88 C1 N_A_96_49#_c_254_n 0.0139059f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_C1_c_72_n N_A_96_49#_c_254_n 0.00534458f $X=0.42 $Y=1.51 $X2=0 $Y2=0
cc_90 N_C1_M1003_g N_VPWR_c_350_n 0.00430884f $X=0.82 $Y=2.465 $X2=0 $Y2=0
cc_91 N_C1_M1003_g N_VPWR_c_354_n 0.00571722f $X=0.82 $Y=2.465 $X2=0 $Y2=0
cc_92 C1 N_VPWR_c_354_n 0.00382558f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_93 N_C1_M1003_g N_VPWR_c_349_n 0.0118478f $X=0.82 $Y=2.465 $X2=0 $Y2=0
cc_94 C1 N_VPWR_c_349_n 0.00660791f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_95 N_C1_M1002_g N_VGND_c_470_n 0.00575161f $X=0.82 $Y=0.665 $X2=0 $Y2=0
cc_96 C1 N_VGND_c_470_n 0.003781f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_97 N_C1_M1002_g N_VGND_c_475_n 0.0121974f $X=0.82 $Y=0.665 $X2=0 $Y2=0
cc_98 C1 N_VGND_c_475_n 0.00656137f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_99 B1 N_B2_M1000_g 0.00115588f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B1_c_111_n N_B2_M1000_g 0.0878918f $X=1.27 $Y=1.375 $X2=0 $Y2=0
cc_101 B1 N_B2_c_150_n 3.0992e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B1_c_111_n N_B2_c_150_n 0.0195963f $X=1.27 $Y=1.375 $X2=0 $Y2=0
cc_103 B1 N_B2_c_151_n 0.0236906f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B1_c_111_n N_B2_c_151_n 0.00197091f $X=1.27 $Y=1.375 $X2=0 $Y2=0
cc_105 N_B1_c_112_n N_B2_c_152_n 0.0325106f $X=1.27 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B1_M1006_g N_A_96_49#_c_264_n 7.25409e-19 $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_107 N_B1_M1006_g N_A_96_49#_c_252_n 0.00225476f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_108 B1 N_A_96_49#_c_252_n 0.0409256f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B1_c_111_n N_A_96_49#_c_252_n 0.00174016f $X=1.27 $Y=1.375 $X2=0 $Y2=0
cc_110 N_B1_c_112_n N_A_96_49#_c_252_n 5.05433e-19 $X=1.27 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B1_M1006_g N_A_96_49#_c_285_n 0.0168914f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_112 B1 N_A_96_49#_c_285_n 0.019074f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B1_c_111_n N_A_96_49#_c_285_n 6.82098e-19 $X=1.27 $Y=1.375 $X2=0 $Y2=0
cc_114 N_B1_c_112_n N_A_96_49#_c_254_n 0.00220526f $X=1.27 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B1_M1006_g N_A_96_49#_c_262_n 0.00427063f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_116 B1 N_A_96_49#_c_262_n 0.0021011f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B1_M1006_g N_VPWR_c_350_n 0.00430884f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_118 N_B1_M1006_g N_VPWR_c_352_n 0.00585385f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B1_M1006_g N_VPWR_c_349_n 0.0108711f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B1_c_112_n N_A_179_49#_c_423_n 0.0111297f $X=1.27 $Y=1.21 $X2=0 $Y2=0
cc_121 B1 N_A_179_49#_c_424_n 0.00420396f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B1_c_111_n N_A_179_49#_c_424_n 5.24871e-19 $X=1.27 $Y=1.375 $X2=0 $Y2=0
cc_123 N_B1_c_112_n N_A_179_49#_c_424_n 0.00574327f $X=1.27 $Y=1.21 $X2=0 $Y2=0
cc_124 N_B1_c_112_n N_A_179_49#_c_422_n 5.41816e-19 $X=1.27 $Y=1.21 $X2=0 $Y2=0
cc_125 N_B1_c_111_n N_A_273_49#_c_447_n 0.00107139f $X=1.27 $Y=1.375 $X2=0 $Y2=0
cc_126 N_B1_c_112_n N_VGND_c_470_n 0.00351205f $X=1.27 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B1_c_112_n N_VGND_c_475_n 0.00544735f $X=1.27 $Y=1.21 $X2=0 $Y2=0
cc_128 N_B2_c_150_n N_A2_M1001_g 2.15658e-19 $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_129 N_B2_c_150_n A2 0.00284984f $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_130 N_B2_c_151_n A2 0.0270658f $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_131 N_B2_c_152_n A2 2.28883e-19 $X=1.815 $Y=1.195 $X2=0 $Y2=0
cc_132 N_B2_c_150_n N_A2_c_188_n 0.0113937f $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_133 N_B2_c_151_n N_A2_c_188_n 2.51591e-19 $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_134 N_B2_c_151_n N_A_96_49#_c_252_n 4.42644e-19 $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_135 N_B2_M1000_g N_A_96_49#_c_285_n 0.0125009f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_136 N_B2_c_151_n N_A_96_49#_c_285_n 0.00783741f $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_137 N_B2_M1000_g N_A_96_49#_c_294_n 0.0211209f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_138 N_B2_M1000_g N_A_96_49#_c_262_n 0.0088708f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_139 N_B2_c_150_n N_A_96_49#_c_262_n 0.00541895f $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_140 N_B2_c_151_n N_A_96_49#_c_262_n 0.00866246f $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_141 N_B2_M1000_g N_VPWR_c_352_n 0.0054895f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_142 N_B2_M1000_g N_VPWR_c_349_n 0.0112391f $X=1.75 $Y=2.465 $X2=0 $Y2=0
cc_143 N_B2_c_152_n N_A_179_49#_c_423_n 0.00832638f $X=1.815 $Y=1.195 $X2=0
+ $Y2=0
cc_144 N_B2_c_152_n N_A_179_49#_c_424_n 4.94307e-19 $X=1.815 $Y=1.195 $X2=0
+ $Y2=0
cc_145 N_B2_c_152_n N_A_179_49#_c_422_n 0.00723256f $X=1.815 $Y=1.195 $X2=0
+ $Y2=0
cc_146 N_B2_c_150_n N_A_273_49#_c_446_n 0.00541116f $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_147 N_B2_c_151_n N_A_273_49#_c_446_n 0.0178187f $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_148 N_B2_c_152_n N_A_273_49#_c_446_n 0.0118728f $X=1.815 $Y=1.195 $X2=0 $Y2=0
cc_149 N_B2_c_151_n N_A_273_49#_c_447_n 0.0022859f $X=1.82 $Y=1.36 $X2=0 $Y2=0
cc_150 N_B2_c_152_n N_VGND_c_468_n 0.00322437f $X=1.815 $Y=1.195 $X2=0 $Y2=0
cc_151 N_B2_c_152_n N_VGND_c_470_n 0.00352686f $X=1.815 $Y=1.195 $X2=0 $Y2=0
cc_152 N_B2_c_152_n N_VGND_c_475_n 0.00662799f $X=1.815 $Y=1.195 $X2=0 $Y2=0
cc_153 N_A2_M1001_g N_A1_M1008_g 0.061607f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_154 A2 A1 0.0262026f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_155 N_A2_c_188_n A1 3.86187e-19 $X=2.515 $Y=1.35 $X2=0 $Y2=0
cc_156 A2 N_A1_c_221_n 0.00201873f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A2_c_188_n N_A1_c_221_n 0.061607f $X=2.515 $Y=1.35 $X2=0 $Y2=0
cc_158 N_A2_c_189_n N_A1_c_222_n 0.0151583f $X=2.525 $Y=1.185 $X2=0 $Y2=0
cc_159 N_A2_M1001_g N_A_96_49#_c_294_n 0.020896f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A2_M1001_g N_A_96_49#_c_260_n 0.0105613f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_161 A2 N_A_96_49#_c_260_n 0.0101292f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_162 N_A2_M1001_g N_A_96_49#_c_262_n 0.00934167f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_163 A2 N_A_96_49#_c_262_n 0.045556f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A2_c_188_n N_A_96_49#_c_262_n 0.00672244f $X=2.515 $Y=1.35 $X2=0 $Y2=0
cc_165 N_A2_M1001_g N_VPWR_c_352_n 0.00533769f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A2_M1001_g N_VPWR_c_349_n 0.0107818f $X=2.67 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A2_c_189_n N_A_179_49#_c_422_n 8.87696e-19 $X=2.525 $Y=1.185 $X2=0
+ $Y2=0
cc_168 A2 N_A_273_49#_c_446_n 0.0495386f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_169 N_A2_c_188_n N_A_273_49#_c_446_n 0.00637691f $X=2.515 $Y=1.35 $X2=0 $Y2=0
cc_170 N_A2_c_189_n N_A_273_49#_c_446_n 0.0117904f $X=2.525 $Y=1.185 $X2=0 $Y2=0
cc_171 N_A2_c_189_n N_VGND_c_468_n 0.0120778f $X=2.525 $Y=1.185 $X2=0 $Y2=0
cc_172 N_A2_c_189_n N_VGND_c_469_n 6.17119e-19 $X=2.525 $Y=1.185 $X2=0 $Y2=0
cc_173 N_A2_c_189_n N_VGND_c_472_n 0.00486043f $X=2.525 $Y=1.185 $X2=0 $Y2=0
cc_174 N_A2_c_189_n N_VGND_c_475_n 0.0045769f $X=2.525 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A1_M1008_g N_A_96_49#_M1009_g 0.0374704f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A1_M1008_g N_A_96_49#_c_260_n 0.015282f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_177 A1 N_A_96_49#_c_260_n 0.0188208f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A1_c_221_n N_A_96_49#_c_260_n 0.00308907f $X=3.12 $Y=1.35 $X2=0 $Y2=0
cc_179 N_A1_M1008_g N_A_96_49#_c_253_n 0.00341786f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A1_M1008_g N_A_96_49#_c_262_n 0.00389301f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_181 A1 N_A_96_49#_c_255_n 0.0258899f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A1_c_221_n N_A_96_49#_c_255_n 0.00210535f $X=3.12 $Y=1.35 $X2=0 $Y2=0
cc_183 A1 N_A_96_49#_c_256_n 3.04982e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A1_c_221_n N_A_96_49#_c_256_n 0.0205073f $X=3.12 $Y=1.35 $X2=0 $Y2=0
cc_185 N_A1_c_222_n N_A_96_49#_c_257_n 0.0142021f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_186 N_A1_M1008_g N_VPWR_c_351_n 0.00986228f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A1_M1008_g N_VPWR_c_352_n 0.00585385f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A1_M1008_g N_VPWR_c_349_n 0.0109986f $X=3.03 $Y=2.465 $X2=0 $Y2=0
cc_189 A1 N_A_273_49#_c_446_n 0.00145093f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A1_c_222_n N_VGND_c_468_n 5.68743e-19 $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_191 A1 N_VGND_c_469_n 0.00374133f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A1_c_221_n N_VGND_c_469_n 0.00251738f $X=3.12 $Y=1.35 $X2=0 $Y2=0
cc_193 N_A1_c_222_n N_VGND_c_469_n 0.0128188f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_194 N_A1_c_222_n N_VGND_c_472_n 0.00486043f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_195 N_A1_c_222_n N_VGND_c_475_n 0.0082726f $X=3.12 $Y=1.185 $X2=0 $Y2=0
cc_196 N_A_96_49#_c_285_n N_VPWR_M1003_d 0.0102231f $X=1.8 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_197 N_A_96_49#_c_260_n N_VPWR_M1008_d 0.00336218f $X=3.395 $Y=1.78 $X2=0
+ $Y2=0
cc_198 N_A_96_49#_c_285_n N_VPWR_c_350_n 0.022455f $X=1.8 $Y=2.015 $X2=0 $Y2=0
cc_199 N_A_96_49#_M1009_g N_VPWR_c_351_n 0.0133011f $X=3.605 $Y=2.465 $X2=0
+ $Y2=0
cc_200 N_A_96_49#_c_260_n N_VPWR_c_351_n 0.0252833f $X=3.395 $Y=1.78 $X2=0 $Y2=0
cc_201 N_A_96_49#_c_294_n N_VPWR_c_352_n 0.0540585f $X=1.965 $Y=2.91 $X2=0 $Y2=0
cc_202 N_A_96_49#_c_264_n N_VPWR_c_354_n 0.0161033f $X=0.605 $Y=2.91 $X2=0 $Y2=0
cc_203 N_A_96_49#_M1009_g N_VPWR_c_355_n 0.0054895f $X=3.605 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_A_96_49#_M1003_s N_VPWR_c_349_n 0.00270818f $X=0.48 $Y=1.835 $X2=0
+ $Y2=0
cc_205 N_A_96_49#_M1000_d N_VPWR_c_349_n 0.00631386f $X=1.825 $Y=1.835 $X2=0
+ $Y2=0
cc_206 N_A_96_49#_M1009_g N_VPWR_c_349_n 0.0113689f $X=3.605 $Y=2.465 $X2=0
+ $Y2=0
cc_207 N_A_96_49#_c_264_n N_VPWR_c_349_n 0.00991608f $X=0.605 $Y=2.91 $X2=0
+ $Y2=0
cc_208 N_A_96_49#_c_294_n N_VPWR_c_349_n 0.031779f $X=1.965 $Y=2.91 $X2=0 $Y2=0
cc_209 N_A_96_49#_c_285_n A_287_367# 0.00844885f $X=1.8 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_210 N_A_96_49#_c_260_n A_549_367# 0.00366293f $X=3.395 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_211 N_A_96_49#_M1009_g X 0.00256752f $X=3.605 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A_96_49#_c_253_n X 0.00557919f $X=3.48 $Y=1.695 $X2=0 $Y2=0
cc_213 N_A_96_49#_c_255_n X 0.0261167f $X=3.67 $Y=1.35 $X2=0 $Y2=0
cc_214 N_A_96_49#_c_256_n X 0.00919167f $X=3.67 $Y=1.35 $X2=0 $Y2=0
cc_215 N_A_96_49#_c_257_n X 0.00391134f $X=3.692 $Y=1.185 $X2=0 $Y2=0
cc_216 N_A_96_49#_M1009_g X 0.0102622f $X=3.605 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_96_49#_M1009_g N_X_c_401_n 0.00853422f $X=3.605 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A_96_49#_c_260_n N_X_c_401_n 0.0134088f $X=3.395 $Y=1.78 $X2=0 $Y2=0
cc_219 N_A_96_49#_c_255_n N_X_c_401_n 0.00325289f $X=3.67 $Y=1.35 $X2=0 $Y2=0
cc_220 N_A_96_49#_c_256_n N_X_c_401_n 0.00449728f $X=3.67 $Y=1.35 $X2=0 $Y2=0
cc_221 N_A_96_49#_c_255_n N_X_c_398_n 0.0062995f $X=3.67 $Y=1.35 $X2=0 $Y2=0
cc_222 N_A_96_49#_c_256_n N_X_c_398_n 0.00646912f $X=3.67 $Y=1.35 $X2=0 $Y2=0
cc_223 N_A_96_49#_c_255_n N_VGND_c_469_n 0.00544187f $X=3.67 $Y=1.35 $X2=0 $Y2=0
cc_224 N_A_96_49#_c_257_n N_VGND_c_469_n 0.00361923f $X=3.692 $Y=1.185 $X2=0
+ $Y2=0
cc_225 N_A_96_49#_c_263_n N_VGND_c_470_n 0.0149547f $X=0.605 $Y=0.42 $X2=0 $Y2=0
cc_226 N_A_96_49#_c_257_n N_VGND_c_474_n 0.00585385f $X=3.692 $Y=1.185 $X2=0
+ $Y2=0
cc_227 N_A_96_49#_M1002_s N_VGND_c_475_n 0.00320142f $X=0.48 $Y=0.245 $X2=0
+ $Y2=0
cc_228 N_A_96_49#_c_263_n N_VGND_c_475_n 0.0090585f $X=0.605 $Y=0.42 $X2=0 $Y2=0
cc_229 N_A_96_49#_c_257_n N_VGND_c_475_n 0.0117644f $X=3.692 $Y=1.185 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_349_n A_287_367# 0.010279f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_231 N_VPWR_c_349_n A_549_367# 0.00899413f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_232 N_VPWR_c_349_n N_X_M1009_d 0.00231914f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_233 N_VPWR_c_351_n X 0.057631f $X=3.305 $Y=2.12 $X2=0 $Y2=0
cc_234 N_VPWR_c_355_n X 0.0389409f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_235 N_VPWR_c_349_n X 0.0222777f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_236 N_VPWR_c_351_n N_X_c_401_n 0.0213412f $X=3.305 $Y=2.12 $X2=0 $Y2=0
cc_237 N_X_c_398_n N_VGND_c_474_n 0.0396611f $X=3.785 $Y=0.42 $X2=0 $Y2=0
cc_238 N_X_M1005_d N_VGND_c_475_n 0.00232552f $X=3.645 $Y=0.235 $X2=0 $Y2=0
cc_239 N_X_c_398_n N_VGND_c_475_n 0.0226657f $X=3.785 $Y=0.42 $X2=0 $Y2=0
cc_240 N_A_179_49#_c_423_n N_A_273_49#_M1010_d 0.00332344f $X=1.77 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_241 N_A_179_49#_M1004_d N_A_273_49#_c_446_n 0.00722294f $X=1.795 $Y=0.245
+ $X2=0 $Y2=0
cc_242 N_A_179_49#_c_423_n N_A_273_49#_c_446_n 0.00347435f $X=1.77 $Y=0.34 $X2=0
+ $Y2=0
cc_243 N_A_179_49#_c_422_n N_A_273_49#_c_446_n 0.0206895f $X=1.935 $Y=0.34 $X2=0
+ $Y2=0
cc_244 N_A_179_49#_c_423_n N_A_273_49#_c_447_n 0.012181f $X=1.77 $Y=0.34 $X2=0
+ $Y2=0
cc_245 N_A_179_49#_c_422_n N_VGND_c_468_n 0.032341f $X=1.935 $Y=0.34 $X2=0 $Y2=0
cc_246 N_A_179_49#_c_423_n N_VGND_c_470_n 0.0305087f $X=1.77 $Y=0.34 $X2=0 $Y2=0
cc_247 N_A_179_49#_c_424_n N_VGND_c_470_n 0.0191643f $X=1.065 $Y=0.39 $X2=0
+ $Y2=0
cc_248 N_A_179_49#_c_422_n N_VGND_c_470_n 0.0204255f $X=1.935 $Y=0.34 $X2=0
+ $Y2=0
cc_249 N_A_179_49#_M1002_d N_VGND_c_475_n 0.00252509f $X=0.895 $Y=0.245 $X2=0
+ $Y2=0
cc_250 N_A_179_49#_M1004_d N_VGND_c_475_n 0.00213105f $X=1.795 $Y=0.245 $X2=0
+ $Y2=0
cc_251 N_A_179_49#_c_423_n N_VGND_c_475_n 0.0191162f $X=1.77 $Y=0.34 $X2=0 $Y2=0
cc_252 N_A_179_49#_c_424_n N_VGND_c_475_n 0.0126354f $X=1.065 $Y=0.39 $X2=0
+ $Y2=0
cc_253 N_A_179_49#_c_422_n N_VGND_c_475_n 0.0124872f $X=1.935 $Y=0.34 $X2=0
+ $Y2=0
cc_254 N_A_273_49#_c_446_n N_VGND_M1007_s 0.00467546f $X=2.79 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_255 N_A_273_49#_c_446_n N_VGND_c_468_n 0.021529f $X=2.79 $Y=0.93 $X2=0 $Y2=0
cc_256 N_A_273_49#_c_463_p N_VGND_c_472_n 0.0124525f $X=2.885 $Y=0.42 $X2=0
+ $Y2=0
cc_257 N_A_273_49#_M1010_d N_VGND_c_475_n 0.00224381f $X=1.365 $Y=0.245 $X2=0
+ $Y2=0
cc_258 N_A_273_49#_M1007_d N_VGND_c_475_n 0.00408812f $X=2.745 $Y=0.235 $X2=0
+ $Y2=0
cc_259 N_A_273_49#_c_446_n N_VGND_c_475_n 0.0134765f $X=2.79 $Y=0.93 $X2=0 $Y2=0
cc_260 N_A_273_49#_c_463_p N_VGND_c_475_n 0.00730901f $X=2.885 $Y=0.42 $X2=0
+ $Y2=0
