# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065000 1.450000 2.345000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.564900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.605000 0.260000 8.075000 1.060000 ;
        RECT 7.620000 1.740000 8.075000 3.075000 ;
        RECT 7.815000 1.060000 8.075000 1.740000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.750000 0.260000 7.055000 2.155000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945000 1.210000 5.470000 2.120000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.995000 0.885000 1.755000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.205000  0.510000 0.535000 0.825000 ;
      RECT 0.205000  0.825000 0.455000 1.925000 ;
      RECT 0.205000  1.925000 1.205000 2.255000 ;
      RECT 0.205000  2.255000 0.500000 3.075000 ;
      RECT 0.670000  2.425000 0.895000 3.245000 ;
      RECT 0.715000  0.085000 1.045000 0.825000 ;
      RECT 1.065000  2.425000 1.545000 2.905000 ;
      RECT 1.065000  2.905000 2.425000 3.075000 ;
      RECT 1.220000  0.510000 1.550000 0.840000 ;
      RECT 1.375000  0.840000 1.545000 2.425000 ;
      RECT 1.725000  1.085000 2.180000 1.110000 ;
      RECT 1.725000  1.110000 2.840000 1.280000 ;
      RECT 1.725000  1.280000 1.895000 2.385000 ;
      RECT 1.725000  2.385000 2.085000 2.735000 ;
      RECT 1.885000  0.640000 2.180000 1.085000 ;
      RECT 2.255000  2.290000 3.195000 2.460000 ;
      RECT 2.255000  2.460000 2.425000 2.905000 ;
      RECT 2.350000  0.085000 2.645000 0.940000 ;
      RECT 2.590000  1.280000 2.840000 2.025000 ;
      RECT 2.595000  2.630000 2.855000 3.245000 ;
      RECT 3.025000  1.125000 3.245000 1.455000 ;
      RECT 3.025000  1.455000 3.195000 2.290000 ;
      RECT 3.025000  2.460000 3.195000 2.905000 ;
      RECT 3.025000  2.905000 4.015000 3.075000 ;
      RECT 3.160000  0.635000 3.585000 0.955000 ;
      RECT 3.365000  2.385000 3.585000 2.735000 ;
      RECT 3.415000  0.955000 3.585000 0.995000 ;
      RECT 3.415000  0.995000 4.775000 1.165000 ;
      RECT 3.415000  1.165000 3.585000 2.385000 ;
      RECT 3.755000  2.135000 4.015000 2.905000 ;
      RECT 3.985000  1.335000 4.355000 1.925000 ;
      RECT 4.005000  0.085000 4.335000 0.825000 ;
      RECT 4.185000  1.925000 4.355000 2.300000 ;
      RECT 4.185000  2.300000 5.810000 2.325000 ;
      RECT 4.185000  2.325000 7.450000 2.470000 ;
      RECT 4.525000  1.165000 4.775000 1.515000 ;
      RECT 4.525000  2.640000 4.825000 3.245000 ;
      RECT 4.545000  0.255000 4.875000 0.655000 ;
      RECT 4.545000  0.655000 5.810000 0.825000 ;
      RECT 4.995000  2.470000 7.450000 2.495000 ;
      RECT 4.995000  2.495000 5.215000 3.060000 ;
      RECT 5.335000  0.085000 5.665000 0.485000 ;
      RECT 5.385000  2.665000 5.715000 3.245000 ;
      RECT 5.640000  0.825000 5.810000 1.295000 ;
      RECT 5.640000  1.295000 6.030000 1.625000 ;
      RECT 5.640000  1.625000 5.810000 2.300000 ;
      RECT 5.980000  0.705000 6.580000 1.035000 ;
      RECT 5.990000  1.805000 6.380000 2.135000 ;
      RECT 6.210000  1.035000 6.580000 1.435000 ;
      RECT 6.210000  1.435000 6.380000 1.805000 ;
      RECT 7.120000  2.665000 7.450000 3.245000 ;
      RECT 7.225000  0.085000 7.435000 1.060000 ;
      RECT 7.225000  1.230000 7.645000 1.560000 ;
      RECT 7.225000  1.560000 7.450000 2.325000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrbp_1
