* File: sky130_fd_sc_lp__and4b_m.spice
* Created: Fri Aug 28 10:08:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4b_m.pex.spice"
.subckt sky130_fd_sc_lp__and4b_m  VNB VPB A_N B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_N_M1007_g N_A_27_55#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_323_73# N_A_27_55#_M1002_g N_A_240_73#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1003 A_395_73# N_B_M1003_g A_323_73# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1004 A_467_73# N_C_M1004_g A_395_73# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75000.9 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_D_M1009_g A_467_73# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0819 PD=0.81 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75001.4 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1011 N_X_M1011_d N_A_240_73#_M1011_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=31.428 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_N_M1008_g N_A_27_55#_M1008_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0651 AS=0.1113 PD=0.73 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1010 N_A_240_73#_M1010_d N_A_27_55#_M1010_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0609 AS=0.0651 PD=0.71 PS=0.73 NRD=0 NRS=14.0658 M=1 R=2.8
+ SA=75000.6 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_A_240_73#_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06195 AS=0.0609 PD=0.715 PS=0.71 NRD=4.6886 NRS=4.6886 M=1 R=2.8
+ SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_240_73#_M1005_d N_C_M1005_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06405 AS=0.06195 PD=0.725 PS=0.715 NRD=11.7215 NRS=2.3443 M=1 R=2.8
+ SA=75001.5 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_D_M1006_g N_A_240_73#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.06405 PD=0.81 PS=0.725 NRD=37.5088 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_240_73#_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=14.0658 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__and4b_m.pxi.spice"
*
.ends
*
*
