* File: sky130_fd_sc_lp__ebufn_lp.spice
* Created: Fri Aug 28 10:32:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ebufn_lp.pex.spice"
.subckt sky130_fd_sc_lp__ebufn_lp  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 A_122_131# N_A_M1004_g N_A_29_483#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g A_122_131# VNB NSHORT L=0.15 W=0.42 AD=0.1015
+ AS=0.0441 PD=0.84 PS=0.63 NRD=34.284 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1009 A_308_47# N_A_242_237#_M1009_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.203 PD=1.08 PS=1.68 NRD=9.276 NRS=2.856 M=1 R=5.6 SA=75000.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_Z_M1008_d N_A_29_483#_M1008_g A_308_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1008 PD=2.25 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 A_708_47# N_TE_B_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_242_237#_M1003_d N_TE_B_M1003_g A_708_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 A_116_483# N_A_M1010_g N_A_29_483#_M1010_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g A_116_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.4384
+ AS=0.0768 PD=2.65 PS=0.88 NRD=123.125 NRS=19.9955 M=1 R=4.26667 SA=75000.6
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 A_515_367# N_A_29_483#_M1002_g N_Z_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.3591 PD=1.5 PS=3.09 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_TE_B_M1007_g A_515_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.284826 AS=0.1512 PD=2.19505 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75000.6
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1011 A_702_401# N_TE_B_M1011_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.144674 PD=0.88 PS=1.11495 NRD=19.9955 NRS=36.1495 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_242_237#_M1006_d N_TE_B_M1006_g A_702_401# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__ebufn_lp.pxi.spice"
*
.ends
*
*
