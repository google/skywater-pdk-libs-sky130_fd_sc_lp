* File: sky130_fd_sc_lp__a32oi_lp.spice
* Created: Wed Sep  2 09:28:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32oi_lp.pex.spice"
.subckt sky130_fd_sc_lp__a32oi_lp  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1008 A_140_47# N_B2_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g A_140_47# VNB NSHORT L=0.15 W=0.42 AD=0.11445
+ AS=0.0504 PD=0.965 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1001 A_357_47# N_A1_M1001_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.11445 PD=0.81 PS=0.965 NRD=39.996 NRS=75.708 M=1 R=2.8 SA=75001.3
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 A_465_47# N_A2_M1004_g A_357_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=39.996 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A3_M1003_g A_465_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.2 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g N_A_56_409#_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1000 N_A_56_409#_M1000_d N_B1_M1000_g N_Y_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_56_409#_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1002 N_A_56_409#_M1002_d N_A2_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A3_M1009_g N_A_56_409#_M1002_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a32oi_lp.pxi.spice"
*
.ends
*
*
