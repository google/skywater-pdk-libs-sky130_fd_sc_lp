* File: sky130_fd_sc_lp__o32a_m.pex.spice
* Created: Fri Aug 28 11:17:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32A_M%A1 2 5 8 10 11 12 13 18 20
c35 10 0 1.83051e-19 $X=1.057 $Y=1.605
r36 18 20 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.057 $Y=1.1
+ $X2=1.057 $Y2=0.935
r37 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.035
+ $Y=1.1 $X2=1.035 $Y2=1.1
r38 12 13 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.877 $Y=1.295
+ $X2=0.877 $Y2=1.665
r39 12 19 4.80898 $w=4.83e-07 $l=1.95e-07 $layer=LI1_cond $X=0.877 $Y=1.295
+ $X2=0.877 $Y2=1.1
r40 11 19 4.31575 $w=4.83e-07 $l=1.75e-07 $layer=LI1_cond $X=0.877 $Y=0.925
+ $X2=0.877 $Y2=1.1
r41 8 10 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.17 $Y=2.225
+ $X2=1.17 $Y2=1.605
r42 5 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.17 $Y=0.615
+ $X2=1.17 $Y2=0.935
r43 2 10 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=1.057 $Y=1.418
+ $X2=1.057 $Y2=1.605
r44 1 18 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=1.057 $Y=1.122
+ $X2=1.057 $Y2=1.1
r45 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=1.057 $Y=1.122
+ $X2=1.057 $Y2=1.418
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_M%A2 3 7 11 12 13 14 15 16 22
r40 15 16 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=2.035
+ $X2=1.65 $Y2=2.405
r41 14 15 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=2.035
r42 13 14 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=1.295
+ $X2=1.65 $Y2=1.665
r43 13 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.62
+ $Y=1.35 $X2=1.62 $Y2=1.35
r44 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.62 $Y=1.69
+ $X2=1.62 $Y2=1.35
r45 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.69
+ $X2=1.62 $Y2=1.855
r46 10 22 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.185
+ $X2=1.62 $Y2=1.35
r47 7 10 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.6 $Y=0.615 $X2=1.6
+ $Y2=1.185
r48 3 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.53 $Y=2.225
+ $X2=1.53 $Y2=1.855
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_M%A_86_55# 1 2 9 12 13 14 15 18 20 23 24 27 30
c71 30 0 1.93692e-19 $X=2.895 $Y=0.7
c72 15 0 1.30319e-19 $X=2.425 $Y=2.94
c73 13 0 1.67781e-19 $X=2.11 $Y=3.03
r74 26 30 8.98746 $w=3.19e-07 $l=3.17884e-07 $layer=LI1_cond $X=3.13 $Y=1.005
+ $X2=2.895 $Y2=0.81
r75 26 27 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.13 $Y=1.005
+ $X2=3.13 $Y2=1.875
r76 25 28 1.09592 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.635 $Y=1.96
+ $X2=2.53 $Y2=1.96
r77 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.045 $Y=1.96
+ $X2=3.13 $Y2=1.875
r78 24 25 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.045 $Y=1.96
+ $X2=2.635 $Y2=1.96
r79 21 23 29.8398 $w=2.08e-07 $l=5.65e-07 $layer=LI1_cond $X=2.53 $Y=2.855
+ $X2=2.53 $Y2=2.29
r80 20 28 15.9521 $w=2.1e-07 $l=2.7e-07 $layer=LI1_cond $X=2.53 $Y=2.23 $X2=2.53
+ $Y2=1.96
r81 20 23 3.16883 $w=2.08e-07 $l=6e-08 $layer=LI1_cond $X=2.53 $Y=2.23 $X2=2.53
+ $Y2=2.29
r82 18 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.275 $Y=2.94
+ $X2=2.275 $Y2=3.03
r83 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.275
+ $Y=2.94 $X2=2.275 $Y2=2.94
r84 15 21 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.425 $Y=2.94
+ $X2=2.53 $Y2=2.855
r85 15 17 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.425 $Y=2.94
+ $X2=2.275 $Y2=2.94
r86 13 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=3.03
+ $X2=2.275 $Y2=3.03
r87 13 14 784.532 $w=1.5e-07 $l=1.53e-06 $layer=POLY_cond $X=2.11 $Y=3.03
+ $X2=0.58 $Y2=3.03
r88 9 12 825.553 $w=1.5e-07 $l=1.61e-06 $layer=POLY_cond $X=0.505 $Y=0.615
+ $X2=0.505 $Y2=2.225
r89 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.505 $Y=2.955
+ $X2=0.58 $Y2=3.03
r90 7 12 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.505 $Y=2.955
+ $X2=0.505 $Y2=2.225
r91 2 23 600 $w=1.7e-07 $l=5.04083e-07 $layer=licon1_PDIFF $count=1 $X=2.145
+ $Y=2.015 $X2=2.53 $Y2=2.29
r92 1 30 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.405 $X2=2.895 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_M%A3 3 7 11 12 13 14 15 16 22
c47 13 0 1.67781e-19 $X=2.16 $Y=1.295
c48 7 0 1.93692e-19 $X=2.25 $Y=0.615
c49 3 0 1.30319e-19 $X=2.07 $Y=2.225
r50 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.405
r51 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=2.035
r52 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.665
r53 13 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.16
+ $Y=1.35 $X2=2.16 $Y2=1.35
r54 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.16 $Y=1.69
+ $X2=2.16 $Y2=1.35
r55 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.69
+ $X2=2.16 $Y2=1.855
r56 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.185
+ $X2=2.16 $Y2=1.35
r57 7 10 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.25 $Y=0.615
+ $X2=2.25 $Y2=1.185
r58 3 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.07 $Y=2.225
+ $X2=2.07 $Y2=1.855
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_M%B2 3 7 11 12 13 16
c43 3 0 3.22814e-20 $X=2.68 $Y=0.615
r44 13 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.7 $Y=1.27
+ $X2=2.7 $Y2=1.27
r45 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.7 $Y=1.61 $X2=2.7
+ $Y2=1.27
r46 11 12 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.61 $X2=2.7
+ $Y2=1.775
r47 10 16 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.105
+ $X2=2.7 $Y2=1.27
r48 7 12 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.755 $Y=2.225
+ $X2=2.755 $Y2=1.775
r49 3 10 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.68 $Y=0.615
+ $X2=2.68 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_M%B1 3 6 8 9 10 15 17
c29 8 0 3.22814e-20 $X=3.6 $Y=0.925
r30 15 18 80.5075 $w=5.7e-07 $l=5.05e-07 $layer=POLY_cond $X=3.36 $Y=1.1
+ $X2=3.36 $Y2=1.605
r31 15 17 48.5934 $w=5.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.36 $Y=1.1
+ $X2=3.36 $Y2=0.935
r32 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.48 $Y=1.1
+ $X2=3.48 $Y2=1.1
r33 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.54 $Y=1.295
+ $X2=3.54 $Y2=1.665
r34 9 16 7.74919 $w=2.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.54 $Y=1.295
+ $X2=3.54 $Y2=1.1
r35 8 16 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=3.54 $Y=0.925
+ $X2=3.54 $Y2=1.1
r36 6 18 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.15 $Y=2.225
+ $X2=3.15 $Y2=1.605
r37 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.15 $Y=0.615
+ $X2=3.15 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_M%X 1 2 8 10 11 12 13 14 15 16 34
r13 15 16 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=2.405
+ $X2=0.275 $Y2=2.775
r14 15 34 5.52212 $w=2.38e-07 $l=1.15e-07 $layer=LI1_cond $X=0.275 $Y=2.405
+ $X2=0.275 $Y2=2.29
r15 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r16 12 13 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r17 11 12 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.295
r18 11 44 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=0.8
r19 10 44 12.7603 $w=2.38e-07 $l=2.45e-07 $layer=LI1_cond $X=0.275 $Y=0.555
+ $X2=0.275 $Y2=0.8
r20 9 14 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=2.125 $X2=0.24
+ $Y2=2.035
r21 8 34 2.16083 $w=2.38e-07 $l=4.5e-08 $layer=LI1_cond $X=0.275 $Y=2.245
+ $X2=0.275 $Y2=2.29
r22 8 9 6.75802 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.275 $Y=2.245
+ $X2=0.275 $Y2=2.125
r23 2 34 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.015 $X2=0.29 $Y2=2.29
r24 1 10 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.405 $X2=0.29 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_M%VPWR 1 2 9 13 16 17 18 20 33 34 37
c41 9 0 1.83051e-19 $X=0.74 $Y=2.29
r42 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 27 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r50 25 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r54 20 22 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 18 31 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 16 30 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.2 $Y=3.33 $X2=3.12
+ $Y2=3.33
r58 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=3.33
+ $X2=3.365 $Y2=3.33
r59 15 33 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.53 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.53 $Y=3.33
+ $X2=3.365 $Y2=3.33
r61 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=3.245
+ $X2=3.365 $Y2=3.33
r62 11 13 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=3.365 $Y=3.245
+ $X2=3.365 $Y2=2.31
r63 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245 $X2=0.74
+ $Y2=3.33
r64 7 9 33.351 $w=3.28e-07 $l=9.55e-07 $layer=LI1_cond $X=0.74 $Y=3.245 $X2=0.74
+ $Y2=2.29
r65 2 13 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=2.015 $X2=3.365 $Y2=2.31
r66 1 9 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.015 $X2=0.74 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_M%VGND 1 2 9 11 15 17 19 29 30 33 36
r40 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r41 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 27 30 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r45 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r46 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r47 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.835
+ $Y2=0
r48 24 26 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.16
+ $Y2=0
r49 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r50 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.74
+ $Y2=0
r52 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.24
+ $Y2=0
r53 17 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r54 17 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r55 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0
r56 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.835 $Y=0.085
+ $X2=1.835 $Y2=0.55
r57 12 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.74
+ $Y2=0
r58 11 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=1.835
+ $Y2=0
r59 11 12 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.67 $Y=0 $X2=0.905
+ $Y2=0
r60 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0
r61 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0.55
r62 2 15 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.675
+ $Y=0.405 $X2=1.835 $Y2=0.55
r63 1 9 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.405 $X2=0.74 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_M%A_249_81# 1 2 3 12 14 15 19 20 21 22
c42 19 0 1.3507e-19 $X=2.465 $Y=0.55
c43 12 0 1.61613e-19 $X=1.385 $Y=0.68
r44 22 25 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.405 $Y=0.35 $X2=3.405
+ $Y2=0.55
r45 20 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0.35
+ $X2=3.405 $Y2=0.35
r46 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.24 $Y=0.35 $X2=2.55
+ $Y2=0.35
r47 17 19 16.6364 $w=1.88e-07 $l=2.85e-07 $layer=LI1_cond $X=2.455 $Y=0.835
+ $X2=2.455 $Y2=0.55
r48 16 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.455 $Y=0.435
+ $X2=2.55 $Y2=0.35
r49 16 19 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=2.455 $Y=0.435
+ $X2=2.455 $Y2=0.55
r50 14 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.36 $Y=0.92
+ $X2=2.455 $Y2=0.835
r51 14 15 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.36 $Y=0.92
+ $X2=1.49 $Y2=0.92
r52 10 15 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.395 $Y=0.835
+ $X2=1.49 $Y2=0.92
r53 10 12 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.395 $Y=0.835
+ $X2=1.395 $Y2=0.68
r54 3 25 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.405 $X2=3.405 $Y2=0.55
r55 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.405 $X2=2.465 $Y2=0.55
r56 1 12 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.245
+ $Y=0.405 $X2=1.385 $Y2=0.68
.ends

