* File: sky130_fd_sc_lp__nand2_1.spice
* Created: Fri Aug 28 10:46:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2_1.pex.spice"
.subckt sky130_fd_sc_lp__nand2_1  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1000 A_112_69# N_B_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.2226 PD=1.08 PS=2.21 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_112_69# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1008 PD=2.21 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75000.6 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
c_127 A_112_69# 0 2.39113e-20 $X=0.56 $Y=0.345
*
.include "sky130_fd_sc_lp__nand2_1.pxi.spice"
*
.ends
*
*
