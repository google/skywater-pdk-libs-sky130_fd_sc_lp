# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__nor4_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.210000 1.450000 1.435000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.345000 0.855000 1.615000 ;
        RECT 0.085000 1.615000 2.185000 1.785000 ;
        RECT 1.855000 1.425000 2.185000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.395000 1.425000 2.725000 1.695000 ;
        RECT 2.395000 1.695000 4.230000 1.865000 ;
        RECT 3.465000 1.425000 4.230000 1.695000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.990000 1.185000 3.295000 1.515000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.293600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.795000 0.265000 1.010000 0.870000 ;
        RECT 0.795000 0.870000 1.950000 1.040000 ;
        RECT 1.620000 1.040000 1.950000 1.085000 ;
        RECT 1.620000 1.085000 2.820000 1.255000 ;
        RECT 1.690000 0.255000 1.950000 0.870000 ;
        RECT 2.650000 0.255000 2.930000 0.845000 ;
        RECT 2.650000 0.845000 3.790000 1.005000 ;
        RECT 2.650000 1.005000 4.715000 1.015000 ;
        RECT 2.650000 1.015000 2.820000 1.085000 ;
        RECT 3.170000 2.035000 4.715000 2.205000 ;
        RECT 3.170000 2.205000 3.500000 2.335000 ;
        RECT 3.590000 1.015000 4.715000 1.175000 ;
        RECT 3.600000 0.255000 3.790000 0.845000 ;
        RECT 4.400000 1.175000 4.715000 2.035000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.330000  0.085000 0.625000 1.095000 ;
      RECT 0.330000  1.955000 2.240000 2.035000 ;
      RECT 0.330000  2.035000 2.530000 2.125000 ;
      RECT 0.330000  2.125000 0.625000 3.075000 ;
      RECT 0.795000  2.295000 1.915000 2.465000 ;
      RECT 0.795000  2.465000 1.020000 3.075000 ;
      RECT 1.190000  0.085000 1.520000 0.700000 ;
      RECT 1.190000  2.635000 1.520000 3.245000 ;
      RECT 1.690000  2.465000 1.915000 3.075000 ;
      RECT 2.085000  2.125000 2.530000 2.905000 ;
      RECT 2.085000  2.905000 4.360000 3.075000 ;
      RECT 2.150000  0.085000 2.480000 0.915000 ;
      RECT 2.740000  2.035000 3.000000 2.505000 ;
      RECT 2.740000  2.505000 3.930000 2.735000 ;
      RECT 3.100000  0.085000 3.430000 0.675000 ;
      RECT 3.960000  0.085000 4.290000 0.835000 ;
      RECT 4.100000  2.375000 4.360000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__nor4_2
END LIBRARY
