* File: sky130_fd_sc_lp__sdfxbp_2.pxi.spice
* Created: Fri Aug 28 11:30:24 2020
* 
x_PM_SKY130_FD_SC_LP__SDFXBP_2%SCD N_SCD_M1035_g N_SCD_M1023_g N_SCD_c_278_n
+ N_SCD_c_279_n N_SCD_c_280_n SCD SCD SCD N_SCD_c_282_n
+ PM_SKY130_FD_SC_LP__SDFXBP_2%SCD
x_PM_SKY130_FD_SC_LP__SDFXBP_2%D N_D_M1006_g N_D_M1014_g N_D_c_310_n N_D_c_315_n
+ D D N_D_c_312_n PM_SKY130_FD_SC_LP__SDFXBP_2%D
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_332_94# N_A_332_94#_M1003_d N_A_332_94#_M1005_s
+ N_A_332_94#_M1026_g N_A_332_94#_M1038_g N_A_332_94#_c_356_n
+ N_A_332_94#_c_357_n N_A_332_94#_c_358_n N_A_332_94#_c_359_n
+ N_A_332_94#_c_360_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_332_94#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%SCE N_SCE_M1020_g N_SCE_c_424_n N_SCE_M1009_g
+ N_SCE_c_414_n N_SCE_c_415_n N_SCE_M1003_g N_SCE_c_417_n N_SCE_M1005_g
+ N_SCE_c_426_n N_SCE_c_419_n N_SCE_c_420_n SCE SCE SCE N_SCE_c_421_n
+ N_SCE_c_422_n PM_SKY130_FD_SC_LP__SDFXBP_2%SCE
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_778_399# N_A_778_399#_M1013_s
+ N_A_778_399#_M1021_s N_A_778_399#_M1004_s N_A_778_399#_M1011_s
+ N_A_778_399#_M1033_g N_A_778_399#_M1031_g N_A_778_399#_c_496_n
+ N_A_778_399#_c_492_n N_A_778_399#_c_498_n N_A_778_399#_c_499_n
+ N_A_778_399#_c_500_n N_A_778_399#_c_501_n N_A_778_399#_c_502_n
+ N_A_778_399#_c_503_n N_A_778_399#_c_504_n N_A_778_399#_c_493_n
+ N_A_778_399#_c_494_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_778_399#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_733_21# N_A_733_21#_M1017_d N_A_733_21#_M1039_d
+ N_A_733_21#_c_605_n N_A_733_21#_c_606_n N_A_733_21#_c_607_n
+ N_A_733_21#_c_608_n N_A_733_21#_c_609_n N_A_733_21#_c_618_n
+ N_A_733_21#_c_619_n N_A_733_21#_c_610_n N_A_733_21#_M1013_g
+ N_A_733_21#_c_620_n N_A_733_21#_M1004_g N_A_733_21#_c_621_n
+ N_A_733_21#_c_622_n N_A_733_21#_c_611_n N_A_733_21#_c_623_n
+ N_A_733_21#_c_624_n N_A_733_21#_c_625_n N_A_733_21#_c_612_n
+ N_A_733_21#_c_613_n N_A_733_21#_c_614_n N_A_733_21#_c_626_n
+ N_A_733_21#_c_615_n N_A_733_21#_c_616_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_733_21#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_1102_93# N_A_1102_93#_M1016_s
+ N_A_1102_93#_M1027_s N_A_1102_93#_M1017_g N_A_1102_93#_c_733_n
+ N_A_1102_93#_c_734_n N_A_1102_93#_M1039_g N_A_1102_93#_c_735_n
+ N_A_1102_93#_M1021_g N_A_1102_93#_c_737_n N_A_1102_93#_M1034_g
+ N_A_1102_93#_c_751_n N_A_1102_93#_c_752_n N_A_1102_93#_c_738_n
+ N_A_1102_93#_c_739_n N_A_1102_93#_c_740_n N_A_1102_93#_c_741_n
+ N_A_1102_93#_c_742_n N_A_1102_93#_c_756_n N_A_1102_93#_c_757_n
+ N_A_1102_93#_c_743_n N_A_1102_93#_c_744_n N_A_1102_93#_c_745_n
+ N_A_1102_93#_c_746_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_1102_93#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_1188_93# N_A_1188_93#_M1018_d
+ N_A_1188_93#_M1001_d N_A_1188_93#_c_880_n N_A_1188_93#_M1010_g
+ N_A_1188_93#_c_881_n N_A_1188_93#_c_882_n N_A_1188_93#_c_898_n
+ N_A_1188_93#_M1024_g N_A_1188_93#_c_899_n N_A_1188_93#_c_900_n
+ N_A_1188_93#_M1027_g N_A_1188_93#_c_883_n N_A_1188_93#_M1016_g
+ N_A_1188_93#_c_902_n N_A_1188_93#_c_884_n N_A_1188_93#_M1011_g
+ N_A_1188_93#_c_886_n N_A_1188_93#_c_887_n N_A_1188_93#_M1015_g
+ N_A_1188_93#_c_889_n N_A_1188_93#_c_890_n N_A_1188_93#_c_891_n
+ N_A_1188_93#_c_892_n N_A_1188_93#_c_893_n N_A_1188_93#_c_907_n
+ N_A_1188_93#_c_894_n N_A_1188_93#_c_895_n N_A_1188_93#_c_896_n
+ N_A_1188_93#_c_897_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_1188_93#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%CLK N_CLK_M1001_g N_CLK_M1018_g CLK CLK CLK
+ N_CLK_c_1033_n N_CLK_c_1034_n PM_SKY130_FD_SC_LP__SDFXBP_2%CLK
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_2122_329# N_A_2122_329#_M1032_d
+ N_A_2122_329#_M1025_d N_A_2122_329#_M1000_g N_A_2122_329#_M1036_g
+ N_A_2122_329#_M1002_g N_A_2122_329#_M1022_g N_A_2122_329#_M1019_g
+ N_A_2122_329#_M1037_g N_A_2122_329#_c_1078_n N_A_2122_329#_c_1079_n
+ N_A_2122_329#_M1029_g N_A_2122_329#_M1007_g N_A_2122_329#_c_1092_n
+ N_A_2122_329#_c_1107_n N_A_2122_329#_c_1081_n N_A_2122_329#_c_1094_n
+ N_A_2122_329#_c_1095_n N_A_2122_329#_c_1190_p N_A_2122_329#_c_1096_n
+ N_A_2122_329#_c_1082_n N_A_2122_329#_c_1083_n N_A_2122_329#_c_1084_n
+ N_A_2122_329#_c_1099_n N_A_2122_329#_c_1085_n N_A_2122_329#_c_1100_n
+ N_A_2122_329#_c_1218_p PM_SKY130_FD_SC_LP__SDFXBP_2%A_2122_329#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_2008_122# N_A_2008_122#_M1021_d
+ N_A_2008_122#_M1011_d N_A_2008_122#_M1025_g N_A_2008_122#_M1032_g
+ N_A_2008_122#_c_1229_n N_A_2008_122#_c_1230_n N_A_2008_122#_c_1241_n
+ N_A_2008_122#_c_1231_n N_A_2008_122#_c_1232_n N_A_2008_122#_c_1233_n
+ N_A_2008_122#_c_1234_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_2008_122#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_2710_56# N_A_2710_56#_M1029_d
+ N_A_2710_56#_M1007_d N_A_2710_56#_c_1296_n N_A_2710_56#_M1012_g
+ N_A_2710_56#_M1008_g N_A_2710_56#_c_1298_n N_A_2710_56#_M1030_g
+ N_A_2710_56#_M1028_g N_A_2710_56#_c_1306_n N_A_2710_56#_c_1300_n
+ N_A_2710_56#_c_1301_n N_A_2710_56#_c_1307_n N_A_2710_56#_c_1302_n
+ N_A_2710_56#_c_1303_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_2710_56#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_27_489# N_A_27_489#_M1023_s N_A_27_489#_M1038_d
+ N_A_27_489#_c_1361_n N_A_27_489#_c_1362_n N_A_27_489#_c_1363_n
+ N_A_27_489#_c_1364_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_27_489#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%VPWR N_VPWR_M1023_d N_VPWR_M1005_d N_VPWR_M1004_d
+ N_VPWR_M1027_d N_VPWR_M1036_d N_VPWR_M1022_d N_VPWR_M1037_d N_VPWR_M1008_d
+ N_VPWR_M1028_d N_VPWR_c_1395_n N_VPWR_c_1396_n N_VPWR_c_1397_n N_VPWR_c_1398_n
+ N_VPWR_c_1399_n N_VPWR_c_1400_n N_VPWR_c_1401_n N_VPWR_c_1402_n
+ N_VPWR_c_1403_n N_VPWR_c_1404_n N_VPWR_c_1405_n N_VPWR_c_1406_n
+ N_VPWR_c_1407_n N_VPWR_c_1408_n VPWR N_VPWR_c_1409_n N_VPWR_c_1410_n
+ N_VPWR_c_1411_n N_VPWR_c_1412_n N_VPWR_c_1413_n N_VPWR_c_1414_n
+ N_VPWR_c_1415_n N_VPWR_c_1416_n N_VPWR_c_1417_n N_VPWR_c_1418_n
+ N_VPWR_c_1419_n N_VPWR_c_1420_n N_VPWR_c_1421_n N_VPWR_c_1394_n
+ PM_SKY130_FD_SC_LP__SDFXBP_2%VPWR
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_182_120# N_A_182_120#_M1020_d
+ N_A_182_120#_M1010_d N_A_182_120#_M1014_d N_A_182_120#_M1039_s
+ N_A_182_120#_c_1560_n N_A_182_120#_c_1583_n N_A_182_120#_c_1570_n
+ N_A_182_120#_c_1584_n N_A_182_120#_c_1561_n N_A_182_120#_c_1572_n
+ N_A_182_120#_c_1601_n N_A_182_120#_c_1562_n N_A_182_120#_c_1563_n
+ N_A_182_120#_c_1564_n N_A_182_120#_c_1574_n N_A_182_120#_c_1565_n
+ N_A_182_120#_c_1566_n N_A_182_120#_c_1567_n N_A_182_120#_c_1568_n
+ N_A_182_120#_c_1569_n N_A_182_120#_c_1575_n N_A_182_120#_c_1576_n
+ N_A_182_120#_c_1577_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_182_120#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%A_993_425# N_A_993_425#_M1033_d
+ N_A_993_425#_M1024_d N_A_993_425#_c_1724_n N_A_993_425#_c_1725_n
+ N_A_993_425#_c_1726_n PM_SKY130_FD_SC_LP__SDFXBP_2%A_993_425#
x_PM_SKY130_FD_SC_LP__SDFXBP_2%Q N_Q_M1002_d N_Q_M1022_s N_Q_c_1759_n
+ N_Q_c_1763_n N_Q_c_1776_n N_Q_c_1760_n Q N_Q_c_1761_n Q
+ PM_SKY130_FD_SC_LP__SDFXBP_2%Q
x_PM_SKY130_FD_SC_LP__SDFXBP_2%Q_N N_Q_N_M1012_d N_Q_N_M1008_s Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1803_n PM_SKY130_FD_SC_LP__SDFXBP_2%Q_N
x_PM_SKY130_FD_SC_LP__SDFXBP_2%VGND N_VGND_M1035_s N_VGND_M1026_d N_VGND_M1013_d
+ N_VGND_M1016_d N_VGND_M1000_d N_VGND_M1002_s N_VGND_M1019_s N_VGND_M1012_s
+ N_VGND_M1030_s N_VGND_c_1821_n N_VGND_c_1822_n N_VGND_c_1823_n N_VGND_c_1824_n
+ N_VGND_c_1825_n N_VGND_c_1826_n N_VGND_c_1827_n N_VGND_c_1828_n
+ N_VGND_c_1829_n N_VGND_c_1830_n N_VGND_c_1831_n N_VGND_c_1832_n
+ N_VGND_c_1833_n N_VGND_c_1834_n N_VGND_c_1835_n N_VGND_c_1836_n
+ N_VGND_c_1837_n N_VGND_c_1838_n N_VGND_c_1839_n VGND N_VGND_c_1840_n
+ N_VGND_c_1841_n N_VGND_c_1842_n N_VGND_c_1843_n N_VGND_c_1844_n
+ N_VGND_c_1845_n N_VGND_c_1846_n N_VGND_c_1847_n
+ PM_SKY130_FD_SC_LP__SDFXBP_2%VGND
cc_1 VNB N_SCD_c_278_n 0.021029f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.13
cc_2 VNB N_SCD_c_279_n 0.0249397f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.635
cc_3 VNB N_SCD_c_280_n 0.00147572f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.8
cc_4 VNB SCD 0.0313198f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_5 VNB N_SCD_c_282_n 0.0172447f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_6 VNB N_D_M1006_g 0.0234194f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.81
cc_7 VNB N_D_c_310_n 0.0101885f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.8
cc_8 VNB D 0.00652322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_D_c_312_n 0.0147056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_332_94#_M1026_g 0.0300461f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.13
cc_11 VNB N_A_332_94#_M1038_g 0.00624234f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_A_332_94#_c_356_n 0.0730893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_332_94#_c_357_n 0.00391059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_332_94#_c_358_n 0.00969211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_332_94#_c_359_n 0.0108476f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_16 VNB N_A_332_94#_c_360_n 0.0085635f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_17 VNB N_SCE_M1020_g 0.0536721f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.8
cc_18 VNB N_SCE_c_414_n 0.0932937f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_19 VNB N_SCE_c_415_n 0.0125232f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.13
cc_20 VNB N_SCE_M1003_g 0.032046f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_21 VNB N_SCE_c_417_n 0.0622702f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_22 VNB N_SCE_M1005_g 0.0419669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_SCE_c_419_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_24 VNB N_SCE_c_420_n 0.0209693f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.295
cc_25 VNB N_SCE_c_421_n 0.0439403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_SCE_c_422_n 0.0106895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_778_399#_M1031_g 0.0415025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_778_399#_c_492_n 0.0100709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_778_399#_c_493_n 0.0161736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_778_399#_c_494_n 0.0183173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_733_21#_c_605_n 0.0557474f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_32 VNB N_A_733_21#_c_606_n 0.00685818f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.635
cc_33 VNB N_A_733_21#_c_607_n 0.214641f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.8
cc_34 VNB N_A_733_21#_c_608_n 0.0102518f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_35 VNB N_A_733_21#_c_609_n 0.0332853f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_36 VNB N_A_733_21#_c_610_n 0.0165399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_733_21#_c_611_n 0.0050611f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.295
cc_38 VNB N_A_733_21#_c_612_n 0.00225276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_733_21#_c_613_n 0.0119289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_733_21#_c_614_n 0.00474004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_733_21#_c_615_n 0.00504555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_733_21#_c_616_n 0.0525418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1102_93#_M1017_g 0.0352358f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.13
cc_44 VNB N_A_1102_93#_c_733_n 0.0116232f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.8
cc_45 VNB N_A_1102_93#_c_734_n 0.00462334f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_46 VNB N_A_1102_93#_c_735_n 0.193401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1102_93#_M1021_g 0.0453169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1102_93#_c_737_n 0.149922f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_49 VNB N_A_1102_93#_c_738_n 0.0775122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1102_93#_c_739_n 0.00494649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1102_93#_c_740_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1102_93#_c_741_n 0.0101845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1102_93#_c_742_n 0.0151945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1102_93#_c_743_n 0.003938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1102_93#_c_744_n 0.0140516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1102_93#_c_745_n 0.0253259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1102_93#_c_746_n 0.0455555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1188_93#_c_880_n 0.0161952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1188_93#_c_881_n 0.0897734f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.635
cc_60 VNB N_A_1188_93#_c_882_n 0.00811513f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.8
cc_61 VNB N_A_1188_93#_c_883_n 0.0173574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1188_93#_c_884_n 0.0729875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1188_93#_M1011_g 0.00797807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1188_93#_c_886_n 0.0126673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1188_93#_c_887_n 0.0253898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1188_93#_M1015_g 0.0153636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1188_93#_c_889_n 0.0112507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1188_93#_c_890_n 0.005457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1188_93#_c_891_n 0.00324239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1188_93#_c_892_n 0.0143825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1188_93#_c_893_n 0.00359793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1188_93#_c_894_n 0.0149409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1188_93#_c_895_n 0.00262989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1188_93#_c_896_n 0.0570187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1188_93#_c_897_n 0.0134162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_CLK_M1001_g 0.0101465f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.81
cc_77 VNB CLK 0.0148626f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.635
cc_78 VNB N_CLK_c_1033_n 0.0301628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_CLK_c_1034_n 0.0198678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_2122_329#_M1000_g 0.0451668f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.13
cc_81 VNB N_A_2122_329#_M1002_g 0.0217101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_2122_329#_M1019_g 0.022462f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.295
cc_83 VNB N_A_2122_329#_c_1078_n 0.0171547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2122_329#_c_1079_n 0.0313678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2122_329#_M1029_g 0.0506526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2122_329#_c_1081_n 0.00311366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2122_329#_c_1082_n 0.00121322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_2122_329#_c_1083_n 0.0295259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2122_329#_c_1084_n 0.00518747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2122_329#_c_1085_n 0.00321009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2008_122#_c_1229_n 0.00301852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2008_122#_c_1230_n 0.00122652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2008_122#_c_1231_n 8.83744e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2008_122#_c_1232_n 0.0289983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2008_122#_c_1233_n 0.0240818f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=1.665
cc_96 VNB N_A_2008_122#_c_1234_n 0.0182003f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.035
cc_97 VNB N_A_2710_56#_c_1296_n 0.0191375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2710_56#_M1008_g 0.00745429f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_99 VNB N_A_2710_56#_c_1298_n 0.0212224f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_100 VNB N_A_2710_56#_M1028_g 0.0106048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_2710_56#_c_1300_n 0.0140355f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=1.295
cc_102 VNB N_A_2710_56#_c_1301_n 0.0159254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2710_56#_c_1302_n 0.00432803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2710_56#_c_1303_n 0.0722985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VPWR_c_1394_n 0.641339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_182_120#_c_1560_n 0.0257828f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_107 VNB N_A_182_120#_c_1561_n 0.00531416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_182_120#_c_1562_n 0.00885119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_182_120#_c_1563_n 0.0160309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_182_120#_c_1564_n 0.00232912f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=1.665
cc_111 VNB N_A_182_120#_c_1565_n 0.00544397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_182_120#_c_1566_n 0.0432245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_182_120#_c_1567_n 0.0043749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_182_120#_c_1568_n 0.00462201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_182_120#_c_1569_n 0.00790202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_Q_c_1759_n 0.0052374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_Q_c_1760_n 0.00205561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_Q_c_1761_n 0.00333592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB Q 0.00867962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_Q_N_c_1803_n 0.00147158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1821_n 0.0115788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1822_n 0.0387756f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.665
cc_123 VNB N_VGND_c_1823_n 0.0124477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1824_n 0.0111835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1825_n 0.0142452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1826_n 0.0212515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1827_n 0.00997922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1828_n 0.0132076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1829_n 0.00879025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1830_n 0.0107404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1831_n 0.0478624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1832_n 0.0407602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1833_n 0.00445561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1834_n 0.0663996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1835_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1836_n 0.0732409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1837_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1838_n 0.0823982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1839_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1840_n 0.0223124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1841_n 0.0152003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1842_n 0.0184941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1843_n 0.015753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1844_n 0.00547551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_1845_n 0.00663599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_1846_n 0.00525267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_1847_n 0.734899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VPB N_SCD_M1023_g 0.0534665f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.765
cc_149 VPB N_SCD_c_280_n 0.0158368f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.8
cc_150 VPB SCD 0.0250073f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_151 VPB N_D_M1014_g 0.0318733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_D_c_310_n 0.00852732f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.8
cc_153 VPB N_D_c_315_n 0.0142741f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_154 VPB D 0.0144358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_332_94#_M1038_g 0.058928f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_156 VPB N_A_332_94#_c_359_n 0.00974341f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.295
cc_157 VPB N_A_332_94#_c_360_n 0.0429013f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.295
cc_158 VPB N_SCE_M1020_g 0.0236537f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.8
cc_159 VPB N_SCE_c_424_n 0.0147674f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.765
cc_160 VPB N_SCE_M1005_g 0.0577478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_SCE_c_426_n 0.0177779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_778_399#_M1033_g 0.0233001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_778_399#_c_496_n 0.00131318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_778_399#_c_492_n 0.00988795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_778_399#_c_498_n 0.00746972f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.295
cc_166 VPB N_A_778_399#_c_499_n 0.00244457f $X=-0.19 $Y=1.655 $X2=0.445
+ $Y2=1.295
cc_167 VPB N_A_778_399#_c_500_n 0.0016651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_778_399#_c_501_n 0.0306144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_778_399#_c_502_n 0.017075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_778_399#_c_503_n 0.0637986f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=2.035
cc_171 VPB N_A_778_399#_c_504_n 0.00173079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_778_399#_c_493_n 0.0272287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_778_399#_c_494_n 0.037161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_733_21#_c_606_n 0.0813478f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.635
cc_175 VPB N_A_733_21#_c_618_n 0.032057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_733_21#_c_619_n 0.0110873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_733_21#_c_620_n 0.0209149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_733_21#_c_621_n 0.0804121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_733_21#_c_622_n 0.0499555f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.295
cc_180 VPB N_A_733_21#_c_623_n 0.00732516f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_733_21#_c_624_n 0.0117802f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.665
cc_182 VPB N_A_733_21#_c_625_n 0.0347977f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=2.035
cc_183 VPB N_A_733_21#_c_626_n 0.00160094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1102_93#_c_733_n 0.00712368f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.8
cc_185 VPB N_A_1102_93#_c_734_n 0.00328182f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_186 VPB N_A_1102_93#_M1039_g 0.0661093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_1102_93#_M1034_g 0.0378441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_1102_93#_c_751_n 0.103062f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1102_93#_c_752_n 0.012806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_1102_93#_c_738_n 0.079655f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_1102_93#_c_741_n 0.00270828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_1102_93#_c_742_n 0.0221066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_1102_93#_c_756_n 0.00552541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_1102_93#_c_757_n 0.00524866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_1102_93#_c_745_n 0.0219821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1188_93#_c_898_n 0.0175264f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_197 VPB N_A_1188_93#_c_899_n 0.170549f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_1188_93#_c_900_n 0.0123088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_1188_93#_M1027_g 0.0239041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_1188_93#_c_902_n 0.108256f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.295
cc_201 VPB N_A_1188_93#_M1011_g 0.0282856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1188_93#_c_891_n 0.00542374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1188_93#_c_892_n 0.0164593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1188_93#_c_893_n 0.00453081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1188_93#_c_907_n 0.00477907f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1188_93#_c_896_n 0.012586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_CLK_M1001_g 0.0277807f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.81
cc_208 VPB N_A_2122_329#_M1036_g 0.0301406f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_209 VPB N_A_2122_329#_M1022_g 0.0213361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_2122_329#_M1037_g 0.0221073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_2122_329#_c_1078_n 0.00617787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_2122_329#_c_1079_n 0.00307407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_2122_329#_M1007_g 0.0254816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_2122_329#_c_1092_n 0.00571877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_2122_329#_c_1081_n 9.52493e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_2122_329#_c_1094_n 0.00662951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_2122_329#_c_1095_n 0.00322351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_2122_329#_c_1096_n 0.00308177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_2122_329#_c_1083_n 0.00666066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_2122_329#_c_1084_n 0.0339255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_2122_329#_c_1099_n 0.0031053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_2122_329#_c_1100_n 0.00184524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_2008_122#_M1025_g 0.0208816f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.13
cc_224 VPB N_A_2008_122#_c_1230_n 0.0111538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_2008_122#_c_1232_n 0.00821442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_2710_56#_M1008_g 0.0243587f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_227 VPB N_A_2710_56#_M1028_g 0.0264965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_2710_56#_c_1306_n 0.0126422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_2710_56#_c_1307_n 0.0148151f $X=-0.19 $Y=1.655 $X2=0.445
+ $Y2=1.665
cc_230 VPB N_A_2710_56#_c_1302_n 0.00267157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_27_489#_c_1361_n 0.0240525f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.13
cc_232 VPB N_A_27_489#_c_1362_n 0.00644385f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.8
cc_233 VPB N_A_27_489#_c_1363_n 0.0101431f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_234 VPB N_A_27_489#_c_1364_n 0.0162501f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_235 VPB N_VPWR_c_1395_n 0.00290961f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.665
cc_236 VPB N_VPWR_c_1396_n 0.0100446f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1397_n 0.00446087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1398_n 0.0179447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1399_n 0.0102458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1400_n 0.0214869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1401_n 0.00738809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1402_n 0.0185012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1403_n 0.0245984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1404_n 0.00441053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1405_n 0.0107145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1406_n 0.0640459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1407_n 0.060386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1408_n 0.00477984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1409_n 0.0178675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1410_n 0.0245063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1411_n 0.0771721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1412_n 0.0834075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1413_n 0.0147084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1414_n 0.0180726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1415_n 0.00433013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1416_n 0.00436966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1417_n 0.00485836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1418_n 0.00629964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1419_n 0.00510939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1420_n 0.00510939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1421_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1394_n 0.107859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_182_120#_c_1570_n 0.00946133f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_182_120#_c_1561_n 0.0287123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_182_120#_c_1572_n 0.0117733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_182_120#_c_1562_n 0.0043808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_182_120#_c_1574_n 0.00772652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_182_120#_c_1575_n 0.0022919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_182_120#_c_1576_n 0.0167686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_182_120#_c_1577_n 0.00659518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_993_425#_c_1724_n 0.00880104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_993_425#_c_1725_n 0.00722605f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.635
cc_273 VPB N_A_993_425#_c_1726_n 0.0119265f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_Q_c_1763_n 0.00374052f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.13
cc_275 VPB Q 0.00429162f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_Q_N_c_1803_n 0.0013826f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 SCD N_D_M1006_g 4.72538e-19 $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_278 SCD D 0.051391f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_279 SCD N_D_c_312_n 9.94214e-19 $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_280 N_SCD_c_278_n N_SCE_M1020_g 0.0584578f $X=0.385 $Y=1.13 $X2=0 $Y2=0
cc_281 SCD N_SCE_M1020_g 0.0251523f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_282 N_SCD_M1023_g N_SCE_c_424_n 0.0187376f $X=0.475 $Y=2.765 $X2=0 $Y2=0
cc_283 N_SCD_c_279_n N_SCE_c_426_n 0.0584578f $X=0.385 $Y=1.635 $X2=0 $Y2=0
cc_284 N_SCD_M1023_g N_A_27_489#_c_1361_n 0.00790455f $X=0.475 $Y=2.765 $X2=0
+ $Y2=0
cc_285 N_SCD_M1023_g N_A_27_489#_c_1362_n 0.0111453f $X=0.475 $Y=2.765 $X2=0
+ $Y2=0
cc_286 SCD N_A_27_489#_c_1362_n 0.0306524f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_287 N_SCD_M1023_g N_A_27_489#_c_1363_n 0.00387142f $X=0.475 $Y=2.765 $X2=0
+ $Y2=0
cc_288 N_SCD_c_280_n N_A_27_489#_c_1363_n 7.12452e-19 $X=0.385 $Y=1.8 $X2=0
+ $Y2=0
cc_289 SCD N_A_27_489#_c_1363_n 0.0306939f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_290 N_SCD_M1023_g N_VPWR_c_1395_n 0.00334503f $X=0.475 $Y=2.765 $X2=0 $Y2=0
cc_291 N_SCD_M1023_g N_VPWR_c_1409_n 0.00539298f $X=0.475 $Y=2.765 $X2=0 $Y2=0
cc_292 N_SCD_M1023_g N_VPWR_c_1394_n 0.0108764f $X=0.475 $Y=2.765 $X2=0 $Y2=0
cc_293 N_SCD_c_278_n N_A_182_120#_c_1569_n 0.00117599f $X=0.385 $Y=1.13 $X2=0
+ $Y2=0
cc_294 SCD N_A_182_120#_c_1569_n 0.00580099f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_295 N_SCD_c_278_n N_VGND_c_1822_n 0.0120977f $X=0.385 $Y=1.13 $X2=0 $Y2=0
cc_296 SCD N_VGND_c_1822_n 0.0266208f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_297 N_SCD_c_282_n N_VGND_c_1822_n 0.00473799f $X=0.385 $Y=1.295 $X2=0 $Y2=0
cc_298 N_SCD_c_278_n N_VGND_c_1832_n 0.00356352f $X=0.385 $Y=1.13 $X2=0 $Y2=0
cc_299 N_SCD_c_278_n N_VGND_c_1847_n 0.00400172f $X=0.385 $Y=1.13 $X2=0 $Y2=0
cc_300 N_D_M1006_g N_A_332_94#_M1026_g 0.0321961f $X=1.265 $Y=0.81 $X2=0 $Y2=0
cc_301 D N_A_332_94#_M1026_g 0.00222335f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_302 N_D_c_312_n N_A_332_94#_M1026_g 0.0145645f $X=1.285 $Y=1.47 $X2=0 $Y2=0
cc_303 N_D_M1014_g N_A_332_94#_M1038_g 0.040072f $X=1.305 $Y=2.765 $X2=0 $Y2=0
cc_304 N_D_c_315_n N_A_332_94#_M1038_g 0.0145645f $X=1.285 $Y=1.975 $X2=0 $Y2=0
cc_305 D N_A_332_94#_M1038_g 0.0244358f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_306 D N_A_332_94#_c_356_n 0.00479585f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_307 N_D_c_310_n N_A_332_94#_c_357_n 0.0145645f $X=1.285 $Y=1.81 $X2=0 $Y2=0
cc_308 D N_A_332_94#_c_357_n 0.00349549f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_309 N_D_M1006_g N_SCE_M1020_g 0.0199612f $X=1.265 $Y=0.81 $X2=0 $Y2=0
cc_310 N_D_M1014_g N_SCE_M1020_g 0.00777143f $X=1.305 $Y=2.765 $X2=0 $Y2=0
cc_311 D N_SCE_M1020_g 0.00547469f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_312 N_D_c_312_n N_SCE_M1020_g 0.0398156f $X=1.285 $Y=1.47 $X2=0 $Y2=0
cc_313 N_D_M1006_g N_SCE_c_414_n 0.0103215f $X=1.265 $Y=0.81 $X2=0 $Y2=0
cc_314 N_D_M1014_g N_SCE_c_426_n 0.0642574f $X=1.305 $Y=2.765 $X2=0 $Y2=0
cc_315 N_D_M1014_g N_A_27_489#_c_1362_n 0.0137915f $X=1.305 $Y=2.765 $X2=0 $Y2=0
cc_316 N_D_c_315_n N_A_27_489#_c_1362_n 8.78229e-19 $X=1.285 $Y=1.975 $X2=0
+ $Y2=0
cc_317 D N_A_27_489#_c_1362_n 0.0603796f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_318 N_D_M1014_g N_A_27_489#_c_1364_n 8.45603e-19 $X=1.305 $Y=2.765 $X2=0
+ $Y2=0
cc_319 D N_A_27_489#_c_1364_n 0.00557574f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_320 N_D_M1014_g N_VPWR_c_1395_n 0.00226509f $X=1.305 $Y=2.765 $X2=0 $Y2=0
cc_321 N_D_M1014_g N_VPWR_c_1407_n 0.00537804f $X=1.305 $Y=2.765 $X2=0 $Y2=0
cc_322 N_D_M1014_g N_VPWR_c_1394_n 0.00981385f $X=1.305 $Y=2.765 $X2=0 $Y2=0
cc_323 N_D_M1006_g N_A_182_120#_c_1560_n 0.0115026f $X=1.265 $Y=0.81 $X2=0 $Y2=0
cc_324 D N_A_182_120#_c_1560_n 0.0508896f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_325 N_D_c_312_n N_A_182_120#_c_1560_n 0.00315953f $X=1.285 $Y=1.47 $X2=0
+ $Y2=0
cc_326 N_D_M1014_g N_A_182_120#_c_1583_n 0.00478342f $X=1.305 $Y=2.765 $X2=0
+ $Y2=0
cc_327 N_D_M1014_g N_A_182_120#_c_1584_n 0.00397311f $X=1.305 $Y=2.765 $X2=0
+ $Y2=0
cc_328 D N_A_182_120#_c_1561_n 0.030481f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_329 N_D_M1006_g N_A_182_120#_c_1569_n 0.0102782f $X=1.265 $Y=0.81 $X2=0 $Y2=0
cc_330 D N_A_182_120#_c_1569_n 0.0155719f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_331 N_D_c_312_n N_A_182_120#_c_1569_n 0.0020554f $X=1.285 $Y=1.47 $X2=0 $Y2=0
cc_332 N_D_M1006_g N_VGND_c_1823_n 0.00148901f $X=1.265 $Y=0.81 $X2=0 $Y2=0
cc_333 N_D_M1006_g N_VGND_c_1847_n 9.33152e-19 $X=1.265 $Y=0.81 $X2=0 $Y2=0
cc_334 N_A_332_94#_M1026_g N_SCE_c_414_n 0.0103186f $X=1.735 $Y=0.81 $X2=0 $Y2=0
cc_335 N_A_332_94#_M1026_g N_SCE_M1003_g 0.0158366f $X=1.735 $Y=0.81 $X2=0 $Y2=0
cc_336 N_A_332_94#_c_356_n N_SCE_M1003_g 0.00765124f $X=2.565 $Y=1.465 $X2=0
+ $Y2=0
cc_337 N_A_332_94#_c_358_n N_SCE_M1003_g 0.00410032f $X=2.635 $Y=0.72 $X2=0
+ $Y2=0
cc_338 N_A_332_94#_c_359_n N_SCE_M1003_g 0.00456309f $X=2.73 $Y=1.555 $X2=0
+ $Y2=0
cc_339 N_A_332_94#_c_358_n N_SCE_c_417_n 0.00869056f $X=2.635 $Y=0.72 $X2=0
+ $Y2=0
cc_340 N_A_332_94#_c_356_n N_SCE_M1005_g 0.0421895f $X=2.565 $Y=1.465 $X2=0
+ $Y2=0
cc_341 N_A_332_94#_c_359_n N_SCE_M1005_g 0.00870426f $X=2.73 $Y=1.555 $X2=0
+ $Y2=0
cc_342 N_A_332_94#_c_359_n N_SCE_c_420_n 8.68405e-19 $X=2.73 $Y=1.555 $X2=0
+ $Y2=0
cc_343 N_A_332_94#_c_358_n N_SCE_c_421_n 0.0034256f $X=2.635 $Y=0.72 $X2=0 $Y2=0
cc_344 N_A_332_94#_c_356_n N_SCE_c_422_n 6.3525e-19 $X=2.565 $Y=1.465 $X2=0
+ $Y2=0
cc_345 N_A_332_94#_c_358_n N_SCE_c_422_n 0.0228359f $X=2.635 $Y=0.72 $X2=0 $Y2=0
cc_346 N_A_332_94#_c_359_n N_SCE_c_422_n 0.0488432f $X=2.73 $Y=1.555 $X2=0 $Y2=0
cc_347 N_A_332_94#_M1038_g N_A_27_489#_c_1362_n 0.00908157f $X=1.735 $Y=2.765
+ $X2=0 $Y2=0
cc_348 N_A_332_94#_M1038_g N_A_27_489#_c_1364_n 0.00884574f $X=1.735 $Y=2.765
+ $X2=0 $Y2=0
cc_349 N_A_332_94#_M1038_g N_VPWR_c_1407_n 0.00351226f $X=1.735 $Y=2.765 $X2=0
+ $Y2=0
cc_350 N_A_332_94#_M1038_g N_VPWR_c_1394_n 0.0066371f $X=1.735 $Y=2.765 $X2=0
+ $Y2=0
cc_351 N_A_332_94#_M1026_g N_A_182_120#_c_1560_n 0.0159225f $X=1.735 $Y=0.81
+ $X2=0 $Y2=0
cc_352 N_A_332_94#_c_356_n N_A_182_120#_c_1560_n 0.014179f $X=2.565 $Y=1.465
+ $X2=0 $Y2=0
cc_353 N_A_332_94#_c_358_n N_A_182_120#_c_1560_n 0.012159f $X=2.635 $Y=0.72
+ $X2=0 $Y2=0
cc_354 N_A_332_94#_c_359_n N_A_182_120#_c_1560_n 0.0158786f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_355 N_A_332_94#_M1038_g N_A_182_120#_c_1570_n 0.0118572f $X=1.735 $Y=2.765
+ $X2=0 $Y2=0
cc_356 N_A_332_94#_M1026_g N_A_182_120#_c_1561_n 0.00419319f $X=1.735 $Y=0.81
+ $X2=0 $Y2=0
cc_357 N_A_332_94#_M1038_g N_A_182_120#_c_1561_n 0.0114846f $X=1.735 $Y=2.765
+ $X2=0 $Y2=0
cc_358 N_A_332_94#_c_356_n N_A_182_120#_c_1561_n 0.0151623f $X=2.565 $Y=1.465
+ $X2=0 $Y2=0
cc_359 N_A_332_94#_c_359_n N_A_182_120#_c_1561_n 0.113287f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_360 N_A_332_94#_c_360_n N_A_182_120#_c_1561_n 0.0126424f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_361 N_A_332_94#_M1005_s N_A_182_120#_c_1572_n 0.0109009f $X=2.64 $Y=2.405
+ $X2=0 $Y2=0
cc_362 N_A_332_94#_c_359_n N_A_182_120#_c_1572_n 0.0162236f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_363 N_A_332_94#_M1005_s N_A_182_120#_c_1601_n 0.0051139f $X=2.64 $Y=2.405
+ $X2=0 $Y2=0
cc_364 N_A_332_94#_c_359_n N_A_182_120#_c_1601_n 0.0140474f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_365 N_A_332_94#_c_359_n N_A_182_120#_c_1562_n 0.0139594f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_366 N_A_332_94#_M1026_g N_A_182_120#_c_1569_n 0.00146767f $X=1.735 $Y=0.81
+ $X2=0 $Y2=0
cc_367 N_A_332_94#_M1005_s N_A_182_120#_c_1576_n 0.00162106f $X=2.64 $Y=2.405
+ $X2=0 $Y2=0
cc_368 N_A_332_94#_c_359_n N_A_182_120#_c_1576_n 0.0430312f $X=2.73 $Y=1.555
+ $X2=0 $Y2=0
cc_369 N_A_332_94#_M1026_g N_VGND_c_1823_n 0.00937155f $X=1.735 $Y=0.81 $X2=0
+ $Y2=0
cc_370 N_A_332_94#_c_358_n N_VGND_c_1823_n 0.0115645f $X=2.635 $Y=0.72 $X2=0
+ $Y2=0
cc_371 N_A_332_94#_c_358_n N_VGND_c_1834_n 0.0120703f $X=2.635 $Y=0.72 $X2=0
+ $Y2=0
cc_372 N_A_332_94#_M1026_g N_VGND_c_1847_n 7.83848e-19 $X=1.735 $Y=0.81 $X2=0
+ $Y2=0
cc_373 N_A_332_94#_c_358_n N_VGND_c_1847_n 0.0148744f $X=2.635 $Y=0.72 $X2=0
+ $Y2=0
cc_374 N_SCE_M1005_g N_A_733_21#_c_605_n 0.0535205f $X=3.18 $Y=2.725 $X2=0 $Y2=0
cc_375 N_SCE_c_421_n N_A_733_21#_c_605_n 0.0126432f $X=3.12 $Y=0.43 $X2=0 $Y2=0
cc_376 N_SCE_c_422_n N_A_733_21#_c_605_n 0.00246702f $X=3.12 $Y=0.43 $X2=0 $Y2=0
cc_377 N_SCE_c_417_n N_A_733_21#_c_608_n 0.0126432f $X=2.955 $Y=0.185 $X2=0
+ $Y2=0
cc_378 N_SCE_c_424_n N_A_27_489#_c_1361_n 8.96335e-19 $X=0.945 $Y=2.335 $X2=0
+ $Y2=0
cc_379 N_SCE_c_424_n N_A_27_489#_c_1362_n 0.0108964f $X=0.945 $Y=2.335 $X2=0
+ $Y2=0
cc_380 N_SCE_c_426_n N_A_27_489#_c_1362_n 0.0131414f $X=0.945 $Y=2.26 $X2=0
+ $Y2=0
cc_381 N_SCE_c_424_n N_VPWR_c_1395_n 0.0118368f $X=0.945 $Y=2.335 $X2=0 $Y2=0
cc_382 N_SCE_c_426_n N_VPWR_c_1395_n 4.97993e-19 $X=0.945 $Y=2.26 $X2=0 $Y2=0
cc_383 N_SCE_M1005_g N_VPWR_c_1396_n 0.00323702f $X=3.18 $Y=2.725 $X2=0 $Y2=0
cc_384 N_SCE_c_424_n N_VPWR_c_1407_n 0.00554242f $X=0.945 $Y=2.335 $X2=0 $Y2=0
cc_385 N_SCE_M1005_g N_VPWR_c_1407_n 0.00416849f $X=3.18 $Y=2.725 $X2=0 $Y2=0
cc_386 N_SCE_c_424_n N_VPWR_c_1394_n 0.00938567f $X=0.945 $Y=2.335 $X2=0 $Y2=0
cc_387 N_SCE_M1005_g N_VPWR_c_1394_n 0.0064031f $X=3.18 $Y=2.725 $X2=0 $Y2=0
cc_388 N_SCE_M1003_g N_A_182_120#_c_1560_n 0.0120983f $X=2.245 $Y=0.81 $X2=0
+ $Y2=0
cc_389 N_SCE_c_424_n N_A_182_120#_c_1583_n 7.57559e-19 $X=0.945 $Y=2.335 $X2=0
+ $Y2=0
cc_390 N_SCE_c_424_n N_A_182_120#_c_1584_n 4.65814e-19 $X=0.945 $Y=2.335 $X2=0
+ $Y2=0
cc_391 N_SCE_M1005_g N_A_182_120#_c_1561_n 9.69243e-19 $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_392 N_SCE_M1005_g N_A_182_120#_c_1572_n 0.00716778f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_393 N_SCE_M1005_g N_A_182_120#_c_1601_n 0.0126671f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_394 N_SCE_M1005_g N_A_182_120#_c_1562_n 0.00732663f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_395 N_SCE_c_421_n N_A_182_120#_c_1562_n 0.00338635f $X=3.12 $Y=0.43 $X2=0
+ $Y2=0
cc_396 N_SCE_c_422_n N_A_182_120#_c_1562_n 0.0613922f $X=3.12 $Y=0.43 $X2=0
+ $Y2=0
cc_397 N_SCE_c_421_n N_A_182_120#_c_1564_n 0.00140172f $X=3.12 $Y=0.43 $X2=0
+ $Y2=0
cc_398 N_SCE_c_422_n N_A_182_120#_c_1564_n 0.011093f $X=3.12 $Y=0.43 $X2=0 $Y2=0
cc_399 N_SCE_M1020_g N_A_182_120#_c_1569_n 0.0124767f $X=0.835 $Y=0.81 $X2=0
+ $Y2=0
cc_400 N_SCE_c_414_n N_A_182_120#_c_1569_n 0.00336476f $X=2.17 $Y=0.185 $X2=0
+ $Y2=0
cc_401 N_SCE_M1005_g N_A_182_120#_c_1576_n 0.0291306f $X=3.18 $Y=2.725 $X2=0
+ $Y2=0
cc_402 N_SCE_c_422_n N_A_182_120#_c_1576_n 0.00925853f $X=3.12 $Y=0.43 $X2=0
+ $Y2=0
cc_403 N_SCE_M1020_g N_VGND_c_1822_n 0.00177543f $X=0.835 $Y=0.81 $X2=0 $Y2=0
cc_404 N_SCE_c_415_n N_VGND_c_1822_n 0.0102212f $X=0.91 $Y=0.185 $X2=0 $Y2=0
cc_405 N_SCE_c_414_n N_VGND_c_1823_n 0.0250258f $X=2.17 $Y=0.185 $X2=0 $Y2=0
cc_406 N_SCE_M1003_g N_VGND_c_1823_n 0.0134549f $X=2.245 $Y=0.81 $X2=0 $Y2=0
cc_407 N_SCE_c_415_n N_VGND_c_1832_n 0.033235f $X=0.91 $Y=0.185 $X2=0 $Y2=0
cc_408 N_SCE_c_414_n N_VGND_c_1834_n 0.0333701f $X=2.17 $Y=0.185 $X2=0 $Y2=0
cc_409 N_SCE_c_422_n N_VGND_c_1834_n 0.0168218f $X=3.12 $Y=0.43 $X2=0 $Y2=0
cc_410 N_SCE_c_414_n N_VGND_c_1847_n 0.0370201f $X=2.17 $Y=0.185 $X2=0 $Y2=0
cc_411 N_SCE_c_415_n N_VGND_c_1847_n 0.0107045f $X=0.91 $Y=0.185 $X2=0 $Y2=0
cc_412 N_SCE_c_417_n N_VGND_c_1847_n 0.0319627f $X=2.955 $Y=0.185 $X2=0 $Y2=0
cc_413 N_SCE_c_419_n N_VGND_c_1847_n 0.00830567f $X=2.245 $Y=0.185 $X2=0 $Y2=0
cc_414 N_SCE_c_422_n N_VGND_c_1847_n 0.00896488f $X=3.12 $Y=0.43 $X2=0 $Y2=0
cc_415 N_A_778_399#_c_492_n N_A_733_21#_c_605_n 0.0053578f $X=4.035 $Y=0.75
+ $X2=0 $Y2=0
cc_416 N_A_778_399#_c_496_n N_A_733_21#_c_606_n 0.0018323f $X=4.035 $Y=2.035
+ $X2=0 $Y2=0
cc_417 N_A_778_399#_c_492_n N_A_733_21#_c_606_n 0.00964795f $X=4.035 $Y=0.75
+ $X2=0 $Y2=0
cc_418 N_A_778_399#_M1031_g N_A_733_21#_c_607_n 0.0104164f $X=5.225 $Y=0.805
+ $X2=0 $Y2=0
cc_419 N_A_778_399#_c_492_n N_A_733_21#_c_609_n 0.0200813f $X=4.035 $Y=0.75
+ $X2=0 $Y2=0
cc_420 N_A_778_399#_c_498_n N_A_733_21#_c_609_n 0.00274637f $X=4.815 $Y=2.12
+ $X2=0 $Y2=0
cc_421 N_A_778_399#_c_492_n N_A_733_21#_c_610_n 0.00979278f $X=4.035 $Y=0.75
+ $X2=0 $Y2=0
cc_422 N_A_778_399#_M1033_g N_A_733_21#_c_620_n 0.0218433f $X=4.89 $Y=2.335
+ $X2=0 $Y2=0
cc_423 N_A_778_399#_c_492_n N_A_733_21#_c_620_n 5.97392e-19 $X=4.035 $Y=0.75
+ $X2=0 $Y2=0
cc_424 N_A_778_399#_c_498_n N_A_733_21#_c_620_n 0.0128224f $X=4.815 $Y=2.12
+ $X2=0 $Y2=0
cc_425 N_A_778_399#_M1033_g N_A_733_21#_c_621_n 0.00458044f $X=4.89 $Y=2.335
+ $X2=0 $Y2=0
cc_426 N_A_778_399#_c_498_n N_A_733_21#_c_624_n 0.0109584f $X=4.815 $Y=2.12
+ $X2=0 $Y2=0
cc_427 N_A_778_399#_c_500_n N_A_733_21#_c_624_n 0.00114423f $X=4.98 $Y=2.035
+ $X2=0 $Y2=0
cc_428 N_A_778_399#_c_501_n N_A_733_21#_c_624_n 0.0798441f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_429 N_A_778_399#_c_502_n N_A_733_21#_c_624_n 0.0154098f $X=6.71 $Y=2.365
+ $X2=0 $Y2=0
cc_430 N_A_778_399#_M1033_g N_A_733_21#_c_625_n 0.020181f $X=4.89 $Y=2.335 $X2=0
+ $Y2=0
cc_431 N_A_778_399#_c_498_n N_A_733_21#_c_625_n 8.05385e-19 $X=4.815 $Y=2.12
+ $X2=0 $Y2=0
cc_432 N_A_778_399#_c_500_n N_A_733_21#_c_625_n 0.00174f $X=4.98 $Y=2.035 $X2=0
+ $Y2=0
cc_433 N_A_778_399#_c_501_n N_A_733_21#_c_625_n 0.00474959f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_434 N_A_778_399#_M1031_g N_A_733_21#_c_612_n 0.00146306f $X=5.225 $Y=0.805
+ $X2=0 $Y2=0
cc_435 N_A_778_399#_c_502_n N_A_733_21#_c_626_n 0.0121085f $X=6.71 $Y=2.365
+ $X2=0 $Y2=0
cc_436 N_A_778_399#_c_504_n N_A_733_21#_c_626_n 0.0123843f $X=6.795 $Y=2.45
+ $X2=0 $Y2=0
cc_437 N_A_778_399#_c_503_n N_A_1102_93#_M1027_s 0.00923247f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_438 N_A_778_399#_M1031_g N_A_1102_93#_M1017_g 0.0380774f $X=5.225 $Y=0.805
+ $X2=0 $Y2=0
cc_439 N_A_778_399#_c_501_n N_A_1102_93#_c_734_n 0.00799427f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_440 N_A_778_399#_c_494_n N_A_1102_93#_c_734_n 0.0380774f $X=4.98 $Y=1.76
+ $X2=0 $Y2=0
cc_441 N_A_778_399#_c_501_n N_A_1102_93#_M1039_g 0.013631f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_442 N_A_778_399#_c_502_n N_A_1102_93#_M1039_g 0.00546306f $X=6.71 $Y=2.365
+ $X2=0 $Y2=0
cc_443 N_A_778_399#_c_494_n N_A_1102_93#_M1039_g 5.45335e-19 $X=4.98 $Y=1.76
+ $X2=0 $Y2=0
cc_444 N_A_778_399#_c_493_n N_A_1102_93#_c_735_n 0.00349749f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_445 N_A_778_399#_c_493_n N_A_1102_93#_M1021_g 0.00323346f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_446 N_A_778_399#_c_501_n N_A_1102_93#_c_741_n 0.0123062f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_447 N_A_778_399#_c_502_n N_A_1102_93#_c_741_n 0.00634272f $X=6.71 $Y=2.365
+ $X2=0 $Y2=0
cc_448 N_A_778_399#_c_501_n N_A_1102_93#_c_742_n 0.00349751f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_449 N_A_778_399#_c_503_n N_A_1102_93#_c_742_n 0.00245236f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_450 N_A_778_399#_c_502_n N_A_1102_93#_c_756_n 0.0187865f $X=6.71 $Y=2.365
+ $X2=0 $Y2=0
cc_451 N_A_778_399#_c_503_n N_A_1102_93#_c_756_n 0.0152028f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_452 N_A_778_399#_c_503_n N_A_1102_93#_c_757_n 0.0255118f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_453 N_A_778_399#_c_501_n N_A_1102_93#_c_745_n 0.0232517f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_454 N_A_778_399#_c_503_n N_A_1188_93#_M1001_d 0.00437555f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_455 N_A_778_399#_c_501_n N_A_1188_93#_c_898_n 0.00224027f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_456 N_A_778_399#_c_504_n N_A_1188_93#_c_898_n 0.00359296f $X=6.795 $Y=2.45
+ $X2=0 $Y2=0
cc_457 N_A_778_399#_c_503_n N_A_1188_93#_c_899_n 0.0238798f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_458 N_A_778_399#_c_504_n N_A_1188_93#_c_899_n 5.36664e-19 $X=6.795 $Y=2.45
+ $X2=0 $Y2=0
cc_459 N_A_778_399#_c_503_n N_A_1188_93#_M1027_g 0.0145366f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_460 N_A_778_399#_c_503_n N_A_1188_93#_c_902_n 0.0163606f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_461 N_A_778_399#_c_493_n N_A_1188_93#_c_884_n 0.0210666f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_462 N_A_778_399#_c_503_n N_A_1188_93#_M1011_g 0.00186686f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_463 N_A_778_399#_c_493_n N_A_1188_93#_M1011_g 0.0111249f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_464 N_A_778_399#_c_493_n N_A_1188_93#_c_887_n 9.04571e-19 $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_465 N_A_778_399#_c_503_n N_A_1188_93#_c_891_n 0.0180356f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_466 N_A_778_399#_c_503_n N_A_1188_93#_c_892_n 0.00261027f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_467 N_A_778_399#_c_503_n N_A_1188_93#_c_893_n 0.0111542f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_468 N_A_778_399#_c_493_n N_A_1188_93#_c_893_n 0.00562536f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_469 N_A_778_399#_c_503_n N_A_1188_93#_c_907_n 0.021804f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_470 N_A_778_399#_c_493_n N_A_1188_93#_c_894_n 0.011712f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_471 N_A_778_399#_c_493_n N_A_1188_93#_c_895_n 0.0184516f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_472 N_A_778_399#_c_503_n N_A_1188_93#_c_896_n 0.00108886f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_473 N_A_778_399#_c_493_n N_A_1188_93#_c_896_n 0.00892582f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_474 N_A_778_399#_c_503_n N_CLK_M1001_g 0.0125255f $X=9.615 $Y=2.45 $X2=0
+ $Y2=0
cc_475 N_A_778_399#_c_493_n N_A_2008_122#_c_1229_n 0.028318f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_476 N_A_778_399#_c_503_n N_A_2008_122#_c_1230_n 0.016921f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_477 N_A_778_399#_c_493_n N_A_2008_122#_c_1230_n 0.0441313f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_478 N_A_778_399#_c_493_n N_A_2008_122#_c_1241_n 0.0134167f $X=9.75 $Y=0.825
+ $X2=0 $Y2=0
cc_479 N_A_778_399#_c_498_n N_VPWR_M1004_d 0.00284683f $X=4.815 $Y=2.12 $X2=0
+ $Y2=0
cc_480 N_A_778_399#_c_503_n N_VPWR_M1027_d 0.00990541f $X=9.615 $Y=2.45 $X2=0
+ $Y2=0
cc_481 N_A_778_399#_c_503_n N_VPWR_c_1398_n 0.0260861f $X=9.615 $Y=2.45 $X2=0
+ $Y2=0
cc_482 N_A_778_399#_c_503_n N_VPWR_c_1412_n 0.00625425f $X=9.615 $Y=2.45 $X2=0
+ $Y2=0
cc_483 N_A_778_399#_M1033_g N_VPWR_c_1394_n 9.73184e-19 $X=4.89 $Y=2.335 $X2=0
+ $Y2=0
cc_484 N_A_778_399#_c_503_n N_VPWR_c_1394_n 0.086009f $X=9.615 $Y=2.45 $X2=0
+ $Y2=0
cc_485 N_A_778_399#_c_504_n N_VPWR_c_1394_n 3.46594e-19 $X=6.795 $Y=2.45 $X2=0
+ $Y2=0
cc_486 N_A_778_399#_c_492_n N_A_182_120#_c_1562_n 0.100547f $X=4.035 $Y=0.75
+ $X2=0 $Y2=0
cc_487 N_A_778_399#_c_492_n N_A_182_120#_c_1563_n 0.0232792f $X=4.035 $Y=0.75
+ $X2=0 $Y2=0
cc_488 N_A_778_399#_M1004_s N_A_182_120#_c_1574_n 0.00797683f $X=3.89 $Y=1.995
+ $X2=0 $Y2=0
cc_489 N_A_778_399#_M1033_g N_A_182_120#_c_1574_n 0.0108672f $X=4.89 $Y=2.335
+ $X2=0 $Y2=0
cc_490 N_A_778_399#_c_496_n N_A_182_120#_c_1574_n 0.0268637f $X=4.035 $Y=2.035
+ $X2=0 $Y2=0
cc_491 N_A_778_399#_c_498_n N_A_182_120#_c_1574_n 0.0524082f $X=4.815 $Y=2.12
+ $X2=0 $Y2=0
cc_492 N_A_778_399#_c_501_n N_A_182_120#_c_1574_n 0.00859654f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_493 N_A_778_399#_c_494_n N_A_182_120#_c_1574_n 0.00126749f $X=4.98 $Y=1.76
+ $X2=0 $Y2=0
cc_494 N_A_778_399#_M1031_g N_A_182_120#_c_1565_n 0.0043702f $X=5.225 $Y=0.805
+ $X2=0 $Y2=0
cc_495 N_A_778_399#_c_492_n N_A_182_120#_c_1565_n 0.0299528f $X=4.035 $Y=0.75
+ $X2=0 $Y2=0
cc_496 N_A_778_399#_M1031_g N_A_182_120#_c_1566_n 0.0166126f $X=5.225 $Y=0.805
+ $X2=0 $Y2=0
cc_497 N_A_778_399#_c_498_n N_A_182_120#_c_1566_n 0.00938636f $X=4.815 $Y=2.12
+ $X2=0 $Y2=0
cc_498 N_A_778_399#_c_499_n N_A_182_120#_c_1566_n 0.0258515f $X=4.98 $Y=1.845
+ $X2=0 $Y2=0
cc_499 N_A_778_399#_c_501_n N_A_182_120#_c_1566_n 0.0886224f $X=6.625 $Y=1.76
+ $X2=0 $Y2=0
cc_500 N_A_778_399#_c_494_n N_A_182_120#_c_1566_n 0.00942401f $X=4.98 $Y=1.76
+ $X2=0 $Y2=0
cc_501 N_A_778_399#_c_492_n N_A_182_120#_c_1567_n 0.0143382f $X=4.035 $Y=0.75
+ $X2=0 $Y2=0
cc_502 N_A_778_399#_c_498_n N_A_182_120#_c_1567_n 0.00624779f $X=4.815 $Y=2.12
+ $X2=0 $Y2=0
cc_503 N_A_778_399#_c_496_n N_A_182_120#_c_1576_n 0.0144085f $X=4.035 $Y=2.035
+ $X2=0 $Y2=0
cc_504 N_A_778_399#_c_498_n N_A_993_425#_M1033_d 0.00219038f $X=4.815 $Y=2.12
+ $X2=-0.19 $Y2=-0.245
cc_505 N_A_778_399#_c_503_n N_A_993_425#_M1024_d 0.00151382f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_506 N_A_778_399#_c_504_n N_A_993_425#_M1024_d 0.00194255f $X=6.795 $Y=2.45
+ $X2=0 $Y2=0
cc_507 N_A_778_399#_c_503_n N_A_993_425#_c_1726_n 0.0120032f $X=9.615 $Y=2.45
+ $X2=0 $Y2=0
cc_508 N_A_778_399#_c_504_n N_A_993_425#_c_1726_n 0.0140604f $X=6.795 $Y=2.45
+ $X2=0 $Y2=0
cc_509 N_A_778_399#_M1031_g N_VGND_c_1824_n 0.0211692f $X=5.225 $Y=0.805 $X2=0
+ $Y2=0
cc_510 N_A_778_399#_c_493_n N_VGND_c_1838_n 0.00434909f $X=9.75 $Y=0.825 $X2=0
+ $Y2=0
cc_511 N_A_778_399#_M1031_g N_VGND_c_1847_n 9.39239e-19 $X=5.225 $Y=0.805 $X2=0
+ $Y2=0
cc_512 N_A_778_399#_c_493_n N_VGND_c_1847_n 0.00667531f $X=9.75 $Y=0.825 $X2=0
+ $Y2=0
cc_513 N_A_733_21#_c_607_n N_A_1102_93#_M1017_g 0.0101494f $X=6.495 $Y=0.18
+ $X2=0 $Y2=0
cc_514 N_A_733_21#_c_612_n N_A_1102_93#_M1017_g 0.0110795f $X=5.8 $Y=0.8 $X2=0
+ $Y2=0
cc_515 N_A_733_21#_c_625_n N_A_1102_93#_c_734_n 0.00898296f $X=5.565 $Y=2.11
+ $X2=0 $Y2=0
cc_516 N_A_733_21#_c_622_n N_A_1102_93#_M1039_g 0.0182664f $X=5.475 $Y=3.075
+ $X2=0 $Y2=0
cc_517 N_A_733_21#_c_624_n N_A_1102_93#_M1039_g 0.0161483f $X=6.115 $Y=2.11
+ $X2=0 $Y2=0
cc_518 N_A_733_21#_c_625_n N_A_1102_93#_M1039_g 0.0171259f $X=5.565 $Y=2.11
+ $X2=0 $Y2=0
cc_519 N_A_733_21#_c_626_n N_A_1102_93#_M1039_g 0.0123806f $X=6.28 $Y=2.65 $X2=0
+ $Y2=0
cc_520 N_A_733_21#_c_615_n N_A_1102_93#_c_744_n 0.0481921f $X=6.66 $Y=0.35 $X2=0
+ $Y2=0
cc_521 N_A_733_21#_c_616_n N_A_1102_93#_c_744_n 0.00911352f $X=6.66 $Y=0.35
+ $X2=0 $Y2=0
cc_522 N_A_733_21#_c_607_n N_A_1102_93#_c_746_n 0.0235678f $X=6.495 $Y=0.18
+ $X2=0 $Y2=0
cc_523 N_A_733_21#_c_607_n N_A_1188_93#_c_880_n 0.00881852f $X=6.495 $Y=0.18
+ $X2=0 $Y2=0
cc_524 N_A_733_21#_c_612_n N_A_1188_93#_c_880_n 0.0018582f $X=5.8 $Y=0.8 $X2=0
+ $Y2=0
cc_525 N_A_733_21#_c_613_n N_A_1188_93#_c_880_n 0.00376655f $X=6.495 $Y=0.35
+ $X2=0 $Y2=0
cc_526 N_A_733_21#_c_615_n N_A_1188_93#_c_880_n 6.61321e-19 $X=6.66 $Y=0.35
+ $X2=0 $Y2=0
cc_527 N_A_733_21#_c_616_n N_A_1188_93#_c_880_n 0.00701551f $X=6.66 $Y=0.35
+ $X2=0 $Y2=0
cc_528 N_A_733_21#_c_613_n N_A_1188_93#_c_881_n 0.00381827f $X=6.495 $Y=0.35
+ $X2=0 $Y2=0
cc_529 N_A_733_21#_c_615_n N_A_1188_93#_c_881_n 0.00205923f $X=6.66 $Y=0.35
+ $X2=0 $Y2=0
cc_530 N_A_733_21#_c_616_n N_A_1188_93#_c_881_n 0.0144912f $X=6.66 $Y=0.35 $X2=0
+ $Y2=0
cc_531 N_A_733_21#_c_626_n N_A_1188_93#_c_898_n 0.0117115f $X=6.28 $Y=2.65 $X2=0
+ $Y2=0
cc_532 N_A_733_21#_c_606_n N_VPWR_c_1396_n 0.0143512f $X=3.74 $Y=3.075 $X2=0
+ $Y2=0
cc_533 N_A_733_21#_c_606_n N_VPWR_c_1397_n 0.00119589f $X=3.74 $Y=3.075 $X2=0
+ $Y2=0
cc_534 N_A_733_21#_c_620_n N_VPWR_c_1397_n 0.0121029f $X=4.365 $Y=3.075 $X2=0
+ $Y2=0
cc_535 N_A_733_21#_c_621_n N_VPWR_c_1397_n 0.0181117f $X=5.4 $Y=3.15 $X2=0 $Y2=0
cc_536 N_A_733_21#_c_623_n N_VPWR_c_1397_n 0.00460513f $X=4.365 $Y=3.15 $X2=0
+ $Y2=0
cc_537 N_A_733_21#_c_619_n N_VPWR_c_1410_n 0.0281095f $X=3.815 $Y=3.15 $X2=0
+ $Y2=0
cc_538 N_A_733_21#_c_621_n N_VPWR_c_1411_n 0.0214856f $X=5.4 $Y=3.15 $X2=0 $Y2=0
cc_539 N_A_733_21#_c_618_n N_VPWR_c_1394_n 0.0140473f $X=4.29 $Y=3.15 $X2=0
+ $Y2=0
cc_540 N_A_733_21#_c_619_n N_VPWR_c_1394_n 0.00617379f $X=3.815 $Y=3.15 $X2=0
+ $Y2=0
cc_541 N_A_733_21#_c_621_n N_VPWR_c_1394_n 0.022739f $X=5.4 $Y=3.15 $X2=0 $Y2=0
cc_542 N_A_733_21#_c_623_n N_VPWR_c_1394_n 0.00364716f $X=4.365 $Y=3.15 $X2=0
+ $Y2=0
cc_543 N_A_733_21#_c_606_n N_A_182_120#_c_1601_n 9.15724e-19 $X=3.74 $Y=3.075
+ $X2=0 $Y2=0
cc_544 N_A_733_21#_c_605_n N_A_182_120#_c_1562_n 0.0194916f $X=3.74 $Y=1.345
+ $X2=0 $Y2=0
cc_545 N_A_733_21#_c_606_n N_A_182_120#_c_1562_n 0.0118281f $X=3.74 $Y=3.075
+ $X2=0 $Y2=0
cc_546 N_A_733_21#_c_610_n N_A_182_120#_c_1562_n 0.00110599f $X=4.25 $Y=1.345
+ $X2=0 $Y2=0
cc_547 N_A_733_21#_c_611_n N_A_182_120#_c_1562_n 0.00394409f $X=3.74 $Y=1.42
+ $X2=0 $Y2=0
cc_548 N_A_733_21#_c_605_n N_A_182_120#_c_1563_n 0.0116028f $X=3.74 $Y=1.345
+ $X2=0 $Y2=0
cc_549 N_A_733_21#_c_607_n N_A_182_120#_c_1563_n 0.0123859f $X=6.495 $Y=0.18
+ $X2=0 $Y2=0
cc_550 N_A_733_21#_c_610_n N_A_182_120#_c_1563_n 0.00349128f $X=4.25 $Y=1.345
+ $X2=0 $Y2=0
cc_551 N_A_733_21#_c_605_n N_A_182_120#_c_1564_n 0.00225865f $X=3.74 $Y=1.345
+ $X2=0 $Y2=0
cc_552 N_A_733_21#_c_606_n N_A_182_120#_c_1574_n 0.0132328f $X=3.74 $Y=3.075
+ $X2=0 $Y2=0
cc_553 N_A_733_21#_c_618_n N_A_182_120#_c_1574_n 0.00693209f $X=4.29 $Y=3.15
+ $X2=0 $Y2=0
cc_554 N_A_733_21#_c_620_n N_A_182_120#_c_1574_n 0.0130435f $X=4.365 $Y=3.075
+ $X2=0 $Y2=0
cc_555 N_A_733_21#_c_621_n N_A_182_120#_c_1574_n 0.00429627f $X=5.4 $Y=3.15
+ $X2=0 $Y2=0
cc_556 N_A_733_21#_c_622_n N_A_182_120#_c_1574_n 0.0115351f $X=5.475 $Y=3.075
+ $X2=0 $Y2=0
cc_557 N_A_733_21#_c_624_n N_A_182_120#_c_1574_n 0.0142205f $X=6.115 $Y=2.11
+ $X2=0 $Y2=0
cc_558 N_A_733_21#_c_625_n N_A_182_120#_c_1574_n 0.00133948f $X=5.565 $Y=2.11
+ $X2=0 $Y2=0
cc_559 N_A_733_21#_c_610_n N_A_182_120#_c_1565_n 0.0196715f $X=4.25 $Y=1.345
+ $X2=0 $Y2=0
cc_560 N_A_733_21#_c_612_n N_A_182_120#_c_1566_n 0.0108774f $X=5.8 $Y=0.8 $X2=0
+ $Y2=0
cc_561 N_A_733_21#_c_610_n N_A_182_120#_c_1567_n 0.00488311f $X=4.25 $Y=1.345
+ $X2=0 $Y2=0
cc_562 N_A_733_21#_c_620_n N_A_182_120#_c_1567_n 0.0015403f $X=4.365 $Y=3.075
+ $X2=0 $Y2=0
cc_563 N_A_733_21#_c_613_n N_A_182_120#_c_1568_n 0.013334f $X=6.495 $Y=0.35
+ $X2=0 $Y2=0
cc_564 N_A_733_21#_c_615_n N_A_182_120#_c_1568_n 0.0158849f $X=6.66 $Y=0.35
+ $X2=0 $Y2=0
cc_565 N_A_733_21#_c_616_n N_A_182_120#_c_1568_n 0.00165505f $X=6.66 $Y=0.35
+ $X2=0 $Y2=0
cc_566 N_A_733_21#_c_606_n N_A_182_120#_c_1576_n 0.0147174f $X=3.74 $Y=3.075
+ $X2=0 $Y2=0
cc_567 N_A_733_21#_c_620_n N_A_182_120#_c_1576_n 8.57872e-19 $X=4.365 $Y=3.075
+ $X2=0 $Y2=0
cc_568 N_A_733_21#_c_622_n N_A_182_120#_c_1577_n 0.00567329f $X=5.475 $Y=3.075
+ $X2=0 $Y2=0
cc_569 N_A_733_21#_c_624_n N_A_182_120#_c_1577_n 0.026043f $X=6.115 $Y=2.11
+ $X2=0 $Y2=0
cc_570 N_A_733_21#_c_625_n N_A_182_120#_c_1577_n 0.00308118f $X=5.565 $Y=2.11
+ $X2=0 $Y2=0
cc_571 N_A_733_21#_c_626_n N_A_182_120#_c_1577_n 0.0180576f $X=6.28 $Y=2.65
+ $X2=0 $Y2=0
cc_572 N_A_733_21#_M1039_d N_A_993_425#_c_1724_n 0.00176461f $X=6.14 $Y=2.505
+ $X2=0 $Y2=0
cc_573 N_A_733_21#_c_622_n N_A_993_425#_c_1724_n 0.0121028f $X=5.475 $Y=3.075
+ $X2=0 $Y2=0
cc_574 N_A_733_21#_c_625_n N_A_993_425#_c_1724_n 2.47351e-19 $X=5.565 $Y=2.11
+ $X2=0 $Y2=0
cc_575 N_A_733_21#_c_626_n N_A_993_425#_c_1724_n 0.0160514f $X=6.28 $Y=2.65
+ $X2=0 $Y2=0
cc_576 N_A_733_21#_c_620_n N_A_993_425#_c_1725_n 9.16525e-19 $X=4.365 $Y=3.075
+ $X2=0 $Y2=0
cc_577 N_A_733_21#_c_621_n N_A_993_425#_c_1725_n 0.0085605f $X=5.4 $Y=3.15 $X2=0
+ $Y2=0
cc_578 N_A_733_21#_c_622_n N_A_993_425#_c_1725_n 0.00969171f $X=5.475 $Y=3.075
+ $X2=0 $Y2=0
cc_579 N_A_733_21#_c_607_n N_VGND_c_1824_n 0.0261591f $X=6.495 $Y=0.18 $X2=0
+ $Y2=0
cc_580 N_A_733_21#_c_612_n N_VGND_c_1824_n 0.0155312f $X=5.8 $Y=0.8 $X2=0 $Y2=0
cc_581 N_A_733_21#_c_614_n N_VGND_c_1824_n 0.00627754f $X=5.92 $Y=0.35 $X2=0
+ $Y2=0
cc_582 N_A_733_21#_c_608_n N_VGND_c_1834_n 0.024949f $X=3.815 $Y=0.18 $X2=0
+ $Y2=0
cc_583 N_A_733_21#_c_607_n N_VGND_c_1836_n 0.0466427f $X=6.495 $Y=0.18 $X2=0
+ $Y2=0
cc_584 N_A_733_21#_c_613_n N_VGND_c_1836_n 0.0347991f $X=6.495 $Y=0.35 $X2=0
+ $Y2=0
cc_585 N_A_733_21#_c_614_n N_VGND_c_1836_n 0.0192498f $X=5.92 $Y=0.35 $X2=0
+ $Y2=0
cc_586 N_A_733_21#_c_615_n N_VGND_c_1836_n 0.0208937f $X=6.66 $Y=0.35 $X2=0
+ $Y2=0
cc_587 N_A_733_21#_c_607_n N_VGND_c_1847_n 0.081423f $X=6.495 $Y=0.18 $X2=0
+ $Y2=0
cc_588 N_A_733_21#_c_608_n N_VGND_c_1847_n 0.0049074f $X=3.815 $Y=0.18 $X2=0
+ $Y2=0
cc_589 N_A_733_21#_c_613_n N_VGND_c_1847_n 0.0191583f $X=6.495 $Y=0.35 $X2=0
+ $Y2=0
cc_590 N_A_733_21#_c_614_n N_VGND_c_1847_n 0.00989952f $X=5.92 $Y=0.35 $X2=0
+ $Y2=0
cc_591 N_A_733_21#_c_615_n N_VGND_c_1847_n 0.0112005f $X=6.66 $Y=0.35 $X2=0
+ $Y2=0
cc_592 N_A_1102_93#_M1017_g N_A_1188_93#_c_880_n 0.0194219f $X=5.585 $Y=0.805
+ $X2=0 $Y2=0
cc_593 N_A_1102_93#_c_739_n N_A_1188_93#_c_881_n 0.0258639f $X=6.065 $Y=1.59
+ $X2=0 $Y2=0
cc_594 N_A_1102_93#_c_741_n N_A_1188_93#_c_881_n 0.0147817f $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_595 N_A_1102_93#_c_742_n N_A_1188_93#_c_881_n 0.02174f $X=7.09 $Y=1.65 $X2=0
+ $Y2=0
cc_596 N_A_1102_93#_c_757_n N_A_1188_93#_c_881_n 0.00281772f $X=7.35 $Y=2.11
+ $X2=0 $Y2=0
cc_597 N_A_1102_93#_c_743_n N_A_1188_93#_c_881_n 0.00628922f $X=7.63 $Y=0.805
+ $X2=0 $Y2=0
cc_598 N_A_1102_93#_c_744_n N_A_1188_93#_c_881_n 0.00577946f $X=7.23 $Y=0.35
+ $X2=0 $Y2=0
cc_599 N_A_1102_93#_c_746_n N_A_1188_93#_c_881_n 0.00410004f $X=7.23 $Y=0.18
+ $X2=0 $Y2=0
cc_600 N_A_1102_93#_c_733_n N_A_1188_93#_c_882_n 0.0258639f $X=5.99 $Y=1.59
+ $X2=0 $Y2=0
cc_601 N_A_1102_93#_M1039_g N_A_1188_93#_c_898_n 0.0153726f $X=6.065 $Y=2.715
+ $X2=0 $Y2=0
cc_602 N_A_1102_93#_c_745_n N_A_1188_93#_c_898_n 0.00158068f $X=6.925 $Y=1.65
+ $X2=0 $Y2=0
cc_603 N_A_1102_93#_c_741_n N_A_1188_93#_M1027_g 0.00324803f $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_604 N_A_1102_93#_c_757_n N_A_1188_93#_M1027_g 0.0108682f $X=7.35 $Y=2.11
+ $X2=0 $Y2=0
cc_605 N_A_1102_93#_c_735_n N_A_1188_93#_c_883_n 0.0104164f $X=9.89 $Y=0.18
+ $X2=0 $Y2=0
cc_606 N_A_1102_93#_c_741_n N_A_1188_93#_c_883_n 0.00308771f $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_607 N_A_1102_93#_c_744_n N_A_1188_93#_c_883_n 0.00212542f $X=7.23 $Y=0.35
+ $X2=0 $Y2=0
cc_608 N_A_1102_93#_c_746_n N_A_1188_93#_c_883_n 0.00148679f $X=7.23 $Y=0.18
+ $X2=0 $Y2=0
cc_609 N_A_1102_93#_M1021_g N_A_1188_93#_c_884_n 0.0124997f $X=9.965 $Y=0.82
+ $X2=0 $Y2=0
cc_610 N_A_1102_93#_M1034_g N_A_1188_93#_M1011_g 0.0146485f $X=10.505 $Y=2.525
+ $X2=0 $Y2=0
cc_611 N_A_1102_93#_M1021_g N_A_1188_93#_M1015_g 0.0124557f $X=9.965 $Y=0.82
+ $X2=0 $Y2=0
cc_612 N_A_1102_93#_c_737_n N_A_1188_93#_M1015_g 0.00959659f $X=11.885 $Y=0.18
+ $X2=0 $Y2=0
cc_613 N_A_1102_93#_c_741_n N_A_1188_93#_c_891_n 0.00753363f $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_614 N_A_1102_93#_c_742_n N_A_1188_93#_c_891_n 9.2068e-19 $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_615 N_A_1102_93#_c_741_n N_A_1188_93#_c_892_n 9.54061e-19 $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_616 N_A_1102_93#_c_742_n N_A_1188_93#_c_892_n 0.0128748f $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_617 N_A_1102_93#_c_735_n N_A_1188_93#_c_894_n 0.0128746f $X=9.89 $Y=0.18
+ $X2=0 $Y2=0
cc_618 N_A_1102_93#_c_741_n N_A_1188_93#_c_897_n 0.0028942f $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_619 N_A_1102_93#_c_741_n CLK 0.0203377f $X=7.09 $Y=1.65 $X2=0 $Y2=0
cc_620 N_A_1102_93#_c_757_n CLK 0.00607042f $X=7.35 $Y=2.11 $X2=0 $Y2=0
cc_621 N_A_1102_93#_c_743_n CLK 0.0260483f $X=7.63 $Y=0.805 $X2=0 $Y2=0
cc_622 N_A_1102_93#_c_744_n CLK 0.00407799f $X=7.23 $Y=0.35 $X2=0 $Y2=0
cc_623 N_A_1102_93#_c_735_n N_CLK_c_1034_n 0.0104164f $X=9.89 $Y=0.18 $X2=0
+ $Y2=0
cc_624 N_A_1102_93#_c_737_n N_A_2122_329#_M1000_g 0.00969975f $X=11.885 $Y=0.18
+ $X2=0 $Y2=0
cc_625 N_A_1102_93#_M1034_g N_A_2122_329#_M1036_g 0.0394756f $X=10.505 $Y=2.525
+ $X2=0 $Y2=0
cc_626 N_A_1102_93#_c_751_n N_A_2122_329#_M1036_g 0.0103107f $X=11.885 $Y=3.15
+ $X2=0 $Y2=0
cc_627 N_A_1102_93#_c_737_n N_A_2122_329#_M1002_g 0.0132414f $X=11.885 $Y=0.18
+ $X2=0 $Y2=0
cc_628 N_A_1102_93#_c_738_n N_A_2122_329#_M1022_g 0.0328052f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_629 N_A_1102_93#_c_738_n N_A_2122_329#_c_1079_n 0.0132414f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_630 N_A_1102_93#_c_738_n N_A_2122_329#_c_1107_n 0.0117989f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_631 N_A_1102_93#_c_738_n N_A_2122_329#_c_1081_n 0.0133704f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_632 N_A_1102_93#_c_738_n N_A_2122_329#_c_1094_n 0.0104965f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_633 N_A_1102_93#_c_751_n N_A_2122_329#_c_1095_n 0.00477364f $X=11.885 $Y=3.15
+ $X2=0 $Y2=0
cc_634 N_A_1102_93#_c_738_n N_A_2122_329#_c_1095_n 0.011358f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_635 N_A_1102_93#_c_737_n N_A_2122_329#_c_1085_n 0.00506133f $X=11.885 $Y=0.18
+ $X2=0 $Y2=0
cc_636 N_A_1102_93#_c_738_n N_A_2122_329#_c_1085_n 0.0193035f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_637 N_A_1102_93#_c_738_n N_A_2122_329#_c_1100_n 0.00484778f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_638 N_A_1102_93#_c_751_n N_A_2008_122#_M1025_g 0.0103107f $X=11.885 $Y=3.15
+ $X2=0 $Y2=0
cc_639 N_A_1102_93#_c_738_n N_A_2008_122#_M1025_g 0.0247514f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_640 N_A_1102_93#_M1021_g N_A_2008_122#_c_1229_n 0.00114485f $X=9.965 $Y=0.82
+ $X2=0 $Y2=0
cc_641 N_A_1102_93#_c_737_n N_A_2008_122#_c_1229_n 0.00362644f $X=11.885 $Y=0.18
+ $X2=0 $Y2=0
cc_642 N_A_1102_93#_M1034_g N_A_2008_122#_c_1230_n 0.00805091f $X=10.505
+ $Y=2.525 $X2=0 $Y2=0
cc_643 N_A_1102_93#_c_738_n N_A_2008_122#_c_1231_n 2.20581e-19 $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_644 N_A_1102_93#_M1034_g N_A_2008_122#_c_1233_n 0.00384891f $X=10.505
+ $Y=2.525 $X2=0 $Y2=0
cc_645 N_A_1102_93#_c_737_n N_A_2008_122#_c_1234_n 0.0095796f $X=11.885 $Y=0.18
+ $X2=0 $Y2=0
cc_646 N_A_1102_93#_c_738_n N_A_2008_122#_c_1234_n 0.0300342f $X=11.96 $Y=3.075
+ $X2=0 $Y2=0
cc_647 N_A_1102_93#_M1034_g N_VPWR_c_1399_n 0.00896412f $X=10.505 $Y=2.525 $X2=0
+ $Y2=0
cc_648 N_A_1102_93#_c_751_n N_VPWR_c_1399_n 0.0333866f $X=11.885 $Y=3.15 $X2=0
+ $Y2=0
cc_649 N_A_1102_93#_c_738_n N_VPWR_c_1399_n 0.00424859f $X=11.96 $Y=3.075 $X2=0
+ $Y2=0
cc_650 N_A_1102_93#_c_751_n N_VPWR_c_1400_n 0.0193276f $X=11.885 $Y=3.15 $X2=0
+ $Y2=0
cc_651 N_A_1102_93#_c_738_n N_VPWR_c_1401_n 0.0122976f $X=11.96 $Y=3.075 $X2=0
+ $Y2=0
cc_652 N_A_1102_93#_M1039_g N_VPWR_c_1411_n 9.15902e-19 $X=6.065 $Y=2.715 $X2=0
+ $Y2=0
cc_653 N_A_1102_93#_c_752_n N_VPWR_c_1412_n 0.0179753f $X=10.58 $Y=3.15 $X2=0
+ $Y2=0
cc_654 N_A_1102_93#_c_751_n N_VPWR_c_1394_n 0.0364792f $X=11.885 $Y=3.15 $X2=0
+ $Y2=0
cc_655 N_A_1102_93#_c_752_n N_VPWR_c_1394_n 0.0116041f $X=10.58 $Y=3.15 $X2=0
+ $Y2=0
cc_656 N_A_1102_93#_M1017_g N_A_182_120#_c_1566_n 0.0152439f $X=5.585 $Y=0.805
+ $X2=0 $Y2=0
cc_657 N_A_1102_93#_c_733_n N_A_182_120#_c_1566_n 0.00770445f $X=5.99 $Y=1.59
+ $X2=0 $Y2=0
cc_658 N_A_1102_93#_c_739_n N_A_182_120#_c_1566_n 0.00203258f $X=6.065 $Y=1.59
+ $X2=0 $Y2=0
cc_659 N_A_1102_93#_c_741_n N_A_182_120#_c_1566_n 0.00543855f $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_660 N_A_1102_93#_c_742_n N_A_182_120#_c_1566_n 3.55289e-19 $X=7.09 $Y=1.65
+ $X2=0 $Y2=0
cc_661 N_A_1102_93#_M1017_g N_A_182_120#_c_1568_n 0.00230997f $X=5.585 $Y=0.805
+ $X2=0 $Y2=0
cc_662 N_A_1102_93#_c_744_n N_A_182_120#_c_1568_n 0.0130718f $X=7.23 $Y=0.35
+ $X2=0 $Y2=0
cc_663 N_A_1102_93#_M1039_g N_A_182_120#_c_1577_n 0.00266623f $X=6.065 $Y=2.715
+ $X2=0 $Y2=0
cc_664 N_A_1102_93#_M1039_g N_A_993_425#_c_1724_n 0.0143033f $X=6.065 $Y=2.715
+ $X2=0 $Y2=0
cc_665 N_A_1102_93#_c_738_n N_Q_c_1763_n 0.00314731f $X=11.96 $Y=3.075 $X2=0
+ $Y2=0
cc_666 N_A_1102_93#_c_738_n N_Q_c_1761_n 0.00158393f $X=11.96 $Y=3.075 $X2=0
+ $Y2=0
cc_667 N_A_1102_93#_c_738_n Q 0.00557573f $X=11.96 $Y=3.075 $X2=0 $Y2=0
cc_668 N_A_1102_93#_c_735_n N_VGND_c_1825_n 0.0215716f $X=9.89 $Y=0.18 $X2=0
+ $Y2=0
cc_669 N_A_1102_93#_c_744_n N_VGND_c_1825_n 0.0124622f $X=7.23 $Y=0.35 $X2=0
+ $Y2=0
cc_670 N_A_1102_93#_c_746_n N_VGND_c_1825_n 0.00376268f $X=7.23 $Y=0.18 $X2=0
+ $Y2=0
cc_671 N_A_1102_93#_c_737_n N_VGND_c_1826_n 0.0261591f $X=11.885 $Y=0.18 $X2=0
+ $Y2=0
cc_672 N_A_1102_93#_c_738_n N_VGND_c_1826_n 0.00360908f $X=11.96 $Y=3.075 $X2=0
+ $Y2=0
cc_673 N_A_1102_93#_c_737_n N_VGND_c_1827_n 0.0156886f $X=11.885 $Y=0.18 $X2=0
+ $Y2=0
cc_674 N_A_1102_93#_c_743_n N_VGND_c_1836_n 0.00629135f $X=7.63 $Y=0.805 $X2=0
+ $Y2=0
cc_675 N_A_1102_93#_c_744_n N_VGND_c_1836_n 0.02743f $X=7.23 $Y=0.35 $X2=0 $Y2=0
cc_676 N_A_1102_93#_c_746_n N_VGND_c_1836_n 0.0227136f $X=7.23 $Y=0.18 $X2=0
+ $Y2=0
cc_677 N_A_1102_93#_c_735_n N_VGND_c_1838_n 0.08763f $X=9.89 $Y=0.18 $X2=0 $Y2=0
cc_678 N_A_1102_93#_c_737_n N_VGND_c_1840_n 0.0207279f $X=11.885 $Y=0.18 $X2=0
+ $Y2=0
cc_679 N_A_1102_93#_M1017_g N_VGND_c_1847_n 7.85159e-19 $X=5.585 $Y=0.805 $X2=0
+ $Y2=0
cc_680 N_A_1102_93#_c_735_n N_VGND_c_1847_n 0.0791327f $X=9.89 $Y=0.18 $X2=0
+ $Y2=0
cc_681 N_A_1102_93#_c_737_n N_VGND_c_1847_n 0.0637807f $X=11.885 $Y=0.18 $X2=0
+ $Y2=0
cc_682 N_A_1102_93#_c_740_n N_VGND_c_1847_n 0.00926736f $X=9.965 $Y=0.18 $X2=0
+ $Y2=0
cc_683 N_A_1102_93#_c_743_n N_VGND_c_1847_n 0.00921962f $X=7.63 $Y=0.805 $X2=0
+ $Y2=0
cc_684 N_A_1102_93#_c_744_n N_VGND_c_1847_n 0.0139792f $X=7.23 $Y=0.35 $X2=0
+ $Y2=0
cc_685 N_A_1102_93#_c_746_n N_VGND_c_1847_n 0.00855357f $X=7.23 $Y=0.18 $X2=0
+ $Y2=0
cc_686 N_A_1188_93#_c_899_n N_CLK_M1001_g 0.00686043f $X=8.705 $Y=3.11 $X2=0
+ $Y2=0
cc_687 N_A_1188_93#_M1027_g N_CLK_M1001_g 0.0260609f $X=7.68 $Y=2.295 $X2=0
+ $Y2=0
cc_688 N_A_1188_93#_c_891_n N_CLK_M1001_g 0.00981289f $X=8.32 $Y=1.667 $X2=0
+ $Y2=0
cc_689 N_A_1188_93#_c_892_n N_CLK_M1001_g 0.016098f $X=7.755 $Y=1.65 $X2=0 $Y2=0
cc_690 N_A_1188_93#_c_893_n N_CLK_M1001_g 0.0036734f $X=8.485 $Y=1.77 $X2=0
+ $Y2=0
cc_691 N_A_1188_93#_c_907_n N_CLK_M1001_g 0.0114805f $X=8.485 $Y=2.11 $X2=0
+ $Y2=0
cc_692 N_A_1188_93#_c_895_n N_CLK_M1001_g 5.9691e-19 $X=8.89 $Y=1.23 $X2=0 $Y2=0
cc_693 N_A_1188_93#_c_896_n N_CLK_M1001_g 0.0374234f $X=8.89 $Y=1.23 $X2=0 $Y2=0
cc_694 N_A_1188_93#_c_897_n N_CLK_M1001_g 7.84456e-19 $X=7.755 $Y=1.485 $X2=0
+ $Y2=0
cc_695 N_A_1188_93#_c_881_n CLK 0.0103638f $X=7.59 $Y=1.2 $X2=0 $Y2=0
cc_696 N_A_1188_93#_c_889_n CLK 0.0152204f $X=7.845 $Y=1.2 $X2=0 $Y2=0
cc_697 N_A_1188_93#_c_891_n CLK 0.0544816f $X=8.32 $Y=1.667 $X2=0 $Y2=0
cc_698 N_A_1188_93#_c_892_n CLK 0.0011723f $X=7.755 $Y=1.65 $X2=0 $Y2=0
cc_699 N_A_1188_93#_c_893_n CLK 0.0190654f $X=8.485 $Y=1.77 $X2=0 $Y2=0
cc_700 N_A_1188_93#_c_894_n CLK 0.013187f $X=8.72 $Y=0.805 $X2=0 $Y2=0
cc_701 N_A_1188_93#_c_895_n CLK 0.0213358f $X=8.89 $Y=1.23 $X2=0 $Y2=0
cc_702 N_A_1188_93#_c_896_n CLK 0.00164146f $X=8.89 $Y=1.23 $X2=0 $Y2=0
cc_703 N_A_1188_93#_c_897_n CLK 0.00788886f $X=7.755 $Y=1.485 $X2=0 $Y2=0
cc_704 N_A_1188_93#_c_889_n N_CLK_c_1033_n 0.00816939f $X=7.845 $Y=1.2 $X2=0
+ $Y2=0
cc_705 N_A_1188_93#_c_891_n N_CLK_c_1033_n 8.51192e-19 $X=8.32 $Y=1.667 $X2=0
+ $Y2=0
cc_706 N_A_1188_93#_c_893_n N_CLK_c_1033_n 0.00366103f $X=8.485 $Y=1.77 $X2=0
+ $Y2=0
cc_707 N_A_1188_93#_c_894_n N_CLK_c_1033_n 0.00307892f $X=8.72 $Y=0.805 $X2=0
+ $Y2=0
cc_708 N_A_1188_93#_c_895_n N_CLK_c_1033_n 8.00949e-19 $X=8.89 $Y=1.23 $X2=0
+ $Y2=0
cc_709 N_A_1188_93#_c_896_n N_CLK_c_1033_n 0.0208555f $X=8.89 $Y=1.23 $X2=0
+ $Y2=0
cc_710 N_A_1188_93#_c_897_n N_CLK_c_1033_n 0.00552291f $X=7.755 $Y=1.485 $X2=0
+ $Y2=0
cc_711 N_A_1188_93#_c_883_n N_CLK_c_1034_n 0.0116351f $X=7.845 $Y=1.125 $X2=0
+ $Y2=0
cc_712 N_A_1188_93#_c_895_n N_CLK_c_1034_n 0.00279514f $X=8.89 $Y=1.23 $X2=0
+ $Y2=0
cc_713 N_A_1188_93#_c_896_n N_CLK_c_1034_n 0.00243234f $X=8.89 $Y=1.23 $X2=0
+ $Y2=0
cc_714 N_A_1188_93#_M1011_g N_A_2122_329#_M1000_g 0.001518f $X=9.995 $Y=2.315
+ $X2=0 $Y2=0
cc_715 N_A_1188_93#_c_887_n N_A_2122_329#_M1000_g 0.0102332f $X=10.41 $Y=1.16
+ $X2=0 $Y2=0
cc_716 N_A_1188_93#_M1015_g N_A_2122_329#_M1000_g 0.0497971f $X=10.41 $Y=0.82
+ $X2=0 $Y2=0
cc_717 N_A_1188_93#_M1011_g N_A_2122_329#_c_1084_n 0.00482746f $X=9.995 $Y=2.315
+ $X2=0 $Y2=0
cc_718 N_A_1188_93#_c_886_n N_A_2008_122#_c_1229_n 0.00301292f $X=10.28 $Y=1.445
+ $X2=0 $Y2=0
cc_719 N_A_1188_93#_c_887_n N_A_2008_122#_c_1229_n 0.0102182f $X=10.41 $Y=1.16
+ $X2=0 $Y2=0
cc_720 N_A_1188_93#_M1015_g N_A_2008_122#_c_1229_n 0.01125f $X=10.41 $Y=0.82
+ $X2=0 $Y2=0
cc_721 N_A_1188_93#_c_890_n N_A_2008_122#_c_1229_n 6.98643e-19 $X=9.995 $Y=1.445
+ $X2=0 $Y2=0
cc_722 N_A_1188_93#_M1011_g N_A_2008_122#_c_1230_n 0.0214964f $X=9.995 $Y=2.315
+ $X2=0 $Y2=0
cc_723 N_A_1188_93#_M1011_g N_A_2008_122#_c_1241_n 8.83771e-19 $X=9.995 $Y=2.315
+ $X2=0 $Y2=0
cc_724 N_A_1188_93#_c_886_n N_A_2008_122#_c_1241_n 0.00784604f $X=10.28 $Y=1.445
+ $X2=0 $Y2=0
cc_725 N_A_1188_93#_c_887_n N_A_2008_122#_c_1241_n 0.00303989f $X=10.41 $Y=1.16
+ $X2=0 $Y2=0
cc_726 N_A_1188_93#_c_890_n N_A_2008_122#_c_1241_n 0.00235901f $X=9.995 $Y=1.445
+ $X2=0 $Y2=0
cc_727 N_A_1188_93#_c_887_n N_A_2008_122#_c_1233_n 0.00908551f $X=10.41 $Y=1.16
+ $X2=0 $Y2=0
cc_728 N_A_1188_93#_c_899_n N_VPWR_c_1398_n 0.0271602f $X=8.705 $Y=3.11 $X2=0
+ $Y2=0
cc_729 N_A_1188_93#_M1027_g N_VPWR_c_1398_n 0.00116328f $X=7.68 $Y=2.295 $X2=0
+ $Y2=0
cc_730 N_A_1188_93#_c_902_n N_VPWR_c_1398_n 0.00720029f $X=8.78 $Y=3.035 $X2=0
+ $Y2=0
cc_731 N_A_1188_93#_c_900_n N_VPWR_c_1411_n 0.0389329f $X=6.57 $Y=3.11 $X2=0
+ $Y2=0
cc_732 N_A_1188_93#_c_899_n N_VPWR_c_1412_n 0.0243183f $X=8.705 $Y=3.11 $X2=0
+ $Y2=0
cc_733 N_A_1188_93#_M1011_g N_VPWR_c_1412_n 0.00414853f $X=9.995 $Y=2.315 $X2=0
+ $Y2=0
cc_734 N_A_1188_93#_c_899_n N_VPWR_c_1394_n 0.056922f $X=8.705 $Y=3.11 $X2=0
+ $Y2=0
cc_735 N_A_1188_93#_c_900_n N_VPWR_c_1394_n 0.00542545f $X=6.57 $Y=3.11 $X2=0
+ $Y2=0
cc_736 N_A_1188_93#_M1027_g N_VPWR_c_1394_n 9.17629e-19 $X=7.68 $Y=2.295 $X2=0
+ $Y2=0
cc_737 N_A_1188_93#_M1011_g N_VPWR_c_1394_n 0.00477801f $X=9.995 $Y=2.315 $X2=0
+ $Y2=0
cc_738 N_A_1188_93#_c_882_n N_A_182_120#_c_1566_n 0.00369183f $X=6.09 $Y=1.2
+ $X2=0 $Y2=0
cc_739 N_A_1188_93#_c_880_n N_A_182_120#_c_1568_n 0.00487552f $X=6.015 $Y=1.125
+ $X2=0 $Y2=0
cc_740 N_A_1188_93#_c_881_n N_A_182_120#_c_1568_n 0.0152059f $X=7.59 $Y=1.2
+ $X2=0 $Y2=0
cc_741 N_A_1188_93#_c_898_n N_A_993_425#_c_1724_n 0.0108593f $X=6.495 $Y=3.035
+ $X2=0 $Y2=0
cc_742 N_A_1188_93#_c_899_n N_A_993_425#_c_1724_n 7.34723e-19 $X=8.705 $Y=3.11
+ $X2=0 $Y2=0
cc_743 N_A_1188_93#_c_900_n N_A_993_425#_c_1724_n 0.00241615f $X=6.57 $Y=3.11
+ $X2=0 $Y2=0
cc_744 N_A_1188_93#_c_898_n N_A_993_425#_c_1726_n 0.00114627f $X=6.495 $Y=3.035
+ $X2=0 $Y2=0
cc_745 N_A_1188_93#_c_899_n N_A_993_425#_c_1726_n 0.011811f $X=8.705 $Y=3.11
+ $X2=0 $Y2=0
cc_746 N_A_1188_93#_M1027_g N_A_993_425#_c_1726_n 9.03897e-19 $X=7.68 $Y=2.295
+ $X2=0 $Y2=0
cc_747 N_A_1188_93#_c_883_n N_VGND_c_1825_n 0.00181767f $X=7.845 $Y=1.125 $X2=0
+ $Y2=0
cc_748 N_A_1188_93#_c_894_n N_VGND_c_1838_n 0.012885f $X=8.72 $Y=0.805 $X2=0
+ $Y2=0
cc_749 N_A_1188_93#_c_883_n N_VGND_c_1847_n 9.39239e-19 $X=7.845 $Y=1.125 $X2=0
+ $Y2=0
cc_750 N_A_1188_93#_M1015_g N_VGND_c_1847_n 9.44905e-19 $X=10.41 $Y=0.82 $X2=0
+ $Y2=0
cc_751 N_A_1188_93#_c_894_n N_VGND_c_1847_n 0.0180329f $X=8.72 $Y=0.805 $X2=0
+ $Y2=0
cc_752 N_CLK_M1001_g N_VPWR_c_1398_n 0.00116328f $X=8.27 $Y=2.295 $X2=0 $Y2=0
cc_753 N_CLK_M1001_g N_VPWR_c_1394_n 9.17629e-19 $X=8.27 $Y=2.295 $X2=0 $Y2=0
cc_754 CLK N_VGND_c_1825_n 0.0173467f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_755 N_CLK_c_1034_n N_VGND_c_1825_n 0.003537f $X=8.325 $Y=1.13 $X2=0 $Y2=0
cc_756 N_CLK_c_1034_n N_VGND_c_1847_n 9.39239e-19 $X=8.325 $Y=1.13 $X2=0 $Y2=0
cc_757 N_A_2122_329#_c_1092_n N_A_2008_122#_M1025_g 0.0148681f $X=11.56 $Y=1.885
+ $X2=0 $Y2=0
cc_758 N_A_2122_329#_c_1081_n N_A_2008_122#_M1025_g 0.00114947f $X=11.815
+ $Y=1.795 $X2=0 $Y2=0
cc_759 N_A_2122_329#_c_1095_n N_A_2008_122#_M1025_g 2.83774e-19 $X=11.94 $Y=2.46
+ $X2=0 $Y2=0
cc_760 N_A_2122_329#_c_1084_n N_A_2008_122#_M1025_g 0.0208448f $X=10.775 $Y=1.81
+ $X2=0 $Y2=0
cc_761 N_A_2122_329#_c_1099_n N_A_2008_122#_M1025_g 4.18325e-19 $X=10.94
+ $Y=1.847 $X2=0 $Y2=0
cc_762 N_A_2122_329#_M1000_g N_A_2008_122#_c_1229_n 0.00253055f $X=10.77 $Y=0.82
+ $X2=0 $Y2=0
cc_763 N_A_2122_329#_M1000_g N_A_2008_122#_c_1230_n 0.00203558f $X=10.77 $Y=0.82
+ $X2=0 $Y2=0
cc_764 N_A_2122_329#_M1036_g N_A_2008_122#_c_1230_n 0.004671f $X=10.865 $Y=2.525
+ $X2=0 $Y2=0
cc_765 N_A_2122_329#_c_1084_n N_A_2008_122#_c_1230_n 0.00294559f $X=10.775
+ $Y=1.81 $X2=0 $Y2=0
cc_766 N_A_2122_329#_c_1099_n N_A_2008_122#_c_1230_n 0.0155933f $X=10.94
+ $Y=1.847 $X2=0 $Y2=0
cc_767 N_A_2122_329#_M1000_g N_A_2008_122#_c_1231_n 4.45865e-19 $X=10.77 $Y=0.82
+ $X2=0 $Y2=0
cc_768 N_A_2122_329#_c_1092_n N_A_2008_122#_c_1231_n 0.0238093f $X=11.56
+ $Y=1.885 $X2=0 $Y2=0
cc_769 N_A_2122_329#_c_1081_n N_A_2008_122#_c_1231_n 0.0188139f $X=11.815
+ $Y=1.795 $X2=0 $Y2=0
cc_770 N_A_2122_329#_M1000_g N_A_2008_122#_c_1232_n 0.0102005f $X=10.77 $Y=0.82
+ $X2=0 $Y2=0
cc_771 N_A_2122_329#_c_1092_n N_A_2008_122#_c_1232_n 0.00558536f $X=11.56
+ $Y=1.885 $X2=0 $Y2=0
cc_772 N_A_2122_329#_c_1084_n N_A_2008_122#_c_1232_n 0.00331559f $X=10.775
+ $Y=1.81 $X2=0 $Y2=0
cc_773 N_A_2122_329#_M1000_g N_A_2008_122#_c_1233_n 0.0154418f $X=10.77 $Y=0.82
+ $X2=0 $Y2=0
cc_774 N_A_2122_329#_c_1092_n N_A_2008_122#_c_1233_n 0.0140105f $X=11.56
+ $Y=1.885 $X2=0 $Y2=0
cc_775 N_A_2122_329#_c_1084_n N_A_2008_122#_c_1233_n 0.00481612f $X=10.775
+ $Y=1.81 $X2=0 $Y2=0
cc_776 N_A_2122_329#_c_1099_n N_A_2008_122#_c_1233_n 0.0237591f $X=10.94
+ $Y=1.847 $X2=0 $Y2=0
cc_777 N_A_2122_329#_M1000_g N_A_2008_122#_c_1234_n 0.013378f $X=10.77 $Y=0.82
+ $X2=0 $Y2=0
cc_778 N_A_2122_329#_c_1081_n N_A_2008_122#_c_1234_n 0.00649599f $X=11.815
+ $Y=1.795 $X2=0 $Y2=0
cc_779 N_A_2122_329#_c_1085_n N_A_2008_122#_c_1234_n 0.00776842f $X=11.685
+ $Y=0.755 $X2=0 $Y2=0
cc_780 N_A_2122_329#_c_1083_n N_A_2710_56#_M1008_g 0.00254964f $X=13.69 $Y=1.49
+ $X2=0 $Y2=0
cc_781 N_A_2122_329#_M1037_g N_A_2710_56#_c_1306_n 2.14085e-19 $X=12.97 $Y=2.465
+ $X2=0 $Y2=0
cc_782 N_A_2122_329#_M1007_g N_A_2710_56#_c_1306_n 0.00733239f $X=13.495
+ $Y=2.155 $X2=0 $Y2=0
cc_783 N_A_2122_329#_c_1094_n N_A_2710_56#_c_1306_n 0.0073373f $X=13.15 $Y=2.46
+ $X2=0 $Y2=0
cc_784 N_A_2122_329#_c_1096_n N_A_2710_56#_c_1306_n 0.0267496f $X=13.235
+ $Y=2.375 $X2=0 $Y2=0
cc_785 N_A_2122_329#_M1029_g N_A_2710_56#_c_1300_n 0.00873812f $X=13.475 $Y=0.49
+ $X2=0 $Y2=0
cc_786 N_A_2122_329#_M1029_g N_A_2710_56#_c_1301_n 0.00573962f $X=13.475 $Y=0.49
+ $X2=0 $Y2=0
cc_787 N_A_2122_329#_c_1082_n N_A_2710_56#_c_1301_n 0.020639f $X=13.69 $Y=1.49
+ $X2=0 $Y2=0
cc_788 N_A_2122_329#_c_1083_n N_A_2710_56#_c_1301_n 0.00741084f $X=13.69 $Y=1.49
+ $X2=0 $Y2=0
cc_789 N_A_2122_329#_M1007_g N_A_2710_56#_c_1307_n 0.00425038f $X=13.495
+ $Y=2.155 $X2=0 $Y2=0
cc_790 N_A_2122_329#_c_1096_n N_A_2710_56#_c_1307_n 0.0107352f $X=13.235
+ $Y=2.375 $X2=0 $Y2=0
cc_791 N_A_2122_329#_c_1082_n N_A_2710_56#_c_1307_n 0.0221699f $X=13.69 $Y=1.49
+ $X2=0 $Y2=0
cc_792 N_A_2122_329#_c_1083_n N_A_2710_56#_c_1307_n 0.00694095f $X=13.69 $Y=1.49
+ $X2=0 $Y2=0
cc_793 N_A_2122_329#_M1029_g N_A_2710_56#_c_1302_n 0.00184291f $X=13.475 $Y=0.49
+ $X2=0 $Y2=0
cc_794 N_A_2122_329#_M1007_g N_A_2710_56#_c_1302_n 0.00275553f $X=13.495
+ $Y=2.155 $X2=0 $Y2=0
cc_795 N_A_2122_329#_c_1082_n N_A_2710_56#_c_1302_n 0.0150034f $X=13.69 $Y=1.49
+ $X2=0 $Y2=0
cc_796 N_A_2122_329#_c_1083_n N_A_2710_56#_c_1302_n 0.0047257f $X=13.69 $Y=1.49
+ $X2=0 $Y2=0
cc_797 N_A_2122_329#_M1029_g N_A_2710_56#_c_1303_n 0.00203187f $X=13.475 $Y=0.49
+ $X2=0 $Y2=0
cc_798 N_A_2122_329#_c_1083_n N_A_2710_56#_c_1303_n 0.00911314f $X=13.69 $Y=1.49
+ $X2=0 $Y2=0
cc_799 N_A_2122_329#_c_1092_n N_VPWR_M1036_d 0.00249921f $X=11.56 $Y=1.885 $X2=0
+ $Y2=0
cc_800 N_A_2122_329#_c_1094_n N_VPWR_M1022_d 0.00502406f $X=13.15 $Y=2.46 $X2=0
+ $Y2=0
cc_801 N_A_2122_329#_c_1094_n N_VPWR_M1037_d 0.00582007f $X=13.15 $Y=2.46 $X2=0
+ $Y2=0
cc_802 N_A_2122_329#_c_1096_n N_VPWR_M1037_d 0.0145898f $X=13.235 $Y=2.375 $X2=0
+ $Y2=0
cc_803 N_A_2122_329#_M1036_g N_VPWR_c_1399_n 0.019363f $X=10.865 $Y=2.525 $X2=0
+ $Y2=0
cc_804 N_A_2122_329#_c_1095_n N_VPWR_c_1399_n 0.0159585f $X=11.94 $Y=2.46 $X2=0
+ $Y2=0
cc_805 N_A_2122_329#_c_1099_n N_VPWR_c_1399_n 0.0341903f $X=10.94 $Y=1.847 $X2=0
+ $Y2=0
cc_806 N_A_2122_329#_c_1095_n N_VPWR_c_1400_n 0.00862229f $X=11.94 $Y=2.46 $X2=0
+ $Y2=0
cc_807 N_A_2122_329#_M1022_g N_VPWR_c_1401_n 0.0118978f $X=12.54 $Y=2.465 $X2=0
+ $Y2=0
cc_808 N_A_2122_329#_M1037_g N_VPWR_c_1401_n 0.00154589f $X=12.97 $Y=2.465 $X2=0
+ $Y2=0
cc_809 N_A_2122_329#_c_1094_n N_VPWR_c_1401_n 0.0214609f $X=13.15 $Y=2.46 $X2=0
+ $Y2=0
cc_810 N_A_2122_329#_c_1095_n N_VPWR_c_1401_n 0.00264707f $X=11.94 $Y=2.46 $X2=0
+ $Y2=0
cc_811 N_A_2122_329#_M1022_g N_VPWR_c_1402_n 0.00154589f $X=12.54 $Y=2.465 $X2=0
+ $Y2=0
cc_812 N_A_2122_329#_M1037_g N_VPWR_c_1402_n 0.0133042f $X=12.97 $Y=2.465 $X2=0
+ $Y2=0
cc_813 N_A_2122_329#_c_1094_n N_VPWR_c_1402_n 0.0204136f $X=13.15 $Y=2.46 $X2=0
+ $Y2=0
cc_814 N_A_2122_329#_M1007_g N_VPWR_c_1403_n 0.00312414f $X=13.495 $Y=2.155
+ $X2=0 $Y2=0
cc_815 N_A_2122_329#_M1007_g N_VPWR_c_1404_n 0.0034616f $X=13.495 $Y=2.155 $X2=0
+ $Y2=0
cc_816 N_A_2122_329#_M1022_g N_VPWR_c_1413_n 0.00486043f $X=12.54 $Y=2.465 $X2=0
+ $Y2=0
cc_817 N_A_2122_329#_M1037_g N_VPWR_c_1413_n 0.00486043f $X=12.97 $Y=2.465 $X2=0
+ $Y2=0
cc_818 N_A_2122_329#_M1036_g N_VPWR_c_1394_n 7.88961e-19 $X=10.865 $Y=2.525
+ $X2=0 $Y2=0
cc_819 N_A_2122_329#_M1022_g N_VPWR_c_1394_n 0.0045039f $X=12.54 $Y=2.465 $X2=0
+ $Y2=0
cc_820 N_A_2122_329#_M1037_g N_VPWR_c_1394_n 0.0045039f $X=12.97 $Y=2.465 $X2=0
+ $Y2=0
cc_821 N_A_2122_329#_M1007_g N_VPWR_c_1394_n 0.00410284f $X=13.495 $Y=2.155
+ $X2=0 $Y2=0
cc_822 N_A_2122_329#_c_1094_n N_VPWR_c_1394_n 0.0270287f $X=13.15 $Y=2.46 $X2=0
+ $Y2=0
cc_823 N_A_2122_329#_c_1095_n N_VPWR_c_1394_n 0.0104591f $X=11.94 $Y=2.46 $X2=0
+ $Y2=0
cc_824 N_A_2122_329#_c_1094_n N_Q_M1022_s 0.00494804f $X=13.15 $Y=2.46 $X2=0
+ $Y2=0
cc_825 N_A_2122_329#_M1002_g N_Q_c_1759_n 0.0142864f $X=12.52 $Y=0.7 $X2=0 $Y2=0
cc_826 N_A_2122_329#_M1019_g N_Q_c_1759_n 0.00286881f $X=12.95 $Y=0.7 $X2=0
+ $Y2=0
cc_827 N_A_2122_329#_c_1079_n N_Q_c_1759_n 0.00263351f $X=13.045 $Y=1.49 $X2=0
+ $Y2=0
cc_828 N_A_2122_329#_c_1190_p N_Q_c_1759_n 0.026813f $X=13.15 $Y=1.53 $X2=0
+ $Y2=0
cc_829 N_A_2122_329#_c_1107_n N_Q_c_1763_n 0.0195449f $X=11.655 $Y=2.04 $X2=0
+ $Y2=0
cc_830 N_A_2122_329#_c_1094_n N_Q_c_1763_n 0.0184933f $X=13.15 $Y=2.46 $X2=0
+ $Y2=0
cc_831 N_A_2122_329#_c_1100_n N_Q_c_1763_n 0.00891438f $X=11.75 $Y=1.885 $X2=0
+ $Y2=0
cc_832 N_A_2122_329#_M1022_g N_Q_c_1776_n 0.0143807f $X=12.54 $Y=2.465 $X2=0
+ $Y2=0
cc_833 N_A_2122_329#_M1037_g N_Q_c_1776_n 0.00468491f $X=12.97 $Y=2.465 $X2=0
+ $Y2=0
cc_834 N_A_2122_329#_c_1079_n N_Q_c_1776_n 0.00228492f $X=13.045 $Y=1.49 $X2=0
+ $Y2=0
cc_835 N_A_2122_329#_c_1094_n N_Q_c_1776_n 0.0306469f $X=13.15 $Y=2.46 $X2=0
+ $Y2=0
cc_836 N_A_2122_329#_c_1190_p N_Q_c_1776_n 0.0217673f $X=13.15 $Y=1.53 $X2=0
+ $Y2=0
cc_837 N_A_2122_329#_c_1096_n N_Q_c_1776_n 0.0203954f $X=13.235 $Y=2.375 $X2=0
+ $Y2=0
cc_838 N_A_2122_329#_M1002_g N_Q_c_1760_n 9.17203e-19 $X=12.52 $Y=0.7 $X2=0
+ $Y2=0
cc_839 N_A_2122_329#_M1019_g N_Q_c_1760_n 9.97884e-19 $X=12.95 $Y=0.7 $X2=0
+ $Y2=0
cc_840 N_A_2122_329#_c_1085_n N_Q_c_1761_n 0.0145637f $X=11.685 $Y=0.755 $X2=0
+ $Y2=0
cc_841 N_A_2122_329#_M1002_g Q 0.00733655f $X=12.52 $Y=0.7 $X2=0 $Y2=0
cc_842 N_A_2122_329#_M1022_g Q 0.00537683f $X=12.54 $Y=2.465 $X2=0 $Y2=0
cc_843 N_A_2122_329#_c_1081_n Q 0.0437081f $X=11.815 $Y=1.795 $X2=0 $Y2=0
cc_844 N_A_2122_329#_c_1190_p Q 0.0202253f $X=13.15 $Y=1.53 $X2=0 $Y2=0
cc_845 N_A_2122_329#_c_1100_n Q 0.00648463f $X=11.75 $Y=1.885 $X2=0 $Y2=0
cc_846 N_A_2122_329#_M1000_g N_VGND_c_1826_n 0.0125252f $X=10.77 $Y=0.82 $X2=0
+ $Y2=0
cc_847 N_A_2122_329#_c_1085_n N_VGND_c_1826_n 0.0238161f $X=11.685 $Y=0.755
+ $X2=0 $Y2=0
cc_848 N_A_2122_329#_M1002_g N_VGND_c_1827_n 0.0103266f $X=12.52 $Y=0.7 $X2=0
+ $Y2=0
cc_849 N_A_2122_329#_M1019_g N_VGND_c_1827_n 5.40855e-19 $X=12.95 $Y=0.7 $X2=0
+ $Y2=0
cc_850 N_A_2122_329#_c_1085_n N_VGND_c_1827_n 0.0206762f $X=11.685 $Y=0.755
+ $X2=0 $Y2=0
cc_851 N_A_2122_329#_M1019_g N_VGND_c_1828_n 0.00480481f $X=12.95 $Y=0.7 $X2=0
+ $Y2=0
cc_852 N_A_2122_329#_c_1078_n N_VGND_c_1828_n 0.00482585f $X=13.4 $Y=1.49 $X2=0
+ $Y2=0
cc_853 N_A_2122_329#_M1029_g N_VGND_c_1828_n 0.00656819f $X=13.475 $Y=0.49 $X2=0
+ $Y2=0
cc_854 N_A_2122_329#_c_1190_p N_VGND_c_1828_n 0.00643401f $X=13.15 $Y=1.53 $X2=0
+ $Y2=0
cc_855 N_A_2122_329#_c_1082_n N_VGND_c_1828_n 0.00370459f $X=13.69 $Y=1.49 $X2=0
+ $Y2=0
cc_856 N_A_2122_329#_c_1218_p N_VGND_c_1828_n 0.0108532f $X=13.235 $Y=1.53 $X2=0
+ $Y2=0
cc_857 N_A_2122_329#_M1029_g N_VGND_c_1829_n 0.00282693f $X=13.475 $Y=0.49 $X2=0
+ $Y2=0
cc_858 N_A_2122_329#_c_1085_n N_VGND_c_1840_n 0.00910089f $X=11.685 $Y=0.755
+ $X2=0 $Y2=0
cc_859 N_A_2122_329#_M1002_g N_VGND_c_1841_n 0.00448994f $X=12.52 $Y=0.7 $X2=0
+ $Y2=0
cc_860 N_A_2122_329#_M1019_g N_VGND_c_1841_n 0.00540763f $X=12.95 $Y=0.7 $X2=0
+ $Y2=0
cc_861 N_A_2122_329#_M1029_g N_VGND_c_1842_n 0.00540763f $X=13.475 $Y=0.49 $X2=0
+ $Y2=0
cc_862 N_A_2122_329#_M1000_g N_VGND_c_1847_n 9.44906e-19 $X=10.77 $Y=0.82 $X2=0
+ $Y2=0
cc_863 N_A_2122_329#_M1002_g N_VGND_c_1847_n 0.00812427f $X=12.52 $Y=0.7 $X2=0
+ $Y2=0
cc_864 N_A_2122_329#_M1019_g N_VGND_c_1847_n 0.0104197f $X=12.95 $Y=0.7 $X2=0
+ $Y2=0
cc_865 N_A_2122_329#_M1029_g N_VGND_c_1847_n 0.0113695f $X=13.475 $Y=0.49 $X2=0
+ $Y2=0
cc_866 N_A_2122_329#_c_1085_n N_VGND_c_1847_n 0.0113231f $X=11.685 $Y=0.755
+ $X2=0 $Y2=0
cc_867 N_A_2008_122#_M1025_g N_VPWR_c_1399_n 0.0160836f $X=11.44 $Y=2.315 $X2=0
+ $Y2=0
cc_868 N_A_2008_122#_c_1230_n N_VPWR_c_1399_n 0.0201144f $X=10.21 $Y=2.02 $X2=0
+ $Y2=0
cc_869 N_A_2008_122#_c_1230_n N_VPWR_c_1412_n 0.00749997f $X=10.21 $Y=2.02 $X2=0
+ $Y2=0
cc_870 N_A_2008_122#_M1025_g N_VPWR_c_1394_n 7.88961e-19 $X=11.44 $Y=2.315 $X2=0
+ $Y2=0
cc_871 N_A_2008_122#_c_1230_n N_VPWR_c_1394_n 0.0100422f $X=10.21 $Y=2.02 $X2=0
+ $Y2=0
cc_872 N_A_2008_122#_c_1229_n N_VGND_c_1826_n 0.0149388f $X=10.195 $Y=0.825
+ $X2=0 $Y2=0
cc_873 N_A_2008_122#_c_1232_n N_VGND_c_1826_n 0.00376832f $X=11.345 $Y=1.53
+ $X2=0 $Y2=0
cc_874 N_A_2008_122#_c_1233_n N_VGND_c_1826_n 0.0268237f $X=11.18 $Y=1.502 $X2=0
+ $Y2=0
cc_875 N_A_2008_122#_c_1234_n N_VGND_c_1826_n 0.00797736f $X=11.362 $Y=1.365
+ $X2=0 $Y2=0
cc_876 N_A_2008_122#_c_1229_n N_VGND_c_1838_n 0.00469744f $X=10.195 $Y=0.825
+ $X2=0 $Y2=0
cc_877 N_A_2008_122#_c_1229_n N_VGND_c_1847_n 0.0080553f $X=10.195 $Y=0.825
+ $X2=0 $Y2=0
cc_878 N_A_2008_122#_c_1234_n N_VGND_c_1847_n 9.44905e-19 $X=11.362 $Y=1.365
+ $X2=0 $Y2=0
cc_879 N_A_2710_56#_c_1307_n N_VPWR_M1008_d 0.0032561f $X=14.2 $Y=1.755 $X2=0
+ $Y2=0
cc_880 N_A_2710_56#_M1008_g N_VPWR_c_1404_n 0.00328509f $X=14.445 $Y=2.465 $X2=0
+ $Y2=0
cc_881 N_A_2710_56#_c_1306_n N_VPWR_c_1404_n 0.0228131f $X=13.71 $Y=1.98 $X2=0
+ $Y2=0
cc_882 N_A_2710_56#_c_1307_n N_VPWR_c_1404_n 0.0145773f $X=14.2 $Y=1.755 $X2=0
+ $Y2=0
cc_883 N_A_2710_56#_M1028_g N_VPWR_c_1406_n 0.00749233f $X=14.875 $Y=2.465 $X2=0
+ $Y2=0
cc_884 N_A_2710_56#_M1008_g N_VPWR_c_1414_n 0.00585385f $X=14.445 $Y=2.465 $X2=0
+ $Y2=0
cc_885 N_A_2710_56#_M1028_g N_VPWR_c_1414_n 0.00564131f $X=14.875 $Y=2.465 $X2=0
+ $Y2=0
cc_886 N_A_2710_56#_M1008_g N_VPWR_c_1394_n 0.0118904f $X=14.445 $Y=2.465 $X2=0
+ $Y2=0
cc_887 N_A_2710_56#_M1028_g N_VPWR_c_1394_n 0.0110509f $X=14.875 $Y=2.465 $X2=0
+ $Y2=0
cc_888 N_A_2710_56#_c_1306_n N_VPWR_c_1394_n 0.0125384f $X=13.71 $Y=1.98 $X2=0
+ $Y2=0
cc_889 N_A_2710_56#_c_1296_n N_Q_N_c_1803_n 0.00145784f $X=14.445 $Y=1.185 $X2=0
+ $Y2=0
cc_890 N_A_2710_56#_M1008_g N_Q_N_c_1803_n 0.0029963f $X=14.445 $Y=2.465 $X2=0
+ $Y2=0
cc_891 N_A_2710_56#_c_1298_n N_Q_N_c_1803_n 0.0146858f $X=14.875 $Y=1.185 $X2=0
+ $Y2=0
cc_892 N_A_2710_56#_M1028_g N_Q_N_c_1803_n 0.0291599f $X=14.875 $Y=2.465 $X2=0
+ $Y2=0
cc_893 N_A_2710_56#_c_1301_n N_Q_N_c_1803_n 0.012289f $X=14.2 $Y=1.225 $X2=0
+ $Y2=0
cc_894 N_A_2710_56#_c_1307_n N_Q_N_c_1803_n 0.00977603f $X=14.2 $Y=1.755 $X2=0
+ $Y2=0
cc_895 N_A_2710_56#_c_1302_n N_Q_N_c_1803_n 0.0384027f $X=14.29 $Y=1.35 $X2=0
+ $Y2=0
cc_896 N_A_2710_56#_c_1303_n N_Q_N_c_1803_n 0.0309185f $X=14.875 $Y=1.35 $X2=0
+ $Y2=0
cc_897 N_A_2710_56#_c_1301_n N_VGND_M1012_s 0.00242368f $X=14.2 $Y=1.225 $X2=0
+ $Y2=0
cc_898 N_A_2710_56#_c_1300_n N_VGND_c_1828_n 0.0293442f $X=13.69 $Y=0.49 $X2=0
+ $Y2=0
cc_899 N_A_2710_56#_c_1301_n N_VGND_c_1828_n 0.007449f $X=14.2 $Y=1.225 $X2=0
+ $Y2=0
cc_900 N_A_2710_56#_c_1296_n N_VGND_c_1829_n 0.0108704f $X=14.445 $Y=1.185 $X2=0
+ $Y2=0
cc_901 N_A_2710_56#_c_1298_n N_VGND_c_1829_n 6.97329e-19 $X=14.875 $Y=1.185
+ $X2=0 $Y2=0
cc_902 N_A_2710_56#_c_1300_n N_VGND_c_1829_n 0.0428127f $X=13.69 $Y=0.49 $X2=0
+ $Y2=0
cc_903 N_A_2710_56#_c_1301_n N_VGND_c_1829_n 0.0221062f $X=14.2 $Y=1.225 $X2=0
+ $Y2=0
cc_904 N_A_2710_56#_c_1303_n N_VGND_c_1829_n 0.00127882f $X=14.875 $Y=1.35 $X2=0
+ $Y2=0
cc_905 N_A_2710_56#_c_1298_n N_VGND_c_1831_n 0.00664252f $X=14.875 $Y=1.185
+ $X2=0 $Y2=0
cc_906 N_A_2710_56#_c_1300_n N_VGND_c_1842_n 0.0132762f $X=13.69 $Y=0.49 $X2=0
+ $Y2=0
cc_907 N_A_2710_56#_c_1296_n N_VGND_c_1843_n 0.00564095f $X=14.445 $Y=1.185
+ $X2=0 $Y2=0
cc_908 N_A_2710_56#_c_1298_n N_VGND_c_1843_n 0.00564131f $X=14.875 $Y=1.185
+ $X2=0 $Y2=0
cc_909 N_A_2710_56#_c_1296_n N_VGND_c_1847_n 0.00948291f $X=14.445 $Y=1.185
+ $X2=0 $Y2=0
cc_910 N_A_2710_56#_c_1298_n N_VGND_c_1847_n 0.0110509f $X=14.875 $Y=1.185 $X2=0
+ $Y2=0
cc_911 N_A_2710_56#_c_1300_n N_VGND_c_1847_n 0.0111688f $X=13.69 $Y=0.49 $X2=0
+ $Y2=0
cc_912 N_A_27_489#_c_1362_n N_VPWR_M1023_d 0.00218982f $X=1.785 $Y=2.375
+ $X2=-0.19 $Y2=1.655
cc_913 N_A_27_489#_c_1362_n N_VPWR_c_1395_n 0.0170224f $X=1.785 $Y=2.375 $X2=0
+ $Y2=0
cc_914 N_A_27_489#_c_1361_n N_VPWR_c_1409_n 0.0210467f $X=0.26 $Y=2.59 $X2=0
+ $Y2=0
cc_915 N_A_27_489#_M1023_s N_VPWR_c_1394_n 0.00212301f $X=0.135 $Y=2.445 $X2=0
+ $Y2=0
cc_916 N_A_27_489#_M1038_d N_VPWR_c_1394_n 0.00213122f $X=1.81 $Y=2.445 $X2=0
+ $Y2=0
cc_917 N_A_27_489#_c_1361_n N_VPWR_c_1394_n 0.0125689f $X=0.26 $Y=2.59 $X2=0
+ $Y2=0
cc_918 N_A_27_489#_c_1362_n A_204_489# 0.00366293f $X=1.785 $Y=2.375 $X2=-0.19
+ $Y2=1.655
cc_919 N_A_27_489#_c_1362_n N_A_182_120#_M1014_d 0.00176461f $X=1.785 $Y=2.375
+ $X2=0 $Y2=0
cc_920 N_A_27_489#_c_1362_n N_A_182_120#_c_1583_n 0.0147769f $X=1.785 $Y=2.375
+ $X2=0 $Y2=0
cc_921 N_A_27_489#_M1038_d N_A_182_120#_c_1570_n 0.00495471f $X=1.81 $Y=2.445
+ $X2=0 $Y2=0
cc_922 N_A_27_489#_c_1362_n N_A_182_120#_c_1570_n 0.00387154f $X=1.785 $Y=2.375
+ $X2=0 $Y2=0
cc_923 N_A_27_489#_c_1364_n N_A_182_120#_c_1570_n 0.0199304f $X=1.95 $Y=2.375
+ $X2=0 $Y2=0
cc_924 N_A_27_489#_c_1364_n N_A_182_120#_c_1561_n 0.0338886f $X=1.95 $Y=2.375
+ $X2=0 $Y2=0
cc_925 N_VPWR_c_1394_n A_204_489# 0.00899413f $X=15.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_926 N_VPWR_c_1394_n N_A_182_120#_M1014_d 0.0022517f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1395_n N_A_182_120#_c_1583_n 0.00858436f $X=0.71 $Y=2.795 $X2=0
+ $Y2=0
cc_928 N_VPWR_c_1407_n N_A_182_120#_c_1570_n 0.0401509f $X=3.36 $Y=3.33 $X2=0
+ $Y2=0
cc_929 N_VPWR_c_1394_n N_A_182_120#_c_1570_n 0.0248759f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1395_n N_A_182_120#_c_1584_n 0.00574666f $X=0.71 $Y=2.795 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1407_n N_A_182_120#_c_1584_n 0.0154229f $X=3.36 $Y=3.33 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1394_n N_A_182_120#_c_1584_n 0.00988605f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1396_n N_A_182_120#_c_1572_n 0.0137731f $X=3.445 $Y=2.88 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1407_n N_A_182_120#_c_1572_n 0.0473678f $X=3.36 $Y=3.33 $X2=0
+ $Y2=0
cc_935 N_VPWR_c_1394_n N_A_182_120#_c_1572_n 0.0270372f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_936 N_VPWR_c_1396_n N_A_182_120#_c_1601_n 0.0137152f $X=3.445 $Y=2.88 $X2=0
+ $Y2=0
cc_937 N_VPWR_M1004_d N_A_182_120#_c_1574_n 0.00537978f $X=4.44 $Y=2.125 $X2=0
+ $Y2=0
cc_938 N_VPWR_c_1397_n N_A_182_120#_c_1574_n 0.0214121f $X=4.58 $Y=2.8 $X2=0
+ $Y2=0
cc_939 N_VPWR_c_1394_n N_A_182_120#_c_1574_n 0.0112542f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_940 N_VPWR_c_1407_n N_A_182_120#_c_1575_n 0.0121143f $X=3.36 $Y=3.33 $X2=0
+ $Y2=0
cc_941 N_VPWR_c_1394_n N_A_182_120#_c_1575_n 0.00659864f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_942 N_VPWR_M1005_d N_A_182_120#_c_1576_n 0.0039281f $X=3.255 $Y=2.405 $X2=0
+ $Y2=0
cc_943 N_VPWR_c_1396_n N_A_182_120#_c_1576_n 0.0212608f $X=3.445 $Y=2.88 $X2=0
+ $Y2=0
cc_944 N_VPWR_c_1394_n N_A_182_120#_c_1576_n 0.0330602f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_945 N_VPWR_c_1411_n N_A_993_425#_c_1724_n 0.0801074f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_946 N_VPWR_c_1394_n N_A_993_425#_c_1724_n 0.0455557f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_947 N_VPWR_c_1397_n N_A_993_425#_c_1725_n 0.0206938f $X=4.58 $Y=2.8 $X2=0
+ $Y2=0
cc_948 N_VPWR_c_1411_n N_A_993_425#_c_1725_n 0.0213714f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_949 N_VPWR_c_1394_n N_A_993_425#_c_1725_n 0.0110524f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_950 N_VPWR_c_1411_n N_A_993_425#_c_1726_n 0.0214121f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_951 N_VPWR_c_1394_n N_A_993_425#_c_1726_n 0.0110604f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_952 N_VPWR_c_1394_n N_Q_M1022_s 0.00387813f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_953 N_VPWR_M1022_d N_Q_c_1763_n 0.00303163f $X=12.2 $Y=1.835 $X2=0 $Y2=0
cc_954 N_VPWR_M1022_d N_Q_c_1776_n 0.00220581f $X=12.2 $Y=1.835 $X2=0 $Y2=0
cc_955 N_VPWR_M1022_d Q 6.40254e-19 $X=12.2 $Y=1.835 $X2=0 $Y2=0
cc_956 N_VPWR_c_1394_n N_Q_N_M1008_s 0.00345315f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_957 N_VPWR_c_1406_n N_Q_N_c_1803_n 0.0463491f $X=15.09 $Y=1.98 $X2=0 $Y2=0
cc_958 N_VPWR_c_1414_n N_Q_N_c_1803_n 0.0153611f $X=14.985 $Y=3.33 $X2=0 $Y2=0
cc_959 N_VPWR_c_1394_n N_Q_N_c_1803_n 0.00989321f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_960 N_A_182_120#_c_1574_n N_A_993_425#_M1033_d 0.00599097f $X=5.605 $Y=2.46
+ $X2=-0.19 $Y2=-0.245
cc_961 N_A_182_120#_M1039_s N_A_993_425#_c_1724_n 0.0032703f $X=5.625 $Y=2.505
+ $X2=0 $Y2=0
cc_962 N_A_182_120#_c_1574_n N_A_993_425#_c_1724_n 0.00832904f $X=5.605 $Y=2.46
+ $X2=0 $Y2=0
cc_963 N_A_182_120#_c_1577_n N_A_993_425#_c_1724_n 0.0237737f $X=5.77 $Y=2.46
+ $X2=0 $Y2=0
cc_964 N_A_182_120#_c_1574_n N_A_993_425#_c_1725_n 0.0248111f $X=5.605 $Y=2.46
+ $X2=0 $Y2=0
cc_965 N_A_182_120#_c_1577_n N_A_993_425#_c_1725_n 0.00130726f $X=5.77 $Y=2.46
+ $X2=0 $Y2=0
cc_966 N_A_182_120#_c_1565_n N_VGND_M1013_d 0.0123126f $X=4.455 $Y=1.335 $X2=0
+ $Y2=0
cc_967 N_A_182_120#_c_1569_n N_VGND_c_1822_n 0.0110667f $X=1.05 $Y=0.81 $X2=0
+ $Y2=0
cc_968 N_A_182_120#_c_1560_n N_VGND_c_1823_n 0.02448f $X=2.295 $Y=1.122 $X2=0
+ $Y2=0
cc_969 N_A_182_120#_c_1569_n N_VGND_c_1823_n 0.00596803f $X=1.05 $Y=0.81 $X2=0
+ $Y2=0
cc_970 N_A_182_120#_c_1563_n N_VGND_c_1824_n 0.0150385f $X=4.37 $Y=0.38 $X2=0
+ $Y2=0
cc_971 N_A_182_120#_c_1565_n N_VGND_c_1824_n 0.0538295f $X=4.455 $Y=1.335 $X2=0
+ $Y2=0
cc_972 N_A_182_120#_c_1566_n N_VGND_c_1824_n 0.0271222f $X=6.09 $Y=1.42 $X2=0
+ $Y2=0
cc_973 N_A_182_120#_c_1569_n N_VGND_c_1832_n 0.00501465f $X=1.05 $Y=0.81 $X2=0
+ $Y2=0
cc_974 N_A_182_120#_c_1563_n N_VGND_c_1834_n 0.044359f $X=4.37 $Y=0.38 $X2=0
+ $Y2=0
cc_975 N_A_182_120#_c_1564_n N_VGND_c_1834_n 0.00963698f $X=3.69 $Y=0.38 $X2=0
+ $Y2=0
cc_976 N_A_182_120#_c_1563_n N_VGND_c_1847_n 0.0279031f $X=4.37 $Y=0.38 $X2=0
+ $Y2=0
cc_977 N_A_182_120#_c_1564_n N_VGND_c_1847_n 0.0063608f $X=3.69 $Y=0.38 $X2=0
+ $Y2=0
cc_978 N_A_182_120#_c_1569_n N_VGND_c_1847_n 0.00841298f $X=1.05 $Y=0.81 $X2=0
+ $Y2=0
cc_979 N_Q_c_1759_n N_VGND_M1002_s 5.5277e-19 $X=12.64 $Y=1.135 $X2=0 $Y2=0
cc_980 N_Q_c_1761_n N_VGND_M1002_s 0.0020446f $X=12.222 $Y=1.22 $X2=0 $Y2=0
cc_981 N_Q_c_1759_n N_VGND_c_1827_n 0.00606161f $X=12.64 $Y=1.135 $X2=0 $Y2=0
cc_982 N_Q_c_1760_n N_VGND_c_1827_n 0.0240123f $X=12.735 $Y=0.425 $X2=0 $Y2=0
cc_983 N_Q_c_1761_n N_VGND_c_1827_n 0.0176293f $X=12.222 $Y=1.22 $X2=0 $Y2=0
cc_984 N_Q_c_1759_n N_VGND_c_1828_n 0.00168489f $X=12.64 $Y=1.135 $X2=0 $Y2=0
cc_985 N_Q_c_1760_n N_VGND_c_1828_n 0.00154423f $X=12.735 $Y=0.425 $X2=0 $Y2=0
cc_986 N_Q_c_1760_n N_VGND_c_1841_n 0.0158441f $X=12.735 $Y=0.425 $X2=0 $Y2=0
cc_987 N_Q_c_1760_n N_VGND_c_1847_n 0.00884325f $X=12.735 $Y=0.425 $X2=0 $Y2=0
cc_988 N_Q_N_c_1803_n N_VGND_c_1831_n 0.0307723f $X=14.66 $Y=0.42 $X2=0 $Y2=0
cc_989 N_Q_N_c_1803_n N_VGND_c_1843_n 0.0153611f $X=14.66 $Y=0.42 $X2=0 $Y2=0
cc_990 N_Q_N_M1012_d N_VGND_c_1847_n 0.00345315f $X=14.52 $Y=0.235 $X2=0 $Y2=0
cc_991 N_Q_N_c_1803_n N_VGND_c_1847_n 0.00989321f $X=14.66 $Y=0.42 $X2=0 $Y2=0
