* File: sky130_fd_sc_lp__a211oi_m.spice
* Created: Fri Aug 28 09:48:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a211oi_m.pex.spice"
.subckt sky130_fd_sc_lp__a211oi_m  VNB VPB A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1005 A_110_47# N_A2_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A1_M1001_g A_110_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=25.704 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_27_369#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_27_369#_M1006_d N_A1_M1006_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0693 AS=0.0819 PD=0.75 PS=0.81 NRD=0 NRS=42.1974 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 A_314_369# N_B1_M1002_g N_A_27_369#_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0567 AS=0.0693 PD=0.69 PS=0.75 NRD=37.5088 NRS=23.443 M=1 R=2.8
+ SA=75001.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_C1_M1000_g A_314_369# VPB PHIGHVT L=0.15 W=0.42 AD=0.1113
+ AS=0.0567 PD=1.37 PS=0.69 NRD=0 NRS=37.5088 M=1 R=2.8 SA=75001.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__a211oi_m.pxi.spice"
*
.ends
*
*
