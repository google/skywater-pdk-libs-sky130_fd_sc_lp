* File: sky130_fd_sc_lp__a311oi_1.spice
* Created: Wed Sep  2 09:25:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a311oi_1  VNB VPB A3 A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1003 A_181_47# N_A3_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.1239
+ AS=0.2226 PD=1.135 PS=2.21 NRD=13.212 NRS=0 M=1 R=5.6 SA=75000.2 SB=75002.2
+ A=0.126 P=1.98 MULT=1
MM1008 A_270_47# N_A2_M1008_g A_181_47# VNB NSHORT L=0.15 W=0.84 AD=0.1281
+ AS=0.1239 PD=1.145 PS=1.135 NRD=13.92 NRS=13.212 M=1 R=5.6 SA=75000.6
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1007 N_Y_M1007_d N_A1_M1007_g A_270_47# VNB NSHORT L=0.15 W=0.84 AD=0.1764
+ AS=0.1281 PD=1.26 PS=1.145 NRD=18.564 NRS=13.92 M=1 R=5.6 SA=75001.1
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1827 AS=0.1764 PD=1.275 PS=1.26 NRD=10.704 NRS=1.428 M=1 R=5.6 SA=75001.7
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1004_d N_C1_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1827 PD=2.21 PS=1.275 NRD=0 NRS=11.424 M=1 R=5.6 SA=75002.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_A_181_367#_M1009_d N_A3_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.19215 AS=0.3339 PD=1.565 PS=3.05 NRD=3.9006 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_181_367#_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.31815 AS=0.19215 PD=1.765 PS=1.565 NRD=19.5424 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.8 A=0.189 P=2.82 MULT=1
MM1001 N_A_181_367#_M1001_d N_A1_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.27405 AS=0.31815 PD=1.695 PS=1.765 NRD=13.2778 NRS=15.6221 M=1
+ R=8.4 SA=75001.3 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 A_520_367# N_B1_M1005_g N_A_181_367#_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.27405 PD=1.47 PS=1.695 NRD=7.8012 NRS=10.9335 M=1 R=8.4
+ SA=75001.9 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_C1_M1006_g A_520_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.3339
+ AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75002.2 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a311oi_1.pxi.spice"
*
.ends
*
*
