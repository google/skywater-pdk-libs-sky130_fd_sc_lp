* File: sky130_fd_sc_lp__iso0p_lp2.pxi.spice
* Created: Fri Aug 28 10:40:47 2020
* 
x_PM_SKY130_FD_SC_LP__ISO0P_LP2%SLEEP N_SLEEP_c_53_n N_SLEEP_M1008_g
+ N_SLEEP_M1007_g N_SLEEP_c_54_n N_SLEEP_M1003_g SLEEP SLEEP N_SLEEP_c_55_n
+ N_SLEEP_c_56_n PM_SKY130_FD_SC_LP__ISO0P_LP2%SLEEP
x_PM_SKY130_FD_SC_LP__ISO0P_LP2%A_27_93# N_A_27_93#_M1008_s N_A_27_93#_M1007_s
+ N_A_27_93#_c_83_n N_A_27_93#_M1009_g N_A_27_93#_c_84_n N_A_27_93#_M1004_g
+ N_A_27_93#_c_85_n N_A_27_93#_c_123_p N_A_27_93#_c_90_n N_A_27_93#_c_86_n
+ N_A_27_93#_c_92_n PM_SKY130_FD_SC_LP__ISO0P_LP2%A_27_93#
x_PM_SKY130_FD_SC_LP__ISO0P_LP2%A N_A_M1000_g N_A_c_142_n N_A_M1005_g
+ N_A_c_144_n N_A_c_145_n A A N_A_c_147_n N_A_c_148_n
+ PM_SKY130_FD_SC_LP__ISO0P_LP2%A
x_PM_SKY130_FD_SC_LP__ISO0P_LP2%A_342_417# N_A_342_417#_M1000_d
+ N_A_342_417#_M1009_d N_A_342_417#_c_188_n N_A_342_417#_M1001_g
+ N_A_342_417#_M1006_g N_A_342_417#_c_189_n N_A_342_417#_M1002_g
+ N_A_342_417#_c_223_p N_A_342_417#_c_196_n N_A_342_417#_c_197_n
+ N_A_342_417#_c_190_n N_A_342_417#_c_191_n N_A_342_417#_c_192_n
+ N_A_342_417#_c_193_n N_A_342_417#_c_198_n N_A_342_417#_c_194_n
+ PM_SKY130_FD_SC_LP__ISO0P_LP2%A_342_417#
x_PM_SKY130_FD_SC_LP__ISO0P_LP2%KAPWR N_KAPWR_M1007_d N_KAPWR_M1005_d KAPWR
+ N_KAPWR_c_253_n N_KAPWR_c_264_n N_KAPWR_c_252_n
+ PM_SKY130_FD_SC_LP__ISO0P_LP2%KAPWR
x_PM_SKY130_FD_SC_LP__ISO0P_LP2%X N_X_M1002_d N_X_M1006_d X X X X X N_X_c_287_n
+ PM_SKY130_FD_SC_LP__ISO0P_LP2%X
x_PM_SKY130_FD_SC_LP__ISO0P_LP2%VGND N_VGND_M1003_d N_VGND_M1001_s
+ N_VGND_c_301_n N_VGND_c_302_n VGND N_VGND_c_303_n N_VGND_c_304_n
+ N_VGND_c_305_n N_VGND_c_306_n N_VGND_c_307_n N_VGND_c_308_n
+ PM_SKY130_FD_SC_LP__ISO0P_LP2%VGND
x_PM_SKY130_FD_SC_LP__ISO0P_LP2%VPWR VPWR N_VPWR_c_343_n VPWR
+ PM_SKY130_FD_SC_LP__ISO0P_LP2%VPWR
cc_1 VNB N_SLEEP_c_53_n 0.0196793f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.01
cc_2 VNB N_SLEEP_c_54_n 0.0184753f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.01
cc_3 VNB N_SLEEP_c_55_n 0.063957f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.175
cc_4 VNB N_SLEEP_c_56_n 0.00122182f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.175
cc_5 VNB N_A_27_93#_c_83_n 0.0700145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_93#_c_84_n 0.0188999f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_A_27_93#_c_85_n 0.042136f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.175
cc_8 VNB N_A_27_93#_c_86_n 0.0032708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_142_n 0.0123327f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.585
cc_10 VNB N_A_M1005_g 5.66077e-19 $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.01
cc_11 VNB N_A_c_144_n 0.017557f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.675
cc_12 VNB N_A_c_145_n 0.0170663f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB A 0.00476803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_c_147_n 0.0377061f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.685
cc_15 VNB N_A_c_148_n 0.0187342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_342_417#_c_188_n 0.0188631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_342_417#_c_189_n 0.020326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_342_417#_c_190_n 0.00555058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_342_417#_c_191_n 0.0211155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_342_417#_c_192_n 0.00104353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_342_417#_c_193_n 0.00122182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_342_417#_c_194_n 0.0685529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_287_n 0.0647669f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.685
cc_24 VNB N_VGND_c_301_n 0.0162715f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.675
cc_25 VNB N_VGND_c_302_n 0.0186777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_303_n 0.0291685f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.175
cc_27 VNB N_VGND_c_304_n 0.0295741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_305_n 0.0303334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_306_n 0.271448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_307_n 0.0130796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_308_n 0.00644364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB VPWR 0.163682f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.01
cc_33 VPB N_SLEEP_M1007_g 0.0536538f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.585
cc_34 VPB N_SLEEP_c_55_n 0.0103677f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.175
cc_35 VPB N_SLEEP_c_56_n 0.00326766f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.175
cc_36 VPB N_A_27_93#_c_83_n 0.00974876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_27_93#_M1009_g 0.049197f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.675
cc_38 VPB N_A_27_93#_c_85_n 0.0141159f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.175
cc_39 VPB N_A_27_93#_c_90_n 0.014596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_27_93#_c_86_n 0.00362611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_27_93#_c_92_n 0.0058727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_M1005_g 0.050667f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.01
cc_43 VPB A 0.00664533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_342_417#_M1006_g 0.0525377f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_45 VPB N_A_342_417#_c_196_n 0.0105624f $X=-0.19 $Y=1.655 $X2=0.732 $Y2=1.665
cc_46 VPB N_A_342_417#_c_197_n 0.00957918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_342_417#_c_198_n 0.00379314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_342_417#_c_194_n 0.0105597f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_KAPWR_c_252_n 0.0220396f $X=-0.19 $Y=1.655 $X2=0.732 $Y2=1.295
cc_50 VPB N_X_c_287_n 0.0609139f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.685
cc_51 VPB VPWR 0.0448742f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.01
cc_52 VPB N_VPWR_c_343_n 0.102188f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.01
cc_53 N_SLEEP_c_55_n N_A_27_93#_c_83_n 0.03063f $X=0.71 $Y=1.175 $X2=0 $Y2=0
cc_54 N_SLEEP_c_56_n N_A_27_93#_c_83_n 0.00282527f $X=0.71 $Y=1.175 $X2=0 $Y2=0
cc_55 N_SLEEP_c_56_n N_A_27_93#_M1009_g 4.09251e-19 $X=0.71 $Y=1.175 $X2=0 $Y2=0
cc_56 N_SLEEP_c_54_n N_A_27_93#_c_84_n 0.00511621f $X=0.845 $Y=1.01 $X2=0 $Y2=0
cc_57 N_SLEEP_c_53_n N_A_27_93#_c_85_n 0.0364623f $X=0.485 $Y=1.01 $X2=0 $Y2=0
cc_58 N_SLEEP_c_56_n N_A_27_93#_c_85_n 0.0595519f $X=0.71 $Y=1.175 $X2=0 $Y2=0
cc_59 N_SLEEP_M1007_g N_A_27_93#_c_90_n 0.023693f $X=0.535 $Y=2.585 $X2=0 $Y2=0
cc_60 N_SLEEP_c_55_n N_A_27_93#_c_90_n 0.00140772f $X=0.71 $Y=1.175 $X2=0 $Y2=0
cc_61 N_SLEEP_c_56_n N_A_27_93#_c_90_n 0.0305572f $X=0.71 $Y=1.175 $X2=0 $Y2=0
cc_62 N_SLEEP_M1007_g N_A_27_93#_c_86_n 0.00501581f $X=0.535 $Y=2.585 $X2=0
+ $Y2=0
cc_63 N_SLEEP_c_55_n N_A_27_93#_c_86_n 0.0028784f $X=0.71 $Y=1.175 $X2=0 $Y2=0
cc_64 N_SLEEP_c_56_n N_A_27_93#_c_86_n 0.0405531f $X=0.71 $Y=1.175 $X2=0 $Y2=0
cc_65 N_SLEEP_M1007_g N_KAPWR_c_253_n 0.0158972f $X=0.535 $Y=2.585 $X2=0 $Y2=0
cc_66 N_SLEEP_M1007_g N_KAPWR_c_252_n 0.00547899f $X=0.535 $Y=2.585 $X2=0 $Y2=0
cc_67 N_SLEEP_c_53_n N_VGND_c_301_n 0.00161762f $X=0.485 $Y=1.01 $X2=0 $Y2=0
cc_68 N_SLEEP_c_54_n N_VGND_c_301_n 0.0124399f $X=0.845 $Y=1.01 $X2=0 $Y2=0
cc_69 N_SLEEP_c_56_n N_VGND_c_301_n 0.00194697f $X=0.71 $Y=1.175 $X2=0 $Y2=0
cc_70 N_SLEEP_c_53_n N_VGND_c_303_n 0.00510437f $X=0.485 $Y=1.01 $X2=0 $Y2=0
cc_71 N_SLEEP_c_54_n N_VGND_c_303_n 0.00424179f $X=0.845 $Y=1.01 $X2=0 $Y2=0
cc_72 N_SLEEP_c_53_n N_VGND_c_306_n 0.00515964f $X=0.485 $Y=1.01 $X2=0 $Y2=0
cc_73 N_SLEEP_c_54_n N_VGND_c_306_n 0.0043341f $X=0.845 $Y=1.01 $X2=0 $Y2=0
cc_74 N_SLEEP_M1007_g VPWR 0.0104709f $X=0.535 $Y=2.585 $X2=-0.19 $Y2=-0.245
cc_75 N_SLEEP_M1007_g N_VPWR_c_343_n 0.00939206f $X=0.535 $Y=2.585 $X2=0 $Y2=0
cc_76 N_A_27_93#_c_83_n N_A_c_142_n 0.00859206f $X=1.585 $Y=1.68 $X2=0 $Y2=0
cc_77 N_A_27_93#_c_86_n N_A_c_142_n 0.00116732f $X=1.43 $Y=1.175 $X2=0 $Y2=0
cc_78 N_A_27_93#_c_83_n N_A_M1005_g 0.0251021f $X=1.585 $Y=1.68 $X2=0 $Y2=0
cc_79 N_A_27_93#_c_86_n N_A_M1005_g 0.00114805f $X=1.43 $Y=1.175 $X2=0 $Y2=0
cc_80 N_A_27_93#_c_84_n N_A_c_144_n 0.0242364f $X=1.625 $Y=1.01 $X2=0 $Y2=0
cc_81 N_A_27_93#_c_83_n N_A_c_145_n 0.0242364f $X=1.585 $Y=1.68 $X2=0 $Y2=0
cc_82 N_A_27_93#_c_86_n N_A_c_145_n 4.15826e-19 $X=1.43 $Y=1.175 $X2=0 $Y2=0
cc_83 N_A_27_93#_c_83_n A 0.00200383f $X=1.585 $Y=1.68 $X2=0 $Y2=0
cc_84 N_A_27_93#_c_86_n A 0.0152129f $X=1.43 $Y=1.175 $X2=0 $Y2=0
cc_85 N_A_27_93#_c_83_n N_A_c_148_n 0.0160243f $X=1.585 $Y=1.68 $X2=0 $Y2=0
cc_86 N_A_27_93#_c_86_n N_A_c_148_n 2.66615e-19 $X=1.43 $Y=1.175 $X2=0 $Y2=0
cc_87 N_A_27_93#_M1009_g N_A_342_417#_c_197_n 0.00114967f $X=1.585 $Y=2.585
+ $X2=0 $Y2=0
cc_88 N_A_27_93#_c_90_n N_A_342_417#_c_197_n 0.0130231f $X=1.2 $Y=2.035 $X2=0
+ $Y2=0
cc_89 N_A_27_93#_c_84_n N_A_342_417#_c_192_n 7.13207e-19 $X=1.625 $Y=1.01 $X2=0
+ $Y2=0
cc_90 N_A_27_93#_c_86_n N_A_342_417#_c_192_n 0.00717322f $X=1.43 $Y=1.175 $X2=0
+ $Y2=0
cc_91 N_A_27_93#_c_90_n N_KAPWR_M1007_d 0.00806642f $X=1.2 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_27_93#_c_83_n N_KAPWR_c_253_n 7.60099e-19 $X=1.585 $Y=1.68 $X2=0 $Y2=0
cc_93 N_A_27_93#_M1009_g N_KAPWR_c_253_n 0.0158374f $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_94 N_A_27_93#_c_123_p N_KAPWR_c_253_n 0.0239452f $X=0.27 $Y=2.23 $X2=0 $Y2=0
cc_95 N_A_27_93#_c_90_n N_KAPWR_c_253_n 0.0596276f $X=1.2 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_27_93#_M1007_s N_KAPWR_c_252_n 0.00156869f $X=0.135 $Y=2.085 $X2=0
+ $Y2=0
cc_97 N_A_27_93#_M1009_g N_KAPWR_c_252_n 0.00893175f $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_98 N_A_27_93#_c_123_p N_KAPWR_c_252_n 0.0285176f $X=0.27 $Y=2.23 $X2=0 $Y2=0
cc_99 N_A_27_93#_c_90_n N_KAPWR_c_252_n 0.0136833f $X=1.2 $Y=2.035 $X2=0 $Y2=0
cc_100 N_A_27_93#_c_83_n N_VGND_c_301_n 0.00255877f $X=1.585 $Y=1.68 $X2=0 $Y2=0
cc_101 N_A_27_93#_c_84_n N_VGND_c_301_n 0.0124399f $X=1.625 $Y=1.01 $X2=0 $Y2=0
cc_102 N_A_27_93#_c_85_n N_VGND_c_301_n 0.00748999f $X=0.27 $Y=0.72 $X2=0 $Y2=0
cc_103 N_A_27_93#_c_86_n N_VGND_c_301_n 0.029924f $X=1.43 $Y=1.175 $X2=0 $Y2=0
cc_104 N_A_27_93#_c_85_n N_VGND_c_303_n 0.00734893f $X=0.27 $Y=0.72 $X2=0 $Y2=0
cc_105 N_A_27_93#_c_84_n N_VGND_c_304_n 0.00424179f $X=1.625 $Y=1.01 $X2=0 $Y2=0
cc_106 N_A_27_93#_c_84_n N_VGND_c_306_n 0.0043341f $X=1.625 $Y=1.01 $X2=0 $Y2=0
cc_107 N_A_27_93#_c_85_n N_VGND_c_306_n 0.00765198f $X=0.27 $Y=0.72 $X2=0 $Y2=0
cc_108 N_A_27_93#_M1007_s VPWR 0.00148697f $X=0.135 $Y=2.085 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A_27_93#_M1009_g VPWR 0.00954039f $X=1.585 $Y=2.585 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_27_93#_c_123_p VPWR 0.00237013f $X=0.27 $Y=2.23 $X2=-0.19 $Y2=-0.245
cc_111 N_A_27_93#_M1009_g N_VPWR_c_343_n 0.00939206f $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_112 N_A_27_93#_c_123_p N_VPWR_c_343_n 0.0145967f $X=0.27 $Y=2.23 $X2=0 $Y2=0
cc_113 A N_A_342_417#_M1006_g 3.21608e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A_M1005_g N_A_342_417#_c_196_n 0.0185631f $X=2.135 $Y=2.585 $X2=0 $Y2=0
cc_115 A N_A_342_417#_c_196_n 0.0521732f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A_c_147_n N_A_342_417#_c_196_n 0.00206682f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_117 N_A_c_144_n N_A_342_417#_c_190_n 0.00656473f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_c_145_n N_A_342_417#_c_190_n 0.00111161f $X=2.02 $Y=1.145 $X2=0 $Y2=0
cc_119 A N_A_342_417#_c_191_n 0.0350828f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_120 N_A_c_147_n N_A_342_417#_c_191_n 0.00855509f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_121 N_A_c_142_n N_A_342_417#_c_192_n 0.0038137f $X=2.055 $Y=1.315 $X2=0 $Y2=0
cc_122 N_A_c_145_n N_A_342_417#_c_192_n 0.00610338f $X=2.02 $Y=1.145 $X2=0 $Y2=0
cc_123 A N_A_342_417#_c_192_n 0.0176014f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A_c_148_n N_A_342_417#_c_192_n 0.00503056f $X=2.145 $Y=1.48 $X2=0 $Y2=0
cc_125 N_A_M1005_g N_A_342_417#_c_198_n 0.00499172f $X=2.135 $Y=2.585 $X2=0
+ $Y2=0
cc_126 A N_A_342_417#_c_198_n 0.029869f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A_c_147_n N_A_342_417#_c_198_n 7.5756e-19 $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_128 N_A_M1005_g N_A_342_417#_c_194_n 5.24053e-19 $X=2.135 $Y=2.585 $X2=0
+ $Y2=0
cc_129 A N_A_342_417#_c_194_n 0.00235212f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A_c_147_n N_A_342_417#_c_194_n 0.02202f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_131 N_A_M1005_g N_KAPWR_c_264_n 0.0154411f $X=2.135 $Y=2.585 $X2=0 $Y2=0
cc_132 N_A_M1005_g N_KAPWR_c_252_n 0.00546148f $X=2.135 $Y=2.585 $X2=0 $Y2=0
cc_133 N_A_c_144_n N_VGND_c_301_n 0.00161762f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_144_n N_VGND_c_302_n 0.00333051f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_144_n N_VGND_c_304_n 0.00510437f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_c_144_n N_VGND_c_306_n 0.00515964f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_M1005_g VPWR 0.00954039f $X=2.135 $Y=2.585 $X2=-0.19 $Y2=-0.245
cc_138 N_A_M1005_g N_VPWR_c_343_n 0.00939206f $X=2.135 $Y=2.585 $X2=0 $Y2=0
cc_139 N_A_342_417#_c_196_n N_KAPWR_M1005_d 0.00890832f $X=2.925 $Y=2.04 $X2=0
+ $Y2=0
cc_140 N_A_342_417#_c_223_p N_KAPWR_c_253_n 0.0223967f $X=1.87 $Y=2.23 $X2=0
+ $Y2=0
cc_141 N_A_342_417#_M1006_g N_KAPWR_c_264_n 0.0157309f $X=3.245 $Y=2.585 $X2=0
+ $Y2=0
cc_142 N_A_342_417#_c_223_p N_KAPWR_c_264_n 0.023792f $X=1.87 $Y=2.23 $X2=0
+ $Y2=0
cc_143 N_A_342_417#_c_196_n N_KAPWR_c_264_n 0.0638026f $X=2.925 $Y=2.04 $X2=0
+ $Y2=0
cc_144 N_A_342_417#_c_194_n N_KAPWR_c_264_n 6.55345e-19 $X=3.06 $Y=1.17 $X2=0
+ $Y2=0
cc_145 N_A_342_417#_M1009_d N_KAPWR_c_252_n 0.00302349f $X=1.71 $Y=2.085 $X2=0
+ $Y2=0
cc_146 N_A_342_417#_M1006_g N_KAPWR_c_252_n 0.00938018f $X=3.245 $Y=2.585 $X2=0
+ $Y2=0
cc_147 N_A_342_417#_c_223_p N_KAPWR_c_252_n 0.0260106f $X=1.87 $Y=2.23 $X2=0
+ $Y2=0
cc_148 N_A_342_417#_c_196_n N_KAPWR_c_252_n 0.013166f $X=2.925 $Y=2.04 $X2=0
+ $Y2=0
cc_149 N_A_342_417#_c_189_n N_X_c_287_n 0.0371006f $X=3.295 $Y=1.005 $X2=0 $Y2=0
cc_150 N_A_342_417#_c_196_n N_X_c_287_n 0.0126104f $X=2.925 $Y=2.04 $X2=0 $Y2=0
cc_151 N_A_342_417#_c_193_n N_X_c_287_n 0.0185607f $X=3.077 $Y=1.225 $X2=0 $Y2=0
cc_152 N_A_342_417#_c_198_n N_X_c_287_n 0.0576603f $X=3.077 $Y=1.955 $X2=0 $Y2=0
cc_153 N_A_342_417#_c_190_n N_VGND_c_301_n 0.00748572f $X=2.2 $Y=0.72 $X2=0
+ $Y2=0
cc_154 N_A_342_417#_c_188_n N_VGND_c_302_n 0.0132056f $X=2.935 $Y=1.005 $X2=0
+ $Y2=0
cc_155 N_A_342_417#_c_189_n N_VGND_c_302_n 0.00168986f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_156 N_A_342_417#_c_190_n N_VGND_c_302_n 0.0247472f $X=2.2 $Y=0.72 $X2=0 $Y2=0
cc_157 N_A_342_417#_c_191_n N_VGND_c_302_n 0.0253566f $X=2.925 $Y=1.115 $X2=0
+ $Y2=0
cc_158 N_A_342_417#_c_190_n N_VGND_c_304_n 0.00701182f $X=2.2 $Y=0.72 $X2=0
+ $Y2=0
cc_159 N_A_342_417#_c_188_n N_VGND_c_305_n 0.00424179f $X=2.935 $Y=1.005 $X2=0
+ $Y2=0
cc_160 N_A_342_417#_c_189_n N_VGND_c_305_n 0.00510437f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_161 N_A_342_417#_c_188_n N_VGND_c_306_n 0.0043341f $X=2.935 $Y=1.005 $X2=0
+ $Y2=0
cc_162 N_A_342_417#_c_189_n N_VGND_c_306_n 0.00515964f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_163 N_A_342_417#_c_190_n N_VGND_c_306_n 0.00730097f $X=2.2 $Y=0.72 $X2=0
+ $Y2=0
cc_164 N_A_342_417#_M1009_d VPWR 0.0017499f $X=1.71 $Y=2.085 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A_342_417#_M1006_g VPWR 0.0105252f $X=3.245 $Y=2.585 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A_342_417#_c_223_p VPWR 0.00225613f $X=1.87 $Y=2.23 $X2=-0.19
+ $Y2=-0.245
cc_167 N_A_342_417#_M1006_g N_VPWR_c_343_n 0.00939206f $X=3.245 $Y=2.585 $X2=0
+ $Y2=0
cc_168 N_A_342_417#_c_223_p N_VPWR_c_343_n 0.0138587f $X=1.87 $Y=2.23 $X2=0
+ $Y2=0
cc_169 N_KAPWR_c_252_n N_X_M1006_d 0.00127496f $X=2.98 $Y=2.775 $X2=0 $Y2=0
cc_170 N_KAPWR_c_264_n N_X_c_287_n 0.0242547f $X=2.98 $Y=2.395 $X2=0 $Y2=0
cc_171 N_KAPWR_c_252_n N_X_c_287_n 0.0402347f $X=2.98 $Y=2.775 $X2=0 $Y2=0
cc_172 N_KAPWR_M1007_d VPWR 0.00358693f $X=0.66 $Y=2.085 $X2=-0.19 $Y2=1.655
cc_173 N_KAPWR_M1005_d VPWR 0.00385662f $X=2.26 $Y=2.085 $X2=-0.19 $Y2=1.655
cc_174 N_KAPWR_c_253_n VPWR 0.00911842f $X=1.32 $Y=2.395 $X2=-0.19 $Y2=1.655
cc_175 N_KAPWR_c_264_n VPWR 0.00977075f $X=2.98 $Y=2.395 $X2=-0.19 $Y2=1.655
cc_176 N_KAPWR_c_252_n VPWR 0.328419f $X=2.98 $Y=2.775 $X2=-0.19 $Y2=1.655
cc_177 N_KAPWR_c_253_n N_VPWR_c_343_n 0.0554861f $X=1.32 $Y=2.395 $X2=0 $Y2=0
cc_178 N_KAPWR_c_264_n N_VPWR_c_343_n 0.0597049f $X=2.98 $Y=2.395 $X2=0 $Y2=0
cc_179 N_KAPWR_c_252_n N_VPWR_c_343_n 0.00754143f $X=2.98 $Y=2.775 $X2=0 $Y2=0
cc_180 N_X_c_287_n N_VGND_c_305_n 0.0101312f $X=3.51 $Y=0.72 $X2=0 $Y2=0
cc_181 N_X_c_287_n N_VGND_c_306_n 0.0121005f $X=3.51 $Y=0.72 $X2=0 $Y2=0
cc_182 N_X_M1006_d VPWR 0.00132346f $X=3.37 $Y=2.085 $X2=-0.19 $Y2=-0.245
cc_183 N_X_c_287_n VPWR 0.00383788f $X=3.51 $Y=0.72 $X2=-0.19 $Y2=-0.245
cc_184 N_X_c_287_n N_VPWR_c_343_n 0.0240782f $X=3.51 $Y=0.72 $X2=0 $Y2=0
