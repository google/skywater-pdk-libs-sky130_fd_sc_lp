* NGSPICE file created from sky130_fd_sc_lp__a311o_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a311o_m A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 VGND B1 a_54_154# VNB nshort w=420000u l=150000u
+  ad=2.982e+11p pd=3.1e+06u as=2.289e+11p ps=2.77e+06u
M1001 VGND a_54_154# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1002 VPWR a_54_154# X VPB phighvt w=420000u l=150000u
+  ad=3.1835e+11p pd=3.23e+06u as=1.113e+11p ps=1.37e+06u
M1003 VPWR A2 a_196_403# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1004 a_486_403# B1 a_196_403# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 a_54_154# C1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_220_48# A3 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 a_54_154# C1 a_486_403# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 a_292_48# A2 a_220_48# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 a_54_154# A1 a_292_48# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_196_403# A1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_196_403# A3 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

