* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4b_4 A B C D_N VGND VNB VPB VPWR X
X0 X a_83_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND C a_83_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_659_367# a_737_315# a_83_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND D_N a_737_315# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_83_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_83_21# a_737_315# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 X a_83_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_551_367# C a_659_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR A a_479_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR a_83_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR D_N a_737_315# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VPWR a_83_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND A a_83_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_83_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_479_367# B a_551_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 X a_83_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 X a_83_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VGND a_83_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
