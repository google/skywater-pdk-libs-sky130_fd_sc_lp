* NGSPICE file created from sky130_fd_sc_lp__clkdlybuf4s25_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
M1000 X a_394_52# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=1.35e+12p ps=7.48e+06u
M1001 VPWR a_282_52# a_394_52# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1002 a_282_52# a_27_52# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1003 VGND A a_27_52# VNB nshort w=420000u l=150000u
+  ad=1.0924e+12p pd=6.44e+06u as=1.113e+11p ps=1.37e+06u
M1004 a_282_52# a_27_52# VGND VNB nshort w=1e+06u l=250000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1005 X a_394_52# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 VGND a_282_52# a_394_52# VNB nshort w=1e+06u l=250000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1007 VPWR A a_27_52# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

