* File: sky130_fd_sc_lp__bufbuf_16.pxi.spice
* Created: Fri Aug 28 10:10:58 2020
* 
x_PM_SKY130_FD_SC_LP__BUFBUF_16%A N_A_M1018_g N_A_M1051_g A N_A_c_242_n
+ N_A_c_243_n PM_SKY130_FD_SC_LP__BUFBUF_16%A
x_PM_SKY130_FD_SC_LP__BUFBUF_16%A_27_49# N_A_27_49#_M1018_s N_A_27_49#_M1051_s
+ N_A_27_49#_M1027_g N_A_27_49#_M1001_g N_A_27_49#_M1032_g N_A_27_49#_M1022_g
+ N_A_27_49#_M1048_g N_A_27_49#_M1039_g N_A_27_49#_c_274_n N_A_27_49#_c_286_n
+ N_A_27_49#_c_287_n N_A_27_49#_c_275_n N_A_27_49#_c_276_n N_A_27_49#_c_300_n
+ N_A_27_49#_c_277_n N_A_27_49#_c_278_n N_A_27_49#_c_279_n N_A_27_49#_c_280_n
+ N_A_27_49#_c_281_n N_A_27_49#_c_282_n PM_SKY130_FD_SC_LP__BUFBUF_16%A_27_49#
x_PM_SKY130_FD_SC_LP__BUFBUF_16%A_196_49# N_A_196_49#_M1027_d
+ N_A_196_49#_M1048_d N_A_196_49#_M1001_s N_A_196_49#_M1039_s
+ N_A_196_49#_M1008_g N_A_196_49#_M1003_g N_A_196_49#_M1011_g
+ N_A_196_49#_M1019_g N_A_196_49#_M1023_g N_A_196_49#_M1025_g
+ N_A_196_49#_M1029_g N_A_196_49#_M1040_g N_A_196_49#_M1033_g
+ N_A_196_49#_M1041_g N_A_196_49#_M1035_g N_A_196_49#_M1042_g
+ N_A_196_49#_c_498_p N_A_196_49#_c_530_p N_A_196_49#_c_386_n
+ N_A_196_49#_c_387_n N_A_196_49#_c_399_n N_A_196_49#_c_400_n
+ N_A_196_49#_c_388_n N_A_196_49#_c_401_n N_A_196_49#_c_389_n
+ N_A_196_49#_c_402_n N_A_196_49#_c_390_n N_A_196_49#_c_440_p
+ N_A_196_49#_c_391_n N_A_196_49#_c_404_n N_A_196_49#_c_392_n
+ PM_SKY130_FD_SC_LP__BUFBUF_16%A_196_49#
x_PM_SKY130_FD_SC_LP__BUFBUF_16%A_610_47# N_A_610_47#_M1008_s
+ N_A_610_47#_M1023_s N_A_610_47#_M1033_s N_A_610_47#_M1003_d
+ N_A_610_47#_M1025_d N_A_610_47#_M1041_d N_A_610_47#_M1002_g
+ N_A_610_47#_M1000_g N_A_610_47#_M1006_g N_A_610_47#_M1004_g
+ N_A_610_47#_M1009_g N_A_610_47#_M1005_g N_A_610_47#_M1012_g
+ N_A_610_47#_M1007_g N_A_610_47#_M1013_g N_A_610_47#_M1010_g
+ N_A_610_47#_M1014_g N_A_610_47#_M1015_g N_A_610_47#_M1016_g
+ N_A_610_47#_M1017_g N_A_610_47#_M1024_g N_A_610_47#_M1020_g
+ N_A_610_47#_M1028_g N_A_610_47#_M1021_g N_A_610_47#_M1030_g
+ N_A_610_47#_M1026_g N_A_610_47#_M1034_g N_A_610_47#_M1031_g
+ N_A_610_47#_M1038_g N_A_610_47#_M1036_g N_A_610_47#_M1043_g
+ N_A_610_47#_M1037_g N_A_610_47#_M1044_g N_A_610_47#_M1045_g
+ N_A_610_47#_M1046_g N_A_610_47#_M1047_g N_A_610_47#_M1049_g
+ N_A_610_47#_M1050_g N_A_610_47#_c_898_p N_A_610_47#_c_724_p
+ N_A_610_47#_c_575_n N_A_610_47#_c_576_n N_A_610_47#_c_607_n
+ N_A_610_47#_c_608_n N_A_610_47#_c_888_p N_A_610_47#_c_714_p
+ N_A_610_47#_c_577_n N_A_610_47#_c_609_n N_A_610_47#_c_889_p
+ N_A_610_47#_c_715_p N_A_610_47#_c_578_n N_A_610_47#_c_610_n
+ N_A_610_47#_c_579_n N_A_610_47#_c_611_n N_A_610_47#_c_580_n
+ N_A_610_47#_c_612_n N_A_610_47#_c_581_n N_A_610_47#_c_582_n
+ N_A_610_47#_c_583_n N_A_610_47#_c_584_n N_A_610_47#_c_585_n
+ N_A_610_47#_c_586_n N_A_610_47#_c_587_n N_A_610_47#_c_588_n
+ N_A_610_47#_c_589_n N_A_610_47#_c_590_n
+ PM_SKY130_FD_SC_LP__BUFBUF_16%A_610_47#
x_PM_SKY130_FD_SC_LP__BUFBUF_16%VPWR N_VPWR_M1051_d N_VPWR_M1022_d
+ N_VPWR_M1003_s N_VPWR_M1019_s N_VPWR_M1040_s N_VPWR_M1042_s N_VPWR_M1004_s
+ N_VPWR_M1007_s N_VPWR_M1015_s N_VPWR_M1020_s N_VPWR_M1026_s N_VPWR_M1036_s
+ N_VPWR_M1045_s N_VPWR_M1050_s N_VPWR_c_926_n N_VPWR_c_927_n N_VPWR_c_928_n
+ N_VPWR_c_929_n N_VPWR_c_930_n N_VPWR_c_931_n N_VPWR_c_932_n N_VPWR_c_933_n
+ N_VPWR_c_934_n N_VPWR_c_935_n N_VPWR_c_936_n N_VPWR_c_937_n N_VPWR_c_938_n
+ N_VPWR_c_939_n N_VPWR_c_940_n N_VPWR_c_941_n N_VPWR_c_942_n N_VPWR_c_943_n
+ N_VPWR_c_944_n N_VPWR_c_945_n N_VPWR_c_946_n N_VPWR_c_947_n N_VPWR_c_948_n
+ N_VPWR_c_949_n N_VPWR_c_950_n N_VPWR_c_951_n N_VPWR_c_952_n N_VPWR_c_953_n
+ N_VPWR_c_954_n N_VPWR_c_955_n VPWR N_VPWR_c_956_n N_VPWR_c_957_n
+ N_VPWR_c_958_n N_VPWR_c_959_n N_VPWR_c_960_n N_VPWR_c_961_n N_VPWR_c_962_n
+ N_VPWR_c_963_n N_VPWR_c_964_n N_VPWR_c_965_n N_VPWR_c_966_n N_VPWR_c_967_n
+ N_VPWR_c_925_n PM_SKY130_FD_SC_LP__BUFBUF_16%VPWR
x_PM_SKY130_FD_SC_LP__BUFBUF_16%X N_X_M1002_d N_X_M1009_d N_X_M1013_d
+ N_X_M1016_d N_X_M1028_d N_X_M1034_d N_X_M1043_d N_X_M1046_d N_X_M1000_d
+ N_X_M1005_d N_X_M1010_d N_X_M1017_d N_X_M1021_d N_X_M1031_d N_X_M1037_d
+ N_X_M1047_d X N_X_c_1158_n N_X_c_1159_n N_X_c_1160_n N_X_c_1161_n N_X_c_1162_n
+ N_X_c_1163_n N_X_c_1164_n N_X_c_1165_n N_X_c_1174_n
+ PM_SKY130_FD_SC_LP__BUFBUF_16%X
x_PM_SKY130_FD_SC_LP__BUFBUF_16%VGND N_VGND_M1018_d N_VGND_M1032_s
+ N_VGND_M1008_d N_VGND_M1011_d N_VGND_M1029_d N_VGND_M1035_d N_VGND_M1006_s
+ N_VGND_M1012_s N_VGND_M1014_s N_VGND_M1024_s N_VGND_M1030_s N_VGND_M1038_s
+ N_VGND_M1044_s N_VGND_M1049_s N_VGND_c_1343_n N_VGND_c_1344_n N_VGND_c_1345_n
+ N_VGND_c_1346_n N_VGND_c_1347_n N_VGND_c_1348_n N_VGND_c_1349_n
+ N_VGND_c_1350_n N_VGND_c_1351_n N_VGND_c_1352_n N_VGND_c_1353_n
+ N_VGND_c_1354_n N_VGND_c_1355_n N_VGND_c_1356_n N_VGND_c_1357_n
+ N_VGND_c_1358_n N_VGND_c_1359_n N_VGND_c_1360_n N_VGND_c_1361_n
+ N_VGND_c_1362_n N_VGND_c_1363_n N_VGND_c_1364_n N_VGND_c_1365_n
+ N_VGND_c_1366_n N_VGND_c_1367_n N_VGND_c_1368_n N_VGND_c_1369_n
+ N_VGND_c_1370_n N_VGND_c_1371_n N_VGND_c_1372_n VGND N_VGND_c_1373_n
+ N_VGND_c_1374_n N_VGND_c_1375_n N_VGND_c_1376_n N_VGND_c_1377_n
+ N_VGND_c_1378_n N_VGND_c_1379_n N_VGND_c_1380_n N_VGND_c_1381_n
+ N_VGND_c_1382_n N_VGND_c_1383_n N_VGND_c_1384_n N_VGND_c_1385_n
+ PM_SKY130_FD_SC_LP__BUFBUF_16%VGND
cc_1 VNB N_A_M1018_g 0.0277822f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.665
cc_2 VNB N_A_M1051_g 0.00183908f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_A_c_242_n 0.0501087f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.46
cc_4 VNB N_A_c_243_n 0.00111806f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.46
cc_5 VNB N_A_27_49#_M1027_g 0.0215698f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_27_49#_M1032_g 0.0213234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_49#_M1048_g 0.0272357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_49#_c_274_n 0.028851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_49#_c_275_n 0.00417409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_49#_c_276_n 0.0110786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_49#_c_277_n 0.0018632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_49#_c_278_n 3.82705e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_49#_c_279_n 0.00138602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_49#_c_280_n 0.0280517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_49#_c_281_n 0.00113095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_49#_c_282_n 0.0443924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_196_49#_M1008_g 0.0263182f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.625
cc_18 VNB N_A_196_49#_M1003_g 5.79352e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_196_49#_M1011_g 0.0214082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_196_49#_M1019_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_196_49#_M1023_g 0.021612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_196_49#_M1025_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_196_49#_M1029_g 0.021612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_196_49#_M1040_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_196_49#_M1033_g 0.0215915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_196_49#_M1041_g 4.57435e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_196_49#_M1035_g 0.0217944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_196_49#_M1042_g 4.70146e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_196_49#_c_386_n 0.00289786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_196_49#_c_387_n 0.00263148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_196_49#_c_388_n 0.0164558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_196_49#_c_389_n 0.0372629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_196_49#_c_390_n 0.00199211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_196_49#_c_391_n 0.00223187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_196_49#_c_392_n 0.131182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_610_47#_M1002_g 0.0217825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_610_47#_M1000_g 3.84315e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_610_47#_M1006_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_610_47#_M1004_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_610_47#_M1009_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_610_47#_M1005_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_610_47#_M1012_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_610_47#_M1007_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_610_47#_M1013_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_610_47#_M1010_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_610_47#_M1014_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_610_47#_M1015_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_610_47#_M1016_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_610_47#_M1017_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_610_47#_M1024_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_610_47#_M1020_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_610_47#_M1028_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_610_47#_M1021_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_610_47#_M1030_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_610_47#_M1026_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_610_47#_M1034_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_610_47#_M1031_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_610_47#_M1038_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_610_47#_M1036_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_610_47#_M1043_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_610_47#_M1037_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_610_47#_M1044_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_610_47#_M1045_g 3.84875e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_610_47#_M1046_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_610_47#_M1047_g 4.18354e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_610_47#_M1049_g 0.0324651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_610_47#_M1050_g 7.21331e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_610_47#_c_575_n 0.00272552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_610_47#_c_576_n 0.003138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_610_47#_c_577_n 0.00240399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_610_47#_c_578_n 0.00133064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_610_47#_c_579_n 0.00210048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_610_47#_c_580_n 0.00210048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_610_47#_c_581_n 0.00367436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_610_47#_c_582_n 0.00189682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_610_47#_c_583_n 0.00112451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_610_47#_c_584_n 0.00112451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_610_47#_c_585_n 0.00112451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_610_47#_c_586_n 0.00112451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_610_47#_c_587_n 0.00112451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_610_47#_c_588_n 0.00112451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_610_47#_c_589_n 0.00112451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_610_47#_c_590_n 0.339545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VPWR_c_925_n 0.521925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_X_c_1158_n 0.00387731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_X_c_1159_n 0.00450559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_X_c_1160_n 0.00450559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_X_c_1161_n 0.00450559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_X_c_1162_n 0.00450559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_X_c_1163_n 0.00450559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_X_c_1164_n 0.00450559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_X_c_1165_n 0.00491613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1343_n 6.09197e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1344_n 6.09197e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1345_n 0.0245316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1346_n 0.0154808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1347_n 0.00194604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1348_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1349_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1350_n 0.00530283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1351_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1352_n 0.00530283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1353_n 0.00530283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1354_n 0.00530283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1355_n 0.00530283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1356_n 0.00530283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1357_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1358_n 0.00530283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1359_n 0.0109056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1360_n 0.0467359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1361_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1362_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1363_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1364_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1365_n 0.0168376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1366_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1367_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1368_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1369_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1370_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1371_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1372_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1373_n 0.0154417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1374_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1375_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1376_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1377_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1378_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1379_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1380_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1381_n 0.00446109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1382_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1383_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1384_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1385_n 0.586406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VPB N_A_M1051_g 0.0263457f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_137 VPB N_A_c_243_n 0.00580632f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.46
cc_138 VPB N_A_27_49#_M1001_g 0.0190447f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.46
cc_139 VPB N_A_27_49#_M1022_g 0.0188982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_27_49#_M1039_g 0.0237962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_27_49#_c_286_n 0.00880428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_27_49#_c_287_n 0.0378753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_27_49#_c_278_n 0.00135782f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_27_49#_c_280_n 0.00793551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_27_49#_c_282_n 0.0046822f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_196_49#_M1003_g 0.0230769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_196_49#_M1019_g 0.0190295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_196_49#_M1025_g 0.0190295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_196_49#_M1040_g 0.0190295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_196_49#_M1041_g 0.0190093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_196_49#_M1042_g 0.0191959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_196_49#_c_399_n 0.00290581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_196_49#_c_400_n 0.00222593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_196_49#_c_401_n 0.0210267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_196_49#_c_402_n 0.0203304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_196_49#_c_390_n 0.00313916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_196_49#_c_404_n 0.00263594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_610_47#_M1000_g 0.0185778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_610_47#_M1004_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_610_47#_M1005_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_610_47#_M1007_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_610_47#_M1010_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_610_47#_M1015_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_610_47#_M1017_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_610_47#_M1020_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_610_47#_M1021_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_610_47#_M1026_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_610_47#_M1031_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_610_47#_M1036_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_610_47#_M1037_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_610_47#_M1045_g 0.0187835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_610_47#_M1047_g 0.0192485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_610_47#_M1050_g 0.0277364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_610_47#_c_607_n 0.00240637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_610_47#_c_608_n 0.00275727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_610_47#_c_609_n 0.00240637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_610_47#_c_610_n 0.00120085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_610_47#_c_611_n 0.00210048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_610_47#_c_612_n 0.00210048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_610_47#_c_581_n 0.00114059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_610_47#_c_582_n 0.0100817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_610_47#_c_583_n 0.00155931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_610_47#_c_584_n 0.00155931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_610_47#_c_585_n 0.00155931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_610_47#_c_586_n 0.00155931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_610_47#_c_587_n 0.00155931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_610_47#_c_588_n 0.00155931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_610_47#_c_589_n 0.00155931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_926_n 0.00457135f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_927_n 4.05231e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_928_n 0.0244658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_929_n 0.0189025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_930_n 0.00396563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_931_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_932_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_933_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_934_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_935_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_936_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_937_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_938_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_939_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_940_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_941_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_942_n 0.0108797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_943_n 0.0508715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_944_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_945_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_946_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_947_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_948_n 0.0168376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_949_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_950_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_951_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_952_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_953_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_954_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_955_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_956_n 0.0172072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_957_n 0.0149122f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_958_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_959_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_960_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_961_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_962_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_963_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_964_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_965_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_966_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_967_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_925_n 0.0644389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_X_c_1158_n 0.00181478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_X_c_1159_n 0.00208793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_X_c_1160_n 0.00208793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_X_c_1161_n 0.00208793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_X_c_1162_n 0.00208793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_X_c_1163_n 0.00208793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_X_c_1164_n 0.00208793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_X_c_1165_n 0.00284596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 N_A_M1018_g N_A_27_49#_M1027_g 0.0242054f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_241 N_A_M1051_g N_A_27_49#_M1001_g 0.0242054f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_242 N_A_c_242_n N_A_27_49#_c_286_n 0.00125014f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_243 N_A_c_243_n N_A_27_49#_c_286_n 0.0185329f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_244 N_A_M1018_g N_A_27_49#_c_275_n 0.0172632f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_245 N_A_c_242_n N_A_27_49#_c_275_n 0.00107988f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_246 N_A_c_243_n N_A_27_49#_c_275_n 0.00952576f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_247 N_A_c_242_n N_A_27_49#_c_276_n 0.00502923f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_248 N_A_c_243_n N_A_27_49#_c_276_n 0.0170721f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_249 N_A_M1051_g N_A_27_49#_c_300_n 0.0149592f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A_c_243_n N_A_27_49#_c_300_n 0.00651388f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_251 N_A_M1018_g N_A_27_49#_c_277_n 0.0041541f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_252 N_A_c_243_n N_A_27_49#_c_277_n 0.00356293f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_253 N_A_c_242_n N_A_27_49#_c_278_n 0.00477895f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_254 N_A_c_243_n N_A_27_49#_c_278_n 0.011445f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_255 N_A_c_242_n N_A_27_49#_c_281_n 0.00152518f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_256 N_A_c_243_n N_A_27_49#_c_281_n 0.0149428f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_257 N_A_c_242_n N_A_27_49#_c_282_n 0.0242054f $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_258 N_A_c_243_n N_A_27_49#_c_282_n 3.4989e-19 $X=0.32 $Y=1.46 $X2=0 $Y2=0
cc_259 N_A_M1051_g N_VPWR_c_926_n 0.00371643f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A_M1051_g N_VPWR_c_956_n 0.00585385f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A_M1051_g N_VPWR_c_925_n 0.0117692f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A_M1018_g N_VGND_c_1343_n 0.0117991f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_263 N_A_M1018_g N_VGND_c_1373_n 0.00477554f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_264 N_A_M1018_g N_VGND_c_1385_n 0.00919076f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_265 N_A_27_49#_M1032_g N_A_196_49#_c_386_n 0.0138902f $X=1.335 $Y=0.665 $X2=0
+ $Y2=0
cc_266 N_A_27_49#_M1048_g N_A_196_49#_c_386_n 0.0160847f $X=1.765 $Y=0.665 $X2=0
+ $Y2=0
cc_267 N_A_27_49#_c_279_n N_A_196_49#_c_386_n 0.0469885f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_268 N_A_27_49#_c_280_n N_A_196_49#_c_386_n 0.00108448f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_269 N_A_27_49#_c_282_n N_A_196_49#_c_386_n 0.00246472f $X=1.84 $Y=1.49 $X2=0
+ $Y2=0
cc_270 N_A_27_49#_M1027_g N_A_196_49#_c_387_n 0.00138043f $X=0.905 $Y=0.665
+ $X2=0 $Y2=0
cc_271 N_A_27_49#_c_275_n N_A_196_49#_c_387_n 0.00892235f $X=0.665 $Y=1.1 $X2=0
+ $Y2=0
cc_272 N_A_27_49#_c_277_n N_A_196_49#_c_387_n 0.00367961f $X=0.75 $Y=1.405 $X2=0
+ $Y2=0
cc_273 N_A_27_49#_c_279_n N_A_196_49#_c_387_n 0.0154155f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_274 N_A_27_49#_c_282_n N_A_196_49#_c_387_n 0.00256759f $X=1.84 $Y=1.49 $X2=0
+ $Y2=0
cc_275 N_A_27_49#_M1022_g N_A_196_49#_c_399_n 0.0134366f $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_276 N_A_27_49#_M1039_g N_A_196_49#_c_399_n 0.0144127f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_277 N_A_27_49#_c_279_n N_A_196_49#_c_399_n 0.0473012f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_278 N_A_27_49#_c_280_n N_A_196_49#_c_399_n 0.00106738f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_279 N_A_27_49#_c_282_n N_A_196_49#_c_399_n 0.00242587f $X=1.84 $Y=1.49 $X2=0
+ $Y2=0
cc_280 N_A_27_49#_M1001_g N_A_196_49#_c_400_n 6.41325e-19 $X=0.905 $Y=2.465
+ $X2=0 $Y2=0
cc_281 N_A_27_49#_c_278_n N_A_196_49#_c_400_n 0.00886392f $X=0.75 $Y=1.92 $X2=0
+ $Y2=0
cc_282 N_A_27_49#_c_279_n N_A_196_49#_c_400_n 0.0170387f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_283 N_A_27_49#_c_282_n N_A_196_49#_c_400_n 0.00252068f $X=1.84 $Y=1.49 $X2=0
+ $Y2=0
cc_284 N_A_27_49#_M1048_g N_A_196_49#_c_389_n 0.00286958f $X=1.765 $Y=0.665
+ $X2=0 $Y2=0
cc_285 N_A_27_49#_c_279_n N_A_196_49#_c_389_n 0.0182127f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_286 N_A_27_49#_c_280_n N_A_196_49#_c_389_n 0.00420971f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_287 N_A_27_49#_c_279_n N_A_196_49#_c_402_n 0.00248104f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_288 N_A_27_49#_c_280_n N_A_196_49#_c_402_n 8.44824e-19 $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_289 N_A_27_49#_M1039_g N_A_196_49#_c_390_n 0.00249373f $X=1.765 $Y=2.465
+ $X2=0 $Y2=0
cc_290 N_A_27_49#_c_280_n N_A_196_49#_c_390_n 0.00174797f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_291 N_A_27_49#_c_279_n N_A_196_49#_c_391_n 0.0210913f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_292 N_A_27_49#_c_280_n N_A_196_49#_c_391_n 0.00667574f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_293 N_A_27_49#_c_279_n N_A_196_49#_c_404_n 0.0210917f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_294 N_A_27_49#_c_280_n N_A_196_49#_c_404_n 0.00655377f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_295 N_A_27_49#_c_280_n N_A_196_49#_c_392_n 0.00468613f $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_296 N_A_27_49#_c_300_n N_VPWR_M1051_d 0.00396488f $X=0.665 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_297 N_A_27_49#_c_278_n N_VPWR_M1051_d 9.43676e-19 $X=0.75 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_298 N_A_27_49#_M1001_g N_VPWR_c_926_n 0.00220476f $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_299 N_A_27_49#_c_300_n N_VPWR_c_926_n 0.0143747f $X=0.665 $Y=2.005 $X2=0
+ $Y2=0
cc_300 N_A_27_49#_M1001_g N_VPWR_c_927_n 7.71921e-19 $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_301 N_A_27_49#_M1022_g N_VPWR_c_927_n 0.0140974f $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_A_27_49#_M1039_g N_VPWR_c_927_n 0.0159861f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_27_49#_M1039_g N_VPWR_c_928_n 0.00486043f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_304 N_A_27_49#_c_287_n N_VPWR_c_956_n 0.0190529f $X=0.26 $Y=2.865 $X2=0 $Y2=0
cc_305 N_A_27_49#_M1001_g N_VPWR_c_957_n 0.00585385f $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_306 N_A_27_49#_M1022_g N_VPWR_c_957_n 0.00486043f $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_27_49#_M1051_s N_VPWR_c_925_n 0.00254229f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_308 N_A_27_49#_M1001_g N_VPWR_c_925_n 0.0107648f $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_27_49#_M1022_g N_VPWR_c_925_n 0.00835506f $X=1.335 $Y=2.465 $X2=0
+ $Y2=0
cc_310 N_A_27_49#_M1039_g N_VPWR_c_925_n 0.00975473f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A_27_49#_c_287_n N_VPWR_c_925_n 0.0113912f $X=0.26 $Y=2.865 $X2=0 $Y2=0
cc_312 N_A_27_49#_c_275_n N_VGND_M1018_d 0.00180108f $X=0.665 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_313 N_A_27_49#_M1027_g N_VGND_c_1343_n 0.0103163f $X=0.905 $Y=0.665 $X2=0
+ $Y2=0
cc_314 N_A_27_49#_M1032_g N_VGND_c_1343_n 5.98801e-19 $X=1.335 $Y=0.665 $X2=0
+ $Y2=0
cc_315 N_A_27_49#_c_275_n N_VGND_c_1343_n 0.0165868f $X=0.665 $Y=1.1 $X2=0 $Y2=0
cc_316 N_A_27_49#_c_279_n N_VGND_c_1343_n 5.31672e-19 $X=2.015 $Y=1.49 $X2=0
+ $Y2=0
cc_317 N_A_27_49#_M1027_g N_VGND_c_1344_n 6.12946e-19 $X=0.905 $Y=0.665 $X2=0
+ $Y2=0
cc_318 N_A_27_49#_M1032_g N_VGND_c_1344_n 0.0106581f $X=1.335 $Y=0.665 $X2=0
+ $Y2=0
cc_319 N_A_27_49#_M1048_g N_VGND_c_1344_n 0.0123675f $X=1.765 $Y=0.665 $X2=0
+ $Y2=0
cc_320 N_A_27_49#_M1048_g N_VGND_c_1345_n 0.00477554f $X=1.765 $Y=0.665 $X2=0
+ $Y2=0
cc_321 N_A_27_49#_c_274_n N_VGND_c_1373_n 0.0178111f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_322 N_A_27_49#_M1027_g N_VGND_c_1374_n 0.00477554f $X=0.905 $Y=0.665 $X2=0
+ $Y2=0
cc_323 N_A_27_49#_M1032_g N_VGND_c_1374_n 0.00477554f $X=1.335 $Y=0.665 $X2=0
+ $Y2=0
cc_324 N_A_27_49#_M1018_s N_VGND_c_1385_n 0.00368844f $X=0.135 $Y=0.245 $X2=0
+ $Y2=0
cc_325 N_A_27_49#_M1027_g N_VGND_c_1385_n 0.00825815f $X=0.905 $Y=0.665 $X2=0
+ $Y2=0
cc_326 N_A_27_49#_M1032_g N_VGND_c_1385_n 0.00825815f $X=1.335 $Y=0.665 $X2=0
+ $Y2=0
cc_327 N_A_27_49#_M1048_g N_VGND_c_1385_n 0.00955784f $X=1.765 $Y=0.665 $X2=0
+ $Y2=0
cc_328 N_A_27_49#_c_274_n N_VGND_c_1385_n 0.0100304f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_329 N_A_196_49#_M1035_g N_A_610_47#_M1002_g 0.0211018f $X=5.125 $Y=0.655
+ $X2=0 $Y2=0
cc_330 N_A_196_49#_M1042_g N_A_610_47#_M1000_g 0.0211018f $X=5.125 $Y=2.465
+ $X2=0 $Y2=0
cc_331 N_A_196_49#_M1011_g N_A_610_47#_c_575_n 0.0138763f $X=3.405 $Y=0.655
+ $X2=0 $Y2=0
cc_332 N_A_196_49#_M1023_g N_A_610_47#_c_575_n 0.0148746f $X=3.835 $Y=0.655
+ $X2=0 $Y2=0
cc_333 N_A_196_49#_c_440_p N_A_610_47#_c_575_n 0.0445941f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_334 N_A_196_49#_c_392_n N_A_610_47#_c_575_n 0.00243542f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_335 N_A_196_49#_M1008_g N_A_610_47#_c_576_n 0.00144226f $X=2.975 $Y=0.655
+ $X2=0 $Y2=0
cc_336 N_A_196_49#_c_389_n N_A_610_47#_c_576_n 0.0112954f $X=2.35 $Y=1.15 $X2=0
+ $Y2=0
cc_337 N_A_196_49#_c_440_p N_A_610_47#_c_576_n 0.0186942f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_338 N_A_196_49#_c_392_n N_A_610_47#_c_576_n 0.00253619f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_339 N_A_196_49#_M1019_g N_A_610_47#_c_607_n 0.0142895f $X=3.405 $Y=2.465
+ $X2=0 $Y2=0
cc_340 N_A_196_49#_M1025_g N_A_610_47#_c_607_n 0.0145185f $X=3.835 $Y=2.465
+ $X2=0 $Y2=0
cc_341 N_A_196_49#_c_440_p N_A_610_47#_c_607_n 0.0422575f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_342 N_A_196_49#_c_392_n N_A_610_47#_c_607_n 0.00243878f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_343 N_A_196_49#_M1003_g N_A_610_47#_c_608_n 0.00144677f $X=2.975 $Y=2.465
+ $X2=0 $Y2=0
cc_344 N_A_196_49#_c_402_n N_A_610_47#_c_608_n 0.00474293f $X=2.35 $Y=1.845
+ $X2=0 $Y2=0
cc_345 N_A_196_49#_c_390_n N_A_610_47#_c_608_n 5.20639e-19 $X=2.435 $Y=1.76
+ $X2=0 $Y2=0
cc_346 N_A_196_49#_c_440_p N_A_610_47#_c_608_n 0.0182878f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_347 N_A_196_49#_c_392_n N_A_610_47#_c_608_n 0.00253619f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_348 N_A_196_49#_M1029_g N_A_610_47#_c_577_n 0.0149212f $X=4.265 $Y=0.655
+ $X2=0 $Y2=0
cc_349 N_A_196_49#_M1033_g N_A_610_47#_c_577_n 0.0149212f $X=4.695 $Y=0.655
+ $X2=0 $Y2=0
cc_350 N_A_196_49#_c_440_p N_A_610_47#_c_577_n 0.0420697f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_351 N_A_196_49#_c_392_n N_A_610_47#_c_577_n 0.00243542f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_352 N_A_196_49#_M1040_g N_A_610_47#_c_609_n 0.0145678f $X=4.265 $Y=2.465
+ $X2=0 $Y2=0
cc_353 N_A_196_49#_M1041_g N_A_610_47#_c_609_n 0.0145678f $X=4.695 $Y=2.465
+ $X2=0 $Y2=0
cc_354 N_A_196_49#_c_440_p N_A_610_47#_c_609_n 0.0422575f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_355 N_A_196_49#_c_392_n N_A_610_47#_c_609_n 0.00243878f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_356 N_A_196_49#_M1035_g N_A_610_47#_c_578_n 0.015598f $X=5.125 $Y=0.655 $X2=0
+ $Y2=0
cc_357 N_A_196_49#_c_440_p N_A_610_47#_c_578_n 0.00649467f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_358 N_A_196_49#_M1042_g N_A_610_47#_c_610_n 0.0151929f $X=5.125 $Y=2.465
+ $X2=0 $Y2=0
cc_359 N_A_196_49#_c_440_p N_A_610_47#_c_610_n 0.00652308f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_360 N_A_196_49#_c_440_p N_A_610_47#_c_579_n 0.021133f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_361 N_A_196_49#_c_392_n N_A_610_47#_c_579_n 0.00253619f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_362 N_A_196_49#_c_440_p N_A_610_47#_c_611_n 0.021133f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_363 N_A_196_49#_c_392_n N_A_610_47#_c_611_n 0.00253619f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_364 N_A_196_49#_c_440_p N_A_610_47#_c_580_n 0.021133f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_365 N_A_196_49#_c_392_n N_A_610_47#_c_580_n 0.00253619f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_366 N_A_196_49#_c_440_p N_A_610_47#_c_612_n 0.021133f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_367 N_A_196_49#_c_392_n N_A_610_47#_c_612_n 0.00253619f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_368 N_A_196_49#_M1035_g N_A_610_47#_c_581_n 0.00889731f $X=5.125 $Y=0.655
+ $X2=0 $Y2=0
cc_369 N_A_196_49#_c_440_p N_A_610_47#_c_581_n 0.0148694f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_370 N_A_196_49#_c_440_p N_A_610_47#_c_582_n 8.54896e-19 $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_371 N_A_196_49#_c_392_n N_A_610_47#_c_582_n 0.00428664f $X=5.125 $Y=1.48
+ $X2=0 $Y2=0
cc_372 N_A_196_49#_c_392_n N_A_610_47#_c_590_n 0.0211018f $X=5.125 $Y=1.48 $X2=0
+ $Y2=0
cc_373 N_A_196_49#_c_399_n N_VPWR_M1022_d 0.00176922f $X=1.885 $Y=1.852 $X2=0
+ $Y2=0
cc_374 N_A_196_49#_c_399_n N_VPWR_c_927_n 0.0171764f $X=1.885 $Y=1.852 $X2=0
+ $Y2=0
cc_375 N_A_196_49#_c_401_n N_VPWR_c_928_n 0.0178111f $X=1.98 $Y=2.025 $X2=0
+ $Y2=0
cc_376 N_A_196_49#_M1003_g N_VPWR_c_929_n 0.0156017f $X=2.975 $Y=2.465 $X2=0
+ $Y2=0
cc_377 N_A_196_49#_M1019_g N_VPWR_c_929_n 7.65361e-19 $X=3.405 $Y=2.465 $X2=0
+ $Y2=0
cc_378 N_A_196_49#_c_401_n N_VPWR_c_929_n 0.0407018f $X=1.98 $Y=2.025 $X2=0
+ $Y2=0
cc_379 N_A_196_49#_c_389_n N_VPWR_c_929_n 0.00974611f $X=2.35 $Y=1.15 $X2=0
+ $Y2=0
cc_380 N_A_196_49#_c_440_p N_VPWR_c_929_n 0.00133115f $X=4.97 $Y=1.48 $X2=0
+ $Y2=0
cc_381 N_A_196_49#_c_392_n N_VPWR_c_929_n 0.00241065f $X=5.125 $Y=1.48 $X2=0
+ $Y2=0
cc_382 N_A_196_49#_M1019_g N_VPWR_c_930_n 0.00158567f $X=3.405 $Y=2.465 $X2=0
+ $Y2=0
cc_383 N_A_196_49#_M1025_g N_VPWR_c_930_n 0.0016342f $X=3.835 $Y=2.465 $X2=0
+ $Y2=0
cc_384 N_A_196_49#_M1040_g N_VPWR_c_931_n 0.0016342f $X=4.265 $Y=2.465 $X2=0
+ $Y2=0
cc_385 N_A_196_49#_M1041_g N_VPWR_c_931_n 0.0016342f $X=4.695 $Y=2.465 $X2=0
+ $Y2=0
cc_386 N_A_196_49#_M1042_g N_VPWR_c_932_n 0.0016342f $X=5.125 $Y=2.465 $X2=0
+ $Y2=0
cc_387 N_A_196_49#_M1025_g N_VPWR_c_944_n 0.00585385f $X=3.835 $Y=2.465 $X2=0
+ $Y2=0
cc_388 N_A_196_49#_M1040_g N_VPWR_c_944_n 0.00585385f $X=4.265 $Y=2.465 $X2=0
+ $Y2=0
cc_389 N_A_196_49#_M1041_g N_VPWR_c_946_n 0.00585385f $X=4.695 $Y=2.465 $X2=0
+ $Y2=0
cc_390 N_A_196_49#_M1042_g N_VPWR_c_946_n 0.00585385f $X=5.125 $Y=2.465 $X2=0
+ $Y2=0
cc_391 N_A_196_49#_c_498_p N_VPWR_c_957_n 0.0131621f $X=1.12 $Y=2.025 $X2=0
+ $Y2=0
cc_392 N_A_196_49#_M1003_g N_VPWR_c_958_n 0.00486043f $X=2.975 $Y=2.465 $X2=0
+ $Y2=0
cc_393 N_A_196_49#_M1019_g N_VPWR_c_958_n 0.00585385f $X=3.405 $Y=2.465 $X2=0
+ $Y2=0
cc_394 N_A_196_49#_M1001_s N_VPWR_c_925_n 0.00475637f $X=0.98 $Y=1.835 $X2=0
+ $Y2=0
cc_395 N_A_196_49#_M1039_s N_VPWR_c_925_n 0.00375985f $X=1.84 $Y=1.835 $X2=0
+ $Y2=0
cc_396 N_A_196_49#_M1003_g N_VPWR_c_925_n 0.00835506f $X=2.975 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_A_196_49#_M1019_g N_VPWR_c_925_n 0.0106302f $X=3.405 $Y=2.465 $X2=0
+ $Y2=0
cc_398 N_A_196_49#_M1025_g N_VPWR_c_925_n 0.0106302f $X=3.835 $Y=2.465 $X2=0
+ $Y2=0
cc_399 N_A_196_49#_M1040_g N_VPWR_c_925_n 0.0106302f $X=4.265 $Y=2.465 $X2=0
+ $Y2=0
cc_400 N_A_196_49#_M1041_g N_VPWR_c_925_n 0.0106302f $X=4.695 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_A_196_49#_M1042_g N_VPWR_c_925_n 0.0106555f $X=5.125 $Y=2.465 $X2=0
+ $Y2=0
cc_402 N_A_196_49#_c_498_p N_VPWR_c_925_n 0.00808656f $X=1.12 $Y=2.025 $X2=0
+ $Y2=0
cc_403 N_A_196_49#_c_401_n N_VPWR_c_925_n 0.0100304f $X=1.98 $Y=2.025 $X2=0
+ $Y2=0
cc_404 N_A_196_49#_M1042_g N_X_c_1174_n 7.3936e-19 $X=5.125 $Y=2.465 $X2=0 $Y2=0
cc_405 N_A_196_49#_c_386_n N_VGND_M1032_s 0.00176461f $X=1.885 $Y=1.15 $X2=0
+ $Y2=0
cc_406 N_A_196_49#_c_389_n N_VGND_M1008_d 0.0023968f $X=2.35 $Y=1.15 $X2=0 $Y2=0
cc_407 N_A_196_49#_c_386_n N_VGND_c_1344_n 0.0170777f $X=1.885 $Y=1.15 $X2=0
+ $Y2=0
cc_408 N_A_196_49#_c_388_n N_VGND_c_1345_n 0.0178111f $X=1.98 $Y=0.42 $X2=0
+ $Y2=0
cc_409 N_A_196_49#_M1008_g N_VGND_c_1346_n 0.0033589f $X=2.975 $Y=0.655 $X2=0
+ $Y2=0
cc_410 N_A_196_49#_c_388_n N_VGND_c_1346_n 0.0264537f $X=1.98 $Y=0.42 $X2=0
+ $Y2=0
cc_411 N_A_196_49#_c_389_n N_VGND_c_1346_n 0.0219388f $X=2.35 $Y=1.15 $X2=0
+ $Y2=0
cc_412 N_A_196_49#_c_392_n N_VGND_c_1346_n 3.8292e-19 $X=5.125 $Y=1.48 $X2=0
+ $Y2=0
cc_413 N_A_196_49#_M1008_g N_VGND_c_1347_n 6.7553e-19 $X=2.975 $Y=0.655 $X2=0
+ $Y2=0
cc_414 N_A_196_49#_M1011_g N_VGND_c_1347_n 0.0104076f $X=3.405 $Y=0.655 $X2=0
+ $Y2=0
cc_415 N_A_196_49#_M1023_g N_VGND_c_1347_n 0.00165155f $X=3.835 $Y=0.655 $X2=0
+ $Y2=0
cc_416 N_A_196_49#_M1029_g N_VGND_c_1348_n 0.0016342f $X=4.265 $Y=0.655 $X2=0
+ $Y2=0
cc_417 N_A_196_49#_M1033_g N_VGND_c_1348_n 0.0016342f $X=4.695 $Y=0.655 $X2=0
+ $Y2=0
cc_418 N_A_196_49#_M1035_g N_VGND_c_1349_n 0.0016342f $X=5.125 $Y=0.655 $X2=0
+ $Y2=0
cc_419 N_A_196_49#_M1023_g N_VGND_c_1361_n 0.00585385f $X=3.835 $Y=0.655 $X2=0
+ $Y2=0
cc_420 N_A_196_49#_M1029_g N_VGND_c_1361_n 0.00585385f $X=4.265 $Y=0.655 $X2=0
+ $Y2=0
cc_421 N_A_196_49#_M1033_g N_VGND_c_1363_n 0.00585385f $X=4.695 $Y=0.655 $X2=0
+ $Y2=0
cc_422 N_A_196_49#_M1035_g N_VGND_c_1363_n 0.00585385f $X=5.125 $Y=0.655 $X2=0
+ $Y2=0
cc_423 N_A_196_49#_c_530_p N_VGND_c_1374_n 0.0124525f $X=1.12 $Y=0.42 $X2=0
+ $Y2=0
cc_424 N_A_196_49#_M1008_g N_VGND_c_1375_n 0.00585385f $X=2.975 $Y=0.655 $X2=0
+ $Y2=0
cc_425 N_A_196_49#_M1011_g N_VGND_c_1375_n 0.00486043f $X=3.405 $Y=0.655 $X2=0
+ $Y2=0
cc_426 N_A_196_49#_M1027_d N_VGND_c_1385_n 0.00536646f $X=0.98 $Y=0.245 $X2=0
+ $Y2=0
cc_427 N_A_196_49#_M1048_d N_VGND_c_1385_n 0.00368844f $X=1.84 $Y=0.245 $X2=0
+ $Y2=0
cc_428 N_A_196_49#_M1008_g N_VGND_c_1385_n 0.0119436f $X=2.975 $Y=0.655 $X2=0
+ $Y2=0
cc_429 N_A_196_49#_M1011_g N_VGND_c_1385_n 0.00835506f $X=3.405 $Y=0.655 $X2=0
+ $Y2=0
cc_430 N_A_196_49#_M1023_g N_VGND_c_1385_n 0.0106302f $X=3.835 $Y=0.655 $X2=0
+ $Y2=0
cc_431 N_A_196_49#_M1029_g N_VGND_c_1385_n 0.0106302f $X=4.265 $Y=0.655 $X2=0
+ $Y2=0
cc_432 N_A_196_49#_M1033_g N_VGND_c_1385_n 0.0106302f $X=4.695 $Y=0.655 $X2=0
+ $Y2=0
cc_433 N_A_196_49#_M1035_g N_VGND_c_1385_n 0.0106555f $X=5.125 $Y=0.655 $X2=0
+ $Y2=0
cc_434 N_A_196_49#_c_530_p N_VGND_c_1385_n 0.00730901f $X=1.12 $Y=0.42 $X2=0
+ $Y2=0
cc_435 N_A_196_49#_c_388_n N_VGND_c_1385_n 0.0100304f $X=1.98 $Y=0.42 $X2=0
+ $Y2=0
cc_436 N_A_610_47#_c_607_n N_VPWR_M1019_s 0.00176773f $X=3.92 $Y=1.835 $X2=0
+ $Y2=0
cc_437 N_A_610_47#_c_609_n N_VPWR_M1040_s 0.00176773f $X=4.78 $Y=1.835 $X2=0
+ $Y2=0
cc_438 N_A_610_47#_c_610_n N_VPWR_M1042_s 0.00180632f $X=5.305 $Y=1.835 $X2=0
+ $Y2=0
cc_439 N_A_610_47#_c_607_n N_VPWR_c_930_n 0.0135577f $X=3.92 $Y=1.835 $X2=0
+ $Y2=0
cc_440 N_A_610_47#_c_609_n N_VPWR_c_931_n 0.0135577f $X=4.78 $Y=1.835 $X2=0
+ $Y2=0
cc_441 N_A_610_47#_M1000_g N_VPWR_c_932_n 0.0016342f $X=5.555 $Y=2.465 $X2=0
+ $Y2=0
cc_442 N_A_610_47#_c_610_n N_VPWR_c_932_n 0.0135581f $X=5.305 $Y=1.835 $X2=0
+ $Y2=0
cc_443 N_A_610_47#_c_582_n N_VPWR_c_932_n 0.0012888f $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_444 N_A_610_47#_M1004_g N_VPWR_c_933_n 0.00211386f $X=5.985 $Y=2.465 $X2=0
+ $Y2=0
cc_445 N_A_610_47#_M1005_g N_VPWR_c_933_n 0.00211386f $X=6.415 $Y=2.465 $X2=0
+ $Y2=0
cc_446 N_A_610_47#_c_582_n N_VPWR_c_933_n 8.57152e-19 $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_447 N_A_610_47#_c_583_n N_VPWR_c_933_n 0.0171417f $X=6.2 $Y=1.48 $X2=0 $Y2=0
cc_448 N_A_610_47#_c_590_n N_VPWR_c_933_n 5.09955e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_449 N_A_610_47#_M1005_g N_VPWR_c_934_n 0.00585385f $X=6.415 $Y=2.465 $X2=0
+ $Y2=0
cc_450 N_A_610_47#_M1007_g N_VPWR_c_934_n 0.00585385f $X=6.845 $Y=2.465 $X2=0
+ $Y2=0
cc_451 N_A_610_47#_M1007_g N_VPWR_c_935_n 0.00211386f $X=6.845 $Y=2.465 $X2=0
+ $Y2=0
cc_452 N_A_610_47#_M1010_g N_VPWR_c_935_n 0.00211386f $X=7.275 $Y=2.465 $X2=0
+ $Y2=0
cc_453 N_A_610_47#_c_582_n N_VPWR_c_935_n 8.57152e-19 $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_454 N_A_610_47#_c_584_n N_VPWR_c_935_n 0.0171417f $X=7.06 $Y=1.48 $X2=0 $Y2=0
cc_455 N_A_610_47#_c_590_n N_VPWR_c_935_n 5.09955e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_456 N_A_610_47#_M1015_g N_VPWR_c_936_n 0.00211386f $X=7.705 $Y=2.465 $X2=0
+ $Y2=0
cc_457 N_A_610_47#_M1017_g N_VPWR_c_936_n 0.00211386f $X=8.135 $Y=2.465 $X2=0
+ $Y2=0
cc_458 N_A_610_47#_c_582_n N_VPWR_c_936_n 8.57152e-19 $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_459 N_A_610_47#_c_585_n N_VPWR_c_936_n 0.0171417f $X=7.92 $Y=1.48 $X2=0 $Y2=0
cc_460 N_A_610_47#_c_590_n N_VPWR_c_936_n 5.09955e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_461 N_A_610_47#_M1020_g N_VPWR_c_937_n 0.00211386f $X=8.565 $Y=2.465 $X2=0
+ $Y2=0
cc_462 N_A_610_47#_M1021_g N_VPWR_c_937_n 0.00211386f $X=8.995 $Y=2.465 $X2=0
+ $Y2=0
cc_463 N_A_610_47#_c_582_n N_VPWR_c_937_n 8.57152e-19 $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_464 N_A_610_47#_c_586_n N_VPWR_c_937_n 0.0171417f $X=8.78 $Y=1.48 $X2=0 $Y2=0
cc_465 N_A_610_47#_c_590_n N_VPWR_c_937_n 5.09955e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_466 N_A_610_47#_M1026_g N_VPWR_c_938_n 0.00211386f $X=9.425 $Y=2.465 $X2=0
+ $Y2=0
cc_467 N_A_610_47#_M1031_g N_VPWR_c_938_n 0.00211386f $X=9.855 $Y=2.465 $X2=0
+ $Y2=0
cc_468 N_A_610_47#_c_582_n N_VPWR_c_938_n 8.57152e-19 $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_469 N_A_610_47#_c_587_n N_VPWR_c_938_n 0.0171417f $X=9.64 $Y=1.48 $X2=0 $Y2=0
cc_470 N_A_610_47#_c_590_n N_VPWR_c_938_n 5.09955e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_471 N_A_610_47#_M1036_g N_VPWR_c_939_n 0.00211386f $X=10.285 $Y=2.465 $X2=0
+ $Y2=0
cc_472 N_A_610_47#_M1037_g N_VPWR_c_939_n 0.00211386f $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_473 N_A_610_47#_c_582_n N_VPWR_c_939_n 8.57152e-19 $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_474 N_A_610_47#_c_588_n N_VPWR_c_939_n 0.0171417f $X=10.5 $Y=1.48 $X2=0 $Y2=0
cc_475 N_A_610_47#_c_590_n N_VPWR_c_939_n 5.09955e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_476 N_A_610_47#_M1037_g N_VPWR_c_940_n 0.00585385f $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_477 N_A_610_47#_M1045_g N_VPWR_c_940_n 0.00585385f $X=11.145 $Y=2.465 $X2=0
+ $Y2=0
cc_478 N_A_610_47#_M1045_g N_VPWR_c_941_n 0.00211386f $X=11.145 $Y=2.465 $X2=0
+ $Y2=0
cc_479 N_A_610_47#_M1047_g N_VPWR_c_941_n 0.00211386f $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_480 N_A_610_47#_c_582_n N_VPWR_c_941_n 8.57152e-19 $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_481 N_A_610_47#_c_589_n N_VPWR_c_941_n 0.0171417f $X=11.36 $Y=1.48 $X2=0
+ $Y2=0
cc_482 N_A_610_47#_c_590_n N_VPWR_c_941_n 5.09955e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_483 N_A_610_47#_M1050_g N_VPWR_c_943_n 0.00414232f $X=12.005 $Y=2.465 $X2=0
+ $Y2=0
cc_484 N_A_610_47#_c_714_p N_VPWR_c_944_n 0.0149362f $X=4.05 $Y=2.045 $X2=0
+ $Y2=0
cc_485 N_A_610_47#_c_715_p N_VPWR_c_946_n 0.0149362f $X=4.91 $Y=2.045 $X2=0
+ $Y2=0
cc_486 N_A_610_47#_M1000_g N_VPWR_c_948_n 0.00585385f $X=5.555 $Y=2.465 $X2=0
+ $Y2=0
cc_487 N_A_610_47#_M1004_g N_VPWR_c_948_n 0.00585385f $X=5.985 $Y=2.465 $X2=0
+ $Y2=0
cc_488 N_A_610_47#_M1017_g N_VPWR_c_950_n 0.00585385f $X=8.135 $Y=2.465 $X2=0
+ $Y2=0
cc_489 N_A_610_47#_M1020_g N_VPWR_c_950_n 0.00585385f $X=8.565 $Y=2.465 $X2=0
+ $Y2=0
cc_490 N_A_610_47#_M1021_g N_VPWR_c_952_n 0.00585385f $X=8.995 $Y=2.465 $X2=0
+ $Y2=0
cc_491 N_A_610_47#_M1026_g N_VPWR_c_952_n 0.00585385f $X=9.425 $Y=2.465 $X2=0
+ $Y2=0
cc_492 N_A_610_47#_M1031_g N_VPWR_c_954_n 0.00585385f $X=9.855 $Y=2.465 $X2=0
+ $Y2=0
cc_493 N_A_610_47#_M1036_g N_VPWR_c_954_n 0.00585385f $X=10.285 $Y=2.465 $X2=0
+ $Y2=0
cc_494 N_A_610_47#_c_724_p N_VPWR_c_958_n 0.0136943f $X=3.19 $Y=2.045 $X2=0
+ $Y2=0
cc_495 N_A_610_47#_M1010_g N_VPWR_c_959_n 0.00585385f $X=7.275 $Y=2.465 $X2=0
+ $Y2=0
cc_496 N_A_610_47#_M1015_g N_VPWR_c_959_n 0.00585385f $X=7.705 $Y=2.465 $X2=0
+ $Y2=0
cc_497 N_A_610_47#_M1047_g N_VPWR_c_960_n 0.00585385f $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_498 N_A_610_47#_M1050_g N_VPWR_c_960_n 0.00585385f $X=12.005 $Y=2.465 $X2=0
+ $Y2=0
cc_499 N_A_610_47#_M1003_d N_VPWR_c_925_n 0.00423456f $X=3.05 $Y=1.835 $X2=0
+ $Y2=0
cc_500 N_A_610_47#_M1025_d N_VPWR_c_925_n 0.003017f $X=3.91 $Y=1.835 $X2=0 $Y2=0
cc_501 N_A_610_47#_M1041_d N_VPWR_c_925_n 0.003017f $X=4.77 $Y=1.835 $X2=0 $Y2=0
cc_502 N_A_610_47#_M1000_g N_VPWR_c_925_n 0.0106555f $X=5.555 $Y=2.465 $X2=0
+ $Y2=0
cc_503 N_A_610_47#_M1004_g N_VPWR_c_925_n 0.0106302f $X=5.985 $Y=2.465 $X2=0
+ $Y2=0
cc_504 N_A_610_47#_M1005_g N_VPWR_c_925_n 0.0106302f $X=6.415 $Y=2.465 $X2=0
+ $Y2=0
cc_505 N_A_610_47#_M1007_g N_VPWR_c_925_n 0.0106302f $X=6.845 $Y=2.465 $X2=0
+ $Y2=0
cc_506 N_A_610_47#_M1010_g N_VPWR_c_925_n 0.0106302f $X=7.275 $Y=2.465 $X2=0
+ $Y2=0
cc_507 N_A_610_47#_M1015_g N_VPWR_c_925_n 0.0106302f $X=7.705 $Y=2.465 $X2=0
+ $Y2=0
cc_508 N_A_610_47#_M1017_g N_VPWR_c_925_n 0.0106302f $X=8.135 $Y=2.465 $X2=0
+ $Y2=0
cc_509 N_A_610_47#_M1020_g N_VPWR_c_925_n 0.0106302f $X=8.565 $Y=2.465 $X2=0
+ $Y2=0
cc_510 N_A_610_47#_M1021_g N_VPWR_c_925_n 0.0106302f $X=8.995 $Y=2.465 $X2=0
+ $Y2=0
cc_511 N_A_610_47#_M1026_g N_VPWR_c_925_n 0.0106302f $X=9.425 $Y=2.465 $X2=0
+ $Y2=0
cc_512 N_A_610_47#_M1031_g N_VPWR_c_925_n 0.0106302f $X=9.855 $Y=2.465 $X2=0
+ $Y2=0
cc_513 N_A_610_47#_M1036_g N_VPWR_c_925_n 0.0106302f $X=10.285 $Y=2.465 $X2=0
+ $Y2=0
cc_514 N_A_610_47#_M1037_g N_VPWR_c_925_n 0.0106302f $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_515 N_A_610_47#_M1045_g N_VPWR_c_925_n 0.0106302f $X=11.145 $Y=2.465 $X2=0
+ $Y2=0
cc_516 N_A_610_47#_M1047_g N_VPWR_c_925_n 0.0104456f $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_517 N_A_610_47#_M1050_g N_VPWR_c_925_n 0.0115628f $X=12.005 $Y=2.465 $X2=0
+ $Y2=0
cc_518 N_A_610_47#_c_724_p N_VPWR_c_925_n 0.00866972f $X=3.19 $Y=2.045 $X2=0
+ $Y2=0
cc_519 N_A_610_47#_c_714_p N_VPWR_c_925_n 0.0100304f $X=4.05 $Y=2.045 $X2=0
+ $Y2=0
cc_520 N_A_610_47#_c_715_p N_VPWR_c_925_n 0.0100304f $X=4.91 $Y=2.045 $X2=0
+ $Y2=0
cc_521 N_A_610_47#_M1002_g N_X_c_1158_n 0.00196849f $X=5.555 $Y=0.655 $X2=0
+ $Y2=0
cc_522 N_A_610_47#_M1000_g N_X_c_1158_n 0.00235242f $X=5.555 $Y=2.465 $X2=0
+ $Y2=0
cc_523 N_A_610_47#_M1006_g N_X_c_1158_n 0.00357508f $X=5.985 $Y=0.655 $X2=0
+ $Y2=0
cc_524 N_A_610_47#_M1004_g N_X_c_1158_n 0.00250971f $X=5.985 $Y=2.465 $X2=0
+ $Y2=0
cc_525 N_A_610_47#_c_578_n N_X_c_1158_n 0.0126773f $X=5.305 $Y=1.13 $X2=0 $Y2=0
cc_526 N_A_610_47#_c_610_n N_X_c_1158_n 0.0107091f $X=5.305 $Y=1.835 $X2=0 $Y2=0
cc_527 N_A_610_47#_c_581_n N_X_c_1158_n 0.0367603f $X=5.4 $Y=1.665 $X2=0 $Y2=0
cc_528 N_A_610_47#_c_582_n N_X_c_1158_n 0.0268818f $X=11.36 $Y=1.665 $X2=0 $Y2=0
cc_529 N_A_610_47#_c_583_n N_X_c_1158_n 0.030908f $X=6.2 $Y=1.48 $X2=0 $Y2=0
cc_530 N_A_610_47#_c_590_n N_X_c_1158_n 0.0199484f $X=12.005 $Y=1.48 $X2=0 $Y2=0
cc_531 N_A_610_47#_M1009_g N_X_c_1159_n 0.00362883f $X=6.415 $Y=0.655 $X2=0
+ $Y2=0
cc_532 N_A_610_47#_M1005_g N_X_c_1159_n 0.00253248f $X=6.415 $Y=2.465 $X2=0
+ $Y2=0
cc_533 N_A_610_47#_M1012_g N_X_c_1159_n 0.00362883f $X=6.845 $Y=0.655 $X2=0
+ $Y2=0
cc_534 N_A_610_47#_M1007_g N_X_c_1159_n 0.00253248f $X=6.845 $Y=2.465 $X2=0
+ $Y2=0
cc_535 N_A_610_47#_c_582_n N_X_c_1159_n 0.029632f $X=11.36 $Y=1.665 $X2=0 $Y2=0
cc_536 N_A_610_47#_c_583_n N_X_c_1159_n 0.0310539f $X=6.2 $Y=1.48 $X2=0 $Y2=0
cc_537 N_A_610_47#_c_584_n N_X_c_1159_n 0.0310539f $X=7.06 $Y=1.48 $X2=0 $Y2=0
cc_538 N_A_610_47#_c_590_n N_X_c_1159_n 0.0209262f $X=12.005 $Y=1.48 $X2=0 $Y2=0
cc_539 N_A_610_47#_M1013_g N_X_c_1160_n 0.00362883f $X=7.275 $Y=0.655 $X2=0
+ $Y2=0
cc_540 N_A_610_47#_M1010_g N_X_c_1160_n 0.00253248f $X=7.275 $Y=2.465 $X2=0
+ $Y2=0
cc_541 N_A_610_47#_M1014_g N_X_c_1160_n 0.00362883f $X=7.705 $Y=0.655 $X2=0
+ $Y2=0
cc_542 N_A_610_47#_M1015_g N_X_c_1160_n 0.00253248f $X=7.705 $Y=2.465 $X2=0
+ $Y2=0
cc_543 N_A_610_47#_c_582_n N_X_c_1160_n 0.029632f $X=11.36 $Y=1.665 $X2=0 $Y2=0
cc_544 N_A_610_47#_c_584_n N_X_c_1160_n 0.0310539f $X=7.06 $Y=1.48 $X2=0 $Y2=0
cc_545 N_A_610_47#_c_585_n N_X_c_1160_n 0.0310539f $X=7.92 $Y=1.48 $X2=0 $Y2=0
cc_546 N_A_610_47#_c_590_n N_X_c_1160_n 0.0209262f $X=12.005 $Y=1.48 $X2=0 $Y2=0
cc_547 N_A_610_47#_M1016_g N_X_c_1161_n 0.00362883f $X=8.135 $Y=0.655 $X2=0
+ $Y2=0
cc_548 N_A_610_47#_M1017_g N_X_c_1161_n 0.00253248f $X=8.135 $Y=2.465 $X2=0
+ $Y2=0
cc_549 N_A_610_47#_M1024_g N_X_c_1161_n 0.00362883f $X=8.565 $Y=0.655 $X2=0
+ $Y2=0
cc_550 N_A_610_47#_M1020_g N_X_c_1161_n 0.00253248f $X=8.565 $Y=2.465 $X2=0
+ $Y2=0
cc_551 N_A_610_47#_c_582_n N_X_c_1161_n 0.029632f $X=11.36 $Y=1.665 $X2=0 $Y2=0
cc_552 N_A_610_47#_c_585_n N_X_c_1161_n 0.0310539f $X=7.92 $Y=1.48 $X2=0 $Y2=0
cc_553 N_A_610_47#_c_586_n N_X_c_1161_n 0.0310539f $X=8.78 $Y=1.48 $X2=0 $Y2=0
cc_554 N_A_610_47#_c_590_n N_X_c_1161_n 0.0209262f $X=12.005 $Y=1.48 $X2=0 $Y2=0
cc_555 N_A_610_47#_M1028_g N_X_c_1162_n 0.00362883f $X=8.995 $Y=0.655 $X2=0
+ $Y2=0
cc_556 N_A_610_47#_M1021_g N_X_c_1162_n 0.00253248f $X=8.995 $Y=2.465 $X2=0
+ $Y2=0
cc_557 N_A_610_47#_M1030_g N_X_c_1162_n 0.00362883f $X=9.425 $Y=0.655 $X2=0
+ $Y2=0
cc_558 N_A_610_47#_M1026_g N_X_c_1162_n 0.00253248f $X=9.425 $Y=2.465 $X2=0
+ $Y2=0
cc_559 N_A_610_47#_c_582_n N_X_c_1162_n 0.029632f $X=11.36 $Y=1.665 $X2=0 $Y2=0
cc_560 N_A_610_47#_c_586_n N_X_c_1162_n 0.0310539f $X=8.78 $Y=1.48 $X2=0 $Y2=0
cc_561 N_A_610_47#_c_587_n N_X_c_1162_n 0.0310539f $X=9.64 $Y=1.48 $X2=0 $Y2=0
cc_562 N_A_610_47#_c_590_n N_X_c_1162_n 0.0209262f $X=12.005 $Y=1.48 $X2=0 $Y2=0
cc_563 N_A_610_47#_M1034_g N_X_c_1163_n 0.00362883f $X=9.855 $Y=0.655 $X2=0
+ $Y2=0
cc_564 N_A_610_47#_M1031_g N_X_c_1163_n 0.00253248f $X=9.855 $Y=2.465 $X2=0
+ $Y2=0
cc_565 N_A_610_47#_M1038_g N_X_c_1163_n 0.00362883f $X=10.285 $Y=0.655 $X2=0
+ $Y2=0
cc_566 N_A_610_47#_M1036_g N_X_c_1163_n 0.00253248f $X=10.285 $Y=2.465 $X2=0
+ $Y2=0
cc_567 N_A_610_47#_c_582_n N_X_c_1163_n 0.029632f $X=11.36 $Y=1.665 $X2=0 $Y2=0
cc_568 N_A_610_47#_c_587_n N_X_c_1163_n 0.0310539f $X=9.64 $Y=1.48 $X2=0 $Y2=0
cc_569 N_A_610_47#_c_588_n N_X_c_1163_n 0.0310539f $X=10.5 $Y=1.48 $X2=0 $Y2=0
cc_570 N_A_610_47#_c_590_n N_X_c_1163_n 0.0209262f $X=12.005 $Y=1.48 $X2=0 $Y2=0
cc_571 N_A_610_47#_M1043_g N_X_c_1164_n 0.00362883f $X=10.715 $Y=0.655 $X2=0
+ $Y2=0
cc_572 N_A_610_47#_M1037_g N_X_c_1164_n 0.00253248f $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_573 N_A_610_47#_M1044_g N_X_c_1164_n 0.00362883f $X=11.145 $Y=0.655 $X2=0
+ $Y2=0
cc_574 N_A_610_47#_M1045_g N_X_c_1164_n 0.00253248f $X=11.145 $Y=2.465 $X2=0
+ $Y2=0
cc_575 N_A_610_47#_c_582_n N_X_c_1164_n 0.0295864f $X=11.36 $Y=1.665 $X2=0 $Y2=0
cc_576 N_A_610_47#_c_588_n N_X_c_1164_n 0.0310539f $X=10.5 $Y=1.48 $X2=0 $Y2=0
cc_577 N_A_610_47#_c_589_n N_X_c_1164_n 0.0310539f $X=11.36 $Y=1.48 $X2=0 $Y2=0
cc_578 N_A_610_47#_c_590_n N_X_c_1164_n 0.0209262f $X=12.005 $Y=1.48 $X2=0 $Y2=0
cc_579 N_A_610_47#_M1046_g N_X_c_1165_n 0.00362883f $X=11.575 $Y=0.655 $X2=0
+ $Y2=0
cc_580 N_A_610_47#_M1047_g N_X_c_1165_n 0.00270348f $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_581 N_A_610_47#_M1049_g N_X_c_1165_n 0.00673525f $X=12.005 $Y=0.655 $X2=0
+ $Y2=0
cc_582 N_A_610_47#_M1050_g N_X_c_1165_n 0.00589224f $X=12.005 $Y=2.465 $X2=0
+ $Y2=0
cc_583 N_A_610_47#_c_582_n N_X_c_1165_n 0.00698543f $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_584 N_A_610_47#_c_589_n N_X_c_1165_n 0.0303505f $X=11.36 $Y=1.48 $X2=0 $Y2=0
cc_585 N_A_610_47#_c_590_n N_X_c_1165_n 0.0308454f $X=12.005 $Y=1.48 $X2=0 $Y2=0
cc_586 N_A_610_47#_M1000_g N_X_c_1174_n 0.00292296f $X=5.555 $Y=2.465 $X2=0
+ $Y2=0
cc_587 N_A_610_47#_M1004_g N_X_c_1174_n 0.00766908f $X=5.985 $Y=2.465 $X2=0
+ $Y2=0
cc_588 N_A_610_47#_M1005_g N_X_c_1174_n 0.00766908f $X=6.415 $Y=2.465 $X2=0
+ $Y2=0
cc_589 N_A_610_47#_M1007_g N_X_c_1174_n 0.00766908f $X=6.845 $Y=2.465 $X2=0
+ $Y2=0
cc_590 N_A_610_47#_M1010_g N_X_c_1174_n 0.00766908f $X=7.275 $Y=2.465 $X2=0
+ $Y2=0
cc_591 N_A_610_47#_M1015_g N_X_c_1174_n 0.00766908f $X=7.705 $Y=2.465 $X2=0
+ $Y2=0
cc_592 N_A_610_47#_M1017_g N_X_c_1174_n 0.00766908f $X=8.135 $Y=2.465 $X2=0
+ $Y2=0
cc_593 N_A_610_47#_M1020_g N_X_c_1174_n 0.00766908f $X=8.565 $Y=2.465 $X2=0
+ $Y2=0
cc_594 N_A_610_47#_M1021_g N_X_c_1174_n 0.00766908f $X=8.995 $Y=2.465 $X2=0
+ $Y2=0
cc_595 N_A_610_47#_M1026_g N_X_c_1174_n 0.00766908f $X=9.425 $Y=2.465 $X2=0
+ $Y2=0
cc_596 N_A_610_47#_M1031_g N_X_c_1174_n 0.00766908f $X=9.855 $Y=2.465 $X2=0
+ $Y2=0
cc_597 N_A_610_47#_M1036_g N_X_c_1174_n 0.00766908f $X=10.285 $Y=2.465 $X2=0
+ $Y2=0
cc_598 N_A_610_47#_M1037_g N_X_c_1174_n 0.00766908f $X=10.715 $Y=2.465 $X2=0
+ $Y2=0
cc_599 N_A_610_47#_M1045_g N_X_c_1174_n 0.00766908f $X=11.145 $Y=2.465 $X2=0
+ $Y2=0
cc_600 N_A_610_47#_M1047_g N_X_c_1174_n 0.0123908f $X=11.575 $Y=2.465 $X2=0
+ $Y2=0
cc_601 N_A_610_47#_M1050_g N_X_c_1174_n 0.002131f $X=12.005 $Y=2.465 $X2=0 $Y2=0
cc_602 N_A_610_47#_c_715_p N_X_c_1174_n 0.00375391f $X=4.91 $Y=2.045 $X2=0 $Y2=0
cc_603 N_A_610_47#_c_582_n N_X_c_1174_n 0.579595f $X=11.36 $Y=1.665 $X2=0 $Y2=0
cc_604 N_A_610_47#_c_583_n N_X_c_1174_n 8.1932e-19 $X=6.2 $Y=1.48 $X2=0 $Y2=0
cc_605 N_A_610_47#_c_584_n N_X_c_1174_n 8.1932e-19 $X=7.06 $Y=1.48 $X2=0 $Y2=0
cc_606 N_A_610_47#_c_585_n N_X_c_1174_n 8.1932e-19 $X=7.92 $Y=1.48 $X2=0 $Y2=0
cc_607 N_A_610_47#_c_586_n N_X_c_1174_n 8.1932e-19 $X=8.78 $Y=1.48 $X2=0 $Y2=0
cc_608 N_A_610_47#_c_587_n N_X_c_1174_n 8.1932e-19 $X=9.64 $Y=1.48 $X2=0 $Y2=0
cc_609 N_A_610_47#_c_588_n N_X_c_1174_n 8.1932e-19 $X=10.5 $Y=1.48 $X2=0 $Y2=0
cc_610 N_A_610_47#_c_589_n N_X_c_1174_n 8.1932e-19 $X=11.36 $Y=1.48 $X2=0 $Y2=0
cc_611 N_A_610_47#_c_575_n N_VGND_M1011_d 0.00176461f $X=3.92 $Y=1.13 $X2=0
+ $Y2=0
cc_612 N_A_610_47#_c_577_n N_VGND_M1029_d 0.00176461f $X=4.78 $Y=1.13 $X2=0
+ $Y2=0
cc_613 N_A_610_47#_c_578_n N_VGND_M1035_d 0.00180544f $X=5.305 $Y=1.13 $X2=0
+ $Y2=0
cc_614 N_A_610_47#_c_575_n N_VGND_c_1347_n 0.0152916f $X=3.92 $Y=1.13 $X2=0
+ $Y2=0
cc_615 N_A_610_47#_c_577_n N_VGND_c_1348_n 0.0135055f $X=4.78 $Y=1.13 $X2=0
+ $Y2=0
cc_616 N_A_610_47#_M1002_g N_VGND_c_1349_n 0.0016342f $X=5.555 $Y=0.655 $X2=0
+ $Y2=0
cc_617 N_A_610_47#_c_578_n N_VGND_c_1349_n 0.0145078f $X=5.305 $Y=1.13 $X2=0
+ $Y2=0
cc_618 N_A_610_47#_M1006_g N_VGND_c_1350_n 0.00190642f $X=5.985 $Y=0.655 $X2=0
+ $Y2=0
cc_619 N_A_610_47#_M1009_g N_VGND_c_1350_n 0.00190642f $X=6.415 $Y=0.655 $X2=0
+ $Y2=0
cc_620 N_A_610_47#_c_582_n N_VGND_c_1350_n 0.00138201f $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_621 N_A_610_47#_c_583_n N_VGND_c_1350_n 0.0125963f $X=6.2 $Y=1.48 $X2=0 $Y2=0
cc_622 N_A_610_47#_c_590_n N_VGND_c_1350_n 7.58855e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_623 N_A_610_47#_M1009_g N_VGND_c_1351_n 0.00585385f $X=6.415 $Y=0.655 $X2=0
+ $Y2=0
cc_624 N_A_610_47#_M1012_g N_VGND_c_1351_n 0.00585385f $X=6.845 $Y=0.655 $X2=0
+ $Y2=0
cc_625 N_A_610_47#_M1012_g N_VGND_c_1352_n 0.00190642f $X=6.845 $Y=0.655 $X2=0
+ $Y2=0
cc_626 N_A_610_47#_M1013_g N_VGND_c_1352_n 0.00190642f $X=7.275 $Y=0.655 $X2=0
+ $Y2=0
cc_627 N_A_610_47#_c_582_n N_VGND_c_1352_n 0.00138201f $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_628 N_A_610_47#_c_584_n N_VGND_c_1352_n 0.0125963f $X=7.06 $Y=1.48 $X2=0
+ $Y2=0
cc_629 N_A_610_47#_c_590_n N_VGND_c_1352_n 7.58855e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_630 N_A_610_47#_M1014_g N_VGND_c_1353_n 0.00190642f $X=7.705 $Y=0.655 $X2=0
+ $Y2=0
cc_631 N_A_610_47#_M1016_g N_VGND_c_1353_n 0.00190642f $X=8.135 $Y=0.655 $X2=0
+ $Y2=0
cc_632 N_A_610_47#_c_582_n N_VGND_c_1353_n 0.00138201f $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_633 N_A_610_47#_c_585_n N_VGND_c_1353_n 0.0125963f $X=7.92 $Y=1.48 $X2=0
+ $Y2=0
cc_634 N_A_610_47#_c_590_n N_VGND_c_1353_n 7.58855e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_635 N_A_610_47#_M1024_g N_VGND_c_1354_n 0.00190642f $X=8.565 $Y=0.655 $X2=0
+ $Y2=0
cc_636 N_A_610_47#_M1028_g N_VGND_c_1354_n 0.00190642f $X=8.995 $Y=0.655 $X2=0
+ $Y2=0
cc_637 N_A_610_47#_c_582_n N_VGND_c_1354_n 0.00138201f $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_638 N_A_610_47#_c_586_n N_VGND_c_1354_n 0.0125963f $X=8.78 $Y=1.48 $X2=0
+ $Y2=0
cc_639 N_A_610_47#_c_590_n N_VGND_c_1354_n 7.58855e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_640 N_A_610_47#_M1030_g N_VGND_c_1355_n 0.00190642f $X=9.425 $Y=0.655 $X2=0
+ $Y2=0
cc_641 N_A_610_47#_M1034_g N_VGND_c_1355_n 0.00190642f $X=9.855 $Y=0.655 $X2=0
+ $Y2=0
cc_642 N_A_610_47#_c_582_n N_VGND_c_1355_n 0.00138201f $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_643 N_A_610_47#_c_587_n N_VGND_c_1355_n 0.0125963f $X=9.64 $Y=1.48 $X2=0
+ $Y2=0
cc_644 N_A_610_47#_c_590_n N_VGND_c_1355_n 7.58855e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_645 N_A_610_47#_M1038_g N_VGND_c_1356_n 0.00190642f $X=10.285 $Y=0.655 $X2=0
+ $Y2=0
cc_646 N_A_610_47#_M1043_g N_VGND_c_1356_n 0.00190642f $X=10.715 $Y=0.655 $X2=0
+ $Y2=0
cc_647 N_A_610_47#_c_582_n N_VGND_c_1356_n 0.00138201f $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_648 N_A_610_47#_c_588_n N_VGND_c_1356_n 0.0125963f $X=10.5 $Y=1.48 $X2=0
+ $Y2=0
cc_649 N_A_610_47#_c_590_n N_VGND_c_1356_n 7.58855e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_650 N_A_610_47#_M1043_g N_VGND_c_1357_n 0.00585385f $X=10.715 $Y=0.655 $X2=0
+ $Y2=0
cc_651 N_A_610_47#_M1044_g N_VGND_c_1357_n 0.00585385f $X=11.145 $Y=0.655 $X2=0
+ $Y2=0
cc_652 N_A_610_47#_M1044_g N_VGND_c_1358_n 0.00190642f $X=11.145 $Y=0.655 $X2=0
+ $Y2=0
cc_653 N_A_610_47#_M1046_g N_VGND_c_1358_n 0.00190642f $X=11.575 $Y=0.655 $X2=0
+ $Y2=0
cc_654 N_A_610_47#_c_582_n N_VGND_c_1358_n 0.00138201f $X=11.36 $Y=1.665 $X2=0
+ $Y2=0
cc_655 N_A_610_47#_c_589_n N_VGND_c_1358_n 0.0125963f $X=11.36 $Y=1.48 $X2=0
+ $Y2=0
cc_656 N_A_610_47#_c_590_n N_VGND_c_1358_n 7.58855e-19 $X=12.005 $Y=1.48 $X2=0
+ $Y2=0
cc_657 N_A_610_47#_M1049_g N_VGND_c_1360_n 0.00462267f $X=12.005 $Y=0.655 $X2=0
+ $Y2=0
cc_658 N_A_610_47#_c_888_p N_VGND_c_1361_n 0.0149362f $X=4.05 $Y=0.45 $X2=0
+ $Y2=0
cc_659 N_A_610_47#_c_889_p N_VGND_c_1363_n 0.0149362f $X=4.91 $Y=0.45 $X2=0
+ $Y2=0
cc_660 N_A_610_47#_M1002_g N_VGND_c_1365_n 0.00585385f $X=5.555 $Y=0.655 $X2=0
+ $Y2=0
cc_661 N_A_610_47#_M1006_g N_VGND_c_1365_n 0.00585385f $X=5.985 $Y=0.655 $X2=0
+ $Y2=0
cc_662 N_A_610_47#_M1016_g N_VGND_c_1367_n 0.00585385f $X=8.135 $Y=0.655 $X2=0
+ $Y2=0
cc_663 N_A_610_47#_M1024_g N_VGND_c_1367_n 0.00585385f $X=8.565 $Y=0.655 $X2=0
+ $Y2=0
cc_664 N_A_610_47#_M1028_g N_VGND_c_1369_n 0.00585385f $X=8.995 $Y=0.655 $X2=0
+ $Y2=0
cc_665 N_A_610_47#_M1030_g N_VGND_c_1369_n 0.00585385f $X=9.425 $Y=0.655 $X2=0
+ $Y2=0
cc_666 N_A_610_47#_M1034_g N_VGND_c_1371_n 0.00585385f $X=9.855 $Y=0.655 $X2=0
+ $Y2=0
cc_667 N_A_610_47#_M1038_g N_VGND_c_1371_n 0.00585385f $X=10.285 $Y=0.655 $X2=0
+ $Y2=0
cc_668 N_A_610_47#_c_898_p N_VGND_c_1375_n 0.0138717f $X=3.19 $Y=0.45 $X2=0
+ $Y2=0
cc_669 N_A_610_47#_M1013_g N_VGND_c_1376_n 0.00585385f $X=7.275 $Y=0.655 $X2=0
+ $Y2=0
cc_670 N_A_610_47#_M1014_g N_VGND_c_1376_n 0.00585385f $X=7.705 $Y=0.655 $X2=0
+ $Y2=0
cc_671 N_A_610_47#_M1046_g N_VGND_c_1377_n 0.00585385f $X=11.575 $Y=0.655 $X2=0
+ $Y2=0
cc_672 N_A_610_47#_M1049_g N_VGND_c_1377_n 0.00585385f $X=12.005 $Y=0.655 $X2=0
+ $Y2=0
cc_673 N_A_610_47#_M1008_s N_VGND_c_1385_n 0.00406062f $X=3.05 $Y=0.235 $X2=0
+ $Y2=0
cc_674 N_A_610_47#_M1023_s N_VGND_c_1385_n 0.003017f $X=3.91 $Y=0.235 $X2=0
+ $Y2=0
cc_675 N_A_610_47#_M1033_s N_VGND_c_1385_n 0.003017f $X=4.77 $Y=0.235 $X2=0
+ $Y2=0
cc_676 N_A_610_47#_M1002_g N_VGND_c_1385_n 0.0106555f $X=5.555 $Y=0.655 $X2=0
+ $Y2=0
cc_677 N_A_610_47#_M1006_g N_VGND_c_1385_n 0.0107375f $X=5.985 $Y=0.655 $X2=0
+ $Y2=0
cc_678 N_A_610_47#_M1009_g N_VGND_c_1385_n 0.0107375f $X=6.415 $Y=0.655 $X2=0
+ $Y2=0
cc_679 N_A_610_47#_M1012_g N_VGND_c_1385_n 0.0107375f $X=6.845 $Y=0.655 $X2=0
+ $Y2=0
cc_680 N_A_610_47#_M1013_g N_VGND_c_1385_n 0.0107375f $X=7.275 $Y=0.655 $X2=0
+ $Y2=0
cc_681 N_A_610_47#_M1014_g N_VGND_c_1385_n 0.0107375f $X=7.705 $Y=0.655 $X2=0
+ $Y2=0
cc_682 N_A_610_47#_M1016_g N_VGND_c_1385_n 0.0107375f $X=8.135 $Y=0.655 $X2=0
+ $Y2=0
cc_683 N_A_610_47#_M1024_g N_VGND_c_1385_n 0.0107375f $X=8.565 $Y=0.655 $X2=0
+ $Y2=0
cc_684 N_A_610_47#_M1028_g N_VGND_c_1385_n 0.0107375f $X=8.995 $Y=0.655 $X2=0
+ $Y2=0
cc_685 N_A_610_47#_M1030_g N_VGND_c_1385_n 0.0107375f $X=9.425 $Y=0.655 $X2=0
+ $Y2=0
cc_686 N_A_610_47#_M1034_g N_VGND_c_1385_n 0.0107375f $X=9.855 $Y=0.655 $X2=0
+ $Y2=0
cc_687 N_A_610_47#_M1038_g N_VGND_c_1385_n 0.0107375f $X=10.285 $Y=0.655 $X2=0
+ $Y2=0
cc_688 N_A_610_47#_M1043_g N_VGND_c_1385_n 0.0107375f $X=10.715 $Y=0.655 $X2=0
+ $Y2=0
cc_689 N_A_610_47#_M1044_g N_VGND_c_1385_n 0.0107375f $X=11.145 $Y=0.655 $X2=0
+ $Y2=0
cc_690 N_A_610_47#_M1046_g N_VGND_c_1385_n 0.0107375f $X=11.575 $Y=0.655 $X2=0
+ $Y2=0
cc_691 N_A_610_47#_M1049_g N_VGND_c_1385_n 0.0117419f $X=12.005 $Y=0.655 $X2=0
+ $Y2=0
cc_692 N_A_610_47#_c_898_p N_VGND_c_1385_n 0.00886411f $X=3.19 $Y=0.45 $X2=0
+ $Y2=0
cc_693 N_A_610_47#_c_888_p N_VGND_c_1385_n 0.0100304f $X=4.05 $Y=0.45 $X2=0
+ $Y2=0
cc_694 N_A_610_47#_c_889_p N_VGND_c_1385_n 0.0100304f $X=4.91 $Y=0.45 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_925_n N_X_M1000_d 0.00388669f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_696 N_VPWR_c_925_n N_X_M1005_d 0.003017f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_697 N_VPWR_c_925_n N_X_M1010_d 0.003017f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_698 N_VPWR_c_925_n N_X_M1017_d 0.003017f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_699 N_VPWR_c_925_n N_X_M1021_d 0.003017f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_700 N_VPWR_c_925_n N_X_M1031_d 0.003017f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_701 N_VPWR_c_925_n N_X_M1037_d 0.003017f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_702 N_VPWR_c_925_n N_X_M1047_d 0.003017f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_703 N_VPWR_c_933_n N_X_c_1158_n 0.0080303f $X=6.2 $Y=2.09 $X2=0 $Y2=0
cc_704 N_VPWR_c_948_n N_X_c_1158_n 0.0140491f $X=6.07 $Y=3.33 $X2=0 $Y2=0
cc_705 N_VPWR_c_925_n N_X_c_1158_n 0.0090585f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_706 N_VPWR_c_933_n N_X_c_1159_n 0.00804307f $X=6.2 $Y=2.09 $X2=0 $Y2=0
cc_707 N_VPWR_c_934_n N_X_c_1159_n 0.0149362f $X=6.93 $Y=3.33 $X2=0 $Y2=0
cc_708 N_VPWR_c_935_n N_X_c_1159_n 0.00804307f $X=7.06 $Y=2.09 $X2=0 $Y2=0
cc_709 N_VPWR_c_925_n N_X_c_1159_n 0.0100304f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_710 N_VPWR_c_935_n N_X_c_1160_n 0.00804307f $X=7.06 $Y=2.09 $X2=0 $Y2=0
cc_711 N_VPWR_c_936_n N_X_c_1160_n 0.00804307f $X=7.92 $Y=2.09 $X2=0 $Y2=0
cc_712 N_VPWR_c_959_n N_X_c_1160_n 0.0149362f $X=7.79 $Y=3.33 $X2=0 $Y2=0
cc_713 N_VPWR_c_925_n N_X_c_1160_n 0.0100304f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_714 N_VPWR_c_936_n N_X_c_1161_n 0.00804307f $X=7.92 $Y=2.09 $X2=0 $Y2=0
cc_715 N_VPWR_c_937_n N_X_c_1161_n 0.00804307f $X=8.78 $Y=2.09 $X2=0 $Y2=0
cc_716 N_VPWR_c_950_n N_X_c_1161_n 0.0149362f $X=8.65 $Y=3.33 $X2=0 $Y2=0
cc_717 N_VPWR_c_925_n N_X_c_1161_n 0.0100304f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_718 N_VPWR_c_937_n N_X_c_1162_n 0.00804307f $X=8.78 $Y=2.09 $X2=0 $Y2=0
cc_719 N_VPWR_c_938_n N_X_c_1162_n 0.00804307f $X=9.64 $Y=2.09 $X2=0 $Y2=0
cc_720 N_VPWR_c_952_n N_X_c_1162_n 0.0149362f $X=9.51 $Y=3.33 $X2=0 $Y2=0
cc_721 N_VPWR_c_925_n N_X_c_1162_n 0.0100304f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_722 N_VPWR_c_938_n N_X_c_1163_n 0.00804307f $X=9.64 $Y=2.09 $X2=0 $Y2=0
cc_723 N_VPWR_c_939_n N_X_c_1163_n 0.00804307f $X=10.5 $Y=2.09 $X2=0 $Y2=0
cc_724 N_VPWR_c_954_n N_X_c_1163_n 0.0149362f $X=10.37 $Y=3.33 $X2=0 $Y2=0
cc_725 N_VPWR_c_925_n N_X_c_1163_n 0.0100304f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_726 N_VPWR_c_939_n N_X_c_1164_n 0.00804307f $X=10.5 $Y=2.09 $X2=0 $Y2=0
cc_727 N_VPWR_c_940_n N_X_c_1164_n 0.0149362f $X=11.23 $Y=3.33 $X2=0 $Y2=0
cc_728 N_VPWR_c_941_n N_X_c_1164_n 0.00804307f $X=11.36 $Y=2.09 $X2=0 $Y2=0
cc_729 N_VPWR_c_925_n N_X_c_1164_n 0.0100304f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_730 N_VPWR_c_941_n N_X_c_1165_n 0.00804307f $X=11.36 $Y=2.09 $X2=0 $Y2=0
cc_731 N_VPWR_c_960_n N_X_c_1165_n 0.0149362f $X=12.09 $Y=3.33 $X2=0 $Y2=0
cc_732 N_VPWR_c_925_n N_X_c_1165_n 0.0100304f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_733 N_VPWR_M1004_s N_X_c_1174_n 0.00192363f $X=6.06 $Y=1.835 $X2=0 $Y2=0
cc_734 N_VPWR_M1007_s N_X_c_1174_n 0.00192363f $X=6.92 $Y=1.835 $X2=0 $Y2=0
cc_735 N_VPWR_M1015_s N_X_c_1174_n 0.00192363f $X=7.78 $Y=1.835 $X2=0 $Y2=0
cc_736 N_VPWR_M1020_s N_X_c_1174_n 0.00192363f $X=8.64 $Y=1.835 $X2=0 $Y2=0
cc_737 N_VPWR_M1026_s N_X_c_1174_n 0.00192363f $X=9.5 $Y=1.835 $X2=0 $Y2=0
cc_738 N_VPWR_M1036_s N_X_c_1174_n 0.00192363f $X=10.36 $Y=1.835 $X2=0 $Y2=0
cc_739 N_VPWR_M1045_s N_X_c_1174_n 0.00192363f $X=11.22 $Y=1.835 $X2=0 $Y2=0
cc_740 N_VPWR_c_932_n N_X_c_1174_n 0.00167362f $X=5.34 $Y=2.26 $X2=0 $Y2=0
cc_741 N_VPWR_c_933_n N_X_c_1174_n 0.0257374f $X=6.2 $Y=2.09 $X2=0 $Y2=0
cc_742 N_VPWR_c_935_n N_X_c_1174_n 0.0257374f $X=7.06 $Y=2.09 $X2=0 $Y2=0
cc_743 N_VPWR_c_936_n N_X_c_1174_n 0.0257374f $X=7.92 $Y=2.09 $X2=0 $Y2=0
cc_744 N_VPWR_c_937_n N_X_c_1174_n 0.0257374f $X=8.78 $Y=2.09 $X2=0 $Y2=0
cc_745 N_VPWR_c_938_n N_X_c_1174_n 0.0257374f $X=9.64 $Y=2.09 $X2=0 $Y2=0
cc_746 N_VPWR_c_939_n N_X_c_1174_n 0.0257374f $X=10.5 $Y=2.09 $X2=0 $Y2=0
cc_747 N_VPWR_c_941_n N_X_c_1174_n 0.0257374f $X=11.36 $Y=2.09 $X2=0 $Y2=0
cc_748 N_VPWR_c_943_n N_X_c_1174_n 0.00676623f $X=12.22 $Y=2.09 $X2=0 $Y2=0
cc_749 N_X_c_1159_n N_VGND_c_1351_n 0.0149362f $X=6.63 $Y=0.45 $X2=0 $Y2=0
cc_750 N_X_c_1164_n N_VGND_c_1357_n 0.0149362f $X=10.93 $Y=0.45 $X2=0 $Y2=0
cc_751 N_X_c_1158_n N_VGND_c_1365_n 0.0140491f $X=5.77 $Y=0.45 $X2=0 $Y2=0
cc_752 N_X_c_1161_n N_VGND_c_1367_n 0.0149362f $X=8.35 $Y=0.45 $X2=0 $Y2=0
cc_753 N_X_c_1162_n N_VGND_c_1369_n 0.0149362f $X=9.21 $Y=0.45 $X2=0 $Y2=0
cc_754 N_X_c_1163_n N_VGND_c_1371_n 0.0149362f $X=10.07 $Y=0.45 $X2=0 $Y2=0
cc_755 N_X_c_1160_n N_VGND_c_1376_n 0.0149362f $X=7.49 $Y=0.45 $X2=0 $Y2=0
cc_756 N_X_c_1165_n N_VGND_c_1377_n 0.0149362f $X=11.79 $Y=0.45 $X2=0 $Y2=0
cc_757 N_X_M1002_d N_VGND_c_1385_n 0.00388669f $X=5.63 $Y=0.235 $X2=0 $Y2=0
cc_758 N_X_M1009_d N_VGND_c_1385_n 0.003017f $X=6.49 $Y=0.235 $X2=0 $Y2=0
cc_759 N_X_M1013_d N_VGND_c_1385_n 0.003017f $X=7.35 $Y=0.235 $X2=0 $Y2=0
cc_760 N_X_M1016_d N_VGND_c_1385_n 0.003017f $X=8.21 $Y=0.235 $X2=0 $Y2=0
cc_761 N_X_M1028_d N_VGND_c_1385_n 0.003017f $X=9.07 $Y=0.235 $X2=0 $Y2=0
cc_762 N_X_M1034_d N_VGND_c_1385_n 0.003017f $X=9.93 $Y=0.235 $X2=0 $Y2=0
cc_763 N_X_M1043_d N_VGND_c_1385_n 0.003017f $X=10.79 $Y=0.235 $X2=0 $Y2=0
cc_764 N_X_M1046_d N_VGND_c_1385_n 0.003017f $X=11.65 $Y=0.235 $X2=0 $Y2=0
cc_765 N_X_c_1158_n N_VGND_c_1385_n 0.0090585f $X=5.77 $Y=0.45 $X2=0 $Y2=0
cc_766 N_X_c_1159_n N_VGND_c_1385_n 0.0100304f $X=6.63 $Y=0.45 $X2=0 $Y2=0
cc_767 N_X_c_1160_n N_VGND_c_1385_n 0.0100304f $X=7.49 $Y=0.45 $X2=0 $Y2=0
cc_768 N_X_c_1161_n N_VGND_c_1385_n 0.0100304f $X=8.35 $Y=0.45 $X2=0 $Y2=0
cc_769 N_X_c_1162_n N_VGND_c_1385_n 0.0100304f $X=9.21 $Y=0.45 $X2=0 $Y2=0
cc_770 N_X_c_1163_n N_VGND_c_1385_n 0.0100304f $X=10.07 $Y=0.45 $X2=0 $Y2=0
cc_771 N_X_c_1164_n N_VGND_c_1385_n 0.0100304f $X=10.93 $Y=0.45 $X2=0 $Y2=0
cc_772 N_X_c_1165_n N_VGND_c_1385_n 0.0100304f $X=11.79 $Y=0.45 $X2=0 $Y2=0
