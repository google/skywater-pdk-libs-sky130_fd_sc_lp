* File: sky130_fd_sc_lp__a41oi_m.pxi.spice
* Created: Wed Sep  2 09:30:01 2020
* 
x_PM_SKY130_FD_SC_LP__A41OI_M%B1 N_B1_c_80_n N_B1_c_81_n N_B1_M1007_g
+ N_B1_M1008_g N_B1_c_83_n N_B1_c_84_n N_B1_c_89_n N_B1_c_90_n N_B1_c_91_n B1 B1
+ B1 B1 B1 N_B1_c_86_n PM_SKY130_FD_SC_LP__A41OI_M%B1
x_PM_SKY130_FD_SC_LP__A41OI_M%A1 N_A1_c_131_n N_A1_M1005_g N_A1_M1001_g
+ N_A1_c_139_n N_A1_c_132_n N_A1_c_133_n A1 A1 A1 N_A1_c_135_n N_A1_c_136_n
+ PM_SKY130_FD_SC_LP__A41OI_M%A1
x_PM_SKY130_FD_SC_LP__A41OI_M%A2 N_A2_M1009_g N_A2_M1003_g N_A2_c_187_n
+ N_A2_c_188_n A2 A2 A2 A2 A2 N_A2_c_190_n PM_SKY130_FD_SC_LP__A41OI_M%A2
x_PM_SKY130_FD_SC_LP__A41OI_M%A3 N_A3_M1006_g N_A3_M1002_g N_A3_c_237_n
+ N_A3_c_238_n A3 A3 A3 A3 N_A3_c_235_n PM_SKY130_FD_SC_LP__A41OI_M%A3
x_PM_SKY130_FD_SC_LP__A41OI_M%A4 N_A4_c_288_n N_A4_M1000_g N_A4_M1004_g
+ N_A4_c_289_n N_A4_c_290_n N_A4_c_282_n N_A4_c_283_n N_A4_c_284_n N_A4_c_285_n
+ A4 A4 A4 A4 A4 N_A4_c_287_n PM_SKY130_FD_SC_LP__A41OI_M%A4
x_PM_SKY130_FD_SC_LP__A41OI_M%Y N_Y_M1008_d N_Y_M1007_s N_Y_c_324_n N_Y_c_325_n
+ Y Y Y Y Y Y PM_SKY130_FD_SC_LP__A41OI_M%Y
x_PM_SKY130_FD_SC_LP__A41OI_M%A_186_531# N_A_186_531#_M1007_d
+ N_A_186_531#_M1009_d N_A_186_531#_M1000_d N_A_186_531#_c_356_n
+ N_A_186_531#_c_357_n N_A_186_531#_c_358_n N_A_186_531#_c_359_n
+ N_A_186_531#_c_360_n N_A_186_531#_c_361_n N_A_186_531#_c_362_n
+ PM_SKY130_FD_SC_LP__A41OI_M%A_186_531#
x_PM_SKY130_FD_SC_LP__A41OI_M%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_c_405_n
+ N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n
+ VPWR N_VPWR_c_411_n N_VPWR_c_404_n PM_SKY130_FD_SC_LP__A41OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A41OI_M%VGND N_VGND_M1008_s N_VGND_M1004_d N_VGND_c_447_n
+ N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n VGND N_VGND_c_451_n
+ N_VGND_c_452_n N_VGND_c_453_n PM_SKY130_FD_SC_LP__A41OI_M%VGND
cc_1 VNB N_B1_c_80_n 0.0216197f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.895
cc_2 VNB N_B1_c_81_n 0.0134079f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.895
cc_3 VNB N_B1_M1008_g 0.0266378f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.445
cc_4 VNB N_B1_c_83_n 0.0158199f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.21
cc_5 VNB N_B1_c_84_n 0.0209297f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.715
cc_6 VNB B1 7.95909e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_B1_c_86_n 0.0147005f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.375
cc_8 VNB N_A1_c_131_n 0.0189444f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.21
cc_9 VNB N_A1_c_132_n 0.0159281f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.445
cc_10 VNB N_A1_c_133_n 0.0136504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A1 0.00162753f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.375
cc_12 VNB N_A1_c_135_n 0.0183239f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_13 VNB N_A1_c_136_n 0.0171941f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_14 VNB N_A2_M1003_g 0.0304458f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.27
cc_15 VNB N_A2_c_187_n 0.0209231f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.82
cc_16 VNB N_A2_c_188_n 0.00154757f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.445
cc_17 VNB A2 0.0125656f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.445
cc_18 VNB N_A2_c_190_n 0.0174836f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_19 VNB N_A3_M1002_g 0.0595584f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.27
cc_20 VNB A3 0.0155328f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.445
cc_21 VNB N_A3_c_235_n 0.0232714f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_22 VNB N_A4_M1004_g 0.0267104f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=2.12
cc_23 VNB N_A4_c_282_n 0.0439887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A4_c_283_n 0.00705639f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.82
cc_25 VNB N_A4_c_284_n 0.00885579f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.445
cc_26 VNB N_A4_c_285_n 0.0253898f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.21
cc_27 VNB A4 0.00912409f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.715
cc_28 VNB N_A4_c_287_n 0.0382913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_324_n 0.0157392f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.27
cc_30 VNB N_Y_c_325_n 0.00244252f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.82
cc_31 VNB Y 0.0138974f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.445
cc_32 VNB Y 0.0342477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_404_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_447_n 0.00495479f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.82
cc_35 VNB N_VGND_c_448_n 0.0127868f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.375
cc_36 VNB N_VGND_c_449_n 0.0520838f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.88
cc_37 VNB N_VGND_c_450_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0.822 $Y2=2.12
cc_38 VNB N_VGND_c_451_n 0.0137583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_452_n 0.201407f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.375
cc_40 VNB N_VGND_c_453_n 0.0276349f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.295
cc_41 VPB N_B1_M1007_g 0.0379122f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.865
cc_42 VPB N_B1_c_84_n 0.004426f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.715
cc_43 VPB N_B1_c_89_n 0.0196803f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.88
cc_44 VPB N_B1_c_90_n 0.0156631f $X=-0.19 $Y=1.655 $X2=0.822 $Y2=2.12
cc_45 VPB N_B1_c_91_n 0.016068f $X=-0.19 $Y=1.655 $X2=0.822 $Y2=2.27
cc_46 VPB B1 0.00727229f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_47 VPB N_A1_c_131_n 0.00333478f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.21
cc_48 VPB N_A1_M1005_g 0.0499803f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=1.88
cc_49 VPB N_A1_c_139_n 0.0190504f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.445
cc_50 VPB A1 0.00297037f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.375
cc_51 VPB N_A2_M1009_g 0.0523751f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.895
cc_52 VPB N_A2_c_188_n 0.0144102f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.445
cc_53 VPB A2 0.00821575f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.445
cc_54 VPB N_A3_M1006_g 0.038303f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.895
cc_55 VPB N_A3_c_237_n 0.0234306f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.82
cc_56 VPB N_A3_c_238_n 0.0302145f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.445
cc_57 VPB A3 0.00613112f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.445
cc_58 VPB N_A3_c_235_n 0.00918679f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_59 VPB N_A4_c_288_n 0.0201018f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.97
cc_60 VPB N_A4_c_289_n 0.0360499f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.865
cc_61 VPB N_A4_c_290_n 0.00720082f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.865
cc_62 VPB N_A4_c_284_n 0.0459522f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.445
cc_63 VPB A4 0.0318983f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.715
cc_64 VPB Y 0.0660314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_186_531#_c_356_n 7.6827e-19 $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.445
cc_66 VPB N_A_186_531#_c_357_n 0.0115551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_186_531#_c_358_n 0.00597734f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.375
cc_68 VPB N_A_186_531#_c_359_n 7.90901e-19 $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.88
cc_69 VPB N_A_186_531#_c_360_n 0.00721802f $X=-0.19 $Y=1.655 $X2=0.822 $Y2=2.27
cc_70 VPB N_A_186_531#_c_361_n 0.00448409f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_71 VPB N_A_186_531#_c_362_n 0.0130318f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_72 VPB N_VPWR_c_405_n 0.00495206f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.865
cc_73 VPB N_VPWR_c_406_n 0.00482547f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.445
cc_74 VPB N_VPWR_c_407_n 0.0410689f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.21
cc_75 VPB N_VPWR_c_408_n 0.00401177f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.715
cc_76 VPB N_VPWR_c_409_n 0.0173909f $X=-0.19 $Y=1.655 $X2=0.822 $Y2=2.12
cc_77 VPB N_VPWR_c_410_n 0.00362723f $X=-0.19 $Y=1.655 $X2=0.822 $Y2=2.27
cc_78 VPB N_VPWR_c_411_n 0.0283708f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.295
cc_79 VPB N_VPWR_c_404_n 0.0748153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 N_B1_c_84_n N_A1_c_131_n 0.0138922f $X=0.7 $Y=1.715 $X2=0 $Y2=0
cc_81 N_B1_c_90_n N_A1_M1005_g 0.00740356f $X=0.822 $Y=2.12 $X2=0 $Y2=0
cc_82 N_B1_c_91_n N_A1_M1005_g 0.0342125f $X=0.822 $Y=2.27 $X2=0 $Y2=0
cc_83 B1 N_A1_M1005_g 0.00200385f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_84 N_B1_c_89_n N_A1_c_139_n 0.0138922f $X=0.7 $Y=1.88 $X2=0 $Y2=0
cc_85 N_B1_M1008_g N_A1_c_132_n 0.0140947f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_86 N_B1_M1008_g N_A1_c_133_n 0.00642957f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_87 N_B1_c_90_n A1 0.00163733f $X=0.822 $Y=2.12 $X2=0 $Y2=0
cc_88 B1 A1 0.0399209f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_89 N_B1_c_86_n A1 0.00228901f $X=0.7 $Y=1.375 $X2=0 $Y2=0
cc_90 B1 N_A1_c_135_n 0.002219f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B1_c_86_n N_A1_c_135_n 0.0138922f $X=0.7 $Y=1.375 $X2=0 $Y2=0
cc_92 N_B1_c_80_n N_A1_c_136_n 0.00642957f $X=0.92 $Y=0.895 $X2=0 $Y2=0
cc_93 N_B1_c_83_n N_A1_c_136_n 0.00560802f $X=0.7 $Y=1.21 $X2=0 $Y2=0
cc_94 B1 N_Y_M1007_s 0.00380424f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_95 N_B1_c_80_n N_Y_c_324_n 0.0154372f $X=0.92 $Y=0.895 $X2=0 $Y2=0
cc_96 N_B1_c_81_n N_Y_c_324_n 0.00745684f $X=0.685 $Y=0.895 $X2=0 $Y2=0
cc_97 N_B1_c_83_n N_Y_c_324_n 0.00668311f $X=0.7 $Y=1.21 $X2=0 $Y2=0
cc_98 B1 N_Y_c_324_n 0.0130189f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_99 N_B1_c_86_n N_Y_c_324_n 0.00163404f $X=0.7 $Y=1.375 $X2=0 $Y2=0
cc_100 N_B1_M1008_g N_Y_c_325_n 0.00461748f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_101 N_B1_M1007_g Y 0.0051606f $X=0.855 $Y=2.865 $X2=0 $Y2=0
cc_102 N_B1_c_83_n Y 0.0243871f $X=0.7 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B1_c_90_n Y 0.0022208f $X=0.822 $Y=2.12 $X2=0 $Y2=0
cc_104 B1 Y 0.121791f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B1_M1007_g N_A_186_531#_c_356_n 3.54603e-19 $X=0.855 $Y=2.865 $X2=0
+ $Y2=0
cc_106 B1 N_A_186_531#_c_356_n 0.0101614f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_107 N_B1_M1007_g N_A_186_531#_c_358_n 0.00140852f $X=0.855 $Y=2.865 $X2=0
+ $Y2=0
cc_108 B1 N_A_186_531#_c_358_n 0.0132332f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B1_M1007_g N_VPWR_c_407_n 0.00536034f $X=0.855 $Y=2.865 $X2=0 $Y2=0
cc_110 B1 N_VPWR_c_407_n 0.0046355f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B1_M1007_g N_VPWR_c_404_n 0.0111323f $X=0.855 $Y=2.865 $X2=0 $Y2=0
cc_112 B1 N_VPWR_c_404_n 0.00630181f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B1_c_81_n N_VGND_c_447_n 0.00393459f $X=0.685 $Y=0.895 $X2=0 $Y2=0
cc_114 N_B1_M1008_g N_VGND_c_447_n 0.00460896f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_115 N_B1_M1008_g N_VGND_c_449_n 0.00585385f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_116 N_B1_c_81_n N_VGND_c_452_n 0.00434699f $X=0.685 $Y=0.895 $X2=0 $Y2=0
cc_117 N_B1_M1008_g N_VGND_c_452_n 0.00760785f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_118 N_A1_M1005_g N_A2_M1009_g 0.0461349f $X=1.285 $Y=2.865 $X2=0 $Y2=0
cc_119 N_A1_c_139_n N_A2_M1009_g 0.0117231f $X=1.252 $Y=1.88 $X2=0 $Y2=0
cc_120 N_A1_c_132_n N_A2_M1003_g 0.050197f $X=1.39 $Y=0.765 $X2=0 $Y2=0
cc_121 N_A1_c_136_n N_A2_M1003_g 0.00847404f $X=1.252 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A1_c_135_n N_A2_c_187_n 0.0117231f $X=1.24 $Y=1.375 $X2=0 $Y2=0
cc_123 N_A1_c_131_n N_A2_c_188_n 0.0117231f $X=1.252 $Y=1.703 $X2=0 $Y2=0
cc_124 N_A1_M1005_g A2 0.00150711f $X=1.285 $Y=2.865 $X2=0 $Y2=0
cc_125 N_A1_c_132_n A2 0.00339156f $X=1.39 $Y=0.765 $X2=0 $Y2=0
cc_126 A1 A2 0.0489131f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A1_c_136_n A2 0.00993345f $X=1.252 $Y=1.21 $X2=0 $Y2=0
cc_128 A1 N_A2_c_190_n 9.49951e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_129 N_A1_c_136_n N_A2_c_190_n 0.0117231f $X=1.252 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A1_c_133_n N_Y_c_324_n 0.00179843f $X=1.39 $Y=0.915 $X2=0 $Y2=0
cc_131 A1 N_Y_c_324_n 0.0154981f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A1_c_135_n N_Y_c_324_n 0.00293277f $X=1.24 $Y=1.375 $X2=0 $Y2=0
cc_133 N_A1_c_136_n N_Y_c_324_n 0.00305007f $X=1.252 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A1_c_132_n N_Y_c_325_n 9.96744e-19 $X=1.39 $Y=0.765 $X2=0 $Y2=0
cc_135 N_A1_c_133_n N_Y_c_325_n 0.00230285f $X=1.39 $Y=0.915 $X2=0 $Y2=0
cc_136 N_A1_M1005_g N_A_186_531#_c_356_n 6.60816e-19 $X=1.285 $Y=2.865 $X2=0
+ $Y2=0
cc_137 N_A1_M1005_g N_A_186_531#_c_357_n 0.0134072f $X=1.285 $Y=2.865 $X2=0
+ $Y2=0
cc_138 N_A1_c_139_n N_A_186_531#_c_357_n 0.00208123f $X=1.252 $Y=1.88 $X2=0
+ $Y2=0
cc_139 A1 N_A_186_531#_c_357_n 0.00718942f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A1_c_139_n N_A_186_531#_c_358_n 0.00153292f $X=1.252 $Y=1.88 $X2=0
+ $Y2=0
cc_141 A1 N_A_186_531#_c_358_n 0.00351692f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_142 N_A1_M1005_g N_VPWR_c_405_n 0.002825f $X=1.285 $Y=2.865 $X2=0 $Y2=0
cc_143 N_A1_M1005_g N_VPWR_c_407_n 0.00420792f $X=1.285 $Y=2.865 $X2=0 $Y2=0
cc_144 N_A1_M1005_g N_VPWR_c_404_n 0.0058978f $X=1.285 $Y=2.865 $X2=0 $Y2=0
cc_145 N_A1_c_132_n N_VGND_c_449_n 0.00585385f $X=1.39 $Y=0.765 $X2=0 $Y2=0
cc_146 N_A1_c_133_n N_VGND_c_449_n 7.95576e-19 $X=1.39 $Y=0.915 $X2=0 $Y2=0
cc_147 N_A1_c_132_n N_VGND_c_452_n 0.0108402f $X=1.39 $Y=0.765 $X2=0 $Y2=0
cc_148 N_A1_c_133_n N_VGND_c_452_n 9.62037e-19 $X=1.39 $Y=0.915 $X2=0 $Y2=0
cc_149 N_A2_M1003_g N_A3_M1002_g 0.0389855f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_150 A2 N_A3_M1002_g 0.00901616f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_151 N_A2_c_190_n N_A3_M1002_g 0.0141403f $X=1.805 $Y=1.29 $X2=0 $Y2=0
cc_152 N_A2_M1009_g N_A3_c_237_n 0.00685108f $X=1.715 $Y=2.865 $X2=0 $Y2=0
cc_153 N_A2_c_188_n N_A3_c_237_n 0.0141403f $X=1.805 $Y=1.795 $X2=0 $Y2=0
cc_154 A2 N_A3_c_237_n 0.00245285f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_155 N_A2_M1009_g N_A3_c_238_n 0.0391733f $X=1.715 $Y=2.865 $X2=0 $Y2=0
cc_156 A2 N_A3_c_238_n 9.58344e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A2_M1009_g A3 4.64094e-19 $X=1.715 $Y=2.865 $X2=0 $Y2=0
cc_158 N_A2_c_187_n A3 6.90611e-19 $X=1.805 $Y=1.63 $X2=0 $Y2=0
cc_159 A2 A3 0.0412059f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_160 N_A2_c_187_n N_A3_c_235_n 0.0141403f $X=1.805 $Y=1.63 $X2=0 $Y2=0
cc_161 A2 N_Y_c_324_n 0.00969313f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_162 A2 N_Y_c_325_n 0.0151242f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_163 N_A2_M1009_g N_A_186_531#_c_357_n 0.0129381f $X=1.715 $Y=2.865 $X2=0
+ $Y2=0
cc_164 A2 N_A_186_531#_c_357_n 0.0112793f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_165 N_A2_M1009_g N_A_186_531#_c_359_n 6.71115e-19 $X=1.715 $Y=2.865 $X2=0
+ $Y2=0
cc_166 N_A2_c_188_n N_A_186_531#_c_361_n 0.00256253f $X=1.805 $Y=1.795 $X2=0
+ $Y2=0
cc_167 A2 N_A_186_531#_c_361_n 0.0038256f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_168 N_A2_M1009_g N_VPWR_c_405_n 0.00153867f $X=1.715 $Y=2.865 $X2=0 $Y2=0
cc_169 N_A2_M1009_g N_VPWR_c_409_n 0.00420792f $X=1.715 $Y=2.865 $X2=0 $Y2=0
cc_170 N_A2_M1009_g N_VPWR_c_404_n 0.0058978f $X=1.715 $Y=2.865 $X2=0 $Y2=0
cc_171 N_A2_M1003_g N_VGND_c_449_n 0.00398598f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_172 A2 N_VGND_c_449_n 0.00709152f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_173 N_A2_M1003_g N_VGND_c_452_n 0.00561906f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_174 A2 N_VGND_c_452_n 0.00925592f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_175 A2 A_300_47# 0.00271508f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_176 N_A3_M1002_g N_A4_M1004_g 0.0558751f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_177 A3 N_A4_c_289_n 7.87816e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_178 N_A3_M1006_g N_A4_c_290_n 0.0224778f $X=2.145 $Y=2.865 $X2=0 $Y2=0
cc_179 N_A3_c_238_n N_A4_c_290_n 0.0121061f $X=2.377 $Y=2.185 $X2=0 $Y2=0
cc_180 A3 N_A4_c_290_n 7.27227e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_181 A3 N_A4_c_282_n 0.00413797f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_182 A3 N_A4_c_283_n 0.00967042f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_183 N_A3_c_235_n N_A4_c_283_n 0.00259152f $X=2.52 $Y=1.68 $X2=0 $Y2=0
cc_184 N_A3_M1006_g N_A4_c_284_n 0.0025741f $X=2.145 $Y=2.865 $X2=0 $Y2=0
cc_185 N_A3_c_235_n N_A4_c_284_n 0.0336069f $X=2.52 $Y=1.68 $X2=0 $Y2=0
cc_186 A3 A4 0.0694605f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_187 N_A3_c_235_n A4 7.11724e-19 $X=2.52 $Y=1.68 $X2=0 $Y2=0
cc_188 N_A3_M1002_g N_A4_c_287_n 0.00515828f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_189 A3 N_A4_c_287_n 0.0089957f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_190 N_A3_M1006_g N_A_186_531#_c_359_n 6.3924e-19 $X=2.145 $Y=2.865 $X2=0
+ $Y2=0
cc_191 N_A3_M1006_g N_A_186_531#_c_360_n 0.0163489f $X=2.145 $Y=2.865 $X2=0
+ $Y2=0
cc_192 N_A3_c_238_n N_A_186_531#_c_360_n 0.00874908f $X=2.377 $Y=2.185 $X2=0
+ $Y2=0
cc_193 A3 N_A_186_531#_c_360_n 0.0107849f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_194 N_A3_M1006_g N_A_186_531#_c_362_n 5.1591e-19 $X=2.145 $Y=2.865 $X2=0
+ $Y2=0
cc_195 A3 N_A_186_531#_c_362_n 0.00612426f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_196 N_A3_M1006_g N_VPWR_c_406_n 0.001525f $X=2.145 $Y=2.865 $X2=0 $Y2=0
cc_197 N_A3_M1006_g N_VPWR_c_409_n 0.00420792f $X=2.145 $Y=2.865 $X2=0 $Y2=0
cc_198 N_A3_M1006_g N_VPWR_c_404_n 0.0058978f $X=2.145 $Y=2.865 $X2=0 $Y2=0
cc_199 N_A3_M1002_g N_VGND_c_448_n 0.00238543f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_200 A3 N_VGND_c_448_n 0.00154085f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_201 N_A3_M1002_g N_VGND_c_449_n 0.00585385f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_202 N_A3_M1002_g N_VGND_c_452_n 0.0109411f $X=2.255 $Y=0.445 $X2=0 $Y2=0
cc_203 A3 N_VGND_c_452_n 0.0083706f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_204 N_A4_c_288_n N_A_186_531#_c_360_n 0.00447878f $X=2.575 $Y=2.545 $X2=0
+ $Y2=0
cc_205 N_A4_c_290_n N_A_186_531#_c_360_n 0.0034668f $X=2.65 $Y=2.47 $X2=0 $Y2=0
cc_206 N_A4_c_288_n N_A_186_531#_c_362_n 0.0069435f $X=2.575 $Y=2.545 $X2=0
+ $Y2=0
cc_207 N_A4_c_289_n N_A_186_531#_c_362_n 0.0174549f $X=2.925 $Y=2.47 $X2=0 $Y2=0
cc_208 N_A4_c_290_n N_A_186_531#_c_362_n 4.38156e-19 $X=2.65 $Y=2.47 $X2=0 $Y2=0
cc_209 A4 N_A_186_531#_c_362_n 0.00357481f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_210 N_A4_c_288_n N_VPWR_c_406_n 0.0026911f $X=2.575 $Y=2.545 $X2=0 $Y2=0
cc_211 N_A4_c_288_n N_VPWR_c_411_n 0.00413299f $X=2.575 $Y=2.545 $X2=0 $Y2=0
cc_212 N_A4_c_288_n N_VPWR_c_404_n 0.00685448f $X=2.575 $Y=2.545 $X2=0 $Y2=0
cc_213 N_A4_c_289_n N_VPWR_c_404_n 0.00316976f $X=2.925 $Y=2.47 $X2=0 $Y2=0
cc_214 A4 N_VPWR_c_404_n 0.007537f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_215 N_A4_M1004_g N_VGND_c_448_n 0.0107012f $X=2.615 $Y=0.445 $X2=0 $Y2=0
cc_216 N_A4_c_282_n N_VGND_c_448_n 0.00880395f $X=2.925 $Y=0.915 $X2=0 $Y2=0
cc_217 N_A4_M1004_g N_VGND_c_449_n 0.00486043f $X=2.615 $Y=0.445 $X2=0 $Y2=0
cc_218 N_A4_M1004_g N_VGND_c_452_n 0.00444929f $X=2.615 $Y=0.445 $X2=0 $Y2=0
cc_219 N_A4_c_282_n N_VGND_c_452_n 0.00159672f $X=2.925 $Y=0.915 $X2=0 $Y2=0
cc_220 A4 N_VGND_c_452_n 0.00703194f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_221 Y N_VPWR_c_407_n 0.0114541f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_222 Y N_VPWR_c_404_n 0.0101742f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_223 N_Y_c_324_n N_VGND_c_447_n 0.00925747f $X=1.105 $Y=0.925 $X2=0 $Y2=0
cc_224 N_Y_c_325_n N_VGND_c_449_n 0.00832735f $X=1.21 $Y=0.51 $X2=0 $Y2=0
cc_225 N_Y_M1008_d N_VGND_c_452_n 0.00296117f $X=1.07 $Y=0.235 $X2=0 $Y2=0
cc_226 N_Y_c_324_n N_VGND_c_452_n 0.0149317f $X=1.105 $Y=0.925 $X2=0 $Y2=0
cc_227 N_Y_c_325_n N_VGND_c_452_n 0.00769932f $X=1.21 $Y=0.51 $X2=0 $Y2=0
cc_228 Y N_VGND_c_452_n 0.0110404f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_229 N_A_186_531#_c_357_n N_VPWR_c_405_n 0.0139569f $X=1.825 $Y=2.52 $X2=0
+ $Y2=0
cc_230 N_A_186_531#_c_360_n N_VPWR_c_406_n 0.0132936f $X=2.625 $Y=2.52 $X2=0
+ $Y2=0
cc_231 N_A_186_531#_c_356_n N_VPWR_c_407_n 0.00662458f $X=1.07 $Y=2.78 $X2=0
+ $Y2=0
cc_232 N_A_186_531#_c_357_n N_VPWR_c_407_n 0.00305343f $X=1.825 $Y=2.52 $X2=0
+ $Y2=0
cc_233 N_A_186_531#_c_357_n N_VPWR_c_409_n 0.00305343f $X=1.825 $Y=2.52 $X2=0
+ $Y2=0
cc_234 N_A_186_531#_c_359_n N_VPWR_c_409_n 0.00758652f $X=1.93 $Y=2.8 $X2=0
+ $Y2=0
cc_235 N_A_186_531#_c_360_n N_VPWR_c_409_n 0.00305343f $X=2.625 $Y=2.52 $X2=0
+ $Y2=0
cc_236 N_A_186_531#_c_360_n N_VPWR_c_411_n 0.00249315f $X=2.625 $Y=2.52 $X2=0
+ $Y2=0
cc_237 N_A_186_531#_c_362_n N_VPWR_c_411_n 0.00955779f $X=2.79 $Y=2.52 $X2=0
+ $Y2=0
cc_238 N_A_186_531#_c_356_n N_VPWR_c_404_n 0.00671925f $X=1.07 $Y=2.78 $X2=0
+ $Y2=0
cc_239 N_A_186_531#_c_357_n N_VPWR_c_404_n 0.0111075f $X=1.825 $Y=2.52 $X2=0
+ $Y2=0
cc_240 N_A_186_531#_c_359_n N_VPWR_c_404_n 0.00754714f $X=1.93 $Y=2.8 $X2=0
+ $Y2=0
cc_241 N_A_186_531#_c_360_n N_VPWR_c_404_n 0.0100892f $X=2.625 $Y=2.52 $X2=0
+ $Y2=0
cc_242 N_A_186_531#_c_362_n N_VPWR_c_404_n 0.0111741f $X=2.79 $Y=2.52 $X2=0
+ $Y2=0
cc_243 N_VGND_c_452_n A_300_47# 0.00518883f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_244 N_VGND_c_452_n A_372_47# 0.0127373f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_245 N_VGND_c_452_n A_466_47# 0.0060645f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
