* File: sky130_fd_sc_lp__busdrivernovlpsleep_20.spice
* Created: Fri Aug 28 10:13:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__busdrivernovlpsleep_20.pex.spice"
.subckt sky130_fd_sc_lp__busdrivernovlpsleep_20  VNB VPB SLEEP TE_B A VPWR KAPWR
+ Z VGND
* 
* VGND	VGND
* Z	Z
* KAPWR	KAPWR
* VPWR	VPWR
* A	A
* TE_B	TE_B
* SLEEP	SLEEP
* VPB	VPB
* VNB	VNB
MM1030 A_110_47# N_SLEEP_M1030_g N_A_27_47#_M1030_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_SLEEP_M1002_g A_110_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0847 AS=0.0441 PD=0.786667 PS=0.63 NRD=17.136 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75002 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1002_d N_SLEEP_M1013_g N_A_280_47#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1694 AS=0.1176 PD=1.57333 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1045 N_VGND_M1045_d N_SLEEP_M1045_g N_A_280_47#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1045_d N_TE_B_M1008_g N_A_280_47#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1040 N_VGND_M1040_d N_TE_B_M1040_g N_A_280_47#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1063 N_VGND_M1063_d N_A_280_47#_M1063_g N_A_407_491#_M1063_s VNB NSHORT L=0.15
+ W=0.42 AD=0.30975 AS=0.1113 PD=1.895 PS=1.37 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1037 A_1053_47# N_A_280_47#_M1037_g N_VGND_M1063_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.30975 PD=0.63 PS=1.895 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_896_367#_M1014_d N_A_705_367#_M1014_g A_1053_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.18275 AS=0.0441 PD=1.86 PS=0.63 NRD=18.564 NRS=14.28 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1038 N_A_1486_47#_M1038_d N_A_407_491#_M1038_g N_VGND_M1038_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.2226 PD=1.37 PS=2.21 NRD=35.712 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75002.9 A=0.126 P=1.98 MULT=1
MM1050 N_A_1486_47#_M1038_d N_A_407_491#_M1050_g N_VGND_M1050_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.2562 PD=1.37 PS=1.45 NRD=0 NRS=47.136 M=1 R=5.6
+ SA=75000.9 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1003 N_A_1486_47#_M1003_d N_A_M1003_g N_VGND_M1050_s VNB NSHORT L=0.15 W=0.84
+ AD=0.212325 AS=0.2562 PD=1.45 PS=1.45 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1071 N_A_1486_47#_M1003_d N_A_M1071_g N_VGND_M1071_s VNB NSHORT L=0.15 W=0.84
+ AD=0.212325 AS=0.2618 PD=1.45 PS=2.03333 NRD=17.136 NRS=0 M=1 R=5.6 SA=75002.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1020 N_A_2063_47#_M1020_d N_A_407_491#_M1020_g N_VGND_M1071_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1309 PD=0.7 PS=1.01667 NRD=0 NRS=0 M=1 R=2.8
+ SA=75003.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1065 N_VGND_M1065_d N_A_1486_47#_M1065_g N_A_2063_47#_M1020_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_2519_47#_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1575 AS=0.2226 PD=1.215 PS=2.21 NRD=7.848 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1041 N_VGND_M1007_d N_A_M1041_g N_A_2519_47#_M1041_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1575 AS=0.1449 PD=1.215 PS=1.185 NRD=5.712 NRS=9.276 M=1 R=5.6 SA=75000.7
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_2519_47#_M1041_s N_A_2063_47#_M1005_g N_A_705_367#_M1005_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1449 AS=0.1176 PD=1.185 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.2 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1055 N_A_2519_47#_M1055_d N_A_2063_47#_M1055_g N_A_705_367#_M1005_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.2604 AS=0.1176 PD=2.3 PS=1.12 NRD=3.564 NRS=0 M=1 R=5.6
+ SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A_1486_47#_M1000_g N_Z_M1000_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75005.8 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1000_d N_A_1486_47#_M1009_g N_Z_M1009_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75005.4 A=0.096 P=1.58 MULT=1
MM1021 N_VGND_M1021_d N_A_1486_47#_M1021_g N_Z_M1009_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75004.9 A=0.096 P=1.58 MULT=1
MM1025 N_VGND_M1021_d N_A_1486_47#_M1025_g N_Z_M1025_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75004.5 A=0.096 P=1.58 MULT=1
MM1029 N_VGND_M1029_d N_A_1486_47#_M1029_g N_Z_M1025_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.9
+ SB=75004.1 A=0.096 P=1.58 MULT=1
MM1032 N_VGND_M1029_d N_A_1486_47#_M1032_g N_Z_M1032_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.4
+ SB=75003.7 A=0.096 P=1.58 MULT=1
MM1047 N_VGND_M1047_d N_A_1486_47#_M1047_g N_Z_M1032_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.8
+ SB=75003.2 A=0.096 P=1.58 MULT=1
MM1048 N_VGND_M1047_d N_A_1486_47#_M1048_g N_Z_M1048_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.2
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1052 N_VGND_M1052_d N_A_1486_47#_M1052_g N_Z_M1048_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.7
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1056 N_VGND_M1052_d N_A_1486_47#_M1056_g N_Z_M1056_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.1
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1058 N_VGND_M1058_d N_A_1486_47#_M1058_g N_Z_M1056_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.5
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1059 N_VGND_M1058_d N_A_1486_47#_M1059_g N_Z_M1059_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.9
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1062 N_VGND_M1062_d N_A_1486_47#_M1062_g N_Z_M1059_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75005.4
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1073 N_VGND_M1062_d N_A_1486_47#_M1073_g N_Z_M1073_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75005.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1026 N_VPWR_M1026_d N_SLEEP_M1026_g N_A_27_47#_M1026_s VPB PHIGHVT L=0.25 W=1
+ AD=0.190854 AS=0.265 PD=1.63415 PS=2.53 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1006 A_228_491# N_SLEEP_M1006_g N_VPWR_M1026_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.122146 PD=0.85 PS=1.04585 NRD=15.3857 NRS=19.2272 M=1 R=4.26667
+ SA=75000.8 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_280_47#_M1001_d N_TE_B_M1001_g A_228_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1035 N_KAPWR_M1035_d N_A_280_47#_M1035_g N_A_407_491#_M1035_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.251621 AS=0.1696 PD=1.472 PS=1.81 NRD=21.5321 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1011 N_KAPWR_M1035_d N_A_280_47#_M1011_g N_A_705_367#_M1011_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.495379 AS=0.23625 PD=2.898 PS=1.635 NRD=0 NRS=14.8341 M=1
+ R=8.4 SA=75000.7 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1042 N_KAPWR_M1042_d N_A_280_47#_M1042_g N_A_705_367#_M1011_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.23625 PD=1.54 PS=1.635 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.3 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1036 N_KAPWR_M1042_d N_A_27_47#_M1036_g N_A_896_367#_M1036_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1066 N_KAPWR_M1066_d N_A_27_47#_M1066_g N_A_896_367#_M1036_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1049 A_1172_451# N_SLEEP_M1049_g N_VPWR_M1049_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1057 N_A_896_367#_M1057_d N_A_280_47#_M1057_g A_1172_451# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1176 AS=0.0882 PD=1.12 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1027 N_VPWR_M1027_d N_A_705_367#_M1027_g N_A_896_367#_M1057_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1023 N_A_1486_47#_M1023_d N_A_896_367#_M1023_g N_A_1492_367#_M1023_s VPB
+ PHIGHVT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1
+ R=8.4 SA=75000.2 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1067 N_A_1486_47#_M1023_d N_A_896_367#_M1067_g N_A_1492_367#_M1067_s VPB
+ PHIGHVT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1
+ R=8.4 SA=75000.6 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1012 N_A_1492_367#_M1067_s N_A_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1044 N_A_1492_367#_M1044_d N_A_M1044_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1018 A_2033_373# N_A_407_491#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=0.84
+ AD=0.0882 AS=0.2394 PD=1.05 PS=2.25 NRD=11.7215 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1068 N_A_2063_47#_M1068_d N_A_1486_47#_M1068_g A_2033_373# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 N_VPWR_M1015_d N_SLEEP_M1015_g N_A_2345_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1046 N_VPWR_M1046_d N_SLEEP_M1046_g N_A_2345_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1016 N_A_705_367#_M1016_d N_A_M1016_g N_A_2345_367#_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1069 N_A_705_367#_M1016_d N_A_M1069_g N_A_2345_367#_M1069_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1004 N_Z_M1004_d N_A_705_367#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75008.4 A=0.189 P=2.82 MULT=1
MM1010 N_Z_M1004_d N_A_705_367#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75007.9 A=0.189 P=2.82 MULT=1
MM1017 N_Z_M1017_d N_A_705_367#_M1017_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75007.5 A=0.189 P=2.82 MULT=1
MM1019 N_Z_M1017_d N_A_705_367#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75007.1 A=0.189 P=2.82 MULT=1
MM1022 N_Z_M1022_d N_A_705_367#_M1022_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75006.7 A=0.189 P=2.82 MULT=1
MM1024 N_Z_M1022_d N_A_705_367#_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75006.2 A=0.189 P=2.82 MULT=1
MM1028 N_Z_M1028_d N_A_705_367#_M1028_g N_VPWR_M1024_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75005.8 A=0.189 P=2.82 MULT=1
MM1031 N_Z_M1028_d N_A_705_367#_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75005.4 A=0.189 P=2.82 MULT=1
MM1033 N_Z_M1033_d N_A_705_367#_M1033_g N_VPWR_M1031_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1034 N_Z_M1033_d N_A_705_367#_M1034_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1039 N_Z_M1039_d N_A_705_367#_M1039_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1043 N_Z_M1039_d N_A_705_367#_M1043_g N_VPWR_M1043_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.9
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1051 N_Z_M1051_d N_A_705_367#_M1051_g N_VPWR_M1043_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.3
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1053 N_Z_M1051_d N_A_705_367#_M1053_g N_VPWR_M1053_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.8
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1054 N_Z_M1054_d N_A_705_367#_M1054_g N_VPWR_M1053_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1060 N_Z_M1054_d N_A_705_367#_M1060_g N_VPWR_M1060_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1061 N_Z_M1061_d N_A_705_367#_M1061_g N_VPWR_M1060_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1064 N_Z_M1061_d N_A_705_367#_M1064_g N_VPWR_M1064_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1070 N_Z_M1070_d N_A_705_367#_M1070_g N_VPWR_M1064_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1072 N_Z_M1070_d N_A_705_367#_M1072_g N_VPWR_M1072_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75008.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX74_noxref VNB VPB NWDIODE A=44.5735 P=51.53
*
.include "sky130_fd_sc_lp__busdrivernovlpsleep_20.pxi.spice"
*
.ends
*
*
