* File: sky130_fd_sc_lp__nor3_1.spice
* Created: Fri Aug 28 10:55:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor3_1.pex.spice"
.subckt sky130_fd_sc_lp__nor3_1  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75001.1 A=0.126
+ P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.84 AD=0.1344
+ AS=0.1176 PD=1.16 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.6 SB=75000.7
+ A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_C_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1344 PD=2.21 PS=1.16 NRD=0 NRS=2.856 M=1 R=5.6 SA=75001.1 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1005 A_110_367# N_A_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26 AD=0.1953
+ AS=0.3339 PD=1.57 PS=3.05 NRD=15.6221 NRS=0 M=1 R=8.4 SA=75000.2 SB=75001.1
+ A=0.189 P=2.82 MULT=1
MM1004 A_202_367# N_B_M1004_g A_110_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.1827
+ AS=0.1953 PD=1.55 PS=1.57 NRD=14.0658 NRS=15.6221 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g A_202_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.3339
+ AS=0.1827 PD=3.05 PS=1.55 NRD=0 NRS=14.0658 M=1 R=8.4 SA=75001.1 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.2895 P=8.33
c_37 VPB 0 1.47358e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__nor3_1.pxi.spice"
*
.ends
*
*
