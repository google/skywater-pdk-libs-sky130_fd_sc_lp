* File: sky130_fd_sc_lp__inv_8.pxi.spice
* Created: Wed Sep  2 09:56:05 2020
* 
x_PM_SKY130_FD_SC_LP__INV_8%A N_A_M1001_g N_A_M1000_g N_A_M1004_g N_A_M1002_g
+ N_A_M1005_g N_A_M1003_g N_A_M1007_g N_A_M1006_g N_A_M1010_g N_A_M1008_g
+ N_A_M1012_g N_A_M1009_g N_A_M1013_g N_A_M1011_g N_A_M1014_g N_A_M1015_g
+ N_A_c_102_n N_A_c_103_n A N_A_c_105_n PM_SKY130_FD_SC_LP__INV_8%A
x_PM_SKY130_FD_SC_LP__INV_8%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_M1006_d
+ N_VPWR_M1009_d N_VPWR_M1015_d N_VPWR_c_229_n N_VPWR_c_230_n N_VPWR_c_231_n
+ N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n
+ N_VPWR_c_237_n N_VPWR_c_238_n N_VPWR_c_239_n VPWR N_VPWR_c_240_n
+ N_VPWR_c_241_n N_VPWR_c_242_n N_VPWR_c_243_n N_VPWR_c_228_n
+ PM_SKY130_FD_SC_LP__INV_8%VPWR
x_PM_SKY130_FD_SC_LP__INV_8%Y N_Y_M1001_s N_Y_M1005_s N_Y_M1010_s N_Y_M1013_s
+ N_Y_M1000_s N_Y_M1003_s N_Y_M1008_s N_Y_M1011_s N_Y_c_291_n N_Y_c_292_n
+ N_Y_c_293_n N_Y_c_304_n N_Y_c_305_n N_Y_c_416_p N_Y_c_387_n N_Y_c_294_n
+ N_Y_c_306_n N_Y_c_411_p N_Y_c_391_n N_Y_c_333_n N_Y_c_307_n N_Y_c_417_p
+ N_Y_c_395_n N_Y_c_295_n N_Y_c_308_n N_Y_c_418_p N_Y_c_399_n N_Y_c_296_n
+ N_Y_c_309_n N_Y_c_297_n N_Y_c_310_n N_Y_c_298_n N_Y_c_311_n N_Y_c_299_n
+ N_Y_c_312_n N_Y_c_300_n N_Y_c_313_n Y Y N_Y_c_301_n Y
+ PM_SKY130_FD_SC_LP__INV_8%Y
x_PM_SKY130_FD_SC_LP__INV_8%VGND N_VGND_M1001_d N_VGND_M1004_d N_VGND_M1007_d
+ N_VGND_M1012_d N_VGND_M1014_d N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n
+ N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n
+ N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n VGND N_VGND_c_439_n
+ N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n
+ PM_SKY130_FD_SC_LP__INV_8%VGND
cc_1 VNB N_A_M1001_g 0.0272298f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.655
cc_2 VNB N_A_M1000_g 5.36722e-19 $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=2.465
cc_3 VNB N_A_M1004_g 0.021612f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=0.655
cc_4 VNB N_A_M1002_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=2.465
cc_5 VNB N_A_M1005_g 0.0216041f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=0.655
cc_6 VNB N_A_M1003_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.465
cc_7 VNB N_A_M1007_g 0.0221104f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=0.655
cc_8 VNB N_A_M1006_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=2.465
cc_9 VNB N_A_M1010_g 0.0227f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=0.655
cc_10 VNB N_A_M1008_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=2.465
cc_11 VNB N_A_M1012_g 0.0216061f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=0.655
cc_12 VNB N_A_M1009_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=2.465
cc_13 VNB N_A_M1013_g 0.0215926f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=0.655
cc_14 VNB N_A_M1011_g 4.57539e-19 $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.465
cc_15 VNB N_A_M1014_g 0.0268386f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=0.655
cc_16 VNB N_A_M1015_g 5.01157e-19 $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=2.465
cc_17 VNB N_A_c_102_n 0.00176541f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.49
cc_18 VNB N_A_c_103_n 0.00185932f $X=-0.19 $Y=-0.245 $X2=3.65 $Y2=1.48
cc_19 VNB A 0.00378912f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_20 VNB N_A_c_105_n 0.180983f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=1.48
cc_21 VNB N_VPWR_c_228_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.48
cc_22 VNB N_Y_c_291_n 0.0214285f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=0.655
cc_23 VNB N_Y_c_292_n 0.00837668f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=0.655
cc_24 VNB N_Y_c_293_n 0.0149163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_294_n 0.00244948f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=1.315
cc_26 VNB N_Y_c_295_n 0.00269389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_296_n 0.00232031f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.48
cc_28 VNB N_Y_c_297_n 0.00214052f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.48
cc_29 VNB N_Y_c_298_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.48
cc_30 VNB N_Y_c_299_n 0.00347338f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=1.48
cc_31 VNB N_Y_c_300_n 0.00210048f $X=-0.19 $Y=-0.245 $X2=2.212 $Y2=1.295
cc_32 VNB N_Y_c_301_n 0.0127485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB Y 0.0230605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_428_n 0.0287407f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=0.655
cc_35 VNB N_VGND_c_429_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.465
cc_36 VNB N_VGND_c_430_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_431_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_432_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_433_n 0.0142549f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=0.655
cc_40 VNB N_VGND_c_434_n 0.0287404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_435_n 0.013281f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=2.465
cc_42 VNB N_VGND_c_436_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_437_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=1.315
cc_44 VNB N_VGND_c_438_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=0.655
cc_45 VNB N_VGND_c_439_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_440_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=1.315
cc_47 VNB N_VGND_c_441_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=2.465
cc_48 VNB N_VGND_c_442_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.49
cc_49 VNB N_VGND_c_443_n 0.242138f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.49
cc_50 VPB N_A_M1000_g 0.0238187f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=2.465
cc_51 VPB N_A_M1002_g 0.0191131f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=2.465
cc_52 VPB N_A_M1003_g 0.0191131f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=2.465
cc_53 VPB N_A_M1006_g 0.0191131f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=2.465
cc_54 VPB N_A_M1008_g 0.0191131f $X=-0.19 $Y=1.655 $X2=2.45 $Y2=2.465
cc_55 VPB N_A_M1009_g 0.0191131f $X=-0.19 $Y=1.655 $X2=2.88 $Y2=2.465
cc_56 VPB N_A_M1011_g 0.0190938f $X=-0.19 $Y=1.655 $X2=3.31 $Y2=2.465
cc_57 VPB N_A_M1015_g 0.0234235f $X=-0.19 $Y=1.655 $X2=3.74 $Y2=2.465
cc_58 VPB N_VPWR_c_229_n 0.0418562f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=0.655
cc_59 VPB N_VPWR_c_230_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_231_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_232_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_233_n 0.00400996f $X=-0.19 $Y=1.655 $X2=2.45 $Y2=2.465
cc_63 VPB N_VPWR_c_234_n 0.014229f $X=-0.19 $Y=1.655 $X2=2.88 $Y2=0.655
cc_64 VPB N_VPWR_c_235_n 0.042227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_236_n 0.013281f $X=-0.19 $Y=1.655 $X2=3.31 $Y2=1.315
cc_66 VPB N_VPWR_c_237_n 0.00564836f $X=-0.19 $Y=1.655 $X2=3.31 $Y2=0.655
cc_67 VPB N_VPWR_c_238_n 0.0166024f $X=-0.19 $Y=1.655 $X2=3.31 $Y2=0.655
cc_68 VPB N_VPWR_c_239_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_240_n 0.0166024f $X=-0.19 $Y=1.655 $X2=3.74 $Y2=2.465
cc_70 VPB N_VPWR_c_241_n 0.0166024f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.48
cc_71 VPB N_VPWR_c_242_n 0.00497514f $X=-0.19 $Y=1.655 $X2=2.365 $Y2=1.485
cc_72 VPB N_VPWR_c_243_n 0.00497514f $X=-0.19 $Y=1.655 $X2=3.65 $Y2=1.48
cc_73 VPB N_VPWR_c_228_n 0.0585537f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.48
cc_74 VPB N_Y_c_291_n 0.00514138f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=0.655
cc_75 VPB N_Y_c_304_n 0.0080617f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=1.645
cc_76 VPB N_Y_c_305_n 0.0148315f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=2.465
cc_77 VPB N_Y_c_306_n 0.00240582f $X=-0.19 $Y=1.655 $X2=2.88 $Y2=0.655
cc_78 VPB N_Y_c_307_n 0.00239258f $X=-0.19 $Y=1.655 $X2=3.74 $Y2=1.315
cc_79 VPB N_Y_c_308_n 0.00240582f $X=-0.19 $Y=1.655 $X2=1.95 $Y2=1.48
cc_80 VPB N_Y_c_309_n 0.0147951f $X=-0.19 $Y=1.655 $X2=1.95 $Y2=1.48
cc_81 VPB N_Y_c_310_n 0.00210233f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.48
cc_82 VPB N_Y_c_311_n 0.00210233f $X=-0.19 $Y=1.655 $X2=2.88 $Y2=1.48
cc_83 VPB N_Y_c_312_n 0.00208355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_Y_c_313_n 0.00210233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB Y 0.00537816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 N_A_M1000_g N_VPWR_c_229_n 0.00343774f $X=0.73 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_VPWR_c_230_n 0.0016342f $X=1.16 $Y=2.465 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_VPWR_c_230_n 0.0016342f $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VPWR_c_231_n 0.00585385f $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A_M1006_g N_VPWR_c_231_n 0.00585385f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_91 N_A_M1006_g N_VPWR_c_232_n 0.0016342f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A_M1008_g N_VPWR_c_232_n 0.0016342f $X=2.45 $Y=2.465 $X2=0 $Y2=0
cc_93 N_A_M1009_g N_VPWR_c_233_n 0.0016342f $X=2.88 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_M1011_g N_VPWR_c_233_n 0.0016342f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A_M1015_g N_VPWR_c_235_n 0.00343774f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A_M1000_g N_VPWR_c_238_n 0.00585385f $X=0.73 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A_M1002_g N_VPWR_c_238_n 0.00585385f $X=1.16 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_M1008_g N_VPWR_c_240_n 0.00585385f $X=2.45 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_M1009_g N_VPWR_c_240_n 0.00585385f $X=2.88 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_M1011_g N_VPWR_c_241_n 0.00585385f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A_M1015_g N_VPWR_c_241_n 0.00585385f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_M1000_g N_VPWR_c_228_n 0.0117311f $X=0.73 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_M1002_g N_VPWR_c_228_n 0.0106302f $X=1.16 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A_M1003_g N_VPWR_c_228_n 0.0106302f $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A_M1006_g N_VPWR_c_228_n 0.0106302f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_M1008_g N_VPWR_c_228_n 0.0106302f $X=2.45 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_M1009_g N_VPWR_c_228_n 0.0106302f $X=2.88 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_M1011_g N_VPWR_c_228_n 0.0106302f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_M1015_g N_VPWR_c_228_n 0.0116481f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A_M1001_g N_Y_c_291_n 0.00265692f $X=0.73 $Y=0.655 $X2=0 $Y2=0
cc_111 N_A_M1000_g N_Y_c_291_n 0.00292529f $X=0.73 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_c_102_n N_Y_c_291_n 0.0150242f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_113 N_A_c_105_n N_Y_c_291_n 0.00720148f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_114 N_A_M1001_g N_Y_c_292_n 0.0170045f $X=0.73 $Y=0.655 $X2=0 $Y2=0
cc_115 N_A_c_102_n N_Y_c_292_n 0.0263361f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_116 N_A_c_105_n N_Y_c_292_n 0.00563276f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_117 N_A_M1000_g N_Y_c_304_n 0.016309f $X=0.73 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_c_102_n N_Y_c_304_n 0.0275222f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_119 N_A_c_105_n N_Y_c_304_n 0.00553508f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_120 N_A_M1004_g N_Y_c_294_n 0.0150885f $X=1.16 $Y=0.655 $X2=0 $Y2=0
cc_121 N_A_M1005_g N_Y_c_294_n 0.0146529f $X=1.59 $Y=0.655 $X2=0 $Y2=0
cc_122 N_A_c_102_n N_Y_c_294_n 0.0402443f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_123 N_A_c_105_n N_Y_c_294_n 0.00244902f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_124 N_A_M1002_g N_Y_c_306_n 0.0144397f $X=1.16 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_M1003_g N_Y_c_306_n 0.0144397f $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_c_102_n N_Y_c_306_n 0.0420698f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_127 N_A_c_105_n N_Y_c_306_n 0.00240656f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_128 N_A_M1007_g N_Y_c_333_n 0.0108185f $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_129 N_A_M1010_g N_Y_c_333_n 0.0110803f $X=2.45 $Y=0.655 $X2=0 $Y2=0
cc_130 N_A_c_102_n N_Y_c_333_n 0.00405943f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_131 N_A_c_103_n N_Y_c_333_n 0.00555683f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_132 A N_Y_c_333_n 0.0202395f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_133 N_A_c_105_n N_Y_c_333_n 4.82597e-19 $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_134 N_A_M1006_g N_Y_c_307_n 0.0144246f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_M1008_g N_Y_c_307_n 0.0144397f $X=2.45 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_c_102_n N_Y_c_307_n 0.00854563f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_137 N_A_c_103_n N_Y_c_307_n 0.0117061f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_138 A N_Y_c_307_n 0.0232084f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A_c_105_n N_Y_c_307_n 0.00240522f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_140 N_A_M1012_g N_Y_c_295_n 0.013601f $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_141 N_A_M1013_g N_Y_c_295_n 0.0150272f $X=3.31 $Y=0.655 $X2=0 $Y2=0
cc_142 N_A_c_103_n N_Y_c_295_n 0.0422712f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_143 N_A_c_105_n N_Y_c_295_n 0.00243542f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_144 N_A_M1009_g N_Y_c_308_n 0.0144397f $X=2.88 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1011_g N_Y_c_308_n 0.0144397f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_c_103_n N_Y_c_308_n 0.0422336f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_147 N_A_c_105_n N_Y_c_308_n 0.00240656f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_148 N_A_M1014_g N_Y_c_296_n 0.0166975f $X=3.74 $Y=0.655 $X2=0 $Y2=0
cc_149 N_A_c_103_n N_Y_c_296_n 0.0109821f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_150 N_A_M1015_g N_Y_c_309_n 0.0160634f $X=3.74 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_c_103_n N_Y_c_309_n 0.0109821f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_152 N_A_c_102_n N_Y_c_297_n 0.020245f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_153 N_A_c_105_n N_Y_c_297_n 0.00255521f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_154 N_A_c_102_n N_Y_c_310_n 0.0211331f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_155 N_A_c_105_n N_Y_c_310_n 0.00250529f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_156 N_A_M1007_g N_Y_c_298_n 0.00197629f $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_157 N_A_c_102_n N_Y_c_298_n 0.0167405f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_158 A N_Y_c_298_n 0.00461278f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A_c_105_n N_Y_c_298_n 0.00255521f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_160 N_A_c_102_n N_Y_c_311_n 0.0211331f $X=2.06 $Y=1.49 $X2=0 $Y2=0
cc_161 N_A_c_105_n N_Y_c_311_n 0.00250529f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_162 N_A_M1010_g N_Y_c_299_n 0.00188389f $X=2.45 $Y=0.655 $X2=0 $Y2=0
cc_163 N_A_M1012_g N_Y_c_299_n 7.32812e-19 $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_164 N_A_c_103_n N_Y_c_299_n 0.0210412f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_165 A N_Y_c_299_n 0.00446821f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_166 N_A_c_105_n N_Y_c_299_n 0.00253619f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_167 N_A_c_103_n N_Y_c_312_n 0.0212044f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_168 N_A_c_105_n N_Y_c_312_n 0.00250529f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_169 N_A_c_103_n N_Y_c_300_n 0.0212043f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_170 N_A_c_105_n N_Y_c_300_n 0.00253619f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_171 N_A_c_103_n N_Y_c_313_n 0.0212044f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_172 N_A_c_105_n N_Y_c_313_n 0.00250529f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_173 N_A_M1014_g Y 0.00658014f $X=3.74 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A_c_103_n Y 0.0162257f $X=3.65 $Y=1.48 $X2=0 $Y2=0
cc_175 N_A_c_105_n Y 0.00792033f $X=3.74 $Y=1.48 $X2=0 $Y2=0
cc_176 N_A_M1001_g N_VGND_c_428_n 0.00343774f $X=0.73 $Y=0.655 $X2=0 $Y2=0
cc_177 N_A_M1004_g N_VGND_c_429_n 0.0016342f $X=1.16 $Y=0.655 $X2=0 $Y2=0
cc_178 N_A_M1005_g N_VGND_c_429_n 0.0016342f $X=1.59 $Y=0.655 $X2=0 $Y2=0
cc_179 N_A_M1005_g N_VGND_c_430_n 0.00585385f $X=1.59 $Y=0.655 $X2=0 $Y2=0
cc_180 N_A_M1007_g N_VGND_c_430_n 0.00585385f $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_181 N_A_M1007_g N_VGND_c_431_n 0.0018833f $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_182 N_A_M1010_g N_VGND_c_431_n 0.0018833f $X=2.45 $Y=0.655 $X2=0 $Y2=0
cc_183 N_A_M1012_g N_VGND_c_432_n 0.0016342f $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_184 N_A_M1013_g N_VGND_c_432_n 0.0016342f $X=3.31 $Y=0.655 $X2=0 $Y2=0
cc_185 N_A_M1014_g N_VGND_c_434_n 0.00343774f $X=3.74 $Y=0.655 $X2=0 $Y2=0
cc_186 N_A_M1001_g N_VGND_c_437_n 0.00585385f $X=0.73 $Y=0.655 $X2=0 $Y2=0
cc_187 N_A_M1004_g N_VGND_c_437_n 0.00585385f $X=1.16 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A_M1010_g N_VGND_c_439_n 0.00585385f $X=2.45 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A_M1012_g N_VGND_c_439_n 0.00585385f $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_190 N_A_M1013_g N_VGND_c_440_n 0.00585385f $X=3.31 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A_M1014_g N_VGND_c_440_n 0.00585385f $X=3.74 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A_M1001_g N_VGND_c_443_n 0.0117311f $X=0.73 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A_M1004_g N_VGND_c_443_n 0.0106302f $X=1.16 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A_M1005_g N_VGND_c_443_n 0.0106302f $X=1.59 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A_M1007_g N_VGND_c_443_n 0.00624036f $X=2.02 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A_M1010_g N_VGND_c_443_n 0.00624036f $X=2.45 $Y=0.655 $X2=0 $Y2=0
cc_197 N_A_M1012_g N_VGND_c_443_n 0.0106302f $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_198 N_A_M1013_g N_VGND_c_443_n 0.0106302f $X=3.31 $Y=0.655 $X2=0 $Y2=0
cc_199 N_A_M1014_g N_VGND_c_443_n 0.0116481f $X=3.74 $Y=0.655 $X2=0 $Y2=0
cc_200 N_VPWR_c_228_n N_Y_M1000_s 0.003017f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_228_n N_Y_M1003_s 0.003017f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_c_228_n N_Y_M1008_s 0.003017f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_203 N_VPWR_c_228_n N_Y_M1011_s 0.003017f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_M1000_d N_Y_c_304_n 0.00299978f $X=0.37 $Y=1.835 $X2=0 $Y2=0
cc_205 N_VPWR_c_229_n N_Y_c_304_n 0.0193144f $X=0.515 $Y=2.27 $X2=0 $Y2=0
cc_206 N_VPWR_c_238_n N_Y_c_387_n 0.0149362f $X=1.245 $Y=3.33 $X2=0 $Y2=0
cc_207 N_VPWR_c_228_n N_Y_c_387_n 0.0100304f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_208 N_VPWR_M1002_d N_Y_c_306_n 0.00176461f $X=1.235 $Y=1.835 $X2=0 $Y2=0
cc_209 N_VPWR_c_230_n N_Y_c_306_n 0.0135055f $X=1.375 $Y=2.26 $X2=0 $Y2=0
cc_210 N_VPWR_c_231_n N_Y_c_391_n 0.0149362f $X=2.105 $Y=3.33 $X2=0 $Y2=0
cc_211 N_VPWR_c_228_n N_Y_c_391_n 0.0100304f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_M1006_d N_Y_c_307_n 0.00176461f $X=2.095 $Y=1.835 $X2=0 $Y2=0
cc_213 N_VPWR_c_232_n N_Y_c_307_n 0.0135055f $X=2.235 $Y=2.26 $X2=0 $Y2=0
cc_214 N_VPWR_c_240_n N_Y_c_395_n 0.0149362f $X=2.965 $Y=3.33 $X2=0 $Y2=0
cc_215 N_VPWR_c_228_n N_Y_c_395_n 0.0100304f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_M1009_d N_Y_c_308_n 0.00176461f $X=2.955 $Y=1.835 $X2=0 $Y2=0
cc_217 N_VPWR_c_233_n N_Y_c_308_n 0.0135055f $X=3.095 $Y=2.26 $X2=0 $Y2=0
cc_218 N_VPWR_c_241_n N_Y_c_399_n 0.0149362f $X=3.825 $Y=3.33 $X2=0 $Y2=0
cc_219 N_VPWR_c_228_n N_Y_c_399_n 0.0100304f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_220 N_VPWR_M1015_d N_Y_c_309_n 0.00298626f $X=3.815 $Y=1.835 $X2=0 $Y2=0
cc_221 N_VPWR_c_235_n N_Y_c_309_n 0.0213059f $X=3.955 $Y=2.26 $X2=0 $Y2=0
cc_222 N_Y_c_292_n N_VGND_M1001_d 0.00259223f $X=0.815 $Y=1.13 $X2=-0.19
+ $Y2=-0.245
cc_223 N_Y_c_294_n N_VGND_M1004_d 0.00176461f $X=1.675 $Y=1.13 $X2=0 $Y2=0
cc_224 N_Y_c_333_n N_VGND_M1007_d 0.00332607f $X=2.535 $Y=0.905 $X2=0 $Y2=0
cc_225 N_Y_c_295_n N_VGND_M1012_d 0.00176461f $X=3.395 $Y=1.13 $X2=0 $Y2=0
cc_226 N_Y_c_296_n N_VGND_M1014_d 0.00119058f $X=3.985 $Y=1.13 $X2=0 $Y2=0
cc_227 N_Y_c_301_n N_VGND_M1014_d 0.00144697f $X=4.105 $Y=1.215 $X2=0 $Y2=0
cc_228 N_Y_c_292_n N_VGND_c_428_n 0.0201545f $X=0.815 $Y=1.13 $X2=0 $Y2=0
cc_229 N_Y_c_294_n N_VGND_c_429_n 0.0135055f $X=1.675 $Y=1.13 $X2=0 $Y2=0
cc_230 N_Y_c_411_p N_VGND_c_430_n 0.0149362f $X=1.805 $Y=0.465 $X2=0 $Y2=0
cc_231 N_Y_c_333_n N_VGND_c_431_n 0.0131862f $X=2.535 $Y=0.905 $X2=0 $Y2=0
cc_232 N_Y_c_295_n N_VGND_c_432_n 0.0135055f $X=3.395 $Y=1.13 $X2=0 $Y2=0
cc_233 N_Y_c_296_n N_VGND_c_434_n 0.00915704f $X=3.985 $Y=1.13 $X2=0 $Y2=0
cc_234 N_Y_c_301_n N_VGND_c_434_n 0.0121489f $X=4.105 $Y=1.215 $X2=0 $Y2=0
cc_235 N_Y_c_416_p N_VGND_c_437_n 0.0149362f $X=0.945 $Y=0.465 $X2=0 $Y2=0
cc_236 N_Y_c_417_p N_VGND_c_439_n 0.0149362f $X=2.665 $Y=0.465 $X2=0 $Y2=0
cc_237 N_Y_c_418_p N_VGND_c_440_n 0.0149362f $X=3.525 $Y=0.465 $X2=0 $Y2=0
cc_238 N_Y_M1001_s N_VGND_c_443_n 0.003017f $X=0.805 $Y=0.235 $X2=0 $Y2=0
cc_239 N_Y_M1005_s N_VGND_c_443_n 0.00268963f $X=1.665 $Y=0.235 $X2=0 $Y2=0
cc_240 N_Y_M1010_s N_VGND_c_443_n 0.00268963f $X=2.525 $Y=0.235 $X2=0 $Y2=0
cc_241 N_Y_M1013_s N_VGND_c_443_n 0.003017f $X=3.385 $Y=0.235 $X2=0 $Y2=0
cc_242 N_Y_c_416_p N_VGND_c_443_n 0.0100304f $X=0.945 $Y=0.465 $X2=0 $Y2=0
cc_243 N_Y_c_411_p N_VGND_c_443_n 0.0100304f $X=1.805 $Y=0.465 $X2=0 $Y2=0
cc_244 N_Y_c_333_n N_VGND_c_443_n 0.0105538f $X=2.535 $Y=0.905 $X2=0 $Y2=0
cc_245 N_Y_c_417_p N_VGND_c_443_n 0.0100304f $X=2.665 $Y=0.465 $X2=0 $Y2=0
cc_246 N_Y_c_418_p N_VGND_c_443_n 0.0100304f $X=3.525 $Y=0.465 $X2=0 $Y2=0
