* File: sky130_fd_sc_lp__mux2i_4.pex.spice
* Created: Wed Sep  2 10:01:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2I_4%A0 3 7 11 15 19 23 27 31 33 34 35 56 57
c77 19 0 4.56457e-20 $X=1.415 $Y=0.765
r78 55 57 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=1.55 $Y=1.51
+ $X2=1.845 $Y2=1.51
r79 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.51 $X2=1.55 $Y2=1.51
r80 53 55 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.415 $Y=1.51
+ $X2=1.55 $Y2=1.51
r81 52 56 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.21 $Y=1.587
+ $X2=1.55 $Y2=1.587
r82 51 53 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.21 $Y=1.51
+ $X2=1.415 $Y2=1.51
r83 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.51 $X2=1.21 $Y2=1.51
r84 49 51 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.985 $Y=1.51
+ $X2=1.21 $Y2=1.51
r85 48 49 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=0.985 $Y2=1.51
r86 46 48 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.87 $Y=1.51
+ $X2=0.905 $Y2=1.51
r87 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.87
+ $Y=1.51 $X2=0.87 $Y2=1.51
r88 44 46 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=0.555 $Y=1.51
+ $X2=0.87 $Y2=1.51
r89 42 44 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.53 $Y=1.51
+ $X2=0.555 $Y2=1.51
r90 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.51 $X2=0.53 $Y2=1.51
r91 39 42 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.475 $Y=1.51
+ $X2=0.53 $Y2=1.51
r92 35 52 0.354598 $w=3.23e-07 $l=1e-08 $layer=LI1_cond $X=1.2 $Y=1.587 $X2=1.21
+ $Y2=1.587
r93 35 47 11.7017 $w=3.23e-07 $l=3.3e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=0.87 $Y2=1.587
r94 34 47 5.31897 $w=3.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=0.87 $Y2=1.587
r95 34 43 6.73736 $w=3.23e-07 $l=1.9e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=0.53 $Y2=1.587
r96 33 43 10.2833 $w=3.23e-07 $l=2.9e-07 $layer=LI1_cond $X=0.24 $Y=1.587
+ $X2=0.53 $Y2=1.587
r97 29 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.675
+ $X2=1.845 $Y2=1.51
r98 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.845 $Y=1.675
+ $X2=1.845 $Y2=2.465
r99 25 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.345
+ $X2=1.845 $Y2=1.51
r100 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.845 $Y=1.345
+ $X2=1.845 $Y2=0.765
r101 21 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.675
+ $X2=1.415 $Y2=1.51
r102 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.415 $Y=1.675
+ $X2=1.415 $Y2=2.465
r103 17 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.345
+ $X2=1.415 $Y2=1.51
r104 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.415 $Y=1.345
+ $X2=1.415 $Y2=0.765
r105 13 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.675
+ $X2=0.985 $Y2=1.51
r106 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.985 $Y=1.675
+ $X2=0.985 $Y2=2.465
r107 9 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=1.51
r108 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=0.765
r109 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.675
+ $X2=0.555 $Y2=1.51
r110 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.555 $Y=1.675
+ $X2=0.555 $Y2=2.465
r111 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=1.51
r112 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%A1 3 7 11 15 19 23 27 31 33 34 35 51 52
c70 3 0 3.64334e-20 $X=2.275 $Y=0.765
r71 50 52 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=3.61 $Y=1.51
+ $X2=3.885 $Y2=1.51
r72 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.61
+ $Y=1.51 $X2=3.61 $Y2=1.51
r73 48 50 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.565 $Y=1.51
+ $X2=3.61 $Y2=1.51
r74 47 48 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.295 $Y=1.51
+ $X2=3.565 $Y2=1.51
r75 46 47 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.135 $Y=1.51
+ $X2=3.295 $Y2=1.51
r76 45 46 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=2.865 $Y=1.51
+ $X2=3.135 $Y2=1.51
r77 44 45 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.705 $Y=1.51
+ $X2=2.865 $Y2=1.51
r78 42 44 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=2.59 $Y=1.51
+ $X2=2.705 $Y2=1.51
r79 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.59
+ $Y=1.51 $X2=2.59 $Y2=1.51
r80 39 42 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=2.275 $Y=1.51
+ $X2=2.59 $Y2=1.51
r81 35 51 0.271163 $w=4.23e-07 $l=1e-08 $layer=LI1_cond $X=3.6 $Y=1.547 $X2=3.61
+ $Y2=1.547
r82 34 35 13.0158 $w=4.23e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.547
+ $X2=3.6 $Y2=1.547
r83 33 34 13.0158 $w=4.23e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.547
+ $X2=3.12 $Y2=1.547
r84 33 43 1.35582 $w=4.23e-07 $l=5e-08 $layer=LI1_cond $X=2.64 $Y=1.547 $X2=2.59
+ $Y2=1.547
r85 29 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.885 $Y=1.345
+ $X2=3.885 $Y2=1.51
r86 29 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.885 $Y=1.345
+ $X2=3.885 $Y2=0.765
r87 25 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=1.675
+ $X2=3.565 $Y2=1.51
r88 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.565 $Y=1.675
+ $X2=3.565 $Y2=2.465
r89 21 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.345
+ $X2=3.295 $Y2=1.51
r90 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.295 $Y=1.345
+ $X2=3.295 $Y2=0.765
r91 17 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.135 $Y=1.675
+ $X2=3.135 $Y2=1.51
r92 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.135 $Y=1.675
+ $X2=3.135 $Y2=2.465
r93 13 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.345
+ $X2=2.865 $Y2=1.51
r94 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.865 $Y=1.345
+ $X2=2.865 $Y2=0.765
r95 9 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.675
+ $X2=2.705 $Y2=1.51
r96 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.705 $Y=1.675
+ $X2=2.705 $Y2=2.465
r97 5 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=1.675
+ $X2=2.275 $Y2=1.51
r98 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.275 $Y=1.675
+ $X2=2.275 $Y2=2.465
r99 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=1.345
+ $X2=2.275 $Y2=1.51
r100 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.275 $Y=1.345
+ $X2=2.275 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%S 3 7 11 15 19 23 27 31 33 35 36 38 40 43 46
+ 47 48 49 50 51 74 96
c132 74 0 1.35208e-19 $X=6.735 $Y=1.51
c133 43 0 2.6512e-20 $X=9.075 $Y=1.5
r134 74 75 1.47401 $w=3.27e-07 $l=1e-08 $layer=POLY_cond $X=6.735 $Y=1.51
+ $X2=6.745 $Y2=1.51
r135 72 74 26.5321 $w=3.27e-07 $l=1.8e-07 $layer=POLY_cond $X=6.555 $Y=1.51
+ $X2=6.735 $Y2=1.51
r136 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.555
+ $Y=1.51 $X2=6.555 $Y2=1.51
r137 70 72 36.8502 $w=3.27e-07 $l=2.5e-07 $layer=POLY_cond $X=6.305 $Y=1.51
+ $X2=6.555 $Y2=1.51
r138 69 70 1.47401 $w=3.27e-07 $l=1e-08 $layer=POLY_cond $X=6.295 $Y=1.51
+ $X2=6.305 $Y2=1.51
r139 67 69 11.792 $w=3.27e-07 $l=8e-08 $layer=POLY_cond $X=6.215 $Y=1.51
+ $X2=6.295 $Y2=1.51
r140 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.215
+ $Y=1.51 $X2=6.215 $Y2=1.51
r141 65 67 50.1162 $w=3.27e-07 $l=3.4e-07 $layer=POLY_cond $X=5.875 $Y=1.51
+ $X2=6.215 $Y2=1.51
r142 64 65 1.47401 $w=3.27e-07 $l=1e-08 $layer=POLY_cond $X=5.865 $Y=1.51
+ $X2=5.875 $Y2=1.51
r143 62 64 48.6422 $w=3.27e-07 $l=3.3e-07 $layer=POLY_cond $X=5.535 $Y=1.51
+ $X2=5.865 $Y2=1.51
r144 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.535
+ $Y=1.51 $X2=5.535 $Y2=1.51
r145 60 62 13.2661 $w=3.27e-07 $l=9e-08 $layer=POLY_cond $X=5.445 $Y=1.51
+ $X2=5.535 $Y2=1.51
r146 59 60 1.47401 $w=3.27e-07 $l=1e-08 $layer=POLY_cond $X=5.435 $Y=1.51
+ $X2=5.445 $Y2=1.51
r147 51 96 7.89897 $w=5.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.96 $Y=1.68
+ $X2=7.045 $Y2=1.68
r148 51 73 7.49725 $w=5.88e-07 $l=3.2e-07 $layer=LI1_cond $X=6.875 $Y=1.625
+ $X2=6.555 $Y2=1.625
r149 50 73 2.05793 $w=4.18e-07 $l=7.5e-08 $layer=LI1_cond $X=6.48 $Y=1.625
+ $X2=6.555 $Y2=1.625
r150 50 68 7.27137 $w=4.18e-07 $l=2.65e-07 $layer=LI1_cond $X=6.48 $Y=1.625
+ $X2=6.215 $Y2=1.625
r151 49 68 5.89941 $w=4.18e-07 $l=2.15e-07 $layer=LI1_cond $X=6 $Y=1.625
+ $X2=6.215 $Y2=1.625
r152 49 63 12.7592 $w=4.18e-07 $l=4.65e-07 $layer=LI1_cond $X=6 $Y=1.625
+ $X2=5.535 $Y2=1.625
r153 48 63 0.411587 $w=4.18e-07 $l=1.5e-08 $layer=LI1_cond $X=5.52 $Y=1.625
+ $X2=5.535 $Y2=1.625
r154 47 48 13.1708 $w=4.18e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.625
+ $X2=5.52 $Y2=1.625
r155 46 47 13.1708 $w=4.18e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.625
+ $X2=5.04 $Y2=1.625
r156 43 45 17.7097 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=9.012 $Y=1.5
+ $X2=9.012 $Y2=1.86
r157 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.075
+ $Y=1.5 $X2=9.075 $Y2=1.5
r158 40 45 2.94836 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=8.855 $Y=1.86
+ $X2=9.012 $Y2=1.86
r159 40 96 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=8.855 $Y=1.86
+ $X2=7.045 $Y2=1.86
r160 36 44 38.924 $w=3.61e-07 $l=1.88348e-07 $layer=POLY_cond $X=9.075 $Y=1.665
+ $X2=9.025 $Y2=1.5
r161 36 38 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=9.075 $Y=1.665
+ $X2=9.075 $Y2=2.465
r162 33 44 58.9517 $w=3.61e-07 $l=3.78583e-07 $layer=POLY_cond $X=8.885 $Y=1.185
+ $X2=9.025 $Y2=1.5
r163 33 35 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.885 $Y=1.185
+ $X2=8.885 $Y2=0.655
r164 29 75 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.745 $Y=1.675
+ $X2=6.745 $Y2=1.51
r165 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.745 $Y=1.675
+ $X2=6.745 $Y2=2.465
r166 25 74 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.345
+ $X2=6.735 $Y2=1.51
r167 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.735 $Y=1.345
+ $X2=6.735 $Y2=0.655
r168 21 70 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.345
+ $X2=6.305 $Y2=1.51
r169 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.305 $Y=1.345
+ $X2=6.305 $Y2=0.655
r170 17 69 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.295 $Y=1.675
+ $X2=6.295 $Y2=1.51
r171 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.295 $Y=1.675
+ $X2=6.295 $Y2=2.465
r172 13 65 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.875 $Y=1.345
+ $X2=5.875 $Y2=1.51
r173 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.875 $Y=1.345
+ $X2=5.875 $Y2=0.655
r174 9 64 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.865 $Y=1.675
+ $X2=5.865 $Y2=1.51
r175 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.865 $Y=1.675
+ $X2=5.865 $Y2=2.465
r176 5 60 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.445 $Y=1.345
+ $X2=5.445 $Y2=1.51
r177 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.445 $Y=1.345
+ $X2=5.445 $Y2=0.655
r178 1 59 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.435 $Y=1.675
+ $X2=5.435 $Y2=1.51
r179 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.435 $Y=1.675
+ $X2=5.435 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%A_1418_21# 1 2 9 11 13 16 18 20 23 25 27 30
+ 32 34 35 44 45 46 49 51 53 60 62 71
c109 35 0 1.35208e-19 $X=8.505 $Y=1.51
c110 30 0 2.6512e-20 $X=8.455 $Y=0.655
r111 68 69 22.7611 $w=3.6e-07 $l=1.7e-07 $layer=POLY_cond $X=8.025 $Y=1.535
+ $X2=8.195 $Y2=1.535
r112 67 68 56.2333 $w=3.6e-07 $l=4.2e-07 $layer=POLY_cond $X=7.605 $Y=1.535
+ $X2=8.025 $Y2=1.535
r113 66 67 1.33889 $w=3.6e-07 $l=1e-08 $layer=POLY_cond $X=7.595 $Y=1.535
+ $X2=7.605 $Y2=1.535
r114 63 64 1.33889 $w=3.6e-07 $l=1e-08 $layer=POLY_cond $X=7.165 $Y=1.535
+ $X2=7.175 $Y2=1.535
r115 59 60 19.7172 $w=1.78e-07 $l=3.2e-07 $layer=LI1_cond $X=9.105 $Y=1.075
+ $X2=9.425 $Y2=1.075
r116 57 60 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.425 $Y=1.165
+ $X2=9.425 $Y2=1.075
r117 57 62 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.425 $Y=1.165
+ $X2=9.425 $Y2=1.845
r118 53 55 32.9269 $w=3.13e-07 $l=9e-07 $layer=LI1_cond $X=9.352 $Y=2.01
+ $X2=9.352 $Y2=2.91
r119 51 62 8.16989 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=9.352 $Y=2.002
+ $X2=9.352 $Y2=1.845
r120 51 53 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=9.352 $Y=2.002
+ $X2=9.352 $Y2=2.01
r121 47 59 0.0633028 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=9.105 $Y=0.985
+ $X2=9.105 $Y2=1.075
r122 47 49 31.3318 $w=1.98e-07 $l=5.65e-07 $layer=LI1_cond $X=9.105 $Y=0.985
+ $X2=9.105 $Y2=0.42
r123 45 59 6.16162 $w=1.78e-07 $l=1e-07 $layer=LI1_cond $X=9.005 $Y=1.075
+ $X2=9.105 $Y2=1.075
r124 45 46 20.3333 $w=1.78e-07 $l=3.3e-07 $layer=LI1_cond $X=9.005 $Y=1.075
+ $X2=8.675 $Y2=1.075
r125 43 46 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=8.59 $Y=1.165
+ $X2=8.675 $Y2=1.075
r126 43 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.59 $Y=1.165
+ $X2=8.59 $Y2=1.415
r127 42 71 6.025 $w=3.6e-07 $l=4.5e-08 $layer=POLY_cond $X=8.41 $Y=1.535
+ $X2=8.455 $Y2=1.535
r128 42 69 28.7861 $w=3.6e-07 $l=2.15e-07 $layer=POLY_cond $X=8.41 $Y=1.535
+ $X2=8.195 $Y2=1.535
r129 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.41
+ $Y=1.51 $X2=8.41 $Y2=1.51
r130 38 66 27.4472 $w=3.6e-07 $l=2.05e-07 $layer=POLY_cond $X=7.39 $Y=1.535
+ $X2=7.595 $Y2=1.535
r131 38 64 28.7861 $w=3.6e-07 $l=2.15e-07 $layer=POLY_cond $X=7.39 $Y=1.535
+ $X2=7.175 $Y2=1.535
r132 37 41 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=7.39 $Y=1.51
+ $X2=8.41 $Y2=1.51
r133 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.39
+ $Y=1.51 $X2=7.39 $Y2=1.51
r134 35 44 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.505 $Y=1.51
+ $X2=8.59 $Y2=1.415
r135 35 41 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=8.505 $Y=1.51
+ $X2=8.41 $Y2=1.51
r136 32 71 22.7611 $w=3.6e-07 $l=2.61534e-07 $layer=POLY_cond $X=8.625 $Y=1.725
+ $X2=8.455 $Y2=1.535
r137 32 34 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.625 $Y=1.725
+ $X2=8.625 $Y2=2.465
r138 28 71 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.455 $Y=1.345
+ $X2=8.455 $Y2=1.535
r139 28 30 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.455 $Y=1.345
+ $X2=8.455 $Y2=0.655
r140 25 69 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.195 $Y=1.725
+ $X2=8.195 $Y2=1.535
r141 25 27 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.195 $Y=1.725
+ $X2=8.195 $Y2=2.465
r142 21 68 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.025 $Y=1.345
+ $X2=8.025 $Y2=1.535
r143 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.025 $Y=1.345
+ $X2=8.025 $Y2=0.655
r144 18 67 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.605 $Y=1.725
+ $X2=7.605 $Y2=1.535
r145 18 20 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.605 $Y=1.725
+ $X2=7.605 $Y2=2.465
r146 14 66 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.595 $Y=1.345
+ $X2=7.595 $Y2=1.535
r147 14 16 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.595 $Y=1.345
+ $X2=7.595 $Y2=0.655
r148 11 64 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.175 $Y=1.725
+ $X2=7.175 $Y2=1.535
r149 11 13 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.175 $Y=1.725
+ $X2=7.175 $Y2=2.465
r150 7 63 23.3057 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.165 $Y=1.345
+ $X2=7.165 $Y2=1.535
r151 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.165 $Y=1.345
+ $X2=7.165 $Y2=0.655
r152 2 55 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.15
+ $Y=1.835 $X2=9.29 $Y2=2.91
r153 2 53 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=9.15
+ $Y=1.835 $X2=9.29 $Y2=2.01
r154 1 49 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.96
+ $Y=0.235 $X2=9.1 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 37 39 40 41 45
+ 53 55 59 60 64 70 73 76
c109 53 0 3.64334e-20 $X=1.895 $Y=1.105
c110 39 0 4.56457e-20 $X=1.035 $Y=1.16
r111 78 79 1.28049 $w=3.58e-07 $l=4e-08 $layer=LI1_cond $X=2.075 $Y=1.065
+ $X2=2.075 $Y2=1.105
r112 76 78 0.160062 $w=3.58e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=1.06
+ $X2=2.075 $Y2=1.065
r113 73 79 6.08234 $w=3.58e-07 $l=1.9e-07 $layer=LI1_cond $X=2.075 $Y=1.295
+ $X2=2.075 $Y2=1.105
r114 66 67 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.2 $Y=1.105
+ $X2=1.2 $Y2=1.16
r115 64 66 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.2 $Y=0.72
+ $X2=1.2 $Y2=1.105
r116 59 72 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.18 $Y=1.165 $X2=4.18
+ $Y2=1.065
r117 59 60 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.18 $Y=1.165
+ $X2=4.18 $Y2=1.93
r118 56 78 4.17751 $w=2e-07 $l=1.8e-07 $layer=LI1_cond $X=2.255 $Y=1.065
+ $X2=2.075 $Y2=1.065
r119 56 58 45.75 $w=1.98e-07 $l=8.25e-07 $layer=LI1_cond $X=2.255 $Y=1.065
+ $X2=3.08 $Y2=1.065
r120 55 72 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.095 $Y=1.065
+ $X2=4.18 $Y2=1.065
r121 55 58 56.2864 $w=1.98e-07 $l=1.015e-06 $layer=LI1_cond $X=4.095 $Y=1.065
+ $X2=3.08 $Y2=1.065
r122 54 66 1.70047 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=1.105
+ $X2=1.2 $Y2=1.105
r123 53 79 2.2115 $w=2.8e-07 $l=1.8e-07 $layer=LI1_cond $X=1.895 $Y=1.105
+ $X2=2.075 $Y2=1.105
r124 53 54 21.8141 $w=2.78e-07 $l=5.3e-07 $layer=LI1_cond $X=1.895 $Y=1.105
+ $X2=1.365 $Y2=1.105
r125 50 52 52.9899 $w=1.78e-07 $l=8.6e-07 $layer=LI1_cond $X=2.92 $Y=2.02
+ $X2=3.78 $Y2=2.02
r126 48 50 52.9899 $w=1.78e-07 $l=8.6e-07 $layer=LI1_cond $X=2.06 $Y=2.02
+ $X2=2.92 $Y2=2.02
r127 46 70 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.02
+ $X2=1.2 $Y2=2.02
r128 46 48 47.7525 $w=1.78e-07 $l=7.75e-07 $layer=LI1_cond $X=1.285 $Y=2.02
+ $X2=2.06 $Y2=2.02
r129 45 60 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.095 $Y=2.02
+ $X2=4.18 $Y2=1.93
r130 45 52 19.4091 $w=1.78e-07 $l=3.15e-07 $layer=LI1_cond $X=4.095 $Y=2.02
+ $X2=3.78 $Y2=2.02
r131 42 62 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.425 $Y=2.015
+ $X2=0.33 $Y2=2.015
r132 41 70 5.04255 $w=1.75e-07 $l=8.74643e-08 $layer=LI1_cond $X=1.115 $Y=2.015
+ $X2=1.2 $Y2=2.02
r133 41 42 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.115 $Y=2.015
+ $X2=0.425 $Y2=2.015
r134 39 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=1.2 $Y2=1.16
r135 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.16
+ $X2=0.345 $Y2=1.16
r136 35 62 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.33 $Y=2.1 $X2=0.33
+ $Y2=2.015
r137 35 37 39.4019 $w=1.88e-07 $l=6.75e-07 $layer=LI1_cond $X=0.33 $Y=2.1
+ $X2=0.33 $Y2=2.775
r138 31 40 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.25 $Y=1.075
+ $X2=0.345 $Y2=1.16
r139 31 33 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=0.25 $Y=1.075
+ $X2=0.25 $Y2=0.49
r140 10 52 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=3.64
+ $Y=1.835 $X2=3.78 $Y2=2.015
r141 9 50 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.835 $X2=2.92 $Y2=2.015
r142 8 48 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=2.015
r143 7 70 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=1.835 $X2=1.2 $Y2=2.095
r144 6 62 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.095
r145 6 37 400 $w=1.7e-07 $l=1.00055e-06 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.775
r146 5 72 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=3.96
+ $Y=0.345 $X2=4.1 $Y2=1.06
r147 4 58 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.345 $X2=3.08 $Y2=1.06
r148 3 76 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.345 $X2=2.06 $Y2=1.06
r149 2 64 91 $w=1.7e-07 $l=4.72361e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.345 $X2=1.2 $Y2=0.72
r150 1 33 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.345 $X2=0.26 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%A_126_367# 1 2 3 4 15 17 18 19 27 31 32
c47 27 0 3.05715e-20 $X=6.51 $Y=2.17
r48 31 32 8.3011 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.445 $Y=2.232
+ $X2=4.615 $Y2=2.232
r49 25 27 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.65 $Y=2.17
+ $X2=6.51 $Y2=2.17
r50 25 32 36.1448 $w=3.28e-07 $l=1.035e-06 $layer=LI1_cond $X=5.65 $Y=2.17
+ $X2=4.615 $Y2=2.17
r51 22 30 3.69874 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=1.735 $Y=2.37
+ $X2=1.63 $Y2=2.37
r52 22 31 166.98 $w=1.78e-07 $l=2.71e-06 $layer=LI1_cond $X=1.735 $Y=2.37
+ $X2=4.445 $Y2=2.37
r53 19 30 3.17035 $w=2.1e-07 $l=9e-08 $layer=LI1_cond $X=1.63 $Y=2.46 $X2=1.63
+ $Y2=2.37
r54 19 20 16.9004 $w=2.08e-07 $l=3.2e-07 $layer=LI1_cond $X=1.63 $Y=2.46
+ $X2=1.63 $Y2=2.78
r55 17 20 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.525 $Y=2.865
+ $X2=1.63 $Y2=2.78
r56 17 18 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.525 $Y=2.865
+ $X2=0.875 $Y2=2.865
r57 13 18 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.77 $Y=2.78
+ $X2=0.875 $Y2=2.865
r58 13 15 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=0.77 $Y=2.78
+ $X2=0.77 $Y2=2.445
r59 4 27 600 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=6.37
+ $Y=1.835 $X2=6.51 $Y2=2.17
r60 3 25 600 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=5.51
+ $Y=1.835 $X2=5.65 $Y2=2.17
r61 2 30 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=1.49
+ $Y=1.835 $X2=1.63 $Y2=2.445
r62 1 15 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=2.445
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%A_470_367# 1 2 3 4 13 17 23 25 27 29 33 34
+ 40 42
r70 41 42 9.2556 $w=5.58e-07 $l=1.35e-07 $layer=LI1_cond $X=7.43 $Y=2.395
+ $X2=7.565 $Y2=2.395
r71 39 41 0.854342 $w=5.58e-07 $l=4e-08 $layer=LI1_cond $X=7.39 $Y=2.395
+ $X2=7.43 $Y2=2.395
r72 39 40 17.2651 $w=5.58e-07 $l=5.1e-07 $layer=LI1_cond $X=7.39 $Y=2.395
+ $X2=6.88 $Y2=2.395
r73 34 36 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.88 $Y=2.59
+ $X2=4.88 $Y2=2.715
r74 32 33 7.30739 $w=4.43e-07 $l=1.05e-07 $layer=LI1_cond $X=3.35 $Y=2.852
+ $X2=3.455 $Y2=2.852
r75 27 44 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=2.285
+ $X2=8.405 $Y2=2.2
r76 27 29 22.8794 $w=3.38e-07 $l=6.75e-07 $layer=LI1_cond $X=8.405 $Y=2.285
+ $X2=8.405 $Y2=2.96
r77 25 44 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.235 $Y=2.2 $X2=8.405
+ $Y2=2.2
r78 25 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.235 $Y=2.2
+ $X2=7.565 $Y2=2.2
r79 21 41 5.0181 $w=2.7e-07 $l=2.8e-07 $layer=LI1_cond $X=7.43 $Y=2.675 $X2=7.43
+ $Y2=2.395
r80 21 23 9.60369 $w=2.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.43 $Y=2.675
+ $X2=7.43 $Y2=2.9
r81 20 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.965 $Y=2.59
+ $X2=4.88 $Y2=2.59
r82 20 40 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=4.965 $Y=2.59
+ $X2=6.88 $Y2=2.59
r83 17 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=2.715
+ $X2=4.88 $Y2=2.715
r84 17 33 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=4.795 $Y=2.715
+ $X2=3.455 $Y2=2.715
r85 13 32 3.03002 $w=4.43e-07 $l=1.17e-07 $layer=LI1_cond $X=3.233 $Y=2.852
+ $X2=3.35 $Y2=2.852
r86 13 15 19.2419 $w=4.43e-07 $l=7.43e-07 $layer=LI1_cond $X=3.233 $Y=2.852
+ $X2=2.49 $Y2=2.852
r87 4 44 400 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=1.835 $X2=8.41 $Y2=2.28
r88 4 29 400 $w=1.7e-07 $l=1.19295e-06 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=1.835 $X2=8.41 $Y2=2.96
r89 3 39 300 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=2 $X=7.25
+ $Y=1.835 $X2=7.39 $Y2=2.2
r90 3 23 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.835 $X2=7.39 $Y2=2.9
r91 2 32 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=1.835 $X2=3.35 $Y2=2.795
r92 1 15 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.835 $X2=2.49 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%VPWR 1 2 3 4 5 18 22 26 30 34 36 44 49 54 59
+ 66 67 70 77 80 83 86
c120 70 0 3.05715e-20 $X=5.105 $Y=3.065
r121 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r122 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r123 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r125 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r126 70 73 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=5.105 $Y=3.065
+ $X2=5.105 $Y2=3.33
r127 67 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r128 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r129 64 86 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=8.885 $Y2=3.33
r130 64 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=9.36 $Y2=3.33
r131 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r132 63 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r133 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r134 60 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.065 $Y=3.33
+ $X2=7.9 $Y2=3.33
r135 60 62 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.065 $Y=3.33
+ $X2=8.4 $Y2=3.33
r136 59 86 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.745 $Y=3.33
+ $X2=8.885 $Y2=3.33
r137 59 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.745 $Y=3.33
+ $X2=8.4 $Y2=3.33
r138 58 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r139 58 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r140 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r141 55 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=3.33
+ $X2=6.96 $Y2=3.33
r142 55 57 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.125 $Y=3.33
+ $X2=7.44 $Y2=3.33
r143 54 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.735 $Y=3.33
+ $X2=7.9 $Y2=3.33
r144 54 57 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.735 $Y=3.33
+ $X2=7.44 $Y2=3.33
r145 53 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r146 53 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r147 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r148 50 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.245 $Y=3.33
+ $X2=6.08 $Y2=3.33
r149 50 52 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.245 $Y=3.33
+ $X2=6.48 $Y2=3.33
r150 49 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=6.96 $Y2=3.33
r151 49 52 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=6.48 $Y2=3.33
r152 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r153 48 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r154 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r155 45 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.105 $Y2=3.33
r156 45 47 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.52 $Y2=3.33
r157 44 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.915 $Y=3.33
+ $X2=6.08 $Y2=3.33
r158 44 47 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.915 $Y=3.33
+ $X2=5.52 $Y2=3.33
r159 42 43 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r160 39 43 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r161 38 42 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r162 38 39 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r163 36 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.94 $Y=3.33
+ $X2=5.105 $Y2=3.33
r164 36 42 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.94 $Y=3.33
+ $X2=4.56 $Y2=3.33
r165 34 74 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r166 34 43 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r167 30 33 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=8.885 $Y=2.29
+ $X2=8.885 $Y2=2.97
r168 28 86 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=3.245
+ $X2=8.885 $Y2=3.33
r169 28 33 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=8.885 $Y=3.245
+ $X2=8.885 $Y2=2.97
r170 24 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=3.245 $X2=7.9
+ $Y2=3.33
r171 24 26 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=7.9 $Y=3.245
+ $X2=7.9 $Y2=2.54
r172 20 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.96 $Y=3.245
+ $X2=6.96 $Y2=3.33
r173 20 22 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=6.96 $Y=3.245
+ $X2=6.96 $Y2=2.945
r174 16 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.08 $Y=3.245
+ $X2=6.08 $Y2=3.33
r175 16 18 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=6.08 $Y=3.245
+ $X2=6.08 $Y2=2.96
r176 5 33 400 $w=1.7e-07 $l=1.21236e-06 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.835 $X2=8.86 $Y2=2.97
r177 5 30 400 $w=1.7e-07 $l=5.28985e-07 $layer=licon1_PDIFF $count=1 $X=8.7
+ $Y=1.835 $X2=8.86 $Y2=2.29
r178 4 26 300 $w=1.7e-07 $l=8.07543e-07 $layer=licon1_PDIFF $count=2 $X=7.68
+ $Y=1.835 $X2=7.9 $Y2=2.54
r179 3 22 600 $w=1.7e-07 $l=1.17792e-06 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.835 $X2=6.96 $Y2=2.945
r180 2 18 600 $w=1.7e-07 $l=1.19295e-06 $layer=licon1_PDIFF $count=1 $X=5.94
+ $Y=1.835 $X2=6.08 $Y2=2.96
r181 1 70 600 $w=1.7e-07 $l=1.30048e-06 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=1.835 $X2=5.105 $Y2=3.065
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%A_110_69# 1 2 3 4 15 17 18 20 21 24 25 26 29
+ 31 35 39
r90 33 35 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=8.24 $Y=1.075
+ $X2=8.24 $Y2=0.42
r91 32 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.475 $Y=1.16
+ $X2=7.38 $Y2=1.16
r92 31 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.145 $Y=1.16
+ $X2=8.24 $Y2=1.075
r93 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.145 $Y=1.16
+ $X2=7.475 $Y2=1.16
r94 27 39 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.38 $Y=1.075
+ $X2=7.38 $Y2=1.16
r95 27 29 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=7.38 $Y=1.075
+ $X2=7.38 $Y2=0.42
r96 25 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.285 $Y=1.16
+ $X2=7.38 $Y2=1.16
r97 25 26 174.193 $w=1.68e-07 $l=2.67e-06 $layer=LI1_cond $X=7.285 $Y=1.16
+ $X2=4.615 $Y2=1.16
r98 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.53 $Y=1.075
+ $X2=4.615 $Y2=1.16
r99 23 24 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.53 $Y=0.795
+ $X2=4.53 $Y2=1.075
r100 22 38 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.795 $Y=0.71
+ $X2=1.665 $Y2=0.71
r101 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.445 $Y=0.71
+ $X2=4.53 $Y2=0.795
r102 21 22 172.888 $w=1.68e-07 $l=2.65e-06 $layer=LI1_cond $X=4.445 $Y=0.71
+ $X2=1.795 $Y2=0.71
r103 20 38 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.625
+ $X2=1.665 $Y2=0.71
r104 19 20 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=1.665 $Y=0.455
+ $X2=1.665 $Y2=0.625
r105 17 19 6.96842 $w=2e-07 $l=1.72916e-07 $layer=LI1_cond $X=1.535 $Y=0.355
+ $X2=1.665 $Y2=0.455
r106 17 18 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=1.535 $Y=0.355
+ $X2=0.855 $Y2=0.355
r107 13 18 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=0.69 $Y=0.455
+ $X2=0.855 $Y2=0.355
r108 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.69 $Y=0.455
+ $X2=0.69 $Y2=0.47
r109 4 35 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.1
+ $Y=0.235 $X2=8.24 $Y2=0.42
r110 3 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.24
+ $Y=0.235 $X2=7.38 $Y2=0.42
r111 2 38 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.345 $X2=1.63 $Y2=0.63
r112 1 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.345 $X2=0.69 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%A_470_69# 1 2 3 4 13 20 21 22 25 27 31 33
r59 29 31 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=6.52 $Y=0.735
+ $X2=6.52 $Y2=0.42
r60 28 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=0.82
+ $X2=5.66 $Y2=0.82
r61 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.355 $Y=0.82
+ $X2=6.52 $Y2=0.735
r62 27 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.355 $Y=0.82
+ $X2=5.825 $Y2=0.82
r63 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.66 $Y=0.735
+ $X2=5.66 $Y2=0.82
r64 23 25 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.66 $Y=0.735
+ $X2=5.66 $Y2=0.45
r65 21 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=0.82
+ $X2=5.66 $Y2=0.82
r66 21 22 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.495 $Y=0.82
+ $X2=4.965 $Y2=0.82
r67 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.88 $Y=0.735
+ $X2=4.965 $Y2=0.82
r68 19 20 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.88 $Y=0.455
+ $X2=4.88 $Y2=0.735
r69 15 18 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=2.57 $Y=0.355
+ $X2=3.59 $Y2=0.355
r70 13 19 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.795 $Y=0.355
+ $X2=4.88 $Y2=0.455
r71 13 18 66.8227 $w=1.98e-07 $l=1.205e-06 $layer=LI1_cond $X=4.795 $Y=0.355
+ $X2=3.59 $Y2=0.355
r72 4 31 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.38
+ $Y=0.235 $X2=6.52 $Y2=0.42
r73 3 25 91 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=2 $X=5.52
+ $Y=0.235 $X2=5.66 $Y2=0.45
r74 2 18 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.345 $X2=3.59 $Y2=0.36
r75 1 15 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.345 $X2=2.57 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_4%VGND 1 2 3 4 5 18 20 24 28 32 36 38 39 41 42
+ 44 45 46 55 68 69 72 75
r109 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r110 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r111 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r112 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r113 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r114 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r115 63 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r116 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r117 60 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.115 $Y=0 $X2=6.985
+ $Y2=0
r118 60 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.115 $Y=0
+ $X2=7.44 $Y2=0
r119 59 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r120 59 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r121 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r122 56 72 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.185 $Y=0 $X2=6.09
+ $Y2=0
r123 56 58 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.185 $Y=0 $X2=6.48
+ $Y2=0
r124 55 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.855 $Y=0 $X2=6.985
+ $Y2=0
r125 55 58 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.855 $Y=0
+ $X2=6.48 $Y2=0
r126 54 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r127 53 54 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r128 49 53 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=5.04
+ $Y2=0
r129 49 50 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r130 46 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r131 46 50 1.27103 $w=4.9e-07 $l=4.56e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=0.24
+ $Y2=0
r132 44 65 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.505 $Y=0 $X2=8.4
+ $Y2=0
r133 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.505 $Y=0 $X2=8.67
+ $Y2=0
r134 43 68 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=8.835 $Y=0
+ $X2=9.36 $Y2=0
r135 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.835 $Y=0 $X2=8.67
+ $Y2=0
r136 41 62 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.645 $Y=0
+ $X2=7.44 $Y2=0
r137 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.645 $Y=0 $X2=7.81
+ $Y2=0
r138 40 65 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.975 $Y=0 $X2=8.4
+ $Y2=0
r139 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.975 $Y=0 $X2=7.81
+ $Y2=0
r140 38 53 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.135 $Y=0 $X2=5.04
+ $Y2=0
r141 38 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.135 $Y=0 $X2=5.23
+ $Y2=0
r142 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.67 $Y=0.085
+ $X2=8.67 $Y2=0
r143 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.67 $Y=0.085
+ $X2=8.67 $Y2=0.36
r144 30 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0
r145 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0.36
r146 26 75 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=0.085
+ $X2=6.985 $Y2=0
r147 26 28 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=6.985 $Y=0.085
+ $X2=6.985 $Y2=0.36
r148 22 72 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=0.085
+ $X2=6.09 $Y2=0
r149 22 24 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=6.09 $Y=0.085
+ $X2=6.09 $Y2=0.4
r150 21 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.325 $Y=0 $X2=5.23
+ $Y2=0
r151 20 72 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.995 $Y=0 $X2=6.09
+ $Y2=0
r152 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.995 $Y=0
+ $X2=5.325 $Y2=0
r153 16 39 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.23 $Y=0.085
+ $X2=5.23 $Y2=0
r154 16 18 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=5.23 $Y=0.085
+ $X2=5.23 $Y2=0.4
r155 5 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=8.53
+ $Y=0.235 $X2=8.67 $Y2=0.36
r156 4 32 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.67
+ $Y=0.235 $X2=7.81 $Y2=0.36
r157 3 28 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.81
+ $Y=0.235 $X2=6.95 $Y2=0.36
r158 2 24 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.95
+ $Y=0.235 $X2=6.09 $Y2=0.4
r159 1 18 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.235 $X2=5.23 $Y2=0.4
.ends

