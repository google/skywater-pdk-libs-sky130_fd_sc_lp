* File: sky130_fd_sc_lp__a22o_0.spice
* Created: Fri Aug 28 09:53:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22o_0.pex.spice"
.subckt sky130_fd_sc_lp__a22o_0  VNB VPB A2 A1 B1 B2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_85_155#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07875 AS=0.1281 PD=0.795 PS=1.45 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1003 A_235_47# N_A2_M1003_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.07875 PD=0.63 PS=0.795 NRD=14.28 NRS=27.132 M=1 R=2.8 SA=75000.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 N_A_85_155#_M1009_d N_A1_M1009_g A_235_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_415_47# N_B1_M1001_g N_A_85_155#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=31.428 M=1 R=2.8 SA=75001.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B2_M1004_g A_415_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_85_155#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.128 AS=0.1824 PD=1.04 PS=1.85 NRD=15.3857 NRS=6.1464 M=1 R=4.26667
+ SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1007 N_A_257_491#_M1007_d N_A2_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.128 PD=0.92 PS=1.04 NRD=0 NRS=21.5321 M=1 R=4.26667
+ SA=75000.8 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1000 N_A_85_155#_M1000_d N_B1_M1000_g N_A_257_491#_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1248 AS=0.0896 PD=1.03 PS=0.92 NRD=21.5321 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1006 N_A_257_491#_M1006_d N_B2_M1006_g N_A_85_155#_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1344 AS=0.1248 PD=1.06 PS=1.03 NRD=24.6053 NRS=12.2928 M=1
+ R=4.26667 SA=75001.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_257_491#_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1344 PD=1.81 PS=1.06 NRD=0 NRS=18.4589 M=1 R=4.26667
+ SA=75002.3 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a22o_0.pxi.spice"
*
.ends
*
*
