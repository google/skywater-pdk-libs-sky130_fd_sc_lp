* File: sky130_fd_sc_lp__clkdlybuf4s50_2.pxi.spice
* Created: Fri Aug 28 10:17:13 2020
* 
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%A N_A_M1005_g N_A_M1009_g A A N_A_c_66_n
+ PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%A
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%A_27_52# N_A_27_52#_M1005_s
+ N_A_27_52#_M1009_s N_A_27_52#_M1000_g N_A_27_52#_c_98_n N_A_27_52#_c_105_n
+ N_A_27_52#_c_106_n N_A_27_52#_c_99_n N_A_27_52#_c_100_n N_A_27_52#_c_107_n
+ N_A_27_52#_c_124_n N_A_27_52#_c_101_n N_A_27_52#_c_102_n N_A_27_52#_M1004_g
+ PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%A_27_52#
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%A_282_52# N_A_282_52#_M1004_d
+ N_A_282_52#_M1000_d N_A_282_52#_M1008_g N_A_282_52#_M1003_g
+ N_A_282_52#_c_162_n N_A_282_52#_c_163_n N_A_282_52#_c_168_n
+ N_A_282_52#_c_164_n N_A_282_52#_c_165_n N_A_282_52#_c_170_n
+ N_A_282_52#_c_166_n PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%A_282_52#
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%A_394_52# N_A_394_52#_M1008_s
+ N_A_394_52#_M1003_s N_A_394_52#_M1001_g N_A_394_52#_M1002_g
+ N_A_394_52#_M1006_g N_A_394_52#_M1007_g N_A_394_52#_c_236_n
+ N_A_394_52#_c_238_n N_A_394_52#_c_240_n N_A_394_52#_c_231_n
+ N_A_394_52#_c_232_n N_A_394_52#_c_226_n N_A_394_52#_c_227_n
+ N_A_394_52#_c_256_n N_A_394_52#_c_228_n
+ PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%A_394_52#
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%VPWR N_VPWR_M1009_d N_VPWR_M1003_d
+ N_VPWR_M1007_s N_VPWR_c_306_n N_VPWR_c_307_n N_VPWR_c_308_n N_VPWR_c_309_n
+ N_VPWR_c_310_n N_VPWR_c_311_n VPWR N_VPWR_c_312_n N_VPWR_c_313_n
+ N_VPWR_c_314_n N_VPWR_c_305_n VPWR PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%VPWR
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%X N_X_M1001_s N_X_M1002_d X X X X X X X
+ N_X_c_366_n N_X_c_355_n X PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%X
x_PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%VGND N_VGND_M1005_d N_VGND_M1008_d
+ N_VGND_M1006_d N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n
+ N_VGND_c_386_n N_VGND_c_387_n VGND N_VGND_c_388_n N_VGND_c_389_n
+ N_VGND_c_390_n N_VGND_c_391_n VGND PM_SKY130_FD_SC_LP__CLKDLYBUF4S50_2%VGND
cc_1 VNB N_A_M1005_g 0.0594522f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.47
cc_2 VNB A 0.0208018f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A_c_66_n 0.0326678f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_4 VNB N_A_27_52#_c_98_n 0.0205357f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_5 VNB N_A_27_52#_c_99_n 0.0050785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_52#_c_100_n 0.0115829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_52#_c_101_n 0.00219081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_52#_c_102_n 0.0108849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_52#_M1004_g 0.0660704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_282_52#_c_162_n 0.011676f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.335
cc_11 VNB N_A_282_52#_c_163_n 0.0150178f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.295
cc_12 VNB N_A_282_52#_c_164_n 0.0124045f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.665
cc_13 VNB N_A_282_52#_c_165_n 0.0396892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_282_52#_c_166_n 0.0419838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_394_52#_M1001_g 0.0450125f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_A_394_52#_M1002_g 0.00156615f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_17 VNB N_A_394_52#_M1006_g 0.0486632f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.665
cc_18 VNB N_A_394_52#_M1007_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.5
cc_19 VNB N_A_394_52#_c_226_n 0.0114279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_394_52#_c_227_n 4.4684e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_394_52#_c_228_n 0.0409209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_305_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB X 0.0402718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_382_n 0.00643581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_383_n 0.0035061f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.335
cc_26 VNB N_VGND_c_384_n 0.0132299f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.295
cc_27 VNB N_VGND_c_385_n 0.0223869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_386_n 0.0503863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_387_n 0.00532387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_388_n 0.0179296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_389_n 0.0223295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_390_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_391_n 0.258584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_A_M1009_g 0.0249089f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_35 VPB A 0.00827303f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_36 VPB N_A_c_66_n 0.00600603f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_37 VPB N_A_27_52#_M1000_g 0.0460129f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_38 VPB N_A_27_52#_c_105_n 0.00794922f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_39 VPB N_A_27_52#_c_106_n 0.0339238f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.665
cc_40 VPB N_A_27_52#_c_107_n 0.00375793f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.5
cc_41 VPB N_A_27_52#_c_101_n 0.00495942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_27_52#_c_102_n 0.0365622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_282_52#_M1003_g 0.0708555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_282_52#_c_168_n 0.0102217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_282_52#_c_165_n 0.011742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_282_52#_c_170_n 0.0138541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_394_52#_M1002_g 0.0208585f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_48 VPB N_A_394_52#_M1007_g 0.0236223f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.5
cc_49 VPB N_A_394_52#_c_231_n 0.00281615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_394_52#_c_232_n 0.0023233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_394_52#_c_227_n 0.00305928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_306_n 0.00284395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_307_n 0.002833f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.335
cc_54 VPB N_VPWR_c_308_n 0.013204f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_309_n 0.063294f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.665
cc_56 VPB N_VPWR_c_310_n 0.0477761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_311_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_312_n 0.0178675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_313_n 0.0217903f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_314_n 0.00516427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_305_n 0.0554067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB X 0.00701467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_X_c_355_n 0.00541438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 A N_A_27_52#_M1009_s 0.00237131f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_M1009_g N_A_27_52#_M1000_g 0.0249332f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_M1005_g N_A_27_52#_c_98_n 0.00946431f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_67 N_A_M1009_g N_A_27_52#_c_105_n 7.4234e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_68 A N_A_27_52#_c_105_n 0.0239868f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_c_66_n N_A_27_52#_c_105_n 7.87914e-19 $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_70 N_A_M1009_g N_A_27_52#_c_106_n 0.0106934f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_71 N_A_M1005_g N_A_27_52#_c_99_n 0.0106533f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_72 A N_A_27_52#_c_99_n 0.0106601f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A_M1005_g N_A_27_52#_c_100_n 0.00435937f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_74 A N_A_27_52#_c_100_n 0.0289379f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_c_66_n N_A_27_52#_c_100_n 0.00100334f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_76 N_A_M1009_g N_A_27_52#_c_107_n 0.0116182f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_77 A N_A_27_52#_c_107_n 0.00941865f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A_M1005_g N_A_27_52#_c_124_n 0.00261224f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_79 A N_A_27_52#_c_124_n 0.017308f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 A N_A_27_52#_c_101_n 0.0114464f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_c_66_n N_A_27_52#_c_101_n 0.00196087f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_82 A N_A_27_52#_c_102_n 3.24068e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A_c_66_n N_A_27_52#_c_102_n 0.0249332f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_84 N_A_M1005_g N_A_27_52#_M1004_g 0.0249332f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_85 A N_A_27_52#_M1004_g 0.00183643f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A_M1009_g N_VPWR_c_306_n 0.0068949f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_M1009_g N_VPWR_c_312_n 0.0054895f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_88 N_A_M1009_g N_VPWR_c_305_n 0.0110277f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_M1005_g N_VGND_c_382_n 0.00322874f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_90 N_A_M1005_g N_VGND_c_388_n 0.00547602f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_91 N_A_M1005_g N_VGND_c_391_n 0.00694827f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_92 N_A_27_52#_c_102_n N_A_282_52#_M1003_g 0.00287905f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_93 N_A_27_52#_c_124_n N_A_282_52#_c_163_n 0.0221959f $X=1.085 $Y=1.535 $X2=0
+ $Y2=0
cc_94 N_A_27_52#_c_101_n N_A_282_52#_c_163_n 0.00828764f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_95 N_A_27_52#_c_102_n N_A_282_52#_c_163_n 0.00414437f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_96 N_A_27_52#_M1004_g N_A_282_52#_c_163_n 0.00567511f $X=1.16 $Y=0.76 $X2=0
+ $Y2=0
cc_97 N_A_27_52#_M1000_g N_A_282_52#_c_168_n 0.00398828f $X=1.16 $Y=2.595 $X2=0
+ $Y2=0
cc_98 N_A_27_52#_c_101_n N_A_282_52#_c_168_n 0.0285056f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_99 N_A_27_52#_c_102_n N_A_282_52#_c_168_n 0.00361912f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_100 N_A_27_52#_c_102_n N_A_282_52#_c_165_n 0.00235448f $X=1.415 $Y=1.765
+ $X2=0 $Y2=0
cc_101 N_A_27_52#_M1004_g N_A_282_52#_c_165_n 0.00316492f $X=1.16 $Y=0.76 $X2=0
+ $Y2=0
cc_102 N_A_27_52#_M1000_g N_A_282_52#_c_170_n 0.0191551f $X=1.16 $Y=2.595 $X2=0
+ $Y2=0
cc_103 N_A_27_52#_c_101_n N_A_282_52#_c_170_n 0.00501863f $X=1.415 $Y=1.765
+ $X2=0 $Y2=0
cc_104 N_A_27_52#_c_102_n N_A_282_52#_c_170_n 0.00392394f $X=1.415 $Y=1.765
+ $X2=0 $Y2=0
cc_105 N_A_27_52#_c_107_n N_VPWR_M1009_d 0.0100392f $X=0.91 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_106 N_A_27_52#_M1000_g N_VPWR_c_306_n 0.0239003f $X=1.16 $Y=2.595 $X2=0 $Y2=0
cc_107 N_A_27_52#_c_107_n N_VPWR_c_306_n 0.0196228f $X=0.91 $Y=2.117 $X2=0 $Y2=0
cc_108 N_A_27_52#_c_101_n N_VPWR_c_306_n 0.0011162f $X=1.415 $Y=1.765 $X2=0
+ $Y2=0
cc_109 N_A_27_52#_M1000_g N_VPWR_c_310_n 0.0185301f $X=1.16 $Y=2.595 $X2=0 $Y2=0
cc_110 N_A_27_52#_c_106_n N_VPWR_c_312_n 0.0210467f $X=0.26 $Y=2.915 $X2=0 $Y2=0
cc_111 N_A_27_52#_M1009_s N_VPWR_c_305_n 0.00215158f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_112 N_A_27_52#_M1000_g N_VPWR_c_305_n 0.0309562f $X=1.16 $Y=2.595 $X2=0 $Y2=0
cc_113 N_A_27_52#_c_106_n N_VPWR_c_305_n 0.0125689f $X=0.26 $Y=2.915 $X2=0 $Y2=0
cc_114 N_A_27_52#_c_99_n N_VGND_M1005_d 0.00954115f $X=0.91 $Y=0.92 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_27_52#_c_99_n N_VGND_c_382_n 0.0207743f $X=0.91 $Y=0.92 $X2=0 $Y2=0
cc_116 N_A_27_52#_M1004_g N_VGND_c_382_n 0.00356758f $X=1.16 $Y=0.76 $X2=0 $Y2=0
cc_117 N_A_27_52#_M1004_g N_VGND_c_386_n 0.0186549f $X=1.16 $Y=0.76 $X2=0 $Y2=0
cc_118 N_A_27_52#_c_98_n N_VGND_c_388_n 0.0152237f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_119 N_A_27_52#_c_98_n N_VGND_c_391_n 0.0118277f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_120 N_A_27_52#_c_99_n N_VGND_c_391_n 0.01767f $X=0.91 $Y=0.92 $X2=0 $Y2=0
cc_121 N_A_27_52#_M1004_g N_VGND_c_391_n 0.0228755f $X=1.16 $Y=0.76 $X2=0 $Y2=0
cc_122 N_A_282_52#_c_166_n N_A_394_52#_M1001_g 0.024387f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_123 N_A_282_52#_M1003_g N_A_394_52#_M1002_g 0.024387f $X=2.485 $Y=2.595 $X2=0
+ $Y2=0
cc_124 N_A_282_52#_c_162_n N_A_394_52#_c_236_n 0.0577683f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_125 N_A_282_52#_c_166_n N_A_394_52#_c_236_n 0.0289245f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_126 N_A_282_52#_c_164_n N_A_394_52#_c_238_n 0.0305669f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_127 N_A_282_52#_c_166_n N_A_394_52#_c_238_n 0.0415495f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_128 N_A_282_52#_c_162_n N_A_394_52#_c_240_n 0.00858119f $X=1.55 $Y=0.435
+ $X2=0 $Y2=0
cc_129 N_A_282_52#_c_163_n N_A_394_52#_c_240_n 0.0121129f $X=1.755 $Y=1.655
+ $X2=0 $Y2=0
cc_130 N_A_282_52#_c_164_n N_A_394_52#_c_240_n 0.0177106f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_131 N_A_282_52#_c_165_n N_A_394_52#_c_240_n 0.00503939f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_132 N_A_282_52#_c_166_n N_A_394_52#_c_240_n 8.78991e-19 $X=2.375 $Y=1.37
+ $X2=0 $Y2=0
cc_133 N_A_282_52#_M1003_g N_A_394_52#_c_231_n 0.0162472f $X=2.485 $Y=2.595
+ $X2=0 $Y2=0
cc_134 N_A_282_52#_c_164_n N_A_394_52#_c_231_n 0.0101562f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_135 N_A_282_52#_M1003_g N_A_394_52#_c_232_n 0.0367464f $X=2.485 $Y=2.595
+ $X2=0 $Y2=0
cc_136 N_A_282_52#_c_168_n N_A_394_52#_c_232_n 0.00990869f $X=1.755 $Y=2.1 $X2=0
+ $Y2=0
cc_137 N_A_282_52#_c_164_n N_A_394_52#_c_232_n 0.0270017f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_138 N_A_282_52#_c_165_n N_A_394_52#_c_232_n 0.00459953f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_139 N_A_282_52#_c_170_n N_A_394_52#_c_232_n 0.0129926f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_140 N_A_282_52#_c_164_n N_A_394_52#_c_226_n 0.0207685f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_141 N_A_282_52#_c_166_n N_A_394_52#_c_226_n 0.00694396f $X=2.375 $Y=1.37
+ $X2=0 $Y2=0
cc_142 N_A_282_52#_c_164_n N_A_394_52#_c_227_n 0.00227963f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_143 N_A_282_52#_c_165_n N_A_394_52#_c_227_n 0.00442182f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_144 N_A_282_52#_M1003_g N_A_394_52#_c_256_n 0.0267868f $X=2.485 $Y=2.595
+ $X2=0 $Y2=0
cc_145 N_A_282_52#_c_170_n N_A_394_52#_c_256_n 0.0679402f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_146 N_A_282_52#_c_165_n N_A_394_52#_c_228_n 0.024387f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_147 N_A_282_52#_c_170_n N_VPWR_c_306_n 0.0233833f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_148 N_A_282_52#_M1003_g N_VPWR_c_307_n 0.0293591f $X=2.485 $Y=2.595 $X2=0
+ $Y2=0
cc_149 N_A_282_52#_M1003_g N_VPWR_c_310_n 0.0181551f $X=2.485 $Y=2.595 $X2=0
+ $Y2=0
cc_150 N_A_282_52#_c_170_n N_VPWR_c_310_n 0.0301474f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_151 N_A_282_52#_M1000_d N_VPWR_c_305_n 0.00215158f $X=1.41 $Y=2.095 $X2=0
+ $Y2=0
cc_152 N_A_282_52#_M1003_g N_VPWR_c_305_n 0.0303754f $X=2.485 $Y=2.595 $X2=0
+ $Y2=0
cc_153 N_A_282_52#_c_170_n N_VPWR_c_305_n 0.0175018f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_154 N_A_282_52#_M1003_g N_X_c_355_n 8.18301e-19 $X=2.485 $Y=2.595 $X2=0 $Y2=0
cc_155 N_A_282_52#_c_166_n N_VGND_c_383_n 0.0176721f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_156 N_A_282_52#_c_162_n N_VGND_c_386_n 0.0250858f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_157 N_A_282_52#_c_166_n N_VGND_c_386_n 0.0173758f $X=2.375 $Y=1.37 $X2=0
+ $Y2=0
cc_158 N_A_282_52#_c_162_n N_VGND_c_391_n 0.0155553f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_159 N_A_282_52#_c_166_n N_VGND_c_391_n 0.030234f $X=2.375 $Y=1.37 $X2=0 $Y2=0
cc_160 N_A_394_52#_c_231_n N_VPWR_M1003_d 0.00441005f $X=2.855 $Y=1.91 $X2=0
+ $Y2=0
cc_161 N_A_394_52#_M1002_g N_VPWR_c_307_n 0.007883f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_394_52#_c_231_n N_VPWR_c_307_n 0.0244283f $X=2.855 $Y=1.91 $X2=0
+ $Y2=0
cc_163 N_A_394_52#_c_232_n N_VPWR_c_307_n 0.00665185f $X=2.54 $Y=1.91 $X2=0
+ $Y2=0
cc_164 N_A_394_52#_c_226_n N_VPWR_c_307_n 5.09408e-19 $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_165 N_A_394_52#_c_256_n N_VPWR_c_307_n 0.0275329f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_166 N_A_394_52#_M1007_g N_VPWR_c_309_n 0.0125713f $X=3.6 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A_394_52#_c_256_n N_VPWR_c_310_n 0.0153681f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_168 N_A_394_52#_M1002_g N_VPWR_c_313_n 0.00564131f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_394_52#_M1007_g N_VPWR_c_313_n 0.00357668f $X=3.6 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_394_52#_M1003_s N_VPWR_c_305_n 0.00357787f $X=1.97 $Y=2.095 $X2=0
+ $Y2=0
cc_171 N_A_394_52#_M1002_g N_VPWR_c_305_n 0.010493f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A_394_52#_M1007_g N_VPWR_c_305_n 0.00653187f $X=3.6 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_394_52#_c_256_n N_VPWR_c_305_n 0.00945867f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_174 N_A_394_52#_M1001_g X 0.00799384f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A_394_52#_M1002_g X 0.0014189f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_394_52#_M1006_g X 0.021587f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_177 N_A_394_52#_M1007_g X 0.00596988f $X=3.6 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_394_52#_c_226_n X 0.0370853f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_179 N_A_394_52#_c_227_n X 0.00685385f $X=2.94 $Y=1.825 $X2=0 $Y2=0
cc_180 N_A_394_52#_c_228_n X 0.0142477f $X=3.6 $Y=1.46 $X2=0 $Y2=0
cc_181 N_A_394_52#_M1002_g X 0.0131738f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A_394_52#_M1007_g X 0.0322293f $X=3.6 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_394_52#_M1001_g N_X_c_366_n 0.00495371f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_184 N_A_394_52#_M1006_g N_X_c_366_n 0.0114044f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_185 N_A_394_52#_c_226_n N_X_c_366_n 0.00268957f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_186 N_A_394_52#_c_228_n N_X_c_366_n 0.00225933f $X=3.6 $Y=1.46 $X2=0 $Y2=0
cc_187 N_A_394_52#_M1002_g N_X_c_355_n 0.00339314f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_394_52#_M1007_g N_X_c_355_n 0.00698802f $X=3.6 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_394_52#_c_231_n N_X_c_355_n 0.0124458f $X=2.855 $Y=1.91 $X2=0 $Y2=0
cc_190 N_A_394_52#_c_226_n N_X_c_355_n 0.00881931f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_191 N_A_394_52#_c_227_n N_X_c_355_n 6.38382e-19 $X=2.94 $Y=1.825 $X2=0 $Y2=0
cc_192 N_A_394_52#_c_228_n N_X_c_355_n 0.00399236f $X=3.6 $Y=1.46 $X2=0 $Y2=0
cc_193 N_A_394_52#_c_238_n N_VGND_M1008_d 0.00205184f $X=2.855 $Y=1.097 $X2=0
+ $Y2=0
cc_194 N_A_394_52#_c_226_n N_VGND_M1008_d 0.00293623f $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_195 N_A_394_52#_M1001_g N_VGND_c_383_n 0.00514775f $X=3.17 $Y=0.47 $X2=0
+ $Y2=0
cc_196 N_A_394_52#_c_236_n N_VGND_c_383_n 0.0133572f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_197 N_A_394_52#_c_238_n N_VGND_c_383_n 0.00446569f $X=2.855 $Y=1.097 $X2=0
+ $Y2=0
cc_198 N_A_394_52#_c_226_n N_VGND_c_383_n 0.0103475f $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_199 N_A_394_52#_M1006_g N_VGND_c_385_n 0.00756872f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_200 N_A_394_52#_c_236_n N_VGND_c_386_n 0.0140261f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_201 N_A_394_52#_M1001_g N_VGND_c_389_n 0.0051159f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_202 N_A_394_52#_M1006_g N_VGND_c_389_n 0.00352007f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_203 N_A_394_52#_M1001_g N_VGND_c_391_n 0.00947564f $X=3.17 $Y=0.47 $X2=0
+ $Y2=0
cc_204 N_A_394_52#_M1006_g N_VGND_c_391_n 0.00613857f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_205 N_A_394_52#_c_236_n N_VGND_c_391_n 0.00945114f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_305_n N_X_M1002_d 0.00223559f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_207 N_VPWR_c_313_n X 0.0278606f $X=3.875 $Y=3.33 $X2=0 $Y2=0
cc_208 N_VPWR_c_305_n X 0.0174924f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_209 N_VPWR_c_309_n N_X_c_355_n 0.0493429f $X=3.96 $Y=1.98 $X2=0 $Y2=0
cc_210 N_X_c_366_n N_VGND_c_389_n 0.0207025f $X=3.61 $Y=0.475 $X2=0 $Y2=0
cc_211 N_X_c_366_n N_VGND_c_391_n 0.0174088f $X=3.61 $Y=0.475 $X2=0 $Y2=0
