* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__buf_16 A VGND VNB VPB VPWR X
X0 a_130_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 X a_130_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR A a_130_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND a_130_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 X a_130_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 X a_130_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 X a_130_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VGND a_130_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR a_130_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR A a_130_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND a_130_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VPWR A a_130_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 X a_130_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 X a_130_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VGND a_130_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR a_130_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 X a_130_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_130_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 X a_130_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VPWR a_130_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VGND A a_130_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_130_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 X a_130_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 X a_130_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VPWR a_130_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VPWR a_130_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 X a_130_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 X a_130_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 VGND A a_130_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 a_130_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 X a_130_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 VPWR a_130_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_130_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 VGND A a_130_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 X a_130_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 a_130_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 VPWR a_130_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 VGND a_130_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 X a_130_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 VGND a_130_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X40 VPWR a_130_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X41 X a_130_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X42 VGND a_130_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X43 VGND a_130_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
