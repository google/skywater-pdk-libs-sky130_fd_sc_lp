* File: sky130_fd_sc_lp__clkinv_1.pex.spice
* Created: Wed Sep  2 09:40:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKINV_1%A 3 7 9 11 13 14 15
r30 20 22 12.5087 $w=5.78e-07 $l=1.5e-07 $layer=POLY_cond $X=0.385 $Y=1.44
+ $X2=0.535 $Y2=1.44
r31 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.27 $X2=0.385 $Y2=1.27
r32 14 15 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r33 14 21 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.27
r34 13 21 10.7458 $w=3.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.29 $Y=0.925
+ $X2=0.29 $Y2=1.27
r35 9 22 35.8581 $w=5.78e-07 $l=4.3e-07 $layer=POLY_cond $X=0.965 $Y=1.44
+ $X2=0.535 $Y2=1.44
r36 9 11 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=0.965 $Y=1.6
+ $X2=0.965 $Y2=2.53
r37 5 9 35.1088 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.965 $Y=1.105
+ $X2=0.965 $Y2=1.44
r38 5 7 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.965 $Y=1.105
+ $X2=0.965 $Y2=0.56
r39 1 22 35.1088 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.535 $Y=1.775
+ $X2=0.535 $Y2=1.44
r40 1 3 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.535 $Y=1.775
+ $X2=0.535 $Y2=2.53
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_1%VPWR 1 2 7 9 11 13 15 17 27
r21 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r22 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 18 23 4.55946 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.237 $Y2=3.33
r24 18 20 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 17 26 4.50146 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=1.242 $Y2=3.33
r26 17 20 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r28 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 11 26 3.01621 $w=3e-07 $l=1.05924e-07 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.242 $Y2=3.33
r31 11 13 34.5733 $w=2.98e-07 $l=9e-07 $layer=LI1_cond $X=1.195 $Y=3.245
+ $X2=1.195 $Y2=2.345
r32 7 23 3.12265 $w=3.2e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.315 $Y=3.245
+ $X2=0.237 $Y2=3.33
r33 7 9 32.4125 $w=3.18e-07 $l=9e-07 $layer=LI1_cond $X=0.315 $Y=3.245 $X2=0.315
+ $Y2=2.345
r34 2 13 300 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.11 $X2=1.18 $Y2=2.345
r35 1 9 300 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=2 $X=0.195
+ $Y=2.11 $X2=0.32 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_1%Y 1 2 9 13 15 16 17
r24 17 32 9.57519 $w=6.38e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=1.665
+ $X2=0.965 $Y2=1.9
r25 16 17 4.76877 $w=8.08e-07 $l=2.85e-07 $layer=LI1_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.58
r26 16 22 2.52298 $w=6.38e-07 $l=1.35e-07 $layer=LI1_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.16
r27 15 22 4.39185 $w=6.38e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=0.925
+ $X2=0.965 $Y2=1.16
r28 15 28 7.75425 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=0.925
+ $X2=0.965 $Y2=0.84
r29 13 32 22.2973 $w=2.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.76 $Y=2.345
+ $X2=0.76 $Y2=1.9
r30 9 28 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=0.745 $Y=0.56
+ $X2=0.745 $Y2=0.84
r31 2 13 300 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=2.11 $X2=0.75 $Y2=2.345
r32 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.35 $X2=0.75 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_1%VGND 1 4 6 8 10 17
r12 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r13 10 16 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.227
+ $Y2=0
r14 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.72
+ $Y2=0
r15 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r16 8 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r17 4 16 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.227 $Y2=0
r18 4 6 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.56
r19 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.35 $X2=1.18 $Y2=0.56
.ends

