* File: sky130_fd_sc_lp__isobufsrc_2.pxi.spice
* Created: Fri Aug 28 10:41:49 2020
* 
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_2%A N_A_c_55_n N_A_M1001_g N_A_M1003_g A
+ N_A_c_58_n PM_SKY130_FD_SC_LP__ISOBUFSRC_2%A
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_2%SLEEP N_SLEEP_M1008_g N_SLEEP_M1000_g
+ N_SLEEP_M1009_g N_SLEEP_M1007_g N_SLEEP_c_82_n N_SLEEP_c_83_n N_SLEEP_c_84_n
+ SLEEP SLEEP N_SLEEP_c_86_n N_SLEEP_c_87_n N_SLEEP_c_88_n N_SLEEP_c_89_n
+ PM_SKY130_FD_SC_LP__ISOBUFSRC_2%SLEEP
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_2%A_40_131# N_A_40_131#_M1001_s
+ N_A_40_131#_M1003_s N_A_40_131#_M1002_g N_A_40_131#_M1004_g
+ N_A_40_131#_M1005_g N_A_40_131#_M1006_g N_A_40_131#_c_162_n
+ N_A_40_131#_c_167_n N_A_40_131#_c_168_n N_A_40_131#_c_169_n
+ N_A_40_131#_c_163_n PM_SKY130_FD_SC_LP__ISOBUFSRC_2%A_40_131#
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_2%VPWR N_VPWR_M1003_d N_VPWR_M1009_d
+ N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n N_VPWR_c_239_n VPWR
+ N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_235_n N_VPWR_c_243_n
+ PM_SKY130_FD_SC_LP__ISOBUFSRC_2%VPWR
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_2%A_283_367# N_A_283_367#_M1008_s
+ N_A_283_367#_M1005_d N_A_283_367#_c_274_n N_A_283_367#_c_269_n
+ N_A_283_367#_c_270_n N_A_283_367#_c_280_p
+ PM_SKY130_FD_SC_LP__ISOBUFSRC_2%A_283_367#
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_2%X N_X_M1000_s N_X_M1006_s N_X_M1002_s
+ N_X_c_288_n N_X_c_290_n N_X_c_291_n N_X_c_284_n N_X_c_335_p N_X_c_295_n
+ N_X_c_298_n N_X_c_299_n X X X X N_X_c_282_n N_X_c_285_n X
+ PM_SKY130_FD_SC_LP__ISOBUFSRC_2%X
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_2%VGND N_VGND_M1001_d N_VGND_M1004_d
+ N_VGND_M1007_d N_VGND_c_344_n N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n
+ N_VGND_c_348_n N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n
+ VGND N_VGND_c_353_n N_VGND_c_354_n N_VGND_c_355_n
+ PM_SKY130_FD_SC_LP__ISOBUFSRC_2%VGND
cc_1 VNB N_A_c_55_n 0.0241138f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.185
cc_2 VNB N_A_M1003_g 0.00876136f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=2.045
cc_3 VNB A 0.00391952f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_c_58_n 0.0435595f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.35
cc_5 VNB N_SLEEP_M1008_g 0.00801208f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.865
cc_6 VNB N_SLEEP_M1009_g 0.00818841f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.35
cc_7 VNB N_SLEEP_c_82_n 0.0154741f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.35
cc_8 VNB N_SLEEP_c_83_n 0.00286312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SLEEP_c_84_n 0.0350185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB SLEEP 0.0094207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_SLEEP_c_86_n 0.0340578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_SLEEP_c_87_n 0.0191036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SLEEP_c_88_n 0.0187962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_SLEEP_c_89_n 0.00242065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_40_131#_M1004_g 0.0217311f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_16 VNB N_A_40_131#_M1006_g 0.0226061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_40_131#_c_162_n 0.0459342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_40_131#_c_163_n 0.0364659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_235_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_282_n 0.0121728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB X 0.0392983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_344_n 0.00125389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_345_n 0.0195879f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_24 VNB N_VGND_c_346_n 3.20903e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_347_n 0.0156518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_348_n 0.0148035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_349_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_350_n 0.0110503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_351_n 0.011684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_352_n 0.0051069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_353_n 0.0207735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_354_n 0.200116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_355_n 0.0124031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_A_M1003_g 0.0290193f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=2.045
cc_35 VPB N_SLEEP_M1008_g 0.0219717f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.865
cc_36 VPB N_SLEEP_M1009_g 0.0231001f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.35
cc_37 VPB N_A_40_131#_M1002_g 0.0175377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_40_131#_M1005_g 0.0183585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_40_131#_c_162_n 0.00248628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_40_131#_c_167_n 0.0118207f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_40_131#_c_168_n 0.0440463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_40_131#_c_169_n 3.91648e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_40_131#_c_163_n 0.00481917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_236_n 0.0352776f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_237_n 0.0312174f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=1.35
cc_46 VPB N_VPWR_c_238_n 0.0338754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_239_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_240_n 0.0296693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_241_n 0.013281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_235_n 0.0861187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_243_n 0.00737949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_X_c_284_n 6.96303e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_X_c_285_n 0.0197554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB X 0.0215822f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 N_A_M1003_g N_SLEEP_M1008_g 0.0211152f $X=0.815 $Y=2.045 $X2=0 $Y2=0
cc_56 N_A_c_55_n SLEEP 0.00112309f $X=0.54 $Y=1.185 $X2=0 $Y2=0
cc_57 A SLEEP 0.0208664f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_58 N_A_c_58_n SLEEP 0.00158838f $X=0.815 $Y=1.35 $X2=0 $Y2=0
cc_59 A N_SLEEP_c_86_n 8.6118e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_60 N_A_c_58_n N_SLEEP_c_86_n 0.0215137f $X=0.815 $Y=1.35 $X2=0 $Y2=0
cc_61 N_A_c_55_n N_SLEEP_c_87_n 0.00315643f $X=0.54 $Y=1.185 $X2=0 $Y2=0
cc_62 N_A_c_55_n N_A_40_131#_c_162_n 0.0127423f $X=0.54 $Y=1.185 $X2=0 $Y2=0
cc_63 N_A_M1003_g N_A_40_131#_c_162_n 0.00528313f $X=0.815 $Y=2.045 $X2=0 $Y2=0
cc_64 A N_A_40_131#_c_162_n 0.0254262f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_M1003_g N_A_40_131#_c_167_n 0.016323f $X=0.815 $Y=2.045 $X2=0 $Y2=0
cc_66 A N_A_40_131#_c_168_n 0.0214592f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A_c_58_n N_A_40_131#_c_168_n 0.0073792f $X=0.815 $Y=1.35 $X2=0 $Y2=0
cc_68 N_A_M1003_g N_VPWR_c_236_n 0.0123802f $X=0.815 $Y=2.045 $X2=0 $Y2=0
cc_69 N_A_c_55_n N_VGND_c_344_n 0.00346565f $X=0.54 $Y=1.185 $X2=0 $Y2=0
cc_70 A N_VGND_c_344_n 0.0195665f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_c_58_n N_VGND_c_344_n 0.00212303f $X=0.815 $Y=1.35 $X2=0 $Y2=0
cc_72 N_A_c_55_n N_VGND_c_345_n 0.00141226f $X=0.54 $Y=1.185 $X2=0 $Y2=0
cc_73 N_A_c_55_n N_VGND_c_353_n 0.00399858f $X=0.54 $Y=1.185 $X2=0 $Y2=0
cc_74 N_A_c_55_n N_VGND_c_354_n 0.0046122f $X=0.54 $Y=1.185 $X2=0 $Y2=0
cc_75 N_SLEEP_c_82_n N_A_40_131#_M1004_g 0.00795531f $X=2.555 $Y=1.16 $X2=0
+ $Y2=0
cc_76 N_SLEEP_c_86_n N_A_40_131#_M1004_g 0.00760371f $X=1.265 $Y=1.35 $X2=0
+ $Y2=0
cc_77 N_SLEEP_c_87_n N_A_40_131#_M1004_g 0.0149247f $X=1.292 $Y=1.185 $X2=0
+ $Y2=0
cc_78 N_SLEEP_c_89_n N_A_40_131#_M1004_g 0.00576973f $X=1.775 $Y=1.255 $X2=0
+ $Y2=0
cc_79 N_SLEEP_M1009_g N_A_40_131#_M1005_g 0.0230507f $X=2.63 $Y=2.465 $X2=0
+ $Y2=0
cc_80 N_SLEEP_c_82_n N_A_40_131#_M1006_g 0.0112303f $X=2.555 $Y=1.16 $X2=0 $Y2=0
cc_81 N_SLEEP_c_83_n N_A_40_131#_M1006_g 0.00164432f $X=2.685 $Y=1.16 $X2=0
+ $Y2=0
cc_82 N_SLEEP_c_84_n N_A_40_131#_M1006_g 0.0179624f $X=2.72 $Y=1.35 $X2=0 $Y2=0
cc_83 N_SLEEP_c_88_n N_A_40_131#_M1006_g 0.014687f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_84 N_SLEEP_c_89_n N_A_40_131#_M1006_g 4.87471e-19 $X=1.775 $Y=1.255 $X2=0
+ $Y2=0
cc_85 SLEEP N_A_40_131#_c_162_n 0.00378826f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_86 N_SLEEP_M1008_g N_A_40_131#_c_167_n 0.0159487f $X=1.34 $Y=2.465 $X2=0
+ $Y2=0
cc_87 N_SLEEP_c_82_n N_A_40_131#_c_167_n 0.00591232f $X=2.555 $Y=1.16 $X2=0
+ $Y2=0
cc_88 SLEEP N_A_40_131#_c_167_n 0.0410064f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_89 N_SLEEP_c_86_n N_A_40_131#_c_167_n 0.00566317f $X=1.265 $Y=1.35 $X2=0
+ $Y2=0
cc_90 N_SLEEP_M1008_g N_A_40_131#_c_169_n 6.23496e-19 $X=1.34 $Y=2.465 $X2=0
+ $Y2=0
cc_91 N_SLEEP_c_82_n N_A_40_131#_c_169_n 0.0249391f $X=2.555 $Y=1.16 $X2=0 $Y2=0
cc_92 N_SLEEP_c_83_n N_A_40_131#_c_169_n 0.00494609f $X=2.685 $Y=1.16 $X2=0
+ $Y2=0
cc_93 N_SLEEP_c_84_n N_A_40_131#_c_169_n 0.0024751f $X=2.72 $Y=1.35 $X2=0 $Y2=0
cc_94 N_SLEEP_c_86_n N_A_40_131#_c_169_n 3.59524e-19 $X=1.265 $Y=1.35 $X2=0
+ $Y2=0
cc_95 N_SLEEP_c_89_n N_A_40_131#_c_169_n 0.00152366f $X=1.775 $Y=1.255 $X2=0
+ $Y2=0
cc_96 N_SLEEP_M1008_g N_A_40_131#_c_163_n 0.0301376f $X=1.34 $Y=2.465 $X2=0
+ $Y2=0
cc_97 N_SLEEP_c_82_n N_A_40_131#_c_163_n 0.00262536f $X=2.555 $Y=1.16 $X2=0
+ $Y2=0
cc_98 N_SLEEP_c_84_n N_A_40_131#_c_163_n 0.0230507f $X=2.72 $Y=1.35 $X2=0 $Y2=0
cc_99 N_SLEEP_c_86_n N_A_40_131#_c_163_n 0.0125098f $X=1.265 $Y=1.35 $X2=0 $Y2=0
cc_100 N_SLEEP_c_89_n N_A_40_131#_c_163_n 0.00783032f $X=1.775 $Y=1.255 $X2=0
+ $Y2=0
cc_101 N_SLEEP_M1008_g N_VPWR_c_236_n 0.00717778f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_102 N_SLEEP_M1009_g N_VPWR_c_237_n 0.0155522f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_103 N_SLEEP_M1008_g N_VPWR_c_238_n 0.00585385f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_104 N_SLEEP_M1009_g N_VPWR_c_238_n 0.00486043f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_105 N_SLEEP_M1008_g N_VPWR_c_235_n 0.0118611f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_106 N_SLEEP_M1009_g N_VPWR_c_235_n 0.0082726f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_107 N_SLEEP_c_83_n N_X_M1006_s 4.81672e-19 $X=2.685 $Y=1.16 $X2=0 $Y2=0
cc_108 SLEEP N_X_c_288_n 0.0192731f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_109 N_SLEEP_c_87_n N_X_c_288_n 0.00232771f $X=1.292 $Y=1.185 $X2=0 $Y2=0
cc_110 N_SLEEP_c_87_n N_X_c_290_n 0.00538866f $X=1.292 $Y=1.185 $X2=0 $Y2=0
cc_111 N_SLEEP_c_89_n N_X_c_291_n 0.0405405f $X=1.775 $Y=1.255 $X2=0 $Y2=0
cc_112 N_SLEEP_M1009_g N_X_c_284_n 0.0178351f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_113 N_SLEEP_c_83_n N_X_c_284_n 0.00703577f $X=2.685 $Y=1.16 $X2=0 $Y2=0
cc_114 N_SLEEP_c_84_n N_X_c_284_n 0.00227463f $X=2.72 $Y=1.35 $X2=0 $Y2=0
cc_115 N_SLEEP_c_83_n N_X_c_295_n 0.0157867f $X=2.685 $Y=1.16 $X2=0 $Y2=0
cc_116 N_SLEEP_c_84_n N_X_c_295_n 0.00261103f $X=2.72 $Y=1.35 $X2=0 $Y2=0
cc_117 N_SLEEP_c_88_n N_X_c_295_n 0.0117068f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_118 N_SLEEP_M1009_g N_X_c_298_n 8.60449e-19 $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_119 N_SLEEP_c_82_n N_X_c_299_n 0.0145842f $X=2.555 $Y=1.16 $X2=0 $Y2=0
cc_120 N_SLEEP_M1009_g X 0.0165174f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_121 N_SLEEP_c_83_n X 0.0343109f $X=2.685 $Y=1.16 $X2=0 $Y2=0
cc_122 N_SLEEP_c_84_n X 0.00814607f $X=2.72 $Y=1.35 $X2=0 $Y2=0
cc_123 N_SLEEP_c_88_n X 0.00645327f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_124 N_SLEEP_c_83_n N_VGND_M1007_d 7.00615e-19 $X=2.685 $Y=1.16 $X2=0 $Y2=0
cc_125 SLEEP N_VGND_c_344_n 0.0164013f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_126 N_SLEEP_c_86_n N_VGND_c_344_n 9.63447e-19 $X=1.265 $Y=1.35 $X2=0 $Y2=0
cc_127 N_SLEEP_c_87_n N_VGND_c_344_n 0.00220188f $X=1.292 $Y=1.185 $X2=0 $Y2=0
cc_128 N_SLEEP_c_87_n N_VGND_c_345_n 0.00330481f $X=1.292 $Y=1.185 $X2=0 $Y2=0
cc_129 N_SLEEP_c_87_n N_VGND_c_346_n 4.78045e-19 $X=1.292 $Y=1.185 $X2=0 $Y2=0
cc_130 N_SLEEP_c_88_n N_VGND_c_346_n 5.37623e-19 $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_131 N_SLEEP_c_88_n N_VGND_c_347_n 0.00873456f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_132 N_SLEEP_c_87_n N_VGND_c_348_n 0.0054895f $X=1.292 $Y=1.185 $X2=0 $Y2=0
cc_133 N_SLEEP_c_88_n N_VGND_c_351_n 0.00365202f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_134 N_SLEEP_c_87_n N_VGND_c_354_n 0.0110907f $X=1.292 $Y=1.185 $X2=0 $Y2=0
cc_135 N_SLEEP_c_88_n N_VGND_c_354_n 0.00434777f $X=2.72 $Y=1.185 $X2=0 $Y2=0
cc_136 N_A_40_131#_c_167_n N_VPWR_M1003_d 0.00279025f $X=1.945 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_40_131#_c_167_n N_VPWR_c_236_n 0.0230207f $X=1.945 $Y=1.77 $X2=0
+ $Y2=0
cc_138 N_A_40_131#_M1005_g N_VPWR_c_237_n 0.00109252f $X=2.2 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_40_131#_M1002_g N_VPWR_c_238_n 0.00357877f $X=1.77 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_40_131#_M1005_g N_VPWR_c_238_n 0.00357877f $X=2.2 $Y=2.465 $X2=0
+ $Y2=0
cc_141 N_A_40_131#_M1002_g N_VPWR_c_235_n 0.00537654f $X=1.77 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_40_131#_M1005_g N_VPWR_c_235_n 0.00537654f $X=2.2 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_40_131#_c_167_n N_A_283_367#_M1008_s 0.00176461f $X=1.945 $Y=1.77
+ $X2=-0.19 $Y2=-0.245
cc_144 N_A_40_131#_c_167_n N_A_283_367#_c_269_n 0.0135055f $X=1.945 $Y=1.77
+ $X2=0 $Y2=0
cc_145 N_A_40_131#_M1002_g N_A_283_367#_c_270_n 0.0117609f $X=1.77 $Y=2.465
+ $X2=0 $Y2=0
cc_146 N_A_40_131#_M1005_g N_A_283_367#_c_270_n 0.0117609f $X=2.2 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_40_131#_c_167_n N_X_M1002_s 5.03153e-19 $X=1.945 $Y=1.77 $X2=0 $Y2=0
cc_148 N_A_40_131#_c_169_n N_X_M1002_s 0.00137738f $X=2.11 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A_40_131#_M1004_g N_X_c_291_n 0.00990046f $X=1.815 $Y=0.655 $X2=0 $Y2=0
cc_150 N_A_40_131#_M1006_g N_X_c_291_n 0.00988678f $X=2.245 $Y=0.655 $X2=0 $Y2=0
cc_151 N_A_40_131#_M1005_g N_X_c_284_n 0.0110405f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_40_131#_c_169_n N_X_c_284_n 0.00907688f $X=2.11 $Y=1.51 $X2=0 $Y2=0
cc_153 N_A_40_131#_M1002_g N_X_c_298_n 0.00896657f $X=1.77 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_40_131#_M1005_g N_X_c_298_n 0.00900398f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_40_131#_c_167_n N_X_c_298_n 0.00536701f $X=1.945 $Y=1.77 $X2=0 $Y2=0
cc_156 N_A_40_131#_c_169_n N_X_c_298_n 0.012676f $X=2.11 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A_40_131#_c_163_n N_X_c_298_n 4.99587e-19 $X=2.2 $Y=1.505 $X2=0 $Y2=0
cc_158 N_A_40_131#_c_167_n N_VGND_c_344_n 3.11277e-19 $X=1.945 $Y=1.77 $X2=0
+ $Y2=0
cc_159 N_A_40_131#_M1004_g N_VGND_c_346_n 0.00772269f $X=1.815 $Y=0.655 $X2=0
+ $Y2=0
cc_160 N_A_40_131#_M1006_g N_VGND_c_346_n 0.00758038f $X=2.245 $Y=0.655 $X2=0
+ $Y2=0
cc_161 N_A_40_131#_M1006_g N_VGND_c_347_n 5.37623e-19 $X=2.245 $Y=0.655 $X2=0
+ $Y2=0
cc_162 N_A_40_131#_M1004_g N_VGND_c_348_n 0.00365202f $X=1.815 $Y=0.655 $X2=0
+ $Y2=0
cc_163 N_A_40_131#_M1006_g N_VGND_c_351_n 0.00365202f $X=2.245 $Y=0.655 $X2=0
+ $Y2=0
cc_164 N_A_40_131#_c_162_n N_VGND_c_353_n 0.00436993f $X=0.325 $Y=0.865 $X2=0
+ $Y2=0
cc_165 N_A_40_131#_M1004_g N_VGND_c_354_n 0.00434777f $X=1.815 $Y=0.655 $X2=0
+ $Y2=0
cc_166 N_A_40_131#_M1006_g N_VGND_c_354_n 0.00434777f $X=2.245 $Y=0.655 $X2=0
+ $Y2=0
cc_167 N_A_40_131#_c_162_n N_VGND_c_354_n 0.00775106f $X=0.325 $Y=0.865 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_235_n N_A_283_367#_M1008_s 0.00220345f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_169 N_VPWR_c_235_n N_A_283_367#_M1005_d 0.00376627f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_238_n N_A_283_367#_c_274_n 0.0139427f $X=2.68 $Y=3.33 $X2=0
+ $Y2=0
cc_171 N_VPWR_c_235_n N_A_283_367#_c_274_n 0.00894187f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_238_n N_A_283_367#_c_270_n 0.0487587f $X=2.68 $Y=3.33 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_235_n N_A_283_367#_c_270_n 0.0310969f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_235_n N_X_M1002_s 0.00225186f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_175 N_VPWR_M1009_d N_X_c_284_n 0.00814988f $X=2.705 $Y=1.835 $X2=0 $Y2=0
cc_176 N_VPWR_c_237_n N_X_c_284_n 0.0199378f $X=2.845 $Y=2.47 $X2=0 $Y2=0
cc_177 N_VPWR_c_237_n N_X_c_285_n 0.00220189f $X=2.845 $Y=2.47 $X2=0 $Y2=0
cc_178 N_A_283_367#_c_270_n N_X_M1002_s 0.00335193f $X=2.32 $Y=2.985 $X2=0 $Y2=0
cc_179 N_A_283_367#_M1005_d N_X_c_284_n 0.00809843f $X=2.275 $Y=1.835 $X2=0
+ $Y2=0
cc_180 N_A_283_367#_c_280_p N_X_c_284_n 0.0135534f $X=2.415 $Y=2.53 $X2=0 $Y2=0
cc_181 N_A_283_367#_c_270_n N_X_c_298_n 0.0152459f $X=2.32 $Y=2.985 $X2=0.295
+ $Y2=1.947
cc_182 N_X_c_291_n N_VGND_M1004_d 0.00335437f $X=2.365 $Y=0.82 $X2=0 $Y2=0
cc_183 N_X_c_295_n N_VGND_M1007_d 0.00707471f $X=2.985 $Y=0.82 $X2=0 $Y2=0
cc_184 N_X_c_282_n N_VGND_M1007_d 6.06399e-19 $X=3.13 $Y=0.905 $X2=0 $Y2=0
cc_185 X N_VGND_M1007_d 0.00243406f $X=3.12 $Y=0.925 $X2=0 $Y2=0
cc_186 N_X_c_288_n N_VGND_c_344_n 6.57844e-19 $X=1.565 $Y=0.735 $X2=0 $Y2=0
cc_187 N_X_c_291_n N_VGND_c_346_n 0.016459f $X=2.365 $Y=0.82 $X2=0 $Y2=0
cc_188 N_X_c_295_n N_VGND_c_347_n 0.0156459f $X=2.985 $Y=0.82 $X2=0 $Y2=0
cc_189 N_X_c_282_n N_VGND_c_347_n 0.00611061f $X=3.13 $Y=0.905 $X2=0 $Y2=0
cc_190 N_X_c_290_n N_VGND_c_348_n 0.0156443f $X=1.6 $Y=0.42 $X2=0 $Y2=0
cc_191 N_X_c_291_n N_VGND_c_348_n 0.00196209f $X=2.365 $Y=0.82 $X2=0 $Y2=0
cc_192 N_X_c_282_n N_VGND_c_350_n 0.00365955f $X=3.13 $Y=0.905 $X2=0 $Y2=0
cc_193 N_X_c_291_n N_VGND_c_351_n 0.00196209f $X=2.365 $Y=0.82 $X2=0 $Y2=0
cc_194 N_X_c_335_p N_VGND_c_351_n 0.0124139f $X=2.46 $Y=0.42 $X2=0 $Y2=0
cc_195 N_X_c_295_n N_VGND_c_351_n 0.00196209f $X=2.985 $Y=0.82 $X2=0 $Y2=0
cc_196 N_X_M1000_s N_VGND_c_354_n 0.00245017f $X=1.46 $Y=0.235 $X2=0 $Y2=0
cc_197 N_X_M1006_s N_VGND_c_354_n 0.00266476f $X=2.32 $Y=0.235 $X2=0 $Y2=0
cc_198 N_X_c_290_n N_VGND_c_354_n 0.00983564f $X=1.6 $Y=0.42 $X2=0 $Y2=0
cc_199 N_X_c_291_n N_VGND_c_354_n 0.00891615f $X=2.365 $Y=0.82 $X2=0 $Y2=0
cc_200 N_X_c_335_p N_VGND_c_354_n 0.00730033f $X=2.46 $Y=0.42 $X2=0 $Y2=0
cc_201 N_X_c_295_n N_VGND_c_354_n 0.00481455f $X=2.985 $Y=0.82 $X2=0 $Y2=0
cc_202 N_X_c_282_n N_VGND_c_354_n 0.00653835f $X=3.13 $Y=0.905 $X2=0 $Y2=0
