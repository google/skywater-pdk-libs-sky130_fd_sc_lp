* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand4_4 A B C D VGND VNB VPB VPWR Y
X0 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_454_65# B a_843_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_843_67# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 Y A a_843_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_454_65# B a_843_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VGND D a_27_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_27_65# D VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_27_65# C a_454_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_454_65# C a_27_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_843_67# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_843_67# B a_454_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 Y A a_843_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VGND D a_27_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_27_65# C a_454_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_27_65# D VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_454_65# C a_27_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_843_67# B a_454_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
