# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__or4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__or4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 0.775000 1.310000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 0.925000 1.920000 1.455000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 0.470000 0.815000 1.435000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.215000 1.405000 4.715000 1.760000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.450000 0.255000 3.695000 2.275000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.160000  0.280000 0.410000 1.625000 ;
      RECT 0.160000  1.625000 2.460000 1.795000 ;
      RECT 0.495000  1.795000 0.790000 2.390000 ;
      RECT 0.960000  2.045000 1.255000 3.245000 ;
      RECT 0.985000  0.085000 1.245000 0.605000 ;
      RECT 1.415000  0.265000 1.650000 0.585000 ;
      RECT 1.415000  0.585000 2.810000 0.595000 ;
      RECT 1.480000  0.595000 2.810000 0.755000 ;
      RECT 1.865000  0.085000 2.195000 0.415000 ;
      RECT 2.130000  0.925000 2.460000 1.625000 ;
      RECT 2.435000  0.280000 2.810000 0.585000 ;
      RECT 2.435000  1.995000 2.810000 2.275000 ;
      RECT 2.475000  2.445000 4.205000 2.615000 ;
      RECT 2.475000  2.615000 2.805000 3.075000 ;
      RECT 2.640000  0.755000 2.810000 1.185000 ;
      RECT 2.640000  1.185000 3.280000 1.515000 ;
      RECT 2.640000  1.515000 2.810000 1.995000 ;
      RECT 2.980000  0.085000 3.280000 1.015000 ;
      RECT 2.985000  2.785000 3.315000 3.245000 ;
      RECT 3.845000  2.785000 4.175000 3.245000 ;
      RECT 3.865000  0.085000 4.140000 0.895000 ;
      RECT 3.865000  1.065000 4.665000 1.235000 ;
      RECT 3.865000  1.235000 4.035000 1.930000 ;
      RECT 3.865000  1.930000 4.700000 2.260000 ;
      RECT 3.865000  2.260000 4.205000 2.445000 ;
      RECT 4.335000  0.700000 4.665000 1.065000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__or4bb_2
END LIBRARY
