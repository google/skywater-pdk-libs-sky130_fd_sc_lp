* File: sky130_fd_sc_lp__or3_1.spice
* Created: Wed Sep  2 10:30:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or3_1.pex.spice"
.subckt sky130_fd_sc_lp__or3_1  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_C_M1007_g N_A_47_47#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1323 AS=0.1113 PD=1.05 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1006 N_A_47_47#_M1006_d N_B_M1006_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1323 PD=0.7 PS=1.05 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_47_47#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0952 AS=0.0588 PD=0.823333 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_47_47#_M1001_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1904 PD=2.21 PS=1.64667 NRD=0 NRS=4.632 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 A_157_462# N_C_M1003_g N_A_47_47#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0609 AS=0.1113 PD=0.71 PS=1.37 NRD=42.1974 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1004 A_245_462# N_B_M1004_g A_157_462# VPB PHIGHVT L=0.15 W=0.42 AD=0.0651
+ AS=0.0609 PD=0.73 PS=0.71 NRD=46.886 NRS=42.1974 M=1 R=2.8 SA=75000.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_245_462# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.123375 AS=0.0651 PD=0.9525 PS=0.73 NRD=111.975 NRS=46.886 M=1 R=2.8
+ SA=75001.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_47_47#_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.370125 PD=3.05 PS=2.8575 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__or3_1.pxi.spice"
*
.ends
*
*
