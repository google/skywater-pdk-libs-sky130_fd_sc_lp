* File: sky130_fd_sc_lp__o21bai_0.spice
* Created: Fri Aug 28 11:06:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21bai_0.pex.spice"
.subckt sky130_fd_sc_lp__o21bai_0  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_B1_N_M1007_g N_A_39_51#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_320_47#_M1005_d N_A_39_51#_M1005_g N_Y_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_320_47#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_320_47#_M1003_d N_A1_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_B1_N_M1002_g N_A_39_51#_M1002_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0863377 AS=0.1113 PD=0.808302 PS=1.37 NRD=24.6053 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_A_39_51#_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.131562 PD=0.92 PS=1.2317 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75000.5 SB=75001 A=0.096 P=1.58 MULT=1
MM1004 A_406_473# N_A2_M1004_g N_Y_M1006_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0896 PD=0.88 PS=0.92 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75001 SB=75000.6
+ A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_406_473# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
c_71 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o21bai_0.pxi.spice"
*
.ends
*
*
