* File: sky130_fd_sc_lp__o21ba_lp.pxi.spice
* Created: Wed Sep  2 10:17:04 2020
* 
x_PM_SKY130_FD_SC_LP__O21BA_LP%A1 N_A1_M1001_g N_A1_M1004_g A1 A1 N_A1_c_82_n
+ PM_SKY130_FD_SC_LP__O21BA_LP%A1
x_PM_SKY130_FD_SC_LP__O21BA_LP%A2 N_A2_M1010_g N_A2_M1002_g N_A2_c_109_n
+ N_A2_c_110_n A2 A2 N_A2_c_112_n PM_SKY130_FD_SC_LP__O21BA_LP%A2
x_PM_SKY130_FD_SC_LP__O21BA_LP%A_317_29# N_A_317_29#_M1007_s N_A_317_29#_M1000_d
+ N_A_317_29#_M1005_g N_A_317_29#_M1008_g N_A_317_29#_c_150_n
+ N_A_317_29#_c_151_n N_A_317_29#_c_152_n N_A_317_29#_c_153_n
+ N_A_317_29#_c_154_n N_A_317_29#_c_155_n N_A_317_29#_c_156_n
+ N_A_317_29#_c_157_n N_A_317_29#_c_160_n PM_SKY130_FD_SC_LP__O21BA_LP%A_317_29#
x_PM_SKY130_FD_SC_LP__O21BA_LP%B1_N N_B1_N_c_222_n N_B1_N_M1000_g N_B1_N_c_223_n
+ N_B1_N_c_224_n N_B1_N_M1007_g N_B1_N_M1003_g N_B1_N_c_225_n N_B1_N_c_218_n
+ N_B1_N_c_219_n B1_N N_B1_N_c_221_n PM_SKY130_FD_SC_LP__O21BA_LP%B1_N
x_PM_SKY130_FD_SC_LP__O21BA_LP%A_253_389# N_A_253_389#_M1005_d
+ N_A_253_389#_M1010_d N_A_253_389#_M1011_g N_A_253_389#_M1006_g
+ N_A_253_389#_M1009_g N_A_253_389#_c_279_n N_A_253_389#_c_285_n
+ N_A_253_389#_c_280_n N_A_253_389#_c_281_n N_A_253_389#_c_287_n
+ N_A_253_389#_c_288_n N_A_253_389#_c_282_n N_A_253_389#_c_289_n
+ PM_SKY130_FD_SC_LP__O21BA_LP%A_253_389#
x_PM_SKY130_FD_SC_LP__O21BA_LP%VPWR N_VPWR_M1004_s N_VPWR_M1008_d N_VPWR_M1006_s
+ N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_371_n
+ N_VPWR_c_372_n VPWR N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_366_n
+ N_VPWR_c_376_n PM_SKY130_FD_SC_LP__O21BA_LP%VPWR
x_PM_SKY130_FD_SC_LP__O21BA_LP%X N_X_M1009_d N_X_M1006_d N_X_c_410_n X X X X X X
+ PM_SKY130_FD_SC_LP__O21BA_LP%X
x_PM_SKY130_FD_SC_LP__O21BA_LP%A_34_55# N_A_34_55#_M1001_s N_A_34_55#_M1002_d
+ N_A_34_55#_c_431_n N_A_34_55#_c_432_n N_A_34_55#_c_433_n N_A_34_55#_c_434_n
+ PM_SKY130_FD_SC_LP__O21BA_LP%A_34_55#
x_PM_SKY130_FD_SC_LP__O21BA_LP%VGND N_VGND_M1001_d N_VGND_M1003_d N_VGND_c_460_n
+ N_VGND_c_461_n VGND N_VGND_c_462_n N_VGND_c_463_n N_VGND_c_464_n
+ N_VGND_c_465_n N_VGND_c_466_n PM_SKY130_FD_SC_LP__O21BA_LP%VGND
cc_1 VNB N_A1_M1001_g 0.0456194f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.485
cc_2 VNB A1 0.0277145f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A1_c_82_n 0.0640531f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.28
cc_4 VNB N_A2_M1002_g 0.0367114f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.445
cc_5 VNB N_A2_c_109_n 0.0254369f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_A2_c_110_n 0.00247565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB A2 0.00170127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_c_112_n 0.0187663f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.28
cc_9 VNB N_A_317_29#_M1005_g 0.028149f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_A_317_29#_M1008_g 0.00575484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_317_29#_c_150_n 0.033944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_317_29#_c_151_n 0.0089078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_317_29#_c_152_n 0.0319919f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=1.28
cc_14 VNB N_A_317_29#_c_153_n 0.0112926f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.28
cc_15 VNB N_A_317_29#_c_154_n 0.00806486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_317_29#_c_155_n 0.0016576f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.45
cc_17 VNB N_A_317_29#_c_156_n 0.0253551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_317_29#_c_157_n 0.0244021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_N_M1007_g 0.0266935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_N_M1003_g 0.0242593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_N_c_218_n 0.026492f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=1.115
cc_22 VNB N_B1_N_c_219_n 0.00564076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB B1_N 0.00782535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_N_c_221_n 0.0231644f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.45
cc_25 VNB N_A_253_389#_M1011_g 0.0203184f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_26 VNB N_A_253_389#_M1009_g 0.0251596f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=1.28
cc_27 VNB N_A_253_389#_c_279_n 0.0101079f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=1.115
cc_28 VNB N_A_253_389#_c_280_n 0.00121962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_253_389#_c_281_n 0.0645421f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.45
cc_30 VNB N_A_253_389#_c_282_n 0.0091298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_366_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_410_n 0.0227724f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_33 VNB X 0.0425768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_34_55#_c_431_n 0.0215063f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_35 VNB N_A_34_55#_c_432_n 0.0222137f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_36 VNB N_A_34_55#_c_433_n 0.00984463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_34_55#_c_434_n 0.0030877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_460_n 0.0068875f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_39 VNB N_VGND_c_461_n 0.0116384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_462_n 0.0576122f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.28
cc_41 VNB N_VGND_c_463_n 0.0282798f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.45
cc_42 VNB N_VGND_c_464_n 0.276363f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.45
cc_43 VNB N_VGND_c_465_n 0.0264409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_466_n 0.00610336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A1_M1004_g 0.0309765f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.445
cc_46 VPB A1 0.0123908f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_47 VPB N_A1_c_82_n 0.0207877f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.28
cc_48 VPB N_A2_M1010_g 0.0253969f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=0.485
cc_49 VPB N_A2_c_110_n 0.0114324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB A2 0.00122131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_317_29#_M1008_g 0.0360247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_317_29#_c_155_n 0.00487629f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.45
cc_53 VPB N_A_317_29#_c_160_n 0.0112916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B1_N_c_222_n 0.0208762f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.115
cc_55 VPB N_B1_N_c_223_n 0.0424036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_B1_N_c_224_n 0.0170002f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.785
cc_57 VPB N_B1_N_c_225_n 0.0824787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_B1_N_c_219_n 0.0140186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB B1_N 0.00494378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_253_389#_M1006_g 0.0514306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_253_389#_c_279_n 0.00397134f $X=-0.19 $Y=1.655 $X2=0.497 $Y2=1.115
cc_62 VPB N_A_253_389#_c_285_n 0.0156084f $X=-0.19 $Y=1.655 $X2=0.497 $Y2=1.785
cc_63 VPB N_A_253_389#_c_281_n 0.00907824f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.45
cc_64 VPB N_A_253_389#_c_287_n 0.00887764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_253_389#_c_288_n 0.0029652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_253_389#_c_289_n 0.00264252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_367_n 0.0154644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_368_n 0.0483861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_369_n 0.00905631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_370_n 0.00655363f $X=-0.19 $Y=1.655 $X2=0.497 $Y2=1.115
cc_71 VPB N_VPWR_c_371_n 0.0315663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_372_n 0.00510584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_373_n 0.038698f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.45
cc_74 VPB N_VPWR_c_374_n 0.0185957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_366_n 0.0776837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_376_n 0.006319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB X 0.021167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB X 0.00899022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB X 0.0314291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 N_A1_M1001_g N_A2_M1002_g 0.0233503f $X=0.53 $Y=0.485 $X2=0 $Y2=0
cc_81 N_A1_M1004_g N_A2_c_110_n 0.0540132f $X=0.65 $Y=2.445 $X2=0 $Y2=0
cc_82 A1 A2 0.0540841f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A1_c_82_n A2 7.48253e-19 $X=0.385 $Y=1.28 $X2=0 $Y2=0
cc_84 A1 N_A2_c_112_n 0.00437388f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A1_c_82_n N_A2_c_112_n 0.0540132f $X=0.385 $Y=1.28 $X2=0 $Y2=0
cc_86 N_A1_M1004_g N_VPWR_c_368_n 0.030952f $X=0.65 $Y=2.445 $X2=0 $Y2=0
cc_87 A1 N_VPWR_c_368_n 0.0247387f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A1_c_82_n N_VPWR_c_368_n 0.00796239f $X=0.385 $Y=1.28 $X2=0 $Y2=0
cc_89 N_A1_M1004_g N_VPWR_c_373_n 0.00849388f $X=0.65 $Y=2.445 $X2=0 $Y2=0
cc_90 N_A1_M1004_g N_VPWR_c_366_n 0.00815197f $X=0.65 $Y=2.445 $X2=0 $Y2=0
cc_91 N_A1_M1001_g N_A_34_55#_c_431_n 0.00948802f $X=0.53 $Y=0.485 $X2=0 $Y2=0
cc_92 N_A1_M1001_g N_A_34_55#_c_432_n 0.00913445f $X=0.53 $Y=0.485 $X2=0 $Y2=0
cc_93 A1 N_A_34_55#_c_432_n 0.0267811f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A1_c_82_n N_A_34_55#_c_432_n 0.00444961f $X=0.385 $Y=1.28 $X2=0 $Y2=0
cc_95 N_A1_M1001_g N_A_34_55#_c_433_n 0.00419293f $X=0.53 $Y=0.485 $X2=0 $Y2=0
cc_96 A1 N_A_34_55#_c_433_n 0.0281902f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A1_c_82_n N_A_34_55#_c_433_n 0.00626078f $X=0.385 $Y=1.28 $X2=0 $Y2=0
cc_98 N_A1_M1001_g N_A_34_55#_c_434_n 8.74762e-19 $X=0.53 $Y=0.485 $X2=0 $Y2=0
cc_99 N_A1_M1001_g N_VGND_c_460_n 0.00493744f $X=0.53 $Y=0.485 $X2=0 $Y2=0
cc_100 N_A1_M1001_g N_VGND_c_464_n 0.00665445f $X=0.53 $Y=0.485 $X2=0 $Y2=0
cc_101 N_A1_M1001_g N_VGND_c_465_n 0.00511657f $X=0.53 $Y=0.485 $X2=0 $Y2=0
cc_102 N_A2_M1002_g N_A_317_29#_M1005_g 0.0198806f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_103 N_A2_M1010_g N_A_317_29#_M1008_g 0.0220665f $X=1.14 $Y=2.445 $X2=0 $Y2=0
cc_104 N_A2_c_110_n N_A_317_29#_M1008_g 0.00961611f $X=1.18 $Y=1.785 $X2=0 $Y2=0
cc_105 N_A2_c_109_n N_A_317_29#_c_153_n 0.00961611f $X=1.18 $Y=1.62 $X2=0 $Y2=0
cc_106 A2 N_A_317_29#_c_153_n 0.00145143f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A2_c_112_n N_A_317_29#_c_157_n 0.00201451f $X=1.18 $Y=1.28 $X2=0 $Y2=0
cc_108 N_A2_M1010_g N_A_253_389#_c_279_n 9.12975e-19 $X=1.14 $Y=2.445 $X2=0
+ $Y2=0
cc_109 N_A2_M1002_g N_A_253_389#_c_279_n 0.00205362f $X=1.12 $Y=0.485 $X2=0
+ $Y2=0
cc_110 N_A2_c_109_n N_A_253_389#_c_279_n 0.00114747f $X=1.18 $Y=1.62 $X2=0 $Y2=0
cc_111 A2 N_A_253_389#_c_279_n 0.0289129f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_112 N_A2_c_112_n N_A_253_389#_c_279_n 0.0041465f $X=1.18 $Y=1.28 $X2=0 $Y2=0
cc_113 N_A2_M1010_g N_A_253_389#_c_288_n 0.0022119f $X=1.14 $Y=2.445 $X2=0 $Y2=0
cc_114 N_A2_c_110_n N_A_253_389#_c_288_n 3.65856e-19 $X=1.18 $Y=1.785 $X2=0
+ $Y2=0
cc_115 A2 N_A_253_389#_c_288_n 0.00353019f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A2_M1002_g N_A_253_389#_c_282_n 3.04252e-19 $X=1.12 $Y=0.485 $X2=0
+ $Y2=0
cc_117 N_A2_M1010_g N_VPWR_c_368_n 0.00479847f $X=1.14 $Y=2.445 $X2=0 $Y2=0
cc_118 N_A2_M1010_g N_VPWR_c_373_n 0.00945281f $X=1.14 $Y=2.445 $X2=0 $Y2=0
cc_119 N_A2_M1010_g N_VPWR_c_366_n 0.00901766f $X=1.14 $Y=2.445 $X2=0 $Y2=0
cc_120 N_A2_M1002_g N_A_34_55#_c_431_n 8.74762e-19 $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_121 N_A2_M1002_g N_A_34_55#_c_432_n 0.0120622f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_122 A2 N_A_34_55#_c_432_n 0.0259718f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_123 N_A2_c_112_n N_A_34_55#_c_432_n 0.00134924f $X=1.18 $Y=1.28 $X2=0 $Y2=0
cc_124 N_A2_M1002_g N_A_34_55#_c_434_n 0.00868064f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_125 N_A2_M1002_g N_VGND_c_460_n 0.00493744f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_126 N_A2_M1002_g N_VGND_c_462_n 0.00511657f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_127 N_A2_M1002_g N_VGND_c_464_n 0.00610588f $X=1.12 $Y=0.485 $X2=0 $Y2=0
cc_128 N_A_317_29#_M1008_g N_B1_N_c_222_n 0.0300255f $X=1.71 $Y=2.445 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_317_29#_c_152_n N_B1_N_c_222_n 0.00482927f $X=2.03 $Y=1.5 $X2=-0.19
+ $Y2=-0.245
cc_130 N_A_317_29#_c_155_n N_B1_N_c_222_n 0.00580017f $X=2.54 $Y=1.925 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_317_29#_c_156_n N_B1_N_c_222_n 0.00490231f $X=2.195 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A_317_29#_c_160_n N_B1_N_c_222_n 0.00969259f $X=2.665 $Y=2.09 $X2=-0.19
+ $Y2=-0.245
cc_133 N_A_317_29#_c_150_n N_B1_N_M1007_g 0.00879168f $X=2.03 $Y=0.98 $X2=0
+ $Y2=0
cc_134 N_A_317_29#_c_154_n N_B1_N_M1007_g 0.0123259f $X=2.46 $Y=0.585 $X2=0
+ $Y2=0
cc_135 N_A_317_29#_c_156_n N_B1_N_M1007_g 0.00484085f $X=2.195 $Y=1.07 $X2=0
+ $Y2=0
cc_136 N_A_317_29#_c_154_n N_B1_N_M1003_g 0.00254015f $X=2.46 $Y=0.585 $X2=0
+ $Y2=0
cc_137 N_A_317_29#_c_155_n N_B1_N_c_225_n 0.00384883f $X=2.54 $Y=1.925 $X2=0
+ $Y2=0
cc_138 N_A_317_29#_c_160_n N_B1_N_c_225_n 0.00425798f $X=2.665 $Y=2.09 $X2=0
+ $Y2=0
cc_139 N_A_317_29#_c_156_n N_B1_N_c_218_n 0.00477548f $X=2.195 $Y=1.07 $X2=0
+ $Y2=0
cc_140 N_A_317_29#_c_157_n N_B1_N_c_218_n 0.00879168f $X=2.195 $Y=1.07 $X2=0
+ $Y2=0
cc_141 N_A_317_29#_c_155_n N_B1_N_c_219_n 0.00135807f $X=2.54 $Y=1.925 $X2=0
+ $Y2=0
cc_142 N_A_317_29#_c_160_n N_B1_N_c_219_n 2.6548e-19 $X=2.665 $Y=2.09 $X2=0
+ $Y2=0
cc_143 N_A_317_29#_c_156_n B1_N 0.0490774f $X=2.195 $Y=1.07 $X2=0 $Y2=0
cc_144 N_A_317_29#_c_157_n B1_N 3.94652e-19 $X=2.195 $Y=1.07 $X2=0 $Y2=0
cc_145 N_A_317_29#_c_160_n B1_N 7.99109e-19 $X=2.665 $Y=2.09 $X2=0 $Y2=0
cc_146 N_A_317_29#_c_156_n N_B1_N_c_221_n 0.00135807f $X=2.195 $Y=1.07 $X2=0
+ $Y2=0
cc_147 N_A_317_29#_c_157_n N_B1_N_c_221_n 0.00782396f $X=2.195 $Y=1.07 $X2=0
+ $Y2=0
cc_148 N_A_317_29#_M1005_g N_A_253_389#_c_279_n 0.0054862f $X=1.66 $Y=0.485
+ $X2=0 $Y2=0
cc_149 N_A_317_29#_M1008_g N_A_253_389#_c_279_n 0.0148618f $X=1.71 $Y=2.445
+ $X2=0 $Y2=0
cc_150 N_A_317_29#_c_150_n N_A_253_389#_c_279_n 0.00804759f $X=2.03 $Y=0.98
+ $X2=0 $Y2=0
cc_151 N_A_317_29#_c_151_n N_A_253_389#_c_279_n 0.00369221f $X=1.735 $Y=0.98
+ $X2=0 $Y2=0
cc_152 N_A_317_29#_c_152_n N_A_253_389#_c_279_n 0.00280474f $X=2.03 $Y=1.5 $X2=0
+ $Y2=0
cc_153 N_A_317_29#_c_153_n N_A_253_389#_c_279_n 0.00607015f $X=1.835 $Y=1.5
+ $X2=0 $Y2=0
cc_154 N_A_317_29#_c_154_n N_A_253_389#_c_279_n 0.00770613f $X=2.46 $Y=0.585
+ $X2=0 $Y2=0
cc_155 N_A_317_29#_c_155_n N_A_253_389#_c_279_n 0.0104673f $X=2.54 $Y=1.925
+ $X2=0 $Y2=0
cc_156 N_A_317_29#_c_156_n N_A_253_389#_c_279_n 0.0492887f $X=2.195 $Y=1.07
+ $X2=0 $Y2=0
cc_157 N_A_317_29#_c_157_n N_A_253_389#_c_279_n 0.00200266f $X=2.195 $Y=1.07
+ $X2=0 $Y2=0
cc_158 N_A_317_29#_c_160_n N_A_253_389#_c_279_n 8.02744e-19 $X=2.665 $Y=2.09
+ $X2=0 $Y2=0
cc_159 N_A_317_29#_M1000_d N_A_253_389#_c_285_n 0.00706364f $X=2.525 $Y=1.945
+ $X2=0 $Y2=0
cc_160 N_A_317_29#_c_160_n N_A_253_389#_c_285_n 0.0229256f $X=2.665 $Y=2.09
+ $X2=0 $Y2=0
cc_161 N_A_317_29#_c_160_n N_A_253_389#_c_287_n 0.0108144f $X=2.665 $Y=2.09
+ $X2=0 $Y2=0
cc_162 N_A_317_29#_M1008_g N_A_253_389#_c_288_n 0.0420989f $X=1.71 $Y=2.445
+ $X2=0 $Y2=0
cc_163 N_A_317_29#_M1005_g N_A_253_389#_c_282_n 0.00729611f $X=1.66 $Y=0.485
+ $X2=0 $Y2=0
cc_164 N_A_317_29#_c_150_n N_A_253_389#_c_282_n 0.00689537f $X=2.03 $Y=0.98
+ $X2=0 $Y2=0
cc_165 N_A_317_29#_c_154_n N_A_253_389#_c_282_n 0.0227533f $X=2.46 $Y=0.585
+ $X2=0 $Y2=0
cc_166 N_A_317_29#_c_156_n N_A_253_389#_c_282_n 6.3398e-19 $X=2.195 $Y=1.07
+ $X2=0 $Y2=0
cc_167 N_A_317_29#_M1008_g N_VPWR_c_369_n 0.00460802f $X=1.71 $Y=2.445 $X2=0
+ $Y2=0
cc_168 N_A_317_29#_M1008_g N_VPWR_c_373_n 0.00713612f $X=1.71 $Y=2.445 $X2=0
+ $Y2=0
cc_169 N_A_317_29#_M1008_g N_VPWR_c_366_n 0.00901766f $X=1.71 $Y=2.445 $X2=0
+ $Y2=0
cc_170 N_A_317_29#_M1005_g N_A_34_55#_c_432_n 0.00160984f $X=1.66 $Y=0.485 $X2=0
+ $Y2=0
cc_171 N_A_317_29#_M1005_g N_A_34_55#_c_434_n 0.00423268f $X=1.66 $Y=0.485 $X2=0
+ $Y2=0
cc_172 N_A_317_29#_c_154_n N_VGND_c_461_n 0.0153904f $X=2.46 $Y=0.585 $X2=0
+ $Y2=0
cc_173 N_A_317_29#_M1005_g N_VGND_c_462_n 0.00469294f $X=1.66 $Y=0.485 $X2=0
+ $Y2=0
cc_174 N_A_317_29#_c_154_n N_VGND_c_462_n 0.0142766f $X=2.46 $Y=0.585 $X2=0
+ $Y2=0
cc_175 N_A_317_29#_M1005_g N_VGND_c_464_n 0.00974404f $X=1.66 $Y=0.485 $X2=0
+ $Y2=0
cc_176 N_A_317_29#_c_154_n N_VGND_c_464_n 0.0119616f $X=2.46 $Y=0.585 $X2=0
+ $Y2=0
cc_177 N_B1_N_M1003_g N_A_253_389#_M1011_g 0.021188f $X=3.035 $Y=0.585 $X2=0
+ $Y2=0
cc_178 N_B1_N_c_219_n N_A_253_389#_M1006_g 0.0245876f $X=2.985 $Y=1.745 $X2=0
+ $Y2=0
cc_179 N_B1_N_c_222_n N_A_253_389#_c_279_n 0.001078f $X=2.4 $Y=3.02 $X2=0 $Y2=0
cc_180 N_B1_N_c_222_n N_A_253_389#_c_285_n 0.0245342f $X=2.4 $Y=3.02 $X2=0 $Y2=0
cc_181 N_B1_N_c_223_n N_A_253_389#_c_285_n 0.00516825f $X=3 $Y=3.095 $X2=0 $Y2=0
cc_182 N_B1_N_c_225_n N_A_253_389#_c_285_n 0.0184367f $X=3.075 $Y=3.02 $X2=0
+ $Y2=0
cc_183 N_B1_N_c_219_n N_A_253_389#_c_285_n 0.00413607f $X=2.985 $Y=1.745 $X2=0
+ $Y2=0
cc_184 N_B1_N_M1003_g N_A_253_389#_c_280_n 4.72661e-19 $X=3.035 $Y=0.585 $X2=0
+ $Y2=0
cc_185 N_B1_N_c_218_n N_A_253_389#_c_280_n 3.03985e-19 $X=3.035 $Y=1.15 $X2=0
+ $Y2=0
cc_186 B1_N N_A_253_389#_c_280_n 0.0517714f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_187 N_B1_N_c_218_n N_A_253_389#_c_281_n 0.0319932f $X=3.035 $Y=1.15 $X2=0
+ $Y2=0
cc_188 B1_N N_A_253_389#_c_281_n 0.00405558f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_189 N_B1_N_c_219_n N_A_253_389#_c_287_n 0.0108574f $X=2.985 $Y=1.745 $X2=0
+ $Y2=0
cc_190 N_B1_N_c_222_n N_A_253_389#_c_288_n 8.64799e-19 $X=2.4 $Y=3.02 $X2=0
+ $Y2=0
cc_191 N_B1_N_M1007_g N_A_253_389#_c_282_n 0.00299393f $X=2.675 $Y=0.585 $X2=0
+ $Y2=0
cc_192 N_B1_N_c_221_n N_A_253_389#_c_289_n 3.03985e-19 $X=2.985 $Y=1.24 $X2=0
+ $Y2=0
cc_193 N_B1_N_c_222_n N_VPWR_c_369_n 0.00880971f $X=2.4 $Y=3.02 $X2=0 $Y2=0
cc_194 N_B1_N_c_225_n N_VPWR_c_370_n 0.00924075f $X=3.075 $Y=3.02 $X2=0 $Y2=0
cc_195 N_B1_N_c_224_n N_VPWR_c_371_n 0.0218672f $X=2.525 $Y=3.095 $X2=0 $Y2=0
cc_196 N_B1_N_c_223_n N_VPWR_c_366_n 0.0192872f $X=3 $Y=3.095 $X2=0 $Y2=0
cc_197 N_B1_N_c_224_n N_VPWR_c_366_n 0.00896019f $X=2.525 $Y=3.095 $X2=0 $Y2=0
cc_198 N_B1_N_M1007_g N_VGND_c_461_n 0.00180376f $X=2.675 $Y=0.585 $X2=0 $Y2=0
cc_199 N_B1_N_M1003_g N_VGND_c_461_n 0.012273f $X=3.035 $Y=0.585 $X2=0 $Y2=0
cc_200 N_B1_N_c_218_n N_VGND_c_461_n 0.00102988f $X=3.035 $Y=1.15 $X2=0 $Y2=0
cc_201 B1_N N_VGND_c_461_n 0.00989998f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_202 N_B1_N_M1007_g N_VGND_c_462_n 0.00430542f $X=2.675 $Y=0.585 $X2=0 $Y2=0
cc_203 N_B1_N_M1003_g N_VGND_c_462_n 0.00379792f $X=3.035 $Y=0.585 $X2=0 $Y2=0
cc_204 N_B1_N_M1007_g N_VGND_c_464_n 0.00544287f $X=2.675 $Y=0.585 $X2=0 $Y2=0
cc_205 N_B1_N_M1003_g N_VGND_c_464_n 0.00457201f $X=3.035 $Y=0.585 $X2=0 $Y2=0
cc_206 N_A_253_389#_c_285_n N_VPWR_M1008_d 0.0166411f $X=3.415 $Y=2.52 $X2=0
+ $Y2=0
cc_207 N_A_253_389#_c_285_n N_VPWR_M1006_s 0.00809225f $X=3.415 $Y=2.52 $X2=0
+ $Y2=0
cc_208 N_A_253_389#_c_287_n N_VPWR_M1006_s 0.0111458f $X=3.5 $Y=2.435 $X2=0
+ $Y2=0
cc_209 N_A_253_389#_c_285_n N_VPWR_c_369_n 0.0242699f $X=3.415 $Y=2.52 $X2=0
+ $Y2=0
cc_210 N_A_253_389#_c_288_n N_VPWR_c_369_n 0.00658467f $X=1.445 $Y=2.13 $X2=0
+ $Y2=0
cc_211 N_A_253_389#_M1006_g N_VPWR_c_370_n 0.0128241f $X=3.775 $Y=2.595 $X2=0
+ $Y2=0
cc_212 N_A_253_389#_c_285_n N_VPWR_c_370_n 0.0190544f $X=3.415 $Y=2.52 $X2=0
+ $Y2=0
cc_213 N_A_253_389#_c_285_n N_VPWR_c_371_n 0.0153401f $X=3.415 $Y=2.52 $X2=0
+ $Y2=0
cc_214 N_A_253_389#_c_288_n N_VPWR_c_373_n 0.0189483f $X=1.445 $Y=2.13 $X2=0
+ $Y2=0
cc_215 N_A_253_389#_M1006_g N_VPWR_c_374_n 0.00840199f $X=3.775 $Y=2.595 $X2=0
+ $Y2=0
cc_216 N_A_253_389#_M1006_g N_VPWR_c_366_n 0.0145244f $X=3.775 $Y=2.595 $X2=0
+ $Y2=0
cc_217 N_A_253_389#_c_285_n N_VPWR_c_366_n 0.0295909f $X=3.415 $Y=2.52 $X2=0
+ $Y2=0
cc_218 N_A_253_389#_c_288_n N_VPWR_c_366_n 0.0191735f $X=1.445 $Y=2.13 $X2=0
+ $Y2=0
cc_219 N_A_253_389#_M1011_g N_X_c_410_n 0.00125204f $X=3.465 $Y=0.585 $X2=0
+ $Y2=0
cc_220 N_A_253_389#_M1009_g N_X_c_410_n 0.0101733f $X=3.825 $Y=0.585 $X2=0 $Y2=0
cc_221 N_A_253_389#_M1009_g X 0.0375896f $X=3.825 $Y=0.585 $X2=0 $Y2=0
cc_222 N_A_253_389#_c_280_n X 0.0425941f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A_253_389#_c_287_n X 0.0180511f $X=3.5 $Y=2.435 $X2=0 $Y2=0
cc_224 N_A_253_389#_M1006_g X 0.00427623f $X=3.775 $Y=2.595 $X2=0 $Y2=0
cc_225 N_A_253_389#_c_287_n X 0.0176154f $X=3.5 $Y=2.435 $X2=0 $Y2=0
cc_226 N_A_253_389#_M1006_g X 0.0244355f $X=3.775 $Y=2.595 $X2=0 $Y2=0
cc_227 N_A_253_389#_c_285_n X 0.00931262f $X=3.415 $Y=2.52 $X2=0 $Y2=0
cc_228 N_A_253_389#_c_279_n N_A_34_55#_c_432_n 0.0131057f $X=1.765 $Y=1.965
+ $X2=0 $Y2=0
cc_229 N_A_253_389#_c_282_n N_A_34_55#_c_434_n 0.03723f $X=1.875 $Y=0.49 $X2=0
+ $Y2=0
cc_230 N_A_253_389#_M1011_g N_VGND_c_461_n 0.0130814f $X=3.465 $Y=0.585 $X2=0
+ $Y2=0
cc_231 N_A_253_389#_M1009_g N_VGND_c_461_n 0.00180376f $X=3.825 $Y=0.585 $X2=0
+ $Y2=0
cc_232 N_A_253_389#_c_282_n N_VGND_c_462_n 0.0235651f $X=1.875 $Y=0.49 $X2=0
+ $Y2=0
cc_233 N_A_253_389#_M1011_g N_VGND_c_463_n 0.00379792f $X=3.465 $Y=0.585 $X2=0
+ $Y2=0
cc_234 N_A_253_389#_M1009_g N_VGND_c_463_n 0.00430542f $X=3.825 $Y=0.585 $X2=0
+ $Y2=0
cc_235 N_A_253_389#_M1011_g N_VGND_c_464_n 0.00457201f $X=3.465 $Y=0.585 $X2=0
+ $Y2=0
cc_236 N_A_253_389#_M1009_g N_VGND_c_464_n 0.00544287f $X=3.825 $Y=0.585 $X2=0
+ $Y2=0
cc_237 N_A_253_389#_c_282_n N_VGND_c_464_n 0.013524f $X=1.875 $Y=0.49 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_366_n N_X_M1006_d 0.0023218f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_c_370_n X 0.0184494f $X=3.51 $Y=2.95 $X2=0 $Y2=0
cc_240 N_VPWR_c_374_n X 0.019758f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_241 N_VPWR_c_366_n X 0.012508f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_242 N_X_c_410_n N_VGND_c_461_n 0.0153904f $X=4.04 $Y=0.585 $X2=0 $Y2=0
cc_243 N_X_c_410_n N_VGND_c_463_n 0.0141724f $X=4.04 $Y=0.585 $X2=0 $Y2=0
cc_244 N_X_c_410_n N_VGND_c_464_n 0.0119193f $X=4.04 $Y=0.585 $X2=0 $Y2=0
cc_245 N_A_34_55#_c_431_n N_VGND_c_460_n 0.0118289f $X=0.315 $Y=0.49 $X2=0 $Y2=0
cc_246 N_A_34_55#_c_432_n N_VGND_c_460_n 0.0249995f $X=1.17 $Y=0.85 $X2=0 $Y2=0
cc_247 N_A_34_55#_c_434_n N_VGND_c_460_n 0.0118289f $X=1.335 $Y=0.49 $X2=0 $Y2=0
cc_248 N_A_34_55#_c_434_n N_VGND_c_462_n 0.0220075f $X=1.335 $Y=0.49 $X2=0 $Y2=0
cc_249 N_A_34_55#_c_431_n N_VGND_c_464_n 0.0125757f $X=0.315 $Y=0.49 $X2=0 $Y2=0
cc_250 N_A_34_55#_c_432_n N_VGND_c_464_n 0.0127264f $X=1.17 $Y=0.85 $X2=0 $Y2=0
cc_251 N_A_34_55#_c_434_n N_VGND_c_464_n 0.0125757f $X=1.335 $Y=0.49 $X2=0 $Y2=0
cc_252 N_A_34_55#_c_431_n N_VGND_c_465_n 0.0220075f $X=0.315 $Y=0.49 $X2=0 $Y2=0
