* File: sky130_fd_sc_lp__fahcon_1.spice
* Created: Wed Sep  2 09:53:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__fahcon_1.pex.spice"
.subckt sky130_fd_sc_lp__fahcon_1  VNB VPB A B CI VPWR COUT_N SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT_N	COUT_N
* VPWR	VPWR
* CI	CI
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_A_M1025_g N_A_33_367#_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.264827 AS=0.2394 PD=1.68 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1003 N_A_247_367#_M1003_d N_A_33_367#_M1003_g N_VGND_M1025_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.201773 PD=0.92 PS=1.28 NRD=0 NRS=68.436 M=1 R=4.26667
+ SA=75001 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1029 N_A_367_119#_M1029_d N_A_329_269#_M1029_g N_A_247_367#_M1003_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1292 AS=0.0896 PD=1.075 PS=0.92 NRD=21.552 NRS=0 M=1
+ R=4.26667 SA=75001.4 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1005 N_A_33_367#_M1005_d N_B_M1005_g N_A_367_119#_M1029_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0976 AS=0.1292 PD=0.945 PS=1.075 NRD=3.744 NRS=0 M=1 R=4.26667
+ SA=75001.9 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1001 N_A_359_367#_M1001_d N_A_329_269#_M1001_g N_A_33_367#_M1005_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1984 AS=0.0976 PD=1.26 PS=0.945 NRD=22.488 NRS=0.936 M=1
+ R=4.26667 SA=75002.3 SB=75001 A=0.096 P=1.58 MULT=1
MM1031 N_A_247_367#_M1031_d N_B_M1031_g N_A_359_367#_M1001_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.1984 PD=1.85 PS=1.26 NRD=0 NRS=41.244 M=1 R=4.26667
+ SA=75003.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_B_M1011_g N_A_329_269#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.322946 AS=0.3066 PD=1.86162 PS=2.41 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.3
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1008 N_A_1034_380#_M1008_d N_B_M1008_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0896 AS=0.246054 PD=0.92 PS=1.41838 NRD=0 NRS=97.968 M=1 R=4.26667
+ SA=75001.2 SB=75004.4 A=0.096 P=1.58 MULT=1
MM1020 N_COUT_N_M1020_d N_A_359_367#_M1020_g N_A_1034_380#_M1008_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1776 AS=0.0896 PD=1.195 PS=0.92 NRD=14.988 NRS=0 M=1
+ R=4.26667 SA=75001.7 SB=75003.9 A=0.096 P=1.58 MULT=1
MM1009 N_A_1340_412#_M1009_d N_A_367_119#_M1009_g N_COUT_N_M1020_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2179 AS=0.1776 PD=1.425 PS=1.195 NRD=40.776 NRS=36.552 M=1
+ R=4.26667 SA=75002.4 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1016 N_VGND_M1016_d N_CI_M1016_g N_A_1340_412#_M1009_d VNB NSHORT L=0.15
+ W=0.64 AD=0.132151 AS=0.2179 PD=1.06378 PS=1.425 NRD=20.148 NRS=20.148 M=1
+ R=4.26667 SA=75002.3 SB=75003.6 A=0.096 P=1.58 MULT=1
MM1012 N_A_1571_367#_M1012_d N_CI_M1012_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.84 AD=0.175832 AS=0.173449 PD=1.40189 PS=1.39622 NRD=0 NRS=0.708 M=1 R=5.6
+ SA=75002.2 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1002 N_A_1758_87#_M1002_d N_A_359_367#_M1002_g N_A_1571_367#_M1012_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1728 AS=0.133968 PD=1.18 PS=1.06811 NRD=0 NRS=22.02
+ M=1 R=4.26667 SA=75003.4 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1019 N_A_1708_411#_M1019_d N_A_367_119#_M1019_g N_A_1758_87#_M1002_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.192 AS=0.1728 PD=1.24 PS=1.18 NRD=60 NRS=48.744 M=1
+ R=4.26667 SA=75004.1 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_A_1571_367#_M1015_g N_A_1708_411#_M1019_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.233859 AS=0.192 PD=1.34919 PS=1.24 NRD=58.2 NRS=0 M=1
+ R=4.26667 SA=75004.8 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1017 N_SUM_M1017_d N_A_1758_87#_M1017_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.306941 PD=2.25 PS=1.77081 NRD=0 NRS=16.428 M=1 R=5.6
+ SA=75004.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1030 N_VPWR_M1030_d N_A_M1030_g N_A_33_367#_M1030_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.323307 AS=0.3591 PD=1.94575 PS=3.09 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1021 N_A_247_367#_M1021_d N_A_33_367#_M1021_g N_VPWR_M1030_d VPB PHIGHVT
+ L=0.15 W=1 AD=0.211957 AS=0.256593 PD=1.53261 PS=1.54425 NRD=0 NRS=24.6053 M=1
+ R=6.66667 SA=75000.8 SB=75002 A=0.15 P=2.3 MULT=1
MM1022 N_A_359_367#_M1022_d N_A_329_269#_M1022_g N_A_247_367#_M1021_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2107 AS=0.178043 PD=1.38 PS=1.28739 NRD=51.5943
+ NRS=31.0669 M=1 R=5.6 SA=75001.4 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1013 N_A_33_367#_M1013_d N_B_M1013_g N_A_359_367#_M1022_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1176 AS=0.2107 PD=1.12 PS=1.38 NRD=0 NRS=0 M=1 R=5.6 SA=75002
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1000 N_A_367_119#_M1000_d N_A_329_269#_M1000_g N_A_33_367#_M1013_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2198 AS=0.1176 PD=1.455 PS=1.12 NRD=19.9167 NRS=0 M=1 R=5.6
+ SA=75002.4 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1018 N_A_247_367#_M1018_d N_B_M1018_g N_A_367_119#_M1000_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2352 AS=0.2198 PD=2.24 PS=1.455 NRD=0 NRS=28.1316 M=1 R=5.6
+ SA=75003 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1027 N_VPWR_M1027_d N_B_M1027_g N_A_329_269#_M1027_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.337245 AS=0.3528 PD=1.97363 PS=3.08 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.5 A=0.189 P=2.82 MULT=1
MM1024 N_A_1034_380#_M1024_d N_B_M1024_g N_VPWR_M1027_d VPB PHIGHVT L=0.15 W=1
+ AD=0.216522 AS=0.267655 PD=1.54348 PS=1.56637 NRD=0 NRS=50.7275 M=1 R=6.66667
+ SA=75000.9 SB=75002.4 A=0.15 P=2.3 MULT=1
MM1010 N_COUT_N_M1010_d N_A_367_119#_M1010_g N_A_1034_380#_M1024_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.3402 AS=0.181878 PD=1.65 PS=1.29652 NRD=37.5088 NRS=33.2142
+ M=1 R=5.6 SA=75001.4 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1014 N_A_1340_412#_M1014_d N_A_359_367#_M1014_g N_COUT_N_M1010_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.226104 AS=0.3402 PD=1.42435 PS=1.65 NRD=24.625 NRS=86.7588
+ M=1 R=5.6 SA=75002.4 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1026 N_VPWR_M1026_d N_CI_M1026_g N_A_1340_412#_M1014_d VPB PHIGHVT L=0.15 W=1
+ AD=0.188053 AS=0.269171 PD=1.43363 PS=1.69565 NRD=0 NRS=21.9852 M=1 R=6.66667
+ SA=75002.4 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1023 N_A_1571_367#_M1023_d N_CI_M1023_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.236947 PD=3.09 PS=1.80637 NRD=0 NRS=12.4898 M=1 R=8.4
+ SA=75002.4 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1006 N_A_1758_87#_M1006_d N_A_359_367#_M1006_g N_A_1708_411#_M1006_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1176 AS=0.4027 PD=1.12 PS=2.94 NRD=0 NRS=99.5244
+ M=1 R=5.6 SA=75000.3 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1028 N_A_1571_367#_M1028_d N_A_367_119#_M1028_g N_A_1758_87#_M1006_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_A_1571_367#_M1007_g N_A_1708_411#_M1007_s VPB PHIGHVT
+ L=0.15 W=1 AD=0.201991 AS=0.285 PD=1.45575 PS=2.57 NRD=20.685 NRS=0 M=1
+ R=6.66667 SA=75000.2 SB=75000.7 A=0.15 P=2.3 MULT=1
MM1004 N_SUM_M1004_d N_A_1758_87#_M1004_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3402 AS=0.254509 PD=3.06 PS=1.83425 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=22.3225 P=27.61
*
.include "sky130_fd_sc_lp__fahcon_1.pxi.spice"
*
.ends
*
*
