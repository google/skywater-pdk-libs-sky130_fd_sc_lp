# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__busdrivernovlpsleep_20
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__busdrivernovlpsleep_20 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  23.52000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.400000 0.440000 12.385000 0.770000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  1.228000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  0.625000 1.920000  0.915000 1.950000 ;
        RECT  0.625000 1.950000 12.010000 2.120000 ;
        RECT  0.625000 2.120000  0.915000 2.150000 ;
        RECT  5.355000 1.920000  5.645000 1.950000 ;
        RECT  5.355000 2.120000  5.645000 2.150000 ;
        RECT 11.720000 1.920000 12.010000 1.950000 ;
        RECT 11.720000 2.120000 12.010000 2.150000 ;
    END
  END SLEEP
  PIN TE_B
    ANTENNAGATEAREA  0.348000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035000 1.200000 2.415000 1.590000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  4.968000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 14.480000 1.920000 22.510000 2.150000 ;
    END
  END Z
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.675000 23.450000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 23.520000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 23.520000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 23.710000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 23.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 23.520000 0.085000 ;
      RECT  0.000000  3.245000 23.520000 3.415000 ;
      RECT  0.095000  0.255000  0.425000 3.075000 ;
      RECT  0.595000  1.200000  0.925000 2.150000 ;
      RECT  0.625000  2.320000  0.955000 3.245000 ;
      RECT  0.945000  0.085000  1.250000 1.020000 ;
      RECT  1.420000  0.255000  1.635000 0.860000 ;
      RECT  1.420000  0.860000  2.550000 1.030000 ;
      RECT  1.420000  1.030000  1.625000 1.760000 ;
      RECT  1.420000  1.760000  3.165000 1.930000 ;
      RECT  1.475000  1.930000  1.805000 3.065000 ;
      RECT  1.805000  0.085000  2.135000 0.690000 ;
      RECT  1.995000  2.100000  3.505000 2.270000 ;
      RECT  1.995000  2.270000  2.325000 3.075000 ;
      RECT  2.305000  0.255000  2.550000 0.860000 ;
      RECT  2.495000  2.440000  3.400000 3.075000 ;
      RECT  2.720000  0.085000  2.995000 1.040000 ;
      RECT  2.900000  1.345000  3.165000 1.760000 ;
      RECT  3.185000  0.275000  3.505000 0.605000 ;
      RECT  3.335000  0.605000  3.505000 0.645000 ;
      RECT  3.335000  0.645000  5.455000 0.815000 ;
      RECT  3.335000  0.815000  3.505000 2.100000 ;
      RECT  3.675000  0.085000  5.110000 0.475000 ;
      RECT  3.675000  0.985000  6.015000 1.155000 ;
      RECT  3.675000  1.155000  3.895000 3.065000 ;
      RECT  4.065000  1.850000  4.315000 3.045000 ;
      RECT  4.485000  1.325000  4.815000 1.815000 ;
      RECT  4.485000  2.060000  4.715000 2.325000 ;
      RECT  4.485000  2.325000  6.525000 2.495000 ;
      RECT  4.485000  2.495000  4.715000 3.070000 ;
      RECT  4.885000  2.665000  5.215000 3.015000 ;
      RECT  5.270000  1.765000  5.675000 2.155000 ;
      RECT  5.285000  0.265000  6.695000 0.435000 ;
      RECT  5.285000  0.435000  5.455000 0.645000 ;
      RECT  5.405000  2.665000  5.735000 3.245000 ;
      RECT  5.660000  0.605000  6.355000 0.815000 ;
      RECT  5.845000  1.155000  6.015000 1.550000 ;
      RECT  5.845000  1.550000  6.760000 1.720000 ;
      RECT  6.185000  0.815000  6.355000 1.200000 ;
      RECT  6.185000  1.200000  7.230000 1.370000 ;
      RECT  6.195000  2.085000  7.230000 2.255000 ;
      RECT  6.195000  2.255000  6.525000 2.325000 ;
      RECT  6.195000  2.495000  6.525000 3.065000 ;
      RECT  6.335000  1.720000  6.760000 1.905000 ;
      RECT  6.525000  0.435000  6.695000 0.850000 ;
      RECT  6.525000  0.850000  7.565000 1.020000 ;
      RECT  6.705000  2.435000  6.955000 3.245000 ;
      RECT  6.970000  1.370000  7.230000 2.085000 ;
      RECT  6.975000  0.085000  7.225000 0.680000 ;
      RECT  7.395000  0.265000  8.245000 0.435000 ;
      RECT  7.395000  0.435000  7.565000 0.850000 ;
      RECT  7.500000  1.815000  7.750000 2.895000 ;
      RECT  7.500000  2.895000  8.610000 3.065000 ;
      RECT  7.735000  0.605000  7.905000 0.995000 ;
      RECT  7.735000  0.995000  9.745000 1.165000 ;
      RECT  7.735000  1.165000  8.110000 1.225000 ;
      RECT  7.920000  1.225000  8.110000 2.715000 ;
      RECT  8.075000  0.435000  8.245000 0.655000 ;
      RECT  8.075000  0.655000 10.155000 0.825000 ;
      RECT  8.280000  1.815000  8.610000 2.320000 ;
      RECT  8.280000  2.320000  9.470000 2.500000 ;
      RECT  8.280000  2.500000  8.610000 2.895000 ;
      RECT  8.415000  0.085000  8.785000 0.465000 ;
      RECT  8.780000  2.670000  9.040000 3.245000 ;
      RECT  9.210000  2.500000  9.470000 3.065000 ;
      RECT  9.455000  0.085000 10.190000 0.485000 ;
      RECT  9.455000  1.165000  9.745000 1.505000 ;
      RECT  9.710000  1.845000 10.040000 3.245000 ;
      RECT  9.985000  0.825000 10.155000 0.995000 ;
      RECT  9.985000  0.995000 10.315000 1.325000 ;
      RECT 10.360000  0.265000 10.550000 0.645000 ;
      RECT 10.360000  0.645000 11.140000 0.815000 ;
      RECT 10.485000  0.995000 10.800000 1.665000 ;
      RECT 10.500000  1.845000 11.140000 2.015000 ;
      RECT 10.500000  2.015000 10.830000 2.725000 ;
      RECT 10.720000  0.085000 11.050000 0.465000 ;
      RECT 10.970000  0.815000 11.140000 0.955000 ;
      RECT 10.970000  0.955000 12.455000 1.130000 ;
      RECT 10.970000  1.130000 11.140000 1.845000 ;
      RECT 11.270000  2.320000 11.530000 3.245000 ;
      RECT 11.445000  1.325000 12.115000 1.615000 ;
      RECT 11.700000  2.320000 12.980000 2.490000 ;
      RECT 11.700000  2.490000 12.030000 3.035000 ;
      RECT 11.710000  1.615000 12.055000 2.150000 ;
      RECT 12.200000  2.735000 12.460000 3.245000 ;
      RECT 12.285000  1.130000 12.455000 1.275000 ;
      RECT 12.285000  1.275000 14.030000 1.605000 ;
      RECT 12.555000  0.295000 12.885000 0.465000 ;
      RECT 12.650000  2.185000 12.980000 2.320000 ;
      RECT 12.650000  2.490000 12.980000 2.775000 ;
      RECT 12.650000  2.775000 13.840000 3.075000 ;
      RECT 12.680000  0.465000 12.885000 0.925000 ;
      RECT 12.680000  0.925000 13.905000 1.095000 ;
      RECT 13.055000  0.085000 13.365000 0.755000 ;
      RECT 13.150000  1.785000 14.370000 1.955000 ;
      RECT 13.150000  1.955000 13.410000 2.605000 ;
      RECT 13.575000  0.265000 14.790000 0.435000 ;
      RECT 13.575000  0.435000 13.905000 0.925000 ;
      RECT 13.590000  2.185000 13.840000 2.775000 ;
      RECT 14.025000  2.135000 14.360000 3.245000 ;
      RECT 14.075000  0.615000 14.370000 1.095000 ;
      RECT 14.200000  1.095000 14.370000 1.550000 ;
      RECT 14.200000  1.550000 14.860000 1.780000 ;
      RECT 14.200000  1.780000 14.370000 1.785000 ;
      RECT 14.540000  0.435000 14.790000 1.095000 ;
      RECT 14.540000  1.950000 15.650000 2.130000 ;
      RECT 14.540000  2.130000 14.710000 3.065000 ;
      RECT 14.890000  2.310000 15.140000 3.245000 ;
      RECT 14.960000  1.035000 15.150000 1.410000 ;
      RECT 15.320000  0.255000 15.650000 1.950000 ;
      RECT 15.320000  2.130000 15.650000 3.065000 ;
      RECT 15.820000  1.035000 16.010000 1.410000 ;
      RECT 15.830000  0.085000 16.000000 0.865000 ;
      RECT 15.830000  2.290000 16.000000 3.245000 ;
      RECT 16.180000  0.255000 16.510000 3.065000 ;
      RECT 16.680000  1.035000 16.870000 1.410000 ;
      RECT 16.690000  0.085000 16.860000 0.865000 ;
      RECT 16.690000  2.290000 16.860000 3.245000 ;
      RECT 17.040000  0.255000 17.370000 3.065000 ;
      RECT 17.540000  1.035000 17.730000 1.410000 ;
      RECT 17.550000  0.085000 17.720000 0.865000 ;
      RECT 17.550000  2.290000 17.720000 3.245000 ;
      RECT 17.900000  0.255000 18.230000 3.065000 ;
      RECT 18.400000  1.035000 18.590000 1.410000 ;
      RECT 18.410000  0.085000 18.580000 0.865000 ;
      RECT 18.410000  2.290000 18.580000 3.245000 ;
      RECT 18.760000  0.255000 19.090000 3.065000 ;
      RECT 19.260000  1.345000 19.450000 1.760000 ;
      RECT 19.270000  0.085000 19.440000 0.865000 ;
      RECT 19.270000  2.290000 19.440000 3.245000 ;
      RECT 19.620000  0.255000 19.950000 3.065000 ;
      RECT 20.120000  1.345000 20.310000 1.760000 ;
      RECT 20.130000  0.085000 20.300000 0.865000 ;
      RECT 20.130000  2.290000 20.300000 3.245000 ;
      RECT 20.480000  0.260000 20.810000 3.065000 ;
      RECT 20.980000  1.345000 21.170000 1.760000 ;
      RECT 20.990000  0.085000 21.160000 0.865000 ;
      RECT 20.990000  2.290000 21.160000 3.245000 ;
      RECT 21.340000  0.255000 21.670000 3.065000 ;
      RECT 21.840000  1.345000 22.430000 1.760000 ;
      RECT 21.850000  2.290000 22.020000 3.245000 ;
      RECT 22.200000  1.940000 22.530000 3.065000 ;
      RECT 22.710000  2.290000 22.960000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  1.580000  0.325000 1.750000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  0.685000  1.950000  0.855000 2.120000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.500000  2.715000  2.670000 2.885000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  2.860000  2.715000  3.030000 2.885000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.220000  2.715000  3.390000 2.885000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.105000  2.715000  4.275000 2.885000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.565000  1.580000  4.735000 1.750000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  2.715000  5.125000 2.885000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.415000  1.950000  5.585000 2.120000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.580000  6.565000 1.750000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.515000  1.210000  9.685000 1.380000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.485000  1.210000 10.655000 1.380000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 11.780000  1.950000 11.950000 2.120000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 14.595000  1.580000 14.765000 1.750000 ;
      RECT 14.980000  1.210000 15.150000 1.380000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.400000  1.950000 15.570000 2.120000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.840000  1.210000 16.010000 1.380000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.260000  1.950000 16.430000 2.120000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.700000  1.210000 16.870000 1.380000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.120000  1.950000 17.290000 2.120000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
      RECT 17.560000  1.210000 17.730000 1.380000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.245000 18.085000 3.415000 ;
      RECT 17.980000  1.950000 18.150000 2.120000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.245000 18.565000 3.415000 ;
      RECT 18.420000  1.210000 18.590000 1.380000 ;
      RECT 18.840000  1.950000 19.010000 2.120000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.245000 19.045000 3.415000 ;
      RECT 19.260000  1.580000 19.430000 1.750000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  3.245000 19.525000 3.415000 ;
      RECT 19.700000  1.950000 19.870000 2.120000 ;
      RECT 19.835000 -0.085000 20.005000 0.085000 ;
      RECT 19.835000  3.245000 20.005000 3.415000 ;
      RECT 20.120000  1.580000 20.290000 1.750000 ;
      RECT 20.315000 -0.085000 20.485000 0.085000 ;
      RECT 20.315000  3.245000 20.485000 3.415000 ;
      RECT 20.560000  1.950000 20.730000 2.120000 ;
      RECT 20.795000 -0.085000 20.965000 0.085000 ;
      RECT 20.795000  3.245000 20.965000 3.415000 ;
      RECT 20.980000  1.580000 21.150000 1.750000 ;
      RECT 21.275000 -0.085000 21.445000 0.085000 ;
      RECT 21.275000  3.245000 21.445000 3.415000 ;
      RECT 21.420000  1.950000 21.590000 2.120000 ;
      RECT 21.755000 -0.085000 21.925000 0.085000 ;
      RECT 21.755000  3.245000 21.925000 3.415000 ;
      RECT 21.840000  1.580000 22.010000 1.750000 ;
      RECT 22.200000  1.580000 22.370000 1.750000 ;
      RECT 22.235000 -0.085000 22.405000 0.085000 ;
      RECT 22.235000  3.245000 22.405000 3.415000 ;
      RECT 22.280000  1.950000 22.450000 2.120000 ;
      RECT 22.715000 -0.085000 22.885000 0.085000 ;
      RECT 22.715000  3.245000 22.885000 3.415000 ;
      RECT 23.195000 -0.085000 23.365000 0.085000 ;
      RECT 23.195000  3.245000 23.365000 3.415000 ;
    LAYER met1 ;
      RECT  0.095000 1.550000  0.385000 1.595000 ;
      RECT  0.095000 1.595000  4.795000 1.735000 ;
      RECT  0.095000 1.735000  0.385000 1.780000 ;
      RECT  4.505000 1.550000  4.795000 1.595000 ;
      RECT  4.505000 1.735000  4.795000 1.780000 ;
      RECT  6.335000 1.550000  6.625000 1.595000 ;
      RECT  6.335000 1.595000 22.465000 1.735000 ;
      RECT  6.335000 1.735000  6.625000 1.780000 ;
      RECT  9.455000 1.180000  9.745000 1.225000 ;
      RECT  9.455000 1.225000 18.695000 1.365000 ;
      RECT  9.455000 1.365000  9.745000 1.410000 ;
      RECT 10.425000 1.180000 10.715000 1.225000 ;
      RECT 10.425000 1.365000 10.715000 1.410000 ;
      RECT 14.500000 1.735000 22.465000 1.780000 ;
      RECT 14.505000 1.550000 22.465000 1.595000 ;
      RECT 14.920000 1.180000 18.695000 1.225000 ;
      RECT 14.920000 1.365000 18.695000 1.410000 ;
  END
END sky130_fd_sc_lp__busdrivernovlpsleep_20
END LIBRARY
