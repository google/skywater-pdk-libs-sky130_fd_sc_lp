* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_lp__sleep_sergate_plv_21 VIRTPWR VPWR SLEEP VPB
*.PININFO VIRTPWR:? VPWR:? SLEEP:? VPB:?
M1000 VIRTPWR SLEEP VPB phighvt w=7e+06u l=150000u ad=3.815e+12p
+ pd=2.909e+07u as=3.815e+12p ps=2.909e+07u
M1001 VIRTPWR SLEEP VPB phighvt w=7e+06u l=150000u ad=0p pd=0u as=0p
+ ps=0u
M1002 VPWR SLEEP VPB phighvt w=7e+06u l=150000u ad=0p pd=0u as=0p
+ ps=0u
.ENDS sky130_fd_sc_lp__sleep_sergate_plv_21
