* File: sky130_fd_sc_lp__a31o_lp.spice
* Created: Wed Sep  2 09:26:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a31o_lp.pex.spice"
.subckt sky130_fd_sc_lp__a31o_lp  VNB VPB B1 A1 A2 A3 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 A_116_56# N_B1_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_48_409#_M1005_d N_B1_M1005_g A_116_56# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1009 A_274_56# N_A1_M1009_g N_A_48_409#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1010 A_352_56# N_A2_M1010_g A_274_56# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A3_M1011_g A_352_56# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.8 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1001 A_516_56# N_A_48_409#_M1001_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_48_409#_M1002_g A_516_56# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_155_409#_M1003_d N_B1_M1003_g N_A_48_409#_M1003_s VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_155_409#_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1004 N_A_155_409#_M1004_d N_A2_M1004_g N_VPWR_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_A3_M1000_g N_A_155_409#_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_X_M1006_d N_A_48_409#_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a31o_lp.pxi.spice"
*
.ends
*
*
