* File: sky130_fd_sc_lp__clkinv_4.spice
* Created: Fri Aug 28 10:18:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkinv_4.pex.spice"
.subckt sky130_fd_sc_lp__clkinv_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.5 A=0.063
+ P=1.14 MULT=1
MM1004 N_Y_M1000_d N_A_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.1 A=0.063
+ P=1.14 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1008 N_Y_M1007_d N_A_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3402 AS=0.1764 PD=3.06 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1002_d N_A_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1005_d N_A_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__clkinv_4.pxi.spice"
*
.ends
*
*
