* File: sky130_fd_sc_lp__ha_2.pxi.spice
* Created: Fri Aug 28 10:36:21 2020
* 
x_PM_SKY130_FD_SC_LP__HA_2%A_270_95# N_A_270_95#_M1004_s N_A_270_95#_M1014_d
+ N_A_270_95#_c_102_n N_A_270_95#_M1011_g N_A_270_95#_c_103_n
+ N_A_270_95#_M1003_g N_A_270_95#_M1005_g N_A_270_95#_M1008_g
+ N_A_270_95#_c_106_n N_A_270_95#_c_107_n N_A_270_95#_M1015_g
+ N_A_270_95#_M1016_g N_A_270_95#_c_109_n N_A_270_95#_c_110_n
+ N_A_270_95#_c_111_n N_A_270_95#_c_112_n N_A_270_95#_c_113_n
+ N_A_270_95#_c_114_n N_A_270_95#_c_115_n N_A_270_95#_c_116_n
+ PM_SKY130_FD_SC_LP__HA_2%A_270_95#
x_PM_SKY130_FD_SC_LP__HA_2%B N_B_M1009_g N_B_M1006_g N_B_c_214_n N_B_c_215_n
+ N_B_M1014_g N_B_M1004_g N_B_c_217_n N_B_c_223_n B N_B_c_219_n N_B_c_220_n
+ PM_SKY130_FD_SC_LP__HA_2%B
x_PM_SKY130_FD_SC_LP__HA_2%A N_A_M1010_g N_A_M1013_g N_A_c_294_n N_A_c_295_n
+ N_A_M1001_g N_A_M1007_g N_A_c_298_n A A N_A_c_292_n PM_SKY130_FD_SC_LP__HA_2%A
x_PM_SKY130_FD_SC_LP__HA_2%A_227_397# N_A_227_397#_M1011_d N_A_227_397#_M1006_d
+ N_A_227_397#_M1002_g N_A_227_397#_c_357_n N_A_227_397#_M1000_g
+ N_A_227_397#_M1017_g N_A_227_397#_M1012_g N_A_227_397#_c_360_n
+ N_A_227_397#_c_367_n N_A_227_397#_c_368_n N_A_227_397#_c_369_n
+ N_A_227_397#_c_370_n N_A_227_397#_c_371_n N_A_227_397#_c_361_n
+ N_A_227_397#_c_373_n N_A_227_397#_c_362_n N_A_227_397#_c_363_n
+ N_A_227_397#_c_364_n PM_SKY130_FD_SC_LP__HA_2%A_227_397#
x_PM_SKY130_FD_SC_LP__HA_2%VPWR N_VPWR_M1013_s N_VPWR_M1003_d N_VPWR_M1007_d
+ N_VPWR_M1016_d N_VPWR_M1017_s N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_490_n
+ N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n VPWR
+ N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_487_n
+ PM_SKY130_FD_SC_LP__HA_2%VPWR
x_PM_SKY130_FD_SC_LP__HA_2%COUT N_COUT_M1005_s N_COUT_M1008_s COUT COUT COUT
+ COUT COUT N_COUT_c_570_n COUT PM_SKY130_FD_SC_LP__HA_2%COUT
x_PM_SKY130_FD_SC_LP__HA_2%SUM N_SUM_M1000_s N_SUM_M1002_d SUM SUM SUM SUM SUM
+ SUM SUM N_SUM_c_586_n SUM N_SUM_c_600_n PM_SKY130_FD_SC_LP__HA_2%SUM
x_PM_SKY130_FD_SC_LP__HA_2%A_45_121# N_A_45_121#_M1010_s N_A_45_121#_M1009_d
+ N_A_45_121#_c_609_n N_A_45_121#_c_610_n N_A_45_121#_c_611_n
+ N_A_45_121#_c_612_n PM_SKY130_FD_SC_LP__HA_2%A_45_121#
x_PM_SKY130_FD_SC_LP__HA_2%VGND N_VGND_M1010_d N_VGND_M1001_d N_VGND_M1015_d
+ N_VGND_M1012_d N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n
+ N_VGND_c_640_n VGND N_VGND_c_641_n N_VGND_c_642_n N_VGND_c_643_n
+ N_VGND_c_644_n N_VGND_c_645_n N_VGND_c_646_n N_VGND_c_647_n
+ PM_SKY130_FD_SC_LP__HA_2%VGND
cc_1 VNB N_A_270_95#_c_102_n 0.0201087f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.135
cc_2 VNB N_A_270_95#_c_103_n 0.0281079f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.515
cc_3 VNB N_A_270_95#_M1003_g 0.00780571f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=2.305
cc_4 VNB N_A_270_95#_M1008_g 0.00799353f $X=-0.19 $Y=-0.245 $X2=3.33 $Y2=2.465
cc_5 VNB N_A_270_95#_c_106_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=3.685 $Y2=1.26
cc_6 VNB N_A_270_95#_c_107_n 0.0172427f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=1.185
cc_7 VNB N_A_270_95#_M1016_g 0.0148417f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=2.465
cc_8 VNB N_A_270_95#_c_109_n 0.00490964f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=1.26
cc_9 VNB N_A_270_95#_c_110_n 0.00496721f $X=-0.19 $Y=-0.245 $X2=2.17 $Y2=0.865
cc_10 VNB N_A_270_95#_c_111_n 0.0012768f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=2.14
cc_11 VNB N_A_270_95#_c_112_n 0.0197565f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=1.35
cc_12 VNB N_A_270_95#_c_113_n 0.008181f $X=-0.19 $Y=-0.245 $X2=3.195 $Y2=1.35
cc_13 VNB N_A_270_95#_c_114_n 0.0415777f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.35
cc_14 VNB N_A_270_95#_c_115_n 0.0374218f $X=-0.19 $Y=-0.245 $X2=3.217 $Y2=1.26
cc_15 VNB N_A_270_95#_c_116_n 0.0195888f $X=-0.19 $Y=-0.245 $X2=3.217 $Y2=1.185
cc_16 VNB N_B_M1009_g 0.0306172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_c_214_n 0.104774f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=2.305
cc_18 VNB N_B_c_215_n 0.0116608f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=2.305
cc_19 VNB N_B_M1004_g 0.0600144f $X=-0.19 $Y=-0.245 $X2=3.33 $Y2=2.465
cc_20 VNB N_B_c_217_n 0.0130647f $X=-0.19 $Y=-0.245 $X2=3.685 $Y2=1.26
cc_21 VNB B 0.00201576f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=0.655
cc_22 VNB N_B_c_219_n 0.0139487f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=2.465
cc_23 VNB N_B_c_220_n 0.0126303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_M1010_g 0.0491461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_M1001_g 0.0365185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB A 0.014856f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=1.26
cc_27 VNB N_A_c_292_n 0.0170888f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=2.465
cc_28 VNB N_A_227_397#_M1002_g 0.00646792f $X=-0.19 $Y=-0.245 $X2=1.425
+ $Y2=0.815
cc_29 VNB N_A_227_397#_c_357_n 0.0176763f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=2.305
cc_30 VNB N_A_227_397#_M1017_g 0.0106048f $X=-0.19 $Y=-0.245 $X2=3.33 $Y2=0.655
cc_31 VNB N_A_227_397#_M1012_g 0.0352088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_227_397#_c_360_n 0.00434432f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=0.655
cc_33 VNB N_A_227_397#_c_361_n 0.00114328f $X=-0.19 $Y=-0.245 $X2=2.155 $Y2=1.15
cc_34 VNB N_A_227_397#_c_362_n 0.00393996f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=2.14
cc_35 VNB N_A_227_397#_c_363_n 0.00311263f $X=-0.19 $Y=-0.245 $X2=3.195 $Y2=1.35
cc_36 VNB N_A_227_397#_c_364_n 0.0569185f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.332
cc_37 VNB N_VPWR_c_487_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB COUT 0.00367737f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.815
cc_39 VNB N_SUM_c_586_n 0.00637058f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=0.655
cc_40 VNB N_A_45_121#_c_609_n 0.0170921f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.815
cc_41 VNB N_A_45_121#_c_610_n 0.0122165f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=2.305
cc_42 VNB N_A_45_121#_c_611_n 0.0104963f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=2.305
cc_43 VNB N_A_45_121#_c_612_n 6.63884e-19 $X=-0.19 $Y=-0.245 $X2=3.33 $Y2=0.655
cc_44 VNB N_VGND_c_636_n 0.0129217f $X=-0.19 $Y=-0.245 $X2=3.33 $Y2=1.515
cc_45 VNB N_VGND_c_637_n 0.00995736f $X=-0.19 $Y=-0.245 $X2=3.685 $Y2=1.26
cc_46 VNB N_VGND_c_638_n 0.00444917f $X=-0.19 $Y=-0.245 $X2=3.76 $Y2=2.465
cc_47 VNB N_VGND_c_639_n 0.0113226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_640_n 0.0482593f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.35
cc_49 VNB N_VGND_c_641_n 0.0544714f $X=-0.19 $Y=-0.245 $X2=2.17 $Y2=0.865
cc_50 VNB N_VGND_c_642_n 0.0180594f $X=-0.19 $Y=-0.245 $X2=3.195 $Y2=1.35
cc_51 VNB N_VGND_c_643_n 0.0163082f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.35
cc_52 VNB N_VGND_c_644_n 0.0262509f $X=-0.19 $Y=-0.245 $X2=3.217 $Y2=1.185
cc_53 VNB N_VGND_c_645_n 0.00817144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_646_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_647_n 0.290673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VPB N_A_270_95#_M1003_g 0.0297576f $X=-0.19 $Y=1.655 $X2=1.6 $Y2=2.305
cc_57 VPB N_A_270_95#_M1008_g 0.0220047f $X=-0.19 $Y=1.655 $X2=3.33 $Y2=2.465
cc_58 VPB N_A_270_95#_M1016_g 0.0191092f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=2.465
cc_59 VPB N_A_270_95#_c_111_n 0.00300547f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=2.14
cc_60 VPB N_B_M1006_g 0.0184954f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.815
cc_61 VPB N_B_M1004_g 0.00399941f $X=-0.19 $Y=1.655 $X2=3.33 $Y2=2.465
cc_62 VPB N_B_c_223_n 0.026006f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=1.185
cc_63 VPB B 0.0017222f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=0.655
cc_64 VPB N_B_c_219_n 0.0141846f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=2.465
cc_65 VPB N_A_M1013_g 0.0421941f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.815
cc_66 VPB N_A_c_294_n 0.160333f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.815
cc_67 VPB N_A_c_295_n 0.011606f $X=-0.19 $Y=1.655 $X2=1.6 $Y2=1.515
cc_68 VPB N_A_M1001_g 0.00349088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_M1007_g 0.0338216f $X=-0.19 $Y=1.655 $X2=3.33 $Y2=2.465
cc_70 VPB N_A_c_298_n 0.0118538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB A 0.0179672f $X=-0.19 $Y=1.655 $X2=3.405 $Y2=1.26
cc_72 VPB N_A_c_292_n 0.0243247f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=2.465
cc_73 VPB N_A_227_397#_M1002_g 0.0188175f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.815
cc_74 VPB N_A_227_397#_M1017_g 0.0264982f $X=-0.19 $Y=1.655 $X2=3.33 $Y2=0.655
cc_75 VPB N_A_227_397#_c_367_n 0.0188963f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=1.335
cc_76 VPB N_A_227_397#_c_368_n 0.00726875f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=2.465
cc_77 VPB N_A_227_397#_c_369_n 0.00120689f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_227_397#_c_370_n 0.00423343f $X=-0.19 $Y=1.655 $X2=1.525 $Y2=1.35
cc_79 VPB N_A_227_397#_c_371_n 0.00140781f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.35
cc_80 VPB N_A_227_397#_c_361_n 0.00119828f $X=-0.19 $Y=1.655 $X2=2.155 $Y2=1.15
cc_81 VPB N_A_227_397#_c_373_n 0.00251952f $X=-0.19 $Y=1.655 $X2=2.17 $Y2=0.865
cc_82 VPB N_VPWR_c_488_n 0.0504022f $X=-0.19 $Y=1.655 $X2=3.33 $Y2=2.465
cc_83 VPB N_VPWR_c_489_n 0.0235727f $X=-0.19 $Y=1.655 $X2=3.405 $Y2=1.26
cc_84 VPB N_VPWR_c_490_n 0.00631261f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=1.335
cc_85 VPB N_VPWR_c_491_n 3.3184e-19 $X=-0.19 $Y=1.655 $X2=1.525 $Y2=1.35
cc_86 VPB N_VPWR_c_492_n 0.0144718f $X=-0.19 $Y=1.655 $X2=3.76 $Y2=1.26
cc_87 VPB N_VPWR_c_493_n 0.012416f $X=-0.19 $Y=1.655 $X2=2.155 $Y2=0.865
cc_88 VPB N_VPWR_c_494_n 0.0123263f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=2.14
cc_89 VPB N_VPWR_c_495_n 0.005715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_496_n 0.0337568f $X=-0.19 $Y=1.655 $X2=3.195 $Y2=1.35
cc_91 VPB N_VPWR_c_497_n 0.00347341f $X=-0.19 $Y=1.655 $X2=3.195 $Y2=1.35
cc_92 VPB N_VPWR_c_498_n 0.0125849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_499_n 0.00436447f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.332
cc_94 VPB N_VPWR_c_500_n 0.0266517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_501_n 0.0170875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_502_n 0.0051042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_487_n 0.0600807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB COUT 0.00206673f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.815
cc_99 VPB SUM 0.00439502f $X=-0.19 $Y=1.655 $X2=1.6 $Y2=1.515
cc_100 VPB N_SUM_c_586_n 2.96492e-19 $X=-0.19 $Y=1.655 $X2=3.76 $Y2=0.655
cc_101 N_A_270_95#_c_102_n N_B_M1009_g 0.0112482f $X=1.425 $Y=1.135 $X2=0 $Y2=0
cc_102 N_A_270_95#_M1003_g N_B_M1006_g 0.0160784f $X=1.6 $Y=2.305 $X2=0 $Y2=0
cc_103 N_A_270_95#_c_102_n N_B_c_214_n 0.0103769f $X=1.425 $Y=1.135 $X2=0 $Y2=0
cc_104 N_A_270_95#_c_110_n N_B_c_214_n 0.00454685f $X=2.17 $Y=0.865 $X2=0 $Y2=0
cc_105 N_A_270_95#_c_103_n N_B_M1004_g 6.01102e-19 $X=1.6 $Y=1.515 $X2=0 $Y2=0
cc_106 N_A_270_95#_M1003_g N_B_M1004_g 0.0037214f $X=1.6 $Y=2.305 $X2=0 $Y2=0
cc_107 N_A_270_95#_c_110_n N_B_M1004_g 0.00970681f $X=2.17 $Y=0.865 $X2=0 $Y2=0
cc_108 N_A_270_95#_c_111_n N_B_M1004_g 0.00519652f $X=2.59 $Y=2.14 $X2=0 $Y2=0
cc_109 N_A_270_95#_c_112_n N_B_M1004_g 0.0241191f $X=2.695 $Y=1.35 $X2=0 $Y2=0
cc_110 N_A_270_95#_c_114_n N_B_M1004_g 0.0213949f $X=1.935 $Y=1.35 $X2=0 $Y2=0
cc_111 N_A_270_95#_c_103_n N_B_c_217_n 0.009865f $X=1.6 $Y=1.515 $X2=0 $Y2=0
cc_112 N_A_270_95#_M1003_g N_B_c_223_n 0.0122988f $X=1.6 $Y=2.305 $X2=0 $Y2=0
cc_113 N_A_270_95#_c_111_n N_B_c_223_n 7.6948e-19 $X=2.59 $Y=2.14 $X2=0 $Y2=0
cc_114 N_A_270_95#_c_103_n B 3.48341e-19 $X=1.6 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A_270_95#_c_103_n N_B_c_219_n 0.0212285f $X=1.6 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A_270_95#_c_103_n N_B_c_220_n 0.00574288f $X=1.6 $Y=1.515 $X2=0 $Y2=0
cc_117 N_A_270_95#_M1003_g N_A_c_294_n 0.00921615f $X=1.6 $Y=2.305 $X2=0 $Y2=0
cc_118 N_A_270_95#_M1008_g N_A_M1001_g 0.00512047f $X=3.33 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_270_95#_c_110_n N_A_M1001_g 0.00152985f $X=2.17 $Y=0.865 $X2=0 $Y2=0
cc_120 N_A_270_95#_c_111_n N_A_M1001_g 0.00530765f $X=2.59 $Y=2.14 $X2=0 $Y2=0
cc_121 N_A_270_95#_c_112_n N_A_M1001_g 0.00515565f $X=2.695 $Y=1.35 $X2=0 $Y2=0
cc_122 N_A_270_95#_c_113_n N_A_M1001_g 0.0174985f $X=3.195 $Y=1.35 $X2=0 $Y2=0
cc_123 N_A_270_95#_c_115_n N_A_M1001_g 0.0213869f $X=3.217 $Y=1.26 $X2=0 $Y2=0
cc_124 N_A_270_95#_c_116_n N_A_M1001_g 0.0100167f $X=3.217 $Y=1.185 $X2=0 $Y2=0
cc_125 N_A_270_95#_c_111_n N_A_M1007_g 0.00272551f $X=2.59 $Y=2.14 $X2=0 $Y2=0
cc_126 N_A_270_95#_M1008_g N_A_c_298_n 0.0392122f $X=3.33 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_270_95#_c_111_n N_A_c_298_n 0.00440004f $X=2.59 $Y=2.14 $X2=0 $Y2=0
cc_128 N_A_270_95#_c_113_n N_A_c_298_n 0.00254969f $X=3.195 $Y=1.35 $X2=0 $Y2=0
cc_129 N_A_270_95#_M1016_g N_A_227_397#_M1002_g 0.0559165f $X=3.76 $Y=2.465
+ $X2=0 $Y2=0
cc_130 N_A_270_95#_c_107_n N_A_227_397#_c_357_n 0.0221802f $X=3.76 $Y=1.185
+ $X2=0 $Y2=0
cc_131 N_A_270_95#_c_102_n N_A_227_397#_c_360_n 0.00361963f $X=1.425 $Y=1.135
+ $X2=0 $Y2=0
cc_132 N_A_270_95#_c_103_n N_A_227_397#_c_360_n 0.0175487f $X=1.6 $Y=1.515 $X2=0
+ $Y2=0
cc_133 N_A_270_95#_M1003_g N_A_227_397#_c_360_n 0.00549973f $X=1.6 $Y=2.305
+ $X2=0 $Y2=0
cc_134 N_A_270_95#_c_110_n N_A_227_397#_c_360_n 0.00869479f $X=2.17 $Y=0.865
+ $X2=0 $Y2=0
cc_135 N_A_270_95#_c_112_n N_A_227_397#_c_360_n 0.0266903f $X=2.695 $Y=1.35
+ $X2=0 $Y2=0
cc_136 N_A_270_95#_c_103_n N_A_227_397#_c_367_n 0.00618152f $X=1.6 $Y=1.515
+ $X2=0 $Y2=0
cc_137 N_A_270_95#_M1003_g N_A_227_397#_c_367_n 0.00474315f $X=1.6 $Y=2.305
+ $X2=0 $Y2=0
cc_138 N_A_270_95#_c_111_n N_A_227_397#_c_367_n 0.0136513f $X=2.59 $Y=2.14 $X2=0
+ $Y2=0
cc_139 N_A_270_95#_c_112_n N_A_227_397#_c_367_n 0.0414188f $X=2.695 $Y=1.35
+ $X2=0 $Y2=0
cc_140 N_A_270_95#_c_114_n N_A_227_397#_c_367_n 0.00183286f $X=1.935 $Y=1.35
+ $X2=0 $Y2=0
cc_141 N_A_270_95#_c_103_n N_A_227_397#_c_368_n 0.00347326f $X=1.6 $Y=1.515
+ $X2=0 $Y2=0
cc_142 N_A_270_95#_M1003_g N_A_227_397#_c_368_n 0.01954f $X=1.6 $Y=2.305 $X2=0
+ $Y2=0
cc_143 N_A_270_95#_M1003_g N_A_227_397#_c_369_n 0.00417356f $X=1.6 $Y=2.305
+ $X2=0 $Y2=0
cc_144 N_A_270_95#_c_111_n N_A_227_397#_c_369_n 0.0201191f $X=2.59 $Y=2.14 $X2=0
+ $Y2=0
cc_145 N_A_270_95#_M1014_d N_A_227_397#_c_370_n 0.00173272f $X=2.45 $Y=1.985
+ $X2=0 $Y2=0
cc_146 N_A_270_95#_M1008_g N_A_227_397#_c_370_n 0.0168313f $X=3.33 $Y=2.465
+ $X2=0 $Y2=0
cc_147 N_A_270_95#_M1016_g N_A_227_397#_c_370_n 0.0151399f $X=3.76 $Y=2.465
+ $X2=0 $Y2=0
cc_148 N_A_270_95#_c_111_n N_A_227_397#_c_370_n 0.0135055f $X=2.59 $Y=2.14 $X2=0
+ $Y2=0
cc_149 N_A_270_95#_M1016_g N_A_227_397#_c_361_n 0.00907112f $X=3.76 $Y=2.465
+ $X2=0 $Y2=0
cc_150 N_A_270_95#_M1003_g N_A_227_397#_c_373_n 0.0068898f $X=1.6 $Y=2.305 $X2=0
+ $Y2=0
cc_151 N_A_270_95#_c_102_n N_A_227_397#_c_362_n 0.00331519f $X=1.425 $Y=1.135
+ $X2=0 $Y2=0
cc_152 N_A_270_95#_c_103_n N_A_227_397#_c_362_n 8.86691e-19 $X=1.6 $Y=1.515
+ $X2=0 $Y2=0
cc_153 N_A_270_95#_c_110_n N_A_227_397#_c_362_n 0.0234154f $X=2.17 $Y=0.865
+ $X2=0 $Y2=0
cc_154 N_A_270_95#_c_114_n N_A_227_397#_c_362_n 0.00481629f $X=1.935 $Y=1.35
+ $X2=0 $Y2=0
cc_155 N_A_270_95#_c_109_n N_A_227_397#_c_363_n 0.00233017f $X=3.76 $Y=1.26
+ $X2=0 $Y2=0
cc_156 N_A_270_95#_c_109_n N_A_227_397#_c_364_n 0.0205281f $X=3.76 $Y=1.26 $X2=0
+ $Y2=0
cc_157 N_A_270_95#_M1003_g N_VPWR_c_489_n 0.0081537f $X=1.6 $Y=2.305 $X2=0 $Y2=0
cc_158 N_A_270_95#_M1008_g N_VPWR_c_490_n 0.00953757f $X=3.33 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A_270_95#_M1016_g N_VPWR_c_490_n 0.00125151f $X=3.76 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_270_95#_M1008_g N_VPWR_c_491_n 0.00125151f $X=3.33 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_270_95#_M1016_g N_VPWR_c_491_n 0.00881515f $X=3.76 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_270_95#_M1008_g N_VPWR_c_498_n 0.00359504f $X=3.33 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_270_95#_M1016_g N_VPWR_c_498_n 0.00359504f $X=3.76 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_270_95#_M1003_g N_VPWR_c_487_n 8.61222e-19 $X=1.6 $Y=2.305 $X2=0
+ $Y2=0
cc_165 N_A_270_95#_M1008_g N_VPWR_c_487_n 0.00429447f $X=3.33 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_270_95#_M1016_g N_VPWR_c_487_n 0.00429447f $X=3.76 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_270_95#_c_106_n COUT 0.0101253f $X=3.685 $Y=1.26 $X2=0 $Y2=0
cc_168 N_A_270_95#_c_107_n COUT 0.00487703f $X=3.76 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A_270_95#_M1016_g COUT 0.0186409f $X=3.76 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_270_95#_c_109_n COUT 0.00190249f $X=3.76 $Y=1.26 $X2=0 $Y2=0
cc_171 N_A_270_95#_c_113_n COUT 0.0265543f $X=3.195 $Y=1.35 $X2=0 $Y2=0
cc_172 N_A_270_95#_c_115_n COUT 0.0104658f $X=3.217 $Y=1.26 $X2=0 $Y2=0
cc_173 N_A_270_95#_c_116_n COUT 0.0030173f $X=3.217 $Y=1.185 $X2=0 $Y2=0
cc_174 N_A_270_95#_c_107_n N_COUT_c_570_n 0.00752715f $X=3.76 $Y=1.185 $X2=0
+ $Y2=0
cc_175 N_A_270_95#_c_116_n N_COUT_c_570_n 0.00638868f $X=3.217 $Y=1.185 $X2=0
+ $Y2=0
cc_176 N_A_270_95#_c_107_n COUT 0.00189571f $X=3.76 $Y=1.185 $X2=0 $Y2=0
cc_177 N_A_270_95#_c_116_n COUT 0.00228561f $X=3.217 $Y=1.185 $X2=0 $Y2=0
cc_178 N_A_270_95#_c_102_n N_A_45_121#_c_610_n 0.00143946f $X=1.425 $Y=1.135
+ $X2=0 $Y2=0
cc_179 N_A_270_95#_c_102_n N_A_45_121#_c_612_n 4.31322e-19 $X=1.425 $Y=1.135
+ $X2=0 $Y2=0
cc_180 N_A_270_95#_c_102_n N_VGND_c_636_n 8.47936e-19 $X=1.425 $Y=1.135 $X2=0
+ $Y2=0
cc_181 N_A_270_95#_c_110_n N_VGND_c_637_n 0.0108177f $X=2.17 $Y=0.865 $X2=0
+ $Y2=0
cc_182 N_A_270_95#_c_113_n N_VGND_c_637_n 0.0321857f $X=3.195 $Y=1.35 $X2=0
+ $Y2=0
cc_183 N_A_270_95#_c_115_n N_VGND_c_637_n 0.00433889f $X=3.217 $Y=1.26 $X2=0
+ $Y2=0
cc_184 N_A_270_95#_c_116_n N_VGND_c_637_n 0.0060935f $X=3.217 $Y=1.185 $X2=0
+ $Y2=0
cc_185 N_A_270_95#_c_107_n N_VGND_c_638_n 0.00906616f $X=3.76 $Y=1.185 $X2=0
+ $Y2=0
cc_186 N_A_270_95#_c_110_n N_VGND_c_641_n 0.00556326f $X=2.17 $Y=0.865 $X2=0
+ $Y2=0
cc_187 N_A_270_95#_c_107_n N_VGND_c_642_n 0.00526178f $X=3.76 $Y=1.185 $X2=0
+ $Y2=0
cc_188 N_A_270_95#_c_116_n N_VGND_c_642_n 0.00564131f $X=3.217 $Y=1.185 $X2=0
+ $Y2=0
cc_189 N_A_270_95#_c_102_n N_VGND_c_647_n 9.27138e-19 $X=1.425 $Y=1.135 $X2=0
+ $Y2=0
cc_190 N_A_270_95#_c_107_n N_VGND_c_647_n 0.00973873f $X=3.76 $Y=1.185 $X2=0
+ $Y2=0
cc_191 N_A_270_95#_c_110_n N_VGND_c_647_n 0.0088989f $X=2.17 $Y=0.865 $X2=0
+ $Y2=0
cc_192 N_A_270_95#_c_116_n N_VGND_c_647_n 0.0114086f $X=3.217 $Y=1.185 $X2=0
+ $Y2=0
cc_193 N_B_M1009_g N_A_M1010_g 0.0206795f $X=0.995 $Y=0.815 $X2=0 $Y2=0
cc_194 N_B_c_220_n N_A_M1010_g 0.00879271f $X=1.15 $Y=1.495 $X2=0 $Y2=0
cc_195 N_B_M1006_g N_A_M1013_g 0.0322233f $X=1.06 $Y=2.305 $X2=0 $Y2=0
cc_196 N_B_M1006_g N_A_c_294_n 0.00909527f $X=1.06 $Y=2.305 $X2=0 $Y2=0
cc_197 N_B_c_223_n N_A_c_294_n 0.00844658f $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_198 N_B_M1004_g N_A_M1001_g 0.0405739f $X=2.385 $Y=0.865 $X2=0 $Y2=0
cc_199 N_B_c_223_n N_A_M1007_g 0.0234305f $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_200 N_B_c_223_n N_A_c_298_n 0.0405739f $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_201 B A 0.0252539f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_202 N_B_c_219_n A 0.00130829f $X=1.15 $Y=1.66 $X2=0 $Y2=0
cc_203 B N_A_c_292_n 3.1873e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_204 N_B_c_219_n N_A_c_292_n 0.039556f $X=1.15 $Y=1.66 $X2=0 $Y2=0
cc_205 N_B_M1004_g N_A_227_397#_c_360_n 0.00135792f $X=2.385 $Y=0.865 $X2=0
+ $Y2=0
cc_206 N_B_c_217_n N_A_227_397#_c_360_n 2.87394e-19 $X=1.03 $Y=1.285 $X2=0 $Y2=0
cc_207 B N_A_227_397#_c_360_n 0.0142682f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_208 N_B_c_219_n N_A_227_397#_c_360_n 5.53018e-19 $X=1.15 $Y=1.66 $X2=0 $Y2=0
cc_209 N_B_c_220_n N_A_227_397#_c_360_n 0.00371265f $X=1.15 $Y=1.495 $X2=0 $Y2=0
cc_210 N_B_M1004_g N_A_227_397#_c_367_n 0.00152906f $X=2.385 $Y=0.865 $X2=0
+ $Y2=0
cc_211 N_B_c_223_n N_A_227_397#_c_367_n 0.00414705f $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_212 N_B_M1006_g N_A_227_397#_c_368_n 0.00599967f $X=1.06 $Y=2.305 $X2=0 $Y2=0
cc_213 N_B_c_223_n N_A_227_397#_c_368_n 2.6931e-19 $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_214 B N_A_227_397#_c_368_n 0.0262792f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_215 N_B_c_219_n N_A_227_397#_c_368_n 0.0054717f $X=1.15 $Y=1.66 $X2=0 $Y2=0
cc_216 N_B_c_223_n N_A_227_397#_c_369_n 0.015818f $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_217 N_B_c_223_n N_A_227_397#_c_370_n 0.0105295f $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_218 N_B_c_223_n N_A_227_397#_c_371_n 0.00325715f $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_219 N_B_M1006_g N_A_227_397#_c_373_n 0.00842377f $X=1.06 $Y=2.305 $X2=0 $Y2=0
cc_220 N_B_c_214_n N_A_227_397#_c_362_n 0.00545514f $X=2.31 $Y=0.19 $X2=0 $Y2=0
cc_221 N_B_M1004_g N_A_227_397#_c_362_n 9.43793e-19 $X=2.385 $Y=0.865 $X2=0
+ $Y2=0
cc_222 N_B_M1006_g N_VPWR_c_488_n 0.00239803f $X=1.06 $Y=2.305 $X2=0 $Y2=0
cc_223 N_B_c_223_n N_VPWR_c_489_n 0.00347834f $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_224 N_B_M1006_g N_VPWR_c_487_n 8.61222e-19 $X=1.06 $Y=2.305 $X2=0 $Y2=0
cc_225 N_B_c_223_n N_VPWR_c_487_n 8.61222e-19 $X=2.38 $Y=1.875 $X2=0 $Y2=0
cc_226 N_B_M1009_g N_A_45_121#_c_609_n 4.47146e-19 $X=0.995 $Y=0.815 $X2=0 $Y2=0
cc_227 N_B_M1009_g N_A_45_121#_c_610_n 0.00825064f $X=0.995 $Y=0.815 $X2=0 $Y2=0
cc_228 N_B_c_217_n N_A_45_121#_c_610_n 0.0105057f $X=1.03 $Y=1.285 $X2=0 $Y2=0
cc_229 B N_A_45_121#_c_610_n 0.0191142f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_230 N_B_c_219_n N_A_45_121#_c_610_n 0.00387498f $X=1.15 $Y=1.66 $X2=0 $Y2=0
cc_231 N_B_M1009_g N_A_45_121#_c_612_n 7.0559e-19 $X=0.995 $Y=0.815 $X2=0 $Y2=0
cc_232 N_B_c_214_n N_A_45_121#_c_612_n 0.00282931f $X=2.31 $Y=0.19 $X2=0 $Y2=0
cc_233 N_B_M1009_g N_VGND_c_636_n 0.0193786f $X=0.995 $Y=0.815 $X2=0 $Y2=0
cc_234 N_B_c_215_n N_VGND_c_636_n 0.00735148f $X=1.07 $Y=0.19 $X2=0 $Y2=0
cc_235 N_B_c_214_n N_VGND_c_637_n 0.0121759f $X=2.31 $Y=0.19 $X2=0 $Y2=0
cc_236 N_B_M1004_g N_VGND_c_637_n 0.00172994f $X=2.385 $Y=0.865 $X2=0 $Y2=0
cc_237 N_B_c_215_n N_VGND_c_641_n 0.0454834f $X=1.07 $Y=0.19 $X2=0 $Y2=0
cc_238 N_B_c_214_n N_VGND_c_647_n 0.0524118f $X=2.31 $Y=0.19 $X2=0 $Y2=0
cc_239 N_B_c_215_n N_VGND_c_647_n 0.00812742f $X=1.07 $Y=0.19 $X2=0 $Y2=0
cc_240 N_A_M1013_g N_A_227_397#_c_368_n 4.84343e-19 $X=0.7 $Y=2.305 $X2=0 $Y2=0
cc_241 A N_A_227_397#_c_368_n 3.51358e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_242 N_A_M1007_g N_A_227_397#_c_369_n 9.10659e-19 $X=2.805 $Y=2.305 $X2=0
+ $Y2=0
cc_243 N_A_c_294_n N_A_227_397#_c_370_n 0.00390741f $X=2.73 $Y=3.07 $X2=0 $Y2=0
cc_244 N_A_M1007_g N_A_227_397#_c_370_n 0.0169731f $X=2.805 $Y=2.305 $X2=0 $Y2=0
cc_245 N_A_c_294_n N_A_227_397#_c_371_n 0.00288504f $X=2.73 $Y=3.07 $X2=0 $Y2=0
cc_246 N_A_M1013_g N_A_227_397#_c_373_n 0.00136182f $X=0.7 $Y=2.305 $X2=0 $Y2=0
cc_247 N_A_c_294_n N_A_227_397#_c_373_n 0.00523019f $X=2.73 $Y=3.07 $X2=0 $Y2=0
cc_248 N_A_M1013_g N_VPWR_c_488_n 0.0309315f $X=0.7 $Y=2.305 $X2=0 $Y2=0
cc_249 N_A_c_295_n N_VPWR_c_488_n 0.00957316f $X=0.775 $Y=3.07 $X2=0 $Y2=0
cc_250 A N_VPWR_c_488_n 0.0275533f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_251 N_A_c_292_n N_VPWR_c_488_n 0.00710657f $X=0.565 $Y=1.66 $X2=0 $Y2=0
cc_252 N_A_c_294_n N_VPWR_c_489_n 0.0233862f $X=2.73 $Y=3.07 $X2=0 $Y2=0
cc_253 N_A_M1007_g N_VPWR_c_490_n 0.0090836f $X=2.805 $Y=2.305 $X2=0 $Y2=0
cc_254 N_A_c_295_n N_VPWR_c_496_n 0.0327282f $X=0.775 $Y=3.07 $X2=0 $Y2=0
cc_255 N_A_c_294_n N_VPWR_c_500_n 0.0212347f $X=2.73 $Y=3.07 $X2=0 $Y2=0
cc_256 N_A_c_294_n N_VPWR_c_487_n 0.0727173f $X=2.73 $Y=3.07 $X2=0 $Y2=0
cc_257 N_A_c_295_n N_VPWR_c_487_n 0.00757253f $X=0.775 $Y=3.07 $X2=0 $Y2=0
cc_258 N_A_M1010_g N_A_45_121#_c_609_n 0.00740567f $X=0.565 $Y=0.815 $X2=0 $Y2=0
cc_259 N_A_M1010_g N_A_45_121#_c_610_n 0.0112726f $X=0.565 $Y=0.815 $X2=0 $Y2=0
cc_260 A N_A_45_121#_c_610_n 0.0168856f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_261 N_A_c_292_n N_A_45_121#_c_610_n 0.00141812f $X=0.565 $Y=1.66 $X2=0 $Y2=0
cc_262 N_A_M1010_g N_A_45_121#_c_611_n 0.00426039f $X=0.565 $Y=0.815 $X2=0 $Y2=0
cc_263 A N_A_45_121#_c_611_n 0.0211374f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_264 N_A_c_292_n N_A_45_121#_c_611_n 0.00309986f $X=0.565 $Y=1.66 $X2=0 $Y2=0
cc_265 N_A_M1010_g N_VGND_c_636_n 0.0033606f $X=0.565 $Y=0.815 $X2=0 $Y2=0
cc_266 N_A_M1001_g N_VGND_c_637_n 0.0114868f $X=2.745 $Y=0.865 $X2=0 $Y2=0
cc_267 N_A_M1001_g N_VGND_c_641_n 0.00332367f $X=2.745 $Y=0.865 $X2=0 $Y2=0
cc_268 N_A_M1010_g N_VGND_c_644_n 0.00410613f $X=0.565 $Y=0.815 $X2=0 $Y2=0
cc_269 N_A_M1010_g N_VGND_c_647_n 0.00474994f $X=0.565 $Y=0.815 $X2=0 $Y2=0
cc_270 N_A_M1001_g N_VGND_c_647_n 0.00387424f $X=2.745 $Y=0.865 $X2=0 $Y2=0
cc_271 N_A_227_397#_c_369_n N_VPWR_M1003_d 0.00601967f $X=2.25 $Y=2.475 $X2=0
+ $Y2=0
cc_272 N_A_227_397#_c_371_n N_VPWR_M1003_d 0.00147391f $X=2.335 $Y=2.56 $X2=0
+ $Y2=0
cc_273 N_A_227_397#_c_370_n N_VPWR_M1007_d 0.0122418f $X=3.97 $Y=2.56 $X2=0
+ $Y2=0
cc_274 N_A_227_397#_c_370_n N_VPWR_M1016_d 0.0046649f $X=3.97 $Y=2.56 $X2=0
+ $Y2=0
cc_275 N_A_227_397#_c_361_n N_VPWR_M1016_d 0.00641385f $X=4.055 $Y=2.475 $X2=0
+ $Y2=0
cc_276 N_A_227_397#_c_368_n N_VPWR_c_488_n 0.0055786f $X=1.66 $Y=1.77 $X2=0
+ $Y2=0
cc_277 N_A_227_397#_c_373_n N_VPWR_c_488_n 0.0165045f $X=1.275 $Y=2.13 $X2=0
+ $Y2=0
cc_278 N_A_227_397#_c_367_n N_VPWR_c_489_n 0.00952809f $X=2.165 $Y=1.77 $X2=0
+ $Y2=0
cc_279 N_A_227_397#_c_369_n N_VPWR_c_489_n 0.0162292f $X=2.25 $Y=2.475 $X2=0
+ $Y2=0
cc_280 N_A_227_397#_c_371_n N_VPWR_c_489_n 0.0141163f $X=2.335 $Y=2.56 $X2=0
+ $Y2=0
cc_281 N_A_227_397#_c_373_n N_VPWR_c_489_n 0.015838f $X=1.275 $Y=2.13 $X2=0
+ $Y2=0
cc_282 N_A_227_397#_c_370_n N_VPWR_c_490_n 0.020926f $X=3.97 $Y=2.56 $X2=0 $Y2=0
cc_283 N_A_227_397#_M1002_g N_VPWR_c_491_n 0.00721913f $X=4.19 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_A_227_397#_M1017_g N_VPWR_c_491_n 5.06813e-19 $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_285 N_A_227_397#_c_370_n N_VPWR_c_491_n 0.0170655f $X=3.97 $Y=2.56 $X2=0
+ $Y2=0
cc_286 N_A_227_397#_M1017_g N_VPWR_c_493_n 0.0288816f $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_A_227_397#_c_364_n N_VPWR_c_493_n 0.00143173f $X=4.62 $Y=1.365 $X2=0
+ $Y2=0
cc_288 N_A_227_397#_c_373_n N_VPWR_c_496_n 0.00492217f $X=1.275 $Y=2.13 $X2=0
+ $Y2=0
cc_289 N_A_227_397#_c_370_n N_VPWR_c_498_n 0.00721067f $X=3.97 $Y=2.56 $X2=0
+ $Y2=0
cc_290 N_A_227_397#_c_370_n N_VPWR_c_500_n 0.00959651f $X=3.97 $Y=2.56 $X2=0
+ $Y2=0
cc_291 N_A_227_397#_c_371_n N_VPWR_c_500_n 0.00301977f $X=2.335 $Y=2.56 $X2=0
+ $Y2=0
cc_292 N_A_227_397#_M1002_g N_VPWR_c_501_n 0.00486043f $X=4.19 $Y=2.465 $X2=0
+ $Y2=0
cc_293 N_A_227_397#_M1017_g N_VPWR_c_501_n 0.00435091f $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_294 N_A_227_397#_M1002_g N_VPWR_c_487_n 0.00824727f $X=4.19 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_227_397#_M1017_g N_VPWR_c_487_n 0.00839005f $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_227_397#_c_370_n N_VPWR_c_487_n 0.0306348f $X=3.97 $Y=2.56 $X2=0
+ $Y2=0
cc_297 N_A_227_397#_c_371_n N_VPWR_c_487_n 0.00425831f $X=2.335 $Y=2.56 $X2=0
+ $Y2=0
cc_298 N_A_227_397#_c_373_n N_VPWR_c_487_n 0.00695091f $X=1.275 $Y=2.13 $X2=0
+ $Y2=0
cc_299 N_A_227_397#_c_370_n N_COUT_M1008_s 0.00481984f $X=3.97 $Y=2.56 $X2=0
+ $Y2=0
cc_300 N_A_227_397#_M1002_g COUT 7.01132e-19 $X=4.19 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A_227_397#_c_370_n COUT 0.0164342f $X=3.97 $Y=2.56 $X2=0 $Y2=0
cc_302 N_A_227_397#_c_361_n COUT 0.0438875f $X=4.055 $Y=2.475 $X2=0 $Y2=0
cc_303 N_A_227_397#_c_363_n COUT 0.0195264f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_304 N_A_227_397#_c_364_n COUT 3.06502e-19 $X=4.62 $Y=1.365 $X2=0 $Y2=0
cc_305 N_A_227_397#_c_357_n N_COUT_c_570_n 9.3465e-19 $X=4.345 $Y=1.185 $X2=0
+ $Y2=0
cc_306 N_A_227_397#_M1002_g SUM 0.00170727f $X=4.19 $Y=2.465 $X2=0 $Y2=0
cc_307 N_A_227_397#_M1017_g SUM 0.00796673f $X=4.62 $Y=2.465 $X2=0 $Y2=0
cc_308 N_A_227_397#_c_361_n SUM 0.0321967f $X=4.055 $Y=2.475 $X2=0 $Y2=0
cc_309 N_A_227_397#_c_364_n SUM 0.00478658f $X=4.62 $Y=1.365 $X2=0 $Y2=0
cc_310 N_A_227_397#_M1002_g N_SUM_c_586_n 0.0012372f $X=4.19 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A_227_397#_c_357_n N_SUM_c_586_n 0.00475043f $X=4.345 $Y=1.185 $X2=0
+ $Y2=0
cc_312 N_A_227_397#_M1017_g N_SUM_c_586_n 0.0092898f $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_313 N_A_227_397#_M1012_g N_SUM_c_586_n 0.00723964f $X=4.775 $Y=0.655 $X2=0
+ $Y2=0
cc_314 N_A_227_397#_c_361_n N_SUM_c_586_n 0.00794286f $X=4.055 $Y=2.475 $X2=0
+ $Y2=0
cc_315 N_A_227_397#_c_363_n N_SUM_c_586_n 0.0242888f $X=4.21 $Y=1.35 $X2=0 $Y2=0
cc_316 N_A_227_397#_c_364_n N_SUM_c_586_n 0.0129031f $X=4.62 $Y=1.365 $X2=0
+ $Y2=0
cc_317 N_A_227_397#_M1017_g N_SUM_c_600_n 0.0211676f $X=4.62 $Y=2.465 $X2=0
+ $Y2=0
cc_318 N_A_227_397#_c_360_n N_A_45_121#_c_610_n 0.0137056f $X=1.572 $Y=1.685
+ $X2=0 $Y2=0
cc_319 N_A_227_397#_c_362_n N_A_45_121#_c_612_n 0.0173889f $X=1.64 $Y=0.815
+ $X2=0 $Y2=0
cc_320 N_A_227_397#_c_357_n N_VGND_c_638_n 0.00660626f $X=4.345 $Y=1.185 $X2=0
+ $Y2=0
cc_321 N_A_227_397#_c_363_n N_VGND_c_638_n 0.0207901f $X=4.21 $Y=1.35 $X2=0
+ $Y2=0
cc_322 N_A_227_397#_c_364_n N_VGND_c_638_n 0.00456632f $X=4.62 $Y=1.365 $X2=0
+ $Y2=0
cc_323 N_A_227_397#_c_357_n N_VGND_c_640_n 7.28716e-19 $X=4.345 $Y=1.185 $X2=0
+ $Y2=0
cc_324 N_A_227_397#_M1012_g N_VGND_c_640_n 0.0186714f $X=4.775 $Y=0.655 $X2=0
+ $Y2=0
cc_325 N_A_227_397#_c_362_n N_VGND_c_641_n 0.00527734f $X=1.64 $Y=0.815 $X2=0
+ $Y2=0
cc_326 N_A_227_397#_c_357_n N_VGND_c_643_n 0.00585385f $X=4.345 $Y=1.185 $X2=0
+ $Y2=0
cc_327 N_A_227_397#_M1012_g N_VGND_c_643_n 0.00486043f $X=4.775 $Y=0.655 $X2=0
+ $Y2=0
cc_328 N_A_227_397#_c_357_n N_VGND_c_647_n 0.011106f $X=4.345 $Y=1.185 $X2=0
+ $Y2=0
cc_329 N_A_227_397#_M1012_g N_VGND_c_647_n 0.00824727f $X=4.775 $Y=0.655 $X2=0
+ $Y2=0
cc_330 N_A_227_397#_c_362_n N_VGND_c_647_n 0.00812674f $X=1.64 $Y=0.815 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_487_n N_COUT_M1008_s 0.00346035f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_332 N_VPWR_c_487_n N_SUM_M1002_d 0.00380103f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_333 N_VPWR_c_493_n SUM 0.0942617f $X=4.9 $Y=1.98 $X2=0 $Y2=0
cc_334 N_VPWR_c_501_n N_SUM_c_600_n 0.020801f $X=4.815 $Y=3.33 $X2=0 $Y2=0
cc_335 N_VPWR_c_487_n N_SUM_c_600_n 0.0124201f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_336 N_COUT_c_570_n N_VGND_c_638_n 0.0590227f $X=3.545 $Y=0.42 $X2=0 $Y2=0
cc_337 N_COUT_c_570_n N_VGND_c_642_n 0.0192645f $X=3.545 $Y=0.42 $X2=0 $Y2=0
cc_338 N_COUT_M1005_s N_VGND_c_647_n 0.00223559f $X=3.405 $Y=0.235 $X2=0 $Y2=0
cc_339 N_COUT_c_570_n N_VGND_c_647_n 0.0125574f $X=3.545 $Y=0.42 $X2=0 $Y2=0
cc_340 N_SUM_c_586_n N_VGND_c_640_n 0.0307993f $X=4.56 $Y=0.42 $X2=0 $Y2=0
cc_341 N_SUM_c_586_n N_VGND_c_643_n 0.0120977f $X=4.56 $Y=0.42 $X2=0 $Y2=0
cc_342 N_SUM_M1000_s N_VGND_c_647_n 0.00571434f $X=4.42 $Y=0.235 $X2=0 $Y2=0
cc_343 N_SUM_c_586_n N_VGND_c_647_n 0.00691495f $X=4.56 $Y=0.42 $X2=0 $Y2=0
cc_344 N_A_45_121#_c_610_n N_VGND_c_636_n 0.0173217f $X=1.105 $Y=1.16 $X2=0
+ $Y2=0
cc_345 N_A_45_121#_c_612_n N_VGND_c_641_n 0.00346302f $X=1.21 $Y=0.815 $X2=0
+ $Y2=0
cc_346 N_A_45_121#_c_609_n N_VGND_c_644_n 0.00554479f $X=0.35 $Y=0.815 $X2=0
+ $Y2=0
cc_347 N_A_45_121#_c_609_n N_VGND_c_647_n 0.0097402f $X=0.35 $Y=0.815 $X2=0
+ $Y2=0
cc_348 N_A_45_121#_c_612_n N_VGND_c_647_n 0.0053872f $X=1.21 $Y=0.815 $X2=0
+ $Y2=0
