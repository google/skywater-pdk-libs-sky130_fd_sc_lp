* File: sky130_fd_sc_lp__dfxtp_1.spice
* Created: Wed Sep  2 09:45:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfxtp_1.pex.spice"
.subckt sky130_fd_sc_lp__dfxtp_1  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1002 N_A_110_70#_M1002_d N_CLK_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_110_70#_M1011_g N_A_217_413#_M1011_s VNB NSHORT L=0.15
+ W=0.42 AD=0.10605 AS=0.1113 PD=0.925 PS=1.37 NRD=34.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004 A=0.063 P=1.14 MULT=1
MM1018 N_A_440_413#_M1018_d N_D_M1018_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.10605 PD=0.7 PS=0.925 NRD=0 NRS=30 M=1 R=2.8 SA=75000.8
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1020 N_A_526_413#_M1020_d N_A_110_70#_M1020_g N_A_440_413#_M1018_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.3 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1016 A_626_163# N_A_217_413#_M1016_g N_A_526_413#_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_668_137#_M1008_g A_626_163# VNB NSHORT L=0.15 W=0.42
+ AD=0.182264 AS=0.0441 PD=1.10943 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8
+ SA=75002.1 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1005 N_A_668_137#_M1005_d N_A_526_413#_M1005_g N_VGND_M1008_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.121419 AS=0.277736 PD=1.1834 PS=1.69057 NRD=2.808 NRS=6.552
+ M=1 R=4.26667 SA=75002.1 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1009 N_A_957_379#_M1009_d N_A_217_413#_M1009_g N_A_668_137#_M1005_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1134 AS=0.0796811 PD=0.96 PS=0.776604 NRD=35.712 NRS=13.56
+ M=1 R=2.8 SA=75002.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1017 A_1116_119# N_A_110_70#_M1017_g N_A_957_379#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1134 PD=0.63 PS=0.96 NRD=14.28 NRS=38.568 M=1 R=2.8
+ SA=75002.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_1158_93#_M1013_g A_1116_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0834849 AS=0.0441 PD=0.788491 PS=0.63 NRD=17.856 NRS=14.28 M=1 R=2.8
+ SA=75003.3 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_1158_93#_M1010_d N_A_957_379#_M1010_g N_VGND_M1013_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.2048 AS=0.127215 PD=1.92 PS=1.20151 NRD=10.308 NRS=2.808
+ M=1 R=4.26667 SA=75002.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_Q_M1007_d N_A_1158_93#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_A_110_70#_M1021_d N_CLK_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_A_110_70#_M1012_g N_A_217_413#_M1012_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.174672 AS=0.1696 PD=1.43698 PS=1.81 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1023 N_A_440_413#_M1023_d N_D_M1023_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.114628 PD=0.7 PS=0.943019 NRD=0 NRS=128.976 M=1 R=2.8
+ SA=75000.9 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1004 N_A_526_413#_M1004_d N_A_217_413#_M1004_g N_A_440_413#_M1023_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1155 AS=0.0588 PD=0.97 PS=0.7 NRD=121.943 NRS=0 M=1
+ R=2.8 SA=75001.3 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1019 A_666_413# N_A_110_70#_M1019_g N_A_526_413#_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1155 PD=0.63 PS=0.97 NRD=23.443 NRS=4.6886 M=1 R=2.8
+ SA=75002 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1022_d N_A_668_137#_M1022_g A_666_413# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.117233 AS=0.0441 PD=0.936667 PS=0.63 NRD=105.119 NRS=23.443 M=1 R=2.8
+ SA=75002.4 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_668_137#_M1000_d N_A_526_413#_M1000_g N_VPWR_M1022_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1512 AS=0.234467 PD=1.2 PS=1.87333 NRD=0 NRS=15.2281 M=1
+ R=5.6 SA=75001.6 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1001 N_A_957_379#_M1001_d N_A_110_70#_M1001_g N_A_668_137#_M1000_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.3304 AS=0.1512 PD=1.98 PS=1.2 NRD=63.3158 NRS=18.7544 M=1
+ R=5.6 SA=75002.1 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1003 A_1116_379# N_A_217_413#_M1003_g N_A_957_379#_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1652 PD=0.63 PS=0.99 NRD=23.443 NRS=44.5417 M=1 R=2.8
+ SA=75003.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_1158_93#_M1006_g A_1116_379# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0952 AS=0.0441 PD=0.823333 PS=0.63 NRD=30.4759 NRS=23.443 M=1 R=2.8
+ SA=75003.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1014 N_A_1158_93#_M1014_d N_A_957_379#_M1014_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1904 PD=2.21 PS=1.64667 NRD=0 NRS=5.8509 M=1
+ R=5.6 SA=75002.1 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 N_Q_M1015_d N_A_1158_93#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.9271 P=20.81
*
.include "sky130_fd_sc_lp__dfxtp_1.pxi.spice"
*
.ends
*
*
