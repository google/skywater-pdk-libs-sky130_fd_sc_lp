* NGSPICE file created from sky130_fd_sc_lp__or2_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or2_2 A B VGND VNB VPB VPWR X
M1000 a_131_390# B a_48_390# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1001 VPWR a_48_390# X VPB phighvt w=1.26e+06u l=150000u
+  ad=7.14e+11p pd=6.32e+06u as=3.528e+11p ps=3.08e+06u
M1002 VGND a_48_390# X VNB nshort w=840000u l=150000u
+  ad=6.027e+11p pd=6.01e+06u as=2.352e+11p ps=2.24e+06u
M1003 VGND A a_48_390# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1004 a_48_390# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_48_390# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_131_390# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_48_390# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

