* File: sky130_fd_sc_lp__nor4bb_lp.pex.spice
* Created: Fri Aug 28 10:59:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%C_N 2 5 7 9 12 14 16 17 18 19 20 24 26
c53 2 0 7.95967e-20 $X=0.607 $Y=1.658
r54 24 26 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.607 $Y=1.34
+ $X2=0.607 $Y2=1.175
r55 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.34 $X2=0.63 $Y2=1.34
r56 20 25 10.1228 $w=3.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.65 $Y=1.665
+ $X2=0.65 $Y2=1.34
r57 19 25 1.40162 $w=3.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.65 $Y=1.295
+ $X2=0.65 $Y2=1.34
r58 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.005 $Y=0.73
+ $X2=1.005 $Y2=0.445
r59 13 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.72 $Y=0.805
+ $X2=0.645 $Y2=0.805
r60 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.93 $Y=0.805
+ $X2=1.005 $Y2=0.73
r61 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.93 $Y=0.805
+ $X2=0.72 $Y2=0.805
r62 10 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.645 $Y=0.88
+ $X2=0.645 $Y2=0.805
r63 10 26 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.645 $Y=0.88
+ $X2=0.645 $Y2=1.175
r64 7 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.645 $Y=0.73
+ $X2=0.645 $Y2=0.805
r65 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.645 $Y=0.73 $X2=0.645
+ $Y2=0.445
r66 5 17 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.545 $Y=2.545
+ $X2=0.545 $Y2=1.845
r67 2 17 33.9275 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.607 $Y=1.658
+ $X2=0.607 $Y2=1.845
r68 1 24 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.607 $Y=1.362
+ $X2=0.607 $Y2=1.34
r69 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.607 $Y=1.362
+ $X2=0.607 $Y2=1.658
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%A_27_409# 1 2 9 13 17 21 25 27 31 35 38 39
+ 44
c82 44 0 1.98942e-19 $X=1.795 $Y=1.455
r83 43 44 12.7768 $w=6.7e-07 $l=1.6e-07 $layer=POLY_cond $X=1.635 $Y=1.455
+ $X2=1.795 $Y2=1.455
r84 42 43 15.971 $w=6.7e-07 $l=2e-07 $layer=POLY_cond $X=1.435 $Y=1.455
+ $X2=1.635 $Y2=1.455
r85 36 42 17.1689 $w=6.7e-07 $l=2.15e-07 $layer=POLY_cond $X=1.22 $Y=1.455
+ $X2=1.435 $Y2=1.455
r86 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.22
+ $Y=1.285 $X2=1.22 $Y2=1.285
r87 33 35 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.22 $Y=0.995
+ $X2=1.22 $Y2=1.285
r88 32 38 3.75155 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.595 $Y=0.91
+ $X2=0.355 $Y2=0.91
r89 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.055 $Y=0.91
+ $X2=1.22 $Y2=0.995
r90 31 32 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.055 $Y=0.91
+ $X2=0.595 $Y2=0.91
r91 27 29 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.24 $Y=2.19
+ $X2=0.24 $Y2=2.9
r92 25 39 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=2.15
+ $X2=0.24 $Y2=2.025
r93 25 27 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=0.24 $Y=2.15 $X2=0.24
+ $Y2=2.19
r94 23 38 2.92809 $w=3.25e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.2 $Y=0.995
+ $X2=0.355 $Y2=0.91
r95 23 39 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.2 $Y=0.995
+ $X2=0.2 $Y2=2.025
r96 19 38 2.92809 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.355 $Y=0.825
+ $X2=0.355 $Y2=0.91
r97 19 21 8.846 $w=4.78e-07 $l=3.55e-07 $layer=LI1_cond $X=0.355 $Y=0.825
+ $X2=0.355 $Y2=0.47
r98 15 44 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.795 $Y=1.12
+ $X2=1.795 $Y2=1.455
r99 15 17 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.795 $Y=1.12
+ $X2=1.795 $Y2=0.445
r100 11 43 25.9839 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.635 $Y=1.79
+ $X2=1.635 $Y2=1.455
r101 11 13 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.635 $Y=1.79
+ $X2=1.635 $Y2=2.545
r102 7 42 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.435 $Y=1.12
+ $X2=1.435 $Y2=1.455
r103 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.435 $Y=1.12
+ $X2=1.435 $Y2=0.445
r104 2 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r105 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r106 1 21 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.285
+ $Y=0.235 $X2=0.43 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%A_430_21# 1 2 9 11 12 15 19 22 23 24 27 32
+ 37 39 41 44
c86 37 0 2.26962e-19 $X=2.89 $Y=1.33
r87 44 45 31.0318 $w=3.4e-07 $l=7.5e-08 $layer=POLY_cond $X=2.68 $Y=1.24
+ $X2=2.68 $Y2=1.165
r88 41 43 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.43 $Y=0.455
+ $X2=5.43 $Y2=0.645
r89 35 47 32.1596 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.33
+ $X2=2.68 $Y2=1.495
r90 35 44 15.2746 $w=3.4e-07 $l=9e-08 $layer=POLY_cond $X=2.68 $Y=1.33 $X2=2.68
+ $Y2=1.24
r91 34 37 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.685 $Y=1.33
+ $X2=2.89 $Y2=1.33
r92 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.685
+ $Y=1.33 $X2=2.685 $Y2=1.33
r93 32 39 2.44685 $w=3.95e-07 $l=2.64102e-07 $layer=LI1_cond $X=5.51 $Y=1.675
+ $X2=5.285 $Y2=1.76
r94 32 43 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=5.51 $Y=1.675
+ $X2=5.51 $Y2=0.645
r95 27 29 13.697 $w=6.18e-07 $l=7.1e-07 $layer=LI1_cond $X=5.285 $Y=2.19
+ $X2=5.285 $Y2=2.9
r96 25 39 2.44685 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=5.285 $Y=1.845
+ $X2=5.285 $Y2=1.76
r97 25 27 6.6556 $w=6.18e-07 $l=3.45e-07 $layer=LI1_cond $X=5.285 $Y=1.845
+ $X2=5.285 $Y2=2.19
r98 23 39 4.49522 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=4.975 $Y=1.76
+ $X2=5.285 $Y2=1.76
r99 23 24 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=4.975 $Y=1.76
+ $X2=2.975 $Y2=1.76
r100 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.89 $Y=1.675
+ $X2=2.975 $Y2=1.76
r101 21 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=1.495
+ $X2=2.89 $Y2=1.33
r102 21 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.89 $Y=1.495
+ $X2=2.89 $Y2=1.675
r103 19 47 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.725 $Y=2.195
+ $X2=2.725 $Y2=1.495
r104 15 45 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.585 $Y=0.445
+ $X2=2.585 $Y2=1.165
r105 11 44 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.51 $Y=1.24
+ $X2=2.68 $Y2=1.24
r106 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.51 $Y=1.24
+ $X2=2.3 $Y2=1.24
r107 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.225 $Y=1.165
+ $X2=2.3 $Y2=1.24
r108 7 9 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.225 $Y=1.165
+ $X2=2.225 $Y2=0.445
r109 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=5
+ $Y=2.045 $X2=5.14 $Y2=2.9
r110 2 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5
+ $Y=2.045 $X2=5.14 $Y2=2.19
r111 1 41 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.235 $X2=5.43 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%B 1 3 4 5 6 8 10 13 15 16 23
c50 15 0 3.21658e-20 $X=3.405 $Y=0.805
c51 5 0 2.802e-20 $X=3.12 $Y=0.805
r52 21 23 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=3.55 $Y=1.33
+ $X2=3.815 $Y2=1.33
r53 18 21 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.405 $Y=1.33
+ $X2=3.55 $Y2=1.33
r54 16 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.33 $X2=3.55 $Y2=1.33
r55 11 23 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.495
+ $X2=3.815 $Y2=1.33
r56 11 13 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=3.815 $Y=1.495
+ $X2=3.815 $Y2=2.545
r57 10 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.405 $Y=1.165
+ $X2=3.405 $Y2=1.33
r58 9 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.405 $Y=0.88
+ $X2=3.405 $Y2=0.805
r59 9 10 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.405 $Y=0.88
+ $X2=3.405 $Y2=1.165
r60 6 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.405 $Y=0.73
+ $X2=3.405 $Y2=0.805
r61 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.405 $Y=0.73 $X2=3.405
+ $Y2=0.445
r62 4 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.33 $Y=0.805
+ $X2=3.405 $Y2=0.805
r63 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.33 $Y=0.805 $X2=3.12
+ $Y2=0.805
r64 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.045 $Y=0.73
+ $X2=3.12 $Y2=0.805
r65 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.045 $Y=0.73 $X2=3.045
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%A 1 3 4 5 6 8 11 14 16 17 18 22
c52 18 0 3.21658e-20 $X=4.56 $Y=1.295
r53 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.345
+ $Y=0.99 $X2=4.345 $Y2=0.99
r54 18 23 3.83816 $w=6.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.56 $Y=1.16
+ $X2=4.345 $Y2=1.16
r55 17 23 4.73076 $w=6.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.08 $Y=1.16
+ $X2=4.345 $Y2=1.16
r56 15 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.345 $Y=1.33
+ $X2=4.345 $Y2=0.99
r57 15 16 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.33
+ $X2=4.345 $Y2=1.495
r58 13 22 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.345 $Y=0.88
+ $X2=4.345 $Y2=0.99
r59 13 14 13.5877 $w=2.4e-07 $l=2.2798e-07 $layer=POLY_cond $X=4.345 $Y=0.88
+ $X2=4.18 $Y2=0.73
r60 11 16 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=4.305 $Y=2.545
+ $X2=4.305 $Y2=1.495
r61 6 14 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.255 $Y=0.73
+ $X2=4.18 $Y2=0.73
r62 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.255 $Y=0.73 $X2=4.255
+ $Y2=0.445
r63 4 14 12.1617 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.18 $Y=0.805
+ $X2=4.18 $Y2=0.73
r64 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.18 $Y=0.805 $X2=3.91
+ $Y2=0.805
r65 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.835 $Y=0.73
+ $X2=3.91 $Y2=0.805
r66 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.835 $Y=0.73 $X2=3.835
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%D_N 3 7 11 13 16 17
r32 16 18 65.5974 $w=5.4e-07 $l=5.05e-07 $layer=POLY_cond $X=5.02 $Y=0.99
+ $X2=5.02 $Y2=1.495
r33 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.02
+ $Y=0.99 $X2=5.02 $Y2=0.99
r34 13 17 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5.02 $Y=1.295
+ $X2=5.02 $Y2=0.99
r35 9 16 31.5348 $w=2.7e-07 $l=2.64953e-07 $layer=POLY_cond $X=5.215 $Y=0.825
+ $X2=5.02 $Y2=0.99
r36 9 11 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=5.215 $Y=0.825
+ $X2=5.215 $Y2=0.445
r37 7 18 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=4.875 $Y=2.545
+ $X2=4.875 $Y2=1.495
r38 1 16 31.5348 $w=2.7e-07 $l=2.64953e-07 $layer=POLY_cond $X=4.825 $Y=0.825
+ $X2=5.02 $Y2=0.99
r39 1 3 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4.825 $Y=0.825
+ $X2=4.825 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%VPWR 1 2 11 17 21 23 33 34 37 40
r42 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r43 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 34 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r45 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r46 31 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=3.33
+ $X2=4.57 $Y2=3.33
r47 31 33 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=4.735 $Y=3.33
+ $X2=5.52 $Y2=3.33
r48 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r49 29 30 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 27 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 26 29 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 26 27 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r54 24 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 23 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=3.33
+ $X2=4.57 $Y2=3.33
r56 23 29 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.405 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 21 30 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 21 27 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 17 20 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.57 $Y=2.19 $X2=4.57
+ $Y2=2.9
r60 15 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=3.245
+ $X2=4.57 $Y2=3.33
r61 15 20 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.57 $Y=3.245
+ $X2=4.57 $Y2=2.9
r62 11 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.19 $X2=0.81
+ $Y2=2.9
r63 9 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245 $X2=0.81
+ $Y2=3.33
r64 9 14 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.9
r65 2 20 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=2.045 $X2=4.57 $Y2=2.9
r66 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=2.045 $X2=4.57 $Y2=2.19
r67 1 14 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.9
r68 1 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%A_245_409# 1 2 7 9 11 18
r33 12 16 4.64076 $w=1.7e-07 $l=2.0106e-07 $layer=LI1_cond $X=1.535 $Y=2.27
+ $X2=1.37 $Y2=2.19
r34 11 18 4.64076 $w=1.7e-07 $l=2.0106e-07 $layer=LI1_cond $X=2.825 $Y=2.27
+ $X2=2.99 $Y2=2.19
r35 11 12 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=2.825 $Y=2.27
+ $X2=1.535 $Y2=2.27
r36 7 16 3.12541 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=2.355
+ $X2=1.37 $Y2=2.19
r37 7 9 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=1.37 $Y=2.355
+ $X2=1.37 $Y2=2.9
r38 2 18 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=2.85
+ $Y=1.695 $X2=2.99 $Y2=2.19
r39 1 16 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.045 $X2=1.37 $Y2=2.19
r40 1 9 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.045 $X2=1.37 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%A_352_409# 1 2 9 11 12 13 15
r28 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.895 $X2=3.55
+ $Y2=2.98
r29 13 15 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=3.55 $Y=2.895
+ $X2=3.55 $Y2=2.19
r30 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=2.98
+ $X2=3.55 $Y2=2.98
r31 11 12 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=3.385 $Y=2.98
+ $X2=2.065 $Y2=2.98
r32 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.9 $Y=2.895
+ $X2=2.065 $Y2=2.98
r33 7 9 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.9 $Y=2.895 $X2=1.9
+ $Y2=2.8
r34 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=2.045 $X2=3.55 $Y2=2.9
r35 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=2.045 $X2=3.55 $Y2=2.19
r36 1 9 600 $w=1.7e-07 $l=8.22025e-07 $layer=licon1_PDIFF $count=1 $X=1.76
+ $Y=2.045 $X2=1.9 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%Y 1 2 3 10 14 18 20 24 25 34 40
r65 34 40 0.168462 $w=7.08e-07 $l=1e-08 $layer=LI1_cond $X=1.92 $Y=1.675
+ $X2=1.92 $Y2=1.665
r66 25 34 2.56161 $w=7.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=1.84
+ $X2=1.92 $Y2=1.675
r67 25 40 0.640155 $w=7.08e-07 $l=3.8e-08 $layer=LI1_cond $X=1.92 $Y=1.627
+ $X2=1.92 $Y2=1.665
r68 24 25 5.59293 $w=7.08e-07 $l=3.32e-07 $layer=LI1_cond $X=1.92 $Y=1.295
+ $X2=1.92 $Y2=1.627
r69 22 23 8.28752 $w=6.33e-07 $l=4.3e-07 $layer=LI1_cond $X=1.92 $Y=0.47
+ $X2=1.92 $Y2=0.9
r70 20 24 5.22231 $w=7.08e-07 $l=3.1e-07 $layer=LI1_cond $X=1.92 $Y=0.985
+ $X2=1.92 $Y2=1.295
r71 20 23 1.6326 $w=7.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=0.985 $X2=1.92
+ $Y2=0.9
r72 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.62 $Y=0.815
+ $X2=3.62 $Y2=0.47
r73 12 25 5.51135 $w=3.3e-07 $l=3.55e-07 $layer=LI1_cond $X=2.275 $Y=1.84
+ $X2=1.92 $Y2=1.84
r74 12 14 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.275 $Y=1.84
+ $X2=2.46 $Y2=1.84
r75 11 23 8.66331 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=2.275 $Y=0.9
+ $X2=1.92 $Y2=0.9
r76 10 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.455 $Y=0.9
+ $X2=3.62 $Y2=0.815
r77 10 11 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=3.455 $Y=0.9
+ $X2=2.275 $Y2=0.9
r78 3 14 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.695 $X2=2.46 $Y2=1.84
r79 2 18 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.48
+ $Y=0.235 $X2=3.62 $Y2=0.47
r80 1 22 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.87
+ $Y=0.235 $X2=2.01 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_LP%VGND 1 2 3 12 16 20 22 24 29 34 44 45 48
+ 51 54
r82 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r83 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r84 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r85 45 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r86 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r87 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.635 $Y=0 $X2=4.47
+ $Y2=0
r88 42 44 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=4.635 $Y=0 $X2=5.52
+ $Y2=0
r89 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r90 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r91 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r92 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r93 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r94 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.8
+ $Y2=0
r95 35 37 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=3.12
+ $Y2=0
r96 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.47
+ $Y2=0
r97 34 40 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.305 $Y=0 $X2=4.08
+ $Y2=0
r98 33 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r99 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r100 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r101 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r102 30 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r103 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=0 $X2=2.8
+ $Y2=0
r104 29 32 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.635 $Y=0
+ $X2=1.68 $Y2=0
r105 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r106 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r107 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r108 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r109 22 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r110 22 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r111 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.47 $Y=0.085
+ $X2=4.47 $Y2=0
r112 18 20 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.47 $Y=0.085
+ $X2=4.47 $Y2=0.43
r113 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0.085 $X2=2.8
+ $Y2=0
r114 14 16 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.8 $Y=0.085
+ $X2=2.8 $Y2=0.425
r115 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r116 10 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.43
r117 3 20 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=4.33
+ $Y=0.235 $X2=4.47 $Y2=0.43
r118 2 16 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=2.66
+ $Y=0.235 $X2=2.8 $Y2=0.425
r119 1 12 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.22 $Y2=0.43
.ends

