* NGSPICE file created from sky130_fd_sc_lp__a2111o_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_86_275# B1 VGND VNB nshort w=840000u l=150000u
+  ad=5.166e+11p pd=4.59e+06u as=1.512e+12p ps=1.032e+07u
M1001 a_607_367# B1 a_499_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=8.253e+11p pd=6.35e+06u as=4.914e+11p ps=3.3e+06u
M1002 VGND A2 a_715_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=3.276e+11p ps=2.46e+06u
M1003 X a_86_275# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1004 a_86_275# D1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_86_275# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.1592e+12p ps=9.4e+06u
M1006 VGND a_86_275# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_607_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_427_367# D1 a_86_275# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=3.339e+11p ps=3.05e+06u
M1009 VGND C1 a_86_275# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_86_275# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_499_367# C1 a_427_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_607_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_715_49# A1 a_86_275# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

