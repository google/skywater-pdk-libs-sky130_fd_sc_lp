* File: sky130_fd_sc_lp__inv_2.pxi.spice
* Created: Wed Sep  2 09:55:52 2020
* 
x_PM_SKY130_FD_SC_LP__INV_2%A N_A_c_25_n N_A_M1000_g N_A_M1001_g N_A_c_27_n
+ N_A_M1002_g N_A_M1003_g A A N_A_c_30_n PM_SKY130_FD_SC_LP__INV_2%A
x_PM_SKY130_FD_SC_LP__INV_2%VPWR N_VPWR_M1001_d N_VPWR_M1003_d N_VPWR_c_59_n
+ N_VPWR_c_60_n N_VPWR_c_61_n N_VPWR_c_62_n VPWR N_VPWR_c_63_n N_VPWR_c_58_n
+ PM_SKY130_FD_SC_LP__INV_2%VPWR
x_PM_SKY130_FD_SC_LP__INV_2%Y N_Y_M1000_d N_Y_M1001_s Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__INV_2%Y
x_PM_SKY130_FD_SC_LP__INV_2%VGND N_VGND_M1000_s N_VGND_M1002_s N_VGND_c_95_n
+ N_VGND_c_96_n N_VGND_c_97_n N_VGND_c_98_n VGND N_VGND_c_99_n N_VGND_c_100_n
+ PM_SKY130_FD_SC_LP__INV_2%VGND
cc_1 VNB N_A_c_25_n 0.0200192f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.295
cc_2 VNB N_A_M1001_g 0.00178952f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_3 VNB N_A_c_27_n 0.020651f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.295
cc_4 VNB N_A_M1003_g 0.00232428f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_5 VNB A 0.0203343f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A_c_30_n 0.0762774f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.46
cc_7 VNB N_VPWR_c_58_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB Y 0.00471356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_VGND_c_95_n 0.0115187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_VGND_c_96_n 0.0353276f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.765
cc_11 VNB N_VGND_c_97_n 0.0124043f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.625
cc_12 VNB N_VGND_c_98_n 0.048351f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_13 VNB N_VGND_c_99_n 0.0158071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_100_n 0.11417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VPB N_A_M1001_g 0.0251188f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_16 VPB N_A_M1003_g 0.0272177f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_17 VPB A 0.00719599f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_18 VPB N_VPWR_c_59_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_19 VPB N_VPWR_c_60_n 0.0483699f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.765
cc_20 VPB N_VPWR_c_61_n 0.0123785f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_21 VPB N_VPWR_c_62_n 0.0583694f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_22 VPB N_VPWR_c_63_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0.33 $Y2=1.46
cc_23 VPB N_VPWR_c_58_n 0.0456603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_24 VPB Y 0.00319138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 N_A_M1001_g N_VPWR_c_60_n 0.0188656f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_26 N_A_M1003_g N_VPWR_c_60_n 7.92904e-19 $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_27 A N_VPWR_c_60_n 0.026915f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_28 N_A_c_30_n N_VPWR_c_60_n 0.00129037f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_29 N_A_M1003_g N_VPWR_c_62_n 0.0076281f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_30 N_A_M1001_g N_VPWR_c_63_n 0.00486043f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_31 N_A_M1003_g N_VPWR_c_63_n 0.00585385f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_32 N_A_M1001_g N_VPWR_c_58_n 0.00824727f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_33 N_A_M1003_g N_VPWR_c_58_n 0.0115127f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_34 N_A_c_25_n Y 0.00230243f $X=0.485 $Y=1.295 $X2=0 $Y2=0
cc_35 N_A_M1001_g Y 0.00356248f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_36 N_A_c_27_n Y 0.00373469f $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_37 N_A_M1003_g Y 0.00580911f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_38 A Y 0.0403576f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_39 N_A_c_30_n Y 0.0297332f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_40 N_A_c_25_n N_VGND_c_96_n 0.0138736f $X=0.485 $Y=1.295 $X2=0 $Y2=0
cc_41 N_A_c_27_n N_VGND_c_96_n 4.88726e-19 $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_42 A N_VGND_c_96_n 0.0269149f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_43 N_A_c_30_n N_VGND_c_96_n 0.00141307f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_44 N_A_c_27_n N_VGND_c_98_n 0.00714464f $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_45 N_A_c_25_n N_VGND_c_99_n 0.00400407f $X=0.485 $Y=1.295 $X2=0 $Y2=0
cc_46 N_A_c_27_n N_VGND_c_99_n 0.00482246f $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_47 N_A_c_25_n N_VGND_c_100_n 0.00774504f $X=0.485 $Y=1.295 $X2=0 $Y2=0
cc_48 N_A_c_27_n N_VGND_c_100_n 0.00965768f $X=0.915 $Y=1.295 $X2=0 $Y2=0
cc_49 N_VPWR_c_58_n N_Y_M1001_s 0.00397496f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_50 N_VPWR_c_62_n Y 0.00152359f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_51 N_VPWR_c_63_n Y 0.0138717f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_52 N_VPWR_c_58_n Y 0.00886411f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_53 N_VPWR_c_62_n N_VGND_c_98_n 0.0110287f $X=1.13 $Y=1.98 $X2=0 $Y2=0
cc_54 Y N_VGND_c_96_n 0.0291152f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_55 Y N_VGND_c_98_n 0.00465095f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_56 Y N_VGND_c_99_n 0.0124036f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_57 Y N_VGND_c_100_n 0.00864148f $X=0.635 $Y=0.47 $X2=0 $Y2=0
