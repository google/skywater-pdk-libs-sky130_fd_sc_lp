* File: sky130_fd_sc_lp__dlxtn_2.pex.spice
* Created: Wed Sep  2 09:48:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXTN_2%D 3 6 8 9 10 15 17
c36 15 0 1.10902e-19 $X=0.655 $Y=1.345
r37 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.345
+ $X2=0.655 $Y2=1.51
r38 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.345
+ $X2=0.655 $Y2=1.18
r39 9 10 19.0749 $w=2.88e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.345 $X2=1.68
+ $Y2=1.345
r40 8 9 21.658 $w=2.88e-07 $l=5.45e-07 $layer=LI1_cond $X=0.655 $Y=1.345 $X2=1.2
+ $Y2=1.345
r41 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.655
+ $Y=1.345 $X2=0.655 $Y2=1.345
r42 6 18 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=0.705 $Y=2.725
+ $X2=0.705 $Y2=1.51
r43 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.625 $Y=0.86
+ $X2=0.625 $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_2%GATE_N 1 3 6 8 11 12 13 14 15 20
c44 8 0 1.22905e-19 $X=1.55 $Y=1.255
r45 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=0.36
+ $X2=1.715 $Y2=0.525
r46 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.715
+ $Y=0.36 $X2=1.715 $Y2=0.36
r47 15 21 14.0503 $w=3.63e-07 $l=4.45e-07 $layer=LI1_cond $X=2.16 $Y=0.457
+ $X2=1.715 $Y2=0.457
r48 14 21 1.10508 $w=3.63e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=0.457
+ $X2=1.715 $Y2=0.457
r49 13 14 15.1554 $w=3.63e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.457
+ $X2=1.68 $Y2=0.457
r50 11 23 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=1.625 $Y=1.18
+ $X2=1.625 $Y2=0.525
r51 9 12 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.21 $Y=1.255
+ $X2=1.135 $Y2=1.255
r52 8 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.55 $Y=1.255
+ $X2=1.625 $Y2=1.18
r53 8 9 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.55 $Y=1.255 $X2=1.21
+ $Y2=1.255
r54 4 12 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.135 $Y=1.33
+ $X2=1.135 $Y2=1.255
r55 4 6 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=1.135 $Y=1.33
+ $X2=1.135 $Y2=2.725
r56 1 12 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.135 $Y=1.18
+ $X2=1.135 $Y2=1.255
r57 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.135 $Y=1.18
+ $X2=1.135 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_2%A_242_130# 1 2 9 11 12 13 15 18 22 26 27 33
+ 35 36 40 41 42 43 45 47 50 51 53 54 57 58
c149 53 0 1.22905e-19 $X=2.175 $Y=0.985
c150 50 0 2.41741e-19 $X=3.87 $Y=2.08
r151 57 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=1.08
+ $X2=3.72 $Y2=0.915
r152 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.72
+ $Y=1.08 $X2=3.72 $Y2=1.08
r153 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.175
+ $Y=0.985 $X2=2.175 $Y2=0.985
r154 51 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.87 $Y=2.08
+ $X2=3.87 $Y2=2.245
r155 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.87
+ $Y=2.08 $X2=3.87 $Y2=2.08
r156 48 50 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.835 $Y=2.375
+ $X2=3.835 $Y2=2.08
r157 47 58 6.06832 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.835 $Y=2.045
+ $X2=3.835 $Y2=1.915
r158 47 50 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=3.835 $Y=2.045
+ $X2=3.835 $Y2=2.08
r159 45 56 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=1.165
+ $X2=3.815 $Y2=1.08
r160 45 58 39.2878 $w=2.18e-07 $l=7.5e-07 $layer=LI1_cond $X=3.815 $Y=1.165
+ $X2=3.815 $Y2=1.915
r161 44 53 7.54205 $w=1.95e-07 $l=4.29273e-07 $layer=LI1_cond $X=2.34 $Y=1.08
+ $X2=2.025 $Y2=0.81
r162 43 56 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.705 $Y=1.08
+ $X2=3.815 $Y2=1.08
r163 43 44 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=3.705 $Y=1.08
+ $X2=2.34 $Y2=1.08
r164 41 48 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.705 $Y=2.46
+ $X2=3.835 $Y2=2.375
r165 41 42 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.705 $Y=2.46
+ $X2=2.305 $Y2=2.46
r166 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.22 $Y=2.545
+ $X2=2.305 $Y2=2.46
r167 39 40 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.22 $Y=2.545
+ $X2=2.22 $Y2=2.905
r168 35 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=2.99
+ $X2=2.22 $Y2=2.905
r169 35 36 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.135 $Y=2.99
+ $X2=1.515 $Y2=2.99
r170 31 36 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.365 $Y=2.905
+ $X2=1.515 $Y2=2.99
r171 31 33 13.2531 $w=2.98e-07 $l=3.45e-07 $layer=LI1_cond $X=1.365 $Y=2.905
+ $X2=1.365 $Y2=2.56
r172 27 53 7.54205 $w=1.95e-07 $l=1.1e-07 $layer=LI1_cond $X=2.025 $Y=0.92
+ $X2=2.025 $Y2=0.81
r173 27 29 35.359 $w=2.18e-07 $l=6.75e-07 $layer=LI1_cond $X=2.025 $Y=0.92
+ $X2=1.35 $Y2=0.92
r174 25 54 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.175 $Y=1.325
+ $X2=2.175 $Y2=0.985
r175 25 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.175 $Y=1.325
+ $X2=2.175 $Y2=1.49
r176 24 54 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.175 $Y=0.915
+ $X2=2.175 $Y2=0.985
r177 22 65 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.78 $Y=2.615
+ $X2=3.78 $Y2=2.245
r178 18 61 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.63 $Y=0.445 $X2=3.63
+ $Y2=0.915
r179 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.84 $Y=0.765
+ $X2=2.84 $Y2=0.445
r180 12 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.34 $Y=0.84
+ $X2=2.175 $Y2=0.915
r181 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.765 $Y=0.84
+ $X2=2.84 $Y2=0.765
r182 11 12 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.765 $Y=0.84
+ $X2=2.34 $Y2=0.84
r183 9 26 633.266 $w=1.5e-07 $l=1.235e-06 $layer=POLY_cond $X=2.085 $Y=2.725
+ $X2=2.085 $Y2=1.49
r184 2 33 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1.21
+ $Y=2.405 $X2=1.35 $Y2=2.56
r185 1 29 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.21
+ $Y=0.65 $X2=1.35 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_2%A_57_130# 1 2 9 11 12 15 19 21 24 26 31 33
+ 35 36
c79 31 0 1.10902e-19 $X=0.41 $Y=0.86
c80 21 0 2.4855e-20 $X=0.225 $Y=1.66
r81 35 38 11.4197 $w=3.28e-07 $l=3.27e-07 $layer=LI1_cond $X=2.76 $Y=1.43
+ $X2=2.76 $Y2=1.757
r82 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.76
+ $Y=1.43 $X2=2.76 $Y2=1.43
r83 28 31 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.225 $Y=0.86
+ $X2=0.41 $Y2=0.86
r84 27 33 3.26102 $w=1.95e-07 $l=2.43e-07 $layer=LI1_cond $X=0.625 $Y=1.757
+ $X2=0.382 $Y2=1.757
r85 26 38 3.83364 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=1.757
+ $X2=2.76 $Y2=1.757
r86 26 27 112.047 $w=1.93e-07 $l=1.97e-06 $layer=LI1_cond $X=2.595 $Y=1.757
+ $X2=0.625 $Y2=1.757
r87 22 33 3.29278 $w=3.27e-07 $l=9.8e-08 $layer=LI1_cond $X=0.382 $Y=1.855
+ $X2=0.382 $Y2=1.757
r88 22 24 17.1397 $w=4.83e-07 $l=6.95e-07 $layer=LI1_cond $X=0.382 $Y=1.855
+ $X2=0.382 $Y2=2.55
r89 21 33 3.29278 $w=3.27e-07 $l=1.99695e-07 $layer=LI1_cond $X=0.225 $Y=1.66
+ $X2=0.382 $Y2=1.757
r90 20 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.225 $Y=1.025
+ $X2=0.225 $Y2=0.86
r91 20 21 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.225 $Y=1.025
+ $X2=0.225 $Y2=1.66
r92 18 36 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=2.775 $Y=1.755
+ $X2=2.775 $Y2=1.43
r93 18 19 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=2.775 $Y=1.755
+ $X2=2.775 $Y2=1.935
r94 17 36 24.8449 $w=3.6e-07 $l=1.55e-07 $layer=POLY_cond $X=2.775 $Y=1.275
+ $X2=2.775 $Y2=1.43
r95 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.27 $Y=1.125
+ $X2=3.27 $Y2=0.445
r96 12 17 150.063 $w=5.6e-08 $l=2.14243e-07 $layer=POLY_cond $X=2.955 $Y=1.2
+ $X2=2.775 $Y2=1.275
r97 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.195 $Y=1.2
+ $X2=3.27 $Y2=1.125
r98 11 12 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.195 $Y=1.2
+ $X2=2.955 $Y2=1.2
r99 9 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.88 $Y=2.725
+ $X2=2.88 $Y2=1.935
r100 2 24 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.365
+ $Y=2.405 $X2=0.49 $Y2=2.55
r101 1 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.285
+ $Y=0.65 $X2=0.41 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_2%A_349_481# 1 2 9 11 12 15 18 21 24 26 27 30
+ 32 33 36 37 39 43
c113 21 0 1.07053e-19 $X=3.33 $Y=2.205
c114 11 0 1.66779e-20 $X=4.095 $Y=1.56
r115 43 48 75.0636 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.26 $Y=1.005
+ $X2=4.26 $Y2=1.335
r116 43 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.26 $Y=1.005
+ $X2=4.26 $Y2=0.84
r117 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.26
+ $Y=1.005 $X2=4.26 $Y2=1.005
r118 39 42 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.26 $Y=0.73
+ $X2=4.26 $Y2=1.005
r119 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.33
+ $Y=1.7 $X2=3.33 $Y2=1.7
r120 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.33 $Y=2.035
+ $X2=3.33 $Y2=1.7
r121 32 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=0.73
+ $X2=4.26 $Y2=0.73
r122 32 33 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=4.095 $Y=0.73
+ $X2=2.72 $Y2=0.73
r123 28 33 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.59 $Y=0.645
+ $X2=2.72 $Y2=0.73
r124 28 30 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=2.59 $Y=0.645
+ $X2=2.59 $Y2=0.44
r125 26 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.165 $Y=2.12
+ $X2=3.33 $Y2=2.035
r126 26 27 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.165 $Y=2.12
+ $X2=1.955 $Y2=2.12
r127 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.83 $Y=2.205
+ $X2=1.955 $Y2=2.12
r128 22 24 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.83 $Y=2.205
+ $X2=1.83 $Y2=2.57
r129 20 37 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.33 $Y=2.04
+ $X2=3.33 $Y2=1.7
r130 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=2.04
+ $X2=3.33 $Y2=2.205
r131 19 37 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.33 $Y=1.635
+ $X2=3.33 $Y2=1.7
r132 18 48 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=4.17 $Y=1.485
+ $X2=4.17 $Y2=1.335
r133 15 47 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.17 $Y=0.445
+ $X2=4.17 $Y2=0.84
r134 12 19 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.495 $Y=1.56
+ $X2=3.33 $Y2=1.635
r135 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.095 $Y=1.56
+ $X2=4.17 $Y2=1.485
r136 11 12 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.095 $Y=1.56
+ $X2=3.495 $Y2=1.56
r137 9 21 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.24 $Y=2.725
+ $X2=3.24 $Y2=2.205
r138 2 24 600 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=2.405 $X2=1.87 $Y2=2.57
r139 1 30 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.235 $X2=2.625 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_2%A_849_419# 1 2 9 13 15 17 20 22 26 30 35 39
+ 40 41 44 48 52 57 60 64 65 66 67
c118 64 0 1.66779e-20 $X=4.65 $Y=1.74
c119 39 0 1.36635e-19 $X=6.21 $Y=1.435
c120 35 0 1.34688e-19 $X=4.65 $Y=2.095
r121 64 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.65
+ $Y=1.74 $X2=4.65 $Y2=1.74
r122 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6
+ $Y=1.435 $X2=6 $Y2=1.435
r123 58 67 2.79962 $w=3.3e-07 $l=3.71147e-07 $layer=LI1_cond $X=5.705 $Y=1.435
+ $X2=5.415 $Y2=1.62
r124 58 60 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.705 $Y=1.435
+ $X2=6 $Y2=1.435
r125 57 67 3.30809 $w=1.7e-07 $l=4.40738e-07 $layer=LI1_cond $X=5.62 $Y=1.27
+ $X2=5.415 $Y2=1.62
r126 57 66 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.62 $Y=1.27
+ $X2=5.62 $Y2=1.09
r127 52 54 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=5.56 $Y=1.825
+ $X2=5.56 $Y2=2.795
r128 50 67 3.30809 $w=2.9e-07 $l=2.31409e-07 $layer=LI1_cond $X=5.56 $Y=1.79
+ $X2=5.415 $Y2=1.62
r129 50 52 1.39088 $w=2.88e-07 $l=3.5e-08 $layer=LI1_cond $X=5.56 $Y=1.79
+ $X2=5.56 $Y2=1.825
r130 46 66 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=5.522 $Y=0.908
+ $X2=5.522 $Y2=1.09
r131 46 48 15.408 $w=3.63e-07 $l=4.88e-07 $layer=LI1_cond $X=5.522 $Y=0.908
+ $X2=5.522 $Y2=0.42
r132 45 64 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=1.705
+ $X2=4.65 $Y2=1.705
r133 44 67 2.79962 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.415 $Y=1.705
+ $X2=5.415 $Y2=1.62
r134 44 45 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.415 $Y=1.705
+ $X2=4.815 $Y2=1.705
r135 39 61 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=6.21 $Y=1.435 $X2=6
+ $Y2=1.435
r136 39 40 6.91837 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.21 $Y=1.435
+ $X2=6.285 $Y2=1.435
r137 38 65 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.65 $Y=1.575
+ $X2=4.65 $Y2=1.74
r138 35 65 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.65 $Y=2.095
+ $X2=4.65 $Y2=1.74
r139 32 35 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.32 $Y=2.17
+ $X2=4.65 $Y2=2.17
r140 28 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.715 $Y=1.57
+ $X2=6.715 $Y2=1.495
r141 28 30 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=6.715 $Y=1.57
+ $X2=6.715 $Y2=2.465
r142 24 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.715 $Y=1.42
+ $X2=6.715 $Y2=1.495
r143 24 26 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.715 $Y=1.42
+ $X2=6.715 $Y2=0.74
r144 23 40 6.91837 $w=1.5e-07 $l=1.00623e-07 $layer=POLY_cond $X=6.36 $Y=1.495
+ $X2=6.285 $Y2=1.435
r145 22 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.64 $Y=1.495
+ $X2=6.715 $Y2=1.495
r146 22 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.64 $Y=1.495
+ $X2=6.36 $Y2=1.495
r147 18 40 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.285 $Y=1.6
+ $X2=6.285 $Y2=1.435
r148 18 20 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=6.285 $Y=1.6
+ $X2=6.285 $Y2=2.465
r149 15 40 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.285 $Y=1.27
+ $X2=6.285 $Y2=1.435
r150 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.285 $Y=1.27
+ $X2=6.285 $Y2=0.74
r151 13 38 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=4.71 $Y=0.445
+ $X2=4.71 $Y2=1.575
r152 7 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.32 $Y=2.245
+ $X2=4.32 $Y2=2.17
r153 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.32 $Y=2.245
+ $X2=4.32 $Y2=2.615
r154 2 54 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.41
+ $Y=1.68 $X2=5.55 $Y2=2.795
r155 2 52 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.41
+ $Y=1.68 $X2=5.55 $Y2=1.825
r156 1 48 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.33
+ $Y=0.235 $X2=5.47 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_2%A_663_481# 1 2 9 12 14 18 23 24 25 27 30 31
+ 33 35
c99 30 0 1.36635e-19 $X=5.19 $Y=1.355
r100 31 36 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=5.217 $Y=1.355
+ $X2=5.217 $Y2=1.52
r101 31 35 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=5.217 $Y=1.355
+ $X2=5.217 $Y2=1.19
r102 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.19
+ $Y=1.355 $X2=5.19 $Y2=1.355
r103 28 33 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.775 $Y=1.355
+ $X2=4.69 $Y2=1.355
r104 28 30 24.2249 $w=1.88e-07 $l=4.15e-07 $layer=LI1_cond $X=4.775 $Y=1.355
+ $X2=5.19 $Y2=1.355
r105 27 33 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.69 $Y=1.26
+ $X2=4.69 $Y2=1.355
r106 26 27 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=4.69 $Y=0.475
+ $X2=4.69 $Y2=1.26
r107 24 33 4.81226 $w=1.85e-07 $l=8.74643e-08 $layer=LI1_cond $X=4.605 $Y=1.36
+ $X2=4.69 $Y2=1.355
r108 24 25 18.4848 $w=1.78e-07 $l=3e-07 $layer=LI1_cond $X=4.605 $Y=1.36
+ $X2=4.305 $Y2=1.36
r109 22 25 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.22 $Y=1.45
+ $X2=4.305 $Y2=1.36
r110 22 23 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=4.22 $Y=1.45
+ $X2=4.22 $Y2=2.715
r111 18 26 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.605 $Y=0.365
+ $X2=4.69 $Y2=0.475
r112 18 20 34.0495 $w=2.18e-07 $l=6.5e-07 $layer=LI1_cond $X=4.605 $Y=0.365
+ $X2=3.955 $Y2=0.365
r113 14 23 7.93686 $w=3.5e-07 $l=2.13307e-07 $layer=LI1_cond $X=4.135 $Y=2.89
+ $X2=4.22 $Y2=2.715
r114 14 16 22.3903 $w=3.48e-07 $l=6.8e-07 $layer=LI1_cond $X=4.135 $Y=2.89
+ $X2=3.455 $Y2=2.89
r115 12 36 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.335 $Y=2.31
+ $X2=5.335 $Y2=1.52
r116 9 35 171.913 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.255 $Y=0.655
+ $X2=5.255 $Y2=1.19
r117 2 16 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=2.405 $X2=3.455 $Y2=2.88
r118 1 20 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.235 $X2=3.955 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_2%VPWR 1 2 3 4 5 18 22 26 30 34 36 41 42 43 49
+ 56 64 69 75 78 87 91
r84 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r85 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r86 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r87 81 83 7.99975 $w=7.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.86 $Y=2.815
+ $X2=4.86 $Y2=3.33
r88 78 81 2.40769 $w=7.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.86 $Y=2.66
+ $X2=4.86 $Y2=2.815
r89 78 79 9.05078 $w=7.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.86 $Y=2.66
+ $X2=4.86 $Y2=2.495
r90 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r91 73 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r92 73 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r93 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r94 70 87 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.2 $Y=3.33
+ $X2=6.052 $Y2=3.33
r95 70 72 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.2 $Y=3.33 $X2=6.48
+ $Y2=3.33
r96 69 90 4.38699 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=7.002 $Y2=3.33
r97 69 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=6.48 $Y2=3.33
r98 68 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r99 68 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r100 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r101 65 83 9.95332 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=5.245 $Y=3.33
+ $X2=4.86 $Y2=3.33
r102 65 67 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.245 $Y=3.33
+ $X2=5.52 $Y2=3.33
r103 64 87 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=5.905 $Y=3.33
+ $X2=6.052 $Y2=3.33
r104 64 67 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.905 $Y=3.33
+ $X2=5.52 $Y2=3.33
r105 63 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 60 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r108 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r109 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r110 57 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.605 $Y2=3.33
r111 57 59 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 56 83 9.95332 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=4.475 $Y=3.33
+ $X2=4.86 $Y2=3.33
r113 56 62 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.475 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 55 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r116 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r118 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 49 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.605 $Y2=3.33
r120 49 54 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.16 $Y2=3.33
r121 47 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 43 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 43 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 41 46 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 41 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.92 $Y2=3.33
r127 40 51 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 40 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=0.92 $Y2=3.33
r129 36 39 37.9511 $w=2.88e-07 $l=9.55e-07 $layer=LI1_cond $X=6.95 $Y=1.98
+ $X2=6.95 $Y2=2.935
r130 34 90 3.05085 $w=2.9e-07 $l=1.07912e-07 $layer=LI1_cond $X=6.95 $Y=3.245
+ $X2=7.002 $Y2=3.33
r131 34 39 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=6.95 $Y=3.245
+ $X2=6.95 $Y2=2.935
r132 30 33 37.3079 $w=2.93e-07 $l=9.55e-07 $layer=LI1_cond $X=6.052 $Y=1.98
+ $X2=6.052 $Y2=2.935
r133 28 87 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.052 $Y=3.245
+ $X2=6.052 $Y2=3.33
r134 28 33 12.1104 $w=2.93e-07 $l=3.1e-07 $layer=LI1_cond $X=6.052 $Y=3.245
+ $X2=6.052 $Y2=2.935
r135 26 79 18.0382 $w=2.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.13 $Y=2.135
+ $X2=5.13 $Y2=2.495
r136 20 75 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=3.245
+ $X2=2.605 $Y2=3.33
r137 20 22 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=2.605 $Y=3.245
+ $X2=2.605 $Y2=2.88
r138 16 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=3.33
r139 16 18 30.655 $w=2.48e-07 $l=6.65e-07 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=2.58
r140 5 39 400 $w=1.7e-07 $l=1.1679e-06 $layer=licon1_PDIFF $count=1 $X=6.79
+ $Y=1.835 $X2=6.93 $Y2=2.935
r141 5 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.79
+ $Y=1.835 $X2=6.93 $Y2=1.98
r142 4 33 400 $w=1.7e-07 $l=1.16082e-06 $layer=licon1_PDIFF $count=1 $X=5.945
+ $Y=1.835 $X2=6.07 $Y2=2.935
r143 4 30 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.945
+ $Y=1.835 $X2=6.07 $Y2=1.98
r144 3 81 600 $w=1.7e-07 $l=9.07125e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=2.405 $X2=5.12 $Y2=2.815
r145 3 78 600 $w=1.7e-07 $l=3.27261e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=2.405 $X2=4.56 $Y2=2.66
r146 3 26 300 $w=1.7e-07 $l=8.49338e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=2.405 $X2=5.12 $Y2=2.135
r147 2 22 600 $w=1.7e-07 $l=6.48363e-07 $layer=licon1_PDIFF $count=1 $X=2.16
+ $Y=2.405 $X2=2.57 $Y2=2.88
r148 1 18 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=0.78
+ $Y=2.405 $X2=0.92 $Y2=2.58
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_2%Q 1 2 7 8 9 10 11 12 13 22
r20 13 40 5.87094 $w=2.63e-07 $l=1.35e-07 $layer=LI1_cond $X=6.502 $Y=2.775
+ $X2=6.502 $Y2=2.91
r21 12 13 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=6.502 $Y=2.405
+ $X2=6.502 $Y2=2.775
r22 11 12 19.3523 $w=2.63e-07 $l=4.45e-07 $layer=LI1_cond $X=6.502 $Y=1.96
+ $X2=6.502 $Y2=2.405
r23 10 11 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=6.502 $Y=1.665
+ $X2=6.502 $Y2=1.96
r24 9 10 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=6.502 $Y=1.295
+ $X2=6.502 $Y2=1.665
r25 8 9 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=6.502 $Y=0.925
+ $X2=6.502 $Y2=1.295
r26 7 8 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=6.502 $Y=0.555
+ $X2=6.502 $Y2=0.925
r27 7 22 3.91396 $w=2.63e-07 $l=9e-08 $layer=LI1_cond $X=6.502 $Y=0.555
+ $X2=6.502 $Y2=0.465
r28 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.36
+ $Y=1.835 $X2=6.5 $Y2=2.91
r29 2 11 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=6.36
+ $Y=1.835 $X2=6.5 $Y2=1.96
r30 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.36
+ $Y=0.32 $X2=6.5 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_2%VGND 1 2 3 4 5 19 22 26 30 32 34 39 41 43 51
+ 59 64 70 73 76 79 83
r87 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r88 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r89 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r90 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r91 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r92 68 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r93 68 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r94 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r95 65 79 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.2 $Y=0 $X2=6.052
+ $Y2=0
r96 65 67 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.2 $Y=0 $X2=6.48
+ $Y2=0
r97 64 82 4.38699 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=6.805 $Y=0 $X2=7.002
+ $Y2=0
r98 64 67 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.805 $Y=0 $X2=6.48
+ $Y2=0
r99 63 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r100 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r101 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r102 60 76 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=5.17 $Y=0 $X2=5.057
+ $Y2=0
r103 60 62 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.17 $Y=0 $X2=5.52
+ $Y2=0
r104 59 79 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=6.052 $Y2=0
r105 59 62 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.905 $Y=0
+ $X2=5.52 $Y2=0
r106 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r107 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r108 54 57 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r109 52 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.055
+ $Y2=0
r110 52 54 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.6
+ $Y2=0
r111 51 76 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=4.945 $Y=0
+ $X2=5.057 $Y2=0
r112 51 57 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.945 $Y=0
+ $X2=4.56 $Y2=0
r113 50 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r114 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r115 47 50 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r116 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r117 46 49 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r118 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r119 44 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=0 $X2=0.76
+ $Y2=0
r120 44 46 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.2
+ $Y2=0
r121 43 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.055
+ $Y2=0
r122 43 49 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.64
+ $Y2=0
r123 41 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r124 41 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r125 41 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r126 32 82 3.05085 $w=2.9e-07 $l=1.07912e-07 $layer=LI1_cond $X=6.95 $Y=0.085
+ $X2=7.002 $Y2=0
r127 32 34 15.101 $w=2.88e-07 $l=3.8e-07 $layer=LI1_cond $X=6.95 $Y=0.085
+ $X2=6.95 $Y2=0.465
r128 28 79 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.052 $Y=0.085
+ $X2=6.052 $Y2=0
r129 28 30 14.845 $w=2.93e-07 $l=3.8e-07 $layer=LI1_cond $X=6.052 $Y=0.085
+ $X2=6.052 $Y2=0.465
r130 24 76 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=5.057 $Y=0.085
+ $X2=5.057 $Y2=0
r131 24 26 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=5.057 $Y=0.085
+ $X2=5.057 $Y2=0.38
r132 20 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0
r133 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.36
r134 19 39 4.28816 $w=2.13e-07 $l=8e-08 $layer=LI1_cond $X=0.76 $Y=0.917
+ $X2=0.84 $Y2=0.917
r135 18 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0
r136 18 19 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=0.76 $Y=0.085
+ $X2=0.76 $Y2=0.81
r137 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.79
+ $Y=0.32 $X2=6.93 $Y2=0.465
r138 4 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.945
+ $Y=0.32 $X2=6.07 $Y2=0.465
r139 3 26 91 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=2 $X=4.785
+ $Y=0.235 $X2=5.04 $Y2=0.38
r140 2 22 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.055 $Y2=0.36
r141 1 39 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=0.7
+ $Y=0.65 $X2=0.84 $Y2=0.915
.ends

