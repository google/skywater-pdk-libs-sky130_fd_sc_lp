* File: sky130_fd_sc_lp__a32oi_m.spice
* Created: Wed Sep  2 09:28:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32oi_m.pex.spice"
.subckt sky130_fd_sc_lp__a32oi_m  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1009 A_152_47# N_B2_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1869 PD=0.63 PS=1.73 NRD=14.28 NRS=51.42 M=1 R=2.8 SA=75000.4 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g A_152_47# VNB NSHORT L=0.15 W=0.42 AD=0.06825
+ AS=0.0441 PD=0.745 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.7 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1001 A_319_47# N_A1_M1001_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.06825 PD=0.81 PS=0.745 NRD=39.996 NRS=12.852 M=1 R=2.8 SA=75001.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 A_427_47# N_A2_M1005_g A_319_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=39.996 M=1 R=2.8 SA=75001.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A3_M1006_g A_427_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g N_A_40_500#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1449 PD=0.7 PS=1.53 NRD=0 NRS=37.5088 M=1 R=2.8 SA=75000.3
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_40_500#_M1002_d N_B1_M1002_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_40_500#_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0756 AS=0.0756 PD=0.78 PS=0.78 NRD=0 NRS=28.1316 M=1 R=2.8 SA=75001.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_A_40_500#_M1004_d N_A2_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=37.5088 M=1 R=2.8 SA=75001.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A3_M1008_g N_A_40_500#_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_70 VPB 0 3.33391e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a32oi_m.pxi.spice"
*
.ends
*
*
