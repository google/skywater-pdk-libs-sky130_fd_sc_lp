* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_8 A0 A1 S VGND VNB VPB VPWR X
X0 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND S a_1179_311# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_1243_47# a_1179_311# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VPWR S a_1179_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_839_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_839_47# A1 a_84_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 VPWR S a_843_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X10 a_1243_419# A1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X11 a_1243_47# A0 a_84_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_84_21# A0 a_1243_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_843_419# A0 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X16 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_84_21# A1 a_1243_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X18 VGND a_1179_311# a_1243_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_1243_419# a_1179_311# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X22 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VGND a_84_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 X a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 VGND S a_839_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 VPWR a_1179_311# a_1243_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X28 VPWR a_84_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_843_419# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X31 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_84_21# A1 a_839_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X33 a_84_21# A0 a_843_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
.ends
