* NGSPICE file created from sky130_fd_sc_lp__nor3b_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor3b_2 A B C_N VGND VNB VPB VPWR Y
M1000 VGND a_27_131# Y VNB nshort w=840000u l=150000u
+  ad=1.2411e+12p pd=1.027e+07u as=7.938e+11p ps=6.93e+06u
M1001 VPWR C_N a_27_131# VPB phighvt w=420000u l=150000u
+  ad=7.791e+11p pd=7.47e+06u as=1.113e+11p ps=1.37e+06u
M1002 a_472_365# B a_217_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=1.0206e+12p ps=9.18e+06u
M1003 VGND B Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_27_131# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_217_365# a_27_131# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1007 Y B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A a_472_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_131# a_217_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_217_365# B a_472_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND C_N a_27_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1013 a_472_365# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

