* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_975_367# A2 a_720_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_101_23# B1 a_528_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_528_65# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 X a_101_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND a_101_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND A1 a_528_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 X a_101_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_101_23# A3 a_720_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_720_367# A3 a_101_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_528_65# B1 a_101_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VGND A3 a_528_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND a_101_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_528_65# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_720_367# A2 a_975_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 X a_101_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_528_65# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VGND A2 a_528_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VPWR a_101_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR A1 a_975_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_975_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VPWR a_101_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_101_23# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 X a_101_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 VPWR B1 a_101_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
