* File: sky130_fd_sc_lp__and2b_4.pxi.spice
* Created: Fri Aug 28 10:05:22 2020
* 
x_PM_SKY130_FD_SC_LP__AND2B_4%A_N N_A_N_M1004_g N_A_N_M1006_g A_N A_N A_N
+ N_A_N_c_73_n N_A_N_c_74_n PM_SKY130_FD_SC_LP__AND2B_4%A_N
x_PM_SKY130_FD_SC_LP__AND2B_4%A_213_23# N_A_213_23#_M1011_d N_A_213_23#_M1009_d
+ N_A_213_23#_M1001_g N_A_213_23#_M1000_g N_A_213_23#_M1007_g
+ N_A_213_23#_M1002_g N_A_213_23#_M1008_g N_A_213_23#_M1005_g
+ N_A_213_23#_M1012_g N_A_213_23#_M1013_g N_A_213_23#_c_176_p
+ N_A_213_23#_c_104_n N_A_213_23#_c_113_n N_A_213_23#_c_105_n
+ N_A_213_23#_c_183_p N_A_213_23#_c_148_p N_A_213_23#_c_122_p
+ N_A_213_23#_c_106_n N_A_213_23#_c_107_n N_A_213_23#_c_108_n
+ PM_SKY130_FD_SC_LP__AND2B_4%A_213_23#
x_PM_SKY130_FD_SC_LP__AND2B_4%B N_B_M1009_g N_B_M1010_g B N_B_c_216_n
+ PM_SKY130_FD_SC_LP__AND2B_4%B
x_PM_SKY130_FD_SC_LP__AND2B_4%A_43_367# N_A_43_367#_M1006_s N_A_43_367#_M1004_s
+ N_A_43_367#_M1011_g N_A_43_367#_M1003_g N_A_43_367#_c_256_n
+ N_A_43_367#_c_263_n N_A_43_367#_c_264_n N_A_43_367#_c_257_n
+ N_A_43_367#_c_258_n N_A_43_367#_c_259_n N_A_43_367#_c_260_n
+ PM_SKY130_FD_SC_LP__AND2B_4%A_43_367#
x_PM_SKY130_FD_SC_LP__AND2B_4%VPWR N_VPWR_M1004_d N_VPWR_M1002_s N_VPWR_M1013_s
+ N_VPWR_M1003_d N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n
+ N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n VPWR
+ N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_322_n
+ PM_SKY130_FD_SC_LP__AND2B_4%VPWR
x_PM_SKY130_FD_SC_LP__AND2B_4%X N_X_M1001_d N_X_M1008_d N_X_M1000_d N_X_M1005_d
+ N_X_c_382_n N_X_c_421_p N_X_c_383_n N_X_c_384_n N_X_c_423_p X X X
+ PM_SKY130_FD_SC_LP__AND2B_4%X
x_PM_SKY130_FD_SC_LP__AND2B_4%VGND N_VGND_M1006_d N_VGND_M1007_s N_VGND_M1012_s
+ N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n N_VGND_c_431_n N_VGND_c_432_n
+ N_VGND_c_433_n VGND N_VGND_c_434_n N_VGND_c_435_n N_VGND_c_436_n
+ N_VGND_c_437_n N_VGND_c_438_n PM_SKY130_FD_SC_LP__AND2B_4%VGND
cc_1 VNB N_A_N_M1004_g 0.0063596f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.045
cc_2 VNB A_N 0.0070705f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_N_c_73_n 0.036925f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.375
cc_4 VNB N_A_N_c_74_n 0.023177f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.21
cc_5 VNB N_A_213_23#_M1001_g 0.0242734f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_6 VNB N_A_213_23#_M1007_g 0.0222247f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.21
cc_7 VNB N_A_213_23#_M1008_g 0.0222366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_213_23#_M1012_g 0.0246709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_213_23#_c_104_n 0.00226813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_213_23#_c_105_n 0.0188925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_213_23#_c_106_n 0.0288914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_213_23#_c_107_n 0.00136909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_213_23#_c_108_n 0.0621182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_M1010_g 0.0245683f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.875
cc_15 VNB B 0.00338553f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_16 VNB N_B_c_216_n 0.0240692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_43_367#_M1011_g 0.0275272f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB N_A_43_367#_M1003_g 0.00155699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_43_367#_c_256_n 0.0321063f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.54
cc_20 VNB N_A_43_367#_c_257_n 0.00125038f $X=-0.19 $Y=-0.245 $X2=0.742 $Y2=1.665
cc_21 VNB N_A_43_367#_c_258_n 0.0141658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_43_367#_c_259_n 0.00626576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_43_367#_c_260_n 0.0503918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_322_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_382_n 0.0038636f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.375
cc_26 VNB N_X_c_383_n 0.00587307f $X=-0.19 $Y=-0.245 $X2=0.742 $Y2=1.295
cc_27 VNB N_X_c_384_n 0.00343442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_428_n 0.0176844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_429_n 0.0146736f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.375
cc_30 VNB N_VGND_c_430_n 4.97822e-19 $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.54
cc_31 VNB N_VGND_c_431_n 0.00534544f $X=-0.19 $Y=-0.245 $X2=0.742 $Y2=1.665
cc_32 VNB N_VGND_c_432_n 0.0248654f $X=-0.19 $Y=-0.245 $X2=0.742 $Y2=2.035
cc_33 VNB N_VGND_c_433_n 0.00577043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_434_n 0.01628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_435_n 0.0294792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_436_n 0.221299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_437_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_438_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A_N_M1004_g 0.0217837f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.045
cc_40 VPB A_N 0.00138518f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_41 VPB N_A_213_23#_M1000_g 0.0199637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_213_23#_M1002_g 0.0183015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_213_23#_M1005_g 0.0183181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_213_23#_M1013_g 0.0189301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_213_23#_c_113_n 0.00137855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_213_23#_c_108_n 0.0107978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B_M1009_g 0.0192007f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.045
cc_48 VPB B 0.0035141f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_49 VPB N_B_c_216_n 0.00616097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_43_367#_M1003_g 0.0226112f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_43_367#_c_256_n 0.0346904f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.54
cc_52 VPB N_A_43_367#_c_263_n 0.0199096f $X=-0.19 $Y=1.655 $X2=0.742 $Y2=1.295
cc_53 VPB N_A_43_367#_c_264_n 0.0126274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_43_367#_c_257_n 0.0284384f $X=-0.19 $Y=1.655 $X2=0.742 $Y2=1.665
cc_55 VPB N_VPWR_c_323_n 0.0150717f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.375
cc_56 VPB N_VPWR_c_324_n 0.0127282f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.21
cc_57 VPB N_VPWR_c_325_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_326_n 0.00431378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_327_n 0.0103375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_328_n 0.0159684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_329_n 0.0241178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_330_n 0.00510611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_331_n 0.0147575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_332_n 0.0148979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_333_n 0.00436638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_334_n 0.00631927f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_322_n 0.0543222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_X_c_382_n 0.0026621f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.375
cc_69 VPB X 0.00646855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 A_N N_A_213_23#_M1001_g 0.00332859f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_N_c_73_n N_A_213_23#_M1001_g 0.0214108f $X=0.69 $Y=1.375 $X2=0 $Y2=0
cc_72 N_A_N_c_74_n N_A_213_23#_M1001_g 0.0126207f $X=0.667 $Y=1.21 $X2=0 $Y2=0
cc_73 A_N N_A_213_23#_M1000_g 0.00142908f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_N_M1004_g N_A_213_23#_c_108_n 0.0213149f $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_75 A_N N_A_43_367#_c_256_n 0.0599817f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_N_c_73_n N_A_43_367#_c_256_n 0.0222126f $X=0.69 $Y=1.375 $X2=0 $Y2=0
cc_77 N_A_N_c_74_n N_A_43_367#_c_256_n 0.00460646f $X=0.667 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A_N_M1004_g N_A_43_367#_c_263_n 0.00678092f $X=0.555 $Y=2.045 $X2=0
+ $Y2=0
cc_79 A_N N_A_43_367#_c_263_n 0.0162397f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A_N_c_73_n N_A_43_367#_c_258_n 0.00147707f $X=0.69 $Y=1.375 $X2=0 $Y2=0
cc_81 N_A_N_c_74_n N_A_43_367#_c_258_n 0.00591014f $X=0.667 $Y=1.21 $X2=0 $Y2=0
cc_82 A_N N_VPWR_M1004_d 0.00720141f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_83 N_A_N_M1004_g N_X_c_382_n 8.32253e-19 $X=0.555 $Y=2.045 $X2=0 $Y2=0
cc_84 A_N N_X_c_382_n 0.0594263f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A_N_c_73_n N_X_c_382_n 8.60081e-19 $X=0.69 $Y=1.375 $X2=0 $Y2=0
cc_86 A_N N_X_c_384_n 0.00471398f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A_N_c_74_n N_X_c_384_n 0.00110154f $X=0.667 $Y=1.21 $X2=0 $Y2=0
cc_88 A_N N_VGND_c_428_n 0.00747239f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A_N_c_73_n N_VGND_c_428_n 6.69949e-19 $X=0.69 $Y=1.375 $X2=0 $Y2=0
cc_90 N_A_N_c_74_n N_VGND_c_428_n 0.00667924f $X=0.667 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A_N_c_74_n N_VGND_c_432_n 0.00380798f $X=0.667 $Y=1.21 $X2=0 $Y2=0
cc_92 N_A_N_c_74_n N_VGND_c_436_n 0.00458517f $X=0.667 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A_213_23#_M1013_g N_B_M1009_g 0.0410473f $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_213_23#_c_113_n N_B_M1009_g 0.00382031f $X=2.57 $Y=1.93 $X2=0 $Y2=0
cc_95 N_A_213_23#_c_122_p N_B_M1009_g 0.0134154f $X=3.15 $Y=2.095 $X2=0 $Y2=0
cc_96 N_A_213_23#_M1012_g N_B_M1010_g 0.0284863f $X=2.43 $Y=0.665 $X2=0 $Y2=0
cc_97 N_A_213_23#_c_104_n N_B_M1010_g 0.00353881f $X=2.57 $Y=1.415 $X2=0 $Y2=0
cc_98 N_A_213_23#_c_105_n N_B_M1010_g 0.0153021f $X=3.415 $Y=1.08 $X2=0 $Y2=0
cc_99 N_A_213_23#_c_106_n N_B_M1010_g 0.00248752f $X=3.58 $Y=0.39 $X2=0 $Y2=0
cc_100 N_A_213_23#_M1013_g B 2.23358e-19 $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A_213_23#_c_104_n B 0.00525729f $X=2.57 $Y=1.415 $X2=0 $Y2=0
cc_102 N_A_213_23#_c_113_n B 0.00906386f $X=2.57 $Y=1.93 $X2=0 $Y2=0
cc_103 N_A_213_23#_c_105_n B 0.0282218f $X=3.415 $Y=1.08 $X2=0 $Y2=0
cc_104 N_A_213_23#_c_122_p B 0.0274848f $X=3.15 $Y=2.095 $X2=0 $Y2=0
cc_105 N_A_213_23#_c_107_n B 0.0196961f $X=2.57 $Y=1.53 $X2=0 $Y2=0
cc_106 N_A_213_23#_c_108_n B 2.80915e-19 $X=2.43 $Y=1.51 $X2=0 $Y2=0
cc_107 N_A_213_23#_c_104_n N_B_c_216_n 4.87449e-19 $X=2.57 $Y=1.415 $X2=0 $Y2=0
cc_108 N_A_213_23#_c_113_n N_B_c_216_n 2.00321e-19 $X=2.57 $Y=1.93 $X2=0 $Y2=0
cc_109 N_A_213_23#_c_105_n N_B_c_216_n 0.00547352f $X=3.415 $Y=1.08 $X2=0 $Y2=0
cc_110 N_A_213_23#_c_122_p N_B_c_216_n 0.00274255f $X=3.15 $Y=2.095 $X2=0 $Y2=0
cc_111 N_A_213_23#_c_107_n N_B_c_216_n 0.00177963f $X=2.57 $Y=1.53 $X2=0 $Y2=0
cc_112 N_A_213_23#_c_108_n N_B_c_216_n 0.0168142f $X=2.43 $Y=1.51 $X2=0 $Y2=0
cc_113 N_A_213_23#_c_105_n N_A_43_367#_M1011_g 0.0159892f $X=3.415 $Y=1.08 $X2=0
+ $Y2=0
cc_114 N_A_213_23#_c_106_n N_A_43_367#_M1011_g 0.0161418f $X=3.58 $Y=0.39 $X2=0
+ $Y2=0
cc_115 N_A_213_23#_M1000_g N_A_43_367#_c_256_n 0.00137173f $X=1.14 $Y=2.465
+ $X2=0 $Y2=0
cc_116 N_A_213_23#_M1009_d N_A_43_367#_c_263_n 0.00494544f $X=3.01 $Y=1.835
+ $X2=0 $Y2=0
cc_117 N_A_213_23#_M1000_g N_A_43_367#_c_263_n 0.0151189f $X=1.14 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_213_23#_M1002_g N_A_43_367#_c_263_n 0.0129623f $X=1.57 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_A_213_23#_M1005_g N_A_43_367#_c_263_n 0.0129623f $X=2 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_213_23#_M1013_g N_A_43_367#_c_263_n 0.0168179f $X=2.43 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_A_213_23#_c_148_p N_A_43_367#_c_263_n 0.00982882f $X=2.66 $Y=2.095
+ $X2=0 $Y2=0
cc_122 N_A_213_23#_c_122_p N_A_43_367#_c_263_n 0.0343902f $X=3.15 $Y=2.095 $X2=0
+ $Y2=0
cc_123 N_A_213_23#_M1001_g N_A_43_367#_c_258_n 3.31931e-19 $X=1.14 $Y=0.665
+ $X2=0 $Y2=0
cc_124 N_A_213_23#_c_105_n N_A_43_367#_c_259_n 0.0222405f $X=3.415 $Y=1.08 $X2=0
+ $Y2=0
cc_125 N_A_213_23#_c_105_n N_A_43_367#_c_260_n 0.00691819f $X=3.415 $Y=1.08
+ $X2=0 $Y2=0
cc_126 N_A_213_23#_c_113_n N_VPWR_M1013_s 0.00112115f $X=2.57 $Y=1.93 $X2=0
+ $Y2=0
cc_127 N_A_213_23#_c_148_p N_VPWR_M1013_s 0.00107607f $X=2.66 $Y=2.095 $X2=0
+ $Y2=0
cc_128 N_A_213_23#_c_122_p N_VPWR_M1013_s 0.00593388f $X=3.15 $Y=2.095 $X2=0
+ $Y2=0
cc_129 N_A_213_23#_M1000_g N_VPWR_c_323_n 0.0105259f $X=1.14 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_A_213_23#_M1002_g N_VPWR_c_323_n 0.00135454f $X=1.57 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_A_213_23#_M1000_g N_VPWR_c_324_n 0.0036352f $X=1.14 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_A_213_23#_M1002_g N_VPWR_c_324_n 0.0036352f $X=1.57 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_213_23#_M1000_g N_VPWR_c_325_n 0.00135454f $X=1.14 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_213_23#_M1002_g N_VPWR_c_325_n 0.0094624f $X=1.57 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_213_23#_M1005_g N_VPWR_c_325_n 0.00970931f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_213_23#_M1013_g N_VPWR_c_325_n 0.00138138f $X=2.43 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A_213_23#_M1013_g N_VPWR_c_326_n 0.00173782f $X=2.43 $Y=2.465 $X2=0
+ $Y2=0
cc_138 N_A_213_23#_M1005_g N_VPWR_c_331_n 0.0036352f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_213_23#_M1013_g N_VPWR_c_331_n 0.00437171f $X=2.43 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_213_23#_M1009_d N_VPWR_c_322_n 0.00360572f $X=3.01 $Y=1.835 $X2=0
+ $Y2=0
cc_141 N_A_213_23#_M1000_g N_VPWR_c_322_n 0.00436741f $X=1.14 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_213_23#_M1002_g N_VPWR_c_322_n 0.00436741f $X=1.57 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_213_23#_M1005_g N_VPWR_c_322_n 0.00436741f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_213_23#_M1013_g N_VPWR_c_322_n 0.00611027f $X=2.43 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_213_23#_M1001_g N_X_c_382_n 0.00254024f $X=1.14 $Y=0.665 $X2=0 $Y2=0
cc_146 N_A_213_23#_M1000_g N_X_c_382_n 0.0134121f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_213_23#_M1007_g N_X_c_382_n 0.00209552f $X=1.57 $Y=0.665 $X2=0 $Y2=0
cc_148 N_A_213_23#_M1002_g N_X_c_382_n 0.00291707f $X=1.57 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_213_23#_c_176_p N_X_c_382_n 0.0149876f $X=2.48 $Y=1.53 $X2=0 $Y2=0
cc_150 N_A_213_23#_c_108_n N_X_c_382_n 0.0161945f $X=2.43 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A_213_23#_M1007_g N_X_c_383_n 0.0140947f $X=1.57 $Y=0.665 $X2=0 $Y2=0
cc_152 N_A_213_23#_M1008_g N_X_c_383_n 0.0137623f $X=2 $Y=0.665 $X2=0 $Y2=0
cc_153 N_A_213_23#_M1012_g N_X_c_383_n 0.00131418f $X=2.43 $Y=0.665 $X2=0 $Y2=0
cc_154 N_A_213_23#_c_176_p N_X_c_383_n 0.0601911f $X=2.48 $Y=1.53 $X2=0 $Y2=0
cc_155 N_A_213_23#_c_104_n N_X_c_383_n 0.00644339f $X=2.57 $Y=1.415 $X2=0 $Y2=0
cc_156 N_A_213_23#_c_183_p N_X_c_383_n 0.00750776f $X=2.66 $Y=1.08 $X2=0 $Y2=0
cc_157 N_A_213_23#_c_108_n N_X_c_383_n 0.00497162f $X=2.43 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A_213_23#_M1001_g N_X_c_384_n 0.0120984f $X=1.14 $Y=0.665 $X2=0 $Y2=0
cc_159 N_A_213_23#_c_108_n N_X_c_384_n 0.00289915f $X=2.43 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A_213_23#_M1002_g X 0.0135296f $X=1.57 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A_213_23#_M1005_g X 0.0135738f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_213_23#_c_176_p X 0.0608575f $X=2.48 $Y=1.53 $X2=0 $Y2=0
cc_163 N_A_213_23#_c_113_n X 0.00451261f $X=2.57 $Y=1.93 $X2=0 $Y2=0
cc_164 N_A_213_23#_c_108_n X 0.00758519f $X=2.43 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A_213_23#_c_105_n N_VGND_M1012_s 0.00262852f $X=3.415 $Y=1.08 $X2=0
+ $Y2=0
cc_166 N_A_213_23#_c_183_p N_VGND_M1012_s 0.00111107f $X=2.66 $Y=1.08 $X2=0
+ $Y2=0
cc_167 N_A_213_23#_M1001_g N_VGND_c_428_n 0.00337808f $X=1.14 $Y=0.665 $X2=0
+ $Y2=0
cc_168 N_A_213_23#_M1001_g N_VGND_c_429_n 0.00575161f $X=1.14 $Y=0.665 $X2=0
+ $Y2=0
cc_169 N_A_213_23#_M1007_g N_VGND_c_429_n 0.00477554f $X=1.57 $Y=0.665 $X2=0
+ $Y2=0
cc_170 N_A_213_23#_M1001_g N_VGND_c_430_n 6.24308e-19 $X=1.14 $Y=0.665 $X2=0
+ $Y2=0
cc_171 N_A_213_23#_M1007_g N_VGND_c_430_n 0.0109133f $X=1.57 $Y=0.665 $X2=0
+ $Y2=0
cc_172 N_A_213_23#_M1008_g N_VGND_c_430_n 0.0109964f $X=2 $Y=0.665 $X2=0 $Y2=0
cc_173 N_A_213_23#_M1012_g N_VGND_c_430_n 6.39121e-19 $X=2.43 $Y=0.665 $X2=0
+ $Y2=0
cc_174 N_A_213_23#_M1012_g N_VGND_c_431_n 0.00518289f $X=2.43 $Y=0.665 $X2=0
+ $Y2=0
cc_175 N_A_213_23#_c_105_n N_VGND_c_431_n 0.0165691f $X=3.415 $Y=1.08 $X2=0
+ $Y2=0
cc_176 N_A_213_23#_c_183_p N_VGND_c_431_n 0.00846382f $X=2.66 $Y=1.08 $X2=0
+ $Y2=0
cc_177 N_A_213_23#_M1008_g N_VGND_c_434_n 0.00477554f $X=2 $Y=0.665 $X2=0 $Y2=0
cc_178 N_A_213_23#_M1012_g N_VGND_c_434_n 0.00575161f $X=2.43 $Y=0.665 $X2=0
+ $Y2=0
cc_179 N_A_213_23#_c_106_n N_VGND_c_435_n 0.0210467f $X=3.58 $Y=0.39 $X2=0 $Y2=0
cc_180 N_A_213_23#_M1011_d N_VGND_c_436_n 0.00212301f $X=3.44 $Y=0.245 $X2=0
+ $Y2=0
cc_181 N_A_213_23#_M1001_g N_VGND_c_436_n 0.0118214f $X=1.14 $Y=0.665 $X2=0
+ $Y2=0
cc_182 N_A_213_23#_M1007_g N_VGND_c_436_n 0.00825815f $X=1.57 $Y=0.665 $X2=0
+ $Y2=0
cc_183 N_A_213_23#_M1008_g N_VGND_c_436_n 0.00825815f $X=2 $Y=0.665 $X2=0 $Y2=0
cc_184 N_A_213_23#_M1012_g N_VGND_c_436_n 0.0110121f $X=2.43 $Y=0.665 $X2=0
+ $Y2=0
cc_185 N_A_213_23#_c_106_n N_VGND_c_436_n 0.0125689f $X=3.58 $Y=0.39 $X2=0 $Y2=0
cc_186 N_A_213_23#_c_105_n A_616_49# 0.00366293f $X=3.415 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_187 N_B_M1010_g N_A_43_367#_M1011_g 0.0479726f $X=3.005 $Y=0.665 $X2=0 $Y2=0
cc_188 N_B_M1009_g N_A_43_367#_M1003_g 0.0522717f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_189 N_B_M1009_g N_A_43_367#_c_263_n 0.0129331f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_190 B N_A_43_367#_c_257_n 0.0105424f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_191 B N_A_43_367#_c_259_n 0.0135906f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_192 B N_A_43_367#_c_260_n 0.00409892f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_193 N_B_c_216_n N_A_43_367#_c_260_n 0.0479726f $X=2.915 $Y=1.51 $X2=0 $Y2=0
cc_194 N_B_M1009_g N_VPWR_c_326_n 0.00172188f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_195 N_B_M1009_g N_VPWR_c_328_n 0.00138516f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_196 N_B_M1009_g N_VPWR_c_332_n 0.00437171f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_197 N_B_M1009_g N_VPWR_c_322_n 0.00615122f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_198 N_B_M1010_g N_VGND_c_431_n 0.00651204f $X=3.005 $Y=0.665 $X2=0 $Y2=0
cc_199 N_B_M1010_g N_VGND_c_435_n 0.00575161f $X=3.005 $Y=0.665 $X2=0 $Y2=0
cc_200 N_B_M1010_g N_VGND_c_436_n 0.010916f $X=3.005 $Y=0.665 $X2=0 $Y2=0
cc_201 N_A_43_367#_c_263_n N_VPWR_M1004_d 0.00890352f $X=3.545 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A_43_367#_c_263_n N_VPWR_M1002_s 0.00396562f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_203 N_A_43_367#_c_263_n N_VPWR_M1013_s 0.00506026f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_204 N_A_43_367#_c_263_n N_VPWR_M1003_d 0.0048548f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_205 N_A_43_367#_c_257_n N_VPWR_M1003_d 0.0108081f $X=3.63 $Y=2.43 $X2=0 $Y2=0
cc_206 N_A_43_367#_c_263_n N_VPWR_c_323_n 0.021205f $X=3.545 $Y=2.52 $X2=0 $Y2=0
cc_207 N_A_43_367#_c_263_n N_VPWR_c_324_n 0.00670101f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_208 N_A_43_367#_c_263_n N_VPWR_c_325_n 0.0164573f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_209 N_A_43_367#_c_263_n N_VPWR_c_326_n 0.0188975f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_210 N_A_43_367#_M1003_g N_VPWR_c_328_n 0.0108072f $X=3.365 $Y=2.465 $X2=0
+ $Y2=0
cc_211 N_A_43_367#_c_263_n N_VPWR_c_328_n 0.0200712f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_212 N_A_43_367#_c_263_n N_VPWR_c_329_n 0.00514951f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_213 N_A_43_367#_c_264_n N_VPWR_c_329_n 0.00426603f $X=0.425 $Y=2.52 $X2=0
+ $Y2=0
cc_214 N_A_43_367#_c_263_n N_VPWR_c_331_n 0.00711846f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_215 N_A_43_367#_M1003_g N_VPWR_c_332_n 0.0036352f $X=3.365 $Y=2.465 $X2=0
+ $Y2=0
cc_216 N_A_43_367#_c_263_n N_VPWR_c_332_n 0.00715773f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_217 N_A_43_367#_M1003_g N_VPWR_c_322_n 0.00439469f $X=3.365 $Y=2.465 $X2=0
+ $Y2=0
cc_218 N_A_43_367#_c_263_n N_VPWR_c_322_n 0.0547224f $X=3.545 $Y=2.52 $X2=0
+ $Y2=0
cc_219 N_A_43_367#_c_264_n N_VPWR_c_322_n 0.00710942f $X=0.425 $Y=2.52 $X2=0
+ $Y2=0
cc_220 N_A_43_367#_c_263_n N_X_M1000_d 0.00541617f $X=3.545 $Y=2.52 $X2=0 $Y2=0
cc_221 N_A_43_367#_c_263_n N_X_M1005_d 0.00541648f $X=3.545 $Y=2.52 $X2=0 $Y2=0
cc_222 N_A_43_367#_c_263_n N_X_c_382_n 0.00827282f $X=3.545 $Y=2.52 $X2=0 $Y2=0
cc_223 N_A_43_367#_c_256_n N_X_c_384_n 0.00373998f $X=0.34 $Y=2.11 $X2=0 $Y2=0
cc_224 N_A_43_367#_c_263_n X 0.0396074f $X=3.545 $Y=2.52 $X2=0 $Y2=0
cc_225 N_A_43_367#_c_258_n N_VGND_c_428_n 0.0129726f $X=0.4 $Y=0.875 $X2=0 $Y2=0
cc_226 N_A_43_367#_c_258_n N_VGND_c_432_n 0.00555476f $X=0.4 $Y=0.875 $X2=0
+ $Y2=0
cc_227 N_A_43_367#_M1011_g N_VGND_c_435_n 0.00539298f $X=3.365 $Y=0.665 $X2=0
+ $Y2=0
cc_228 N_A_43_367#_M1011_g N_VGND_c_436_n 0.0107491f $X=3.365 $Y=0.665 $X2=0
+ $Y2=0
cc_229 N_A_43_367#_c_258_n N_VGND_c_436_n 0.0106454f $X=0.4 $Y=0.875 $X2=0 $Y2=0
cc_230 N_VPWR_c_322_n N_X_M1000_d 0.00360572f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_231 N_VPWR_c_322_n N_X_M1005_d 0.00360572f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_232 N_VPWR_M1002_s X 0.00228699f $X=1.645 $Y=1.835 $X2=0 $Y2=0
cc_233 N_X_c_383_n N_VGND_M1007_s 0.00180746f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_234 N_X_c_421_p N_VGND_c_429_n 0.0135169f $X=1.355 $Y=0.42 $X2=0 $Y2=0
cc_235 N_X_c_383_n N_VGND_c_430_n 0.0163515f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_236 N_X_c_423_p N_VGND_c_434_n 0.0124525f $X=2.215 $Y=0.42 $X2=0 $Y2=0
cc_237 N_X_M1001_d N_VGND_c_436_n 0.00432284f $X=1.215 $Y=0.245 $X2=0 $Y2=0
cc_238 N_X_M1008_d N_VGND_c_436_n 0.00536646f $X=2.075 $Y=0.245 $X2=0 $Y2=0
cc_239 N_X_c_421_p N_VGND_c_436_n 0.00847534f $X=1.355 $Y=0.42 $X2=0 $Y2=0
cc_240 N_X_c_423_p N_VGND_c_436_n 0.00730901f $X=2.215 $Y=0.42 $X2=0 $Y2=0
cc_241 N_VGND_c_436_n A_616_49# 0.00899413f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
