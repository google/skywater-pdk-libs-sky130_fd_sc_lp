* File: sky130_fd_sc_lp__or2b_2.pex.spice
* Created: Fri Aug 28 11:22:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2B_2%B_N 3 7 12 13 14 17 18
r27 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.04 $X2=0.385 $Y2=1.04
r28 14 18 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.21
+ $X2=0.385 $Y2=1.21
r29 12 17 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.385 $Y=1.395
+ $X2=0.385 $Y2=1.04
r30 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.417 $Y=1.395
+ $X2=0.417 $Y2=1.545
r31 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=0.875
+ $X2=0.385 $Y2=1.04
r32 7 13 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.54 $Y=2.045 $X2=0.54
+ $Y2=1.545
r33 3 10 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.475 $Y=0.455
+ $X2=0.475 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_2%A_191_254# 1 2 9 11 13 16 18 20 24 26 28 30
+ 31 32 40
r81 39 40 5.15902 $w=3.27e-07 $l=3.5e-08 $layer=POLY_cond $X=1.46 $Y=1.36
+ $X2=1.495 $Y2=1.36
r82 38 39 58.2232 $w=3.27e-07 $l=3.95e-07 $layer=POLY_cond $X=1.065 $Y=1.36
+ $X2=1.46 $Y2=1.36
r83 37 38 5.15902 $w=3.27e-07 $l=3.5e-08 $layer=POLY_cond $X=1.03 $Y=1.36
+ $X2=1.065 $Y2=1.36
r84 32 35 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.895 $Y=2.015
+ $X2=2.895 $Y2=2.095
r85 30 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=2.015
+ $X2=2.895 $Y2=2.015
r86 30 31 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.73 $Y=2.015 $X2=1.83
+ $Y2=2.015
r87 26 28 23.2705 $w=2.58e-07 $l=5.25e-07 $layer=LI1_cond $X=1.83 $Y=0.995
+ $X2=2.355 $Y2=0.995
r88 25 40 25.0581 $w=3.27e-07 $l=1.7e-07 $layer=POLY_cond $X=1.665 $Y=1.36
+ $X2=1.495 $Y2=1.36
r89 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.665
+ $Y=1.36 $X2=1.665 $Y2=1.36
r90 22 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.705 $Y=1.93
+ $X2=1.83 $Y2=2.015
r91 22 24 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=1.705 $Y=1.93
+ $X2=1.705 $Y2=1.36
r92 21 26 4.55389 $w=3.81e-07 $l=3.41833e-07 $layer=LI1_cond $X=1.705 $Y=1.28
+ $X2=1.83 $Y2=0.995
r93 21 24 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.705 $Y=1.28
+ $X2=1.705 $Y2=1.36
r94 18 40 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.195
+ $X2=1.495 $Y2=1.36
r95 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.495 $Y=1.195
+ $X2=1.495 $Y2=0.665
r96 14 39 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.46 $Y=1.525
+ $X2=1.46 $Y2=1.36
r97 14 16 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.46 $Y=1.525 $X2=1.46
+ $Y2=2.465
r98 11 38 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.195
+ $X2=1.065 $Y2=1.36
r99 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.065 $Y=1.195
+ $X2=1.065 $Y2=0.665
r100 7 37 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.525
+ $X2=1.03 $Y2=1.36
r101 7 9 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.03 $Y=1.525 $X2=1.03
+ $Y2=2.465
r102 2 35 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=1.835 $X2=2.895 $Y2=2.095
r103 1 28 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.665 $X2=2.355 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_2%A 3 7 9 10 14
c37 3 0 1.10516e-19 $X=2.14 $Y=0.875
r38 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.51
+ $X2=2.23 $Y2=1.675
r39 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.51
+ $X2=2.23 $Y2=1.345
r40 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.51 $X2=2.23 $Y2=1.51
r41 10 15 13.6957 $w=3.43e-07 $l=4.1e-07 $layer=LI1_cond $X=2.64 $Y=1.587
+ $X2=2.23 $Y2=1.587
r42 9 15 2.33829 $w=3.43e-07 $l=7e-08 $layer=LI1_cond $X=2.16 $Y=1.587 $X2=2.23
+ $Y2=1.587
r43 7 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.32 $Y=2.045
+ $X2=2.32 $Y2=1.675
r44 3 16 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.14 $Y=0.875 $X2=2.14
+ $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_2%A_27_49# 1 2 7 9 12 15 16 19 20 23 25 30 32
+ 35 39
r83 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.47
+ $Y=1.36 $X2=3.47 $Y2=1.36
r84 36 39 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=3.03 $Y=1.36 $X2=3.47
+ $Y2=1.36
r85 35 38 14.3529 $w=3.74e-07 $l=4.4e-07 $layer=LI1_cond $X=3.03 $Y=1.3 $X2=3.47
+ $Y2=1.3
r86 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=1.36 $X2=3.03 $Y2=1.36
r87 25 27 5.49627 $w=3.23e-07 $l=1.55e-07 $layer=LI1_cond $X=0.257 $Y=0.455
+ $X2=0.257 $Y2=0.61
r88 23 35 8.31818 $w=3.74e-07 $l=3.49857e-07 $layer=LI1_cond $X=2.775 $Y=1.075
+ $X2=3.03 $Y2=1.3
r89 22 23 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.775 $Y=0.695
+ $X2=2.775 $Y2=1.075
r90 21 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=0.61
+ $X2=0.735 $Y2=0.61
r91 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.69 $Y=0.61
+ $X2=2.775 $Y2=0.695
r92 20 21 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=2.69 $Y=0.61 $X2=0.82
+ $Y2=0.61
r93 19 30 15.0663 $w=3.32e-07 $l=5.19009e-07 $layer=LI1_cond $X=0.735 $Y=1.715
+ $X2=0.325 $Y2=1.962
r94 18 32 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.695
+ $X2=0.735 $Y2=0.61
r95 18 19 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.735 $Y=0.695
+ $X2=0.735 $Y2=1.715
r96 17 27 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=0.42 $Y=0.61
+ $X2=0.257 $Y2=0.61
r97 16 32 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=0.61
+ $X2=0.735 $Y2=0.61
r98 16 17 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.65 $Y=0.61
+ $X2=0.42 $Y2=0.61
r99 14 36 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=2.755 $Y=1.36
+ $X2=3.03 $Y2=1.36
r100 14 15 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.755 $Y=1.36
+ $X2=2.68 $Y2=1.36
r101 10 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.525
+ $X2=2.68 $Y2=1.36
r102 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.68 $Y=1.525
+ $X2=2.68 $Y2=2.045
r103 7 15 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.195
+ $X2=2.68 $Y2=1.36
r104 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.68 $Y=1.195
+ $X2=2.68 $Y2=0.875
r105 2 30 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.835 $X2=0.325 $Y2=2.045
r106 1 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.245 $X2=0.26 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_2%VPWR 1 2 11 17 19 21 31 32 35 38
r26 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r29 29 32 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r30 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r31 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 26 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.84 $Y=3.33 $X2=1.71
+ $Y2=3.33
r33 26 28 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.84 $Y=3.33 $X2=2.16
+ $Y2=3.33
r34 25 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 25 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r37 22 35 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.797 $Y2=3.33
r38 22 24 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33 $X2=1.2
+ $Y2=3.33
r39 21 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.58 $Y=3.33 $X2=1.71
+ $Y2=3.33
r40 21 24 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.58 $Y=3.33 $X2=1.2
+ $Y2=3.33
r41 19 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 19 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 15 38 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=3.33
r44 15 17 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=2.435
r45 11 14 37.3904 $w=2.23e-07 $l=7.3e-07 $layer=LI1_cond $X=0.797 $Y=2.22
+ $X2=0.797 $Y2=2.95
r46 9 35 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.797 $Y=3.245
+ $X2=0.797 $Y2=3.33
r47 9 14 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=0.797 $Y=3.245
+ $X2=0.797 $Y2=2.95
r48 2 17 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=1.835 $X2=1.675 $Y2=2.435
r49 1 14 400 $w=1.7e-07 $l=1.21088e-06 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.835 $X2=0.815 $Y2=2.95
r50 1 11 400 $w=1.7e-07 $l=4.74579e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.835 $X2=0.815 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_2%X 1 2 9 12 13 14 15 16
c19 9 0 1.10516e-19 $X=1.28 $Y=0.96
r20 16 34 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.245 $Y=2.775
+ $X2=1.245 $Y2=2.91
r21 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.245 $Y=2.405
+ $X2=1.245 $Y2=2.775
r22 14 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.245 $Y=1.96
+ $X2=1.245 $Y2=2.405
r23 13 14 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.245 $Y=1.665
+ $X2=1.245 $Y2=1.96
r24 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.245 $Y=1.295
+ $X2=1.245 $Y2=1.665
r25 11 12 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.245 $Y=1.045
+ $X2=1.245 $Y2=1.295
r26 9 11 2.8139 $w=3.63e-07 $l=8.5e-08 $layer=LI1_cond $X=1.262 $Y=0.96
+ $X2=1.262 $Y2=1.045
r27 2 34 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.835 $X2=1.245 $Y2=2.91
r28 2 14 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.835 $X2=1.245 $Y2=1.96
r29 1 9 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.245 $X2=1.28 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_2%VGND 1 2 3 10 14 16 18 23 30 31 42 48
r46 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 42 45 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=1.79 $Y=0 $X2=1.79
+ $Y2=0.26
r48 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r49 36 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r50 31 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r51 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r52 28 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.195
+ $Y2=0
r53 28 30 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r54 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r55 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r56 24 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=1.79
+ $Y2=0
r57 24 26 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=2.64
+ $Y2=0
r58 23 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=3.195
+ $Y2=0
r59 23 26 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.64
+ $Y2=0
r60 21 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r61 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r62 18 38 8.68508 $w=3.43e-07 $l=2.6e-07 $layer=LI1_cond $X=0.762 $Y=0 $X2=0.762
+ $Y2=0.26
r63 18 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r64 18 20 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.59 $Y=0 $X2=0.24
+ $Y2=0
r65 16 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r66 16 43 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r67 12 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=0.085
+ $X2=3.195 $Y2=0
r68 12 14 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=3.195 $Y=0.085
+ $X2=3.195 $Y2=0.81
r69 11 18 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.762
+ $Y2=0
r70 10 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.79
+ $Y2=0
r71 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=0.935
+ $Y2=0
r72 3 14 182 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.665 $X2=3.195 $Y2=0.81
r73 2 45 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.245 $X2=1.79 $Y2=0.26
r74 1 38 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.245 $X2=0.77 $Y2=0.26
.ends

