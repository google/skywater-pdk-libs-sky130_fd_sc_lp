* File: sky130_fd_sc_lp__a32o_4.pex.spice
* Created: Fri Aug 28 10:01:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32O_4%A_101_21# 1 2 3 4 15 19 23 27 31 35 39 43 45
+ 51 53 54 58 60 63 68 70 77 78 79 80 82 84 95
c183 80 0 3.17863e-20 $X=6.507 $Y=1.09
c184 78 0 5.60522e-20 $X=4.52 $Y=1.17
c185 63 0 4.33649e-20 $X=6.345 $Y=1.92
r186 92 93 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.62 $Y=1.48
+ $X2=1.87 $Y2=1.48
r187 91 92 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.44 $Y=1.48
+ $X2=1.62 $Y2=1.48
r188 90 91 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.19 $Y=1.48
+ $X2=1.44 $Y2=1.48
r189 89 90 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.01 $Y=1.48
+ $X2=1.19 $Y2=1.48
r190 88 89 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.76 $Y=1.48
+ $X2=1.01 $Y2=1.48
r191 77 78 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=4.35 $Y=1.17
+ $X2=4.52 $Y2=1.17
r192 76 95 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.03 $Y=1.48 $X2=2.05
+ $Y2=1.48
r193 76 93 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.03 $Y=1.48
+ $X2=1.87 $Y2=1.48
r194 75 76 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.03
+ $Y=1.48 $X2=2.03 $Y2=1.48
r195 71 82 2.23839 $w=1.8e-07 $l=1.4e-07 $layer=LI1_cond $X=6.535 $Y=2.01
+ $X2=6.395 $Y2=2.01
r196 70 84 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.28 $Y=2.01
+ $X2=7.445 $Y2=2.01
r197 70 71 45.904 $w=1.78e-07 $l=7.45e-07 $layer=LI1_cond $X=7.28 $Y=2.01
+ $X2=6.535 $Y2=2.01
r198 66 80 3.64284 $w=2.55e-07 $l=1.23386e-07 $layer=LI1_cond $X=6.595 $Y=1.005
+ $X2=6.507 $Y2=1.09
r199 66 68 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6.595 $Y=1.005
+ $X2=6.595 $Y2=0.685
r200 63 82 4.19361 $w=2.3e-07 $l=1.1225e-07 $layer=LI1_cond $X=6.345 $Y=1.92
+ $X2=6.395 $Y2=2.01
r201 62 80 3.64284 $w=2.55e-07 $l=2.00035e-07 $layer=LI1_cond $X=6.345 $Y=1.175
+ $X2=6.507 $Y2=1.09
r202 62 63 45.904 $w=1.78e-07 $l=7.45e-07 $layer=LI1_cond $X=6.345 $Y=1.175
+ $X2=6.345 $Y2=1.92
r203 61 79 6.92067 $w=1.7e-07 $l=2.84341e-07 $layer=LI1_cond $X=5.31 $Y=1.09
+ $X2=5.065 $Y2=1.005
r204 60 80 2.83584 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=6.255 $Y=1.09
+ $X2=6.507 $Y2=1.09
r205 60 61 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=6.255 $Y=1.09
+ $X2=5.31 $Y2=1.09
r206 56 79 0.066131 $w=2.45e-07 $l=1.22e-07 $layer=LI1_cond $X=5.187 $Y=1.005
+ $X2=5.065 $Y2=1.005
r207 56 58 10.5837 $w=2.43e-07 $l=2.25e-07 $layer=LI1_cond $X=5.187 $Y=1.005
+ $X2=5.187 $Y2=0.78
r208 54 79 6.92067 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=5.065 $Y=1.18
+ $X2=5.065 $Y2=1.005
r209 54 78 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.065 $Y=1.18
+ $X2=4.52 $Y2=1.18
r210 53 77 140.594 $w=1.68e-07 $l=2.155e-06 $layer=LI1_cond $X=2.195 $Y=1.16
+ $X2=4.35 $Y2=1.16
r211 51 75 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.11 $Y=1.385 $X2=2.11
+ $Y2=1.485
r212 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=1.245
+ $X2=2.195 $Y2=1.16
r213 50 51 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.11 $Y=1.245
+ $X2=2.11 $Y2=1.385
r214 48 88 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.67 $Y=1.48 $X2=0.76
+ $Y2=1.48
r215 48 85 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.67 $Y=1.48 $X2=0.58
+ $Y2=1.48
r216 47 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.67
+ $Y=1.48 $X2=0.67 $Y2=1.48
r217 45 75 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=1.485
+ $X2=2.11 $Y2=1.485
r218 45 47 75.1409 $w=1.98e-07 $l=1.355e-06 $layer=LI1_cond $X=2.025 $Y=1.485
+ $X2=0.67 $Y2=1.485
r219 41 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.645
+ $X2=2.05 $Y2=1.48
r220 41 43 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.05 $Y=1.645
+ $X2=2.05 $Y2=2.465
r221 37 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.315
+ $X2=1.87 $Y2=1.48
r222 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.87 $Y=1.315
+ $X2=1.87 $Y2=0.655
r223 33 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.645
+ $X2=1.62 $Y2=1.48
r224 33 35 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.62 $Y=1.645
+ $X2=1.62 $Y2=2.465
r225 29 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.44 $Y=1.315
+ $X2=1.44 $Y2=1.48
r226 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.44 $Y=1.315
+ $X2=1.44 $Y2=0.655
r227 25 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.645
+ $X2=1.19 $Y2=1.48
r228 25 27 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.19 $Y=1.645
+ $X2=1.19 $Y2=2.465
r229 21 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.315
+ $X2=1.01 $Y2=1.48
r230 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.01 $Y=1.315
+ $X2=1.01 $Y2=0.655
r231 17 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.76 $Y=1.645
+ $X2=0.76 $Y2=1.48
r232 17 19 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.76 $Y=1.645
+ $X2=0.76 $Y2=2.465
r233 13 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.315
+ $X2=0.58 $Y2=1.48
r234 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.58 $Y=1.315
+ $X2=0.58 $Y2=0.655
r235 4 84 300 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=2 $X=7.305
+ $Y=1.835 $X2=7.445 $Y2=2.035
r236 3 82 300 $w=1.7e-07 $l=3.28481e-07 $layer=licon1_PDIFF $count=2 $X=6.215
+ $Y=1.835 $X2=6.37 $Y2=2.095
r237 2 68 91 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_NDIFF $count=2 $X=6.455
+ $Y=0.325 $X2=6.595 $Y2=0.685
r238 1 58 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=5.075
+ $Y=0.235 $X2=5.215 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%A3 3 7 11 15 17 18 26
r51 24 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.82 $Y=1.51 $X2=2.91
+ $Y2=1.51
r52 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.51 $X2=2.82 $Y2=1.51
r53 21 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.48 $Y=1.51
+ $X2=2.82 $Y2=1.51
r54 18 25 10.6379 $w=3.23e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.587 $X2=2.82
+ $Y2=1.587
r55 17 25 6.38276 $w=3.23e-07 $l=1.8e-07 $layer=LI1_cond $X=2.64 $Y=1.587
+ $X2=2.82 $Y2=1.587
r56 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.91 $Y=1.675
+ $X2=2.91 $Y2=1.51
r57 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.91 $Y=1.675
+ $X2=2.91 $Y2=2.465
r58 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.91 $Y=1.345
+ $X2=2.91 $Y2=1.51
r59 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.91 $Y=1.345
+ $X2=2.91 $Y2=0.655
r60 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.48 $Y=1.675
+ $X2=2.48 $Y2=1.51
r61 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.48 $Y=1.675 $X2=2.48
+ $Y2=2.465
r62 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.48 $Y=1.345
+ $X2=2.48 $Y2=1.51
r63 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.48 $Y=1.345 $X2=2.48
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%A2 3 5 7 10 12 14 15 18 20 21
r54 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.005
+ $Y=1.51 $X2=4.005 $Y2=1.51
r55 21 26 2.5801 $w=3.33e-07 $l=7.5e-08 $layer=LI1_cond $X=4.08 $Y=1.582
+ $X2=4.005 $Y2=1.582
r56 20 26 13.9325 $w=3.33e-07 $l=4.05e-07 $layer=LI1_cond $X=3.6 $Y=1.582
+ $X2=4.005 $Y2=1.582
r57 17 18 32.0316 $w=3.16e-07 $l=2.1e-07 $layer=POLY_cond $X=4.36 $Y=1.535
+ $X2=4.57 $Y2=1.535
r58 16 17 33.557 $w=3.16e-07 $l=2.2e-07 $layer=POLY_cond $X=4.14 $Y=1.535
+ $X2=4.36 $Y2=1.535
r59 15 25 8.78138 $w=3.8e-07 $l=6e-08 $layer=POLY_cond $X=4.065 $Y=1.535
+ $X2=4.005 $Y2=1.535
r60 15 16 11.0227 $w=3.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.065 $Y=1.535
+ $X2=4.14 $Y2=1.535
r61 12 18 33.557 $w=3.16e-07 $l=3.00333e-07 $layer=POLY_cond $X=4.79 $Y=1.725
+ $X2=4.57 $Y2=1.535
r62 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.79 $Y=1.725
+ $X2=4.79 $Y2=2.465
r63 8 18 20.1942 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.57 $Y=1.345
+ $X2=4.57 $Y2=1.535
r64 8 10 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.57 $Y=1.345
+ $X2=4.57 $Y2=0.655
r65 5 17 20.1942 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.36 $Y=1.725
+ $X2=4.36 $Y2=1.535
r66 5 7 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.36 $Y=1.725 $X2=4.36
+ $Y2=2.465
r67 1 16 20.1942 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.14 $Y=1.345
+ $X2=4.14 $Y2=1.535
r68 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.14 $Y=1.345 $X2=4.14
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%A1 1 3 6 8 10 13 15 16 23 26
c58 13 0 4.33649e-20 $X=5.71 $Y=2.465
c59 1 0 5.60522e-20 $X=5 $Y=1.185
r60 24 26 1.40044 $w=3.93e-07 $l=4.8e-08 $layer=LI1_cond $X=5.67 $Y=1.552
+ $X2=5.622 $Y2=1.552
r61 23 25 5.44633 $w=3.54e-07 $l=4e-08 $layer=POLY_cond $X=5.67 $Y=1.395
+ $X2=5.71 $Y2=1.395
r62 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.67
+ $Y=1.44 $X2=5.67 $Y2=1.44
r63 21 23 32.678 $w=3.54e-07 $l=2.4e-07 $layer=POLY_cond $X=5.43 $Y=1.395
+ $X2=5.67 $Y2=1.395
r64 20 21 28.5932 $w=3.54e-07 $l=2.1e-07 $layer=POLY_cond $X=5.22 $Y=1.395
+ $X2=5.43 $Y2=1.395
r65 16 24 9.62801 $w=3.93e-07 $l=3.3e-07 $layer=LI1_cond $X=6 $Y=1.552 $X2=5.67
+ $Y2=1.552
r66 15 26 3.33842 $w=3.95e-07 $l=1.02e-07 $layer=LI1_cond $X=5.52 $Y=1.552
+ $X2=5.622 $Y2=1.552
r67 11 25 22.9014 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.71 $Y=1.605
+ $X2=5.71 $Y2=1.395
r68 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.71 $Y=1.605
+ $X2=5.71 $Y2=2.465
r69 8 21 22.9014 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.43 $Y=1.185
+ $X2=5.43 $Y2=1.395
r70 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.43 $Y=1.185
+ $X2=5.43 $Y2=0.655
r71 4 20 22.9014 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.22 $Y=1.605
+ $X2=5.22 $Y2=1.395
r72 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.22 $Y=1.605 $X2=5.22
+ $Y2=2.465
r73 1 20 29.9548 $w=3.54e-07 $l=3.07571e-07 $layer=POLY_cond $X=5 $Y=1.185
+ $X2=5.22 $Y2=1.395
r74 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5 $Y=1.185 $X2=5
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%B1 3 7 11 15 17 26
c58 11 0 1.15065e-19 $X=6.65 $Y=2.465
r59 24 26 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.78 $Y=1.51 $X2=6.81
+ $Y2=1.51
r60 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.78
+ $Y=1.51 $X2=6.78 $Y2=1.51
r61 22 24 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=6.65 $Y=1.51 $X2=6.78
+ $Y2=1.51
r62 21 22 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=6.38 $Y=1.51
+ $X2=6.65 $Y2=1.51
r63 19 21 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=6.14 $Y=1.51
+ $X2=6.38 $Y2=1.51
r64 17 25 6.38276 $w=3.23e-07 $l=1.8e-07 $layer=LI1_cond $X=6.96 $Y=1.587
+ $X2=6.78 $Y2=1.587
r65 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.81 $Y=1.345
+ $X2=6.81 $Y2=1.51
r66 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.81 $Y=1.345 $X2=6.81
+ $Y2=0.745
r67 9 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.65 $Y=1.675
+ $X2=6.65 $Y2=1.51
r68 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.65 $Y=1.675
+ $X2=6.65 $Y2=2.465
r69 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.38 $Y=1.345
+ $X2=6.38 $Y2=1.51
r70 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.38 $Y=1.345 $X2=6.38
+ $Y2=0.745
r71 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.14 $Y=1.675
+ $X2=6.14 $Y2=1.51
r72 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.14 $Y=1.675 $X2=6.14
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%B2 3 7 11 15 17 18 26
c38 7 0 3.17863e-20 $X=7.24 $Y=0.745
r39 26 27 1.47853 $w=3.26e-07 $l=1e-08 $layer=POLY_cond $X=7.66 $Y=1.51 $X2=7.67
+ $Y2=1.51
r40 24 26 20.6994 $w=3.26e-07 $l=1.4e-07 $layer=POLY_cond $X=7.52 $Y=1.51
+ $X2=7.66 $Y2=1.51
r41 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.52
+ $Y=1.51 $X2=7.52 $Y2=1.51
r42 22 24 41.3988 $w=3.26e-07 $l=2.8e-07 $layer=POLY_cond $X=7.24 $Y=1.51
+ $X2=7.52 $Y2=1.51
r43 21 22 1.47853 $w=3.26e-07 $l=1e-08 $layer=POLY_cond $X=7.23 $Y=1.51 $X2=7.24
+ $Y2=1.51
r44 18 25 14.1839 $w=3.23e-07 $l=4e-07 $layer=LI1_cond $X=7.92 $Y=1.587 $X2=7.52
+ $Y2=1.587
r45 17 25 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=7.44 $Y=1.587 $X2=7.52
+ $Y2=1.587
r46 13 27 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=1.345
+ $X2=7.67 $Y2=1.51
r47 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.67 $Y=1.345 $X2=7.67
+ $Y2=0.745
r48 9 26 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.66 $Y=1.675
+ $X2=7.66 $Y2=1.51
r49 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.66 $Y=1.675
+ $X2=7.66 $Y2=2.465
r50 5 22 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.24 $Y=1.345
+ $X2=7.24 $Y2=1.51
r51 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.24 $Y=1.345 $X2=7.24
+ $Y2=0.745
r52 1 21 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.23 $Y=1.675
+ $X2=7.23 $Y2=1.51
r53 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.23 $Y=1.675 $X2=7.23
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%VPWR 1 2 3 4 5 6 21 27 31 35 41 45 49 52 53
+ 54 55 56 65 70 75 82 83 86 89 92 95
r110 95 96 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r111 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r113 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r114 83 96 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=5.52 $Y2=3.33
r115 82 83 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r116 80 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.6 $Y=3.33
+ $X2=5.435 $Y2=3.33
r117 80 82 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=5.6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 79 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 79 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r120 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r121 76 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=3.33
+ $X2=4.575 $Y2=3.33
r122 76 78 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.74 $Y=3.33 $X2=5.04
+ $Y2=3.33
r123 75 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.435 $Y2=3.33
r124 75 78 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 71 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=3.33
+ $X2=3.125 $Y2=3.33
r126 71 73 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.29 $Y=3.33
+ $X2=4.08 $Y2=3.33
r127 70 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.41 $Y=3.33
+ $X2=4.575 $Y2=3.33
r128 70 73 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.41 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 69 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r130 69 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r131 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r132 66 86 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.255 $Y2=3.33
r133 66 68 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.64 $Y2=3.33
r134 65 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.96 $Y=3.33
+ $X2=3.125 $Y2=3.33
r135 65 68 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.96 $Y=3.33
+ $X2=2.64 $Y2=3.33
r136 64 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 60 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r139 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r140 56 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r141 56 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r142 56 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r143 54 63 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r144 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=3.33
+ $X2=1.405 $Y2=3.33
r145 52 59 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.24 $Y2=3.33
r146 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.545 $Y2=3.33
r147 51 63 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=0.71 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=3.33
+ $X2=0.545 $Y2=3.33
r149 47 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=3.245
+ $X2=5.435 $Y2=3.33
r150 47 49 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=5.435 $Y=3.245
+ $X2=5.435 $Y2=2.375
r151 43 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=3.245
+ $X2=4.575 $Y2=3.33
r152 43 45 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=4.575 $Y=3.245
+ $X2=4.575 $Y2=2.375
r153 39 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=3.245
+ $X2=3.125 $Y2=3.33
r154 39 41 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3.125 $Y=3.245
+ $X2=3.125 $Y2=2.375
r155 35 38 48.603 $w=2.28e-07 $l=9.7e-07 $layer=LI1_cond $X=2.255 $Y=1.98
+ $X2=2.255 $Y2=2.95
r156 33 86 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=3.245
+ $X2=2.255 $Y2=3.33
r157 33 38 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.255 $Y=3.245
+ $X2=2.255 $Y2=2.95
r158 32 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=1.405 $Y2=3.33
r159 31 86 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.14 $Y=3.33
+ $X2=2.255 $Y2=3.33
r160 31 32 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.14 $Y=3.33
+ $X2=1.57 $Y2=3.33
r161 27 30 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.405 $Y=2.18
+ $X2=1.405 $Y2=2.95
r162 25 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.405 $Y=3.245
+ $X2=1.405 $Y2=3.33
r163 25 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.405 $Y=3.245
+ $X2=1.405 $Y2=2.95
r164 21 24 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.545 $Y=2.18
+ $X2=0.545 $Y2=2.95
r165 19 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.545 $Y=3.245
+ $X2=0.545 $Y2=3.33
r166 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.545 $Y=3.245
+ $X2=0.545 $Y2=2.95
r167 6 49 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=5.295
+ $Y=1.835 $X2=5.435 $Y2=2.375
r168 5 45 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=4.435
+ $Y=1.835 $X2=4.575 $Y2=2.375
r169 4 41 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.835 $X2=3.125 $Y2=2.375
r170 3 38 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=1.835 $X2=2.265 $Y2=2.95
r171 3 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=1.835 $X2=2.265 $Y2=1.98
r172 2 30 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=1.835 $X2=1.405 $Y2=2.95
r173 2 27 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=1.835 $X2=1.405 $Y2=2.18
r174 1 24 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.42
+ $Y=1.835 $X2=0.545 $Y2=2.95
r175 1 21 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.42
+ $Y=1.835 $X2=0.545 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%X 1 2 3 4 13 15 16 19 23 27 29 33 37 42 43 44
+ 45 49 51
r61 49 51 3.92321 $w=2.33e-07 $l=8e-08 $layer=LI1_cond $X=0.217 $Y=1.215
+ $X2=0.217 $Y2=1.295
r62 44 49 2.95087 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=1.13
+ $X2=0.217 $Y2=1.215
r63 44 45 18.0468 $w=2.33e-07 $l=3.68e-07 $layer=LI1_cond $X=0.217 $Y=1.297
+ $X2=0.217 $Y2=1.665
r64 44 51 0.0980803 $w=2.33e-07 $l=2e-09 $layer=LI1_cond $X=0.217 $Y=1.297
+ $X2=0.217 $Y2=1.295
r65 41 45 4.41361 $w=2.33e-07 $l=9e-08 $layer=LI1_cond $X=0.217 $Y=1.755
+ $X2=0.217 $Y2=1.665
r66 37 39 46.5988 $w=2.28e-07 $l=9.3e-07 $layer=LI1_cond $X=1.855 $Y=1.98
+ $X2=1.855 $Y2=2.91
r67 35 37 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.855 $Y=1.925
+ $X2=1.855 $Y2=1.98
r68 31 33 27.703 $w=2.58e-07 $l=6.25e-07 $layer=LI1_cond $X=1.69 $Y=1.045
+ $X2=1.69 $Y2=0.42
r69 30 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.07 $Y=1.84
+ $X2=0.975 $Y2=1.84
r70 29 35 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.74 $Y=1.84
+ $X2=1.855 $Y2=1.925
r71 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.74 $Y=1.84
+ $X2=1.07 $Y2=1.84
r72 28 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.89 $Y=1.13
+ $X2=0.795 $Y2=1.13
r73 27 31 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.56 $Y=1.13
+ $X2=1.69 $Y2=1.045
r74 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.56 $Y=1.13
+ $X2=0.89 $Y2=1.13
r75 23 25 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.975 $Y=1.98
+ $X2=0.975 $Y2=2.91
r76 21 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=1.925
+ $X2=0.975 $Y2=1.84
r77 21 23 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=0.975 $Y=1.925
+ $X2=0.975 $Y2=1.98
r78 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=1.045
+ $X2=0.795 $Y2=1.13
r79 17 19 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=0.795 $Y=1.045
+ $X2=0.795 $Y2=0.42
r80 16 41 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.335 $Y=1.84
+ $X2=0.217 $Y2=1.755
r81 15 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.88 $Y=1.84
+ $X2=0.975 $Y2=1.84
r82 15 16 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=0.88 $Y=1.84
+ $X2=0.335 $Y2=1.84
r83 14 44 4.0965 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=0.335 $Y=1.13
+ $X2=0.217 $Y2=1.13
r84 13 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.7 $Y=1.13 $X2=0.795
+ $Y2=1.13
r85 13 14 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.7 $Y=1.13
+ $X2=0.335 $Y2=1.13
r86 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.695
+ $Y=1.835 $X2=1.835 $Y2=2.91
r87 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.695
+ $Y=1.835 $X2=1.835 $Y2=1.98
r88 3 25 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.835
+ $Y=1.835 $X2=0.975 $Y2=2.91
r89 3 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.835
+ $Y=1.835 $X2=0.975 $Y2=1.98
r90 2 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.235 $X2=1.655 $Y2=0.42
r91 1 19 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.655
+ $Y=0.235 $X2=0.795 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%A_511_367# 1 2 3 4 5 6 19 21 23 27 29 33 35
+ 37 38 39 43 45 47 49 54 56 61
c80 37 0 1.15065e-19 $X=5.927 $Y=2.09
r81 47 63 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=2.905
+ $X2=7.91 $Y2=2.99
r82 47 49 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=7.91 $Y=2.905
+ $X2=7.91 $Y2=2.085
r83 46 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.105 $Y=2.99
+ $X2=6.94 $Y2=2.99
r84 45 63 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.78 $Y=2.99 $X2=7.91
+ $Y2=2.99
r85 45 46 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.78 $Y=2.99
+ $X2=7.105 $Y2=2.99
r86 41 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.94 $Y=2.905
+ $X2=6.94 $Y2=2.99
r87 41 43 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=6.94 $Y=2.905
+ $X2=6.94 $Y2=2.38
r88 40 60 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=6.085 $Y=2.99
+ $X2=5.927 $Y2=2.99
r89 39 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=2.99
+ $X2=6.94 $Y2=2.99
r90 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.775 $Y=2.99
+ $X2=6.085 $Y2=2.99
r91 38 60 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.927 $Y=2.905
+ $X2=5.927 $Y2=2.99
r92 37 58 2.68365 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.927 $Y=2.09
+ $X2=5.927 $Y2=2.005
r93 37 38 29.8172 $w=3.13e-07 $l=8.15e-07 $layer=LI1_cond $X=5.927 $Y=2.09
+ $X2=5.927 $Y2=2.905
r94 36 56 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.1 $Y=2.005
+ $X2=5.005 $Y2=2.005
r95 35 58 4.95685 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=5.77 $Y=2.005
+ $X2=5.927 $Y2=2.005
r96 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.77 $Y=2.005
+ $X2=5.1 $Y2=2.005
r97 31 56 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=2.09
+ $X2=5.005 $Y2=2.005
r98 31 33 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=5.005 $Y=2.09
+ $X2=5.005 $Y2=2.91
r99 30 54 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=4.24 $Y=2.005
+ $X2=4.052 $Y2=2.005
r100 29 56 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.91 $Y=2.005
+ $X2=5.005 $Y2=2.005
r101 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.91 $Y=2.005
+ $X2=4.24 $Y2=2.005
r102 25 54 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.052 $Y=2.09
+ $X2=4.052 $Y2=2.005
r103 25 27 25.2001 $w=3.73e-07 $l=8.2e-07 $layer=LI1_cond $X=4.052 $Y=2.09
+ $X2=4.052 $Y2=2.91
r104 24 52 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.79 $Y=2.005
+ $X2=2.665 $Y2=2.005
r105 23 54 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=3.865 $Y=2.005
+ $X2=4.052 $Y2=2.005
r106 23 24 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=3.865 $Y=2.005
+ $X2=2.79 $Y2=2.005
r107 19 52 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=2.09
+ $X2=2.665 $Y2=2.005
r108 19 21 37.8001 $w=2.48e-07 $l=8.2e-07 $layer=LI1_cond $X=2.665 $Y=2.09
+ $X2=2.665 $Y2=2.91
r109 6 63 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=1.835 $X2=7.875 $Y2=2.91
r110 6 49 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=7.735
+ $Y=1.835 $X2=7.875 $Y2=2.085
r111 5 43 300 $w=1.7e-07 $l=6.43584e-07 $layer=licon1_PDIFF $count=2 $X=6.725
+ $Y=1.835 $X2=6.94 $Y2=2.38
r112 4 60 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.835 $X2=5.925 $Y2=2.91
r113 4 58 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.835 $X2=5.925 $Y2=2.085
r114 3 56 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.835 $X2=5.005 $Y2=2.085
r115 3 33 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.835 $X2=5.005 $Y2=2.91
r116 2 54 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.835 $X2=4.145 $Y2=2.085
r117 2 27 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=4.02
+ $Y=1.835 $X2=4.145 $Y2=2.91
r118 1 52 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=1.835 $X2=2.695 $Y2=2.085
r119 1 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.555
+ $Y=1.835 $X2=2.695 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 53 63 64 70 73 76 79
r113 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r114 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r115 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r116 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r118 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r119 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r120 61 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.62 $Y=0 $X2=7.455
+ $Y2=0
r121 61 63 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.62 $Y=0 $X2=7.92
+ $Y2=0
r122 60 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r123 59 60 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r124 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r125 56 59 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6.96
+ $Y2=0
r126 56 57 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r127 54 76 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.135
+ $Y2=0
r128 54 56 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.6
+ $Y2=0
r129 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=7.455
+ $Y2=0
r130 53 59 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=6.96
+ $Y2=0
r131 52 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r132 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r133 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r134 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.175
+ $Y2=0
r135 49 51 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.64
+ $Y2=0
r136 48 76 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=3.135
+ $Y2=0
r137 48 51 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.64
+ $Y2=0
r138 47 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r139 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r140 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r141 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.225
+ $Y2=0
r142 44 46 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.39 $Y=0 $X2=1.68
+ $Y2=0
r143 43 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.175
+ $Y2=0
r144 43 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.68
+ $Y2=0
r145 42 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r146 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r147 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r148 39 67 4.57341 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.265
+ $Y2=0
r149 39 41 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.72
+ $Y2=0
r150 38 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=1.225
+ $Y2=0
r151 38 41 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=0.72
+ $Y2=0
r152 36 60 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=6.96 $Y2=0
r153 36 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r154 32 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.455 $Y=0.085
+ $X2=7.455 $Y2=0
r155 32 34 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.455 $Y=0.085
+ $X2=7.455 $Y2=0.45
r156 28 76 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=0.085
+ $X2=3.135 $Y2=0
r157 28 30 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=3.135 $Y=0.085
+ $X2=3.135 $Y2=0.4
r158 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0
r159 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0.38
r160 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0
r161 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.225 $Y=0.085
+ $X2=1.225 $Y2=0.36
r162 16 67 3.19276 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.365 $Y=0.085
+ $X2=0.265 $Y2=0
r163 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.365 $Y=0.085
+ $X2=0.365 $Y2=0.38
r164 5 34 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.315
+ $Y=0.325 $X2=7.455 $Y2=0.45
r165 4 30 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.985
+ $Y=0.235 $X2=3.125 $Y2=0.4
r166 3 26 91 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=2 $X=1.945
+ $Y=0.235 $X2=2.175 $Y2=0.38
r167 2 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.235 $X2=1.225 $Y2=0.36
r168 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.24
+ $Y=0.235 $X2=0.365 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%A_511_47# 1 2 9 11 12 14 15 17
r38 15 17 34.3517 $w=2.58e-07 $l=7.75e-07 $layer=LI1_cond $X=3.58 $Y=0.385
+ $X2=4.355 $Y2=0.385
r39 13 15 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.495 $Y=0.515
+ $X2=3.58 $Y2=0.385
r40 13 14 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.495 $Y=0.515
+ $X2=3.495 $Y2=0.735
r41 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.41 $Y=0.82
+ $X2=3.495 $Y2=0.735
r42 11 12 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.41 $Y=0.82
+ $X2=2.86 $Y2=0.82
r43 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.695 $Y=0.735
+ $X2=2.86 $Y2=0.82
r44 7 9 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.695 $Y=0.735
+ $X2=2.695 $Y2=0.36
r45 2 17 182 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=1 $X=4.215
+ $Y=0.235 $X2=4.355 $Y2=0.375
r46 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.555
+ $Y=0.235 $X2=2.695 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%A_760_47# 1 2 3 10 14 16 23
r35 17 21 3.55261 $w=1.9e-07 $l=1.03e-07 $layer=LI1_cond $X=4.895 $Y=0.35
+ $X2=4.792 $Y2=0.35
r36 16 23 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.48 $Y=0.35
+ $X2=5.645 $Y2=0.35
r37 16 17 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=5.48 $Y=0.35
+ $X2=4.895 $Y2=0.35
r38 14 21 3.27668 $w=2.05e-07 $l=9.5e-08 $layer=LI1_cond $X=4.792 $Y=0.445
+ $X2=4.792 $Y2=0.35
r39 14 15 12.9845 $w=2.03e-07 $l=2.4e-07 $layer=LI1_cond $X=4.792 $Y=0.445
+ $X2=4.792 $Y2=0.685
r40 10 15 6.81778 $w=2.1e-07 $l=1.47428e-07 $layer=LI1_cond $X=4.69 $Y=0.79
+ $X2=4.792 $Y2=0.685
r41 10 12 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=4.69 $Y=0.79
+ $X2=3.925 $Y2=0.79
r42 3 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.505
+ $Y=0.235 $X2=5.645 $Y2=0.38
r43 2 21 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.645
+ $Y=0.235 $X2=4.785 $Y2=0.42
r44 1 12 182 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_NDIFF $count=1 $X=3.8
+ $Y=0.235 $X2=3.925 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_4%A_1208_65# 1 2 3 12 14 15 20 21 24
r41 22 24 26.8165 $w=2.58e-07 $l=6.05e-07 $layer=LI1_cond $X=7.92 $Y=1.075
+ $X2=7.92 $Y2=0.47
r42 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.79 $Y=1.16
+ $X2=7.92 $Y2=1.075
r43 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.79 $Y=1.16
+ $X2=7.12 $Y2=1.16
r44 17 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.025 $Y=1.075
+ $X2=7.12 $Y2=1.16
r45 17 19 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=7.025 $Y=1.075
+ $X2=7.025 $Y2=0.47
r46 16 19 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=7.025 $Y=0.425
+ $X2=7.025 $Y2=0.47
r47 14 16 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.93 $Y=0.34
+ $X2=7.025 $Y2=0.425
r48 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.93 $Y=0.34
+ $X2=6.26 $Y2=0.34
r49 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.13 $Y=0.425
+ $X2=6.26 $Y2=0.34
r50 10 12 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=6.13 $Y=0.425
+ $X2=6.13 $Y2=0.67
r51 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.745
+ $Y=0.325 $X2=7.885 $Y2=0.47
r52 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.885
+ $Y=0.325 $X2=7.025 $Y2=0.47
r53 1 12 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.325 $X2=6.165 $Y2=0.67
.ends

