* File: sky130_fd_sc_lp__o21ai_2.pex.spice
* Created: Fri Aug 28 11:04:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21AI_2%A1 3 7 11 15 20 26 27 28 29 34 37
c78 37 0 1.05768e-19 $X=1.955 $Y=1.51
c79 20 0 1.09305e-19 $X=0.29 $Y=1.46
c80 15 0 1.84841e-19 $X=1.975 $Y=0.655
r81 37 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.51
+ $X2=1.955 $Y2=1.675
r82 37 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.51
+ $X2=1.955 $Y2=1.345
r83 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=1.51 $X2=1.955 $Y2=1.51
r84 29 38 5.83335 $w=4.03e-07 $l=2.05e-07 $layer=LI1_cond $X=2.16 $Y=1.547
+ $X2=1.955 $Y2=1.547
r85 28 38 7.82523 $w=4.03e-07 $l=2.75e-07 $layer=LI1_cond $X=1.68 $Y=1.547
+ $X2=1.955 $Y2=1.547
r86 27 28 7.54068 $w=4.03e-07 $l=2.65e-07 $layer=LI1_cond $X=1.415 $Y=1.547
+ $X2=1.68 $Y2=1.547
r87 26 27 8.81108 $w=4.03e-07 $l=1.7e-07 $layer=LI1_cond $X=1.245 $Y=1.605
+ $X2=1.415 $Y2=1.605
r88 21 34 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.29 $Y=1.46 $X2=0.49
+ $Y2=1.46
r89 20 23 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.29 $Y=1.46
+ $X2=0.29 $Y2=1.78
r90 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.46 $X2=0.29 $Y2=1.46
r91 18 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=1.78
+ $X2=0.29 $Y2=1.78
r92 18 26 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.455 $Y=1.78
+ $X2=1.245 $Y2=1.78
r93 15 39 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.975 $Y=0.655
+ $X2=1.975 $Y2=1.345
r94 11 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.935 $Y=2.465
+ $X2=1.935 $Y2=1.675
r95 5 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.625
+ $X2=0.49 $Y2=1.46
r96 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.49 $Y=1.625 $X2=0.49
+ $Y2=2.465
r97 1 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.295
+ $X2=0.49 $Y2=1.46
r98 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.49 $Y=1.295 $X2=0.49
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_2%A2 1 3 6 8 10 13 15 21 22
c53 22 0 1.09305e-19 $X=1.35 $Y=1.35
r54 20 22 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.94 $Y=1.35
+ $X2=1.35 $Y2=1.35
r55 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.35 $X2=0.94 $Y2=1.35
r56 17 20 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.92 $Y=1.35 $X2=0.94
+ $Y2=1.35
r57 15 21 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.72 $Y=1.35
+ $X2=0.94 $Y2=1.35
r58 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.515
+ $X2=1.35 $Y2=1.35
r59 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.35 $Y=1.515
+ $X2=1.35 $Y2=2.465
r60 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.185
+ $X2=1.35 $Y2=1.35
r61 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.35 $Y=1.185
+ $X2=1.35 $Y2=0.655
r62 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.515
+ $X2=0.92 $Y2=1.35
r63 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.92 $Y=1.515 $X2=0.92
+ $Y2=2.465
r64 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.185
+ $X2=0.92 $Y2=1.35
r65 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.92 $Y=1.185 $X2=0.92
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_2%B1 3 7 9 11 14 16 17 21
c44 9 0 6.40318e-20 $X=2.835 $Y=1.185
r45 21 23 35.6195 $w=3.18e-07 $l=2.35e-07 $layer=POLY_cond $X=2.835 $Y=1.35
+ $X2=3.07 $Y2=1.35
r46 16 17 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.085 $Y=1.295
+ $X2=3.085 $Y2=1.665
r47 16 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.35 $X2=3.07 $Y2=1.35
r48 12 21 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.515
+ $X2=2.835 $Y2=1.35
r49 12 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.835 $Y=1.515
+ $X2=2.835 $Y2=2.465
r50 9 21 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.185
+ $X2=2.835 $Y2=1.35
r51 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.835 $Y=1.185
+ $X2=2.835 $Y2=0.655
r52 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.405 $Y=1.515
+ $X2=2.405 $Y2=2.465
r53 1 21 65.1761 $w=3.18e-07 $l=4.3e-07 $layer=POLY_cond $X=2.405 $Y=1.35
+ $X2=2.835 $Y2=1.35
r54 1 5 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.35
+ $X2=2.405 $Y2=1.515
r55 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.405 $Y=1.21
+ $X2=2.405 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_2%VPWR 1 2 3 10 12 18 20 22 26 28 36 45 49
r46 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 40 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 40 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 37 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.165 $Y2=3.33
r53 37 39 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 36 48 4.49223 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=3.132 $Y2=3.33
r55 36 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 32 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r58 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 29 42 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r60 29 31 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 28 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=2.165
+ $Y2=3.33
r62 28 34 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r63 26 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r64 26 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 26 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 22 25 32.1569 $w=3.08e-07 $l=8.65e-07 $layer=LI1_cond $X=3.06 $Y=2.085
+ $X2=3.06 $Y2=2.95
r67 20 48 3.10696 $w=3.1e-07 $l=1.15521e-07 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.132 $Y2=3.33
r68 20 25 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=2.95
r69 16 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=3.33
r70 16 18 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=2.165 $Y=3.245
+ $X2=2.165 $Y2=2.49
r71 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.275 $Y=2.12
+ $X2=0.275 $Y2=2.95
r72 10 42 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r73 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.95
r74 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.91
+ $Y=1.835 $X2=3.05 $Y2=2.95
r75 3 22 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=2.91
+ $Y=1.835 $X2=3.05 $Y2=2.085
r76 2 18 300 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_PDIFF $count=2 $X=2.01
+ $Y=1.835 $X2=2.165 $Y2=2.49
r77 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.95
r78 1 12 400 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_2%A_113_367# 1 2 7 9 11 15
r16 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.64 $Y=2.905
+ $X2=1.64 $Y2=2.49
r17 12 18 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.83 $Y=2.99 $X2=0.72
+ $Y2=2.99
r18 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.475 $Y=2.99
+ $X2=1.64 $Y2=2.905
r19 11 12 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.475 $Y=2.99
+ $X2=0.83 $Y2=2.99
r20 7 18 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=2.905 $X2=0.72
+ $Y2=2.99
r21 7 9 36.9306 $w=2.18e-07 $l=7.05e-07 $layer=LI1_cond $X=0.72 $Y=2.905
+ $X2=0.72 $Y2=2.2
r22 2 15 300 $w=1.7e-07 $l=7.54884e-07 $layer=licon1_PDIFF $count=2 $X=1.425
+ $Y=1.835 $X2=1.64 $Y2=2.49
r23 1 18 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.91
r24 1 9 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_2%Y 1 2 3 14 18 22 23 24 25 31 32 41
c38 18 0 1.05768e-19 $X=2.62 $Y=0.76
r39 32 41 2.30489 $w=2.83e-07 $l=5.7e-08 $layer=LI1_cond $X=1.737 $Y=2.062
+ $X2=1.68 $Y2=2.062
r40 25 31 0.468231 $w=2.85e-07 $l=1.17e-07 $layer=LI1_cond $X=2.617 $Y=2.062
+ $X2=2.5 $Y2=2.062
r41 24 31 13.7484 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=2.16 $Y=2.062
+ $X2=2.5 $Y2=2.062
r42 23 41 0.566112 $w=2.83e-07 $l=1.4e-08 $layer=LI1_cond $X=1.666 $Y=2.062
+ $X2=1.68 $Y2=2.062
r43 23 24 16.5386 $w=2.83e-07 $l=4.09e-07 $layer=LI1_cond $X=1.751 $Y=2.062
+ $X2=2.16 $Y2=2.062
r44 23 32 0.566112 $w=2.83e-07 $l=1.4e-08 $layer=LI1_cond $X=1.751 $Y=2.062
+ $X2=1.737 $Y2=2.062
r45 20 23 14.6157 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.3 $Y=2.12
+ $X2=1.595 $Y2=2.12
r46 20 22 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.3 $Y=2.12 $X2=1.15
+ $Y2=2.12
r47 16 25 6.31478 $w=2.22e-07 $l=1.48358e-07 $layer=LI1_cond $X=2.63 $Y=1.92
+ $X2=2.617 $Y2=2.062
r48 16 18 61.2641 $w=2.08e-07 $l=1.16e-06 $layer=LI1_cond $X=2.63 $Y=1.92
+ $X2=2.63 $Y2=0.76
r49 12 25 6.31478 $w=2.22e-07 $l=1.43e-07 $layer=LI1_cond $X=2.617 $Y=2.205
+ $X2=2.617 $Y2=2.062
r50 12 14 11.5244 $w=2.33e-07 $l=2.35e-07 $layer=LI1_cond $X=2.617 $Y=2.205
+ $X2=2.617 $Y2=2.44
r51 3 25 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=1.98
r52 3 14 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2.44
r53 2 22 300 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=2 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.2
r54 1 18 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.62 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_2%A_30_47# 1 2 3 4 13 15 17 21 23 25 26 27 34
+ 39
c60 39 0 6.40318e-20 $X=3.05 $Y=0.42
c61 21 0 1.84841e-19 $X=1.135 $Y=0.42
r62 34 35 7.83936 $w=2.49e-07 $l=1.6e-07 $layer=LI1_cond $X=1.202 $Y=0.93
+ $X2=1.202 $Y2=1.09
r63 28 37 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.355 $Y=0.34
+ $X2=2.195 $Y2=0.34
r64 27 39 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.905 $Y=0.34
+ $X2=3.06 $Y2=0.34
r65 27 28 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.905 $Y=0.34
+ $X2=2.355 $Y2=0.34
r66 25 37 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0.425
+ $X2=2.195 $Y2=0.34
r67 25 26 20.888 $w=3.18e-07 $l=5.8e-07 $layer=LI1_cond $X=2.195 $Y=0.425
+ $X2=2.195 $Y2=1.005
r68 24 35 2.97181 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=1.365 $Y=1.09
+ $X2=1.202 $Y2=1.09
r69 23 26 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=2.035 $Y=1.09
+ $X2=2.195 $Y2=1.005
r70 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.035 $Y=1.09
+ $X2=1.365 $Y2=1.09
r71 19 34 3.88855 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.202 $Y=0.845
+ $X2=1.202 $Y2=0.93
r72 19 21 15.0704 $w=3.23e-07 $l=4.25e-07 $layer=LI1_cond $X=1.202 $Y=0.845
+ $X2=1.202 $Y2=0.42
r73 18 32 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.37 $Y=0.93 $X2=0.24
+ $Y2=0.93
r74 17 34 2.97181 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=1.04 $Y=0.93
+ $X2=1.202 $Y2=0.93
r75 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.04 $Y=0.93
+ $X2=0.37 $Y2=0.93
r76 13 32 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=0.845
+ $X2=0.24 $Y2=0.93
r77 13 15 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=0.24 $Y=0.845
+ $X2=0.24 $Y2=0.42
r78 4 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.91
+ $Y=0.235 $X2=3.05 $Y2=0.42
r79 3 37 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.05
+ $Y=0.235 $X2=2.19 $Y2=0.42
r80 2 34 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.235 $X2=1.135 $Y2=0.93
r81 2 21 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.235 $X2=1.135 $Y2=0.42
r82 1 32 182 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.93
r83 1 15 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r46 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r49 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r50 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r51 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.7
+ $Y2=0
r52 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r53 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r54 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r55 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=0 $X2=0.705
+ $Y2=0
r56 23 25 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.87 $Y=0 $X2=1.2
+ $Y2=0
r57 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.7
+ $Y2=0
r58 22 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.2
+ $Y2=0
r59 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r60 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r61 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=0.705
+ $Y2=0
r62 17 19 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=0.24
+ $Y2=0
r63 15 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r64 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r65 15 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r66 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r67 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.7 $Y=0.085
+ $X2=1.7 $Y2=0.38
r68 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r69 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.55
r70 2 13 91 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=2 $X=1.425
+ $Y=0.235 $X2=1.7 $Y2=0.38
r71 1 9 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.705 $Y2=0.55
.ends

