* File: sky130_fd_sc_lp__a32oi_1.pxi.spice
* Created: Fri Aug 28 10:01:37 2020
* 
x_PM_SKY130_FD_SC_LP__A32OI_1%B2 N_B2_c_50_n N_B2_M1006_g N_B2_M1000_g B2 B2
+ N_B2_c_53_n PM_SKY130_FD_SC_LP__A32OI_1%B2
x_PM_SKY130_FD_SC_LP__A32OI_1%B1 N_B1_M1004_g N_B1_M1002_g B1 B1 N_B1_c_78_n
+ N_B1_c_79_n PM_SKY130_FD_SC_LP__A32OI_1%B1
x_PM_SKY130_FD_SC_LP__A32OI_1%A1 N_A1_M1001_g N_A1_M1005_g A1 A1 A1 A1
+ N_A1_c_112_n N_A1_c_113_n PM_SKY130_FD_SC_LP__A32OI_1%A1
x_PM_SKY130_FD_SC_LP__A32OI_1%A2 N_A2_c_149_n N_A2_M1008_g N_A2_M1007_g A2 A2 A2
+ A2 N_A2_c_152_n PM_SKY130_FD_SC_LP__A32OI_1%A2
x_PM_SKY130_FD_SC_LP__A32OI_1%A3 N_A3_M1009_g N_A3_M1003_g A3 A3 N_A3_c_190_n
+ N_A3_c_191_n PM_SKY130_FD_SC_LP__A32OI_1%A3
x_PM_SKY130_FD_SC_LP__A32OI_1%A_58_367# N_A_58_367#_M1000_s N_A_58_367#_M1002_d
+ N_A_58_367#_M1007_d N_A_58_367#_c_214_n N_A_58_367#_c_215_n
+ N_A_58_367#_c_218_n N_A_58_367#_c_227_p N_A_58_367#_c_220_n
+ N_A_58_367#_c_223_n N_A_58_367#_c_232_p PM_SKY130_FD_SC_LP__A32OI_1%A_58_367#
x_PM_SKY130_FD_SC_LP__A32OI_1%Y N_Y_M1004_d N_Y_M1000_d N_Y_c_240_n N_Y_c_252_n
+ N_Y_c_247_n N_Y_c_241_n N_Y_c_248_n Y Y Y PM_SKY130_FD_SC_LP__A32OI_1%Y
x_PM_SKY130_FD_SC_LP__A32OI_1%VPWR N_VPWR_M1005_d N_VPWR_M1003_d N_VPWR_c_287_n
+ N_VPWR_c_288_n VPWR N_VPWR_c_289_n N_VPWR_c_290_n N_VPWR_c_291_n
+ N_VPWR_c_286_n PM_SKY130_FD_SC_LP__A32OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A32OI_1%VGND N_VGND_M1006_s N_VGND_M1009_d N_VGND_c_324_n
+ N_VGND_c_325_n N_VGND_c_326_n N_VGND_c_327_n N_VGND_c_328_n N_VGND_c_329_n
+ VGND N_VGND_c_330_n PM_SKY130_FD_SC_LP__A32OI_1%VGND
cc_1 VNB N_B2_c_50_n 0.0182255f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_2 VNB N_B2_M1000_g 0.00146484f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.465
cc_3 VNB B2 0.0235771f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B2_c_53_n 0.0475398f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.46
cc_5 VNB N_B1_M1002_g 0.00146768f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.465
cc_6 VNB B1 0.00541326f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_B1_c_78_n 0.0317804f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.46
cc_8 VNB N_B1_c_79_n 0.0177051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_M1005_g 0.00172813f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.465
cc_10 VNB A1 0.00289143f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A1_c_112_n 0.0306676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_c_113_n 0.0189785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_149_n 0.0186615f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_14 VNB N_A2_M1007_g 0.00166373f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.465
cc_15 VNB A2 0.00380017f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_A2_c_152_n 0.036647f $X=-0.19 $Y=-0.245 $X2=0.332 $Y2=1.46
cc_17 VNB N_A3_M1003_g 0.00167964f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.465
cc_18 VNB A3 0.0381205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A3_c_190_n 0.0346344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A3_c_191_n 0.0212673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_240_n 0.0028212f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_Y_c_241_n 0.00294489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_286_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_324_n 0.0151766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_325_n 0.0375479f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_VGND_c_326_n 0.0358924f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.46
cc_27 VNB N_VGND_c_327_n 0.0115308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_328_n 0.0634279f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.46
cc_29 VNB N_VGND_c_329_n 0.00596836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_330_n 0.233291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_B2_M1000_g 0.0246363f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_32 VPB B2 0.0102988f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_33 VPB N_B1_M1002_g 0.0206822f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_34 VPB B1 0.00273154f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_35 VPB N_A1_M1005_g 0.0233987f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_36 VPB A1 0.00257255f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_37 VPB N_A2_M1007_g 0.0226713f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_38 VPB A2 0.00293638f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_39 VPB N_A3_M1003_g 0.0250078f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_40 VPB A3 0.0162725f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_58_367#_c_214_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_58_367#_c_215_n 0.0373161f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.46
cc_43 VPB N_Y_c_240_n 0.0013607f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_44 VPB N_VPWR_c_287_n 0.0144866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_288_n 0.0481737f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_46 VPB N_VPWR_c_289_n 0.04078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_290_n 0.0129657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_291_n 0.0123114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_286_n 0.0558779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 N_B2_M1000_g N_B1_M1002_g 0.0363863f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_51 N_B2_c_50_n B1 4.641e-19 $X=0.63 $Y=1.295 $X2=0 $Y2=0
cc_52 N_B2_c_53_n N_B1_c_78_n 0.039024f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_53 N_B2_c_50_n N_B1_c_79_n 0.039024f $X=0.63 $Y=1.295 $X2=0 $Y2=0
cc_54 B2 N_A_58_367#_c_215_n 0.0228788f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_55 N_B2_c_53_n N_A_58_367#_c_215_n 0.0014231f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_56 N_B2_M1000_g N_A_58_367#_c_218_n 0.0114565f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_57 N_B2_c_50_n N_Y_c_240_n 0.00921929f $X=0.63 $Y=1.295 $X2=0 $Y2=0
cc_58 N_B2_M1000_g N_Y_c_240_n 0.00970296f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_59 B2 N_Y_c_240_n 0.0395886f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_60 N_B2_c_53_n N_Y_c_240_n 0.00721317f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_61 N_B2_c_50_n N_Y_c_247_n 0.00435494f $X=0.63 $Y=1.295 $X2=0 $Y2=0
cc_62 N_B2_M1000_g N_Y_c_248_n 0.0113015f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_63 N_B2_M1000_g N_VPWR_c_289_n 0.00357877f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_64 N_B2_M1000_g N_VPWR_c_286_n 0.00642834f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_65 N_B2_c_50_n N_VGND_c_325_n 0.0049025f $X=0.63 $Y=1.295 $X2=0 $Y2=0
cc_66 B2 N_VGND_c_325_n 0.0228787f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B2_c_53_n N_VGND_c_325_n 0.0015566f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_68 N_B2_c_50_n N_VGND_c_328_n 0.00482246f $X=0.63 $Y=1.295 $X2=0 $Y2=0
cc_69 N_B2_c_50_n N_VGND_c_330_n 0.008955f $X=0.63 $Y=1.295 $X2=0 $Y2=0
cc_70 N_B1_M1002_g N_A1_M1005_g 0.0290799f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_71 B1 A1 0.0381267f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_72 N_B1_c_78_n A1 3.0655e-19 $X=1.105 $Y=1.46 $X2=0 $Y2=0
cc_73 N_B1_c_79_n A1 8.35611e-19 $X=1.1 $Y=1.295 $X2=0 $Y2=0
cc_74 N_B1_c_78_n N_A1_c_112_n 0.0204825f $X=1.105 $Y=1.46 $X2=0 $Y2=0
cc_75 B1 N_A1_c_113_n 0.00388205f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B1_c_79_n N_A1_c_113_n 0.0177752f $X=1.1 $Y=1.295 $X2=0 $Y2=0
cc_77 N_B1_M1002_g N_A_58_367#_c_218_n 0.0114565f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_78 N_B1_M1002_g N_Y_c_240_n 0.00410365f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_79 B1 N_Y_c_240_n 0.0406434f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B1_c_79_n N_Y_c_240_n 0.00646802f $X=1.1 $Y=1.295 $X2=0 $Y2=0
cc_81 B1 N_Y_c_252_n 0.0275498f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_B1_c_78_n N_Y_c_252_n 9.83929e-19 $X=1.105 $Y=1.46 $X2=0 $Y2=0
cc_83 N_B1_c_79_n N_Y_c_252_n 0.0124879f $X=1.1 $Y=1.295 $X2=0 $Y2=0
cc_84 N_B1_c_79_n N_Y_c_241_n 3.07349e-19 $X=1.1 $Y=1.295 $X2=0 $Y2=0
cc_85 N_B1_M1002_g N_Y_c_248_n 0.0120927f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_86 N_B1_M1002_g Y 0.0126458f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_87 B1 Y 0.0253649f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B1_c_78_n Y 6.02193e-19 $X=1.105 $Y=1.46 $X2=0 $Y2=0
cc_89 N_B1_M1002_g N_VPWR_c_289_n 0.00357877f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_90 N_B1_M1002_g N_VPWR_c_291_n 0.0010514f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B1_M1002_g N_VPWR_c_286_n 0.00555273f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_92 N_B1_c_79_n N_VGND_c_328_n 0.00482246f $X=1.1 $Y=1.295 $X2=0 $Y2=0
cc_93 N_B1_c_79_n N_VGND_c_330_n 0.00518737f $X=1.1 $Y=1.295 $X2=0 $Y2=0
cc_94 A1 N_A2_c_149_n 0.00435278f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_95 N_A1_c_113_n N_A2_c_149_n 0.0320864f $X=1.645 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_96 N_A1_M1005_g N_A2_M1007_g 0.0205255f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_97 A1 N_A2_M1007_g 3.02778e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_98 N_A1_M1005_g A2 3.40421e-19 $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_99 A1 A2 0.0783179f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_100 N_A1_c_112_n A2 0.00103129f $X=1.645 $Y=1.46 $X2=0 $Y2=0
cc_101 N_A1_c_113_n A2 8.03333e-19 $X=1.645 $Y=1.295 $X2=0 $Y2=0
cc_102 N_A1_c_112_n N_A2_c_152_n 0.0214281f $X=1.645 $Y=1.46 $X2=0 $Y2=0
cc_103 N_A1_M1005_g N_A_58_367#_c_220_n 0.0135479f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_104 A1 N_Y_c_252_n 0.0147293f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_105 N_A1_c_113_n N_Y_c_252_n 0.00160472f $X=1.645 $Y=1.295 $X2=0 $Y2=0
cc_106 A1 N_Y_c_241_n 0.037115f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_107 N_A1_c_113_n N_Y_c_241_n 0.00524161f $X=1.645 $Y=1.295 $X2=0 $Y2=0
cc_108 N_A1_M1005_g N_Y_c_248_n 7.33113e-19 $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A1_M1005_g Y 0.0160746f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_110 A1 Y 0.020327f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_111 N_A1_c_112_n Y 8.36724e-19 $X=1.645 $Y=1.46 $X2=0 $Y2=0
cc_112 N_A1_M1005_g N_VPWR_c_289_n 0.00487821f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A1_M1005_g N_VPWR_c_291_n 0.0139259f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A1_M1005_g N_VPWR_c_286_n 0.00842155f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_115 A1 N_VGND_c_328_n 0.00976442f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_116 N_A1_c_113_n N_VGND_c_328_n 0.00402307f $X=1.645 $Y=1.295 $X2=0 $Y2=0
cc_117 A1 N_VGND_c_330_n 0.00962478f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_118 N_A1_c_113_n N_VGND_c_330_n 0.00715227f $X=1.645 $Y=1.295 $X2=0 $Y2=0
cc_119 A1 A_326_69# 0.00975772f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_120 N_A2_M1007_g N_A3_M1003_g 0.0202745f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A2_c_149_n A3 2.47212e-19 $X=2.095 $Y=1.295 $X2=0 $Y2=0
cc_122 A2 A3 0.0458168f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_123 N_A2_c_152_n A3 0.00314725f $X=2.325 $Y=1.46 $X2=0 $Y2=0
cc_124 A2 N_A3_c_190_n 3.17196e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_125 N_A2_c_152_n N_A3_c_190_n 0.0206996f $X=2.325 $Y=1.46 $X2=0 $Y2=0
cc_126 N_A2_c_149_n N_A3_c_191_n 0.0246644f $X=2.095 $Y=1.295 $X2=0 $Y2=0
cc_127 A2 N_A3_c_191_n 0.00998065f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A2_M1007_g N_A_58_367#_c_220_n 0.0163409f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_129 A2 N_A_58_367#_c_220_n 0.00276744f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_130 N_A2_M1007_g Y 0.00574272f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_131 A2 Y 0.0187578f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_132 N_A2_c_152_n Y 0.00108735f $X=2.325 $Y=1.46 $X2=0 $Y2=0
cc_133 N_A2_M1007_g N_VPWR_c_288_n 7.81248e-19 $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A2_M1007_g N_VPWR_c_290_n 0.00487821f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A2_M1007_g N_VPWR_c_291_n 0.0126214f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A2_M1007_g N_VPWR_c_286_n 0.00827265f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A2_c_149_n N_VGND_c_326_n 0.00132803f $X=2.095 $Y=1.295 $X2=0 $Y2=0
cc_138 A2 N_VGND_c_326_n 0.0278396f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_139 N_A2_c_149_n N_VGND_c_328_n 0.00308465f $X=2.095 $Y=1.295 $X2=0 $Y2=0
cc_140 A2 N_VGND_c_328_n 0.0121702f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_141 N_A2_c_149_n N_VGND_c_330_n 0.00421028f $X=2.095 $Y=1.295 $X2=0 $Y2=0
cc_142 A2 N_VGND_c_330_n 0.0117847f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_143 A2 A_434_69# 0.0118277f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_144 A3 N_A_58_367#_c_223_n 0.00975719f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_145 N_A3_M1003_g N_VPWR_c_288_n 0.0202307f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_146 A3 N_VPWR_c_288_n 0.0262295f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A3_c_190_n N_VPWR_c_288_n 5.0317e-19 $X=2.775 $Y=1.46 $X2=0 $Y2=0
cc_148 N_A3_M1003_g N_VPWR_c_290_n 0.00486043f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A3_M1003_g N_VPWR_c_291_n 5.90548e-19 $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A3_M1003_g N_VPWR_c_286_n 0.0082726f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_151 A3 N_VGND_c_326_n 0.0267908f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A3_c_190_n N_VGND_c_326_n 9.95955e-19 $X=2.775 $Y=1.46 $X2=0 $Y2=0
cc_153 N_A3_c_191_n N_VGND_c_326_n 0.0184425f $X=2.775 $Y=1.295 $X2=0 $Y2=0
cc_154 N_A3_c_191_n N_VGND_c_328_n 0.00400407f $X=2.775 $Y=1.295 $X2=0 $Y2=0
cc_155 N_A3_c_191_n N_VGND_c_330_n 0.0078287f $X=2.775 $Y=1.295 $X2=0 $Y2=0
cc_156 N_A_58_367#_c_218_n N_Y_M1000_d 0.00332344f $X=1.18 $Y=2.99 $X2=0 $Y2=0
cc_157 N_A_58_367#_c_218_n N_Y_c_248_n 0.0159805f $X=1.18 $Y=2.99 $X2=0 $Y2=0
cc_158 N_A_58_367#_M1002_d Y 0.00645472f $X=1.135 $Y=1.835 $X2=0 $Y2=0
cc_159 N_A_58_367#_c_227_p Y 0.0190017f $X=1.307 $Y=2.46 $X2=0 $Y2=0
cc_160 N_A_58_367#_c_220_n Y 0.0478108f $X=2.425 $Y=2.375 $X2=0 $Y2=0
cc_161 N_A_58_367#_c_220_n N_VPWR_M1005_d 0.0129627f $X=2.425 $Y=2.375 $X2=-0.19
+ $Y2=1.655
cc_162 N_A_58_367#_c_214_n N_VPWR_c_289_n 0.0179183f $X=0.38 $Y=2.905 $X2=0
+ $Y2=0
cc_163 N_A_58_367#_c_218_n N_VPWR_c_289_n 0.0532109f $X=1.18 $Y=2.99 $X2=0 $Y2=0
cc_164 N_A_58_367#_c_232_p N_VPWR_c_290_n 0.0124525f $X=2.54 $Y=2.495 $X2=0
+ $Y2=0
cc_165 N_A_58_367#_c_220_n N_VPWR_c_291_n 0.0447396f $X=2.425 $Y=2.375 $X2=0
+ $Y2=0
cc_166 N_A_58_367#_M1000_s N_VPWR_c_286_n 0.00215161f $X=0.29 $Y=1.835 $X2=0
+ $Y2=0
cc_167 N_A_58_367#_M1002_d N_VPWR_c_286_n 0.00428898f $X=1.135 $Y=1.835 $X2=0
+ $Y2=0
cc_168 N_A_58_367#_M1007_d N_VPWR_c_286_n 0.00536646f $X=2.4 $Y=1.835 $X2=0
+ $Y2=0
cc_169 N_A_58_367#_c_214_n N_VPWR_c_286_n 0.0101029f $X=0.38 $Y=2.905 $X2=0
+ $Y2=0
cc_170 N_A_58_367#_c_218_n N_VPWR_c_286_n 0.0335898f $X=1.18 $Y=2.99 $X2=0 $Y2=0
cc_171 N_A_58_367#_c_232_p N_VPWR_c_286_n 0.00730901f $X=2.54 $Y=2.495 $X2=0
+ $Y2=0
cc_172 Y N_VPWR_M1005_d 0.0179733f $X=2.075 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_173 N_Y_M1000_d N_VPWR_c_286_n 0.00225186f $X=0.705 $Y=1.835 $X2=0 $Y2=0
cc_174 N_Y_c_241_n N_VGND_c_325_n 6.37773e-19 $X=1.265 $Y=0.49 $X2=0 $Y2=0
cc_175 N_Y_c_241_n N_VGND_c_328_n 0.0143328f $X=1.265 $Y=0.49 $X2=0 $Y2=0
cc_176 N_Y_c_252_n N_VGND_c_330_n 0.00740192f $X=1.1 $Y=0.95 $X2=0 $Y2=0
cc_177 N_Y_c_247_n N_VGND_c_330_n 0.00639544f $X=0.85 $Y=0.95 $X2=0 $Y2=0
cc_178 N_Y_c_241_n N_VGND_c_330_n 0.0108117f $X=1.265 $Y=0.49 $X2=0 $Y2=0
cc_179 N_Y_c_240_n A_141_69# 0.00159394f $X=0.765 $Y=1.92 $X2=-0.19 $Y2=-0.245
cc_180 N_Y_c_252_n A_141_69# 0.00129817f $X=1.1 $Y=0.95 $X2=-0.19 $Y2=-0.245
cc_181 N_Y_c_247_n A_141_69# 0.00212536f $X=0.85 $Y=0.95 $X2=-0.19 $Y2=-0.245
