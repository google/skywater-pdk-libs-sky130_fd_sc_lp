* File: sky130_fd_sc_lp__dfrtp_4.pxi.spice
* Created: Wed Sep  2 09:43:54 2020
* 
x_PM_SKY130_FD_SC_LP__DFRTP_4%CLK N_CLK_M1020_g N_CLK_M1036_g N_CLK_c_264_n
+ N_CLK_c_269_n CLK CLK CLK N_CLK_c_266_n PM_SKY130_FD_SC_LP__DFRTP_4%CLK
x_PM_SKY130_FD_SC_LP__DFRTP_4%A_27_90# N_A_27_90#_M1020_s N_A_27_90#_M1036_s
+ N_A_27_90#_M1013_g N_A_27_90#_M1021_g N_A_27_90#_M1008_g N_A_27_90#_M1001_g
+ N_A_27_90#_M1014_g N_A_27_90#_M1002_g N_A_27_90#_c_303_n N_A_27_90#_c_304_n
+ N_A_27_90#_c_305_n N_A_27_90#_c_337_n N_A_27_90#_c_306_n N_A_27_90#_c_307_n
+ N_A_27_90#_c_338_n N_A_27_90#_c_359_n N_A_27_90#_c_308_n N_A_27_90#_c_309_n
+ N_A_27_90#_c_310_n N_A_27_90#_c_311_n N_A_27_90#_c_312_n N_A_27_90#_c_313_n
+ N_A_27_90#_c_314_n N_A_27_90#_c_315_n N_A_27_90#_c_316_n N_A_27_90#_c_317_n
+ N_A_27_90#_c_318_n N_A_27_90#_c_319_n N_A_27_90#_c_320_n N_A_27_90#_c_321_n
+ N_A_27_90#_c_341_n N_A_27_90#_c_322_n N_A_27_90#_c_323_n N_A_27_90#_c_324_n
+ N_A_27_90#_c_325_n N_A_27_90#_c_326_n N_A_27_90#_c_327_n N_A_27_90#_c_328_n
+ N_A_27_90#_c_329_n N_A_27_90#_c_386_p N_A_27_90#_c_330_n N_A_27_90#_c_331_n
+ N_A_27_90#_c_332_n N_A_27_90#_c_333_n PM_SKY130_FD_SC_LP__DFRTP_4%A_27_90#
x_PM_SKY130_FD_SC_LP__DFRTP_4%D N_D_M1023_g N_D_M1018_g N_D_c_595_n N_D_c_600_n
+ N_D_c_601_n N_D_c_596_n D D PM_SKY130_FD_SC_LP__DFRTP_4%D
x_PM_SKY130_FD_SC_LP__DFRTP_4%A_216_462# N_A_216_462#_M1021_d
+ N_A_216_462#_M1013_d N_A_216_462#_M1009_g N_A_216_462#_M1031_g
+ N_A_216_462#_M1012_g N_A_216_462#_c_649_n N_A_216_462#_c_650_n
+ N_A_216_462#_c_651_n N_A_216_462#_M1028_g N_A_216_462#_c_658_n
+ N_A_216_462#_c_652_n N_A_216_462#_c_660_n N_A_216_462#_c_661_n
+ N_A_216_462#_c_662_n N_A_216_462#_c_663_n N_A_216_462#_c_664_n
+ N_A_216_462#_c_665_n N_A_216_462#_c_780_p N_A_216_462#_c_666_n
+ N_A_216_462#_c_653_n N_A_216_462#_c_654_n N_A_216_462#_c_669_n
+ N_A_216_462#_c_670_n PM_SKY130_FD_SC_LP__DFRTP_4%A_216_462#
x_PM_SKY130_FD_SC_LP__DFRTP_4%A_731_405# N_A_731_405#_M1025_d
+ N_A_731_405#_M1027_d N_A_731_405#_M1000_g N_A_731_405#_c_877_n
+ N_A_731_405#_c_878_n N_A_731_405#_M1033_g N_A_731_405#_c_879_n
+ N_A_731_405#_c_869_n N_A_731_405#_c_870_n N_A_731_405#_c_871_n
+ N_A_731_405#_c_872_n N_A_731_405#_c_881_n N_A_731_405#_c_915_n
+ N_A_731_405#_c_873_n N_A_731_405#_c_874_n N_A_731_405#_c_875_n
+ N_A_731_405#_c_882_n PM_SKY130_FD_SC_LP__DFRTP_4%A_731_405#
x_PM_SKY130_FD_SC_LP__DFRTP_4%RESET_B N_RESET_B_M1034_g N_RESET_B_c_979_n
+ N_RESET_B_c_980_n N_RESET_B_M1022_g N_RESET_B_c_982_n N_RESET_B_M1007_g
+ N_RESET_B_c_995_n N_RESET_B_c_996_n N_RESET_B_M1010_g N_RESET_B_M1024_g
+ N_RESET_B_M1003_g N_RESET_B_c_985_n N_RESET_B_c_986_n N_RESET_B_c_1000_n
+ N_RESET_B_c_1001_n N_RESET_B_c_1002_n N_RESET_B_c_987_n N_RESET_B_c_988_n
+ N_RESET_B_c_989_n N_RESET_B_c_1004_n N_RESET_B_c_1005_n N_RESET_B_c_1027_n
+ RESET_B RESET_B N_RESET_B_c_990_n N_RESET_B_c_991_n RESET_B
+ PM_SKY130_FD_SC_LP__DFRTP_4%RESET_B
x_PM_SKY130_FD_SC_LP__DFRTP_4%A_595_535# N_A_595_535#_M1008_d
+ N_A_595_535#_M1009_d N_A_595_535#_M1007_d N_A_595_535#_c_1187_n
+ N_A_595_535#_c_1188_n N_A_595_535#_M1025_g N_A_595_535#_M1027_g
+ N_A_595_535#_c_1209_n N_A_595_535#_c_1195_n N_A_595_535#_c_1196_n
+ N_A_595_535#_c_1197_n N_A_595_535#_c_1189_n N_A_595_535#_c_1198_n
+ N_A_595_535#_c_1199_n N_A_595_535#_c_1200_n N_A_595_535#_c_1201_n
+ N_A_595_535#_c_1202_n N_A_595_535#_c_1190_n N_A_595_535#_c_1191_n
+ N_A_595_535#_c_1203_n N_A_595_535#_c_1204_n N_A_595_535#_c_1192_n
+ PM_SKY130_FD_SC_LP__DFRTP_4%A_595_535#
x_PM_SKY130_FD_SC_LP__DFRTP_4%A_1475_426# N_A_1475_426#_M1032_d
+ N_A_1475_426#_M1024_d N_A_1475_426#_M1016_g N_A_1475_426#_M1019_g
+ N_A_1475_426#_c_1339_n N_A_1475_426#_c_1340_n N_A_1475_426#_c_1341_n
+ N_A_1475_426#_c_1369_n N_A_1475_426#_c_1342_n N_A_1475_426#_c_1335_n
+ N_A_1475_426#_c_1336_n N_A_1475_426#_c_1344_n N_A_1475_426#_c_1345_n
+ PM_SKY130_FD_SC_LP__DFRTP_4%A_1475_426#
x_PM_SKY130_FD_SC_LP__DFRTP_4%A_1255_449# N_A_1255_449#_M1012_d
+ N_A_1255_449#_M1014_d N_A_1255_449#_c_1422_n N_A_1255_449#_M1032_g
+ N_A_1255_449#_M1030_g N_A_1255_449#_c_1423_n N_A_1255_449#_c_1424_n
+ N_A_1255_449#_M1035_g N_A_1255_449#_M1011_g N_A_1255_449#_c_1426_n
+ N_A_1255_449#_c_1435_n N_A_1255_449#_c_1427_n N_A_1255_449#_c_1428_n
+ N_A_1255_449#_c_1429_n N_A_1255_449#_c_1436_n N_A_1255_449#_c_1430_n
+ N_A_1255_449#_c_1438_n N_A_1255_449#_c_1439_n N_A_1255_449#_c_1431_n
+ N_A_1255_449#_c_1432_n PM_SKY130_FD_SC_LP__DFRTP_4%A_1255_449#
x_PM_SKY130_FD_SC_LP__DFRTP_4%A_1891_47# N_A_1891_47#_M1035_s
+ N_A_1891_47#_M1011_s N_A_1891_47#_M1004_g N_A_1891_47#_M1005_g
+ N_A_1891_47#_M1006_g N_A_1891_47#_M1017_g N_A_1891_47#_M1015_g
+ N_A_1891_47#_M1026_g N_A_1891_47#_M1029_g N_A_1891_47#_M1037_g
+ N_A_1891_47#_c_1545_n N_A_1891_47#_c_1546_n N_A_1891_47#_c_1547_n
+ N_A_1891_47#_c_1548_n N_A_1891_47#_c_1549_n
+ PM_SKY130_FD_SC_LP__DFRTP_4%A_1891_47#
x_PM_SKY130_FD_SC_LP__DFRTP_4%VPWR N_VPWR_M1036_d N_VPWR_M1034_d N_VPWR_M1000_d
+ N_VPWR_M1027_s N_VPWR_M1016_d N_VPWR_M1030_d N_VPWR_M1011_d N_VPWR_M1017_d
+ N_VPWR_M1037_d N_VPWR_c_1641_n N_VPWR_c_1642_n N_VPWR_c_1643_n N_VPWR_c_1644_n
+ N_VPWR_c_1645_n N_VPWR_c_1646_n N_VPWR_c_1647_n N_VPWR_c_1648_n
+ N_VPWR_c_1649_n N_VPWR_c_1650_n N_VPWR_c_1651_n N_VPWR_c_1652_n VPWR
+ N_VPWR_c_1653_n N_VPWR_c_1654_n N_VPWR_c_1655_n N_VPWR_c_1656_n
+ N_VPWR_c_1657_n N_VPWR_c_1658_n N_VPWR_c_1659_n N_VPWR_c_1660_n
+ N_VPWR_c_1661_n N_VPWR_c_1662_n N_VPWR_c_1663_n N_VPWR_c_1664_n
+ N_VPWR_c_1665_n N_VPWR_c_1666_n N_VPWR_c_1640_n
+ PM_SKY130_FD_SC_LP__DFRTP_4%VPWR
x_PM_SKY130_FD_SC_LP__DFRTP_4%A_340_535# N_A_340_535#_M1018_d
+ N_A_340_535#_M1034_s N_A_340_535#_M1023_d N_A_340_535#_c_1807_n
+ N_A_340_535#_c_1808_n N_A_340_535#_c_1809_n N_A_340_535#_c_1810_n
+ N_A_340_535#_c_1811_n N_A_340_535#_c_1805_n N_A_340_535#_c_1813_n
+ N_A_340_535#_c_1814_n N_A_340_535#_c_1806_n N_A_340_535#_c_1815_n
+ PM_SKY130_FD_SC_LP__DFRTP_4%A_340_535#
x_PM_SKY130_FD_SC_LP__DFRTP_4%Q N_Q_M1004_d N_Q_M1015_d N_Q_M1005_s N_Q_M1026_s
+ N_Q_c_1941_p N_Q_c_1927_n N_Q_c_1886_n N_Q_c_1887_n N_Q_c_1891_n N_Q_c_1892_n
+ N_Q_c_1932_n N_Q_c_1888_n N_Q_c_1893_n N_Q_c_1889_n N_Q_c_1890_n N_Q_c_1895_n
+ Q N_Q_c_1923_n PM_SKY130_FD_SC_LP__DFRTP_4%Q
x_PM_SKY130_FD_SC_LP__DFRTP_4%VGND N_VGND_M1020_d N_VGND_M1022_s N_VGND_M1010_d
+ N_VGND_M1019_d N_VGND_M1035_d N_VGND_M1006_s N_VGND_M1029_s N_VGND_c_1947_n
+ N_VGND_c_1948_n N_VGND_c_1949_n N_VGND_c_1950_n N_VGND_c_1951_n
+ N_VGND_c_1952_n N_VGND_c_1953_n N_VGND_c_1954_n N_VGND_c_1955_n
+ N_VGND_c_1956_n N_VGND_c_1957_n N_VGND_c_1958_n N_VGND_c_1959_n VGND
+ N_VGND_c_1960_n N_VGND_c_1961_n N_VGND_c_1962_n N_VGND_c_1963_n
+ N_VGND_c_1964_n N_VGND_c_1965_n N_VGND_c_1966_n N_VGND_c_1967_n
+ PM_SKY130_FD_SC_LP__DFRTP_4%VGND
cc_1 VNB N_CLK_M1020_g 0.0497375f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.66
cc_2 VNB N_CLK_c_264_n 0.00971656f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.89
cc_3 VNB CLK 0.0205061f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_CLK_c_266_n 0.0185755f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.535
cc_5 VNB N_A_27_90#_M1008_g 0.0202499f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_6 VNB N_A_27_90#_M1001_g 0.00513137f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.535
cc_7 VNB N_A_27_90#_c_303_n 0.0141221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_90#_c_304_n 0.00764055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_90#_c_305_n 0.00973086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_90#_c_306_n 0.00360493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_90#_c_307_n 0.0903283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_90#_c_308_n 0.0135882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_90#_c_309_n 0.00269017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_90#_c_310_n 0.00549724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_90#_c_311_n 0.0138316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_90#_c_312_n 0.00412132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_90#_c_313_n 8.63915e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_90#_c_314_n 0.00852359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_90#_c_315_n 0.00120345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_90#_c_316_n 0.0122223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_90#_c_317_n 0.00161333f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_90#_c_318_n 0.00414135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_90#_c_319_n 0.0104681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_90#_c_320_n 0.00161919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_90#_c_321_n 0.00121758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_90#_c_322_n 6.54343e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_90#_c_323_n 0.00286788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_90#_c_324_n 0.00242282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_90#_c_325_n 0.0348187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_90#_c_326_n 0.0027664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_90#_c_327_n 9.32761e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_90#_c_328_n 0.00328252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_90#_c_329_n 0.00557231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_90#_c_330_n 9.82692e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_90#_c_331_n 0.0479345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_90#_c_332_n 0.0194631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_90#_c_333_n 0.0169996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_D_M1018_g 0.0339627f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.535
cc_39 VNB N_D_c_595_n 0.00951706f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.89
cc_40 VNB N_D_c_596_n 0.0223791f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_41 VNB D 0.00246631f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_42 VNB N_A_216_462#_M1031_g 0.0155049f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=2.04
cc_43 VNB N_A_216_462#_M1012_g 0.0283739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_216_462#_c_649_n 0.03328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_216_462#_c_650_n 0.00823988f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.535
cc_46 VNB N_A_216_462#_c_651_n 0.0271485f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.535
cc_47 VNB N_A_216_462#_c_652_n 0.0125938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_216_462#_c_653_n 0.0376319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_216_462#_c_654_n 0.00303931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_731_405#_M1033_g 0.0158512f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_51 VNB N_A_731_405#_c_869_n 0.0219605f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.535
cc_52 VNB N_A_731_405#_c_870_n 2.57998e-19 $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.535
cc_53 VNB N_A_731_405#_c_871_n 0.0160001f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.295
cc_54 VNB N_A_731_405#_c_872_n 0.00918377f $X=-0.19 $Y=-0.245 $X2=0.277
+ $Y2=1.535
cc_55 VNB N_A_731_405#_c_873_n 0.0158062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_731_405#_c_874_n 0.00196249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_731_405#_c_875_n 0.00250639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_M1034_g 0.089689f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.66
cc_59 VNB N_RESET_B_c_979_n 0.0245735f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.04
cc_60 VNB N_RESET_B_c_980_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.63
cc_61 VNB N_RESET_B_M1022_g 0.0298982f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.535
cc_62 VNB N_RESET_B_c_982_n 0.166329f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.89
cc_63 VNB N_RESET_B_M1010_g 0.0544458f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.535
cc_64 VNB N_RESET_B_M1003_g 0.0321758f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=2.035
cc_65 VNB N_RESET_B_c_985_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_RESET_B_c_986_n 0.00251358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_RESET_B_c_987_n 7.90281e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_RESET_B_c_988_n 0.0144745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_RESET_B_c_989_n 0.00417218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_RESET_B_c_990_n 0.0153375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_RESET_B_c_991_n 0.00349668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB RESET_B 2.04008e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_595_535#_c_1187_n 0.0147931f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.89
cc_74 VNB N_A_595_535#_c_1188_n 0.0200232f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.89
cc_75 VNB N_A_595_535#_c_1189_n 0.0136084f $X=-0.19 $Y=-0.245 $X2=0.277
+ $Y2=1.665
cc_76 VNB N_A_595_535#_c_1190_n 0.00377241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_595_535#_c_1191_n 3.13343e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_595_535#_c_1192_n 0.0450959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1475_426#_M1019_g 0.0528885f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=2.04
cc_80 VNB N_A_1475_426#_c_1335_n 0.00969516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1475_426#_c_1336_n 0.00778772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1255_449#_c_1422_n 0.0189046f $X=-0.19 $Y=-0.245 $X2=0.575
+ $Y2=2.63
cc_83 VNB N_A_1255_449#_c_1423_n 0.0494803f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_84 VNB N_A_1255_449#_c_1424_n 0.0200415f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_85 VNB N_A_1255_449#_M1011_g 0.017708f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.535
cc_86 VNB N_A_1255_449#_c_1426_n 0.00981073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1255_449#_c_1427_n 0.00539297f $X=-0.19 $Y=-0.245 $X2=0.277
+ $Y2=1.665
cc_88 VNB N_A_1255_449#_c_1428_n 0.00325236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1255_449#_c_1429_n 0.0525326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1255_449#_c_1430_n 0.0248113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1255_449#_c_1431_n 0.00241414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1255_449#_c_1432_n 0.00265534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1891_47#_M1004_g 0.0237277f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.535
cc_94 VNB N_A_1891_47#_M1006_g 0.0217542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1891_47#_M1015_g 0.0219461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1891_47#_M1029_g 0.0265001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1891_47#_c_1545_n 0.0029066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1891_47#_c_1546_n 0.00132235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1891_47#_c_1547_n 0.00777331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1891_47#_c_1548_n 0.00144472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1891_47#_c_1549_n 0.0711048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VPWR_c_1640_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_340_535#_c_1805_n 0.00393894f $X=-0.19 $Y=-0.245 $X2=0.277
+ $Y2=1.295
cc_104 VNB N_A_340_535#_c_1806_n 0.00230898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_Q_c_1886_n 0.00264117f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.295
cc_106 VNB N_Q_c_1887_n 0.00369286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_Q_c_1888_n 0.00854411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_Q_c_1889_n 0.0194203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_Q_c_1890_n 0.00186402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1947_n 0.0119538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1948_n 0.00822193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1949_n 0.0273867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1950_n 0.00803802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1951_n 0.0017733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1952_n 0.0106846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1953_n 0.029659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1954_n 0.0334322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1955_n 0.00326264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1956_n 0.013185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1957_n 0.0667911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1958_n 0.0483521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1959_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1960_n 0.0173343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1961_n 0.0644213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1962_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1963_n 0.0151002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1964_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1965_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1966_n 0.00407307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1967_n 0.62173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VPB N_CLK_M1036_g 0.0327465f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.63
cc_132 VPB N_CLK_c_264_n 0.0202328f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.89
cc_133 VPB N_CLK_c_269_n 0.0275411f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.04
cc_134 VPB CLK 0.0256406f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_135 VPB N_A_27_90#_M1013_g 0.0493113f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.535
cc_136 VPB N_A_27_90#_M1001_g 0.0640404f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.535
cc_137 VPB N_A_27_90#_M1014_g 0.0287137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_27_90#_c_337_n 0.00431702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_27_90#_c_338_n 0.00499926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_27_90#_c_318_n 4.50957e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_27_90#_c_319_n 0.0294053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_27_90#_c_341_n 0.0302303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_D_M1023_g 0.0337944f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.04
cc_144 VPB N_D_c_595_n 0.00363283f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.89
cc_145 VPB N_D_c_600_n 0.0153624f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.89
cc_146 VPB N_D_c_601_n 0.00747013f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.04
cc_147 VPB N_D_c_596_n 0.019041f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_148 VPB D 0.0047331f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_149 VPB N_A_216_462#_M1009_g 0.0267098f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.535
cc_150 VPB N_A_216_462#_c_651_n 0.0128136f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.535
cc_151 VPB N_A_216_462#_M1028_g 0.027867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_216_462#_c_658_n 0.0114211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_216_462#_c_652_n 0.00582215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_216_462#_c_660_n 0.013772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_216_462#_c_661_n 0.0289972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_216_462#_c_662_n 0.0333467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_216_462#_c_663_n 0.0011327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_216_462#_c_664_n 0.0285852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_216_462#_c_665_n 0.00110575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_216_462#_c_666_n 0.00173429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_216_462#_c_653_n 0.014313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_216_462#_c_654_n 0.00861567f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_216_462#_c_669_n 0.0490388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_216_462#_c_670_n 0.0291399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_731_405#_M1000_g 0.0368349f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.535
cc_166 VPB N_A_731_405#_c_877_n 0.0398609f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.89
cc_167 VPB N_A_731_405#_c_878_n 0.00954399f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.89
cc_168 VPB N_A_731_405#_c_879_n 0.0128103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_731_405#_c_870_n 0.0160307f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.535
cc_170 VPB N_A_731_405#_c_881_n 0.00724852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_731_405#_c_882_n 0.00157769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_RESET_B_M1034_g 0.0722879f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.66
cc_173 VPB N_RESET_B_M1007_g 0.0220246f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_174 VPB N_RESET_B_c_995_n 0.0276477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_RESET_B_c_996_n 0.00784683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_RESET_B_M1010_g 0.0272671f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.535
cc_177 VPB N_RESET_B_M1024_g 0.0304223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_RESET_B_c_986_n 0.0202717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_RESET_B_c_1000_n 0.0153055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_RESET_B_c_1001_n 0.00640675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_RESET_B_c_1002_n 0.00567208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_RESET_B_c_987_n 0.0124126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_RESET_B_c_1004_n 0.0120713f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_RESET_B_c_1005_n 0.0415184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB RESET_B 0.00608824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_595_535#_c_1187_n 0.00608052f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.89
cc_187 VPB N_A_595_535#_M1027_g 0.0226284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_595_535#_c_1195_n 4.64252e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_595_535#_c_1196_n 0.00606564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_595_535#_c_1197_n 0.00196479f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.535
cc_191 VPB N_A_595_535#_c_1198_n 0.0033323f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=2.035
cc_192 VPB N_A_595_535#_c_1199_n 0.00960199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_595_535#_c_1200_n 0.00548296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_595_535#_c_1201_n 0.0102141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_595_535#_c_1202_n 7.07762e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_595_535#_c_1203_n 0.0027461f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_595_535#_c_1204_n 0.0487713f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_1475_426#_M1016_g 0.0232264f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.535
cc_199 VPB N_A_1475_426#_M1019_g 0.0178552f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.04
cc_200 VPB N_A_1475_426#_c_1339_n 0.00225931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1475_426#_c_1340_n 0.00772911f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.535
cc_202 VPB N_A_1475_426#_c_1341_n 8.55813e-19 $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.535
cc_203 VPB N_A_1475_426#_c_1342_n 0.0100699f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.535
cc_204 VPB N_A_1475_426#_c_1336_n 0.013937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1475_426#_c_1344_n 0.00646219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1475_426#_c_1345_n 0.0571377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_1255_449#_M1030_g 0.0447953f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.89
cc_208 VPB N_A_1255_449#_M1011_g 0.0247994f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.535
cc_209 VPB N_A_1255_449#_c_1435_n 0.0185786f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.535
cc_210 VPB N_A_1255_449#_c_1436_n 0.00151731f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_1255_449#_c_1430_n 0.00353037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_1255_449#_c_1438_n 0.00110935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_1255_449#_c_1439_n 0.0102915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_1255_449#_c_1431_n 0.0017132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_1891_47#_M1005_g 0.0200793f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.04
cc_216 VPB N_A_1891_47#_M1017_g 0.0188632f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.535
cc_217 VPB N_A_1891_47#_M1026_g 0.0188424f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=2.035
cc_218 VPB N_A_1891_47#_M1037_g 0.0224211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1891_47#_c_1546_n 0.00379559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_1891_47#_c_1549_n 0.00700947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1641_n 0.0044612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1642_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1643_n 0.00493254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1644_n 0.0181921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1645_n 0.0244837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1646_n 0.0171037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1647_n 0.00716337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1648_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1649_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1650_n 0.0428114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1651_n 0.0191301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1652_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1653_n 0.0199635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1654_n 0.0304606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1655_n 0.0355296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1656_n 0.0306443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1657_n 0.0532488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1658_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1659_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1660_n 0.00576489f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1661_n 0.00436557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1662_n 0.00410386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1663_n 0.0155544f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1664_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1665_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1666_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1640_n 0.114987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_340_535#_c_1807_n 0.00573108f $X=-0.19 $Y=1.655 $X2=0.435
+ $Y2=1.89
cc_249 VPB N_A_340_535#_c_1808_n 0.00643975f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.21
cc_250 VPB N_A_340_535#_c_1809_n 0.00444617f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.58
cc_251 VPB N_A_340_535#_c_1810_n 8.6141e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_340_535#_c_1811_n 0.00519929f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.535
cc_253 VPB N_A_340_535#_c_1805_n 0.00124526f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.295
cc_254 VPB N_A_340_535#_c_1813_n 0.00623484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_340_535#_c_1814_n 0.00147472f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.535
cc_256 VPB N_A_340_535#_c_1815_n 0.00748114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_Q_c_1891_n 0.00304705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_Q_c_1892_n 0.00267972f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.535
cc_259 VPB N_Q_c_1893_n 0.0050492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_Q_c_1889_n 0.00459979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_Q_c_1895_n 0.00144314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 N_CLK_c_264_n N_A_27_90#_M1013_g 0.00675255f $X=0.435 $Y=1.89 $X2=0 $Y2=0
cc_263 N_CLK_c_269_n N_A_27_90#_M1013_g 0.0362579f $X=0.435 $Y=2.04 $X2=0 $Y2=0
cc_264 CLK N_A_27_90#_M1013_g 3.40845e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_265 N_CLK_M1020_g N_A_27_90#_c_304_n 0.0164653f $X=0.475 $Y=0.66 $X2=0 $Y2=0
cc_266 CLK N_A_27_90#_c_304_n 0.00901884f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_267 N_CLK_c_266_n N_A_27_90#_c_304_n 2.06494e-19 $X=0.385 $Y=1.535 $X2=0
+ $Y2=0
cc_268 CLK N_A_27_90#_c_305_n 0.0239327f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_269 N_CLK_c_266_n N_A_27_90#_c_305_n 6.88568e-19 $X=0.385 $Y=1.535 $X2=0
+ $Y2=0
cc_270 N_CLK_M1036_g N_A_27_90#_c_337_n 0.014063f $X=0.575 $Y=2.63 $X2=0 $Y2=0
cc_271 N_CLK_c_269_n N_A_27_90#_c_337_n 0.00124348f $X=0.435 $Y=2.04 $X2=0 $Y2=0
cc_272 CLK N_A_27_90#_c_337_n 0.00114453f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_273 N_CLK_M1020_g N_A_27_90#_c_306_n 0.0030181f $X=0.475 $Y=0.66 $X2=0 $Y2=0
cc_274 CLK N_A_27_90#_c_306_n 0.0478888f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_275 N_CLK_M1020_g N_A_27_90#_c_307_n 0.0347731f $X=0.475 $Y=0.66 $X2=0 $Y2=0
cc_276 CLK N_A_27_90#_c_307_n 4.87302e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_277 N_CLK_c_264_n N_A_27_90#_c_338_n 0.0030181f $X=0.435 $Y=1.89 $X2=0 $Y2=0
cc_278 N_CLK_c_269_n N_A_27_90#_c_338_n 0.00575181f $X=0.435 $Y=2.04 $X2=0 $Y2=0
cc_279 N_CLK_M1020_g N_A_27_90#_c_359_n 0.0024761f $X=0.475 $Y=0.66 $X2=0 $Y2=0
cc_280 N_CLK_M1020_g N_A_27_90#_c_309_n 3.43542e-19 $X=0.475 $Y=0.66 $X2=0 $Y2=0
cc_281 N_CLK_M1036_g N_A_27_90#_c_341_n 4.46816e-19 $X=0.575 $Y=2.63 $X2=0 $Y2=0
cc_282 N_CLK_c_269_n N_A_27_90#_c_341_n 0.00145305f $X=0.435 $Y=2.04 $X2=0 $Y2=0
cc_283 CLK N_A_27_90#_c_341_n 0.0243321f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_284 N_CLK_c_266_n N_A_27_90#_c_323_n 0.0030181f $X=0.385 $Y=1.535 $X2=0 $Y2=0
cc_285 N_CLK_M1020_g N_A_27_90#_c_332_n 0.00459421f $X=0.475 $Y=0.66 $X2=0 $Y2=0
cc_286 N_CLK_M1036_g N_VPWR_c_1641_n 0.010596f $X=0.575 $Y=2.63 $X2=0 $Y2=0
cc_287 N_CLK_M1036_g N_VPWR_c_1653_n 0.0047441f $X=0.575 $Y=2.63 $X2=0 $Y2=0
cc_288 N_CLK_M1036_g N_VPWR_c_1640_n 0.00455844f $X=0.575 $Y=2.63 $X2=0 $Y2=0
cc_289 N_CLK_M1020_g N_VGND_c_1947_n 0.0127451f $X=0.475 $Y=0.66 $X2=0 $Y2=0
cc_290 N_CLK_M1020_g N_VGND_c_1960_n 0.00432588f $X=0.475 $Y=0.66 $X2=0 $Y2=0
cc_291 N_CLK_M1020_g N_VGND_c_1967_n 0.00437282f $X=0.475 $Y=0.66 $X2=0 $Y2=0
cc_292 N_A_27_90#_M1008_g N_D_M1018_g 0.0208168f $X=3.37 $Y=0.805 $X2=0 $Y2=0
cc_293 N_A_27_90#_c_311_n N_D_M1018_g 0.00300275f $X=2.65 $Y=1.17 $X2=0 $Y2=0
cc_294 N_A_27_90#_c_313_n N_D_M1018_g 0.00250038f $X=2.735 $Y=1.085 $X2=0 $Y2=0
cc_295 N_A_27_90#_c_314_n N_D_M1018_g 0.00896519f $X=3.42 $Y=0.45 $X2=0 $Y2=0
cc_296 N_A_27_90#_c_324_n N_D_M1018_g 2.81886e-19 $X=3.46 $Y=1.4 $X2=0 $Y2=0
cc_297 N_A_27_90#_c_326_n N_D_M1018_g 7.75834e-19 $X=3.477 $Y=1.235 $X2=0 $Y2=0
cc_298 N_A_27_90#_c_311_n N_D_c_595_n 0.00456036f $X=2.65 $Y=1.17 $X2=0 $Y2=0
cc_299 N_A_27_90#_c_311_n N_D_c_596_n 0.00382277f $X=2.65 $Y=1.17 $X2=0 $Y2=0
cc_300 N_A_27_90#_c_325_n N_D_c_596_n 0.0208168f $X=3.46 $Y=1.4 $X2=0 $Y2=0
cc_301 N_A_27_90#_M1001_g D 3.60455e-19 $X=3.37 $Y=2.885 $X2=0 $Y2=0
cc_302 N_A_27_90#_c_311_n D 0.0530913f $X=2.65 $Y=1.17 $X2=0 $Y2=0
cc_303 N_A_27_90#_c_312_n D 0.00638629f $X=2.065 $Y=1.17 $X2=0 $Y2=0
cc_304 N_A_27_90#_c_308_n N_A_216_462#_M1021_d 0.00247599f $X=1.895 $Y=0.375
+ $X2=-0.19 $Y2=-0.245
cc_305 N_A_27_90#_M1001_g N_A_216_462#_M1009_g 0.0188069f $X=3.37 $Y=2.885 $X2=0
+ $Y2=0
cc_306 N_A_27_90#_M1008_g N_A_216_462#_M1031_g 0.00818352f $X=3.37 $Y=0.805
+ $X2=0 $Y2=0
cc_307 N_A_27_90#_c_316_n N_A_216_462#_M1031_g 0.00594267f $X=4.14 $Y=0.45 $X2=0
+ $Y2=0
cc_308 N_A_27_90#_c_326_n N_A_216_462#_M1031_g 0.00346734f $X=3.477 $Y=1.235
+ $X2=0 $Y2=0
cc_309 N_A_27_90#_c_328_n N_A_216_462#_M1031_g 0.00455389f $X=4.225 $Y=0.45
+ $X2=0 $Y2=0
cc_310 N_A_27_90#_c_317_n N_A_216_462#_M1012_g 0.00770122f $X=6.315 $Y=0.61
+ $X2=0 $Y2=0
cc_311 N_A_27_90#_c_320_n N_A_216_462#_M1012_g 0.0143476f $X=6.4 $Y=1.245 $X2=0
+ $Y2=0
cc_312 N_A_27_90#_c_386_p N_A_216_462#_M1012_g 0.00588544f $X=6.4 $Y=0.61 $X2=0
+ $Y2=0
cc_313 N_A_27_90#_c_331_n N_A_216_462#_M1012_g 0.0126393f $X=7.26 $Y=0.39 $X2=0
+ $Y2=0
cc_314 N_A_27_90#_c_320_n N_A_216_462#_c_649_n 0.00453387f $X=6.4 $Y=1.245 $X2=0
+ $Y2=0
cc_315 N_A_27_90#_c_321_n N_A_216_462#_c_649_n 0.00500592f $X=7.095 $Y=0.61
+ $X2=0 $Y2=0
cc_316 N_A_27_90#_c_329_n N_A_216_462#_c_649_n 0.00341138f $X=6.4 $Y=1.33 $X2=0
+ $Y2=0
cc_317 N_A_27_90#_c_333_n N_A_216_462#_c_649_n 0.00302283f $X=7.26 $Y=0.555
+ $X2=0 $Y2=0
cc_318 N_A_27_90#_c_319_n N_A_216_462#_c_650_n 0.00573836f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_319 N_A_27_90#_c_320_n N_A_216_462#_c_650_n 0.00174074f $X=6.4 $Y=1.245 $X2=0
+ $Y2=0
cc_320 N_A_27_90#_c_329_n N_A_216_462#_c_650_n 0.00488499f $X=6.4 $Y=1.33 $X2=0
+ $Y2=0
cc_321 N_A_27_90#_c_318_n N_A_216_462#_c_651_n 0.00132033f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_322 N_A_27_90#_c_319_n N_A_216_462#_c_651_n 0.0110177f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_323 N_A_27_90#_c_329_n N_A_216_462#_c_651_n 6.83995e-19 $X=6.4 $Y=1.33 $X2=0
+ $Y2=0
cc_324 N_A_27_90#_M1014_g N_A_216_462#_M1028_g 0.0166905f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_325 N_A_27_90#_M1013_g N_A_216_462#_c_658_n 8.02494e-19 $X=1.005 $Y=2.63
+ $X2=0 $Y2=0
cc_326 N_A_27_90#_c_337_n N_A_216_462#_c_658_n 0.00752788f $X=0.765 $Y=2.385
+ $X2=0 $Y2=0
cc_327 N_A_27_90#_c_338_n N_A_216_462#_c_658_n 0.0010832f $X=0.85 $Y=2.3 $X2=0
+ $Y2=0
cc_328 N_A_27_90#_M1013_g N_A_216_462#_c_652_n 0.0042405f $X=1.005 $Y=2.63 $X2=0
+ $Y2=0
cc_329 N_A_27_90#_c_306_n N_A_216_462#_c_652_n 0.0453681f $X=0.955 $Y=1.145
+ $X2=0 $Y2=0
cc_330 N_A_27_90#_c_307_n N_A_216_462#_c_652_n 0.0206281f $X=0.955 $Y=1.145
+ $X2=0 $Y2=0
cc_331 N_A_27_90#_c_338_n N_A_216_462#_c_652_n 0.00803483f $X=0.85 $Y=2.3 $X2=0
+ $Y2=0
cc_332 N_A_27_90#_c_308_n N_A_216_462#_c_652_n 0.020835f $X=1.895 $Y=0.375 $X2=0
+ $Y2=0
cc_333 N_A_27_90#_c_310_n N_A_216_462#_c_652_n 0.034609f $X=1.98 $Y=1.085 $X2=0
+ $Y2=0
cc_334 N_A_27_90#_c_312_n N_A_216_462#_c_652_n 0.0144391f $X=2.065 $Y=1.17 $X2=0
+ $Y2=0
cc_335 N_A_27_90#_c_322_n N_A_216_462#_c_652_n 0.0129747f $X=0.985 $Y=0.945
+ $X2=0 $Y2=0
cc_336 N_A_27_90#_c_332_n N_A_216_462#_c_652_n 0.00504962f $X=1.09 $Y=0.98 $X2=0
+ $Y2=0
cc_337 N_A_27_90#_M1001_g N_A_216_462#_c_660_n 2.41914e-19 $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_338 N_A_27_90#_M1001_g N_A_216_462#_c_661_n 0.0213414f $X=3.37 $Y=2.885 $X2=0
+ $Y2=0
cc_339 N_A_27_90#_M1001_g N_A_216_462#_c_662_n 0.00247126f $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_340 N_A_27_90#_c_324_n N_A_216_462#_c_662_n 0.00619362f $X=3.46 $Y=1.4 $X2=0
+ $Y2=0
cc_341 N_A_27_90#_c_325_n N_A_216_462#_c_662_n 7.59047e-19 $X=3.46 $Y=1.4 $X2=0
+ $Y2=0
cc_342 N_A_27_90#_M1013_g N_A_216_462#_c_663_n 0.00655112f $X=1.005 $Y=2.63
+ $X2=0 $Y2=0
cc_343 N_A_27_90#_c_338_n N_A_216_462#_c_663_n 0.00660298f $X=0.85 $Y=2.3 $X2=0
+ $Y2=0
cc_344 N_A_27_90#_c_323_n N_A_216_462#_c_663_n 0.00287475f $X=0.985 $Y=1.65
+ $X2=0 $Y2=0
cc_345 N_A_27_90#_M1014_g N_A_216_462#_c_664_n 0.00947506f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_346 N_A_27_90#_c_318_n N_A_216_462#_c_664_n 0.00949841f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_347 N_A_27_90#_c_319_n N_A_216_462#_c_664_n 0.00374175f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_348 N_A_27_90#_c_329_n N_A_216_462#_c_664_n 0.00544468f $X=6.4 $Y=1.33 $X2=0
+ $Y2=0
cc_349 N_A_27_90#_M1008_g N_A_216_462#_c_653_n 0.00245237f $X=3.37 $Y=0.805
+ $X2=0 $Y2=0
cc_350 N_A_27_90#_M1001_g N_A_216_462#_c_653_n 0.00713267f $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_351 N_A_27_90#_c_316_n N_A_216_462#_c_653_n 2.21082e-19 $X=4.14 $Y=0.45 $X2=0
+ $Y2=0
cc_352 N_A_27_90#_c_324_n N_A_216_462#_c_653_n 0.00109024f $X=3.46 $Y=1.4 $X2=0
+ $Y2=0
cc_353 N_A_27_90#_c_325_n N_A_216_462#_c_653_n 0.0202055f $X=3.46 $Y=1.4 $X2=0
+ $Y2=0
cc_354 N_A_27_90#_c_326_n N_A_216_462#_c_653_n 0.00158769f $X=3.477 $Y=1.235
+ $X2=0 $Y2=0
cc_355 N_A_27_90#_M1001_g N_A_216_462#_c_654_n 0.00462832f $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_356 N_A_27_90#_c_325_n N_A_216_462#_c_654_n 0.00117945f $X=3.46 $Y=1.4 $X2=0
+ $Y2=0
cc_357 N_A_27_90#_c_326_n N_A_216_462#_c_654_n 0.0192254f $X=3.477 $Y=1.235
+ $X2=0 $Y2=0
cc_358 N_A_27_90#_M1014_g N_A_216_462#_c_669_n 0.00641221f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_359 N_A_27_90#_c_333_n N_A_216_462#_c_669_n 9.33169e-19 $X=7.26 $Y=0.555
+ $X2=0 $Y2=0
cc_360 N_A_27_90#_M1013_g N_A_216_462#_c_670_n 0.00907032f $X=1.005 $Y=2.63
+ $X2=0 $Y2=0
cc_361 N_A_27_90#_c_307_n N_A_216_462#_c_670_n 0.00853627f $X=0.955 $Y=1.145
+ $X2=0 $Y2=0
cc_362 N_A_27_90#_c_338_n N_A_216_462#_c_670_n 0.0294605f $X=0.85 $Y=2.3 $X2=0
+ $Y2=0
cc_363 N_A_27_90#_c_323_n N_A_216_462#_c_670_n 0.0061886f $X=0.985 $Y=1.65 $X2=0
+ $Y2=0
cc_364 N_A_27_90#_c_317_n N_A_731_405#_M1025_d 0.0117926f $X=6.315 $Y=0.61
+ $X2=-0.19 $Y2=-0.245
cc_365 N_A_27_90#_M1001_g N_A_731_405#_c_878_n 0.0752242f $X=3.37 $Y=2.885 $X2=0
+ $Y2=0
cc_366 N_A_27_90#_c_317_n N_A_731_405#_M1033_g 0.00929099f $X=6.315 $Y=0.61
+ $X2=0 $Y2=0
cc_367 N_A_27_90#_c_328_n N_A_731_405#_M1033_g 0.00165271f $X=4.225 $Y=0.45
+ $X2=0 $Y2=0
cc_368 N_A_27_90#_c_318_n N_A_731_405#_c_872_n 0.00527837f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_369 N_A_27_90#_c_320_n N_A_731_405#_c_872_n 0.00732032f $X=6.4 $Y=1.245 $X2=0
+ $Y2=0
cc_370 N_A_27_90#_c_329_n N_A_731_405#_c_872_n 0.0134739f $X=6.4 $Y=1.33 $X2=0
+ $Y2=0
cc_371 N_A_27_90#_M1014_g N_A_731_405#_c_881_n 0.00204163f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_372 N_A_27_90#_c_318_n N_A_731_405#_c_881_n 0.0215932f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_373 N_A_27_90#_c_319_n N_A_731_405#_c_881_n 0.00296902f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_374 N_A_27_90#_c_317_n N_A_731_405#_c_874_n 0.0264705f $X=6.315 $Y=0.61 $X2=0
+ $Y2=0
cc_375 N_A_27_90#_c_319_n N_A_731_405#_c_874_n 0.00179944f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_376 N_A_27_90#_c_320_n N_A_731_405#_c_874_n 0.0150106f $X=6.4 $Y=1.245 $X2=0
+ $Y2=0
cc_377 N_A_27_90#_c_329_n N_A_731_405#_c_874_n 0.00146464f $X=6.4 $Y=1.33 $X2=0
+ $Y2=0
cc_378 N_A_27_90#_c_318_n N_A_731_405#_c_875_n 0.0143526f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_379 N_A_27_90#_c_319_n N_A_731_405#_c_875_n 3.75974e-19 $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_380 N_A_27_90#_M1014_g N_A_731_405#_c_882_n 0.00456756f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_381 N_A_27_90#_c_318_n N_A_731_405#_c_882_n 8.76771e-19 $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_382 N_A_27_90#_c_319_n N_A_731_405#_c_882_n 0.00252782f $X=6.22 $Y=1.79 $X2=0
+ $Y2=0
cc_383 N_A_27_90#_c_308_n N_RESET_B_M1034_g 0.00700064f $X=1.895 $Y=0.375 $X2=0
+ $Y2=0
cc_384 N_A_27_90#_c_310_n N_RESET_B_M1034_g 0.0174909f $X=1.98 $Y=1.085 $X2=0
+ $Y2=0
cc_385 N_A_27_90#_c_311_n N_RESET_B_M1034_g 0.00715579f $X=2.65 $Y=1.17 $X2=0
+ $Y2=0
cc_386 N_A_27_90#_c_312_n N_RESET_B_M1034_g 0.00531447f $X=2.065 $Y=1.17 $X2=0
+ $Y2=0
cc_387 N_A_27_90#_c_313_n N_RESET_B_M1034_g 5.81808e-19 $X=2.735 $Y=1.085 $X2=0
+ $Y2=0
cc_388 N_A_27_90#_c_332_n N_RESET_B_M1034_g 0.0167945f $X=1.09 $Y=0.98 $X2=0
+ $Y2=0
cc_389 N_A_27_90#_c_310_n N_RESET_B_M1022_g 6.36046e-19 $X=1.98 $Y=1.085 $X2=0
+ $Y2=0
cc_390 N_A_27_90#_c_311_n N_RESET_B_M1022_g 0.00949336f $X=2.65 $Y=1.17 $X2=0
+ $Y2=0
cc_391 N_A_27_90#_c_313_n N_RESET_B_M1022_g 0.00966786f $X=2.735 $Y=1.085 $X2=0
+ $Y2=0
cc_392 N_A_27_90#_c_315_n N_RESET_B_M1022_g 0.00463873f $X=2.82 $Y=0.45 $X2=0
+ $Y2=0
cc_393 N_A_27_90#_M1008_g N_RESET_B_c_982_n 0.0088477f $X=3.37 $Y=0.805 $X2=0
+ $Y2=0
cc_394 N_A_27_90#_c_314_n N_RESET_B_c_982_n 0.00898236f $X=3.42 $Y=0.45 $X2=0
+ $Y2=0
cc_395 N_A_27_90#_c_315_n N_RESET_B_c_982_n 0.00175967f $X=2.82 $Y=0.45 $X2=0
+ $Y2=0
cc_396 N_A_27_90#_c_316_n N_RESET_B_c_982_n 0.00985751f $X=4.14 $Y=0.45 $X2=0
+ $Y2=0
cc_397 N_A_27_90#_c_317_n N_RESET_B_c_982_n 0.00755335f $X=6.315 $Y=0.61 $X2=0
+ $Y2=0
cc_398 N_A_27_90#_c_327_n N_RESET_B_c_982_n 0.00360993f $X=3.505 $Y=0.45 $X2=0
+ $Y2=0
cc_399 N_A_27_90#_c_328_n N_RESET_B_c_982_n 0.00373296f $X=4.225 $Y=0.45 $X2=0
+ $Y2=0
cc_400 N_A_27_90#_c_317_n N_RESET_B_M1010_g 0.0129039f $X=6.315 $Y=0.61 $X2=0
+ $Y2=0
cc_401 N_A_27_90#_c_328_n N_RESET_B_M1010_g 0.00230727f $X=4.225 $Y=0.45 $X2=0
+ $Y2=0
cc_402 N_A_27_90#_M1014_g N_RESET_B_c_1002_n 0.0145844f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_403 N_A_27_90#_M1014_g N_RESET_B_c_1027_n 0.00328972f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_404 N_A_27_90#_c_326_n N_A_595_535#_M1008_d 0.00445368f $X=3.477 $Y=1.235
+ $X2=-0.19 $Y2=-0.245
cc_405 N_A_27_90#_c_319_n N_A_595_535#_c_1187_n 0.00149267f $X=6.22 $Y=1.79
+ $X2=0 $Y2=0
cc_406 N_A_27_90#_c_317_n N_A_595_535#_c_1188_n 0.0168781f $X=6.315 $Y=0.61
+ $X2=0 $Y2=0
cc_407 N_A_27_90#_c_320_n N_A_595_535#_c_1188_n 9.07542e-19 $X=6.4 $Y=1.245
+ $X2=0 $Y2=0
cc_408 N_A_27_90#_M1001_g N_A_595_535#_c_1209_n 0.0104101f $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_409 N_A_27_90#_M1001_g N_A_595_535#_c_1195_n 0.00343186f $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_410 N_A_27_90#_M1001_g N_A_595_535#_c_1197_n 9.92233e-19 $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_411 N_A_27_90#_c_316_n N_A_595_535#_c_1189_n 0.00643524f $X=4.14 $Y=0.45
+ $X2=0 $Y2=0
cc_412 N_A_27_90#_c_317_n N_A_595_535#_c_1189_n 0.0498434f $X=6.315 $Y=0.61
+ $X2=0 $Y2=0
cc_413 N_A_27_90#_c_328_n N_A_595_535#_c_1189_n 0.00814735f $X=4.225 $Y=0.45
+ $X2=0 $Y2=0
cc_414 N_A_27_90#_M1008_g N_A_595_535#_c_1190_n 9.16601e-19 $X=3.37 $Y=0.805
+ $X2=0 $Y2=0
cc_415 N_A_27_90#_c_316_n N_A_595_535#_c_1190_n 0.0134126f $X=4.14 $Y=0.45 $X2=0
+ $Y2=0
cc_416 N_A_27_90#_c_326_n N_A_595_535#_c_1190_n 0.0243457f $X=3.477 $Y=1.235
+ $X2=0 $Y2=0
cc_417 N_A_27_90#_c_317_n N_A_595_535#_c_1191_n 0.0202488f $X=6.315 $Y=0.61
+ $X2=0 $Y2=0
cc_418 N_A_27_90#_M1014_g N_A_595_535#_c_1204_n 0.0427077f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_419 N_A_27_90#_c_319_n N_A_595_535#_c_1204_n 0.00480366f $X=6.22 $Y=1.79
+ $X2=0 $Y2=0
cc_420 N_A_27_90#_c_317_n N_A_595_535#_c_1192_n 0.00126839f $X=6.315 $Y=0.61
+ $X2=0 $Y2=0
cc_421 N_A_27_90#_c_330_n N_A_1475_426#_M1019_g 0.00146618f $X=7.26 $Y=0.39
+ $X2=0 $Y2=0
cc_422 N_A_27_90#_c_331_n N_A_1475_426#_M1019_g 0.00120831f $X=7.26 $Y=0.39
+ $X2=0 $Y2=0
cc_423 N_A_27_90#_c_333_n N_A_1475_426#_M1019_g 0.0201722f $X=7.26 $Y=0.555
+ $X2=0 $Y2=0
cc_424 N_A_27_90#_c_320_n N_A_1255_449#_M1012_d 0.00363786f $X=6.4 $Y=1.245
+ $X2=-0.19 $Y2=-0.245
cc_425 N_A_27_90#_c_321_n N_A_1255_449#_M1012_d 0.0174342f $X=7.095 $Y=0.61
+ $X2=-0.19 $Y2=-0.245
cc_426 N_A_27_90#_c_386_p N_A_1255_449#_M1012_d 6.65705e-19 $X=6.4 $Y=0.61
+ $X2=-0.19 $Y2=-0.245
cc_427 N_A_27_90#_c_318_n N_A_1255_449#_c_1428_n 0.00853212f $X=6.22 $Y=1.79
+ $X2=0 $Y2=0
cc_428 N_A_27_90#_c_321_n N_A_1255_449#_c_1429_n 0.00328962f $X=7.095 $Y=0.61
+ $X2=0 $Y2=0
cc_429 N_A_27_90#_c_330_n N_A_1255_449#_c_1429_n 0.0118309f $X=7.26 $Y=0.39
+ $X2=0 $Y2=0
cc_430 N_A_27_90#_c_331_n N_A_1255_449#_c_1429_n 8.14936e-19 $X=7.26 $Y=0.39
+ $X2=0 $Y2=0
cc_431 N_A_27_90#_c_333_n N_A_1255_449#_c_1429_n 0.00964702f $X=7.26 $Y=0.555
+ $X2=0 $Y2=0
cc_432 N_A_27_90#_c_319_n N_A_1255_449#_c_1438_n 0.00167795f $X=6.22 $Y=1.79
+ $X2=0 $Y2=0
cc_433 N_A_27_90#_M1014_g N_A_1255_449#_c_1439_n 0.0034027f $X=6.2 $Y=2.665
+ $X2=0 $Y2=0
cc_434 N_A_27_90#_c_318_n N_A_1255_449#_c_1439_n 0.0136457f $X=6.22 $Y=1.79
+ $X2=0 $Y2=0
cc_435 N_A_27_90#_c_319_n N_A_1255_449#_c_1439_n 0.00146541f $X=6.22 $Y=1.79
+ $X2=0 $Y2=0
cc_436 N_A_27_90#_c_318_n N_A_1255_449#_c_1431_n 0.0130492f $X=6.22 $Y=1.79
+ $X2=0 $Y2=0
cc_437 N_A_27_90#_c_319_n N_A_1255_449#_c_1431_n 0.00113649f $X=6.22 $Y=1.79
+ $X2=0 $Y2=0
cc_438 N_A_27_90#_c_320_n N_A_1255_449#_c_1432_n 0.0290152f $X=6.4 $Y=1.245
+ $X2=0 $Y2=0
cc_439 N_A_27_90#_c_321_n N_A_1255_449#_c_1432_n 0.0255886f $X=7.095 $Y=0.61
+ $X2=0 $Y2=0
cc_440 N_A_27_90#_c_329_n N_A_1255_449#_c_1432_n 0.0131101f $X=6.4 $Y=1.33 $X2=0
+ $Y2=0
cc_441 N_A_27_90#_c_333_n N_A_1255_449#_c_1432_n 0.00722415f $X=7.26 $Y=0.555
+ $X2=0 $Y2=0
cc_442 N_A_27_90#_c_337_n N_VPWR_M1036_d 0.00177916f $X=0.765 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_443 N_A_27_90#_M1013_g N_VPWR_c_1641_n 0.00945254f $X=1.005 $Y=2.63 $X2=0
+ $Y2=0
cc_444 N_A_27_90#_c_337_n N_VPWR_c_1641_n 0.0161463f $X=0.765 $Y=2.385 $X2=0
+ $Y2=0
cc_445 N_A_27_90#_c_341_n N_VPWR_c_1641_n 0.0130269f $X=0.36 $Y=2.465 $X2=0
+ $Y2=0
cc_446 N_A_27_90#_c_341_n N_VPWR_c_1653_n 0.0110559f $X=0.36 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_A_27_90#_M1013_g N_VPWR_c_1654_n 0.00550536f $X=1.005 $Y=2.63 $X2=0
+ $Y2=0
cc_448 N_A_27_90#_M1001_g N_VPWR_c_1655_n 0.00357877f $X=3.37 $Y=2.885 $X2=0
+ $Y2=0
cc_449 N_A_27_90#_M1014_g N_VPWR_c_1657_n 0.00374419f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_450 N_A_27_90#_M1013_g N_VPWR_c_1640_n 0.005282f $X=1.005 $Y=2.63 $X2=0 $Y2=0
cc_451 N_A_27_90#_M1001_g N_VPWR_c_1640_n 0.0053023f $X=3.37 $Y=2.885 $X2=0
+ $Y2=0
cc_452 N_A_27_90#_M1014_g N_VPWR_c_1640_n 0.00672312f $X=6.2 $Y=2.665 $X2=0
+ $Y2=0
cc_453 N_A_27_90#_c_337_n N_VPWR_c_1640_n 0.00636177f $X=0.765 $Y=2.385 $X2=0
+ $Y2=0
cc_454 N_A_27_90#_c_341_n N_VPWR_c_1640_n 0.00946638f $X=0.36 $Y=2.465 $X2=0
+ $Y2=0
cc_455 N_A_27_90#_M1013_g N_A_340_535#_c_1807_n 0.00271682f $X=1.005 $Y=2.63
+ $X2=0 $Y2=0
cc_456 N_A_27_90#_M1001_g N_A_340_535#_c_1811_n 0.00696726f $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_457 N_A_27_90#_M1008_g N_A_340_535#_c_1805_n 0.00584287f $X=3.37 $Y=0.805
+ $X2=0 $Y2=0
cc_458 N_A_27_90#_c_311_n N_A_340_535#_c_1805_n 0.0138832f $X=2.65 $Y=1.17 $X2=0
+ $Y2=0
cc_459 N_A_27_90#_c_324_n N_A_340_535#_c_1805_n 0.0244517f $X=3.46 $Y=1.4 $X2=0
+ $Y2=0
cc_460 N_A_27_90#_c_326_n N_A_340_535#_c_1805_n 0.0105421f $X=3.477 $Y=1.235
+ $X2=0 $Y2=0
cc_461 N_A_27_90#_M1001_g N_A_340_535#_c_1813_n 0.0153914f $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_462 N_A_27_90#_M1008_g N_A_340_535#_c_1806_n 2.93951e-19 $X=3.37 $Y=0.805
+ $X2=0 $Y2=0
cc_463 N_A_27_90#_c_313_n N_A_340_535#_c_1806_n 0.0155081f $X=2.735 $Y=1.085
+ $X2=0 $Y2=0
cc_464 N_A_27_90#_c_314_n N_A_340_535#_c_1806_n 0.015741f $X=3.42 $Y=0.45 $X2=0
+ $Y2=0
cc_465 N_A_27_90#_c_326_n N_A_340_535#_c_1806_n 0.0127488f $X=3.477 $Y=1.235
+ $X2=0 $Y2=0
cc_466 N_A_27_90#_M1001_g N_A_340_535#_c_1815_n 0.0113483f $X=3.37 $Y=2.885
+ $X2=0 $Y2=0
cc_467 N_A_27_90#_c_324_n N_A_340_535#_c_1815_n 0.00382326f $X=3.46 $Y=1.4 $X2=0
+ $Y2=0
cc_468 N_A_27_90#_c_304_n N_VGND_M1020_d 0.00164866f $X=0.765 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_469 N_A_27_90#_c_359_n N_VGND_M1020_d 0.0062739f $X=1.12 $Y=0.86 $X2=-0.19
+ $Y2=-0.245
cc_470 N_A_27_90#_c_322_n N_VGND_M1020_d 0.00521218f $X=0.985 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_471 N_A_27_90#_c_317_n N_VGND_M1010_d 0.00955367f $X=6.315 $Y=0.61 $X2=0
+ $Y2=0
cc_472 N_A_27_90#_c_304_n N_VGND_c_1947_n 0.0143081f $X=0.765 $Y=0.945 $X2=0
+ $Y2=0
cc_473 N_A_27_90#_c_307_n N_VGND_c_1947_n 4.30879e-19 $X=0.955 $Y=1.145 $X2=0
+ $Y2=0
cc_474 N_A_27_90#_c_359_n N_VGND_c_1947_n 0.0175818f $X=1.12 $Y=0.86 $X2=0 $Y2=0
cc_475 N_A_27_90#_c_309_n N_VGND_c_1947_n 0.0150371f $X=1.205 $Y=0.375 $X2=0
+ $Y2=0
cc_476 N_A_27_90#_c_322_n N_VGND_c_1947_n 0.00872686f $X=0.985 $Y=0.945 $X2=0
+ $Y2=0
cc_477 N_A_27_90#_c_332_n N_VGND_c_1947_n 7.97449e-19 $X=1.09 $Y=0.98 $X2=0
+ $Y2=0
cc_478 N_A_27_90#_c_308_n N_VGND_c_1948_n 0.0139514f $X=1.895 $Y=0.375 $X2=0
+ $Y2=0
cc_479 N_A_27_90#_c_310_n N_VGND_c_1948_n 0.0334845f $X=1.98 $Y=1.085 $X2=0
+ $Y2=0
cc_480 N_A_27_90#_c_311_n N_VGND_c_1948_n 0.0187093f $X=2.65 $Y=1.17 $X2=0 $Y2=0
cc_481 N_A_27_90#_c_313_n N_VGND_c_1948_n 0.0151908f $X=2.735 $Y=1.085 $X2=0
+ $Y2=0
cc_482 N_A_27_90#_c_315_n N_VGND_c_1948_n 0.0139503f $X=2.82 $Y=0.45 $X2=0 $Y2=0
cc_483 N_A_27_90#_c_330_n N_VGND_c_1949_n 0.0167408f $X=7.26 $Y=0.39 $X2=0 $Y2=0
cc_484 N_A_27_90#_c_331_n N_VGND_c_1949_n 0.00584021f $X=7.26 $Y=0.39 $X2=0
+ $Y2=0
cc_485 N_A_27_90#_c_308_n N_VGND_c_1954_n 0.0460633f $X=1.895 $Y=0.375 $X2=0
+ $Y2=0
cc_486 N_A_27_90#_c_309_n N_VGND_c_1954_n 0.00997274f $X=1.205 $Y=0.375 $X2=0
+ $Y2=0
cc_487 N_A_27_90#_c_332_n N_VGND_c_1954_n 8.46661e-19 $X=1.09 $Y=0.98 $X2=0
+ $Y2=0
cc_488 N_A_27_90#_c_317_n N_VGND_c_1956_n 0.0240775f $X=6.315 $Y=0.61 $X2=0
+ $Y2=0
cc_489 N_A_27_90#_c_314_n N_VGND_c_1957_n 0.0227929f $X=3.42 $Y=0.45 $X2=0 $Y2=0
cc_490 N_A_27_90#_c_315_n N_VGND_c_1957_n 0.00713683f $X=2.82 $Y=0.45 $X2=0
+ $Y2=0
cc_491 N_A_27_90#_c_316_n N_VGND_c_1957_n 0.0209072f $X=4.14 $Y=0.45 $X2=0 $Y2=0
cc_492 N_A_27_90#_c_317_n N_VGND_c_1957_n 0.0178722f $X=6.315 $Y=0.61 $X2=0
+ $Y2=0
cc_493 N_A_27_90#_c_327_n N_VGND_c_1957_n 0.00714759f $X=3.505 $Y=0.45 $X2=0
+ $Y2=0
cc_494 N_A_27_90#_c_328_n N_VGND_c_1957_n 0.00671135f $X=4.225 $Y=0.45 $X2=0
+ $Y2=0
cc_495 N_A_27_90#_c_303_n N_VGND_c_1960_n 0.00675374f $X=0.26 $Y=0.66 $X2=0
+ $Y2=0
cc_496 N_A_27_90#_c_317_n N_VGND_c_1961_n 0.0169129f $X=6.315 $Y=0.61 $X2=0
+ $Y2=0
cc_497 N_A_27_90#_c_321_n N_VGND_c_1961_n 0.0139155f $X=7.095 $Y=0.61 $X2=0
+ $Y2=0
cc_498 N_A_27_90#_c_386_p N_VGND_c_1961_n 0.00348025f $X=6.4 $Y=0.61 $X2=0 $Y2=0
cc_499 N_A_27_90#_c_330_n N_VGND_c_1961_n 0.0216732f $X=7.26 $Y=0.39 $X2=0 $Y2=0
cc_500 N_A_27_90#_c_331_n N_VGND_c_1961_n 0.00603306f $X=7.26 $Y=0.39 $X2=0
+ $Y2=0
cc_501 N_A_27_90#_c_303_n N_VGND_c_1967_n 0.00857643f $X=0.26 $Y=0.66 $X2=0
+ $Y2=0
cc_502 N_A_27_90#_c_304_n N_VGND_c_1967_n 0.00610431f $X=0.765 $Y=0.945 $X2=0
+ $Y2=0
cc_503 N_A_27_90#_c_308_n N_VGND_c_1967_n 0.0314089f $X=1.895 $Y=0.375 $X2=0
+ $Y2=0
cc_504 N_A_27_90#_c_309_n N_VGND_c_1967_n 0.00649523f $X=1.205 $Y=0.375 $X2=0
+ $Y2=0
cc_505 N_A_27_90#_c_314_n N_VGND_c_1967_n 0.0185806f $X=3.42 $Y=0.45 $X2=0 $Y2=0
cc_506 N_A_27_90#_c_315_n N_VGND_c_1967_n 0.00550964f $X=2.82 $Y=0.45 $X2=0
+ $Y2=0
cc_507 N_A_27_90#_c_316_n N_VGND_c_1967_n 0.0170364f $X=4.14 $Y=0.45 $X2=0 $Y2=0
cc_508 N_A_27_90#_c_317_n N_VGND_c_1967_n 0.0495454f $X=6.315 $Y=0.61 $X2=0
+ $Y2=0
cc_509 N_A_27_90#_c_321_n N_VGND_c_1967_n 0.0189663f $X=7.095 $Y=0.61 $X2=0
+ $Y2=0
cc_510 N_A_27_90#_c_322_n N_VGND_c_1967_n 0.0069759f $X=0.985 $Y=0.945 $X2=0
+ $Y2=0
cc_511 N_A_27_90#_c_327_n N_VGND_c_1967_n 0.00553982f $X=3.505 $Y=0.45 $X2=0
+ $Y2=0
cc_512 N_A_27_90#_c_328_n N_VGND_c_1967_n 0.00532856f $X=4.225 $Y=0.45 $X2=0
+ $Y2=0
cc_513 N_A_27_90#_c_386_p N_VGND_c_1967_n 0.00524566f $X=6.4 $Y=0.61 $X2=0 $Y2=0
cc_514 N_A_27_90#_c_330_n N_VGND_c_1967_n 0.0111121f $X=7.26 $Y=0.39 $X2=0 $Y2=0
cc_515 N_A_27_90#_c_331_n N_VGND_c_1967_n 0.00818129f $X=7.26 $Y=0.39 $X2=0
+ $Y2=0
cc_516 N_A_27_90#_c_317_n A_829_119# 3.26187e-19 $X=6.315 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_517 N_A_27_90#_c_328_n A_829_119# 0.00140072f $X=4.225 $Y=0.45 $X2=-0.19
+ $Y2=-0.245
cc_518 N_A_27_90#_c_317_n A_905_119# 0.00547248f $X=6.315 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_519 N_A_27_90#_c_330_n A_1449_133# 0.00243029f $X=7.26 $Y=0.39 $X2=-0.19
+ $Y2=-0.245
cc_520 N_D_M1023_g N_A_216_462#_M1009_g 0.0222577f $X=2.47 $Y=2.885 $X2=0 $Y2=0
cc_521 D N_A_216_462#_c_652_n 0.023968f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_522 N_D_M1023_g N_A_216_462#_c_660_n 0.00582071f $X=2.47 $Y=2.885 $X2=0 $Y2=0
cc_523 N_D_c_601_n N_A_216_462#_c_660_n 0.00540663f $X=2.455 $Y=2.175 $X2=0
+ $Y2=0
cc_524 N_D_c_596_n N_A_216_462#_c_660_n 0.0030127f $X=2.865 $Y=1.62 $X2=0 $Y2=0
cc_525 D N_A_216_462#_c_660_n 0.0393474f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_526 N_D_c_601_n N_A_216_462#_c_661_n 0.022034f $X=2.455 $Y=2.175 $X2=0 $Y2=0
cc_527 N_D_c_596_n N_A_216_462#_c_661_n 0.0154363f $X=2.865 $Y=1.62 $X2=0 $Y2=0
cc_528 D N_A_216_462#_c_661_n 3.93966e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_529 N_D_c_600_n N_A_216_462#_c_662_n 0.00258899f $X=2.455 $Y=2.025 $X2=0
+ $Y2=0
cc_530 N_D_c_601_n N_A_216_462#_c_662_n 6.51071e-19 $X=2.455 $Y=2.175 $X2=0
+ $Y2=0
cc_531 N_D_c_596_n N_A_216_462#_c_662_n 0.00224147f $X=2.865 $Y=1.62 $X2=0 $Y2=0
cc_532 D N_A_216_462#_c_662_n 0.0229994f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_533 N_D_M1023_g N_RESET_B_M1034_g 0.0310534f $X=2.47 $Y=2.885 $X2=0 $Y2=0
cc_534 N_D_c_595_n N_RESET_B_M1034_g 0.0382716f $X=2.515 $Y=1.62 $X2=0 $Y2=0
cc_535 D N_RESET_B_M1034_g 0.0165715f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_536 N_D_M1018_g N_RESET_B_M1022_g 0.0399708f $X=2.94 $Y=0.805 $X2=0 $Y2=0
cc_537 N_D_c_595_n N_RESET_B_M1022_g 0.00569352f $X=2.515 $Y=1.62 $X2=0 $Y2=0
cc_538 N_D_M1018_g N_RESET_B_c_982_n 0.00884409f $X=2.94 $Y=0.805 $X2=0 $Y2=0
cc_539 N_D_M1023_g N_VPWR_c_1642_n 0.00849262f $X=2.47 $Y=2.885 $X2=0 $Y2=0
cc_540 N_D_M1023_g N_VPWR_c_1655_n 0.00361815f $X=2.47 $Y=2.885 $X2=0 $Y2=0
cc_541 N_D_M1023_g N_VPWR_c_1640_n 0.00436335f $X=2.47 $Y=2.885 $X2=0 $Y2=0
cc_542 N_D_M1023_g N_A_340_535#_c_1808_n 0.0117308f $X=2.47 $Y=2.885 $X2=0 $Y2=0
cc_543 N_D_M1023_g N_A_340_535#_c_1810_n 7.41928e-19 $X=2.47 $Y=2.885 $X2=0
+ $Y2=0
cc_544 N_D_M1018_g N_A_340_535#_c_1805_n 0.0134995f $X=2.94 $Y=0.805 $X2=0 $Y2=0
cc_545 N_D_c_596_n N_A_340_535#_c_1805_n 0.00705165f $X=2.865 $Y=1.62 $X2=0
+ $Y2=0
cc_546 D N_A_340_535#_c_1805_n 0.0223022f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_547 N_D_M1018_g N_A_340_535#_c_1806_n 0.00398809f $X=2.94 $Y=0.805 $X2=0
+ $Y2=0
cc_548 N_D_c_600_n N_A_340_535#_c_1815_n 0.00206655f $X=2.455 $Y=2.025 $X2=0
+ $Y2=0
cc_549 N_D_c_596_n N_A_340_535#_c_1815_n 0.00133386f $X=2.865 $Y=1.62 $X2=0
+ $Y2=0
cc_550 D N_A_340_535#_c_1815_n 0.00899463f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_551 N_A_216_462#_c_662_n N_A_731_405#_c_877_n 5.4917e-19 $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_552 N_A_216_462#_c_664_n N_A_731_405#_c_877_n 0.00275295f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_553 N_A_216_462#_c_665_n N_A_731_405#_c_877_n 7.75352e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_554 N_A_216_462#_c_653_n N_A_731_405#_c_877_n 0.0214173f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_555 N_A_216_462#_c_654_n N_A_731_405#_c_877_n 0.0167426f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_556 N_A_216_462#_c_662_n N_A_731_405#_c_878_n 0.00370358f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_557 N_A_216_462#_M1031_g N_A_731_405#_M1033_g 0.0389088f $X=4.07 $Y=0.805
+ $X2=0 $Y2=0
cc_558 N_A_216_462#_c_664_n N_A_731_405#_c_879_n 9.50914e-19 $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_559 N_A_216_462#_c_654_n N_A_731_405#_c_879_n 7.52708e-19 $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_560 N_A_216_462#_c_653_n N_A_731_405#_c_869_n 0.0213085f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_561 N_A_216_462#_c_664_n N_A_731_405#_c_871_n 0.0119112f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_562 N_A_216_462#_M1012_g N_A_731_405#_c_872_n 0.00161585f $X=6.31 $Y=0.625
+ $X2=0 $Y2=0
cc_563 N_A_216_462#_c_664_n N_A_731_405#_c_881_n 0.0181967f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_564 N_A_216_462#_c_664_n N_A_731_405#_c_915_n 0.00228499f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_565 N_A_216_462#_c_653_n N_A_731_405#_c_915_n 6.0972e-19 $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_566 N_A_216_462#_c_654_n N_A_731_405#_c_915_n 0.0422537f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_567 N_A_216_462#_c_653_n N_A_731_405#_c_873_n 0.0213085f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_568 N_A_216_462#_c_654_n N_A_731_405#_c_873_n 0.00842986f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_569 N_A_216_462#_M1012_g N_A_731_405#_c_874_n 0.00189642f $X=6.31 $Y=0.625
+ $X2=0 $Y2=0
cc_570 N_A_216_462#_c_664_n N_A_731_405#_c_882_n 0.0105047f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_571 N_A_216_462#_c_658_n N_RESET_B_M1034_g 0.00531969f $X=1.22 $Y=2.455 $X2=0
+ $Y2=0
cc_572 N_A_216_462#_c_652_n N_RESET_B_M1034_g 0.0131685f $X=1.55 $Y=0.725 $X2=0
+ $Y2=0
cc_573 N_A_216_462#_c_660_n N_RESET_B_M1034_g 0.0135358f $X=2.92 $Y=2.19 $X2=0
+ $Y2=0
cc_574 N_A_216_462#_c_662_n N_RESET_B_M1034_g 0.00436989f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_575 N_A_216_462#_c_670_n N_RESET_B_M1034_g 0.0065429f $X=1.715 $Y=2.077 $X2=0
+ $Y2=0
cc_576 N_A_216_462#_M1031_g N_RESET_B_c_982_n 0.008856f $X=4.07 $Y=0.805 $X2=0
+ $Y2=0
cc_577 N_A_216_462#_c_664_n N_RESET_B_c_995_n 0.00270504f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_578 N_A_216_462#_c_664_n N_RESET_B_c_996_n 7.70517e-19 $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_579 N_A_216_462#_c_654_n N_RESET_B_c_996_n 3.45673e-19 $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_580 N_A_216_462#_c_664_n N_RESET_B_M1010_g 0.00157056f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_581 N_A_216_462#_c_664_n N_RESET_B_c_1001_n 0.0161882f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_582 N_A_216_462#_M1028_g N_RESET_B_c_1002_n 0.0148089f $X=6.825 $Y=2.65 $X2=0
+ $Y2=0
cc_583 N_A_216_462#_c_666_n N_RESET_B_c_1002_n 0.00816793f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_A_216_462#_c_669_n N_RESET_B_c_1002_n 0.00411986f $X=7 $Y=2.03 $X2=0
+ $Y2=0
cc_585 N_A_216_462#_c_651_n N_RESET_B_c_987_n 0.00465793f $X=6.78 $Y=1.865 $X2=0
+ $Y2=0
cc_586 N_A_216_462#_M1028_g N_RESET_B_c_987_n 0.00506574f $X=6.825 $Y=2.65 $X2=0
+ $Y2=0
cc_587 N_A_216_462#_c_780_p N_RESET_B_c_987_n 0.00200557f $X=6.96 $Y=2.035 $X2=0
+ $Y2=0
cc_588 N_A_216_462#_c_666_n N_RESET_B_c_987_n 0.0173071f $X=6.96 $Y=2.035 $X2=0
+ $Y2=0
cc_589 N_A_216_462#_c_669_n N_RESET_B_c_987_n 0.00254013f $X=7 $Y=2.03 $X2=0
+ $Y2=0
cc_590 N_A_216_462#_c_651_n N_RESET_B_c_989_n 0.00283039f $X=6.78 $Y=1.865 $X2=0
+ $Y2=0
cc_591 N_A_216_462#_c_664_n N_RESET_B_c_1004_n 0.00797342f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_592 N_A_216_462#_c_664_n N_RESET_B_c_1005_n 0.00462978f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_593 N_A_216_462#_M1012_g N_A_595_535#_c_1188_n 0.0121311f $X=6.31 $Y=0.625
+ $X2=0 $Y2=0
cc_594 N_A_216_462#_c_664_n N_A_595_535#_M1027_g 0.00144728f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_595 N_A_216_462#_c_662_n N_A_595_535#_c_1196_n 0.00289247f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_596 N_A_216_462#_c_664_n N_A_595_535#_c_1196_n 0.00289106f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_597 N_A_216_462#_c_665_n N_A_595_535#_c_1196_n 0.00250042f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_598 N_A_216_462#_c_654_n N_A_595_535#_c_1196_n 0.0192919f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_599 N_A_216_462#_c_662_n N_A_595_535#_c_1197_n 0.00659821f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_600 N_A_216_462#_M1031_g N_A_595_535#_c_1189_n 0.00897924f $X=4.07 $Y=0.805
+ $X2=0 $Y2=0
cc_601 N_A_216_462#_c_653_n N_A_595_535#_c_1189_n 0.0015492f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_602 N_A_216_462#_c_654_n N_A_595_535#_c_1189_n 0.0190812f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_603 N_A_216_462#_c_664_n N_A_595_535#_c_1198_n 0.00281881f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_604 N_A_216_462#_c_664_n N_A_595_535#_c_1200_n 0.00566363f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_605 N_A_216_462#_c_665_n N_A_595_535#_c_1200_n 0.00111983f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_606 N_A_216_462#_c_654_n N_A_595_535#_c_1200_n 0.00616652f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_607 N_A_216_462#_c_664_n N_A_595_535#_c_1201_n 0.0247979f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_608 N_A_216_462#_c_664_n N_A_595_535#_c_1202_n 0.00531685f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_609 N_A_216_462#_c_665_n N_A_595_535#_c_1202_n 0.00133654f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_610 N_A_216_462#_c_654_n N_A_595_535#_c_1202_n 0.0117081f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_611 N_A_216_462#_c_653_n N_A_595_535#_c_1190_n 0.00356584f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_612 N_A_216_462#_c_654_n N_A_595_535#_c_1190_n 0.0103718f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_613 N_A_216_462#_c_664_n N_A_595_535#_c_1203_n 0.0128638f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_614 N_A_216_462#_c_664_n N_A_595_535#_c_1204_n 0.00503982f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_615 N_A_216_462#_c_650_n N_A_595_535#_c_1192_n 0.0121311f $X=6.385 $Y=1.235
+ $X2=0 $Y2=0
cc_616 N_A_216_462#_c_669_n N_A_1475_426#_M1019_g 0.00153365f $X=7 $Y=2.03 $X2=0
+ $Y2=0
cc_617 N_A_216_462#_M1028_g N_A_1475_426#_c_1345_n 0.0166692f $X=6.825 $Y=2.65
+ $X2=0 $Y2=0
cc_618 N_A_216_462#_c_669_n N_A_1475_426#_c_1345_n 0.00970227f $X=7 $Y=2.03
+ $X2=0 $Y2=0
cc_619 N_A_216_462#_c_649_n N_A_1255_449#_c_1428_n 0.00362162f $X=6.705 $Y=1.235
+ $X2=0 $Y2=0
cc_620 N_A_216_462#_c_651_n N_A_1255_449#_c_1428_n 0.0156304f $X=6.78 $Y=1.865
+ $X2=0 $Y2=0
cc_621 N_A_216_462#_c_649_n N_A_1255_449#_c_1429_n 3.59505e-19 $X=6.705 $Y=1.235
+ $X2=0 $Y2=0
cc_622 N_A_216_462#_c_666_n N_A_1255_449#_c_1429_n 0.00381486f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_623 N_A_216_462#_c_669_n N_A_1255_449#_c_1429_n 0.00232869f $X=7 $Y=2.03
+ $X2=0 $Y2=0
cc_624 N_A_216_462#_c_664_n N_A_1255_449#_c_1438_n 0.00682612f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_625 N_A_216_462#_c_651_n N_A_1255_449#_c_1439_n 0.00681613f $X=6.78 $Y=1.865
+ $X2=0 $Y2=0
cc_626 N_A_216_462#_M1028_g N_A_1255_449#_c_1439_n 0.0113602f $X=6.825 $Y=2.65
+ $X2=0 $Y2=0
cc_627 N_A_216_462#_c_664_n N_A_1255_449#_c_1439_n 0.0178597f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_628 N_A_216_462#_c_780_p N_A_1255_449#_c_1439_n 0.0025982f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_629 N_A_216_462#_c_666_n N_A_1255_449#_c_1439_n 0.0176016f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_630 N_A_216_462#_c_649_n N_A_1255_449#_c_1431_n 0.00534936f $X=6.705 $Y=1.235
+ $X2=0 $Y2=0
cc_631 N_A_216_462#_c_651_n N_A_1255_449#_c_1431_n 0.00895237f $X=6.78 $Y=1.865
+ $X2=0 $Y2=0
cc_632 N_A_216_462#_c_664_n N_A_1255_449#_c_1431_n 0.00681182f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_633 N_A_216_462#_c_780_p N_A_1255_449#_c_1431_n 9.64342e-19 $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_634 N_A_216_462#_c_666_n N_A_1255_449#_c_1431_n 8.70491e-19 $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_635 N_A_216_462#_M1012_g N_A_1255_449#_c_1432_n 0.00105668f $X=6.31 $Y=0.625
+ $X2=0 $Y2=0
cc_636 N_A_216_462#_c_649_n N_A_1255_449#_c_1432_n 0.00909294f $X=6.705 $Y=1.235
+ $X2=0 $Y2=0
cc_637 N_A_216_462#_c_666_n N_A_1255_449#_c_1432_n 0.00285448f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_638 N_A_216_462#_c_669_n N_A_1255_449#_c_1432_n 0.00233868f $X=7 $Y=2.03
+ $X2=0 $Y2=0
cc_639 N_A_216_462#_c_658_n N_VPWR_c_1641_n 0.012258f $X=1.22 $Y=2.455 $X2=0
+ $Y2=0
cc_640 N_A_216_462#_M1009_g N_VPWR_c_1642_n 0.00121243f $X=2.9 $Y=2.885 $X2=0
+ $Y2=0
cc_641 N_A_216_462#_c_658_n N_VPWR_c_1654_n 0.0114755f $X=1.22 $Y=2.455 $X2=0
+ $Y2=0
cc_642 N_A_216_462#_M1009_g N_VPWR_c_1655_n 0.00435108f $X=2.9 $Y=2.885 $X2=0
+ $Y2=0
cc_643 N_A_216_462#_M1028_g N_VPWR_c_1657_n 0.00364575f $X=6.825 $Y=2.65 $X2=0
+ $Y2=0
cc_644 N_A_216_462#_M1009_g N_VPWR_c_1640_n 0.00626675f $X=2.9 $Y=2.885 $X2=0
+ $Y2=0
cc_645 N_A_216_462#_M1028_g N_VPWR_c_1640_n 0.00514438f $X=6.825 $Y=2.65 $X2=0
+ $Y2=0
cc_646 N_A_216_462#_c_658_n N_VPWR_c_1640_n 0.0101402f $X=1.22 $Y=2.455 $X2=0
+ $Y2=0
cc_647 N_A_216_462#_c_658_n N_A_340_535#_c_1807_n 0.0193427f $X=1.22 $Y=2.455
+ $X2=0 $Y2=0
cc_648 N_A_216_462#_c_660_n N_A_340_535#_c_1808_n 0.0458919f $X=2.92 $Y=2.19
+ $X2=0 $Y2=0
cc_649 N_A_216_462#_c_662_n N_A_340_535#_c_1808_n 0.00329091f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_650 N_A_216_462#_c_658_n N_A_340_535#_c_1809_n 0.0106235f $X=1.22 $Y=2.455
+ $X2=0 $Y2=0
cc_651 N_A_216_462#_c_662_n N_A_340_535#_c_1809_n 0.00147305f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_652 N_A_216_462#_c_670_n N_A_340_535#_c_1809_n 0.0207437f $X=1.715 $Y=2.077
+ $X2=0 $Y2=0
cc_653 N_A_216_462#_M1009_g N_A_340_535#_c_1810_n 0.00137287f $X=2.9 $Y=2.885
+ $X2=0 $Y2=0
cc_654 N_A_216_462#_M1009_g N_A_340_535#_c_1811_n 0.0122106f $X=2.9 $Y=2.885
+ $X2=0 $Y2=0
cc_655 N_A_216_462#_c_660_n N_A_340_535#_c_1811_n 0.0174756f $X=2.92 $Y=2.19
+ $X2=0 $Y2=0
cc_656 N_A_216_462#_c_661_n N_A_340_535#_c_1811_n 0.00279821f $X=2.92 $Y=2.19
+ $X2=0 $Y2=0
cc_657 N_A_216_462#_c_662_n N_A_340_535#_c_1811_n 0.00546278f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_658 N_A_216_462#_c_654_n N_A_340_535#_c_1805_n 0.00499609f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_659 N_A_216_462#_M1009_g N_A_340_535#_c_1813_n 0.00182823f $X=2.9 $Y=2.885
+ $X2=0 $Y2=0
cc_660 N_A_216_462#_c_660_n N_A_340_535#_c_1813_n 0.0156068f $X=2.92 $Y=2.19
+ $X2=0 $Y2=0
cc_661 N_A_216_462#_c_661_n N_A_340_535#_c_1813_n 0.00298967f $X=2.92 $Y=2.19
+ $X2=0 $Y2=0
cc_662 N_A_216_462#_c_662_n N_A_340_535#_c_1813_n 0.0194476f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_663 N_A_216_462#_c_665_n N_A_340_535#_c_1813_n 4.48468e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_664 N_A_216_462#_c_654_n N_A_340_535#_c_1813_n 0.00744978f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_665 N_A_216_462#_c_660_n N_A_340_535#_c_1814_n 0.0179514f $X=2.92 $Y=2.19
+ $X2=0 $Y2=0
cc_666 N_A_216_462#_c_661_n N_A_340_535#_c_1814_n 0.00163896f $X=2.92 $Y=2.19
+ $X2=0 $Y2=0
cc_667 N_A_216_462#_c_662_n N_A_340_535#_c_1814_n 0.00130575f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_668 N_A_216_462#_c_660_n N_A_340_535#_c_1815_n 0.00586662f $X=2.92 $Y=2.19
+ $X2=0 $Y2=0
cc_669 N_A_216_462#_c_661_n N_A_340_535#_c_1815_n 0.00146366f $X=2.92 $Y=2.19
+ $X2=0 $Y2=0
cc_670 N_A_216_462#_c_662_n N_A_340_535#_c_1815_n 0.0105559f $X=3.935 $Y=2.035
+ $X2=0 $Y2=0
cc_671 N_A_216_462#_c_653_n N_A_340_535#_c_1815_n 2.81172e-19 $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_672 N_A_216_462#_c_654_n N_A_340_535#_c_1815_n 0.00682387f $X=4 $Y=1.31 $X2=0
+ $Y2=0
cc_673 N_A_216_462#_M1012_g N_VGND_c_1961_n 0.00355775f $X=6.31 $Y=0.625 $X2=0
+ $Y2=0
cc_674 N_A_216_462#_M1012_g N_VGND_c_1967_n 0.00586935f $X=6.31 $Y=0.625 $X2=0
+ $Y2=0
cc_675 N_A_731_405#_M1033_g N_RESET_B_c_982_n 0.00961525f $X=4.45 $Y=0.805 $X2=0
+ $Y2=0
cc_676 N_A_731_405#_c_870_n N_RESET_B_c_995_n 0.00252959f $X=4.54 $Y=1.815 $X2=0
+ $Y2=0
cc_677 N_A_731_405#_M1000_g N_RESET_B_c_996_n 0.022092f $X=3.73 $Y=2.885 $X2=0
+ $Y2=0
cc_678 N_A_731_405#_c_877_n N_RESET_B_c_996_n 0.0236706f $X=4.375 $Y=2.1 $X2=0
+ $Y2=0
cc_679 N_A_731_405#_M1033_g N_RESET_B_M1010_g 0.0223058f $X=4.45 $Y=0.805 $X2=0
+ $Y2=0
cc_680 N_A_731_405#_c_879_n N_RESET_B_M1010_g 0.0111798f $X=4.45 $Y=2.025 $X2=0
+ $Y2=0
cc_681 N_A_731_405#_c_871_n N_RESET_B_M1010_g 0.0113516f $X=5.785 $Y=1.57 $X2=0
+ $Y2=0
cc_682 N_A_731_405#_c_915_n N_RESET_B_M1010_g 0.00224225f $X=4.54 $Y=1.31 $X2=0
+ $Y2=0
cc_683 N_A_731_405#_c_873_n N_RESET_B_M1010_g 0.0433603f $X=4.54 $Y=1.31 $X2=0
+ $Y2=0
cc_684 N_A_731_405#_M1027_d N_RESET_B_c_1002_n 0.00335981f $X=5.845 $Y=2.245
+ $X2=0 $Y2=0
cc_685 N_A_731_405#_c_882_n N_RESET_B_c_1002_n 0.00633894f $X=5.985 $Y=2.37
+ $X2=0 $Y2=0
cc_686 N_A_731_405#_M1027_d N_RESET_B_c_1027_n 0.00334094f $X=5.845 $Y=2.245
+ $X2=0 $Y2=0
cc_687 N_A_731_405#_c_882_n N_RESET_B_c_1027_n 0.00816299f $X=5.985 $Y=2.37
+ $X2=0 $Y2=0
cc_688 N_A_731_405#_c_871_n N_A_595_535#_c_1187_n 0.0116174f $X=5.785 $Y=1.57
+ $X2=0 $Y2=0
cc_689 N_A_731_405#_c_872_n N_A_595_535#_c_1187_n 0.00276977f $X=5.87 $Y=1.485
+ $X2=0 $Y2=0
cc_690 N_A_731_405#_c_881_n N_A_595_535#_c_1187_n 0.0018697f $X=5.87 $Y=2.205
+ $X2=0 $Y2=0
cc_691 N_A_731_405#_c_874_n N_A_595_535#_c_1188_n 0.002238f $X=5.98 $Y=0.96
+ $X2=0 $Y2=0
cc_692 N_A_731_405#_c_881_n N_A_595_535#_M1027_g 0.00572294f $X=5.87 $Y=2.205
+ $X2=0 $Y2=0
cc_693 N_A_731_405#_c_882_n N_A_595_535#_M1027_g 0.0134996f $X=5.985 $Y=2.37
+ $X2=0 $Y2=0
cc_694 N_A_731_405#_M1000_g N_A_595_535#_c_1209_n 0.00790632f $X=3.73 $Y=2.885
+ $X2=0 $Y2=0
cc_695 N_A_731_405#_M1000_g N_A_595_535#_c_1195_n 0.00453842f $X=3.73 $Y=2.885
+ $X2=0 $Y2=0
cc_696 N_A_731_405#_M1000_g N_A_595_535#_c_1196_n 0.00463674f $X=3.73 $Y=2.885
+ $X2=0 $Y2=0
cc_697 N_A_731_405#_c_877_n N_A_595_535#_c_1196_n 0.00369757f $X=4.375 $Y=2.1
+ $X2=0 $Y2=0
cc_698 N_A_731_405#_M1000_g N_A_595_535#_c_1197_n 0.00454166f $X=3.73 $Y=2.885
+ $X2=0 $Y2=0
cc_699 N_A_731_405#_M1033_g N_A_595_535#_c_1189_n 0.0106254f $X=4.45 $Y=0.805
+ $X2=0 $Y2=0
cc_700 N_A_731_405#_c_871_n N_A_595_535#_c_1189_n 0.0211049f $X=5.785 $Y=1.57
+ $X2=0 $Y2=0
cc_701 N_A_731_405#_c_915_n N_A_595_535#_c_1189_n 0.0251397f $X=4.54 $Y=1.31
+ $X2=0 $Y2=0
cc_702 N_A_731_405#_c_873_n N_A_595_535#_c_1189_n 0.0050863f $X=4.54 $Y=1.31
+ $X2=0 $Y2=0
cc_703 N_A_731_405#_c_877_n N_A_595_535#_c_1198_n 3.05872e-19 $X=4.375 $Y=2.1
+ $X2=0 $Y2=0
cc_704 N_A_731_405#_M1000_g N_A_595_535#_c_1200_n 0.00491689f $X=3.73 $Y=2.885
+ $X2=0 $Y2=0
cc_705 N_A_731_405#_c_877_n N_A_595_535#_c_1200_n 0.00420999f $X=4.375 $Y=2.1
+ $X2=0 $Y2=0
cc_706 N_A_731_405#_c_870_n N_A_595_535#_c_1201_n 0.00198381f $X=4.54 $Y=1.815
+ $X2=0 $Y2=0
cc_707 N_A_731_405#_c_871_n N_A_595_535#_c_1201_n 0.0266744f $X=5.785 $Y=1.57
+ $X2=0 $Y2=0
cc_708 N_A_731_405#_c_915_n N_A_595_535#_c_1201_n 0.0113328f $X=4.54 $Y=1.31
+ $X2=0 $Y2=0
cc_709 N_A_731_405#_c_877_n N_A_595_535#_c_1202_n 0.0022207f $X=4.375 $Y=2.1
+ $X2=0 $Y2=0
cc_710 N_A_731_405#_c_879_n N_A_595_535#_c_1202_n 0.00533284f $X=4.45 $Y=2.025
+ $X2=0 $Y2=0
cc_711 N_A_731_405#_c_870_n N_A_595_535#_c_1202_n 2.6621e-19 $X=4.54 $Y=1.815
+ $X2=0 $Y2=0
cc_712 N_A_731_405#_c_915_n N_A_595_535#_c_1202_n 0.0129823f $X=4.54 $Y=1.31
+ $X2=0 $Y2=0
cc_713 N_A_731_405#_c_871_n N_A_595_535#_c_1191_n 0.0247682f $X=5.785 $Y=1.57
+ $X2=0 $Y2=0
cc_714 N_A_731_405#_c_872_n N_A_595_535#_c_1191_n 0.0179942f $X=5.87 $Y=1.485
+ $X2=0 $Y2=0
cc_715 N_A_731_405#_c_915_n N_A_595_535#_c_1191_n 0.00275057f $X=4.54 $Y=1.31
+ $X2=0 $Y2=0
cc_716 N_A_731_405#_c_874_n N_A_595_535#_c_1191_n 0.0143485f $X=5.98 $Y=0.96
+ $X2=0 $Y2=0
cc_717 N_A_731_405#_c_871_n N_A_595_535#_c_1203_n 0.0222142f $X=5.785 $Y=1.57
+ $X2=0 $Y2=0
cc_718 N_A_731_405#_c_881_n N_A_595_535#_c_1203_n 0.0172928f $X=5.87 $Y=2.205
+ $X2=0 $Y2=0
cc_719 N_A_731_405#_c_871_n N_A_595_535#_c_1204_n 0.00621637f $X=5.785 $Y=1.57
+ $X2=0 $Y2=0
cc_720 N_A_731_405#_c_881_n N_A_595_535#_c_1204_n 0.0071268f $X=5.87 $Y=2.205
+ $X2=0 $Y2=0
cc_721 N_A_731_405#_c_871_n N_A_595_535#_c_1192_n 0.00496465f $X=5.785 $Y=1.57
+ $X2=0 $Y2=0
cc_722 N_A_731_405#_c_872_n N_A_595_535#_c_1192_n 0.00609901f $X=5.87 $Y=1.485
+ $X2=0 $Y2=0
cc_723 N_A_731_405#_c_881_n N_A_1255_449#_c_1439_n 0.00663504f $X=5.87 $Y=2.205
+ $X2=0 $Y2=0
cc_724 N_A_731_405#_c_882_n N_A_1255_449#_c_1439_n 0.00620546f $X=5.985 $Y=2.37
+ $X2=0 $Y2=0
cc_725 N_A_731_405#_M1000_g N_VPWR_c_1643_n 0.00480066f $X=3.73 $Y=2.885 $X2=0
+ $Y2=0
cc_726 N_A_731_405#_M1000_g N_VPWR_c_1655_n 0.00378318f $X=3.73 $Y=2.885 $X2=0
+ $Y2=0
cc_727 N_A_731_405#_M1027_d N_VPWR_c_1640_n 0.00238545f $X=5.845 $Y=2.245 $X2=0
+ $Y2=0
cc_728 N_A_731_405#_M1000_g N_VPWR_c_1640_n 0.00567109f $X=3.73 $Y=2.885 $X2=0
+ $Y2=0
cc_729 N_A_731_405#_c_878_n N_A_340_535#_c_1813_n 0.00242012f $X=3.805 $Y=2.1
+ $X2=0 $Y2=0
cc_730 N_A_731_405#_M1033_g N_VGND_c_1967_n 9.39239e-19 $X=4.45 $Y=0.805 $X2=0
+ $Y2=0
cc_731 N_RESET_B_c_982_n N_A_595_535#_c_1188_n 0.0200893f $X=4.915 $Y=0.18 $X2=0
+ $Y2=0
cc_732 N_RESET_B_M1010_g N_A_595_535#_M1027_g 0.00779598f $X=4.99 $Y=0.735 $X2=0
+ $Y2=0
cc_733 N_RESET_B_c_1001_n N_A_595_535#_M1027_g 0.00975122f $X=5.785 $Y=2.72
+ $X2=0 $Y2=0
cc_734 N_RESET_B_c_1002_n N_A_595_535#_M1027_g 2.26329e-19 $X=7.345 $Y=2.87
+ $X2=0 $Y2=0
cc_735 N_RESET_B_c_1004_n N_A_595_535#_M1027_g 0.00350029f $X=4.9 $Y=2.35 $X2=0
+ $Y2=0
cc_736 N_RESET_B_c_1027_n N_A_595_535#_M1027_g 0.0116451f $X=5.87 $Y=2.72 $X2=0
+ $Y2=0
cc_737 N_RESET_B_M1007_g N_A_595_535#_c_1195_n 5.23904e-19 $X=4.235 $Y=2.885
+ $X2=0 $Y2=0
cc_738 N_RESET_B_M1007_g N_A_595_535#_c_1196_n 0.00787741f $X=4.235 $Y=2.885
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_995_n N_A_595_535#_c_1196_n 2.32245e-19 $X=4.735 $Y=2.46
+ $X2=0 $Y2=0
cc_740 N_RESET_B_c_996_n N_A_595_535#_c_1196_n 0.00321245f $X=4.31 $Y=2.46 $X2=0
+ $Y2=0
cc_741 N_RESET_B_M1010_g N_A_595_535#_c_1189_n 0.0126679f $X=4.99 $Y=0.735 $X2=0
+ $Y2=0
cc_742 N_RESET_B_M1007_g N_A_595_535#_c_1198_n 0.00176517f $X=4.235 $Y=2.885
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_995_n N_A_595_535#_c_1198_n 0.00952325f $X=4.735 $Y=2.46
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_1004_n N_A_595_535#_c_1198_n 0.0175529f $X=4.9 $Y=2.35 $X2=0
+ $Y2=0
cc_745 N_RESET_B_c_1004_n N_A_595_535#_c_1199_n 0.0027251f $X=4.9 $Y=2.35 $X2=0
+ $Y2=0
cc_746 N_RESET_B_c_995_n N_A_595_535#_c_1200_n 0.00497734f $X=4.735 $Y=2.46
+ $X2=0 $Y2=0
cc_747 N_RESET_B_M1010_g N_A_595_535#_c_1200_n 0.00168632f $X=4.99 $Y=0.735
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_1004_n N_A_595_535#_c_1200_n 0.0135891f $X=4.9 $Y=2.35 $X2=0
+ $Y2=0
cc_749 N_RESET_B_c_1005_n N_A_595_535#_c_1200_n 0.00346821f $X=4.9 $Y=2.35 $X2=0
+ $Y2=0
cc_750 N_RESET_B_c_995_n N_A_595_535#_c_1201_n 0.00295943f $X=4.735 $Y=2.46
+ $X2=0 $Y2=0
cc_751 N_RESET_B_M1010_g N_A_595_535#_c_1201_n 0.0101089f $X=4.99 $Y=0.735 $X2=0
+ $Y2=0
cc_752 N_RESET_B_c_1001_n N_A_595_535#_c_1201_n 0.00406494f $X=5.785 $Y=2.72
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_1004_n N_A_595_535#_c_1201_n 0.0215683f $X=4.9 $Y=2.35 $X2=0
+ $Y2=0
cc_754 N_RESET_B_c_1005_n N_A_595_535#_c_1201_n 0.00435516f $X=4.9 $Y=2.35 $X2=0
+ $Y2=0
cc_755 N_RESET_B_M1010_g N_A_595_535#_c_1191_n 0.0019628f $X=4.99 $Y=0.735 $X2=0
+ $Y2=0
cc_756 N_RESET_B_M1010_g N_A_595_535#_c_1203_n 7.15624e-19 $X=4.99 $Y=0.735
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_1001_n N_A_595_535#_c_1203_n 0.00501365f $X=5.785 $Y=2.72
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_1001_n N_A_595_535#_c_1204_n 0.00274098f $X=5.785 $Y=2.72
+ $X2=0 $Y2=0
cc_759 N_RESET_B_M1010_g N_A_595_535#_c_1192_n 0.0669714f $X=4.99 $Y=0.735 $X2=0
+ $Y2=0
cc_760 N_RESET_B_M1024_g N_A_1475_426#_M1016_g 0.00816694f $X=8.315 $Y=2.65
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_1002_n N_A_1475_426#_M1016_g 0.00730333f $X=7.345 $Y=2.87
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_987_n N_A_1475_426#_M1016_g 0.0184554f $X=7.43 $Y=2.785 $X2=0
+ $Y2=0
cc_763 N_RESET_B_M1003_g N_A_1475_426#_M1019_g 0.0172596f $X=8.41 $Y=0.875 $X2=0
+ $Y2=0
cc_764 N_RESET_B_c_987_n N_A_1475_426#_M1019_g 0.00733387f $X=7.43 $Y=2.785
+ $X2=0 $Y2=0
cc_765 N_RESET_B_c_988_n N_A_1475_426#_M1019_g 0.0144035f $X=8.155 $Y=1.535
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_990_n N_A_1475_426#_M1019_g 0.0155453f $X=8.32 $Y=1.615 $X2=0
+ $Y2=0
cc_767 RESET_B N_A_1475_426#_M1019_g 0.00129968f $X=8.4 $Y=1.665 $X2=0 $Y2=0
cc_768 N_RESET_B_M1024_g N_A_1475_426#_c_1339_n 0.00142613f $X=8.315 $Y=2.65
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_986_n N_A_1475_426#_c_1339_n 5.89898e-19 $X=8.32 $Y=1.955
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_987_n N_A_1475_426#_c_1339_n 0.0248195f $X=7.43 $Y=2.785
+ $X2=0 $Y2=0
cc_771 N_RESET_B_c_988_n N_A_1475_426#_c_1339_n 0.011884f $X=8.155 $Y=1.535
+ $X2=0 $Y2=0
cc_772 RESET_B N_A_1475_426#_c_1339_n 0.0107294f $X=8.4 $Y=1.665 $X2=0 $Y2=0
cc_773 N_RESET_B_M1024_g N_A_1475_426#_c_1340_n 0.00991442f $X=8.315 $Y=2.65
+ $X2=0 $Y2=0
cc_774 N_RESET_B_c_1000_n N_A_1475_426#_c_1340_n 5.77883e-19 $X=8.32 $Y=2.12
+ $X2=0 $Y2=0
cc_775 RESET_B N_A_1475_426#_c_1340_n 0.0154686f $X=8.4 $Y=1.665 $X2=0 $Y2=0
cc_776 N_RESET_B_c_987_n N_A_1475_426#_c_1341_n 0.0136635f $X=7.43 $Y=2.785
+ $X2=0 $Y2=0
cc_777 N_RESET_B_M1024_g N_A_1475_426#_c_1369_n 0.0102199f $X=8.315 $Y=2.65
+ $X2=0 $Y2=0
cc_778 N_RESET_B_M1003_g N_A_1475_426#_c_1335_n 7.84234e-19 $X=8.41 $Y=0.875
+ $X2=0 $Y2=0
cc_779 RESET_B N_A_1475_426#_c_1336_n 0.0089151f $X=8.4 $Y=1.665 $X2=0 $Y2=0
cc_780 N_RESET_B_M1024_g N_A_1475_426#_c_1344_n 0.00269254f $X=8.315 $Y=2.65
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_1000_n N_A_1475_426#_c_1344_n 7.15723e-19 $X=8.32 $Y=2.12
+ $X2=0 $Y2=0
cc_782 RESET_B N_A_1475_426#_c_1344_n 0.0168569f $X=8.4 $Y=1.665 $X2=0 $Y2=0
cc_783 N_RESET_B_M1024_g N_A_1475_426#_c_1345_n 0.00756567f $X=8.315 $Y=2.65
+ $X2=0 $Y2=0
cc_784 N_RESET_B_c_986_n N_A_1475_426#_c_1345_n 0.0105218f $X=8.32 $Y=1.955
+ $X2=0 $Y2=0
cc_785 N_RESET_B_c_987_n N_A_1475_426#_c_1345_n 0.00995407f $X=7.43 $Y=2.785
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_988_n N_A_1475_426#_c_1345_n 0.00473588f $X=8.155 $Y=1.535
+ $X2=0 $Y2=0
cc_787 RESET_B N_A_1475_426#_c_1345_n 6.18247e-19 $X=8.4 $Y=1.665 $X2=0 $Y2=0
cc_788 N_RESET_B_c_1002_n N_A_1255_449#_M1014_d 0.00927087f $X=7.345 $Y=2.87
+ $X2=0 $Y2=0
cc_789 N_RESET_B_M1003_g N_A_1255_449#_c_1422_n 0.0244711f $X=8.41 $Y=0.875
+ $X2=0 $Y2=0
cc_790 N_RESET_B_M1024_g N_A_1255_449#_M1030_g 0.0203265f $X=8.315 $Y=2.65 $X2=0
+ $Y2=0
cc_791 N_RESET_B_c_990_n N_A_1255_449#_c_1426_n 0.0244711f $X=8.32 $Y=1.615
+ $X2=0 $Y2=0
cc_792 N_RESET_B_c_1000_n N_A_1255_449#_c_1435_n 0.0244711f $X=8.32 $Y=2.12
+ $X2=0 $Y2=0
cc_793 N_RESET_B_c_989_n N_A_1255_449#_c_1428_n 0.00527277f $X=7.515 $Y=1.535
+ $X2=0 $Y2=0
cc_794 N_RESET_B_M1003_g N_A_1255_449#_c_1429_n 0.0154293f $X=8.41 $Y=0.875
+ $X2=0 $Y2=0
cc_795 N_RESET_B_c_988_n N_A_1255_449#_c_1429_n 0.0450798f $X=8.155 $Y=1.535
+ $X2=0 $Y2=0
cc_796 N_RESET_B_c_989_n N_A_1255_449#_c_1429_n 0.0137879f $X=7.515 $Y=1.535
+ $X2=0 $Y2=0
cc_797 N_RESET_B_c_990_n N_A_1255_449#_c_1429_n 0.00123753f $X=8.32 $Y=1.615
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_991_n N_A_1255_449#_c_1429_n 0.0311349f $X=8.36 $Y=1.62 $X2=0
+ $Y2=0
cc_799 N_RESET_B_M1003_g N_A_1255_449#_c_1436_n 0.00108447f $X=8.41 $Y=0.875
+ $X2=0 $Y2=0
cc_800 N_RESET_B_c_990_n N_A_1255_449#_c_1436_n 4.16621e-19 $X=8.32 $Y=1.615
+ $X2=0 $Y2=0
cc_801 N_RESET_B_c_991_n N_A_1255_449#_c_1436_n 0.0139495f $X=8.36 $Y=1.62 $X2=0
+ $Y2=0
cc_802 RESET_B N_A_1255_449#_c_1436_n 0.0190958f $X=8.4 $Y=1.665 $X2=0 $Y2=0
cc_803 N_RESET_B_c_986_n N_A_1255_449#_c_1430_n 0.0244711f $X=8.32 $Y=1.955
+ $X2=0 $Y2=0
cc_804 N_RESET_B_c_991_n N_A_1255_449#_c_1430_n 0.00112971f $X=8.36 $Y=1.62
+ $X2=0 $Y2=0
cc_805 RESET_B N_A_1255_449#_c_1430_n 0.00431657f $X=8.4 $Y=1.665 $X2=0 $Y2=0
cc_806 N_RESET_B_c_1002_n N_A_1255_449#_c_1438_n 0.0246499f $X=7.345 $Y=2.87
+ $X2=0 $Y2=0
cc_807 N_RESET_B_c_987_n N_A_1255_449#_c_1431_n 0.00483145f $X=7.43 $Y=2.785
+ $X2=0 $Y2=0
cc_808 N_RESET_B_c_989_n N_A_1255_449#_c_1431_n 9.0989e-19 $X=7.515 $Y=1.535
+ $X2=0 $Y2=0
cc_809 N_RESET_B_c_1001_n N_VPWR_M1027_s 0.0106562f $X=5.785 $Y=2.72 $X2=0 $Y2=0
cc_810 N_RESET_B_M1034_g N_VPWR_c_1642_n 0.00952242f $X=2.04 $Y=2.885 $X2=0
+ $Y2=0
cc_811 N_RESET_B_M1007_g N_VPWR_c_1643_n 0.00315825f $X=4.235 $Y=2.885 $X2=0
+ $Y2=0
cc_812 N_RESET_B_M1024_g N_VPWR_c_1644_n 0.00662613f $X=8.315 $Y=2.65 $X2=0
+ $Y2=0
cc_813 N_RESET_B_c_1002_n N_VPWR_c_1644_n 0.0124986f $X=7.345 $Y=2.87 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_987_n N_VPWR_c_1644_n 0.00943999f $X=7.43 $Y=2.785 $X2=0
+ $Y2=0
cc_815 N_RESET_B_M1024_g N_VPWR_c_1645_n 0.00486495f $X=8.315 $Y=2.65 $X2=0
+ $Y2=0
cc_816 N_RESET_B_M1034_g N_VPWR_c_1654_n 0.00361815f $X=2.04 $Y=2.885 $X2=0
+ $Y2=0
cc_817 N_RESET_B_M1007_g N_VPWR_c_1656_n 0.00435108f $X=4.235 $Y=2.885 $X2=0
+ $Y2=0
cc_818 N_RESET_B_c_1001_n N_VPWR_c_1656_n 0.00492061f $X=5.785 $Y=2.72 $X2=0
+ $Y2=0
cc_819 N_RESET_B_c_1004_n N_VPWR_c_1656_n 0.00434441f $X=4.9 $Y=2.35 $X2=0 $Y2=0
cc_820 N_RESET_B_c_1001_n N_VPWR_c_1657_n 0.0034313f $X=5.785 $Y=2.72 $X2=0
+ $Y2=0
cc_821 N_RESET_B_c_1002_n N_VPWR_c_1657_n 0.0545587f $X=7.345 $Y=2.87 $X2=0
+ $Y2=0
cc_822 N_RESET_B_c_1027_n N_VPWR_c_1657_n 0.00525588f $X=5.87 $Y=2.72 $X2=0
+ $Y2=0
cc_823 N_RESET_B_c_1001_n N_VPWR_c_1663_n 0.0240991f $X=5.785 $Y=2.72 $X2=0
+ $Y2=0
cc_824 N_RESET_B_M1034_g N_VPWR_c_1640_n 0.00573574f $X=2.04 $Y=2.885 $X2=0
+ $Y2=0
cc_825 N_RESET_B_M1007_g N_VPWR_c_1640_n 0.00747288f $X=4.235 $Y=2.885 $X2=0
+ $Y2=0
cc_826 N_RESET_B_c_995_n N_VPWR_c_1640_n 0.00692031f $X=4.735 $Y=2.46 $X2=0
+ $Y2=0
cc_827 N_RESET_B_M1024_g N_VPWR_c_1640_n 0.00514438f $X=8.315 $Y=2.65 $X2=0
+ $Y2=0
cc_828 N_RESET_B_c_1001_n N_VPWR_c_1640_n 0.0135999f $X=5.785 $Y=2.72 $X2=0
+ $Y2=0
cc_829 N_RESET_B_c_1002_n N_VPWR_c_1640_n 0.0535018f $X=7.345 $Y=2.87 $X2=0
+ $Y2=0
cc_830 N_RESET_B_c_1004_n N_VPWR_c_1640_n 0.0108826f $X=4.9 $Y=2.35 $X2=0 $Y2=0
cc_831 N_RESET_B_c_1027_n N_VPWR_c_1640_n 0.00567106f $X=5.87 $Y=2.72 $X2=0
+ $Y2=0
cc_832 N_RESET_B_M1034_g N_A_340_535#_c_1807_n 0.00173473f $X=2.04 $Y=2.885
+ $X2=0 $Y2=0
cc_833 N_RESET_B_M1034_g N_A_340_535#_c_1808_n 0.013175f $X=2.04 $Y=2.885 $X2=0
+ $Y2=0
cc_834 N_RESET_B_M1022_g N_A_340_535#_c_1806_n 3.25009e-19 $X=2.58 $Y=0.805
+ $X2=0 $Y2=0
cc_835 N_RESET_B_c_1002_n A_1380_488# 0.00984044f $X=7.345 $Y=2.87 $X2=-0.19
+ $Y2=-0.245
cc_836 N_RESET_B_M1034_g N_VGND_c_1948_n 0.00558518f $X=2.04 $Y=2.885 $X2=0
+ $Y2=0
cc_837 N_RESET_B_c_979_n N_VGND_c_1948_n 0.0192892f $X=2.505 $Y=0.18 $X2=0 $Y2=0
cc_838 N_RESET_B_M1022_g N_VGND_c_1948_n 0.00518327f $X=2.58 $Y=0.805 $X2=0
+ $Y2=0
cc_839 N_RESET_B_M1003_g N_VGND_c_1949_n 0.00755774f $X=8.41 $Y=0.875 $X2=0
+ $Y2=0
cc_840 N_RESET_B_c_980_n N_VGND_c_1954_n 0.00891616f $X=2.115 $Y=0.18 $X2=0
+ $Y2=0
cc_841 N_RESET_B_c_982_n N_VGND_c_1956_n 0.00732771f $X=4.915 $Y=0.18 $X2=0
+ $Y2=0
cc_842 N_RESET_B_c_979_n N_VGND_c_1957_n 0.0613898f $X=2.505 $Y=0.18 $X2=0 $Y2=0
cc_843 N_RESET_B_M1003_g N_VGND_c_1958_n 0.00394852f $X=8.41 $Y=0.875 $X2=0
+ $Y2=0
cc_844 N_RESET_B_c_979_n N_VGND_c_1967_n 0.00836734f $X=2.505 $Y=0.18 $X2=0
+ $Y2=0
cc_845 N_RESET_B_c_980_n N_VGND_c_1967_n 0.00790479f $X=2.115 $Y=0.18 $X2=0
+ $Y2=0
cc_846 N_RESET_B_c_982_n N_VGND_c_1967_n 0.0606359f $X=4.915 $Y=0.18 $X2=0 $Y2=0
cc_847 N_RESET_B_M1003_g N_VGND_c_1967_n 0.00458517f $X=8.41 $Y=0.875 $X2=0
+ $Y2=0
cc_848 N_RESET_B_c_985_n N_VGND_c_1967_n 0.00888218f $X=2.58 $Y=0.18 $X2=0 $Y2=0
cc_849 N_A_595_535#_c_1209_n N_VPWR_c_1643_n 0.0223735f $X=3.595 $Y=2.935 $X2=0
+ $Y2=0
cc_850 N_A_595_535#_c_1196_n N_VPWR_c_1643_n 0.0147984f $X=4.32 $Y=2.54 $X2=0
+ $Y2=0
cc_851 N_A_595_535#_c_1209_n N_VPWR_c_1655_n 0.0441653f $X=3.595 $Y=2.935 $X2=0
+ $Y2=0
cc_852 N_A_595_535#_c_1196_n N_VPWR_c_1655_n 0.00259904f $X=4.32 $Y=2.54 $X2=0
+ $Y2=0
cc_853 N_A_595_535#_c_1196_n N_VPWR_c_1656_n 0.00239314f $X=4.32 $Y=2.54 $X2=0
+ $Y2=0
cc_854 N_A_595_535#_c_1199_n N_VPWR_c_1656_n 0.014492f $X=4.45 $Y=2.885 $X2=0
+ $Y2=0
cc_855 N_A_595_535#_M1027_g N_VPWR_c_1657_n 0.00391071f $X=5.77 $Y=2.665 $X2=0
+ $Y2=0
cc_856 N_A_595_535#_M1027_g N_VPWR_c_1663_n 0.0086829f $X=5.77 $Y=2.665 $X2=0
+ $Y2=0
cc_857 N_A_595_535#_M1009_d N_VPWR_c_1640_n 0.00262203f $X=2.975 $Y=2.675 $X2=0
+ $Y2=0
cc_858 N_A_595_535#_M1007_d N_VPWR_c_1640_n 0.00220662f $X=4.31 $Y=2.675 $X2=0
+ $Y2=0
cc_859 N_A_595_535#_M1027_g N_VPWR_c_1640_n 0.00684688f $X=5.77 $Y=2.665 $X2=0
+ $Y2=0
cc_860 N_A_595_535#_c_1209_n N_VPWR_c_1640_n 0.0283119f $X=3.595 $Y=2.935 $X2=0
+ $Y2=0
cc_861 N_A_595_535#_c_1196_n N_VPWR_c_1640_n 0.00908072f $X=4.32 $Y=2.54 $X2=0
+ $Y2=0
cc_862 N_A_595_535#_c_1199_n N_VPWR_c_1640_n 0.0100734f $X=4.45 $Y=2.885 $X2=0
+ $Y2=0
cc_863 N_A_595_535#_c_1209_n N_A_340_535#_c_1811_n 0.0287254f $X=3.595 $Y=2.935
+ $X2=0 $Y2=0
cc_864 N_A_595_535#_c_1197_n N_A_340_535#_c_1811_n 0.0151558f $X=3.765 $Y=2.54
+ $X2=0 $Y2=0
cc_865 N_A_595_535#_c_1209_n A_689_535# 0.00460588f $X=3.595 $Y=2.935 $X2=-0.19
+ $Y2=-0.245
cc_866 N_A_595_535#_c_1195_n A_689_535# 0.0013628f $X=3.68 $Y=2.795 $X2=-0.19
+ $Y2=-0.245
cc_867 N_A_595_535#_c_1189_n N_VGND_M1010_d 0.00184417f $X=5.275 $Y=0.96 $X2=0
+ $Y2=0
cc_868 N_A_595_535#_c_1191_n N_VGND_M1010_d 0.00288274f $X=5.44 $Y=0.96 $X2=0
+ $Y2=0
cc_869 N_A_595_535#_c_1188_n N_VGND_c_1956_n 0.0047158f $X=5.65 $Y=1.055 $X2=0
+ $Y2=0
cc_870 N_A_595_535#_c_1188_n N_VGND_c_1961_n 0.0035584f $X=5.65 $Y=1.055 $X2=0
+ $Y2=0
cc_871 N_A_595_535#_c_1188_n N_VGND_c_1967_n 0.00549001f $X=5.65 $Y=1.055 $X2=0
+ $Y2=0
cc_872 N_A_595_535#_c_1189_n A_829_119# 0.00114952f $X=5.275 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_873 N_A_595_535#_c_1189_n A_905_119# 0.00302501f $X=5.275 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_874 N_A_1475_426#_c_1335_n N_A_1255_449#_c_1422_n 0.00510922f $X=9.125
+ $Y=0.79 $X2=0 $Y2=0
cc_875 N_A_1475_426#_c_1336_n N_A_1255_449#_c_1422_n 0.00446533f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_876 N_A_1475_426#_c_1342_n N_A_1255_449#_M1030_g 0.0137807f $X=9.125 $Y=2.385
+ $X2=0 $Y2=0
cc_877 N_A_1475_426#_c_1336_n N_A_1255_449#_M1030_g 0.0105713f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_878 N_A_1475_426#_c_1344_n N_A_1255_449#_M1030_g 0.00194069f $X=8.53 $Y=2.385
+ $X2=0 $Y2=0
cc_879 N_A_1475_426#_c_1336_n N_A_1255_449#_c_1423_n 0.0142983f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_880 N_A_1475_426#_c_1336_n N_A_1255_449#_M1011_g 0.00147278f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_881 N_A_1475_426#_c_1335_n N_A_1255_449#_c_1426_n 0.00668046f $X=9.125
+ $Y=0.79 $X2=0 $Y2=0
cc_882 N_A_1475_426#_c_1342_n N_A_1255_449#_c_1435_n 0.0028218f $X=9.125
+ $Y=2.385 $X2=0 $Y2=0
cc_883 N_A_1475_426#_M1019_g N_A_1255_449#_c_1429_n 0.0169171f $X=7.71 $Y=0.875
+ $X2=0 $Y2=0
cc_884 N_A_1475_426#_c_1335_n N_A_1255_449#_c_1429_n 0.00757266f $X=9.125
+ $Y=0.79 $X2=0 $Y2=0
cc_885 N_A_1475_426#_c_1336_n N_A_1255_449#_c_1429_n 0.0137362f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_886 N_A_1475_426#_c_1342_n N_A_1255_449#_c_1436_n 0.00816017f $X=9.125
+ $Y=2.385 $X2=0 $Y2=0
cc_887 N_A_1475_426#_c_1336_n N_A_1255_449#_c_1436_n 0.0429824f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_888 N_A_1475_426#_c_1336_n N_A_1255_449#_c_1430_n 0.00633309f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_889 N_A_1475_426#_c_1335_n N_A_1891_47#_c_1545_n 0.0230901f $X=9.125 $Y=0.79
+ $X2=0 $Y2=0
cc_890 N_A_1475_426#_c_1336_n N_A_1891_47#_c_1545_n 0.0353452f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_891 N_A_1475_426#_c_1342_n N_A_1891_47#_c_1546_n 0.0144806f $X=9.125 $Y=2.385
+ $X2=0 $Y2=0
cc_892 N_A_1475_426#_c_1336_n N_A_1891_47#_c_1546_n 0.0546285f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_893 N_A_1475_426#_c_1336_n N_A_1891_47#_c_1548_n 0.0152023f $X=9.21 $Y=2.3
+ $X2=0 $Y2=0
cc_894 N_A_1475_426#_c_1340_n N_VPWR_M1016_d 0.00392776f $X=8.365 $Y=2.385 $X2=0
+ $Y2=0
cc_895 N_A_1475_426#_c_1341_n N_VPWR_M1016_d 0.00357315f $X=7.945 $Y=2.385 $X2=0
+ $Y2=0
cc_896 N_A_1475_426#_c_1342_n N_VPWR_M1030_d 0.00324566f $X=9.125 $Y=2.385 $X2=0
+ $Y2=0
cc_897 N_A_1475_426#_M1016_g N_VPWR_c_1644_n 0.00404179f $X=7.45 $Y=2.65 $X2=0
+ $Y2=0
cc_898 N_A_1475_426#_c_1340_n N_VPWR_c_1644_n 0.00785623f $X=8.365 $Y=2.385
+ $X2=0 $Y2=0
cc_899 N_A_1475_426#_c_1341_n N_VPWR_c_1644_n 0.0198034f $X=7.945 $Y=2.385 $X2=0
+ $Y2=0
cc_900 N_A_1475_426#_c_1369_n N_VPWR_c_1644_n 0.00836453f $X=8.53 $Y=2.65 $X2=0
+ $Y2=0
cc_901 N_A_1475_426#_c_1345_n N_VPWR_c_1644_n 0.00115639f $X=7.71 $Y=2.115 $X2=0
+ $Y2=0
cc_902 N_A_1475_426#_c_1369_n N_VPWR_c_1645_n 0.00688941f $X=8.53 $Y=2.65 $X2=0
+ $Y2=0
cc_903 N_A_1475_426#_c_1342_n N_VPWR_c_1646_n 0.0247696f $X=9.125 $Y=2.385 $X2=0
+ $Y2=0
cc_904 N_A_1475_426#_M1016_g N_VPWR_c_1657_n 0.00373981f $X=7.45 $Y=2.65 $X2=0
+ $Y2=0
cc_905 N_A_1475_426#_M1016_g N_VPWR_c_1640_n 0.00514438f $X=7.45 $Y=2.65 $X2=0
+ $Y2=0
cc_906 N_A_1475_426#_c_1340_n N_VPWR_c_1640_n 0.0107762f $X=8.365 $Y=2.385 $X2=0
+ $Y2=0
cc_907 N_A_1475_426#_c_1341_n N_VPWR_c_1640_n 0.00195944f $X=7.945 $Y=2.385
+ $X2=0 $Y2=0
cc_908 N_A_1475_426#_c_1369_n N_VPWR_c_1640_n 0.0106935f $X=8.53 $Y=2.65 $X2=0
+ $Y2=0
cc_909 N_A_1475_426#_c_1342_n N_VPWR_c_1640_n 0.0101904f $X=9.125 $Y=2.385 $X2=0
+ $Y2=0
cc_910 N_A_1475_426#_M1019_g N_VGND_c_1949_n 0.00881468f $X=7.71 $Y=0.875 $X2=0
+ $Y2=0
cc_911 N_A_1475_426#_c_1335_n N_VGND_c_1949_n 0.0080256f $X=9.125 $Y=0.79 $X2=0
+ $Y2=0
cc_912 N_A_1475_426#_c_1335_n N_VGND_c_1958_n 0.0085396f $X=9.125 $Y=0.79 $X2=0
+ $Y2=0
cc_913 N_A_1475_426#_M1019_g N_VGND_c_1961_n 0.00394852f $X=7.71 $Y=0.875 $X2=0
+ $Y2=0
cc_914 N_A_1475_426#_M1019_g N_VGND_c_1967_n 0.00458517f $X=7.71 $Y=0.875 $X2=0
+ $Y2=0
cc_915 N_A_1475_426#_c_1335_n N_VGND_c_1967_n 0.0133035f $X=9.125 $Y=0.79 $X2=0
+ $Y2=0
cc_916 N_A_1255_449#_c_1424_n N_A_1891_47#_M1004_g 0.0205954f $X=9.795 $Y=1.195
+ $X2=0 $Y2=0
cc_917 N_A_1255_449#_M1011_g N_A_1891_47#_M1005_g 0.0205954f $X=9.795 $Y=2.465
+ $X2=0 $Y2=0
cc_918 N_A_1255_449#_c_1422_n N_A_1891_47#_c_1545_n 0.0029119f $X=8.77 $Y=1.195
+ $X2=0 $Y2=0
cc_919 N_A_1255_449#_c_1423_n N_A_1891_47#_c_1545_n 0.0158953f $X=9.72 $Y=1.27
+ $X2=0 $Y2=0
cc_920 N_A_1255_449#_c_1424_n N_A_1891_47#_c_1545_n 0.00583853f $X=9.795
+ $Y=1.195 $X2=0 $Y2=0
cc_921 N_A_1255_449#_M1011_g N_A_1891_47#_c_1545_n 0.00189228f $X=9.795 $Y=2.465
+ $X2=0 $Y2=0
cc_922 N_A_1255_449#_M1030_g N_A_1891_47#_c_1546_n 0.00428866f $X=8.77 $Y=2.65
+ $X2=0 $Y2=0
cc_923 N_A_1255_449#_M1011_g N_A_1891_47#_c_1546_n 0.00985911f $X=9.795 $Y=2.465
+ $X2=0 $Y2=0
cc_924 N_A_1255_449#_M1011_g N_A_1891_47#_c_1547_n 0.0208169f $X=9.795 $Y=2.465
+ $X2=0 $Y2=0
cc_925 N_A_1255_449#_c_1427_n N_A_1891_47#_c_1549_n 0.0205954f $X=9.795 $Y=1.27
+ $X2=0 $Y2=0
cc_926 N_A_1255_449#_M1030_g N_VPWR_c_1645_n 0.00507111f $X=8.77 $Y=2.65 $X2=0
+ $Y2=0
cc_927 N_A_1255_449#_M1030_g N_VPWR_c_1646_n 0.00559613f $X=8.77 $Y=2.65 $X2=0
+ $Y2=0
cc_928 N_A_1255_449#_M1011_g N_VPWR_c_1646_n 0.00224407f $X=9.795 $Y=2.465 $X2=0
+ $Y2=0
cc_929 N_A_1255_449#_M1011_g N_VPWR_c_1647_n 0.00286085f $X=9.795 $Y=2.465 $X2=0
+ $Y2=0
cc_930 N_A_1255_449#_M1011_g N_VPWR_c_1651_n 0.00585385f $X=9.795 $Y=2.465 $X2=0
+ $Y2=0
cc_931 N_A_1255_449#_M1014_d N_VPWR_c_1640_n 0.00295077f $X=6.275 $Y=2.245 $X2=0
+ $Y2=0
cc_932 N_A_1255_449#_M1030_g N_VPWR_c_1640_n 0.00514438f $X=8.77 $Y=2.65 $X2=0
+ $Y2=0
cc_933 N_A_1255_449#_M1011_g N_VPWR_c_1640_n 0.0118474f $X=9.795 $Y=2.465 $X2=0
+ $Y2=0
cc_934 N_A_1255_449#_c_1429_n N_VGND_c_1949_n 0.0271222f $X=8.735 $Y=1.185 $X2=0
+ $Y2=0
cc_935 N_A_1255_449#_c_1424_n N_VGND_c_1950_n 0.00408645f $X=9.795 $Y=1.195
+ $X2=0 $Y2=0
cc_936 N_A_1255_449#_c_1422_n N_VGND_c_1958_n 0.00391917f $X=8.77 $Y=1.195 $X2=0
+ $Y2=0
cc_937 N_A_1255_449#_c_1424_n N_VGND_c_1958_n 0.00585385f $X=9.795 $Y=1.195
+ $X2=0 $Y2=0
cc_938 N_A_1255_449#_c_1422_n N_VGND_c_1967_n 0.00458517f $X=8.77 $Y=1.195 $X2=0
+ $Y2=0
cc_939 N_A_1255_449#_c_1424_n N_VGND_c_1967_n 0.0118474f $X=9.795 $Y=1.195 $X2=0
+ $Y2=0
cc_940 N_A_1891_47#_c_1546_n N_VPWR_c_1646_n 0.0256778f $X=9.58 $Y=1.98 $X2=0
+ $Y2=0
cc_941 N_A_1891_47#_M1005_g N_VPWR_c_1647_n 0.00271318f $X=10.225 $Y=2.465 $X2=0
+ $Y2=0
cc_942 N_A_1891_47#_c_1546_n N_VPWR_c_1647_n 0.00151807f $X=9.58 $Y=1.98 $X2=0
+ $Y2=0
cc_943 N_A_1891_47#_c_1547_n N_VPWR_c_1647_n 0.0176917f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_944 N_A_1891_47#_M1005_g N_VPWR_c_1648_n 7.4139e-19 $X=10.225 $Y=2.465 $X2=0
+ $Y2=0
cc_945 N_A_1891_47#_M1017_g N_VPWR_c_1648_n 0.0144199f $X=10.655 $Y=2.465 $X2=0
+ $Y2=0
cc_946 N_A_1891_47#_M1026_g N_VPWR_c_1648_n 0.0143393f $X=11.085 $Y=2.465 $X2=0
+ $Y2=0
cc_947 N_A_1891_47#_M1037_g N_VPWR_c_1648_n 7.27171e-19 $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_948 N_A_1891_47#_M1026_g N_VPWR_c_1650_n 7.27171e-19 $X=11.085 $Y=2.465 $X2=0
+ $Y2=0
cc_949 N_A_1891_47#_M1037_g N_VPWR_c_1650_n 0.0153838f $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_950 N_A_1891_47#_c_1546_n N_VPWR_c_1651_n 0.0154837f $X=9.58 $Y=1.98 $X2=0
+ $Y2=0
cc_951 N_A_1891_47#_M1005_g N_VPWR_c_1658_n 0.00585385f $X=10.225 $Y=2.465 $X2=0
+ $Y2=0
cc_952 N_A_1891_47#_M1017_g N_VPWR_c_1658_n 0.00486043f $X=10.655 $Y=2.465 $X2=0
+ $Y2=0
cc_953 N_A_1891_47#_M1026_g N_VPWR_c_1659_n 0.00486043f $X=11.085 $Y=2.465 $X2=0
+ $Y2=0
cc_954 N_A_1891_47#_M1037_g N_VPWR_c_1659_n 0.00486043f $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_955 N_A_1891_47#_M1011_s N_VPWR_c_1640_n 0.00288212f $X=9.455 $Y=1.835 $X2=0
+ $Y2=0
cc_956 N_A_1891_47#_M1005_g N_VPWR_c_1640_n 0.0105477f $X=10.225 $Y=2.465 $X2=0
+ $Y2=0
cc_957 N_A_1891_47#_M1017_g N_VPWR_c_1640_n 0.00824727f $X=10.655 $Y=2.465 $X2=0
+ $Y2=0
cc_958 N_A_1891_47#_M1026_g N_VPWR_c_1640_n 0.00824727f $X=11.085 $Y=2.465 $X2=0
+ $Y2=0
cc_959 N_A_1891_47#_M1037_g N_VPWR_c_1640_n 0.00824727f $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_960 N_A_1891_47#_c_1546_n N_VPWR_c_1640_n 0.00944728f $X=9.58 $Y=1.98 $X2=0
+ $Y2=0
cc_961 N_A_1891_47#_M1006_g N_Q_c_1886_n 0.0138529f $X=10.655 $Y=0.655 $X2=0
+ $Y2=0
cc_962 N_A_1891_47#_M1015_g N_Q_c_1886_n 0.0122095f $X=11.085 $Y=0.655 $X2=0
+ $Y2=0
cc_963 N_A_1891_47#_c_1547_n N_Q_c_1886_n 0.0430173f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_964 N_A_1891_47#_c_1549_n N_Q_c_1886_n 0.00246472f $X=11.515 $Y=1.49 $X2=0
+ $Y2=0
cc_965 N_A_1891_47#_M1004_g N_Q_c_1887_n 0.00255478f $X=10.225 $Y=0.655 $X2=0
+ $Y2=0
cc_966 N_A_1891_47#_c_1545_n N_Q_c_1887_n 0.0048f $X=9.58 $Y=0.42 $X2=0 $Y2=0
cc_967 N_A_1891_47#_c_1547_n N_Q_c_1887_n 0.0182231f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_968 N_A_1891_47#_c_1549_n N_Q_c_1887_n 0.00256759f $X=11.515 $Y=1.49 $X2=0
+ $Y2=0
cc_969 N_A_1891_47#_M1017_g N_Q_c_1891_n 0.013053f $X=10.655 $Y=2.465 $X2=0
+ $Y2=0
cc_970 N_A_1891_47#_M1026_g N_Q_c_1891_n 0.013144f $X=11.085 $Y=2.465 $X2=0
+ $Y2=0
cc_971 N_A_1891_47#_c_1547_n N_Q_c_1891_n 0.0469272f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_972 N_A_1891_47#_c_1549_n N_Q_c_1891_n 0.00243542f $X=11.515 $Y=1.49 $X2=0
+ $Y2=0
cc_973 N_A_1891_47#_M1005_g N_Q_c_1892_n 0.00119404f $X=10.225 $Y=2.465 $X2=0
+ $Y2=0
cc_974 N_A_1891_47#_c_1546_n N_Q_c_1892_n 0.00211984f $X=9.58 $Y=1.98 $X2=0
+ $Y2=0
cc_975 N_A_1891_47#_c_1547_n N_Q_c_1892_n 0.0182232f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_976 N_A_1891_47#_c_1549_n N_Q_c_1892_n 0.00253619f $X=11.515 $Y=1.49 $X2=0
+ $Y2=0
cc_977 N_A_1891_47#_M1029_g N_Q_c_1888_n 0.0164167f $X=11.515 $Y=0.655 $X2=0
+ $Y2=0
cc_978 N_A_1891_47#_c_1547_n N_Q_c_1888_n 0.00727995f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_979 N_A_1891_47#_M1037_g N_Q_c_1893_n 0.0154536f $X=11.515 $Y=2.465 $X2=0
+ $Y2=0
cc_980 N_A_1891_47#_c_1547_n N_Q_c_1893_n 0.00727995f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_981 N_A_1891_47#_M1029_g N_Q_c_1889_n 0.0190786f $X=11.515 $Y=0.655 $X2=0
+ $Y2=0
cc_982 N_A_1891_47#_c_1547_n N_Q_c_1889_n 0.013618f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_983 N_A_1891_47#_M1015_g N_Q_c_1890_n 0.00215913f $X=11.085 $Y=0.655 $X2=0
+ $Y2=0
cc_984 N_A_1891_47#_c_1547_n N_Q_c_1890_n 0.0197979f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_985 N_A_1891_47#_c_1549_n N_Q_c_1890_n 0.00256759f $X=11.515 $Y=1.49 $X2=0
+ $Y2=0
cc_986 N_A_1891_47#_c_1547_n N_Q_c_1895_n 0.0153881f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_987 N_A_1891_47#_c_1549_n N_Q_c_1895_n 0.00253619f $X=11.515 $Y=1.49 $X2=0
+ $Y2=0
cc_988 N_A_1891_47#_M1006_g N_Q_c_1923_n 4.39679e-19 $X=10.655 $Y=0.655 $X2=0
+ $Y2=0
cc_989 N_A_1891_47#_M1015_g N_Q_c_1923_n 0.0101821f $X=11.085 $Y=0.655 $X2=0
+ $Y2=0
cc_990 N_A_1891_47#_M1004_g N_VGND_c_1950_n 0.00257443f $X=10.225 $Y=0.655 $X2=0
+ $Y2=0
cc_991 N_A_1891_47#_c_1545_n N_VGND_c_1950_n 0.00151807f $X=9.58 $Y=0.42 $X2=0
+ $Y2=0
cc_992 N_A_1891_47#_c_1547_n N_VGND_c_1950_n 0.0143994f $X=11.335 $Y=1.49 $X2=0
+ $Y2=0
cc_993 N_A_1891_47#_M1004_g N_VGND_c_1951_n 6.41689e-19 $X=10.225 $Y=0.655 $X2=0
+ $Y2=0
cc_994 N_A_1891_47#_M1006_g N_VGND_c_1951_n 0.0105525f $X=10.655 $Y=0.655 $X2=0
+ $Y2=0
cc_995 N_A_1891_47#_M1015_g N_VGND_c_1951_n 0.00153679f $X=11.085 $Y=0.655 $X2=0
+ $Y2=0
cc_996 N_A_1891_47#_M1015_g N_VGND_c_1953_n 7.16758e-19 $X=11.085 $Y=0.655 $X2=0
+ $Y2=0
cc_997 N_A_1891_47#_M1029_g N_VGND_c_1953_n 0.0127834f $X=11.515 $Y=0.655 $X2=0
+ $Y2=0
cc_998 N_A_1891_47#_c_1545_n N_VGND_c_1958_n 0.0154837f $X=9.58 $Y=0.42 $X2=0
+ $Y2=0
cc_999 N_A_1891_47#_M1004_g N_VGND_c_1962_n 0.00585385f $X=10.225 $Y=0.655 $X2=0
+ $Y2=0
cc_1000 N_A_1891_47#_M1006_g N_VGND_c_1962_n 0.00486043f $X=10.655 $Y=0.655
+ $X2=0 $Y2=0
cc_1001 N_A_1891_47#_M1015_g N_VGND_c_1963_n 0.00571722f $X=11.085 $Y=0.655
+ $X2=0 $Y2=0
cc_1002 N_A_1891_47#_M1029_g N_VGND_c_1963_n 0.00486043f $X=11.515 $Y=0.655
+ $X2=0 $Y2=0
cc_1003 N_A_1891_47#_M1035_s N_VGND_c_1967_n 0.00288212f $X=9.455 $Y=0.235 $X2=0
+ $Y2=0
cc_1004 N_A_1891_47#_M1004_g N_VGND_c_1967_n 0.0105477f $X=10.225 $Y=0.655 $X2=0
+ $Y2=0
cc_1005 N_A_1891_47#_M1006_g N_VGND_c_1967_n 0.00824727f $X=10.655 $Y=0.655
+ $X2=0 $Y2=0
cc_1006 N_A_1891_47#_M1015_g N_VGND_c_1967_n 0.0102806f $X=11.085 $Y=0.655 $X2=0
+ $Y2=0
cc_1007 N_A_1891_47#_M1029_g N_VGND_c_1967_n 0.00824727f $X=11.515 $Y=0.655
+ $X2=0 $Y2=0
cc_1008 N_A_1891_47#_c_1545_n N_VGND_c_1967_n 0.00944728f $X=9.58 $Y=0.42 $X2=0
+ $Y2=0
cc_1009 N_VPWR_c_1640_n N_A_340_535#_M1034_s 0.00236684f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_1010 N_VPWR_c_1640_n N_A_340_535#_M1023_d 0.00247422f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_1011 N_VPWR_c_1654_n N_A_340_535#_c_1807_n 0.0152041f $X=2.09 $Y=3.33 $X2=0
+ $Y2=0
cc_1012 N_VPWR_c_1640_n N_A_340_535#_c_1807_n 0.00987105f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_1013 N_VPWR_c_1642_n N_A_340_535#_c_1808_n 0.020497f $X=2.255 $Y=2.915 $X2=0
+ $Y2=0
cc_1014 N_VPWR_c_1654_n N_A_340_535#_c_1808_n 0.00243952f $X=2.09 $Y=3.33 $X2=0
+ $Y2=0
cc_1015 N_VPWR_c_1655_n N_A_340_535#_c_1808_n 0.00243952f $X=3.935 $Y=3.33 $X2=0
+ $Y2=0
cc_1016 N_VPWR_c_1640_n N_A_340_535#_c_1808_n 0.00928579f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_1017 N_VPWR_c_1655_n N_A_340_535#_c_1810_n 0.0118741f $X=3.935 $Y=3.33 $X2=0
+ $Y2=0
cc_1018 N_VPWR_c_1640_n N_A_340_535#_c_1810_n 0.00872326f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_1019 N_VPWR_c_1655_n N_A_340_535#_c_1811_n 0.0024013f $X=3.935 $Y=3.33 $X2=0
+ $Y2=0
cc_1020 N_VPWR_c_1640_n N_A_340_535#_c_1811_n 0.00426746f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_1021 N_VPWR_c_1640_n A_689_535# 0.00168885f $X=11.76 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1022 N_VPWR_c_1640_n N_Q_M1005_s 0.0041489f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_1023 N_VPWR_c_1640_n N_Q_M1026_s 0.00536646f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_1024 N_VPWR_c_1658_n N_Q_c_1927_n 0.0136943f $X=10.705 $Y=3.33 $X2=0 $Y2=0
cc_1025 N_VPWR_c_1640_n N_Q_c_1927_n 0.00866972f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_1026 N_VPWR_M1017_d N_Q_c_1891_n 0.00176461f $X=10.73 $Y=1.835 $X2=0 $Y2=0
cc_1027 N_VPWR_c_1648_n N_Q_c_1891_n 0.0170777f $X=10.87 $Y=2.18 $X2=0 $Y2=0
cc_1028 N_VPWR_c_1647_n N_Q_c_1892_n 0.0016514f $X=10.01 $Y=1.98 $X2=0 $Y2=0
cc_1029 N_VPWR_c_1659_n N_Q_c_1932_n 0.0124525f $X=11.565 $Y=3.33 $X2=0 $Y2=0
cc_1030 N_VPWR_c_1640_n N_Q_c_1932_n 0.00730901f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_1031 N_VPWR_M1037_d N_Q_c_1893_n 0.0066799f $X=11.59 $Y=1.835 $X2=0 $Y2=0
cc_1032 N_VPWR_c_1650_n N_Q_c_1893_n 0.0197619f $X=11.73 $Y=2.18 $X2=0 $Y2=0
cc_1033 N_Q_c_1886_n N_VGND_M1006_s 0.00176461f $X=11.15 $Y=1.15 $X2=0 $Y2=0
cc_1034 N_Q_c_1888_n N_VGND_M1029_s 0.00271681f $X=11.68 $Y=1.15 $X2=0 $Y2=0
cc_1035 N_Q_c_1887_n N_VGND_c_1950_n 0.0016514f $X=10.535 $Y=1.15 $X2=0 $Y2=0
cc_1036 N_Q_c_1886_n N_VGND_c_1951_n 0.0152916f $X=11.15 $Y=1.15 $X2=0 $Y2=0
cc_1037 N_Q_c_1888_n N_VGND_c_1953_n 0.0197619f $X=11.68 $Y=1.15 $X2=0 $Y2=0
cc_1038 N_Q_c_1941_p N_VGND_c_1962_n 0.0136943f $X=10.44 $Y=0.42 $X2=0 $Y2=0
cc_1039 N_Q_c_1923_n N_VGND_c_1963_n 0.0146655f $X=11.3 $Y=0.42 $X2=0 $Y2=0
cc_1040 N_Q_M1004_d N_VGND_c_1967_n 0.0041489f $X=10.3 $Y=0.235 $X2=0 $Y2=0
cc_1041 N_Q_M1015_d N_VGND_c_1967_n 0.00380103f $X=11.16 $Y=0.235 $X2=0 $Y2=0
cc_1042 N_Q_c_1941_p N_VGND_c_1967_n 0.00866972f $X=10.44 $Y=0.42 $X2=0 $Y2=0
cc_1043 N_Q_c_1923_n N_VGND_c_1967_n 0.00933292f $X=11.3 $Y=0.42 $X2=0 $Y2=0
