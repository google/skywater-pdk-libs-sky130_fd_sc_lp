* File: sky130_fd_sc_lp__nor4_0.spice
* Created: Wed Sep  2 10:10:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4_0.pex.spice"
.subckt sky130_fd_sc_lp__nor4_0  VNB VPB A B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1155 PD=0.7 PS=1.39 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.8 A=0.063
+ P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_B_M1007_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.1302
+ AS=0.0588 PD=1.04 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.4 A=0.063
+ P=1.14 MULT=1
MM1004 N_Y_M1004_d N_C_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1302 PD=0.7 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_D_M1001_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1003 A_174_483# N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.1696 PD=0.88 PS=1.81 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1005 A_252_483# N_B_M1005_g A_174_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0768 PD=0.88 PS=0.88 NRD=19.9955 NRS=19.9955 M=1 R=4.26667 SA=75000.6
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1000 A_330_483# N_C_M1000_g A_252_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0768 PD=0.88 PS=0.88 NRD=19.9955 NRS=19.9955 M=1 R=4.26667 SA=75001
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_Y_M1002_d N_D_M1002_g A_330_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.1696
+ AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__nor4_0.pxi.spice"
*
.ends
*
*
