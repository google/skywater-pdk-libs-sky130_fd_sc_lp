* NGSPICE file created from sky130_fd_sc_lp__mux4_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_27_519# VPB phighvt w=420000u l=150000u
+  ad=8.547e+11p pd=8.89e+06u as=2.226e+11p ps=2.74e+06u
M1001 a_1635_149# S1 a_793_117# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=3.423e+11p ps=3.31e+06u
M1002 X a_1635_149# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1003 a_793_117# S0 a_799_501# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.226e+11p ps=2.74e+06u
M1004 a_1245_21# S1 VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=7.35e+11p ps=8.01e+06u
M1005 a_284_81# a_254_55# a_27_519# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1006 a_284_81# a_1245_21# a_1635_149# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1007 a_879_117# a_254_55# a_793_117# VNB nshort w=420000u l=150000u
+  ad=2.226e+11p pd=2.74e+06u as=0p ps=0u
M1008 a_212_81# A0 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 a_284_81# a_254_55# a_212_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1245_21# S1 VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND S0 a_254_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.10925e+11p ps=1.37e+06u
M1012 VGND A3 a_710_117# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.74e+06u
M1013 a_196_519# A0 VPWR VPB phighvt w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=0p ps=0u
M1014 VGND A1 a_33_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.52e+11p ps=2.88e+06u
M1015 a_879_117# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_793_117# S0 a_710_117# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1635_149# S1 a_284_81# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1018 a_33_81# S0 a_284_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A3 a_968_501# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1020 X a_1635_149# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1021 VPWR S0 a_254_55# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1022 a_793_117# a_1245_21# a_1635_149# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_196_519# S0 a_284_81# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_968_501# a_254_55# a_793_117# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_799_501# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

