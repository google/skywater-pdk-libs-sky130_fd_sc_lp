# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__fah_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__fah_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.125000 1.550000 12.590000 1.880000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.759000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.705000 2.290000 8.035000 2.960000 ;
    END
  END B
  PIN CI
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.520000 1.315000 1.850000 ;
    END
  END CI
  PIN COUT
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 0.740000 1.685000 0.910000 ;
        RECT 0.635000 0.910000 0.805000 2.030000 ;
        RECT 0.635000 2.030000 1.145000 2.200000 ;
        RECT 0.975000 2.200000 1.145000 2.895000 ;
        RECT 0.975000 2.895000 2.585000 3.065000 ;
        RECT 1.515000 0.440000 2.090000 0.670000 ;
        RECT 1.515000 0.670000 1.685000 0.740000 ;
        RECT 1.760000 0.280000 2.090000 0.440000 ;
        RECT 2.335000 2.680000 2.585000 2.895000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.440000 0.445000 3.065000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.440000 0.085000 ;
        RECT  0.660000  0.085000  0.990000 0.560000 ;
        RECT  2.270000  0.085000  2.440000 0.670000 ;
        RECT  7.615000  0.085000  7.865000 0.710000 ;
        RECT 11.655000  0.085000 11.905000 0.670000 ;
        RECT 12.645000  0.085000 12.815000 1.020000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.440000 3.415000 ;
        RECT  0.625000 2.380000  0.795000 3.245000 ;
        RECT  2.845000 2.965000  3.175000 3.245000 ;
        RECT  7.105000 2.310000  7.435000 3.245000 ;
        RECT 11.620000 2.860000 11.870000 3.245000 ;
        RECT 12.645000 2.060000 12.815000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  1.170000 1.090000  1.665000 1.340000 ;
      RECT  1.325000 2.075000  1.665000 2.330000 ;
      RECT  1.325000 2.330000  2.935000 2.500000 ;
      RECT  1.325000 2.500000  1.665000 2.715000 ;
      RECT  1.495000 1.340000  1.665000 2.075000 ;
      RECT  1.865000 0.850000  2.790000 1.020000 ;
      RECT  1.865000 1.020000  2.195000 1.980000 ;
      RECT  1.865000 1.980000  3.285000 2.150000 ;
      RECT  2.375000 1.200000  3.140000 1.370000 ;
      RECT  2.375000 1.370000  2.705000 1.580000 ;
      RECT  2.620000 0.265000  4.190000 0.435000 ;
      RECT  2.620000 0.435000  2.790000 0.850000 ;
      RECT  2.765000 2.500000  2.935000 2.615000 ;
      RECT  2.765000 2.615000  3.525000 2.785000 ;
      RECT  2.970000 0.615000  3.840000 0.785000 ;
      RECT  2.970000 0.785000  3.140000 1.200000 ;
      RECT  3.005000 1.550000  3.490000 1.610000 ;
      RECT  3.005000 1.610000  3.635000 1.780000 ;
      RECT  3.115000 2.150000  3.285000 2.265000 ;
      RECT  3.115000 2.265000  4.525000 2.435000 ;
      RECT  3.320000 0.965000  3.490000 1.550000 ;
      RECT  3.355000 2.785000  3.525000 2.895000 ;
      RECT  3.355000 2.895000  6.575000 3.065000 ;
      RECT  3.465000 1.780000  3.635000 1.915000 ;
      RECT  3.465000 1.915000  3.980000 2.085000 ;
      RECT  3.670000 0.785000  3.840000 0.965000 ;
      RECT  3.670000 0.965000  5.160000 1.135000 ;
      RECT  3.815000 1.350000  4.330000 1.680000 ;
      RECT  4.020000 0.435000  4.190000 0.615000 ;
      RECT  4.020000 0.615000  6.215000 0.785000 ;
      RECT  4.160000 1.680000  4.330000 1.810000 ;
      RECT  4.160000 1.810000  4.875000 1.980000 ;
      RECT  4.195000 2.160000  4.525000 2.265000 ;
      RECT  4.195000 2.435000  4.525000 2.715000 ;
      RECT  4.370000 0.265000  7.435000 0.435000 ;
      RECT  4.705000 1.980000  4.875000 2.680000 ;
      RECT  4.705000 2.680000  5.680000 2.895000 ;
      RECT  4.910000 1.135000  5.160000 1.295000 ;
      RECT  4.990000 1.295000  5.160000 1.405000 ;
      RECT  4.990000 1.405000  5.225000 1.575000 ;
      RECT  5.055000 1.575000  5.225000 2.330000 ;
      RECT  5.055000 2.330000  6.225000 2.500000 ;
      RECT  5.340000 0.965000  5.670000 1.055000 ;
      RECT  5.340000 1.055000  6.215000 1.225000 ;
      RECT  5.405000 1.405000  5.865000 2.150000 ;
      RECT  5.885000 0.785000  6.215000 0.875000 ;
      RECT  5.895000 2.500000  6.225000 2.715000 ;
      RECT  6.045000 1.225000  6.215000 1.960000 ;
      RECT  6.045000 1.960000  6.575000 2.130000 ;
      RECT  6.395000 0.615000  6.575000 1.780000 ;
      RECT  6.405000 2.130000  6.575000 2.895000 ;
      RECT  6.755000 0.665000  7.085000 1.780000 ;
      RECT  6.755000 1.960000  7.435000 2.130000 ;
      RECT  6.755000 2.130000  6.925000 3.065000 ;
      RECT  7.265000 0.435000  7.435000 0.890000 ;
      RECT  7.265000 0.890000  8.360000 1.060000 ;
      RECT  7.265000 1.060000  7.435000 1.960000 ;
      RECT  8.045000 0.390000  8.360000 0.890000 ;
      RECT  8.335000 1.240000  8.710000 1.410000 ;
      RECT  8.335000 1.410000  8.505000 2.875000 ;
      RECT  8.335000 2.875000 10.070000 3.045000 ;
      RECT  8.540000 0.265000 11.475000 0.435000 ;
      RECT  8.540000 0.435000  8.710000 1.240000 ;
      RECT  8.685000 1.590000  9.060000 1.760000 ;
      RECT  8.685000 1.760000  9.015000 2.330000 ;
      RECT  8.685000 2.330000 11.090000 2.500000 ;
      RECT  8.685000 2.500000  9.015000 2.695000 ;
      RECT  8.890000 0.615000  9.060000 1.590000 ;
      RECT  9.195000 1.940000  9.920000 2.150000 ;
      RECT  9.240000 0.615000  9.570000 1.760000 ;
      RECT  9.740000 2.680000 11.440000 2.850000 ;
      RECT  9.740000 2.850000 10.070000 2.875000 ;
      RECT  9.750000 1.260000 10.500000 1.430000 ;
      RECT  9.750000 1.430000  9.920000 1.940000 ;
      RECT  9.785000 0.435000 10.115000 1.080000 ;
      RECT 10.250000 1.610000 10.915000 1.780000 ;
      RECT 10.250000 1.780000 10.580000 2.150000 ;
      RECT 10.330000 0.615000 10.660000 1.255000 ;
      RECT 10.330000 1.255000 10.500000 1.260000 ;
      RECT 10.685000 1.550000 10.915000 1.610000 ;
      RECT 10.760000 1.960000 11.265000 2.130000 ;
      RECT 10.760000 2.130000 11.090000 2.330000 ;
      RECT 10.875000 0.615000 11.125000 1.200000 ;
      RECT 10.875000 1.200000 11.265000 1.370000 ;
      RECT 11.095000 1.370000 11.265000 1.960000 ;
      RECT 11.270000 2.510000 12.465000 2.680000 ;
      RECT 11.305000 0.435000 11.475000 0.850000 ;
      RECT 11.305000 0.850000 12.465000 1.020000 ;
      RECT 11.445000 1.200000 13.325000 1.370000 ;
      RECT 11.445000 1.370000 11.775000 1.675000 ;
      RECT 12.135000 0.340000 12.465000 0.850000 ;
      RECT 12.135000 2.060000 12.465000 2.510000 ;
      RECT 12.135000 2.680000 12.465000 3.065000 ;
      RECT 12.995000 0.340000 13.325000 1.200000 ;
      RECT 12.995000 1.370000 13.325000 3.065000 ;
    LAYER mcon ;
      RECT  3.035000 1.580000  3.205000 1.750000 ;
      RECT  5.435000 1.950000  5.605000 2.120000 ;
      RECT  6.395000 1.580000  6.565000 1.750000 ;
      RECT  6.875000 1.580000  7.045000 1.750000 ;
      RECT  9.275000 1.580000  9.445000 1.750000 ;
      RECT  9.275000 1.950000  9.445000 2.120000 ;
      RECT 10.715000 1.580000 10.885000 1.750000 ;
    LAYER met1 ;
      RECT  2.975000 1.550000  3.265000 1.595000 ;
      RECT  2.975000 1.595000  6.625000 1.735000 ;
      RECT  2.975000 1.735000  3.265000 1.780000 ;
      RECT  5.375000 1.920000  5.665000 1.965000 ;
      RECT  5.375000 1.965000  9.505000 2.105000 ;
      RECT  5.375000 2.105000  5.665000 2.150000 ;
      RECT  6.335000 1.550000  6.625000 1.595000 ;
      RECT  6.335000 1.735000  6.625000 1.780000 ;
      RECT  6.815000 1.550000  7.105000 1.595000 ;
      RECT  6.815000 1.595000 10.945000 1.735000 ;
      RECT  6.815000 1.735000  7.105000 1.780000 ;
      RECT  9.215000 1.550000  9.505000 1.595000 ;
      RECT  9.215000 1.735000  9.505000 1.780000 ;
      RECT  9.215000 1.920000  9.505000 1.965000 ;
      RECT  9.215000 2.105000  9.505000 2.150000 ;
      RECT 10.655000 1.550000 10.945000 1.595000 ;
      RECT 10.655000 1.735000 10.945000 1.780000 ;
  END
END sky130_fd_sc_lp__fah_1
