* File: sky130_fd_sc_lp__a311o_lp.spice
* Created: Wed Sep  2 09:25:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311o_lp.pex.spice"
.subckt sky130_fd_sc_lp__a311o_lp  VNB VPB A3 A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1014 A_115_47# N_A_85_21#_M1014_g N_X_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_85_21#_M1007_g A_115_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.08085 AS=0.0441 PD=0.805 PS=0.63 NRD=30 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1004 A_294_47# N_A3_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.08085 PD=0.66 PS=0.805 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.1 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1001 A_372_47# N_A2_M1001_g A_294_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_85_21#_M1002_d N_A1_M1002_g A_372_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.9
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1010 A_536_47# N_B1_M1010_g N_A_85_21#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_B1_M1005_g A_536_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.7 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1012 A_694_47# N_C1_M1012_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1013 N_A_85_21#_M1013_d N_C1_M1013_g A_694_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_85_21#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1003 N_A_257_414#_M1003_d N_A3_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_257_414#_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.1925 AS=0.14 PD=1.385 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1000 N_A_257_414#_M1000_d N_A1_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.1925 PD=1.28 PS=1.385 NRD=0 NRS=20.685 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1011 A_596_414# N_B1_M1011_g N_A_257_414#_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.2625 AS=0.14 PD=1.525 PS=1.28 NRD=40.8578 NRS=0 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1009 N_A_85_21#_M1009_d N_C1_M1009_g A_596_414# VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.2625 PD=2.57 PS=1.525 NRD=0 NRS=40.8578 M=1 R=4 SA=125003
+ SB=125000 A=0.25 P=2.5 MULT=1
DX15_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__a311o_lp.pxi.spice"
*
.ends
*
*
