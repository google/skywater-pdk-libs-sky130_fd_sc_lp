* File: sky130_fd_sc_lp__sdfstp_lp.spice
* Created: Wed Sep  2 10:36:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfstp_lp.pex.spice"
.subckt sky130_fd_sc_lp__sdfstp_lp  VNB VPB SCE D SCD CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1017 A_144_47# N_SCE_M1017_g N_A_27_409#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_SCE_M1004_g A_144_47# VNB NSHORT L=0.15 W=0.42 AD=0.1281
+ AS=0.0441 PD=1.03 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1022 A_368_47# N_A_27_409#_M1022_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1281 PD=0.66 PS=1.03 NRD=18.564 NRS=94.284 M=1 R=2.8 SA=75001.3
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1023 N_A_352_406#_M1023_d N_D_M1023_g A_368_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1044 A_532_47# N_SCE_M1044_g N_A_352_406#_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_SCD_M1024_g A_532_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1041 A_837_108# N_CLK_M1041_g N_A_750_108#_M1041_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_CLK_M1029_g A_837_108# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1031 A_1001_108# N_A_750_108#_M1031_g N_VGND_M1029_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1030 N_A_986_409#_M1030_d N_A_750_108#_M1030_g A_1001_108# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_A_1199_419#_M1020_d N_A_750_108#_M1020_g N_A_352_406#_M1020_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0861 AS=0.1197 PD=0.83 PS=1.41 NRD=18.564 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1045 A_1383_125# N_A_986_409#_M1045_g N_A_1199_419#_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0861 PD=0.63 PS=0.83 NRD=14.28 NRS=18.564 M=1 R=2.8
+ SA=75000.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_A_1425_99#_M1034_g A_1383_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.21575 AS=0.0441 PD=2.04 PS=0.63 NRD=131.052 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1025 A_1736_125# N_A_1199_419#_M1025_g N_A_1425_99#_M1025_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_SET_B_M1014_g A_1736_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=11.424 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 A_1928_125# N_A_1199_419#_M1008_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=28.56 M=1 R=2.8 SA=75001.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1042 N_A_2006_125#_M1042_d N_A_986_409#_M1042_g A_1928_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.135175 AS=0.0504 PD=1.155 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1039 A_2124_66# N_A_750_108#_M1039_g N_A_2006_125#_M1042_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.135175 PD=0.66 PS=1.155 NRD=18.564 NRS=22.848 M=1 R=2.8
+ SA=75000.8 SB=75001 A=0.063 P=1.14 MULT=1
MM1040 A_2202_66# N_A_2172_40#_M1040_g A_2124_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1038 N_VGND_M1038_d N_SET_B_M1038_g A_2202_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_2584_57# N_A_2006_125#_M1005_g N_A_2172_40#_M1005_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_2006_125#_M1007_g A_2584_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 A_2854_57# N_A_2006_125#_M1027_g N_A_2767_57#_M1027_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_2006_125#_M1012_g A_2854_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1032 A_3012_57# N_A_2767_57#_M1032_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1026 N_Q_M1026_d N_A_2767_57#_M1026_g A_3012_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_SCE_M1006_g N_A_27_409#_M1006_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1016 N_A_352_406#_M1016_d N_A_27_409#_M1016_g N_A_245_406#_M1016_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1001 A_458_406# N_D_M1001_g N_A_352_406#_M1016_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.14 PD=1.24 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1018 N_VPWR_M1018_d N_SCE_M1018_g A_458_406# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1000 N_A_245_406#_M1000_d N_SCD_M1000_g N_VPWR_M1018_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_CLK_M1002_g N_A_750_108#_M1002_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1035 N_A_986_409#_M1035_d N_A_750_108#_M1035_g N_VPWR_M1002_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.27 AS=0.14 PD=2.54 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1019 N_A_1199_419#_M1019_d N_A_986_409#_M1019_g N_A_352_406#_M1019_s VPB
+ PHIGHVT L=0.25 W=1 AD=0.305 AS=0.275 PD=1.61 PS=2.55 NRD=65.01 NRS=0 M=1 R=4
+ SA=125000 SB=125007 A=0.25 P=2.5 MULT=1
MM1028 A_1371_419# N_A_750_108#_M1028_g N_A_1199_419#_M1019_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.305 PD=1.28 PS=1.61 NRD=16.7253 NRS=0 M=1 R=4 SA=125001
+ SB=125006 A=0.25 P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A_1425_99#_M1009_g A_1371_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.33515 AS=0.14 PD=1.72 PS=1.28 NRD=16.7253 NRS=16.7253 M=1 R=4 SA=125002
+ SB=125005 A=0.25 P=2.5 MULT=1
MM1036 N_A_1425_99#_M1036_d N_A_1199_419#_M1036_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.33515 PD=1.28 PS=1.72 NRD=0 NRS=58.115 M=1 R=4
+ SA=125002 SB=125004 A=0.25 P=2.5 MULT=1
MM1010 N_VPWR_M1010_d N_SET_B_M1010_g N_A_1425_99#_M1036_d VPB PHIGHVT L=0.25
+ W=1 AD=0.2875 AS=0.14 PD=1.575 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125004
+ A=0.25 P=2.5 MULT=1
MM1043 A_1928_419# N_A_1199_419#_M1043_g N_VPWR_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.2875 PD=1.24 PS=1.575 NRD=12.7853 NRS=58.0953 M=1 R=4 SA=125004
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1011 N_A_2006_125#_M1011_d N_A_750_108#_M1011_g A_1928_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.325 AS=0.12 PD=1.65 PS=1.24 NRD=26.5753 NRS=12.7853 M=1 R=4 SA=125004
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1013 A_2206_419# N_A_986_409#_M1013_g N_A_2006_125#_M1011_d VPB PHIGHVT L=0.25
+ W=1 AD=0.145 AS=0.325 PD=1.29 PS=1.65 NRD=17.7103 NRS=46.2753 M=1 R=4
+ SA=125005 SB=125001 A=0.25 P=2.5 MULT=1
MM1033 N_VPWR_M1033_d N_A_2172_40#_M1033_g A_2206_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.265 AS=0.145 PD=1.53 PS=1.29 NRD=0 NRS=17.7103 M=1 R=4 SA=125006
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1021 N_A_2006_125#_M1021_d N_SET_B_M1021_g N_VPWR_M1033_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.265 PD=2.57 PS=1.53 NRD=0 NRS=49.2303 M=1 R=4 SA=125007
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1015 N_VPWR_M1015_d N_A_2006_125#_M1015_g N_A_2172_40#_M1015_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.455 AS=0.285 PD=2.91 PS=2.57 NRD=33.4703 NRS=0 M=1 R=4
+ SA=125000 SB=125000 A=0.25 P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_A_2006_125#_M1003_g N_A_2767_57#_M1003_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1037 N_Q_M1037_d N_A_2767_57#_M1037_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX46_noxref VNB VPB NWDIODE A=30.3853 P=36.37
c_186 VNB 0 3.13631e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__sdfstp_lp.pxi.spice"
*
.ends
*
*
