* File: sky130_fd_sc_lp__mux2_0.spice
* Created: Wed Sep  2 09:59:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2_0.pex.spice"
.subckt sky130_fd_sc_lp__mux2_0  VNB VPB S A1 A0 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_89_200#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1197 PD=0.78 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1004 A_257_94# N_S_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42 AD=0.08645
+ AS=0.0756 PD=0.935 PS=0.78 NRD=43.092 NRS=0 M=1 R=2.8 SA=75000.7 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_89_200#_M1008_d N_A1_M1008_g A_257_94# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.08645 PD=0.81 PS=0.935 NRD=21.42 NRS=43.092 M=1 R=2.8
+ SA=75000.8 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1003 A_467_125# N_A0_M1003_g N_A_89_200#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=9.996 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_509_99#_M1010_g A_467_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0861 AS=0.0441 PD=0.83 PS=0.63 NRD=18.564 NRS=14.28 M=1 R=2.8 SA=75001.7
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_509_99#_M1007_d N_S_M1007_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.0861 PD=1.38 PS=0.83 NRD=1.428 NRS=18.564 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_89_200#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.134098 AS=0.1696 PD=1.24377 PS=1.81 NRD=16.9223 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1002 A_227_491# N_S_M1002_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0880019 PD=0.63 PS=0.816226 NRD=23.443 NRS=26.9693 M=1 R=2.8 SA=75000.7
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1005 N_A_89_200#_M1005_d N_A0_M1005_g A_227_491# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1137 AS=0.0441 PD=1.01 PS=0.63 NRD=44.5417 NRS=23.443 M=1 R=2.8
+ SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 A_423_515# N_A1_M1006_g N_A_89_200#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.105 AS=0.1137 PD=0.92 PS=1.01 NRD=91.4474 NRS=46.886 M=1 R=2.8 SA=75001.3
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_509_99#_M1011_g A_423_515# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09555 AS=0.105 PD=0.875 PS=0.92 NRD=82.0702 NRS=91.4474 M=1 R=2.8
+ SA=75002 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1000 N_A_509_99#_M1000_d N_S_M1000_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.09555 PD=1.37 PS=0.875 NRD=0 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__mux2_0.pxi.spice"
*
.ends
*
*
