* NGSPICE file created from sky130_fd_sc_lp__dfrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_811_341# a_793_463# VPB phighvt w=420000u l=150000u
+  ad=2.6097e+12p pd=2.302e+07u as=8.82e+10p ps=1.26e+06u
M1001 a_427_191# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.0883e+12p ps=1.851e+07u
M1002 a_784_191# a_196_79# a_637_191# VNB nshort w=420000u l=150000u
+  ad=9.87e+10p pd=1.31e+06u as=2.457e+11p ps=2.01e+06u
M1003 a_1582_128# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 VGND a_1272_128# a_2028_367# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VPWR CLK a_27_79# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1006 a_196_79# a_27_79# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 a_811_341# a_637_191# VGND VNB nshort w=640000u l=150000u
+  ad=2.528e+11p pd=2.07e+06u as=0p ps=0u
M1008 a_308_463# D VPWR VPB phighvt w=420000u l=150000u
+  ad=3.465e+11p pd=4.17e+06u as=0p ps=0u
M1009 VPWR a_1272_128# Q_N VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1010 Q_N a_1272_128# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1011 a_1444_320# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1012 a_637_191# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1013 a_1272_128# a_196_79# a_811_341# VNB nshort w=640000u l=150000u
+  ad=3.662e+11p pd=2.5e+06u as=0p ps=0u
M1014 VPWR a_1272_128# a_2028_367# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1015 a_1424_128# a_27_79# a_1272_128# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1016 VPWR RESET_B a_308_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_1272_128# a_1444_320# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_2028_367# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1019 a_637_191# a_196_79# a_308_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_196_79# a_27_79# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1021 Q a_2028_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1022 VGND a_1272_128# Q_N VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q_N a_1272_128# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1272_128# a_27_79# a_811_341# VPB phighvt w=840000u l=150000u
+  ad=2.688e+11p pd=2.43e+06u as=4.82025e+11p ps=3.03e+06u
M1025 a_811_341# a_637_191# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q a_2028_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_308_463# D a_427_191# VNB nshort w=420000u l=150000u
+  ad=2.268e+11p pd=1.92e+06u as=0p ps=0u
M1028 a_637_191# a_27_79# a_308_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1444_320# a_1272_128# a_1582_128# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1030 VGND a_2028_367# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1402_496# a_196_79# a_1272_128# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1032 VGND RESET_B a_861_191# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1033 VGND CLK a_27_79# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1034 a_861_191# a_811_341# a_784_191# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_793_463# a_27_79# a_637_191# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_1444_320# a_1402_496# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_1444_320# a_1424_128# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

