* File: sky130_fd_sc_lp__a21o_4.pxi.spice
* Created: Wed Sep  2 09:20:07 2020
* 
x_PM_SKY130_FD_SC_LP__A21O_4%A_134_269# N_A_134_269#_M1009_s
+ N_A_134_269#_M1000_s N_A_134_269#_M1005_s N_A_134_269#_M1001_g
+ N_A_134_269#_M1002_g N_A_134_269#_M1004_g N_A_134_269#_M1008_g
+ N_A_134_269#_M1012_g N_A_134_269#_M1010_g N_A_134_269#_M1019_g
+ N_A_134_269#_M1017_g N_A_134_269#_c_99_n N_A_134_269#_c_100_n
+ N_A_134_269#_c_101_n N_A_134_269#_c_125_p N_A_134_269#_c_201_p
+ N_A_134_269#_c_110_p N_A_134_269#_c_218_p N_A_134_269#_c_113_p
+ N_A_134_269#_c_111_p N_A_134_269#_c_102_n N_A_134_269#_c_115_p
+ N_A_134_269#_c_147_p PM_SKY130_FD_SC_LP__A21O_4%A_134_269#
x_PM_SKY130_FD_SC_LP__A21O_4%B1 N_B1_M1009_g N_B1_M1005_g N_B1_c_234_n
+ N_B1_c_235_n N_B1_M1018_g N_B1_M1011_g N_B1_c_237_n B1 B1 N_B1_c_239_n
+ N_B1_c_240_n PM_SKY130_FD_SC_LP__A21O_4%B1
x_PM_SKY130_FD_SC_LP__A21O_4%A2 N_A2_M1014_g N_A2_M1003_g N_A2_M1006_g
+ N_A2_M1016_g N_A2_c_298_n N_A2_c_299_n N_A2_c_300_n N_A2_c_301_n A2 A2 A2
+ PM_SKY130_FD_SC_LP__A21O_4%A2
x_PM_SKY130_FD_SC_LP__A21O_4%A1 N_A1_c_378_n N_A1_M1000_g N_A1_M1007_g
+ N_A1_c_380_n N_A1_M1015_g N_A1_M1013_g A1 A1 N_A1_c_383_n
+ PM_SKY130_FD_SC_LP__A21O_4%A1
x_PM_SKY130_FD_SC_LP__A21O_4%VPWR N_VPWR_M1001_d N_VPWR_M1004_d N_VPWR_M1019_d
+ N_VPWR_M1014_s N_VPWR_M1013_d N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n
+ N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n
+ N_VPWR_c_438_n N_VPWR_c_439_n VPWR N_VPWR_c_440_n N_VPWR_c_441_n
+ N_VPWR_c_442_n N_VPWR_c_429_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n
+ PM_SKY130_FD_SC_LP__A21O_4%VPWR
x_PM_SKY130_FD_SC_LP__A21O_4%X N_X_M1002_d N_X_M1010_d N_X_M1001_s N_X_M1012_s
+ N_X_c_559_n N_X_c_573_p N_X_c_527_n N_X_c_522_n N_X_c_528_n N_X_c_564_n
+ N_X_c_574_p N_X_c_529_n N_X_c_523_n N_X_c_524_n X N_X_c_525_n X
+ PM_SKY130_FD_SC_LP__A21O_4%X
x_PM_SKY130_FD_SC_LP__A21O_4%A_529_367# N_A_529_367#_M1005_d
+ N_A_529_367#_M1011_d N_A_529_367#_M1007_s N_A_529_367#_M1016_d
+ N_A_529_367#_c_579_n N_A_529_367#_c_580_n N_A_529_367#_c_584_n
+ N_A_529_367#_c_581_n N_A_529_367#_c_597_n N_A_529_367#_c_602_n
+ N_A_529_367#_c_582_n N_A_529_367#_c_628_n N_A_529_367#_c_609_n
+ N_A_529_367#_c_631_n PM_SKY130_FD_SC_LP__A21O_4%A_529_367#
x_PM_SKY130_FD_SC_LP__A21O_4%VGND N_VGND_M1002_s N_VGND_M1008_s N_VGND_M1017_s
+ N_VGND_M1018_d N_VGND_M1006_s N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n
+ N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n VGND
+ N_VGND_c_640_n N_VGND_c_641_n N_VGND_c_642_n N_VGND_c_643_n N_VGND_c_644_n
+ N_VGND_c_645_n N_VGND_c_646_n PM_SKY130_FD_SC_LP__A21O_4%VGND
x_PM_SKY130_FD_SC_LP__A21O_4%A_792_49# N_A_792_49#_M1003_d N_A_792_49#_M1015_d
+ N_A_792_49#_c_718_n N_A_792_49#_c_721_n N_A_792_49#_c_716_n
+ PM_SKY130_FD_SC_LP__A21O_4%A_792_49#
cc_1 VNB N_A_134_269#_M1002_g 0.0277571f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.665
cc_2 VNB N_A_134_269#_M1008_g 0.0222385f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=0.665
cc_3 VNB N_A_134_269#_M1010_g 0.0222554f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=0.665
cc_4 VNB N_A_134_269#_M1017_g 0.0262275f $X=-0.19 $Y=-0.245 $X2=2.155 $Y2=0.665
cc_5 VNB N_A_134_269#_c_99_n 0.00177186f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.512
cc_6 VNB N_A_134_269#_c_100_n 0.0835514f $X=-0.19 $Y=-0.245 $X2=2.17 $Y2=1.51
cc_7 VNB N_A_134_269#_c_101_n 0.00299669f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.415
cc_8 VNB N_A_134_269#_c_102_n 0.00309679f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=1.91
cc_9 VNB N_B1_M1005_g 0.00623664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_c_234_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_c_235_n 0.016897f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.675
cc_12 VNB N_B1_M1011_g 0.0134297f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.665
cc_13 VNB N_B1_c_237_n 0.00531178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB B1 0.00639597f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.675
cc_15 VNB N_B1_c_239_n 0.0347676f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.345
cc_16 VNB N_B1_c_240_n 0.0200579f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=0.665
cc_17 VNB N_A2_M1014_g 0.00144794f $X=-0.19 $Y=-0.245 $X2=3.06 $Y2=1.835
cc_18 VNB N_A2_M1003_g 0.0223453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_M1006_g 0.0341123f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.465
cc_20 VNB N_A2_c_298_n 0.0280206f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=2.465
cc_21 VNB N_A2_c_299_n 0.00534272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_c_300_n 0.0160398f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.465
cc_23 VNB N_A2_c_301_n 0.0288725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB A2 3.3633e-19 $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=0.665
cc_25 VNB A2 4.83569e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A1_c_378_n 0.0164424f $X=-0.19 $Y=-0.245 $X2=3.06 $Y2=0.245
cc_27 VNB N_A1_M1007_g 0.00595127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_c_380_n 0.0163115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A1_M1013_g 0.00666377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB A1 9.22189e-19 $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.665
cc_31 VNB N_A1_c_383_n 0.0379491f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=0.665
cc_32 VNB N_VPWR_c_429_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_522_n 0.00568134f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=0.665
cc_34 VNB N_X_c_523_n 5.78398e-19 $X=-0.19 $Y=-0.245 $X2=2.035 $Y2=2.465
cc_35 VNB N_X_c_524_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_525_n 0.0232444f $X=-0.19 $Y=-0.245 $X2=2.17 $Y2=1.512
cc_37 VNB X 0.0216127f $X=-0.19 $Y=-0.245 $X2=2.17 $Y2=1.51
cc_38 VNB N_VGND_c_633_n 0.0289266f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.675
cc_39 VNB N_VGND_c_634_n 4.81113e-19 $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.345
cc_40 VNB N_VGND_c_635_n 6.22396e-19 $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=1.675
cc_41 VNB N_VGND_c_636_n 0.0144144f $X=-0.19 $Y=-0.245 $X2=1.605 $Y2=2.465
cc_42 VNB N_VGND_c_637_n 0.0452016f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=1.345
cc_43 VNB N_VGND_c_638_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_639_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=2.035 $Y2=1.675
cc_45 VNB N_VGND_c_640_n 0.017577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_641_n 0.0343292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_642_n 0.015205f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.04
cc_48 VNB N_VGND_c_643_n 0.034267f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=2.65
cc_49 VNB N_VGND_c_644_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=4.405 $Y2=0.945
cc_50 VNB N_VGND_c_645_n 0.0046535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_646_n 0.307879f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.51
cc_52 VNB N_A_792_49#_c_716_n 0.00709086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_A_134_269#_M1001_g 0.0219892f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=2.465
cc_54 VPB N_A_134_269#_M1004_g 0.0180232f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=2.465
cc_55 VPB N_A_134_269#_M1012_g 0.0180551f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=2.465
cc_56 VPB N_A_134_269#_M1019_g 0.0231454f $X=-0.19 $Y=1.655 $X2=2.035 $Y2=2.465
cc_57 VPB N_A_134_269#_c_100_n 0.0178729f $X=-0.19 $Y=1.655 $X2=2.17 $Y2=1.51
cc_58 VPB N_A_134_269#_c_102_n 0.00144531f $X=-0.19 $Y=1.655 $X2=3.2 $Y2=1.91
cc_59 VPB N_B1_M1005_g 0.0252965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_B1_M1011_g 0.0193884f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.665
cc_61 VPB B1 0.00784116f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=1.675
cc_62 VPB N_A2_M1014_g 0.0196905f $X=-0.19 $Y=1.655 $X2=3.06 $Y2=1.835
cc_63 VPB N_A2_M1016_g 0.0247289f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.665
cc_64 VPB N_A2_c_301_n 0.00666853f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB A2 0.00138467f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=0.665
cc_66 VPB A2 0.00148627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A1_M1007_g 0.0199351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A1_M1013_g 0.0198468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB A1 0.00331821f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.665
cc_70 VPB N_VPWR_c_430_n 0.0392658f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=1.675
cc_71 VPB N_VPWR_c_431_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.295 $Y2=0.665
cc_72 VPB N_VPWR_c_432_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.605 $Y2=2.465
cc_73 VPB N_VPWR_c_433_n 0.0162454f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=0.665
cc_74 VPB N_VPWR_c_434_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=2.155 $Y2=1.345
cc_75 VPB N_VPWR_c_435_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=2.205 $Y2=1.512
cc_76 VPB N_VPWR_c_436_n 0.0137583f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.51
cc_77 VPB N_VPWR_c_437_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_438_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.17 $Y2=1.512
cc_79 VPB N_VPWR_c_439_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.17 $Y2=1.51
cc_80 VPB N_VPWR_c_440_n 0.0366813f $X=-0.19 $Y=1.655 $X2=3.185 $Y2=0.86
cc_81 VPB N_VPWR_c_441_n 0.0133881f $X=-0.19 $Y=1.655 $X2=3.2 $Y2=1.97
cc_82 VPB N_VPWR_c_442_n 0.0194407f $X=-0.19 $Y=1.655 $X2=4.515 $Y2=0.945
cc_83 VPB N_VPWR_c_429_n 0.0709945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_444_n 0.00453137f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=1.51
cc_85 VPB N_VPWR_c_445_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.295 $Y2=1.51
cc_86 VPB N_VPWR_c_446_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.035 $Y2=1.51
cc_87 VPB N_X_c_527_n 0.00305784f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_X_c_528_n 0.00201033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_X_c_529_n 0.0216725f $X=-0.19 $Y=1.655 $X2=2.035 $Y2=2.465
cc_90 VPB X 0.0065525f $X=-0.19 $Y=1.655 $X2=2.17 $Y2=1.51
cc_91 VPB N_A_529_367#_c_579_n 0.0018941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_529_367#_c_580_n 0.00939686f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.665
cc_93 VPB N_A_529_367#_c_581_n 0.00732196f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_529_367#_c_582_n 0.00430689f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 N_A_134_269#_c_100_n N_B1_M1005_g 0.00202262f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_96 N_A_134_269#_c_110_p N_B1_M1005_g 0.00734841f $X=3.2 $Y=2.65 $X2=0 $Y2=0
cc_97 N_A_134_269#_c_111_p N_B1_M1005_g 0.00317783f $X=3.2 $Y=1.97 $X2=0 $Y2=0
cc_98 N_A_134_269#_c_102_n N_B1_c_234_n 0.0102007f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_99 N_A_134_269#_c_113_p N_B1_c_235_n 0.0125122f $X=4.405 $Y=0.945 $X2=0 $Y2=0
cc_100 N_A_134_269#_c_102_n N_B1_c_235_n 0.00448257f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_101 N_A_134_269#_c_115_p N_B1_c_235_n 0.00127672f $X=3.215 $Y=0.95 $X2=0
+ $Y2=0
cc_102 N_A_134_269#_c_110_p N_B1_M1011_g 0.00696765f $X=3.2 $Y=2.65 $X2=0 $Y2=0
cc_103 N_A_134_269#_c_111_p N_B1_M1011_g 0.00166729f $X=3.2 $Y=1.97 $X2=0 $Y2=0
cc_104 N_A_134_269#_c_102_n N_B1_M1011_g 0.0123091f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_105 N_A_134_269#_c_102_n N_B1_c_237_n 0.00244642f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_106 N_A_134_269#_M1019_g B1 0.00238924f $X=2.035 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_134_269#_M1017_g B1 3.96121e-19 $X=2.155 $Y=0.665 $X2=0 $Y2=0
cc_108 N_A_134_269#_c_99_n B1 0.0167299f $X=2.205 $Y=1.512 $X2=0 $Y2=0
cc_109 N_A_134_269#_c_100_n B1 0.0027606f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_110 N_A_134_269#_c_101_n B1 0.0157494f $X=2.29 $Y=1.415 $X2=0 $Y2=0
cc_111 N_A_134_269#_c_125_p B1 0.0276354f $X=3.065 $Y=0.955 $X2=0 $Y2=0
cc_112 N_A_134_269#_c_102_n B1 0.042528f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_113 N_A_134_269#_M1017_g N_B1_c_239_n 0.00306192f $X=2.155 $Y=0.665 $X2=0
+ $Y2=0
cc_114 N_A_134_269#_c_99_n N_B1_c_239_n 3.95876e-19 $X=2.205 $Y=1.512 $X2=0
+ $Y2=0
cc_115 N_A_134_269#_c_100_n N_B1_c_239_n 0.00662571f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_116 N_A_134_269#_c_101_n N_B1_c_239_n 5.28517e-19 $X=2.29 $Y=1.415 $X2=0
+ $Y2=0
cc_117 N_A_134_269#_c_125_p N_B1_c_239_n 0.00146176f $X=3.065 $Y=0.955 $X2=0
+ $Y2=0
cc_118 N_A_134_269#_c_102_n N_B1_c_239_n 0.0050905f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_119 N_A_134_269#_M1017_g N_B1_c_240_n 0.00961873f $X=2.155 $Y=0.665 $X2=0
+ $Y2=0
cc_120 N_A_134_269#_c_101_n N_B1_c_240_n 0.0026365f $X=2.29 $Y=1.415 $X2=0 $Y2=0
cc_121 N_A_134_269#_c_125_p N_B1_c_240_n 0.0182337f $X=3.065 $Y=0.955 $X2=0
+ $Y2=0
cc_122 N_A_134_269#_c_102_n N_B1_c_240_n 0.00335804f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_123 N_A_134_269#_c_102_n N_A2_M1014_g 6.99845e-19 $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_124 N_A_134_269#_c_113_p N_A2_M1003_g 0.0125555f $X=4.405 $Y=0.945 $X2=0
+ $Y2=0
cc_125 N_A_134_269#_c_102_n N_A2_M1003_g 0.00121843f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_126 N_A_134_269#_c_113_p N_A2_c_298_n 0.0036114f $X=4.405 $Y=0.945 $X2=0
+ $Y2=0
cc_127 N_A_134_269#_c_102_n N_A2_c_298_n 3.46374e-19 $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_128 N_A_134_269#_c_113_p N_A2_c_299_n 0.0171012f $X=4.405 $Y=0.945 $X2=0
+ $Y2=0
cc_129 N_A_134_269#_c_102_n N_A2_c_299_n 0.0142261f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_130 N_A_134_269#_c_102_n A2 0.00506182f $X=3.2 $Y=1.91 $X2=0 $Y2=0
cc_131 N_A_134_269#_c_113_p N_A1_c_378_n 0.0107739f $X=4.405 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A_134_269#_c_113_p A1 0.00943072f $X=4.405 $Y=0.945 $X2=0 $Y2=0
cc_133 N_A_134_269#_c_147_p A1 0.0151905f $X=4.53 $Y=0.77 $X2=0 $Y2=0
cc_134 N_A_134_269#_c_147_p N_A1_c_383_n 0.00232209f $X=4.53 $Y=0.77 $X2=0 $Y2=0
cc_135 N_A_134_269#_M1001_g N_VPWR_c_430_n 0.0146751f $X=0.745 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A_134_269#_M1004_g N_VPWR_c_430_n 7.10197e-19 $X=1.175 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A_134_269#_M1001_g N_VPWR_c_431_n 7.10197e-19 $X=0.745 $Y=2.465 $X2=0
+ $Y2=0
cc_138 N_A_134_269#_M1004_g N_VPWR_c_431_n 0.0136126f $X=1.175 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_134_269#_M1012_g N_VPWR_c_431_n 0.0136126f $X=1.605 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_134_269#_M1019_g N_VPWR_c_431_n 7.10197e-19 $X=2.035 $Y=2.465 $X2=0
+ $Y2=0
cc_141 N_A_134_269#_M1012_g N_VPWR_c_432_n 0.00486043f $X=1.605 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_134_269#_M1019_g N_VPWR_c_432_n 0.00486043f $X=2.035 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_134_269#_M1012_g N_VPWR_c_433_n 8.13892e-19 $X=1.605 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_134_269#_M1019_g N_VPWR_c_433_n 0.0222283f $X=2.035 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_134_269#_c_99_n N_VPWR_c_433_n 0.021583f $X=2.205 $Y=1.512 $X2=0
+ $Y2=0
cc_146 N_A_134_269#_c_100_n N_VPWR_c_433_n 0.00605835f $X=2.17 $Y=1.51 $X2=0
+ $Y2=0
cc_147 N_A_134_269#_c_111_p N_VPWR_c_433_n 5.66793e-19 $X=3.2 $Y=1.97 $X2=0
+ $Y2=0
cc_148 N_A_134_269#_M1001_g N_VPWR_c_438_n 0.00486043f $X=0.745 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_134_269#_M1004_g N_VPWR_c_438_n 0.00486043f $X=1.175 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_134_269#_M1005_s N_VPWR_c_429_n 0.00225186f $X=3.06 $Y=1.835 $X2=0
+ $Y2=0
cc_151 N_A_134_269#_M1001_g N_VPWR_c_429_n 0.00824727f $X=0.745 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_134_269#_M1004_g N_VPWR_c_429_n 0.00824727f $X=1.175 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A_134_269#_M1012_g N_VPWR_c_429_n 0.00824727f $X=1.605 $Y=2.465 $X2=0
+ $Y2=0
cc_154 N_A_134_269#_M1019_g N_VPWR_c_429_n 0.00824727f $X=2.035 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_134_269#_M1004_g N_X_c_527_n 0.0139048f $X=1.175 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A_134_269#_M1012_g N_X_c_527_n 0.0138193f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_134_269#_c_99_n N_X_c_527_n 0.0479079f $X=2.205 $Y=1.512 $X2=0 $Y2=0
cc_158 N_A_134_269#_c_100_n N_X_c_527_n 0.00285479f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A_134_269#_M1008_g N_X_c_522_n 0.0141287f $X=1.295 $Y=0.665 $X2=0 $Y2=0
cc_160 N_A_134_269#_M1010_g N_X_c_522_n 0.0137525f $X=1.725 $Y=0.665 $X2=0 $Y2=0
cc_161 N_A_134_269#_M1017_g N_X_c_522_n 0.00131587f $X=2.155 $Y=0.665 $X2=0
+ $Y2=0
cc_162 N_A_134_269#_c_99_n N_X_c_522_n 0.0626799f $X=2.205 $Y=1.512 $X2=0 $Y2=0
cc_163 N_A_134_269#_c_100_n N_X_c_522_n 0.00582235f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A_134_269#_c_101_n N_X_c_522_n 0.0132012f $X=2.29 $Y=1.415 $X2=0 $Y2=0
cc_165 N_A_134_269#_M1019_g N_X_c_528_n 0.00128229f $X=2.035 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_134_269#_c_99_n N_X_c_528_n 0.015469f $X=2.205 $Y=1.512 $X2=0 $Y2=0
cc_167 N_A_134_269#_c_100_n N_X_c_528_n 0.00294396f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_168 N_A_134_269#_M1001_g N_X_c_529_n 0.0152346f $X=0.745 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_134_269#_c_99_n N_X_c_529_n 0.00569942f $X=2.205 $Y=1.512 $X2=0 $Y2=0
cc_170 N_A_134_269#_c_100_n N_X_c_529_n 0.0033896f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_171 N_A_134_269#_M1002_g N_X_c_523_n 0.0129151f $X=0.865 $Y=0.665 $X2=0 $Y2=0
cc_172 N_A_134_269#_c_99_n N_X_c_524_n 0.0154689f $X=2.205 $Y=1.512 $X2=0 $Y2=0
cc_173 N_A_134_269#_c_100_n N_X_c_524_n 0.00296179f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_174 N_A_134_269#_M1002_g N_X_c_525_n 0.00444783f $X=0.865 $Y=0.665 $X2=0
+ $Y2=0
cc_175 N_A_134_269#_M1001_g X 0.00520054f $X=0.745 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_134_269#_M1002_g X 0.0041585f $X=0.865 $Y=0.665 $X2=0 $Y2=0
cc_177 N_A_134_269#_M1004_g X 6.21626e-19 $X=1.175 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_134_269#_M1008_g X 4.66784e-19 $X=1.295 $Y=0.665 $X2=0 $Y2=0
cc_179 N_A_134_269#_c_99_n X 0.0154705f $X=2.205 $Y=1.512 $X2=0 $Y2=0
cc_180 N_A_134_269#_c_100_n X 0.0239422f $X=2.17 $Y=1.51 $X2=0 $Y2=0
cc_181 N_A_134_269#_M1019_g N_A_529_367#_c_580_n 0.00208923f $X=2.035 $Y=2.465
+ $X2=0 $Y2=0
cc_182 N_A_134_269#_M1005_s N_A_529_367#_c_584_n 0.00332344f $X=3.06 $Y=1.835
+ $X2=0 $Y2=0
cc_183 N_A_134_269#_c_110_p N_A_529_367#_c_584_n 0.0159805f $X=3.2 $Y=2.65 $X2=0
+ $Y2=0
cc_184 N_A_134_269#_c_102_n N_A_529_367#_c_581_n 0.018735f $X=3.2 $Y=1.91 $X2=0
+ $Y2=0
cc_185 N_A_134_269#_c_101_n N_VGND_M1017_s 6.98698e-19 $X=2.29 $Y=1.415 $X2=0
+ $Y2=0
cc_186 N_A_134_269#_c_125_p N_VGND_M1017_s 0.0175764f $X=3.065 $Y=0.955 $X2=0
+ $Y2=0
cc_187 N_A_134_269#_c_201_p N_VGND_M1017_s 9.73829e-19 $X=2.375 $Y=0.955 $X2=0
+ $Y2=0
cc_188 N_A_134_269#_c_113_p N_VGND_M1018_d 0.00855116f $X=4.405 $Y=0.945 $X2=0
+ $Y2=0
cc_189 N_A_134_269#_M1002_g N_VGND_c_633_n 0.0126333f $X=0.865 $Y=0.665 $X2=0
+ $Y2=0
cc_190 N_A_134_269#_M1008_g N_VGND_c_633_n 6.15775e-19 $X=1.295 $Y=0.665 $X2=0
+ $Y2=0
cc_191 N_A_134_269#_c_100_n N_VGND_c_633_n 4.14599e-19 $X=2.17 $Y=1.51 $X2=0
+ $Y2=0
cc_192 N_A_134_269#_M1002_g N_VGND_c_634_n 6.15775e-19 $X=0.865 $Y=0.665 $X2=0
+ $Y2=0
cc_193 N_A_134_269#_M1008_g N_VGND_c_634_n 0.0112407f $X=1.295 $Y=0.665 $X2=0
+ $Y2=0
cc_194 N_A_134_269#_M1010_g N_VGND_c_634_n 0.0113159f $X=1.725 $Y=0.665 $X2=0
+ $Y2=0
cc_195 N_A_134_269#_M1017_g N_VGND_c_634_n 6.29009e-19 $X=2.155 $Y=0.665 $X2=0
+ $Y2=0
cc_196 N_A_134_269#_c_113_p N_VGND_c_635_n 0.0176789f $X=4.405 $Y=0.945 $X2=0
+ $Y2=0
cc_197 N_A_134_269#_M1002_g N_VGND_c_638_n 0.00477554f $X=0.865 $Y=0.665 $X2=0
+ $Y2=0
cc_198 N_A_134_269#_M1008_g N_VGND_c_638_n 0.00477554f $X=1.295 $Y=0.665 $X2=0
+ $Y2=0
cc_199 N_A_134_269#_M1010_g N_VGND_c_641_n 0.00477554f $X=1.725 $Y=0.665 $X2=0
+ $Y2=0
cc_200 N_A_134_269#_M1017_g N_VGND_c_641_n 0.00887456f $X=2.155 $Y=0.665 $X2=0
+ $Y2=0
cc_201 N_A_134_269#_c_100_n N_VGND_c_641_n 2.31128e-19 $X=2.17 $Y=1.51 $X2=0
+ $Y2=0
cc_202 N_A_134_269#_c_125_p N_VGND_c_641_n 0.0388529f $X=3.065 $Y=0.955 $X2=0
+ $Y2=0
cc_203 N_A_134_269#_c_201_p N_VGND_c_641_n 0.00793424f $X=2.375 $Y=0.955 $X2=0
+ $Y2=0
cc_204 N_A_134_269#_c_218_p N_VGND_c_642_n 0.0142265f $X=3.2 $Y=0.42 $X2=0 $Y2=0
cc_205 N_A_134_269#_M1009_s N_VGND_c_646_n 0.00263665f $X=3.06 $Y=0.245 $X2=0
+ $Y2=0
cc_206 N_A_134_269#_M1000_s N_VGND_c_646_n 0.00224381f $X=4.39 $Y=0.245 $X2=0
+ $Y2=0
cc_207 N_A_134_269#_M1002_g N_VGND_c_646_n 0.00825815f $X=0.865 $Y=0.665 $X2=0
+ $Y2=0
cc_208 N_A_134_269#_M1008_g N_VGND_c_646_n 0.00825815f $X=1.295 $Y=0.665 $X2=0
+ $Y2=0
cc_209 N_A_134_269#_M1010_g N_VGND_c_646_n 0.00825815f $X=1.725 $Y=0.665 $X2=0
+ $Y2=0
cc_210 N_A_134_269#_M1017_g N_VGND_c_646_n 0.0112971f $X=2.155 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_134_269#_c_218_p N_VGND_c_646_n 0.00925289f $X=3.2 $Y=0.42 $X2=0
+ $Y2=0
cc_212 N_A_134_269#_c_113_p N_VGND_c_646_n 0.00961405f $X=4.405 $Y=0.945 $X2=0
+ $Y2=0
cc_213 N_A_134_269#_c_115_p N_VGND_c_646_n 0.00206327f $X=3.215 $Y=0.95 $X2=0
+ $Y2=0
cc_214 N_A_134_269#_c_113_p N_A_792_49#_M1003_d 0.00632021f $X=4.405 $Y=0.945
+ $X2=-0.19 $Y2=-0.245
cc_215 N_A_134_269#_M1000_s N_A_792_49#_c_718_n 0.00332931f $X=4.39 $Y=0.245
+ $X2=0 $Y2=0
cc_216 N_A_134_269#_c_113_p N_A_792_49#_c_718_n 0.00414135f $X=4.405 $Y=0.945
+ $X2=0 $Y2=0
cc_217 N_A_134_269#_c_147_p N_A_792_49#_c_718_n 0.0122693f $X=4.53 $Y=0.77 $X2=0
+ $Y2=0
cc_218 N_A_134_269#_c_113_p N_A_792_49#_c_721_n 0.0127538f $X=4.405 $Y=0.945
+ $X2=0 $Y2=0
cc_219 N_B1_M1011_g N_A2_M1014_g 0.0201675f $X=3.415 $Y=2.465 $X2=0 $Y2=0
cc_220 N_B1_c_235_n N_A2_M1003_g 0.0312519f $X=3.415 $Y=1.21 $X2=0 $Y2=0
cc_221 N_B1_c_237_n N_A2_c_298_n 0.0200945f $X=3.415 $Y=1.285 $X2=0 $Y2=0
cc_222 N_B1_c_237_n N_A2_c_299_n 0.00116067f $X=3.415 $Y=1.285 $X2=0 $Y2=0
cc_223 N_B1_M1011_g A2 5.80338e-19 $X=3.415 $Y=2.465 $X2=0 $Y2=0
cc_224 N_B1_M1005_g N_VPWR_c_433_n 0.00616008f $X=2.985 $Y=2.465 $X2=0 $Y2=0
cc_225 N_B1_M1011_g N_VPWR_c_434_n 0.00105139f $X=3.415 $Y=2.465 $X2=0 $Y2=0
cc_226 N_B1_M1005_g N_VPWR_c_440_n 0.00357877f $X=2.985 $Y=2.465 $X2=0 $Y2=0
cc_227 N_B1_M1011_g N_VPWR_c_440_n 0.00357877f $X=3.415 $Y=2.465 $X2=0 $Y2=0
cc_228 N_B1_M1005_g N_VPWR_c_429_n 0.00665089f $X=2.985 $Y=2.465 $X2=0 $Y2=0
cc_229 N_B1_M1011_g N_VPWR_c_429_n 0.00537654f $X=3.415 $Y=2.465 $X2=0 $Y2=0
cc_230 B1 N_A_529_367#_c_580_n 0.0229114f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_231 N_B1_c_239_n N_A_529_367#_c_580_n 8.37334e-19 $X=2.872 $Y=1.285 $X2=0
+ $Y2=0
cc_232 N_B1_M1005_g N_A_529_367#_c_584_n 0.0114565f $X=2.985 $Y=2.465 $X2=0
+ $Y2=0
cc_233 N_B1_M1011_g N_A_529_367#_c_584_n 0.0115031f $X=3.415 $Y=2.465 $X2=0
+ $Y2=0
cc_234 N_B1_M1011_g N_A_529_367#_c_581_n 4.86312e-19 $X=3.415 $Y=2.465 $X2=0
+ $Y2=0
cc_235 N_B1_c_235_n N_VGND_c_635_n 0.00922894f $X=3.415 $Y=1.21 $X2=0 $Y2=0
cc_236 N_B1_c_240_n N_VGND_c_635_n 5.60082e-19 $X=2.872 $Y=1.21 $X2=0 $Y2=0
cc_237 N_B1_c_240_n N_VGND_c_641_n 0.00310779f $X=2.872 $Y=1.21 $X2=0 $Y2=0
cc_238 N_B1_c_235_n N_VGND_c_642_n 0.00515898f $X=3.415 $Y=1.21 $X2=0 $Y2=0
cc_239 N_B1_c_240_n N_VGND_c_642_n 0.00575161f $X=2.872 $Y=1.21 $X2=0 $Y2=0
cc_240 N_B1_c_235_n N_VGND_c_646_n 0.00491861f $X=3.415 $Y=1.21 $X2=0 $Y2=0
cc_241 N_B1_c_240_n N_VGND_c_646_n 0.0113107f $X=2.872 $Y=1.21 $X2=0 $Y2=0
cc_242 N_A2_M1003_g N_A1_c_378_n 0.0375621f $X=3.885 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_243 N_A2_M1014_g N_A1_M1007_g 0.0445769f $X=3.845 $Y=2.465 $X2=0 $Y2=0
cc_244 A2 N_A1_M1007_g 0.00506297f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_245 A2 N_A1_M1007_g 0.0116154f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_246 N_A2_M1006_g N_A1_c_380_n 0.0298999f $X=5.175 $Y=0.665 $X2=0 $Y2=0
cc_247 N_A2_M1016_g N_A1_M1013_g 0.0298999f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_248 A2 N_A1_M1013_g 0.0201882f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_249 N_A2_M1003_g A1 5.01353e-19 $X=3.885 $Y=0.665 $X2=0 $Y2=0
cc_250 N_A2_M1006_g A1 6.02537e-19 $X=5.175 $Y=0.665 $X2=0 $Y2=0
cc_251 N_A2_c_298_n A1 3.51547e-19 $X=3.865 $Y=1.46 $X2=0 $Y2=0
cc_252 N_A2_c_299_n A1 0.0255119f $X=4 $Y=1.46 $X2=0 $Y2=0
cc_253 N_A2_c_300_n A1 0.0162403f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_254 A2 A1 0.00909599f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_255 A2 A1 0.0292363f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_256 N_A2_c_298_n N_A1_c_383_n 0.020855f $X=3.865 $Y=1.46 $X2=0 $Y2=0
cc_257 N_A2_c_299_n N_A1_c_383_n 0.00202953f $X=4 $Y=1.46 $X2=0 $Y2=0
cc_258 N_A2_c_300_n N_A1_c_383_n 0.00282183f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_259 N_A2_c_301_n N_A1_c_383_n 0.0298999f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_260 A2 N_A1_c_383_n 4.18706e-19 $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_261 A2 N_VPWR_M1014_s 0.00251378f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_262 A2 N_VPWR_M1014_s 0.00475975f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_263 A2 N_VPWR_M1013_d 0.00605046f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_264 N_A2_M1014_g N_VPWR_c_434_n 0.00977642f $X=3.845 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A2_M1016_g N_VPWR_c_435_n 0.0114867f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A2_M1014_g N_VPWR_c_440_n 0.00564095f $X=3.845 $Y=2.465 $X2=0 $Y2=0
cc_267 N_A2_M1016_g N_VPWR_c_442_n 0.00486043f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A2_M1014_g N_VPWR_c_429_n 0.00525728f $X=3.845 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A2_M1016_g N_VPWR_c_429_n 0.00560393f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_270 A2 N_A_529_367#_M1007_s 0.00354228f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_271 N_A2_M1014_g N_A_529_367#_c_581_n 5.07161e-19 $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_272 N_A2_c_298_n N_A_529_367#_c_581_n 0.00101414f $X=3.865 $Y=1.46 $X2=0
+ $Y2=0
cc_273 N_A2_c_299_n N_A_529_367#_c_581_n 0.00341088f $X=4 $Y=1.46 $X2=0 $Y2=0
cc_274 A2 N_A_529_367#_c_581_n 0.00527944f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_275 N_A2_M1014_g N_A_529_367#_c_597_n 0.0122628f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_276 N_A2_c_298_n N_A_529_367#_c_597_n 2.36954e-19 $X=3.865 $Y=1.46 $X2=0
+ $Y2=0
cc_277 N_A2_c_299_n N_A_529_367#_c_597_n 0.00358007f $X=4 $Y=1.46 $X2=0 $Y2=0
cc_278 A2 N_A_529_367#_c_597_n 0.00848019f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_279 A2 N_A_529_367#_c_597_n 0.0164663f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_280 N_A2_M1016_g N_A_529_367#_c_602_n 0.0115788f $X=5.175 $Y=2.465 $X2=0
+ $Y2=0
cc_281 N_A2_c_300_n N_A_529_367#_c_602_n 0.00343351f $X=5.265 $Y=1.51 $X2=0
+ $Y2=0
cc_282 A2 N_A_529_367#_c_602_n 0.0234241f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_283 N_A2_M1016_g N_A_529_367#_c_582_n 0.0019927f $X=5.175 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_A2_c_300_n N_A_529_367#_c_582_n 0.011227f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_285 N_A2_c_301_n N_A_529_367#_c_582_n 0.00323663f $X=5.265 $Y=1.51 $X2=0
+ $Y2=0
cc_286 A2 N_A_529_367#_c_582_n 0.00527401f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_287 A2 N_A_529_367#_c_609_n 0.0129403f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_288 N_A2_M1003_g N_VGND_c_635_n 0.00935939f $X=3.885 $Y=0.665 $X2=0 $Y2=0
cc_289 N_A2_M1006_g N_VGND_c_637_n 0.00851669f $X=5.175 $Y=0.665 $X2=0 $Y2=0
cc_290 N_A2_c_300_n N_VGND_c_637_n 0.0109469f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_291 N_A2_c_301_n N_VGND_c_637_n 0.00379112f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_292 N_A2_M1003_g N_VGND_c_643_n 0.00554242f $X=3.885 $Y=0.665 $X2=0 $Y2=0
cc_293 N_A2_M1006_g N_VGND_c_643_n 0.00575161f $X=5.175 $Y=0.665 $X2=0 $Y2=0
cc_294 N_A2_M1003_g N_VGND_c_646_n 0.00528667f $X=3.885 $Y=0.665 $X2=0 $Y2=0
cc_295 N_A2_M1006_g N_VGND_c_646_n 0.011582f $X=5.175 $Y=0.665 $X2=0 $Y2=0
cc_296 N_A2_M1006_g N_A_792_49#_c_716_n 7.59749e-19 $X=5.175 $Y=0.665 $X2=0
+ $Y2=0
cc_297 N_A2_c_300_n N_A_792_49#_c_716_n 0.00924462f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_298 N_A1_M1007_g N_VPWR_c_434_n 0.00857011f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A1_M1013_g N_VPWR_c_434_n 5.52668e-19 $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A1_M1007_g N_VPWR_c_435_n 5.81151e-19 $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A1_M1013_g N_VPWR_c_435_n 0.00985142f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A1_M1007_g N_VPWR_c_441_n 0.00564095f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A1_M1013_g N_VPWR_c_441_n 0.00486043f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A1_M1007_g N_VPWR_c_429_n 0.00523194f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A1_M1013_g N_VPWR_c_429_n 0.00458264f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_306 N_A1_M1007_g N_A_529_367#_c_597_n 0.0101892f $X=4.315 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A1_M1013_g N_A_529_367#_c_602_n 0.00980163f $X=4.745 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A1_c_378_n N_VGND_c_635_n 0.00101612f $X=4.315 $Y=1.195 $X2=0 $Y2=0
cc_309 N_A1_c_378_n N_VGND_c_643_n 0.00351226f $X=4.315 $Y=1.195 $X2=0 $Y2=0
cc_310 N_A1_c_380_n N_VGND_c_643_n 0.00351191f $X=4.745 $Y=1.195 $X2=0 $Y2=0
cc_311 N_A1_c_378_n N_VGND_c_646_n 0.0053374f $X=4.315 $Y=1.195 $X2=0 $Y2=0
cc_312 N_A1_c_380_n N_VGND_c_646_n 0.0053283f $X=4.745 $Y=1.195 $X2=0 $Y2=0
cc_313 N_A1_c_378_n N_A_792_49#_c_718_n 0.00944203f $X=4.315 $Y=1.195 $X2=0
+ $Y2=0
cc_314 N_A1_c_380_n N_A_792_49#_c_718_n 0.0107153f $X=4.745 $Y=1.195 $X2=0 $Y2=0
cc_315 N_A1_c_378_n N_A_792_49#_c_716_n 8.82819e-19 $X=4.315 $Y=1.195 $X2=0
+ $Y2=0
cc_316 N_A1_c_380_n N_A_792_49#_c_716_n 0.0120117f $X=4.745 $Y=1.195 $X2=0 $Y2=0
cc_317 N_VPWR_c_429_n N_X_M1001_s 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_318 N_VPWR_c_429_n N_X_M1012_s 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_319 N_VPWR_c_438_n N_X_c_559_n 0.0124525f $X=1.225 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_c_429_n N_X_c_559_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_321 N_VPWR_M1004_d N_X_c_527_n 0.00177483f $X=1.25 $Y=1.835 $X2=0 $Y2=0
cc_322 N_VPWR_c_431_n N_X_c_527_n 0.0172978f $X=1.39 $Y=2.24 $X2=0 $Y2=0
cc_323 N_VPWR_c_433_n N_X_c_528_n 0.007202f $X=2.25 $Y=1.98 $X2=0 $Y2=0
cc_324 N_VPWR_c_432_n N_X_c_564_n 0.0124525f $X=2.085 $Y=3.33 $X2=0 $Y2=0
cc_325 N_VPWR_c_429_n N_X_c_564_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_326 N_VPWR_M1001_d N_X_c_529_n 0.00300749f $X=0.405 $Y=1.835 $X2=0 $Y2=0
cc_327 N_VPWR_c_430_n N_X_c_529_n 0.0243971f $X=0.53 $Y=2.24 $X2=0 $Y2=0
cc_328 N_VPWR_c_429_n N_A_529_367#_M1005_d 0.00215161f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_329 N_VPWR_c_429_n N_A_529_367#_M1011_d 0.00247114f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_429_n N_A_529_367#_M1007_s 0.00269085f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_429_n N_A_529_367#_M1016_d 0.00317907f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_433_n N_A_529_367#_c_579_n 0.0124586f $X=2.25 $Y=1.98 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_440_n N_A_529_367#_c_579_n 0.0179183f $X=3.915 $Y=3.33 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_429_n N_A_529_367#_c_579_n 0.0101082f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_335 N_VPWR_c_433_n N_A_529_367#_c_580_n 0.0660668f $X=2.25 $Y=1.98 $X2=0
+ $Y2=0
cc_336 N_VPWR_c_440_n N_A_529_367#_c_584_n 0.0489954f $X=3.915 $Y=3.33 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_429_n N_A_529_367#_c_584_n 0.0314463f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_338 N_VPWR_M1014_s N_A_529_367#_c_597_n 0.00435712f $X=3.92 $Y=1.835 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_434_n N_A_529_367#_c_597_n 0.0169326f $X=4.08 $Y=2.805 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_429_n N_A_529_367#_c_597_n 0.0103991f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_341 N_VPWR_M1013_d N_A_529_367#_c_602_n 0.00354175f $X=4.82 $Y=1.835 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_435_n N_A_529_367#_c_602_n 0.0167297f $X=4.96 $Y=2.805 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_429_n N_A_529_367#_c_602_n 0.0106723f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_429_n N_A_529_367#_c_628_n 3.66188e-19 $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_441_n N_A_529_367#_c_609_n 0.0131621f $X=4.795 $Y=3.33 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_429_n N_A_529_367#_c_609_n 0.00808656f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_442_n N_A_529_367#_c_631_n 0.0135387f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_429_n N_A_529_367#_c_631_n 0.00769778f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_349 N_X_c_525_n N_VGND_M1002_s 0.00234883f $X=0.48 $Y=1.245 $X2=-0.19
+ $Y2=-0.245
cc_350 N_X_c_522_n N_VGND_M1008_s 0.00176461f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_351 N_X_c_523_n N_VGND_c_633_n 6.51526e-19 $X=0.985 $Y=1.16 $X2=0 $Y2=0
cc_352 N_X_c_525_n N_VGND_c_633_n 0.0236353f $X=0.48 $Y=1.245 $X2=0 $Y2=0
cc_353 N_X_c_522_n N_VGND_c_634_n 0.0170777f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_354 N_X_c_573_p N_VGND_c_638_n 0.0124525f $X=1.08 $Y=0.42 $X2=0 $Y2=0
cc_355 N_X_c_574_p N_VGND_c_641_n 0.0124525f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_356 N_X_M1002_d N_VGND_c_646_n 0.00536646f $X=0.94 $Y=0.245 $X2=0 $Y2=0
cc_357 N_X_M1010_d N_VGND_c_646_n 0.00536646f $X=1.8 $Y=0.245 $X2=0 $Y2=0
cc_358 N_X_c_573_p N_VGND_c_646_n 0.00730901f $X=1.08 $Y=0.42 $X2=0 $Y2=0
cc_359 N_X_c_574_p N_VGND_c_646_n 0.00730901f $X=1.94 $Y=0.42 $X2=0 $Y2=0
cc_360 N_VGND_c_646_n N_A_792_49#_M1003_d 0.00242385f $X=5.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_361 N_VGND_c_646_n N_A_792_49#_M1015_d 0.00254868f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_362 N_VGND_c_643_n N_A_792_49#_c_718_n 0.0317113f $X=5.26 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_646_n N_A_792_49#_c_718_n 0.019825f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_643_n N_A_792_49#_c_721_n 0.0142106f $X=5.26 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_646_n N_A_792_49#_c_721_n 0.00953265f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_637_n N_A_792_49#_c_716_n 0.00155436f $X=5.39 $Y=0.39 $X2=0
+ $Y2=0
cc_367 N_VGND_c_643_n N_A_792_49#_c_716_n 0.0170335f $X=5.26 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_646_n N_A_792_49#_c_716_n 0.0112813f $X=5.52 $Y=0 $X2=0 $Y2=0
