* File: sky130_fd_sc_lp__o221ai_1.pex.spice
* Created: Wed Sep  2 10:19:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221AI_1%C1 3 7 9 13 14
r30 12 14 35.5432 $w=2.78e-07 $l=2.05e-07 $layer=POLY_cond $X=0.29 $Y=1.46
+ $X2=0.495 $Y2=1.46
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.46 $X2=0.29 $Y2=1.46
r32 9 13 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=1.46
r33 5 14 31.2086 $w=2.78e-07 $l=2.49199e-07 $layer=POLY_cond $X=0.675 $Y=1.625
+ $X2=0.495 $Y2=1.46
r34 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.675 $Y=1.625
+ $X2=0.675 $Y2=2.465
r35 1 14 17.1848 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.46
r36 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_1%B1 3 7 9 13 15
c37 13 0 2.89154e-20 $X=1.25 $Y=1.51
r38 12 15 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.25 $Y=1.51
+ $X2=1.445 $Y2=1.51
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.51 $X2=1.25 $Y2=1.51
r40 9 13 5.58215 $w=3.18e-07 $l=1.55e-07 $layer=LI1_cond $X=1.215 $Y=1.665
+ $X2=1.215 $Y2=1.51
r41 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=1.51
r42 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=2.465
r43 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.345
+ $X2=1.445 $Y2=1.51
r44 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.445 $Y=1.345
+ $X2=1.445 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_1%B2 3 7 9 12 13
c38 3 0 2.89154e-20 $X=1.805 $Y=2.465
r39 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.51
+ $X2=1.895 $Y2=1.675
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.51
+ $X2=1.895 $Y2=1.345
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.895
+ $Y=1.51 $X2=1.895 $Y2=1.51
r42 9 13 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.56
+ $X2=1.895 $Y2=1.56
r43 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.985 $Y=0.665
+ $X2=1.985 $Y2=1.345
r44 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.805 $Y=2.465
+ $X2=1.805 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_1%A2 3 7 9 10 11 12 19
c41 7 0 6.2624e-20 $X=2.525 $Y=2.465
r42 23 34 2.50173 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=2.612 $Y=1.675
+ $X2=2.612 $Y2=1.51
r43 20 34 6.18129 $w=3.28e-07 $l=1.77e-07 $layer=LI1_cond $X=2.435 $Y=1.51
+ $X2=2.612 $Y2=1.51
r44 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.51
+ $X2=2.435 $Y2=1.675
r45 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.51
+ $X2=2.435 $Y2=1.345
r46 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=1.51 $X2=2.435 $Y2=1.51
r47 11 12 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.612 $Y=2.405
+ $X2=2.612 $Y2=2.775
r48 10 11 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.612 $Y=2.035
+ $X2=2.612 $Y2=2.405
r49 9 34 0.97783 $w=3.28e-07 $l=2.8e-08 $layer=LI1_cond $X=2.64 $Y=1.51
+ $X2=2.612 $Y2=1.51
r50 9 10 15.1934 $w=2.43e-07 $l=3.23e-07 $layer=LI1_cond $X=2.612 $Y=1.712
+ $X2=2.612 $Y2=2.035
r51 9 23 1.74042 $w=2.43e-07 $l=3.7e-08 $layer=LI1_cond $X=2.612 $Y=1.712
+ $X2=2.612 $Y2=1.675
r52 7 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.525 $Y=2.465
+ $X2=2.525 $Y2=1.675
r53 3 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.415 $Y=0.665
+ $X2=2.415 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_1%A1 3 7 9 14 15
c24 15 0 6.2624e-20 $X=3.07 $Y=1.46
r25 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.46 $X2=3.07 $Y2=1.46
r26 11 14 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.885 $Y=1.46
+ $X2=3.07 $Y2=1.46
r27 9 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.46
r28 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.625
+ $X2=2.885 $Y2=1.46
r29 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.885 $Y=1.625
+ $X2=2.885 $Y2=2.465
r30 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.295
+ $X2=2.885 $Y2=1.46
r31 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.885 $Y=1.295
+ $X2=2.885 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_1%Y 1 2 3 12 14 16 18 20 25 26 27 28 29 36 38
+ 44 58
r59 45 58 7.73671 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=0.755 $Y=2.025
+ $X2=0.885 $Y2=2.025
r60 36 44 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=0.245 $Y=1.005
+ $X2=0.245 $Y2=0.925
r61 29 45 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=0.72 $Y=2.025
+ $X2=0.755 $Y2=2.025
r62 29 54 15.177 $w=1.88e-07 $l=2.6e-07 $layer=LI1_cond $X=0.72 $Y=2.025
+ $X2=0.46 $Y2=2.025
r63 28 45 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=0.755 $Y=1.665
+ $X2=0.755 $Y2=1.93
r64 27 28 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.755 $Y=1.295
+ $X2=0.755 $Y2=1.665
r65 26 36 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=1.09
+ $X2=0.245 $Y2=1.005
r66 26 44 0.132974 $w=2.58e-07 $l=3e-09 $layer=LI1_cond $X=0.245 $Y=0.922
+ $X2=0.245 $Y2=0.925
r67 25 26 16.2672 $w=2.58e-07 $l=3.67e-07 $layer=LI1_cond $X=0.245 $Y=0.555
+ $X2=0.245 $Y2=0.922
r68 25 38 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.245 $Y=0.555
+ $X2=0.245 $Y2=0.42
r69 22 27 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=0.755 $Y=1.175
+ $X2=0.755 $Y2=1.295
r70 18 24 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=2.12
+ $X2=2.155 $Y2=2.035
r71 18 20 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.155 $Y=2.12
+ $X2=2.155 $Y2=2.48
r72 16 24 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=2.035
+ $X2=2.155 $Y2=2.035
r73 16 58 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=1.99 $Y=2.035
+ $X2=0.885 $Y2=2.035
r74 15 26 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.375 $Y=1.09
+ $X2=0.245 $Y2=1.09
r75 14 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.625 $Y=1.09
+ $X2=0.755 $Y2=1.175
r76 14 15 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.625 $Y=1.09
+ $X2=0.375 $Y2=1.09
r77 10 54 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=0.425 $Y=2.025
+ $X2=0.46 $Y2=2.025
r78 10 12 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.425 $Y=2.12
+ $X2=0.425 $Y2=2.48
r79 3 24 600 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=1.88
+ $Y=1.835 $X2=2.155 $Y2=2.035
r80 3 20 300 $w=1.7e-07 $l=7.70325e-07 $layer=licon1_PDIFF $count=2 $X=1.88
+ $Y=1.835 $X2=2.155 $Y2=2.48
r81 2 54 600 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.335
+ $Y=1.835 $X2=0.46 $Y2=2.015
r82 2 12 300 $w=1.7e-07 $l=7.04734e-07 $layer=licon1_PDIFF $count=2 $X=0.335
+ $Y=1.835 $X2=0.46 $Y2=2.48
r83 1 38 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.235 $X2=0.28 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_1%VPWR 1 2 9 11 13 17 19 24 33 37
r42 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 31 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r47 25 33 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.06 $Y2=3.33
r48 25 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 24 36 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.935 $Y=3.33
+ $X2=3.147 $Y2=3.33
r50 24 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 19 33 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=1.06 $Y2=3.33
r54 19 21 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 17 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 17 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 17 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 13 16 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=3.1 $Y=2.005
+ $X2=3.1 $Y2=2.95
r59 11 36 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.1 $Y=3.245
+ $X2=3.147 $Y2=3.33
r60 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.1 $Y=3.245
+ $X2=3.1 $Y2=2.95
r61 7 33 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=3.245 $X2=1.06
+ $Y2=3.33
r62 7 9 15.0849 $w=6.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.06 $Y=3.245
+ $X2=1.06 $Y2=2.4
r63 2 16 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.95
r64 2 13 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.005
r65 1 9 150 $w=1.7e-07 $l=7.68391e-07 $layer=licon1_PDIFF $count=4 $X=0.75
+ $Y=1.835 $X2=1.23 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_1%A_114_47# 1 2 9 14 16
r23 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0.34
+ $X2=0.71 $Y2=0.34
r24 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=0.34
+ $X2=1.715 $Y2=0.34
r25 9 10 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.55 $Y=0.34
+ $X2=0.875 $Y2=0.34
r26 2 16 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=1.52
+ $Y=0.245 $X2=1.715 $Y2=0.37
r27 1 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_1%A_221_49# 1 2 3 12 14 15 18 20 24 26
r45 22 24 24.9696 $w=2.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.13 $Y=1.005
+ $X2=3.13 $Y2=0.42
r46 21 26 7.38875 $w=1.75e-07 $l=1.40478e-07 $layer=LI1_cond $X=2.325 $Y=1.09
+ $X2=2.187 $Y2=1.085
r47 20 22 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.995 $Y=1.09
+ $X2=3.13 $Y2=1.005
r48 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.995 $Y=1.09
+ $X2=2.325 $Y2=1.09
r49 16 26 0.221902 $w=2.75e-07 $l=9e-08 $layer=LI1_cond $X=2.187 $Y=0.995
+ $X2=2.187 $Y2=1.085
r50 16 18 24.0965 $w=2.73e-07 $l=5.75e-07 $layer=LI1_cond $X=2.187 $Y=0.995
+ $X2=2.187 $Y2=0.42
r51 14 26 7.38875 $w=1.75e-07 $l=1.37e-07 $layer=LI1_cond $X=2.05 $Y=1.085
+ $X2=2.187 $Y2=1.085
r52 14 15 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.05 $Y=1.085
+ $X2=1.38 $Y2=1.085
r53 10 15 7.49754 $w=1.8e-07 $l=1.97949e-07 $layer=LI1_cond $X=1.222 $Y=0.995
+ $X2=1.38 $Y2=1.085
r54 10 12 8.59759 $w=3.13e-07 $l=2.35e-07 $layer=LI1_cond $X=1.222 $Y=0.995
+ $X2=1.222 $Y2=0.76
r55 3 24 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.96
+ $Y=0.245 $X2=3.1 $Y2=0.42
r56 2 18 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.06
+ $Y=0.245 $X2=2.2 $Y2=0.42
r57 1 12 182 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_NDIFF $count=1 $X=1.105
+ $Y=0.245 $X2=1.23 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_1%VGND 1 6 8 10 20 21 24
r37 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r39 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.66
+ $Y2=0
r41 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=3.12
+ $Y2=0
r42 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r43 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 12 16 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r45 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.66
+ $Y2=0
r47 10 16 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.16
+ $Y2=0
r48 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r49 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r50 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=0.085 $X2=2.66
+ $Y2=0
r51 4 6 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0.37
r52 1 6 91 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=2 $X=2.49
+ $Y=0.245 $X2=2.66 $Y2=0.37
.ends

