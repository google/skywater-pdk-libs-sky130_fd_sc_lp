* File: sky130_fd_sc_lp__fah_1.pxi.spice
* Created: Wed Sep  2 09:53:43 2020
* 
x_PM_SKY130_FD_SC_LP__FAH_1%CI N_CI_M1008_g N_CI_M1011_g CI N_CI_c_267_n
+ PM_SKY130_FD_SC_LP__FAH_1%CI
x_PM_SKY130_FD_SC_LP__FAH_1%A_84_21# N_A_84_21#_M1023_d N_A_84_21#_M1013_d
+ N_A_84_21#_M1006_g N_A_84_21#_M1018_g N_A_84_21#_c_309_n N_A_84_21#_c_310_n
+ N_A_84_21#_c_311_n N_A_84_21#_c_312_n N_A_84_21#_c_313_n N_A_84_21#_c_314_n
+ N_A_84_21#_c_339_p N_A_84_21#_c_340_p N_A_84_21#_c_324_n N_A_84_21#_c_315_n
+ N_A_84_21#_c_316_n N_A_84_21#_c_317_n N_A_84_21#_c_325_n N_A_84_21#_c_318_n
+ N_A_84_21#_c_319_n N_A_84_21#_c_326_n N_A_84_21#_c_345_p N_A_84_21#_c_389_p
+ N_A_84_21#_c_320_n PM_SKY130_FD_SC_LP__FAH_1%A_84_21#
x_PM_SKY130_FD_SC_LP__FAH_1%A_413_34# N_A_413_34#_M1024_d N_A_413_34#_M1020_d
+ N_A_413_34#_c_464_n N_A_413_34#_M1004_g N_A_413_34#_M1007_g
+ N_A_413_34#_c_466_n N_A_413_34#_c_467_n N_A_413_34#_c_468_n
+ N_A_413_34#_c_469_n N_A_413_34#_c_470_n N_A_413_34#_c_500_n
+ N_A_413_34#_c_471_n N_A_413_34#_c_472_n N_A_413_34#_c_473_n
+ N_A_413_34#_c_474_n N_A_413_34#_c_475_n N_A_413_34#_c_508_p
+ N_A_413_34#_c_535_p N_A_413_34#_c_476_n N_A_413_34#_c_537_p
+ PM_SKY130_FD_SC_LP__FAH_1%A_413_34#
x_PM_SKY130_FD_SC_LP__FAH_1%A_239_135# N_A_239_135#_M1008_d N_A_239_135#_M1002_d
+ N_A_239_135#_M1011_d N_A_239_135#_M1001_d N_A_239_135#_M1027_g
+ N_A_239_135#_c_600_n N_A_239_135#_c_601_n N_A_239_135#_M1012_g
+ N_A_239_135#_c_602_n N_A_239_135#_c_603_n N_A_239_135#_c_610_n
+ N_A_239_135#_c_646_n N_A_239_135#_c_611_n N_A_239_135#_c_604_n
+ N_A_239_135#_c_605_n N_A_239_135#_c_614_n N_A_239_135#_c_615_n
+ N_A_239_135#_c_616_n N_A_239_135#_c_657_n N_A_239_135#_c_617_n
+ N_A_239_135#_c_606_n N_A_239_135#_c_701_n N_A_239_135#_c_703_n
+ N_A_239_135#_c_619_n N_A_239_135#_c_620_n N_A_239_135#_c_607_n
+ N_A_239_135#_c_664_n N_A_239_135#_c_622_n N_A_239_135#_c_623_n
+ N_A_239_135#_c_669_n N_A_239_135#_c_624_n PM_SKY130_FD_SC_LP__FAH_1%A_239_135#
x_PM_SKY130_FD_SC_LP__FAH_1%A_814_384# N_A_814_384#_M1014_d N_A_814_384#_M1003_d
+ N_A_814_384#_c_835_n N_A_814_384#_M1013_g N_A_814_384#_c_836_n
+ N_A_814_384#_c_837_n N_A_814_384#_c_822_n N_A_814_384#_c_823_n
+ N_A_814_384#_c_824_n N_A_814_384#_M1024_g N_A_814_384#_c_826_n
+ N_A_814_384#_c_827_n N_A_814_384#_M1023_g N_A_814_384#_M1020_g
+ N_A_814_384#_c_829_n N_A_814_384#_c_830_n N_A_814_384#_c_831_n
+ N_A_814_384#_c_832_n N_A_814_384#_c_950_p N_A_814_384#_c_928_p
+ N_A_814_384#_c_841_n N_A_814_384#_c_862_n N_A_814_384#_c_938_p
+ N_A_814_384#_c_833_n N_A_814_384#_c_834_n PM_SKY130_FD_SC_LP__FAH_1%A_814_384#
x_PM_SKY130_FD_SC_LP__FAH_1%A_1022_362# N_A_1022_362#_M1005_d
+ N_A_1022_362#_M1029_d N_A_1022_362#_M1001_g N_A_1022_362#_c_1022_n
+ N_A_1022_362#_M1002_g N_A_1022_362#_c_1024_n N_A_1022_362#_c_1025_n
+ N_A_1022_362#_M1017_g N_A_1022_362#_M1015_g N_A_1022_362#_c_1009_n
+ N_A_1022_362#_c_1010_n N_A_1022_362#_c_1011_n N_A_1022_362#_c_1012_n
+ N_A_1022_362#_c_1029_n N_A_1022_362#_c_1013_n N_A_1022_362#_c_1014_n
+ N_A_1022_362#_c_1015_n N_A_1022_362#_c_1016_n N_A_1022_362#_c_1017_n
+ N_A_1022_362#_c_1018_n N_A_1022_362#_c_1019_n N_A_1022_362#_c_1020_n
+ PM_SKY130_FD_SC_LP__FAH_1%A_1022_362#
x_PM_SKY130_FD_SC_LP__FAH_1%A_878_41# N_A_878_41#_M1024_s N_A_878_41#_M1028_s
+ N_A_878_41#_M1015_d N_A_878_41#_c_1205_n N_A_878_41#_c_1206_n
+ N_A_878_41#_M1003_g N_A_878_41#_M1005_g N_A_878_41#_c_1209_n
+ N_A_878_41#_M1029_g N_A_878_41#_M1014_g N_A_878_41#_c_1212_n
+ N_A_878_41#_c_1213_n N_A_878_41#_c_1214_n N_A_878_41#_c_1215_n
+ N_A_878_41#_c_1227_n N_A_878_41#_c_1228_n N_A_878_41#_c_1221_n
+ N_A_878_41#_c_1344_p N_A_878_41#_c_1271_n N_A_878_41#_c_1216_n
+ N_A_878_41#_c_1217_n N_A_878_41#_c_1288_p N_A_878_41#_c_1218_n
+ N_A_878_41#_c_1279_n PM_SKY130_FD_SC_LP__FAH_1%A_878_41#
x_PM_SKY130_FD_SC_LP__FAH_1%B N_B_c_1363_n N_B_M1022_g N_B_c_1356_n N_B_c_1357_n
+ N_B_M1028_g N_B_c_1366_n N_B_M1021_g N_B_M1025_g N_B_c_1368_n N_B_M1009_g
+ N_B_M1031_g N_B_c_1361_n N_B_c_1371_n N_B_c_1372_n N_B_c_1362_n N_B_c_1374_n B
+ B N_B_c_1376_n PM_SKY130_FD_SC_LP__FAH_1%B
x_PM_SKY130_FD_SC_LP__FAH_1%A_2229_269# N_A_2229_269#_M1010_d
+ N_A_2229_269#_M1016_d N_A_2229_269#_M1000_g N_A_2229_269#_c_1483_n
+ N_A_2229_269#_M1019_g N_A_2229_269#_c_1484_n N_A_2229_269#_c_1485_n
+ N_A_2229_269#_c_1486_n N_A_2229_269#_c_1487_n N_A_2229_269#_c_1488_n
+ N_A_2229_269#_c_1489_n N_A_2229_269#_c_1490_n
+ PM_SKY130_FD_SC_LP__FAH_1%A_2229_269#
x_PM_SKY130_FD_SC_LP__FAH_1%A N_A_M1026_g N_A_M1030_g N_A_c_1553_n N_A_M1010_g
+ N_A_M1016_g N_A_c_1555_n A N_A_c_1556_n N_A_c_1557_n
+ PM_SKY130_FD_SC_LP__FAH_1%A
x_PM_SKY130_FD_SC_LP__FAH_1%SUM N_SUM_M1006_s N_SUM_M1018_s SUM SUM SUM SUM SUM
+ SUM SUM PM_SKY130_FD_SC_LP__FAH_1%SUM
x_PM_SKY130_FD_SC_LP__FAH_1%VPWR N_VPWR_M1018_d N_VPWR_M1007_d N_VPWR_M1022_d
+ N_VPWR_M1000_d N_VPWR_M1030_d N_VPWR_c_1621_n N_VPWR_c_1622_n N_VPWR_c_1623_n
+ N_VPWR_c_1624_n N_VPWR_c_1625_n N_VPWR_c_1626_n N_VPWR_c_1627_n VPWR
+ N_VPWR_c_1628_n N_VPWR_c_1629_n N_VPWR_c_1630_n N_VPWR_c_1631_n
+ N_VPWR_c_1620_n N_VPWR_c_1633_n N_VPWR_c_1634_n N_VPWR_c_1635_n
+ N_VPWR_c_1636_n PM_SKY130_FD_SC_LP__FAH_1%VPWR
x_PM_SKY130_FD_SC_LP__FAH_1%COUT N_COUT_M1004_s N_COUT_M1007_s N_COUT_c_1751_n
+ N_COUT_c_1752_n N_COUT_c_1777_n N_COUT_c_1765_n N_COUT_c_1755_n
+ N_COUT_c_1767_n N_COUT_c_1756_n N_COUT_c_1757_n COUT
+ PM_SKY130_FD_SC_LP__FAH_1%COUT
x_PM_SKY130_FD_SC_LP__FAH_1%A_630_100# N_A_630_100#_M1027_d N_A_630_100#_M1017_d
+ N_A_630_100#_M1012_d N_A_630_100#_c_1828_n N_A_630_100#_c_1834_n
+ N_A_630_100#_c_1835_n N_A_630_100#_c_1829_n N_A_630_100#_c_1830_n
+ N_A_630_100#_c_1831_n N_A_630_100#_c_1832_n N_A_630_100#_c_1833_n
+ PM_SKY130_FD_SC_LP__FAH_1%A_630_100#
x_PM_SKY130_FD_SC_LP__FAH_1%A_1741_367# N_A_1741_367#_M1005_s
+ N_A_1741_367#_M1009_d N_A_1741_367#_M1003_s N_A_1741_367#_M1031_d
+ N_A_1741_367#_c_1926_n N_A_1741_367#_c_1922_n N_A_1741_367#_c_1934_n
+ N_A_1741_367#_c_1965_n N_A_1741_367#_c_1938_n N_A_1741_367#_c_1923_n
+ N_A_1741_367#_c_1924_n N_A_1741_367#_c_1929_n N_A_1741_367#_c_1956_n
+ N_A_1741_367#_c_1925_n PM_SKY130_FD_SC_LP__FAH_1%A_1741_367#
x_PM_SKY130_FD_SC_LP__FAH_1%A_1930_367# N_A_1930_367#_M1025_d
+ N_A_1930_367#_M1026_s N_A_1930_367#_M1021_d N_A_1930_367#_M1030_s
+ N_A_1930_367#_c_2000_n N_A_1930_367#_c_2011_n N_A_1930_367#_c_2012_n
+ N_A_1930_367#_c_2001_n N_A_1930_367#_c_2002_n N_A_1930_367#_c_2003_n
+ N_A_1930_367#_c_2004_n N_A_1930_367#_c_2013_n N_A_1930_367#_c_2005_n
+ N_A_1930_367#_c_2066_n N_A_1930_367#_c_2014_n N_A_1930_367#_c_2006_n
+ N_A_1930_367#_c_2079_n N_A_1930_367#_c_2007_n N_A_1930_367#_c_2015_n
+ N_A_1930_367#_c_2008_n N_A_1930_367#_c_2016_n N_A_1930_367#_c_2009_n
+ N_A_1930_367#_c_2071_n N_A_1930_367#_c_2017_n
+ PM_SKY130_FD_SC_LP__FAH_1%A_1930_367#
x_PM_SKY130_FD_SC_LP__FAH_1%VGND N_VGND_M1006_d N_VGND_M1004_d N_VGND_M1028_d
+ N_VGND_M1019_d N_VGND_M1026_d N_VGND_c_2147_n N_VGND_c_2148_n N_VGND_c_2149_n
+ N_VGND_c_2150_n N_VGND_c_2151_n N_VGND_c_2152_n N_VGND_c_2153_n
+ N_VGND_c_2154_n N_VGND_c_2155_n N_VGND_c_2156_n VGND N_VGND_c_2157_n
+ N_VGND_c_2158_n N_VGND_c_2159_n N_VGND_c_2160_n N_VGND_c_2161_n
+ N_VGND_c_2162_n PM_SKY130_FD_SC_LP__FAH_1%VGND
cc_1 VNB N_CI_M1008_g 0.024487f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.995
cc_2 VNB CI 0.00185942f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_3 VNB N_CI_c_267_n 0.0143665f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.685
cc_4 VNB N_A_84_21#_M1006_g 0.0411252f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_5 VNB N_A_84_21#_c_309_n 0.0797622f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.685
cc_6 VNB N_A_84_21#_c_310_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.52
cc_7 VNB N_A_84_21#_c_311_n 0.0552117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_84_21#_c_312_n 0.016609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_84_21#_c_313_n 0.0171892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_84_21#_c_314_n 0.00450873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_84_21#_c_315_n 0.00147423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_84_21#_c_316_n 0.0325466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_84_21#_c_317_n 0.00353434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_84_21#_c_318_n 0.00970198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_84_21#_c_319_n 0.00406933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_84_21#_c_320_n 0.0109275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_413_34#_c_464_n 0.0204297f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=2.595
cc_18 VNB N_A_413_34#_M1007_g 0.00528893f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.685
cc_19 VNB N_A_413_34#_c_466_n 0.0111821f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.52
cc_20 VNB N_A_413_34#_c_467_n 0.0525128f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.85
cc_21 VNB N_A_413_34#_c_468_n 0.011091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_413_34#_c_469_n 0.00199251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_413_34#_c_470_n 0.00747962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_413_34#_c_471_n 0.00895258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_413_34#_c_472_n 0.0138862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_413_34#_c_473_n 0.00322861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_413_34#_c_474_n 0.00637085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_413_34#_c_475_n 0.00101641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_413_34#_c_476_n 0.00699069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_239_135#_M1027_g 0.027028f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.85
cc_31 VNB N_A_239_135#_c_600_n 0.0177564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_239_135#_c_601_n 0.00882722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_239_135#_c_602_n 0.0130156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_239_135#_c_603_n 0.00789537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_239_135#_c_604_n 0.006014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_239_135#_c_605_n 0.0380908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_239_135#_c_606_n 0.00318286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_239_135#_c_607_n 0.00516931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_814_384#_c_822_n 0.00694278f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.685
cc_40 VNB N_A_814_384#_c_823_n 0.0258635f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.52
cc_41 VNB N_A_814_384#_c_824_n 0.00919885f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.85
cc_42 VNB N_A_814_384#_M1024_g 0.0333609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_814_384#_c_826_n 0.0588869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_814_384#_c_827_n 0.0130185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_814_384#_M1023_g 0.0302196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_814_384#_c_829_n 0.00460379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_814_384#_c_830_n 0.00568446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_814_384#_c_831_n 0.0020247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_814_384#_c_832_n 0.00405378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_814_384#_c_833_n 0.0215463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_814_384#_c_834_n 0.00429545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1022_362#_M1002_g 0.0287524f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.685
cc_53 VNB N_A_1022_362#_c_1009_n 0.0294391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1022_362#_c_1010_n 0.0390282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1022_362#_c_1011_n 0.0172805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1022_362#_c_1012_n 0.00331769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1022_362#_c_1013_n 0.00710536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1022_362#_c_1014_n 9.26429e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1022_362#_c_1015_n 0.00605749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1022_362#_c_1016_n 3.03424e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1022_362#_c_1017_n 0.00463712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1022_362#_c_1018_n 0.0512078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1022_362#_c_1019_n 0.00676478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1022_362#_c_1020_n 0.00246025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_878_41#_c_1205_n 0.051482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_878_41#_c_1206_n 0.0192253f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.685
cc_67 VNB N_A_878_41#_M1003_g 0.00752413f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.52
cc_68 VNB N_A_878_41#_M1005_g 0.0310193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_878_41#_c_1209_n 0.0749731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_878_41#_M1029_g 0.00919397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_878_41#_M1014_g 0.0293345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_878_41#_c_1212_n 0.0121702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_878_41#_c_1213_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_878_41#_c_1214_n 0.0134918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_878_41#_c_1215_n 0.0505178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_878_41#_c_1216_n 0.00922307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_878_41#_c_1217_n 0.0113557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_878_41#_c_1218_n 0.0751487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_B_c_1356_n 0.0164768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_B_c_1357_n 0.00592898f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.85
cc_81 VNB N_B_M1028_g 0.0510365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_B_M1025_g 0.0271058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_B_M1009_g 0.0346228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_B_c_1361_n 0.0129944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_B_c_1362_n 0.00562388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2229_269#_c_1483_n 0.0193918f $X=-0.19 $Y=-0.245 $X2=1.15
+ $Y2=1.685
cc_87 VNB N_A_2229_269#_c_1484_n 0.0121115f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.85
cc_88 VNB N_A_2229_269#_c_1485_n 0.0343003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2229_269#_c_1486_n 0.0360316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2229_269#_c_1487_n 0.0118868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2229_269#_c_1488_n 9.33493e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2229_269#_c_1489_n 0.0362402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2229_269#_c_1490_n 0.00770964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_M1026_g 0.0499471f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.995
cc_95 VNB N_A_c_1553_n 0.00534052f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_96 VNB N_A_M1010_g 0.0481231f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.685
cc_97 VNB N_A_c_1555_n 0.00466812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_c_1556_n 0.0101121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_c_1557_n 0.00218029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB SUM 0.0506213f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=2.595
cc_101 VNB N_VPWR_c_1620_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_COUT_c_1751_n 0.00699949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_COUT_c_1752_n 8.11109e-19 $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_104 VNB COUT 0.0101428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_630_100#_c_1828_n 0.00361539f $X=-0.19 $Y=-0.245 $X2=1.15
+ $Y2=1.685
cc_106 VNB N_A_630_100#_c_1829_n 0.00424986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_630_100#_c_1830_n 0.00709765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_630_100#_c_1831_n 0.00444177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_630_100#_c_1832_n 9.71013e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_630_100#_c_1833_n 8.96325e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1741_367#_c_1922_n 0.00879914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1741_367#_c_1923_n 0.00259993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1741_367#_c_1924_n 0.00895234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1741_367#_c_1925_n 0.0043329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1930_367#_c_2000_n 0.00753676f $X=-0.19 $Y=-0.245 $X2=1.15
+ $Y2=1.52
cc_116 VNB N_A_1930_367#_c_2001_n 0.0218773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_1930_367#_c_2002_n 0.0248103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_1930_367#_c_2003_n 0.00342366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_1930_367#_c_2004_n 0.0051068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_1930_367#_c_2005_n 0.021787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_1930_367#_c_2006_n 0.0107992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_1930_367#_c_2007_n 0.00911522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_1930_367#_c_2008_n 0.0156508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_1930_367#_c_2009_n 0.00303914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2147_n 0.00691573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2148_n 0.0068452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2149_n 0.00240024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2150_n 0.0123441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2151_n 0.0208716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2152_n 0.0094787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2153_n 0.0331732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2154_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2155_n 0.12005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2156_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2157_n 0.0912446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2158_n 0.019419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2159_n 0.674331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2160_n 0.0242321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2161_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2162_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VPB N_CI_M1011_g 0.0301781f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=2.595
cc_142 VPB CI 0.002692f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_143 VPB N_CI_c_267_n 0.019211f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.685
cc_144 VPB N_A_84_21#_M1006_g 0.0266086f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_145 VPB N_A_84_21#_c_312_n 0.00961431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_84_21#_c_314_n 0.00635688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_84_21#_c_324_n 0.00334919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_84_21#_c_325_n 0.00191164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_84_21#_c_326_n 0.0569254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_413_34#_M1007_g 0.0288173f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.685
cc_151 VPB N_A_413_34#_c_475_n 0.00389446f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_239_135#_M1012_g 0.0242951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_239_135#_c_602_n 9.61058e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_239_135#_c_610_n 0.018552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_239_135#_c_611_n 0.0109021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_239_135#_c_604_n 0.00443506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_239_135#_c_605_n 0.0196026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_239_135#_c_614_n 0.0113313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_239_135#_c_615_n 0.00377976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_239_135#_c_616_n 0.00358628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_239_135#_c_617_n 0.0185092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_239_135#_c_606_n 0.00308106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_239_135#_c_619_n 0.00262887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_239_135#_c_620_n 0.025699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_239_135#_c_607_n 0.00847804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_239_135#_c_622_n 0.00365339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_239_135#_c_623_n 0.00223413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_239_135#_c_624_n 0.00474308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_814_384#_c_835_n 0.0236561f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=2.595
cc_170 VPB N_A_814_384#_c_836_n 0.0210147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_814_384#_c_837_n 0.00983547f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.685
cc_172 VPB N_A_814_384#_c_822_n 0.0175017f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.685
cc_173 VPB N_A_814_384#_M1020_g 0.02082f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_814_384#_c_829_n 0.0031259f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_814_384#_c_841_n 0.0358972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_814_384#_c_833_n 0.0114095f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_814_384#_c_834_n 0.00125253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_1022_362#_M1001_g 0.0191859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_1022_362#_c_1022_n 0.025247f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.685
cc_180 VPB N_A_1022_362#_M1002_g 7.0385e-19 $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.685
cc_181 VPB N_A_1022_362#_c_1024_n 0.0888675f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.85
cc_182 VPB N_A_1022_362#_c_1025_n 0.012806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_1022_362#_M1015_g 0.0300274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1022_362#_c_1010_n 0.010104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1022_362#_c_1012_n 0.00175116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_1022_362#_c_1029_n 4.62205e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_1022_362#_c_1013_n 0.00864616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_1022_362#_c_1014_n 6.16823e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1022_362#_c_1015_n 0.00306016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_1022_362#_c_1016_n 9.62012e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_1022_362#_c_1017_n 0.00210339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_1022_362#_c_1019_n 0.00187028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_1022_362#_c_1020_n 0.00147179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_878_41#_M1003_g 0.0214228f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.52
cc_195 VPB N_A_878_41#_M1029_g 0.0183575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_878_41#_c_1221_n 0.00248889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_878_41#_c_1216_n 0.00326277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_B_c_1363_n 0.0198206f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=1.52
cc_199 VPB N_B_c_1356_n 0.0108499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_B_c_1357_n 0.00233037f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=1.85
cc_201 VPB N_B_c_1366_n 0.106063f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.685
cc_202 VPB N_B_M1021_g 0.0322428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_B_c_1368_n 0.0785243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_B_M1009_g 0.0314238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_B_c_1361_n 0.00934522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_B_c_1371_n 0.0400916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_B_c_1372_n 0.0676772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_B_c_1362_n 0.00524511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_B_c_1374_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB B 0.00395253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_B_c_1376_n 0.0196649f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_2229_269#_M1000_g 0.0268417f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_213 VPB N_A_2229_269#_c_1484_n 0.0026525f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.85
cc_214 VPB N_A_2229_269#_c_1487_n 0.0573842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_2229_269#_c_1488_n 0.0127877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_2229_269#_c_1489_n 0.0167241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_M1030_g 0.0264267f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=2.595
cc_218 VPB N_A_c_1553_n 0.00387248f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_219 VPB N_A_M1016_g 0.0348695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_c_1555_n 0.00200062f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_c_1556_n 0.0208582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_c_1557_n 0.011021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB SUM 0.0543794f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=2.595
cc_224 VPB N_VPWR_c_1621_n 0.00472864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1622_n 0.0101576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1623_n 0.0061343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1624_n 0.0204211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1625_n 0.00589518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1626_n 0.0917945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1627_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1628_n 0.019006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1629_n 0.0499566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1630_n 0.1062f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1631_n 0.019006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1620_n 0.0990978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1633_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1634_n 0.012939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1635_n 0.00477762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1636_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_COUT_c_1751_n 0.00330126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_COUT_c_1755_n 0.0205296f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.685
cc_242 VPB N_COUT_c_1756_n 0.00678125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_COUT_c_1757_n 0.00818298f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_630_100#_c_1834_n 0.00187307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_630_100#_c_1835_n 0.00355719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_630_100#_c_1829_n 0.00424969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_630_100#_c_1830_n 0.0152359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_630_100#_c_1831_n 0.0041063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_630_100#_c_1832_n 0.00146889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_630_100#_c_1833_n 4.816e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_1741_367#_c_1926_n 0.00633645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_1741_367#_c_1923_n 0.00118214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_1741_367#_c_1924_n 0.00283953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_1741_367#_c_1929_n 0.00555065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_1930_367#_c_2000_n 0.0309923f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.52
cc_256 VPB N_A_1930_367#_c_2011_n 0.0268673f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.85
cc_257 VPB N_A_1930_367#_c_2012_n 0.0028212f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_1930_367#_c_2013_n 0.0104552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_1930_367#_c_2014_n 0.0149747f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_1930_367#_c_2015_n 0.0172311f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_1930_367#_c_2016_n 0.00670573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_1930_367#_c_2017_n 0.0115202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 N_CI_M1008_g N_A_84_21#_M1006_g 0.01808f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_264 N_CI_M1011_g N_A_84_21#_M1006_g 0.0161189f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_265 N_CI_c_267_n N_A_84_21#_M1006_g 0.00756426f $X=1.15 $Y=1.685 $X2=0 $Y2=0
cc_266 N_CI_M1008_g N_A_84_21#_c_309_n 0.00677271f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_267 N_CI_M1008_g N_A_84_21#_c_311_n 0.0212569f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_268 N_CI_M1008_g N_A_84_21#_c_312_n 0.00251755f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_269 N_CI_c_267_n N_A_84_21#_c_312_n 0.00939838f $X=1.15 $Y=1.685 $X2=0 $Y2=0
cc_270 N_CI_M1011_g N_A_84_21#_c_326_n 0.00679631f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_271 N_CI_M1008_g N_A_239_135#_c_603_n 0.00475569f $X=1.12 $Y=0.995 $X2=0
+ $Y2=0
cc_272 CI N_A_239_135#_c_603_n 0.0106549f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_273 N_CI_c_267_n N_A_239_135#_c_603_n 0.00299079f $X=1.15 $Y=1.685 $X2=0
+ $Y2=0
cc_274 N_CI_M1011_g N_A_239_135#_c_620_n 0.00385022f $X=1.195 $Y=2.595 $X2=0
+ $Y2=0
cc_275 N_CI_M1008_g N_A_239_135#_c_607_n 0.00342756f $X=1.12 $Y=0.995 $X2=0
+ $Y2=0
cc_276 N_CI_M1011_g N_A_239_135#_c_607_n 0.00405083f $X=1.195 $Y=2.595 $X2=0
+ $Y2=0
cc_277 CI N_A_239_135#_c_607_n 0.0237223f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_278 N_CI_c_267_n N_A_239_135#_c_607_n 0.00111728f $X=1.15 $Y=1.685 $X2=0
+ $Y2=0
cc_279 N_CI_M1008_g SUM 0.00103349f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_280 N_CI_M1011_g SUM 3.97314e-19 $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_281 N_CI_M1011_g N_VPWR_c_1621_n 0.00416667f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_282 N_CI_M1011_g N_VPWR_c_1629_n 0.0035993f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_283 N_CI_M1011_g N_VPWR_c_1620_n 0.0074086f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_284 N_CI_M1008_g N_COUT_c_1751_n 0.00956473f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_285 N_CI_M1011_g N_COUT_c_1751_n 0.00349088f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_286 CI N_COUT_c_1751_n 0.0237036f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_287 N_CI_c_267_n N_COUT_c_1751_n 0.00116619f $X=1.15 $Y=1.685 $X2=0 $Y2=0
cc_288 N_CI_M1008_g N_COUT_c_1752_n 0.0139357f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_289 CI N_COUT_c_1752_n 0.0039212f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_290 N_CI_c_267_n N_COUT_c_1752_n 7.78415e-19 $X=1.15 $Y=1.685 $X2=0 $Y2=0
cc_291 N_CI_M1011_g N_COUT_c_1765_n 0.0213813f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_292 N_CI_M1011_g N_COUT_c_1755_n 0.0126174f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_293 N_CI_M1011_g N_COUT_c_1767_n 0.00269071f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_294 N_CI_M1011_g N_COUT_c_1756_n 0.00535606f $X=1.195 $Y=2.595 $X2=0 $Y2=0
cc_295 CI N_COUT_c_1756_n 0.0114238f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_296 N_CI_c_267_n N_COUT_c_1756_n 0.00329966f $X=1.15 $Y=1.685 $X2=0 $Y2=0
cc_297 N_CI_M1008_g COUT 0.00389706f $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_298 N_CI_M1008_g N_VGND_c_2147_n 2.26657e-19 $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_299 N_CI_M1008_g N_VGND_c_2159_n 9.62932e-19 $X=1.12 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A_84_21#_c_320_n N_A_413_34#_M1024_d 0.00180746f $X=5.885 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_301 N_A_84_21#_c_309_n N_A_413_34#_c_464_n 0.0267621f $X=1.555 $Y=0.18 $X2=0
+ $Y2=0
cc_302 N_A_84_21#_c_313_n N_A_413_34#_c_464_n 0.00912851f $X=1.75 $Y=1.29 $X2=0
+ $Y2=0
cc_303 N_A_84_21#_c_314_n N_A_413_34#_c_464_n 0.0124006f $X=2.03 $Y=1.98 $X2=0
+ $Y2=0
cc_304 N_A_84_21#_c_339_p N_A_413_34#_c_464_n 0.00544507f $X=2.62 $Y=0.935 $X2=0
+ $Y2=0
cc_305 N_A_84_21#_c_340_p N_A_413_34#_c_464_n 0.00718881f $X=2.195 $Y=0.935
+ $X2=0 $Y2=0
cc_306 N_A_84_21#_c_315_n N_A_413_34#_c_464_n 0.00513999f $X=2.705 $Y=0.85 $X2=0
+ $Y2=0
cc_307 N_A_84_21#_c_314_n N_A_413_34#_M1007_g 0.00753769f $X=2.03 $Y=1.98 $X2=0
+ $Y2=0
cc_308 N_A_84_21#_c_324_n N_A_413_34#_M1007_g 0.0135342f $X=3.115 $Y=2.065 $X2=0
+ $Y2=0
cc_309 N_A_84_21#_c_326_n N_A_413_34#_M1007_g 0.00896958f $X=2.03 $Y=1.985 $X2=0
+ $Y2=0
cc_310 N_A_84_21#_c_345_p N_A_413_34#_M1007_g 0.00404575f $X=3.2 $Y=2.065 $X2=0
+ $Y2=0
cc_311 N_A_84_21#_c_312_n N_A_413_34#_c_466_n 0.00912851f $X=1.75 $Y=1.82 $X2=0
+ $Y2=0
cc_312 N_A_84_21#_c_314_n N_A_413_34#_c_466_n 0.0126376f $X=2.03 $Y=1.98 $X2=0
+ $Y2=0
cc_313 N_A_84_21#_c_324_n N_A_413_34#_c_466_n 0.00536233f $X=3.115 $Y=2.065
+ $X2=0 $Y2=0
cc_314 N_A_84_21#_c_326_n N_A_413_34#_c_466_n 0.007194f $X=2.03 $Y=1.985 $X2=0
+ $Y2=0
cc_315 N_A_84_21#_c_339_p N_A_413_34#_c_467_n 0.00677785f $X=2.62 $Y=0.935 $X2=0
+ $Y2=0
cc_316 N_A_84_21#_c_324_n N_A_413_34#_c_467_n 0.00135989f $X=3.115 $Y=2.065
+ $X2=0 $Y2=0
cc_317 N_A_84_21#_c_339_p N_A_413_34#_c_468_n 0.00669828f $X=2.62 $Y=0.935 $X2=0
+ $Y2=0
cc_318 N_A_84_21#_c_324_n N_A_413_34#_c_468_n 0.00731606f $X=3.115 $Y=2.065
+ $X2=0 $Y2=0
cc_319 N_A_84_21#_c_316_n N_A_413_34#_c_470_n 0.0461774f $X=4.02 $Y=0.35 $X2=0
+ $Y2=0
cc_320 N_A_84_21#_c_319_n N_A_413_34#_c_470_n 0.015292f $X=4.19 $Y=0.7 $X2=0
+ $Y2=0
cc_321 N_A_84_21#_c_316_n N_A_413_34#_c_500_n 0.0105755f $X=4.02 $Y=0.35 $X2=0
+ $Y2=0
cc_322 N_A_84_21#_c_316_n N_A_413_34#_c_472_n 0.00613197f $X=4.02 $Y=0.35 $X2=0
+ $Y2=0
cc_323 N_A_84_21#_c_319_n N_A_413_34#_c_472_n 0.0134868f $X=4.19 $Y=0.7 $X2=0
+ $Y2=0
cc_324 N_A_84_21#_c_320_n N_A_413_34#_c_472_n 0.0460187f $X=5.885 $Y=0.745 $X2=0
+ $Y2=0
cc_325 N_A_84_21#_c_320_n N_A_413_34#_c_474_n 0.0158737f $X=5.885 $Y=0.745 $X2=0
+ $Y2=0
cc_326 N_A_84_21#_c_314_n N_A_413_34#_c_476_n 0.02741f $X=2.03 $Y=1.98 $X2=0
+ $Y2=0
cc_327 N_A_84_21#_c_339_p N_A_413_34#_c_476_n 0.0255534f $X=2.62 $Y=0.935 $X2=0
+ $Y2=0
cc_328 N_A_84_21#_c_324_n N_A_413_34#_c_476_n 0.0114125f $X=3.115 $Y=2.065 $X2=0
+ $Y2=0
cc_329 N_A_84_21#_c_320_n N_A_239_135#_M1002_d 0.00179584f $X=5.885 $Y=0.745
+ $X2=0 $Y2=0
cc_330 N_A_84_21#_c_339_p N_A_239_135#_M1027_g 0.00125042f $X=2.62 $Y=0.935
+ $X2=0 $Y2=0
cc_331 N_A_84_21#_c_315_n N_A_239_135#_M1027_g 0.00742395f $X=2.705 $Y=0.85
+ $X2=0 $Y2=0
cc_332 N_A_84_21#_c_316_n N_A_239_135#_M1027_g 0.00836486f $X=4.02 $Y=0.35 $X2=0
+ $Y2=0
cc_333 N_A_84_21#_c_324_n N_A_239_135#_c_601_n 2.64639e-19 $X=3.115 $Y=2.065
+ $X2=0 $Y2=0
cc_334 N_A_84_21#_c_325_n N_A_239_135#_M1012_g 0.014071f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_335 N_A_84_21#_c_345_p N_A_239_135#_M1012_g 0.00598582f $X=3.2 $Y=2.065 $X2=0
+ $Y2=0
cc_336 N_A_84_21#_c_311_n N_A_239_135#_c_603_n 0.00546274f $X=1.63 $Y=1.215
+ $X2=0 $Y2=0
cc_337 N_A_84_21#_c_313_n N_A_239_135#_c_603_n 0.00425009f $X=1.75 $Y=1.29 $X2=0
+ $Y2=0
cc_338 N_A_84_21#_c_314_n N_A_239_135#_c_603_n 0.0180049f $X=2.03 $Y=1.98 $X2=0
+ $Y2=0
cc_339 N_A_84_21#_c_314_n N_A_239_135#_c_610_n 0.02525f $X=2.03 $Y=1.98 $X2=0
+ $Y2=0
cc_340 N_A_84_21#_c_324_n N_A_239_135#_c_610_n 0.0355007f $X=3.115 $Y=2.065
+ $X2=0 $Y2=0
cc_341 N_A_84_21#_c_326_n N_A_239_135#_c_610_n 0.00994314f $X=2.03 $Y=1.985
+ $X2=0 $Y2=0
cc_342 N_A_84_21#_c_324_n N_A_239_135#_c_646_n 0.00621732f $X=3.115 $Y=2.065
+ $X2=0 $Y2=0
cc_343 N_A_84_21#_c_325_n N_A_239_135#_c_646_n 0.00473359f $X=4.195 $Y=2.35
+ $X2=0 $Y2=0
cc_344 N_A_84_21#_c_345_p N_A_239_135#_c_646_n 0.0126782f $X=3.2 $Y=2.065 $X2=0
+ $Y2=0
cc_345 N_A_84_21#_M1013_d N_A_239_135#_c_611_n 0.0101919f $X=4.22 $Y=2.18 $X2=0
+ $Y2=0
cc_346 N_A_84_21#_c_325_n N_A_239_135#_c_611_n 0.0391726f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_347 N_A_84_21#_c_325_n N_A_239_135#_c_604_n 0.0139378f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_348 N_A_84_21#_c_325_n N_A_239_135#_c_605_n 0.00139764f $X=4.195 $Y=2.35
+ $X2=0 $Y2=0
cc_349 N_A_84_21#_c_325_n N_A_239_135#_c_614_n 0.0138936f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_350 N_A_84_21#_M1013_d N_A_239_135#_c_615_n 0.0154493f $X=4.22 $Y=2.18 $X2=0
+ $Y2=0
cc_351 N_A_84_21#_c_325_n N_A_239_135#_c_615_n 0.0390286f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_352 N_A_84_21#_M1013_d N_A_239_135#_c_616_n 0.00813852f $X=4.22 $Y=2.18 $X2=0
+ $Y2=0
cc_353 N_A_84_21#_M1023_d N_A_239_135#_c_657_n 0.00586748f $X=5.795 $Y=0.635
+ $X2=0 $Y2=0
cc_354 N_A_84_21#_c_389_p N_A_239_135#_c_657_n 0.0203695f $X=6.05 $Y=0.705 $X2=0
+ $Y2=0
cc_355 N_A_84_21#_c_320_n N_A_239_135#_c_657_n 0.00753374f $X=5.885 $Y=0.745
+ $X2=0 $Y2=0
cc_356 N_A_84_21#_c_326_n N_A_239_135#_c_620_n 0.00420399f $X=2.03 $Y=1.985
+ $X2=0 $Y2=0
cc_357 N_A_84_21#_c_312_n N_A_239_135#_c_607_n 0.00420399f $X=1.75 $Y=1.82 $X2=0
+ $Y2=0
cc_358 N_A_84_21#_c_313_n N_A_239_135#_c_607_n 0.00337045f $X=1.75 $Y=1.29 $X2=0
+ $Y2=0
cc_359 N_A_84_21#_c_314_n N_A_239_135#_c_607_n 0.0566542f $X=2.03 $Y=1.98 $X2=0
+ $Y2=0
cc_360 N_A_84_21#_c_324_n N_A_239_135#_c_664_n 0.00825407f $X=3.115 $Y=2.065
+ $X2=0 $Y2=0
cc_361 N_A_84_21#_c_345_p N_A_239_135#_c_664_n 0.00730917f $X=3.2 $Y=2.065 $X2=0
+ $Y2=0
cc_362 N_A_84_21#_c_325_n N_A_239_135#_c_622_n 0.0102862f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_363 N_A_84_21#_M1013_d N_A_239_135#_c_623_n 0.0057469f $X=4.22 $Y=2.18 $X2=0
+ $Y2=0
cc_364 N_A_84_21#_c_325_n N_A_239_135#_c_623_n 0.00286911f $X=4.195 $Y=2.35
+ $X2=0 $Y2=0
cc_365 N_A_84_21#_c_320_n N_A_239_135#_c_669_n 0.015151f $X=5.885 $Y=0.745 $X2=0
+ $Y2=0
cc_366 N_A_84_21#_c_325_n N_A_814_384#_c_835_n 0.0230835f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_367 N_A_84_21#_c_325_n N_A_814_384#_c_836_n 0.0077669f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_368 N_A_84_21#_c_316_n N_A_814_384#_M1024_g 5.82496e-19 $X=4.02 $Y=0.35 $X2=0
+ $Y2=0
cc_369 N_A_84_21#_c_318_n N_A_814_384#_M1024_g 0.00394112f $X=4.105 $Y=0.615
+ $X2=0 $Y2=0
cc_370 N_A_84_21#_c_320_n N_A_814_384#_M1024_g 0.0125784f $X=5.885 $Y=0.745
+ $X2=0 $Y2=0
cc_371 N_A_84_21#_c_389_p N_A_814_384#_M1023_g 0.00243626f $X=6.05 $Y=0.705
+ $X2=0 $Y2=0
cc_372 N_A_84_21#_c_320_n N_A_814_384#_M1023_g 0.0114977f $X=5.885 $Y=0.745
+ $X2=0 $Y2=0
cc_373 N_A_84_21#_c_325_n N_A_1022_362#_M1001_g 3.51891e-19 $X=4.195 $Y=2.35
+ $X2=0 $Y2=0
cc_374 N_A_84_21#_c_320_n N_A_1022_362#_M1002_g 0.0131777f $X=5.885 $Y=0.745
+ $X2=0 $Y2=0
cc_375 N_A_84_21#_c_389_p N_A_1022_362#_c_1011_n 0.00343372f $X=6.05 $Y=0.705
+ $X2=0 $Y2=0
cc_376 N_A_84_21#_c_320_n N_A_878_41#_M1024_s 0.00834201f $X=5.885 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_377 N_A_84_21#_c_316_n N_A_878_41#_c_1215_n 0.015112f $X=4.02 $Y=0.35 $X2=0
+ $Y2=0
cc_378 N_A_84_21#_c_320_n N_A_878_41#_c_1215_n 0.119979f $X=5.885 $Y=0.745 $X2=0
+ $Y2=0
cc_379 N_A_84_21#_M1006_g SUM 0.0495654f $X=0.495 $Y=0.895 $X2=0 $Y2=0
cc_380 N_A_84_21#_c_324_n N_VPWR_M1007_d 0.0099129f $X=3.115 $Y=2.065 $X2=0
+ $Y2=0
cc_381 N_A_84_21#_c_325_n N_VPWR_M1007_d 0.00234735f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_382 N_A_84_21#_c_345_p N_VPWR_M1007_d 0.0137375f $X=3.2 $Y=2.065 $X2=0 $Y2=0
cc_383 N_A_84_21#_M1006_g N_VPWR_c_1621_n 0.00318456f $X=0.495 $Y=0.895 $X2=0
+ $Y2=0
cc_384 N_A_84_21#_M1006_g N_VPWR_c_1628_n 0.00549284f $X=0.495 $Y=0.895 $X2=0
+ $Y2=0
cc_385 N_A_84_21#_M1006_g N_VPWR_c_1620_n 0.0112878f $X=0.495 $Y=0.895 $X2=0
+ $Y2=0
cc_386 N_A_84_21#_c_314_n N_COUT_M1004_s 0.00142984f $X=2.03 $Y=1.98 $X2=-0.19
+ $Y2=-0.245
cc_387 N_A_84_21#_c_340_p N_COUT_M1004_s 0.00380799f $X=2.195 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_388 N_A_84_21#_c_324_n N_COUT_M1007_s 0.00630559f $X=3.115 $Y=2.065 $X2=0
+ $Y2=0
cc_389 N_A_84_21#_M1006_g N_COUT_c_1751_n 0.0105151f $X=0.495 $Y=0.895 $X2=0
+ $Y2=0
cc_390 N_A_84_21#_c_309_n N_COUT_c_1752_n 0.00522411f $X=1.555 $Y=0.18 $X2=0
+ $Y2=0
cc_391 N_A_84_21#_M1006_g N_COUT_c_1777_n 0.00181036f $X=0.495 $Y=0.895 $X2=0
+ $Y2=0
cc_392 N_A_84_21#_c_309_n N_COUT_c_1777_n 6.01197e-19 $X=1.555 $Y=0.18 $X2=0
+ $Y2=0
cc_393 N_A_84_21#_M1006_g N_COUT_c_1765_n 0.00205192f $X=0.495 $Y=0.895 $X2=0
+ $Y2=0
cc_394 N_A_84_21#_M1006_g N_COUT_c_1756_n 0.00186964f $X=0.495 $Y=0.895 $X2=0
+ $Y2=0
cc_395 N_A_84_21#_c_311_n COUT 0.028129f $X=1.63 $Y=1.215 $X2=0 $Y2=0
cc_396 N_A_84_21#_c_313_n COUT 0.00358026f $X=1.75 $Y=1.29 $X2=0 $Y2=0
cc_397 N_A_84_21#_c_340_p COUT 0.0183828f $X=2.195 $Y=0.935 $X2=0 $Y2=0
cc_398 N_A_84_21#_c_325_n N_A_630_100#_M1012_d 0.0122961f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_399 N_A_84_21#_c_325_n N_A_630_100#_c_1834_n 0.023122f $X=4.195 $Y=2.35 $X2=0
+ $Y2=0
cc_400 N_A_84_21#_c_325_n N_A_630_100#_c_1835_n 0.0117061f $X=4.195 $Y=2.35
+ $X2=0 $Y2=0
cc_401 N_A_84_21#_c_345_p N_A_630_100#_c_1835_n 0.00771996f $X=3.2 $Y=2.065
+ $X2=0 $Y2=0
cc_402 N_A_84_21#_c_324_n N_A_630_100#_c_1829_n 0.00606409f $X=3.115 $Y=2.065
+ $X2=0 $Y2=0
cc_403 N_A_84_21#_c_325_n N_A_630_100#_c_1829_n 0.00101346f $X=4.195 $Y=2.35
+ $X2=0 $Y2=0
cc_404 N_A_84_21#_c_345_p N_A_630_100#_c_1829_n 0.0100815f $X=3.2 $Y=2.065 $X2=0
+ $Y2=0
cc_405 N_A_84_21#_c_325_n N_A_630_100#_c_1830_n 0.00721722f $X=4.195 $Y=2.35
+ $X2=0 $Y2=0
cc_406 N_A_84_21#_c_324_n N_A_630_100#_c_1831_n 0.00394086f $X=3.115 $Y=2.065
+ $X2=0 $Y2=0
cc_407 N_A_84_21#_c_345_p N_A_630_100#_c_1831_n 0.00413369f $X=3.2 $Y=2.065
+ $X2=0 $Y2=0
cc_408 N_A_84_21#_c_339_p N_VGND_M1004_d 0.0156168f $X=2.62 $Y=0.935 $X2=0 $Y2=0
cc_409 N_A_84_21#_c_315_n N_VGND_M1004_d 0.0107692f $X=2.705 $Y=0.85 $X2=0 $Y2=0
cc_410 N_A_84_21#_M1006_g N_VGND_c_2147_n 0.00994265f $X=0.495 $Y=0.895 $X2=0
+ $Y2=0
cc_411 N_A_84_21#_c_309_n N_VGND_c_2147_n 0.0244116f $X=1.555 $Y=0.18 $X2=0
+ $Y2=0
cc_412 N_A_84_21#_c_311_n N_VGND_c_2147_n 0.00512344f $X=1.63 $Y=1.215 $X2=0
+ $Y2=0
cc_413 N_A_84_21#_c_309_n N_VGND_c_2148_n 0.00116299f $X=1.555 $Y=0.18 $X2=0
+ $Y2=0
cc_414 N_A_84_21#_c_339_p N_VGND_c_2148_n 0.0126932f $X=2.62 $Y=0.935 $X2=0
+ $Y2=0
cc_415 N_A_84_21#_c_315_n N_VGND_c_2148_n 0.0164107f $X=2.705 $Y=0.85 $X2=0
+ $Y2=0
cc_416 N_A_84_21#_c_317_n N_VGND_c_2148_n 0.0136044f $X=2.79 $Y=0.35 $X2=0 $Y2=0
cc_417 N_A_84_21#_c_309_n N_VGND_c_2153_n 0.0185787f $X=1.555 $Y=0.18 $X2=0
+ $Y2=0
cc_418 N_A_84_21#_c_316_n N_VGND_c_2155_n 0.0857601f $X=4.02 $Y=0.35 $X2=0 $Y2=0
cc_419 N_A_84_21#_c_317_n N_VGND_c_2155_n 0.0114622f $X=2.79 $Y=0.35 $X2=0 $Y2=0
cc_420 N_A_84_21#_c_320_n N_VGND_c_2155_n 0.00341774f $X=5.885 $Y=0.745 $X2=0
+ $Y2=0
cc_421 N_A_84_21#_c_309_n N_VGND_c_2159_n 0.0256835f $X=1.555 $Y=0.18 $X2=0
+ $Y2=0
cc_422 N_A_84_21#_c_310_n N_VGND_c_2159_n 0.0102634f $X=0.57 $Y=0.18 $X2=0 $Y2=0
cc_423 N_A_84_21#_c_339_p N_VGND_c_2159_n 0.00917716f $X=2.62 $Y=0.935 $X2=0
+ $Y2=0
cc_424 N_A_84_21#_c_340_p N_VGND_c_2159_n 0.00371697f $X=2.195 $Y=0.935 $X2=0
+ $Y2=0
cc_425 N_A_84_21#_c_316_n N_VGND_c_2159_n 0.0524914f $X=4.02 $Y=0.35 $X2=0 $Y2=0
cc_426 N_A_84_21#_c_317_n N_VGND_c_2159_n 0.00657784f $X=2.79 $Y=0.35 $X2=0
+ $Y2=0
cc_427 N_A_84_21#_c_320_n N_VGND_c_2159_n 0.00903773f $X=5.885 $Y=0.745 $X2=0
+ $Y2=0
cc_428 N_A_84_21#_c_310_n N_VGND_c_2160_n 0.00878687f $X=0.57 $Y=0.18 $X2=0
+ $Y2=0
cc_429 N_A_413_34#_c_508_p N_A_239_135#_M1001_d 0.00934241f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_430 N_A_413_34#_c_467_n N_A_239_135#_M1027_g 0.00798237f $X=2.64 $Y=1.415
+ $X2=0 $Y2=0
cc_431 N_A_413_34#_c_468_n N_A_239_135#_M1027_g 0.00493827f $X=2.97 $Y=1.285
+ $X2=0 $Y2=0
cc_432 N_A_413_34#_c_469_n N_A_239_135#_M1027_g 0.0151722f $X=3.055 $Y=1.2 $X2=0
+ $Y2=0
cc_433 N_A_413_34#_c_470_n N_A_239_135#_M1027_g 0.00465567f $X=3.67 $Y=0.7 $X2=0
+ $Y2=0
cc_434 N_A_413_34#_c_500_n N_A_239_135#_M1027_g 0.0067697f $X=3.14 $Y=0.7 $X2=0
+ $Y2=0
cc_435 N_A_413_34#_c_471_n N_A_239_135#_M1027_g 0.00268188f $X=3.755 $Y=0.965
+ $X2=0 $Y2=0
cc_436 N_A_413_34#_c_476_n N_A_239_135#_M1027_g 2.60688e-19 $X=2.54 $Y=1.285
+ $X2=0 $Y2=0
cc_437 N_A_413_34#_c_470_n N_A_239_135#_c_600_n 0.00374308f $X=3.67 $Y=0.7 $X2=0
+ $Y2=0
cc_438 N_A_413_34#_c_467_n N_A_239_135#_c_601_n 0.0051484f $X=2.64 $Y=1.415
+ $X2=0 $Y2=0
cc_439 N_A_413_34#_c_468_n N_A_239_135#_c_601_n 0.00198625f $X=2.97 $Y=1.285
+ $X2=0 $Y2=0
cc_440 N_A_413_34#_c_476_n N_A_239_135#_c_601_n 5.96225e-19 $X=2.54 $Y=1.285
+ $X2=0 $Y2=0
cc_441 N_A_413_34#_M1007_g N_A_239_135#_M1012_g 0.00996f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_442 N_A_413_34#_c_467_n N_A_239_135#_c_602_n 0.00996f $X=2.64 $Y=1.415 $X2=0
+ $Y2=0
cc_443 N_A_413_34#_c_470_n N_A_239_135#_c_602_n 0.00466623f $X=3.67 $Y=0.7 $X2=0
+ $Y2=0
cc_444 N_A_413_34#_c_464_n N_A_239_135#_c_603_n 2.02782e-19 $X=2.14 $Y=1.25
+ $X2=0 $Y2=0
cc_445 N_A_413_34#_M1007_g N_A_239_135#_c_610_n 0.0112872f $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_446 N_A_413_34#_M1007_g N_A_239_135#_c_646_n 3.63963e-19 $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_447 N_A_413_34#_c_472_n N_A_239_135#_c_604_n 0.0300196f $X=4.91 $Y=1.05 $X2=0
+ $Y2=0
cc_448 N_A_413_34#_c_473_n N_A_239_135#_c_604_n 0.00159986f $X=3.84 $Y=1.05
+ $X2=0 $Y2=0
cc_449 N_A_413_34#_c_474_n N_A_239_135#_c_604_n 0.00659115f $X=5.14 $Y=1.575
+ $X2=0 $Y2=0
cc_450 N_A_413_34#_c_472_n N_A_239_135#_c_605_n 0.00663482f $X=4.91 $Y=1.05
+ $X2=0 $Y2=0
cc_451 N_A_413_34#_c_473_n N_A_239_135#_c_605_n 0.00646281f $X=3.84 $Y=1.05
+ $X2=0 $Y2=0
cc_452 N_A_413_34#_c_472_n N_A_239_135#_c_614_n 0.00538793f $X=4.91 $Y=1.05
+ $X2=0 $Y2=0
cc_453 N_A_413_34#_c_475_n N_A_239_135#_c_614_n 0.0133285f $X=5.14 $Y=2.33 $X2=0
+ $Y2=0
cc_454 N_A_413_34#_c_475_n N_A_239_135#_c_615_n 0.014994f $X=5.14 $Y=2.33 $X2=0
+ $Y2=0
cc_455 N_A_413_34#_c_508_p N_A_239_135#_c_616_n 0.0275461f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_456 N_A_413_34#_c_535_p N_A_239_135#_c_616_n 0.0085493f $X=5.225 $Y=2.415
+ $X2=0 $Y2=0
cc_457 N_A_413_34#_c_508_p N_A_239_135#_c_617_n 0.00650443f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_458 N_A_413_34#_c_537_p N_A_239_135#_c_617_n 0.0212041f $X=6.06 $Y=2.415
+ $X2=0 $Y2=0
cc_459 N_A_413_34#_M1020_d N_A_239_135#_c_606_n 0.00189078f $X=5.92 $Y=1.895
+ $X2=0 $Y2=0
cc_460 N_A_413_34#_M1020_d N_A_239_135#_c_701_n 0.00705353f $X=5.92 $Y=1.895
+ $X2=0 $Y2=0
cc_461 N_A_413_34#_c_537_p N_A_239_135#_c_701_n 5.15915e-19 $X=6.06 $Y=2.415
+ $X2=0 $Y2=0
cc_462 N_A_413_34#_M1020_d N_A_239_135#_c_703_n 0.0045457f $X=5.92 $Y=1.895
+ $X2=0 $Y2=0
cc_463 N_A_413_34#_c_537_p N_A_239_135#_c_703_n 0.0115951f $X=6.06 $Y=2.415
+ $X2=0 $Y2=0
cc_464 N_A_413_34#_M1007_g N_A_239_135#_c_664_n 0.0160859f $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_465 N_A_413_34#_M1007_g N_A_239_135#_c_622_n 0.00196294f $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_466 N_A_413_34#_c_537_p N_A_239_135#_c_624_n 0.0023425f $X=6.06 $Y=2.415
+ $X2=0 $Y2=0
cc_467 N_A_413_34#_c_474_n N_A_814_384#_c_822_n 3.52734e-19 $X=5.14 $Y=1.575
+ $X2=0 $Y2=0
cc_468 N_A_413_34#_c_475_n N_A_814_384#_c_822_n 0.00313711f $X=5.14 $Y=2.33
+ $X2=0 $Y2=0
cc_469 N_A_413_34#_c_472_n N_A_814_384#_c_824_n 0.00926189f $X=4.91 $Y=1.05
+ $X2=0 $Y2=0
cc_470 N_A_413_34#_c_472_n N_A_814_384#_M1024_g 0.0105745f $X=4.91 $Y=1.05 $X2=0
+ $Y2=0
cc_471 N_A_413_34#_c_474_n N_A_814_384#_M1024_g 0.0120978f $X=5.14 $Y=1.575
+ $X2=0 $Y2=0
cc_472 N_A_413_34#_c_475_n N_A_814_384#_M1020_g 0.00120918f $X=5.14 $Y=2.33
+ $X2=0 $Y2=0
cc_473 N_A_413_34#_c_508_p N_A_814_384#_M1020_g 0.00945637f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_474 N_A_413_34#_c_537_p N_A_814_384#_M1020_g 0.00584239f $X=6.06 $Y=2.415
+ $X2=0 $Y2=0
cc_475 N_A_413_34#_M1020_d N_A_814_384#_c_841_n 0.00224221f $X=5.92 $Y=1.895
+ $X2=0 $Y2=0
cc_476 N_A_413_34#_c_508_p N_A_814_384#_c_841_n 0.0024191f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_477 N_A_413_34#_c_537_p N_A_814_384#_c_841_n 0.00812057f $X=6.06 $Y=2.415
+ $X2=0 $Y2=0
cc_478 N_A_413_34#_c_475_n N_A_814_384#_c_862_n 0.00730974f $X=5.14 $Y=2.33
+ $X2=0 $Y2=0
cc_479 N_A_413_34#_c_508_p N_A_814_384#_c_862_n 0.00342731f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_480 N_A_413_34#_c_508_p N_A_814_384#_c_833_n 5.21532e-19 $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_481 N_A_413_34#_c_474_n N_A_814_384#_c_834_n 0.0129882f $X=5.14 $Y=1.575
+ $X2=0 $Y2=0
cc_482 N_A_413_34#_c_475_n N_A_814_384#_c_834_n 0.0376745f $X=5.14 $Y=2.33 $X2=0
+ $Y2=0
cc_483 N_A_413_34#_c_508_p N_A_814_384#_c_834_n 0.0256061f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_484 N_A_413_34#_c_475_n N_A_1022_362#_M1001_g 0.0129338f $X=5.14 $Y=2.33
+ $X2=0 $Y2=0
cc_485 N_A_413_34#_c_508_p N_A_1022_362#_M1001_g 0.00481824f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_486 N_A_413_34#_c_535_p N_A_1022_362#_M1001_g 0.00611372f $X=5.225 $Y=2.415
+ $X2=0 $Y2=0
cc_487 N_A_413_34#_c_537_p N_A_1022_362#_M1001_g 8.87795e-19 $X=6.06 $Y=2.415
+ $X2=0 $Y2=0
cc_488 N_A_413_34#_c_475_n N_A_1022_362#_c_1022_n 0.0101083f $X=5.14 $Y=2.33
+ $X2=0 $Y2=0
cc_489 N_A_413_34#_c_508_p N_A_1022_362#_c_1022_n 0.00176769f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_490 N_A_413_34#_c_474_n N_A_1022_362#_M1002_g 0.00680228f $X=5.14 $Y=1.575
+ $X2=0 $Y2=0
cc_491 N_A_413_34#_c_475_n N_A_1022_362#_M1002_g 0.00194007f $X=5.14 $Y=2.33
+ $X2=0 $Y2=0
cc_492 N_A_413_34#_c_537_p N_A_1022_362#_M1015_g 0.00150204f $X=6.06 $Y=2.415
+ $X2=0 $Y2=0
cc_493 N_A_413_34#_c_472_n N_A_878_41#_M1024_s 0.010474f $X=4.91 $Y=1.05
+ $X2=-0.19 $Y2=-0.245
cc_494 N_A_413_34#_M1007_g N_VPWR_c_1629_n 0.00557495f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_495 N_A_413_34#_M1007_g N_VPWR_c_1620_n 0.00906012f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_496 N_A_413_34#_M1007_g N_VPWR_c_1634_n 0.00682443f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_497 N_A_413_34#_c_464_n COUT 0.00613463f $X=2.14 $Y=1.25 $X2=0 $Y2=0
cc_498 N_A_413_34#_c_470_n N_A_630_100#_M1027_d 0.0101306f $X=3.67 $Y=0.7
+ $X2=-0.19 $Y2=-0.245
cc_499 N_A_413_34#_c_467_n N_A_630_100#_c_1828_n 7.83949e-19 $X=2.64 $Y=1.415
+ $X2=0 $Y2=0
cc_500 N_A_413_34#_c_468_n N_A_630_100#_c_1828_n 0.0123497f $X=2.97 $Y=1.285
+ $X2=0 $Y2=0
cc_501 N_A_413_34#_c_469_n N_A_630_100#_c_1828_n 0.0157539f $X=3.055 $Y=1.2
+ $X2=0 $Y2=0
cc_502 N_A_413_34#_c_470_n N_A_630_100#_c_1828_n 0.0130962f $X=3.67 $Y=0.7 $X2=0
+ $Y2=0
cc_503 N_A_413_34#_c_473_n N_A_630_100#_c_1828_n 0.0135573f $X=3.84 $Y=1.05
+ $X2=0 $Y2=0
cc_504 N_A_413_34#_c_476_n N_A_630_100#_c_1828_n 0.00462246f $X=2.54 $Y=1.285
+ $X2=0 $Y2=0
cc_505 N_A_413_34#_M1007_g N_A_630_100#_c_1835_n 9.09487e-19 $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_506 N_A_413_34#_c_467_n N_A_630_100#_c_1829_n 0.00446779f $X=2.64 $Y=1.415
+ $X2=0 $Y2=0
cc_507 N_A_413_34#_c_468_n N_A_630_100#_c_1829_n 0.008899f $X=2.97 $Y=1.285
+ $X2=0 $Y2=0
cc_508 N_A_413_34#_c_476_n N_A_630_100#_c_1829_n 0.00106557f $X=2.54 $Y=1.285
+ $X2=0 $Y2=0
cc_509 N_A_413_34#_c_472_n N_A_630_100#_c_1830_n 0.0151468f $X=4.91 $Y=1.05
+ $X2=0 $Y2=0
cc_510 N_A_413_34#_c_473_n N_A_630_100#_c_1830_n 0.0052377f $X=3.84 $Y=1.05
+ $X2=0 $Y2=0
cc_511 N_A_413_34#_c_474_n N_A_630_100#_c_1830_n 0.0072787f $X=5.14 $Y=1.575
+ $X2=0 $Y2=0
cc_512 N_A_413_34#_c_475_n N_A_630_100#_c_1830_n 0.0252167f $X=5.14 $Y=2.33
+ $X2=0 $Y2=0
cc_513 N_A_413_34#_c_508_p N_A_630_100#_c_1830_n 0.00401661f $X=5.895 $Y=2.415
+ $X2=0 $Y2=0
cc_514 N_A_413_34#_c_467_n N_A_630_100#_c_1831_n 0.0045856f $X=2.64 $Y=1.415
+ $X2=0 $Y2=0
cc_515 N_A_413_34#_c_468_n N_A_630_100#_c_1831_n 0.0048122f $X=2.97 $Y=1.285
+ $X2=0 $Y2=0
cc_516 N_A_413_34#_c_476_n N_A_630_100#_c_1831_n 8.30352e-19 $X=2.54 $Y=1.285
+ $X2=0 $Y2=0
cc_517 N_A_413_34#_c_464_n N_VGND_c_2148_n 0.00428593f $X=2.14 $Y=1.25 $X2=0
+ $Y2=0
cc_518 N_A_413_34#_c_464_n N_VGND_c_2153_n 0.00488547f $X=2.14 $Y=1.25 $X2=0
+ $Y2=0
cc_519 N_A_413_34#_c_464_n N_VGND_c_2159_n 0.00639623f $X=2.14 $Y=1.25 $X2=0
+ $Y2=0
cc_520 N_A_239_135#_c_611_n N_A_814_384#_c_835_n 0.0142046f $X=4.705 $Y=2.98
+ $X2=0 $Y2=0
cc_521 N_A_239_135#_c_615_n N_A_814_384#_c_835_n 0.00317834f $X=4.79 $Y=2.68
+ $X2=0 $Y2=0
cc_522 N_A_239_135#_c_622_n N_A_814_384#_c_835_n 0.00149307f $X=3.44 $Y=2.7
+ $X2=0 $Y2=0
cc_523 N_A_239_135#_c_623_n N_A_814_384#_c_835_n 0.00546129f $X=4.79 $Y=2.872
+ $X2=0 $Y2=0
cc_524 N_A_239_135#_c_604_n N_A_814_384#_c_836_n 0.004123f $X=4.16 $Y=1.515
+ $X2=0 $Y2=0
cc_525 N_A_239_135#_c_614_n N_A_814_384#_c_836_n 0.00522187f $X=4.705 $Y=1.895
+ $X2=0 $Y2=0
cc_526 N_A_239_135#_c_615_n N_A_814_384#_c_836_n 0.00225935f $X=4.79 $Y=2.68
+ $X2=0 $Y2=0
cc_527 N_A_239_135#_M1012_g N_A_814_384#_c_837_n 0.0232483f $X=3.485 $Y=2.355
+ $X2=0 $Y2=0
cc_528 N_A_239_135#_c_604_n N_A_814_384#_c_837_n 0.00406923f $X=4.16 $Y=1.515
+ $X2=0 $Y2=0
cc_529 N_A_239_135#_c_605_n N_A_814_384#_c_837_n 0.00447514f $X=3.98 $Y=1.515
+ $X2=0 $Y2=0
cc_530 N_A_239_135#_c_604_n N_A_814_384#_c_822_n 9.67199e-19 $X=4.16 $Y=1.515
+ $X2=0 $Y2=0
cc_531 N_A_239_135#_c_614_n N_A_814_384#_c_822_n 0.00813083f $X=4.705 $Y=1.895
+ $X2=0 $Y2=0
cc_532 N_A_239_135#_c_614_n N_A_814_384#_c_823_n 0.0081019f $X=4.705 $Y=1.895
+ $X2=0 $Y2=0
cc_533 N_A_239_135#_c_604_n N_A_814_384#_c_824_n 0.00946908f $X=4.16 $Y=1.515
+ $X2=0 $Y2=0
cc_534 N_A_239_135#_c_605_n N_A_814_384#_c_824_n 0.0159641f $X=3.98 $Y=1.515
+ $X2=0 $Y2=0
cc_535 N_A_239_135#_c_604_n N_A_814_384#_M1024_g 2.88674e-19 $X=4.16 $Y=1.515
+ $X2=0 $Y2=0
cc_536 N_A_239_135#_c_605_n N_A_814_384#_M1024_g 4.29061e-19 $X=3.98 $Y=1.515
+ $X2=0 $Y2=0
cc_537 N_A_239_135#_c_657_n N_A_814_384#_M1023_g 0.00895042f $X=6.045 $Y=1.14
+ $X2=0 $Y2=0
cc_538 N_A_239_135#_c_606_n N_A_814_384#_M1023_g 0.00354331f $X=6.13 $Y=1.96
+ $X2=0 $Y2=0
cc_539 N_A_239_135#_c_669_n N_A_814_384#_M1023_g 0.00333487f $X=5.505 $Y=1.055
+ $X2=0 $Y2=0
cc_540 N_A_239_135#_c_617_n N_A_814_384#_M1020_g 0.0015962f $X=6.405 $Y=2.98
+ $X2=0 $Y2=0
cc_541 N_A_239_135#_c_703_n N_A_814_384#_M1020_g 0.00131905f $X=6.215 $Y=2.045
+ $X2=0 $Y2=0
cc_542 N_A_239_135#_c_619_n N_A_814_384#_M1020_g 0.00208853f $X=6.49 $Y=2.895
+ $X2=0 $Y2=0
cc_543 N_A_239_135#_c_624_n N_A_814_384#_M1020_g 0.00530899f $X=5.68 $Y=2.872
+ $X2=0 $Y2=0
cc_544 N_A_239_135#_c_701_n N_A_814_384#_c_841_n 0.0259204f $X=6.405 $Y=2.045
+ $X2=0 $Y2=0
cc_545 N_A_239_135#_c_703_n N_A_814_384#_c_841_n 0.00890646f $X=6.215 $Y=2.045
+ $X2=0 $Y2=0
cc_546 N_A_239_135#_M1001_d N_A_814_384#_c_862_n 0.00468123f $X=5.26 $Y=2.07
+ $X2=0 $Y2=0
cc_547 N_A_239_135#_c_657_n N_A_814_384#_c_833_n 0.00264494f $X=6.045 $Y=1.14
+ $X2=0 $Y2=0
cc_548 N_A_239_135#_c_606_n N_A_814_384#_c_833_n 0.00506921f $X=6.13 $Y=1.96
+ $X2=0 $Y2=0
cc_549 N_A_239_135#_c_669_n N_A_814_384#_c_833_n 3.62853e-19 $X=5.505 $Y=1.055
+ $X2=0 $Y2=0
cc_550 N_A_239_135#_M1001_d N_A_814_384#_c_834_n 0.0056104f $X=5.26 $Y=2.07
+ $X2=0 $Y2=0
cc_551 N_A_239_135#_c_657_n N_A_814_384#_c_834_n 0.011734f $X=6.045 $Y=1.14
+ $X2=0 $Y2=0
cc_552 N_A_239_135#_c_606_n N_A_814_384#_c_834_n 0.0389823f $X=6.13 $Y=1.96
+ $X2=0 $Y2=0
cc_553 N_A_239_135#_c_703_n N_A_814_384#_c_834_n 0.0112195f $X=6.215 $Y=2.045
+ $X2=0 $Y2=0
cc_554 N_A_239_135#_c_669_n N_A_814_384#_c_834_n 0.0175584f $X=5.505 $Y=1.055
+ $X2=0 $Y2=0
cc_555 N_A_239_135#_c_615_n N_A_1022_362#_M1001_g 0.00867629f $X=4.79 $Y=2.68
+ $X2=0 $Y2=0
cc_556 N_A_239_135#_c_616_n N_A_1022_362#_M1001_g 0.0253469f $X=5.488 $Y=2.872
+ $X2=0 $Y2=0
cc_557 N_A_239_135#_c_614_n N_A_1022_362#_c_1022_n 6.89735e-19 $X=4.705 $Y=1.895
+ $X2=0 $Y2=0
cc_558 N_A_239_135#_c_669_n N_A_1022_362#_M1002_g 0.00345054f $X=5.505 $Y=1.055
+ $X2=0 $Y2=0
cc_559 N_A_239_135#_c_616_n N_A_1022_362#_c_1024_n 0.0209681f $X=5.488 $Y=2.872
+ $X2=0 $Y2=0
cc_560 N_A_239_135#_c_617_n N_A_1022_362#_M1015_g 0.00650554f $X=6.405 $Y=2.98
+ $X2=0 $Y2=0
cc_561 N_A_239_135#_c_606_n N_A_1022_362#_M1015_g 0.0038818f $X=6.13 $Y=1.96
+ $X2=0 $Y2=0
cc_562 N_A_239_135#_c_701_n N_A_1022_362#_M1015_g 0.00719214f $X=6.405 $Y=2.045
+ $X2=0 $Y2=0
cc_563 N_A_239_135#_c_619_n N_A_1022_362#_M1015_g 0.0202874f $X=6.49 $Y=2.895
+ $X2=0 $Y2=0
cc_564 N_A_239_135#_c_657_n N_A_1022_362#_c_1010_n 0.00129324f $X=6.045 $Y=1.14
+ $X2=0 $Y2=0
cc_565 N_A_239_135#_c_606_n N_A_1022_362#_c_1010_n 0.0111594f $X=6.13 $Y=1.96
+ $X2=0 $Y2=0
cc_566 N_A_239_135#_c_701_n N_A_1022_362#_c_1010_n 0.00497291f $X=6.405 $Y=2.045
+ $X2=0 $Y2=0
cc_567 N_A_239_135#_c_657_n N_A_1022_362#_c_1011_n 0.00370043f $X=6.045 $Y=1.14
+ $X2=0 $Y2=0
cc_568 N_A_239_135#_c_669_n N_A_1022_362#_c_1011_n 4.98336e-19 $X=5.505 $Y=1.055
+ $X2=0 $Y2=0
cc_569 N_A_239_135#_c_701_n N_A_878_41#_c_1227_n 0.0115322f $X=6.405 $Y=2.045
+ $X2=0 $Y2=0
cc_570 N_A_239_135#_c_617_n N_A_878_41#_c_1228_n 0.0127796f $X=6.405 $Y=2.98
+ $X2=0 $Y2=0
cc_571 N_A_239_135#_c_619_n N_A_878_41#_c_1228_n 0.0512899f $X=6.49 $Y=2.895
+ $X2=0 $Y2=0
cc_572 N_A_239_135#_c_646_n N_VPWR_M1007_d 0.0137348f $X=3.355 $Y=2.7 $X2=0
+ $Y2=0
cc_573 N_A_239_135#_c_664_n N_VPWR_M1007_d 0.00605391f $X=2.85 $Y=2.415 $X2=0
+ $Y2=0
cc_574 N_A_239_135#_M1012_g N_VPWR_c_1626_n 7.59499e-19 $X=3.485 $Y=2.355 $X2=0
+ $Y2=0
cc_575 N_A_239_135#_c_646_n N_VPWR_c_1626_n 0.00386308f $X=3.355 $Y=2.7 $X2=0
+ $Y2=0
cc_576 N_A_239_135#_c_611_n N_VPWR_c_1626_n 0.0710919f $X=4.705 $Y=2.98 $X2=0
+ $Y2=0
cc_577 N_A_239_135#_c_616_n N_VPWR_c_1626_n 0.0950512f $X=5.488 $Y=2.872 $X2=0
+ $Y2=0
cc_578 N_A_239_135#_c_617_n N_VPWR_c_1626_n 0.0109469f $X=6.405 $Y=2.98 $X2=0
+ $Y2=0
cc_579 N_A_239_135#_c_622_n N_VPWR_c_1626_n 0.0109843f $X=3.44 $Y=2.7 $X2=0
+ $Y2=0
cc_580 N_A_239_135#_c_623_n N_VPWR_c_1626_n 0.0114622f $X=4.79 $Y=2.872 $X2=0
+ $Y2=0
cc_581 N_A_239_135#_c_664_n N_VPWR_c_1629_n 0.00120838f $X=2.85 $Y=2.415 $X2=0
+ $Y2=0
cc_582 N_A_239_135#_M1011_d N_VPWR_c_1620_n 0.00233022f $X=1.27 $Y=2.095 $X2=0
+ $Y2=0
cc_583 N_A_239_135#_c_610_n N_VPWR_c_1620_n 0.00790482f $X=2.765 $Y=2.415 $X2=0
+ $Y2=0
cc_584 N_A_239_135#_c_646_n N_VPWR_c_1620_n 0.00685476f $X=3.355 $Y=2.7 $X2=0
+ $Y2=0
cc_585 N_A_239_135#_c_611_n N_VPWR_c_1620_n 0.0434094f $X=4.705 $Y=2.98 $X2=0
+ $Y2=0
cc_586 N_A_239_135#_c_616_n N_VPWR_c_1620_n 0.0524588f $X=5.488 $Y=2.872 $X2=0
+ $Y2=0
cc_587 N_A_239_135#_c_617_n N_VPWR_c_1620_n 0.00577923f $X=6.405 $Y=2.98 $X2=0
+ $Y2=0
cc_588 N_A_239_135#_c_664_n N_VPWR_c_1620_n 0.00292075f $X=2.85 $Y=2.415 $X2=0
+ $Y2=0
cc_589 N_A_239_135#_c_622_n N_VPWR_c_1620_n 0.00642982f $X=3.44 $Y=2.7 $X2=0
+ $Y2=0
cc_590 N_A_239_135#_c_623_n N_VPWR_c_1620_n 0.00657784f $X=4.79 $Y=2.872 $X2=0
+ $Y2=0
cc_591 N_A_239_135#_c_646_n N_VPWR_c_1634_n 0.0167866f $X=3.355 $Y=2.7 $X2=0
+ $Y2=0
cc_592 N_A_239_135#_c_664_n N_VPWR_c_1634_n 0.00654128f $X=2.85 $Y=2.415 $X2=0
+ $Y2=0
cc_593 N_A_239_135#_c_622_n N_VPWR_c_1634_n 0.00761521f $X=3.44 $Y=2.7 $X2=0
+ $Y2=0
cc_594 N_A_239_135#_c_610_n N_COUT_M1007_s 0.00591054f $X=2.765 $Y=2.415 $X2=0
+ $Y2=0
cc_595 N_A_239_135#_c_603_n N_COUT_c_1751_n 0.0105534f $X=1.495 $Y=1.215 $X2=0
+ $Y2=0
cc_596 N_A_239_135#_M1008_d N_COUT_c_1752_n 0.00610812f $X=1.195 $Y=0.675 $X2=0
+ $Y2=0
cc_597 N_A_239_135#_c_603_n N_COUT_c_1752_n 0.0206421f $X=1.495 $Y=1.215 $X2=0
+ $Y2=0
cc_598 N_A_239_135#_M1011_d N_COUT_c_1755_n 0.00564752f $X=1.27 $Y=2.095 $X2=0
+ $Y2=0
cc_599 N_A_239_135#_c_610_n N_COUT_c_1755_n 0.0242771f $X=2.765 $Y=2.415 $X2=0
+ $Y2=0
cc_600 N_A_239_135#_c_620_n N_COUT_c_1755_n 0.0247377f $X=1.41 $Y=2.395 $X2=0
+ $Y2=0
cc_601 N_A_239_135#_c_620_n N_COUT_c_1756_n 0.00554002f $X=1.41 $Y=2.395 $X2=0
+ $Y2=0
cc_602 N_A_239_135#_c_607_n N_COUT_c_1756_n 0.00197416f $X=1.495 $Y=2.075 $X2=0
+ $Y2=0
cc_603 N_A_239_135#_c_610_n N_COUT_c_1757_n 0.0179331f $X=2.765 $Y=2.415 $X2=0
+ $Y2=0
cc_604 N_A_239_135#_c_620_n N_COUT_c_1757_n 0.00109764f $X=1.41 $Y=2.395 $X2=0
+ $Y2=0
cc_605 N_A_239_135#_c_603_n COUT 0.0121475f $X=1.495 $Y=1.215 $X2=0 $Y2=0
cc_606 N_A_239_135#_c_611_n N_A_630_100#_M1012_d 0.00695534f $X=4.705 $Y=2.98
+ $X2=0 $Y2=0
cc_607 N_A_239_135#_M1027_g N_A_630_100#_c_1828_n 0.00737702f $X=3.075 $Y=0.82
+ $X2=0 $Y2=0
cc_608 N_A_239_135#_c_600_n N_A_630_100#_c_1828_n 0.00782804f $X=3.41 $Y=1.425
+ $X2=0 $Y2=0
cc_609 N_A_239_135#_c_602_n N_A_630_100#_c_1828_n 0.00757945f $X=3.485 $Y=1.515
+ $X2=0 $Y2=0
cc_610 N_A_239_135#_c_604_n N_A_630_100#_c_1828_n 0.00849355f $X=4.16 $Y=1.515
+ $X2=0 $Y2=0
cc_611 N_A_239_135#_c_604_n N_A_630_100#_c_1834_n 0.011944f $X=4.16 $Y=1.515
+ $X2=0 $Y2=0
cc_612 N_A_239_135#_c_605_n N_A_630_100#_c_1834_n 0.00788454f $X=3.98 $Y=1.515
+ $X2=0 $Y2=0
cc_613 N_A_239_135#_M1012_g N_A_630_100#_c_1835_n 0.019466f $X=3.485 $Y=2.355
+ $X2=0 $Y2=0
cc_614 N_A_239_135#_c_602_n N_A_630_100#_c_1835_n 0.00627423f $X=3.485 $Y=1.515
+ $X2=0 $Y2=0
cc_615 N_A_239_135#_c_604_n N_A_630_100#_c_1835_n 0.0141151f $X=4.16 $Y=1.515
+ $X2=0 $Y2=0
cc_616 N_A_239_135#_c_605_n N_A_630_100#_c_1835_n 0.00419253f $X=3.98 $Y=1.515
+ $X2=0 $Y2=0
cc_617 N_A_239_135#_c_601_n N_A_630_100#_c_1829_n 0.0109334f $X=3.15 $Y=1.425
+ $X2=0 $Y2=0
cc_618 N_A_239_135#_c_602_n N_A_630_100#_c_1830_n 0.00254133f $X=3.485 $Y=1.515
+ $X2=0 $Y2=0
cc_619 N_A_239_135#_c_604_n N_A_630_100#_c_1830_n 0.0266955f $X=4.16 $Y=1.515
+ $X2=0 $Y2=0
cc_620 N_A_239_135#_c_605_n N_A_630_100#_c_1830_n 0.00945717f $X=3.98 $Y=1.515
+ $X2=0 $Y2=0
cc_621 N_A_239_135#_c_614_n N_A_630_100#_c_1830_n 0.0193364f $X=4.705 $Y=1.895
+ $X2=0 $Y2=0
cc_622 N_A_239_135#_c_657_n N_A_630_100#_c_1830_n 0.00746439f $X=6.045 $Y=1.14
+ $X2=0 $Y2=0
cc_623 N_A_239_135#_c_606_n N_A_630_100#_c_1830_n 0.0166317f $X=6.13 $Y=1.96
+ $X2=0 $Y2=0
cc_624 N_A_239_135#_c_701_n N_A_630_100#_c_1830_n 0.0029992f $X=6.405 $Y=2.045
+ $X2=0 $Y2=0
cc_625 N_A_239_135#_c_669_n N_A_630_100#_c_1830_n 0.00367822f $X=5.505 $Y=1.055
+ $X2=0 $Y2=0
cc_626 N_A_239_135#_c_601_n N_A_630_100#_c_1831_n 0.00758452f $X=3.15 $Y=1.425
+ $X2=0 $Y2=0
cc_627 N_A_239_135#_c_606_n N_A_630_100#_c_1832_n 0.00253958f $X=6.13 $Y=1.96
+ $X2=0 $Y2=0
cc_628 N_A_239_135#_c_701_n N_A_630_100#_c_1832_n 0.0023193f $X=6.405 $Y=2.045
+ $X2=0 $Y2=0
cc_629 N_A_239_135#_c_657_n N_A_630_100#_c_1833_n 0.0105958f $X=6.045 $Y=1.14
+ $X2=0 $Y2=0
cc_630 N_A_239_135#_c_606_n N_A_630_100#_c_1833_n 0.0351819f $X=6.13 $Y=1.96
+ $X2=0 $Y2=0
cc_631 N_A_239_135#_c_701_n N_A_630_100#_c_1833_n 0.00988184f $X=6.405 $Y=2.045
+ $X2=0 $Y2=0
cc_632 N_A_239_135#_M1027_g N_VGND_c_2148_n 4.23728e-19 $X=3.075 $Y=0.82 $X2=0
+ $Y2=0
cc_633 N_A_239_135#_M1027_g N_VGND_c_2155_n 7.1892e-19 $X=3.075 $Y=0.82 $X2=0
+ $Y2=0
cc_634 N_A_814_384#_c_836_n N_A_1022_362#_M1001_g 0.00190428f $X=4.385 $Y=1.995
+ $X2=0 $Y2=0
cc_635 N_A_814_384#_M1020_g N_A_1022_362#_M1001_g 0.0180924f $X=5.845 $Y=2.315
+ $X2=0 $Y2=0
cc_636 N_A_814_384#_c_862_n N_A_1022_362#_M1001_g 0.00391384f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_637 N_A_814_384#_c_834_n N_A_1022_362#_M1001_g 0.00152435f $X=5.74 $Y=1.57
+ $X2=0 $Y2=0
cc_638 N_A_814_384#_c_822_n N_A_1022_362#_c_1022_n 0.00396018f $X=4.46 $Y=1.92
+ $X2=0 $Y2=0
cc_639 N_A_814_384#_M1020_g N_A_1022_362#_c_1022_n 0.00466275f $X=5.845 $Y=2.315
+ $X2=0 $Y2=0
cc_640 N_A_814_384#_c_862_n N_A_1022_362#_c_1022_n 7.15705e-19 $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_641 N_A_814_384#_c_834_n N_A_1022_362#_c_1022_n 0.00129254f $X=5.74 $Y=1.57
+ $X2=0 $Y2=0
cc_642 N_A_814_384#_c_822_n N_A_1022_362#_M1002_g 0.00161997f $X=4.46 $Y=1.92
+ $X2=0 $Y2=0
cc_643 N_A_814_384#_M1024_g N_A_1022_362#_M1002_g 0.0312663f $X=4.86 $Y=0.955
+ $X2=0 $Y2=0
cc_644 N_A_814_384#_c_826_n N_A_1022_362#_M1002_g 0.00737859f $X=5.645 $Y=0.19
+ $X2=0 $Y2=0
cc_645 N_A_814_384#_M1023_g N_A_1022_362#_M1002_g 0.023463f $X=5.72 $Y=0.955
+ $X2=0 $Y2=0
cc_646 N_A_814_384#_c_833_n N_A_1022_362#_M1002_g 0.0204803f $X=5.74 $Y=1.57
+ $X2=0 $Y2=0
cc_647 N_A_814_384#_c_834_n N_A_1022_362#_M1002_g 0.00305925f $X=5.74 $Y=1.57
+ $X2=0 $Y2=0
cc_648 N_A_814_384#_M1020_g N_A_1022_362#_c_1024_n 0.00881852f $X=5.845 $Y=2.315
+ $X2=0 $Y2=0
cc_649 N_A_814_384#_M1020_g N_A_1022_362#_M1015_g 0.0158818f $X=5.845 $Y=2.315
+ $X2=0 $Y2=0
cc_650 N_A_814_384#_c_841_n N_A_1022_362#_M1015_g 0.00166343f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_651 N_A_814_384#_c_841_n N_A_1022_362#_c_1009_n 0.00259406f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_652 N_A_814_384#_c_833_n N_A_1022_362#_c_1010_n 0.0131153f $X=5.74 $Y=1.57
+ $X2=0 $Y2=0
cc_653 N_A_814_384#_c_834_n N_A_1022_362#_c_1010_n 2.99611e-19 $X=5.74 $Y=1.57
+ $X2=0 $Y2=0
cc_654 N_A_814_384#_M1023_g N_A_1022_362#_c_1011_n 0.0251389f $X=5.72 $Y=0.955
+ $X2=0 $Y2=0
cc_655 N_A_814_384#_c_829_n N_A_1022_362#_c_1012_n 0.00635973f $X=9.835 $Y=1.94
+ $X2=0 $Y2=0
cc_656 N_A_814_384#_c_830_n N_A_1022_362#_c_1012_n 0.00472011f $X=10.33 $Y=1.345
+ $X2=0 $Y2=0
cc_657 N_A_814_384#_c_832_n N_A_1022_362#_c_1012_n 0.017372f $X=10.495 $Y=1.09
+ $X2=0 $Y2=0
cc_658 N_A_814_384#_c_829_n N_A_1022_362#_c_1029_n 0.00713156f $X=9.835 $Y=1.94
+ $X2=0 $Y2=0
cc_659 N_A_814_384#_c_928_p N_A_1022_362#_c_1029_n 0.0104168f $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_660 N_A_814_384#_c_928_p N_A_1022_362#_c_1013_n 4.44129e-19 $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_661 N_A_814_384#_c_841_n N_A_1022_362#_c_1013_n 0.156924f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_662 N_A_814_384#_c_841_n N_A_1022_362#_c_1014_n 0.0229758f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_663 N_A_814_384#_c_829_n N_A_1022_362#_c_1015_n 0.0140153f $X=9.835 $Y=1.94
+ $X2=0 $Y2=0
cc_664 N_A_814_384#_c_830_n N_A_1022_362#_c_1015_n 0.0160161f $X=10.33 $Y=1.345
+ $X2=0 $Y2=0
cc_665 N_A_814_384#_c_832_n N_A_1022_362#_c_1015_n 0.00815323f $X=10.495 $Y=1.09
+ $X2=0 $Y2=0
cc_666 N_A_814_384#_c_928_p N_A_1022_362#_c_1015_n 0.00791615f $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_667 N_A_814_384#_c_829_n N_A_1022_362#_c_1016_n 0.00127234f $X=9.835 $Y=1.94
+ $X2=0 $Y2=0
cc_668 N_A_814_384#_c_928_p N_A_1022_362#_c_1016_n 0.00109387f $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_669 N_A_814_384#_c_938_p N_A_1022_362#_c_1016_n 0.0296715f $X=9.36 $Y=2.035
+ $X2=0 $Y2=0
cc_670 N_A_814_384#_c_841_n N_A_1022_362#_c_1019_n 9.67352e-19 $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_671 N_A_814_384#_c_829_n N_A_1022_362#_c_1020_n 0.0221113f $X=9.835 $Y=1.94
+ $X2=0 $Y2=0
cc_672 N_A_814_384#_c_831_n N_A_1022_362#_c_1020_n 0.0134616f $X=9.92 $Y=1.345
+ $X2=0 $Y2=0
cc_673 N_A_814_384#_c_928_p N_A_1022_362#_c_1020_n 0.0207121f $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_674 N_A_814_384#_c_938_p N_A_1022_362#_c_1020_n 8.53876e-19 $X=9.36 $Y=2.035
+ $X2=0 $Y2=0
cc_675 N_A_814_384#_c_841_n N_A_878_41#_M1015_d 0.00915843f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_676 N_A_814_384#_c_928_p N_A_878_41#_M1003_g 0.00235239f $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_677 N_A_814_384#_c_841_n N_A_878_41#_M1003_g 0.00477774f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_678 N_A_814_384#_c_928_p N_A_878_41#_M1029_g 0.00212754f $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_679 N_A_814_384#_c_830_n N_A_878_41#_M1014_g 0.00783832f $X=10.33 $Y=1.345
+ $X2=0 $Y2=0
cc_680 N_A_814_384#_c_832_n N_A_878_41#_M1014_g 0.00600568f $X=10.495 $Y=1.09
+ $X2=0 $Y2=0
cc_681 N_A_814_384#_c_950_p N_A_878_41#_M1014_g 0.00737259f $X=10.495 $Y=0.935
+ $X2=0 $Y2=0
cc_682 N_A_814_384#_c_928_p N_A_878_41#_c_1212_n 5.66282e-19 $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_683 N_A_814_384#_c_829_n N_A_878_41#_c_1214_n 0.00633026f $X=9.835 $Y=1.94
+ $X2=0 $Y2=0
cc_684 N_A_814_384#_c_830_n N_A_878_41#_c_1214_n 0.00674818f $X=10.33 $Y=1.345
+ $X2=0 $Y2=0
cc_685 N_A_814_384#_c_832_n N_A_878_41#_c_1214_n 9.88721e-19 $X=10.495 $Y=1.09
+ $X2=0 $Y2=0
cc_686 N_A_814_384#_M1024_g N_A_878_41#_c_1215_n 0.0130319f $X=4.86 $Y=0.955
+ $X2=0 $Y2=0
cc_687 N_A_814_384#_c_826_n N_A_878_41#_c_1215_n 0.0100998f $X=5.645 $Y=0.19
+ $X2=0 $Y2=0
cc_688 N_A_814_384#_M1023_g N_A_878_41#_c_1215_n 0.0125866f $X=5.72 $Y=0.955
+ $X2=0 $Y2=0
cc_689 N_A_814_384#_c_841_n N_A_878_41#_c_1227_n 0.0143713f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_690 N_A_814_384#_c_841_n N_A_878_41#_c_1221_n 0.0290967f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_691 N_A_814_384#_c_841_n N_B_c_1356_n 9.50688e-19 $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_692 N_A_814_384#_c_829_n N_B_M1021_g 0.00471774f $X=9.835 $Y=1.94 $X2=0 $Y2=0
cc_693 N_A_814_384#_c_928_p N_B_M1021_g 0.0100401f $X=9.75 $Y=2.045 $X2=0 $Y2=0
cc_694 N_A_814_384#_c_829_n N_B_M1025_g 0.00250732f $X=9.835 $Y=1.94 $X2=0 $Y2=0
cc_695 N_A_814_384#_c_831_n N_B_M1025_g 0.00177717f $X=9.92 $Y=1.345 $X2=0 $Y2=0
cc_696 N_A_814_384#_c_832_n N_B_M1025_g 7.39382e-19 $X=10.495 $Y=1.09 $X2=0
+ $Y2=0
cc_697 N_A_814_384#_c_832_n N_B_M1009_g 0.00573733f $X=10.495 $Y=1.09 $X2=0
+ $Y2=0
cc_698 N_A_814_384#_c_950_p N_B_M1009_g 0.00707263f $X=10.495 $Y=0.935 $X2=0
+ $Y2=0
cc_699 N_A_814_384#_c_841_n N_B_c_1371_n 0.00763906f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_700 N_A_814_384#_c_841_n B 0.0151101f $X=9.215 $Y=2.035 $X2=0 $Y2=0
cc_701 N_A_814_384#_c_841_n N_VPWR_c_1622_n 0.00264062f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_702 N_A_814_384#_c_835_n N_VPWR_c_1626_n 0.00312768f $X=4.145 $Y=2.07 $X2=0
+ $Y2=0
cc_703 N_A_814_384#_c_835_n N_VPWR_c_1620_n 0.00589073f $X=4.145 $Y=2.07 $X2=0
+ $Y2=0
cc_704 N_A_814_384#_c_837_n N_A_630_100#_c_1834_n 0.00410288f $X=4.22 $Y=1.995
+ $X2=0 $Y2=0
cc_705 N_A_814_384#_c_837_n N_A_630_100#_c_1830_n 0.00146129f $X=4.22 $Y=1.995
+ $X2=0 $Y2=0
cc_706 N_A_814_384#_c_822_n N_A_630_100#_c_1830_n 0.00638205f $X=4.46 $Y=1.92
+ $X2=0 $Y2=0
cc_707 N_A_814_384#_c_823_n N_A_630_100#_c_1830_n 0.0100896f $X=4.785 $Y=1.46
+ $X2=0 $Y2=0
cc_708 N_A_814_384#_c_841_n N_A_630_100#_c_1830_n 0.0480473f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_709 N_A_814_384#_c_862_n N_A_630_100#_c_1830_n 0.0232331f $X=5.665 $Y=2.035
+ $X2=0 $Y2=0
cc_710 N_A_814_384#_c_833_n N_A_630_100#_c_1830_n 0.00232651f $X=5.74 $Y=1.57
+ $X2=0 $Y2=0
cc_711 N_A_814_384#_c_834_n N_A_630_100#_c_1830_n 0.0237868f $X=5.74 $Y=1.57
+ $X2=0 $Y2=0
cc_712 N_A_814_384#_c_841_n N_A_630_100#_c_1832_n 0.023676f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_713 N_A_814_384#_c_841_n N_A_630_100#_c_1833_n 4.03614e-19 $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_714 N_A_814_384#_c_841_n N_A_1741_367#_M1003_s 7.83122e-19 $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_715 N_A_814_384#_c_928_p N_A_1741_367#_c_1926_n 0.00946877f $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_716 N_A_814_384#_c_841_n N_A_1741_367#_c_1926_n 0.0312685f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_717 N_A_814_384#_c_938_p N_A_1741_367#_c_1926_n 0.00148843f $X=9.36 $Y=2.035
+ $X2=0 $Y2=0
cc_718 N_A_814_384#_M1003_d N_A_1741_367#_c_1934_n 0.00390077f $X=9.22 $Y=1.835
+ $X2=0 $Y2=0
cc_719 N_A_814_384#_c_928_p N_A_1741_367#_c_1934_n 0.0387289f $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_720 N_A_814_384#_c_841_n N_A_1741_367#_c_1934_n 0.0062855f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_721 N_A_814_384#_c_938_p N_A_1741_367#_c_1934_n 0.00779657f $X=9.36 $Y=2.035
+ $X2=0 $Y2=0
cc_722 N_A_814_384#_c_832_n N_A_1741_367#_c_1938_n 0.0070059f $X=10.495 $Y=1.09
+ $X2=0 $Y2=0
cc_723 N_A_814_384#_c_950_p N_A_1741_367#_c_1938_n 0.0301001f $X=10.495 $Y=0.935
+ $X2=0 $Y2=0
cc_724 N_A_814_384#_c_832_n N_A_1741_367#_c_1923_n 0.0020935f $X=10.495 $Y=1.09
+ $X2=0 $Y2=0
cc_725 N_A_814_384#_c_841_n N_A_1741_367#_c_1924_n 6.03531e-19 $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_726 N_A_814_384#_c_832_n N_A_1741_367#_c_1925_n 0.00946378f $X=10.495 $Y=1.09
+ $X2=0 $Y2=0
cc_727 N_A_814_384#_c_830_n N_A_1930_367#_M1025_d 0.00189457f $X=10.33 $Y=1.345
+ $X2=-0.19 $Y2=-0.245
cc_728 N_A_814_384#_c_831_n N_A_1930_367#_M1025_d 0.00309948f $X=9.92 $Y=1.345
+ $X2=-0.19 $Y2=-0.245
cc_729 N_A_814_384#_c_829_n N_A_1930_367#_M1021_d 0.00269637f $X=9.835 $Y=1.94
+ $X2=0 $Y2=0
cc_730 N_A_814_384#_c_928_p N_A_1930_367#_M1021_d 0.00643661f $X=9.75 $Y=2.045
+ $X2=0 $Y2=0
cc_731 N_A_814_384#_c_841_n N_A_1930_367#_c_2000_n 0.0206376f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_732 N_A_814_384#_c_830_n N_A_1930_367#_c_2004_n 0.014472f $X=10.33 $Y=1.345
+ $X2=0 $Y2=0
cc_733 N_A_814_384#_c_831_n N_A_1930_367#_c_2004_n 0.0111341f $X=9.92 $Y=1.345
+ $X2=0 $Y2=0
cc_734 N_A_814_384#_c_950_p N_A_1930_367#_c_2004_n 0.0301335f $X=10.495 $Y=0.935
+ $X2=0 $Y2=0
cc_735 N_A_814_384#_c_950_p N_A_1930_367#_c_2005_n 0.0197285f $X=10.495 $Y=0.935
+ $X2=0 $Y2=0
cc_736 N_A_814_384#_c_827_n N_VGND_c_2155_n 0.0218034f $X=4.935 $Y=0.19 $X2=0
+ $Y2=0
cc_737 N_A_814_384#_c_826_n N_VGND_c_2159_n 0.0227149f $X=5.645 $Y=0.19 $X2=0
+ $Y2=0
cc_738 N_A_814_384#_c_827_n N_VGND_c_2159_n 0.00589247f $X=4.935 $Y=0.19 $X2=0
+ $Y2=0
cc_739 N_A_1022_362#_c_1013_n N_A_878_41#_M1003_g 0.00915327f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_740 N_A_1022_362#_c_1016_n N_A_878_41#_M1003_g 0.00237424f $X=9.505 $Y=1.665
+ $X2=0 $Y2=0
cc_741 N_A_1022_362#_c_1020_n N_A_878_41#_M1003_g 0.00169207f $X=9.405 $Y=0.78
+ $X2=0 $Y2=0
cc_742 N_A_1022_362#_c_1020_n N_A_878_41#_M1005_g 0.0100023f $X=9.405 $Y=0.78
+ $X2=0 $Y2=0
cc_743 N_A_1022_362#_c_1012_n N_A_878_41#_M1029_g 0.00498114f $X=10.415 $Y=1.78
+ $X2=0 $Y2=0
cc_744 N_A_1022_362#_c_1029_n N_A_878_41#_M1029_g 0.00619893f $X=10.415 $Y=1.98
+ $X2=0 $Y2=0
cc_745 N_A_1022_362#_c_1015_n N_A_878_41#_M1029_g 0.00459419f $X=10.655 $Y=1.665
+ $X2=0 $Y2=0
cc_746 N_A_1022_362#_c_1017_n N_A_878_41#_M1029_g 2.28326e-19 $X=10.8 $Y=1.665
+ $X2=0 $Y2=0
cc_747 N_A_1022_362#_c_1020_n N_A_878_41#_M1014_g 9.29645e-19 $X=9.405 $Y=0.78
+ $X2=0 $Y2=0
cc_748 N_A_1022_362#_c_1016_n N_A_878_41#_c_1212_n 6.7721e-19 $X=9.505 $Y=1.665
+ $X2=0 $Y2=0
cc_749 N_A_1022_362#_c_1020_n N_A_878_41#_c_1212_n 0.00402834f $X=9.405 $Y=0.78
+ $X2=0 $Y2=0
cc_750 N_A_1022_362#_c_1012_n N_A_878_41#_c_1214_n 0.00224861f $X=10.415 $Y=1.78
+ $X2=0 $Y2=0
cc_751 N_A_1022_362#_c_1015_n N_A_878_41#_c_1214_n 0.00232278f $X=10.655
+ $Y=1.665 $X2=0 $Y2=0
cc_752 N_A_1022_362#_M1002_g N_A_878_41#_c_1215_n 0.00118849f $X=5.29 $Y=0.955
+ $X2=0 $Y2=0
cc_753 N_A_1022_362#_c_1011_n N_A_878_41#_c_1215_n 0.0132428f $X=6.387 $Y=1.185
+ $X2=0 $Y2=0
cc_754 N_A_1022_362#_c_1018_n N_A_878_41#_c_1215_n 0.00214585f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_755 N_A_1022_362#_c_1019_n N_A_878_41#_c_1215_n 0.0189956f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_756 N_A_1022_362#_M1015_g N_A_878_41#_c_1227_n 0.00103487f $X=6.51 $Y=2.315
+ $X2=0 $Y2=0
cc_757 N_A_1022_362#_c_1009_n N_A_878_41#_c_1227_n 5.43684e-19 $X=6.755 $Y=1.26
+ $X2=0 $Y2=0
cc_758 N_A_1022_362#_c_1014_n N_A_878_41#_c_1227_n 4.92868e-19 $X=7.105 $Y=1.665
+ $X2=0 $Y2=0
cc_759 N_A_1022_362#_c_1019_n N_A_878_41#_c_1227_n 0.0122756f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_760 N_A_1022_362#_M1015_g N_A_878_41#_c_1228_n 0.00653202f $X=6.51 $Y=2.315
+ $X2=0 $Y2=0
cc_761 N_A_1022_362#_c_1013_n N_A_878_41#_c_1221_n 0.00390101f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_762 N_A_1022_362#_c_1014_n N_A_878_41#_c_1221_n 9.76192e-19 $X=7.105 $Y=1.665
+ $X2=0 $Y2=0
cc_763 N_A_1022_362#_c_1019_n N_A_878_41#_c_1221_n 0.00782151f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_764 N_A_1022_362#_c_1018_n N_A_878_41#_c_1271_n 0.0017258f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_765 N_A_1022_362#_c_1019_n N_A_878_41#_c_1271_n 0.0158604f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_766 N_A_1022_362#_c_1013_n N_A_878_41#_c_1216_n 0.0195727f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_767 N_A_1022_362#_c_1014_n N_A_878_41#_c_1216_n 0.00235613f $X=7.105 $Y=1.665
+ $X2=0 $Y2=0
cc_768 N_A_1022_362#_c_1018_n N_A_878_41#_c_1216_n 0.00226257f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_769 N_A_1022_362#_c_1019_n N_A_878_41#_c_1216_n 0.0500072f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_770 N_A_1022_362#_c_1013_n N_A_878_41#_c_1217_n 0.0271897f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_771 N_A_1022_362#_c_1013_n N_A_878_41#_c_1218_n 2.24941e-19 $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_772 N_A_1022_362#_c_1018_n N_A_878_41#_c_1279_n 0.00145746f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_773 N_A_1022_362#_c_1019_n N_A_878_41#_c_1279_n 0.0134305f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_774 N_A_1022_362#_M1015_g N_B_c_1363_n 0.0150416f $X=6.51 $Y=2.315 $X2=-0.19
+ $Y2=-0.245
cc_775 N_A_1022_362#_c_1013_n N_B_c_1363_n 2.55573e-19 $X=9.215 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_776 N_A_1022_362#_c_1014_n N_B_c_1363_n 0.0011088f $X=7.105 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_777 N_A_1022_362#_c_1019_n N_B_c_1363_n 0.00208916f $X=6.92 $Y=0.83 $X2=-0.19
+ $Y2=-0.245
cc_778 N_A_1022_362#_c_1013_n N_B_c_1356_n 0.0062048f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_779 N_A_1022_362#_c_1009_n N_B_c_1357_n 0.00583005f $X=6.755 $Y=1.26 $X2=0
+ $Y2=0
cc_780 N_A_1022_362#_c_1010_n N_B_c_1357_n 0.0150416f $X=6.387 $Y=1.26 $X2=0
+ $Y2=0
cc_781 N_A_1022_362#_c_1013_n N_B_c_1357_n 8.48463e-19 $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_782 N_A_1022_362#_c_1014_n N_B_c_1357_n 3.54396e-19 $X=7.105 $Y=1.665 $X2=0
+ $Y2=0
cc_783 N_A_1022_362#_c_1019_n N_B_c_1357_n 0.00547135f $X=6.92 $Y=0.83 $X2=0
+ $Y2=0
cc_784 N_A_1022_362#_c_1018_n N_B_M1028_g 0.0114829f $X=6.92 $Y=0.83 $X2=0 $Y2=0
cc_785 N_A_1022_362#_c_1029_n N_B_M1021_g 2.1608e-19 $X=10.415 $Y=1.98 $X2=0
+ $Y2=0
cc_786 N_A_1022_362#_c_1015_n N_B_M1021_g 8.37019e-19 $X=10.655 $Y=1.665 $X2=0
+ $Y2=0
cc_787 N_A_1022_362#_c_1016_n N_B_M1021_g 3.3325e-19 $X=9.505 $Y=1.665 $X2=0
+ $Y2=0
cc_788 N_A_1022_362#_c_1020_n N_B_M1021_g 0.00175765f $X=9.405 $Y=0.78 $X2=0
+ $Y2=0
cc_789 N_A_1022_362#_c_1020_n N_B_M1025_g 0.0164737f $X=9.405 $Y=0.78 $X2=0
+ $Y2=0
cc_790 N_A_1022_362#_c_1012_n N_B_M1009_g 0.0144343f $X=10.415 $Y=1.78 $X2=0
+ $Y2=0
cc_791 N_A_1022_362#_c_1029_n N_B_M1009_g 0.00238163f $X=10.415 $Y=1.98 $X2=0
+ $Y2=0
cc_792 N_A_1022_362#_c_1015_n N_B_M1009_g 3.23708e-19 $X=10.655 $Y=1.665 $X2=0
+ $Y2=0
cc_793 N_A_1022_362#_c_1017_n N_B_M1009_g 0.00797203f $X=10.8 $Y=1.665 $X2=0
+ $Y2=0
cc_794 N_A_1022_362#_c_1013_n N_B_c_1361_n 0.00965144f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_795 N_A_1022_362#_c_1013_n N_B_c_1371_n 0.00155641f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_796 N_A_1022_362#_c_1015_n N_B_c_1362_n 0.00667625f $X=10.655 $Y=1.665 $X2=0
+ $Y2=0
cc_797 N_A_1022_362#_c_1020_n N_B_c_1362_n 0.00436369f $X=9.405 $Y=0.78 $X2=0
+ $Y2=0
cc_798 N_A_1022_362#_c_1012_n N_A_2229_269#_c_1484_n 6.26817e-19 $X=10.415
+ $Y=1.78 $X2=0 $Y2=0
cc_799 N_A_1022_362#_M1015_g N_VPWR_c_1622_n 0.00124657f $X=6.51 $Y=2.315 $X2=0
+ $Y2=0
cc_800 N_A_1022_362#_c_1025_n N_VPWR_c_1626_n 0.0317937f $X=5.26 $Y=3.15 $X2=0
+ $Y2=0
cc_801 N_A_1022_362#_c_1024_n N_VPWR_c_1620_n 0.0328469f $X=6.435 $Y=3.15 $X2=0
+ $Y2=0
cc_802 N_A_1022_362#_c_1025_n N_VPWR_c_1620_n 0.00604685f $X=5.26 $Y=3.15 $X2=0
+ $Y2=0
cc_803 N_A_1022_362#_c_1022_n N_A_630_100#_c_1830_n 0.00218039f $X=5.29 $Y=1.67
+ $X2=0 $Y2=0
cc_804 N_A_1022_362#_M1002_g N_A_630_100#_c_1830_n 0.00544428f $X=5.29 $Y=0.955
+ $X2=0 $Y2=0
cc_805 N_A_1022_362#_c_1010_n N_A_630_100#_c_1830_n 0.00597627f $X=6.387 $Y=1.26
+ $X2=0 $Y2=0
cc_806 N_A_1022_362#_M1015_g N_A_630_100#_c_1832_n 0.00110962f $X=6.51 $Y=2.315
+ $X2=0 $Y2=0
cc_807 N_A_1022_362#_c_1009_n N_A_630_100#_c_1832_n 8.82398e-19 $X=6.755 $Y=1.26
+ $X2=0 $Y2=0
cc_808 N_A_1022_362#_c_1010_n N_A_630_100#_c_1832_n 0.00440691f $X=6.387 $Y=1.26
+ $X2=0 $Y2=0
cc_809 N_A_1022_362#_c_1014_n N_A_630_100#_c_1832_n 0.021167f $X=7.105 $Y=1.665
+ $X2=0 $Y2=0
cc_810 N_A_1022_362#_c_1019_n N_A_630_100#_c_1832_n 0.00185619f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_811 N_A_1022_362#_M1015_g N_A_630_100#_c_1833_n 0.00245619f $X=6.51 $Y=2.315
+ $X2=0 $Y2=0
cc_812 N_A_1022_362#_c_1010_n N_A_630_100#_c_1833_n 0.0217446f $X=6.387 $Y=1.26
+ $X2=0 $Y2=0
cc_813 N_A_1022_362#_c_1011_n N_A_630_100#_c_1833_n 0.00193644f $X=6.387
+ $Y=1.185 $X2=0 $Y2=0
cc_814 N_A_1022_362#_c_1014_n N_A_630_100#_c_1833_n 4.22712e-19 $X=7.105
+ $Y=1.665 $X2=0 $Y2=0
cc_815 N_A_1022_362#_c_1018_n N_A_630_100#_c_1833_n 0.00406277f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_816 N_A_1022_362#_c_1019_n N_A_630_100#_c_1833_n 0.0770115f $X=6.92 $Y=0.83
+ $X2=0 $Y2=0
cc_817 N_A_1022_362#_c_1016_n N_A_1741_367#_c_1926_n 9.06535e-19 $X=9.505
+ $Y=1.665 $X2=0 $Y2=0
cc_818 N_A_1022_362#_c_1016_n N_A_1741_367#_c_1922_n 0.00114119f $X=9.505
+ $Y=1.665 $X2=0 $Y2=0
cc_819 N_A_1022_362#_c_1020_n N_A_1741_367#_c_1922_n 0.0581629f $X=9.405 $Y=0.78
+ $X2=0 $Y2=0
cc_820 N_A_1022_362#_M1029_d N_A_1741_367#_c_1934_n 0.00505597f $X=10.275
+ $Y=1.835 $X2=0 $Y2=0
cc_821 N_A_1022_362#_c_1012_n N_A_1741_367#_c_1934_n 0.00280575f $X=10.415
+ $Y=1.78 $X2=0 $Y2=0
cc_822 N_A_1022_362#_c_1029_n N_A_1741_367#_c_1934_n 0.0199532f $X=10.415
+ $Y=1.98 $X2=0 $Y2=0
cc_823 N_A_1022_362#_c_1015_n N_A_1741_367#_c_1934_n 0.0116526f $X=10.655
+ $Y=1.665 $X2=0 $Y2=0
cc_824 N_A_1022_362#_c_1017_n N_A_1741_367#_c_1934_n 5.70787e-19 $X=10.8
+ $Y=1.665 $X2=0 $Y2=0
cc_825 N_A_1022_362#_c_1012_n N_A_1741_367#_c_1923_n 0.0145454f $X=10.415
+ $Y=1.78 $X2=0 $Y2=0
cc_826 N_A_1022_362#_c_1029_n N_A_1741_367#_c_1923_n 0.00195321f $X=10.415
+ $Y=1.98 $X2=0 $Y2=0
cc_827 N_A_1022_362#_c_1017_n N_A_1741_367#_c_1923_n 0.00742586f $X=10.8
+ $Y=1.665 $X2=0 $Y2=0
cc_828 N_A_1022_362#_c_1013_n N_A_1741_367#_c_1924_n 0.0316461f $X=9.215
+ $Y=1.665 $X2=0 $Y2=0
cc_829 N_A_1022_362#_c_1016_n N_A_1741_367#_c_1924_n 6.47585e-19 $X=9.505
+ $Y=1.665 $X2=0 $Y2=0
cc_830 N_A_1022_362#_c_1012_n N_A_1741_367#_c_1956_n 0.00785169f $X=10.415
+ $Y=1.78 $X2=0 $Y2=0
cc_831 N_A_1022_362#_c_1017_n N_A_1741_367#_c_1956_n 0.00214633f $X=10.8
+ $Y=1.665 $X2=0 $Y2=0
cc_832 N_A_1022_362#_c_1012_n N_A_1741_367#_c_1925_n 0.00251257f $X=10.415
+ $Y=1.78 $X2=0 $Y2=0
cc_833 N_A_1022_362#_c_1017_n N_A_1741_367#_c_1925_n 0.00128645f $X=10.8
+ $Y=1.665 $X2=0 $Y2=0
cc_834 N_A_1022_362#_c_1013_n N_A_1930_367#_c_2000_n 0.0136751f $X=9.215
+ $Y=1.665 $X2=0 $Y2=0
cc_835 N_A_1022_362#_c_1020_n N_A_1930_367#_c_2002_n 0.0244976f $X=9.405 $Y=0.78
+ $X2=0 $Y2=0
cc_836 N_A_1022_362#_c_1015_n N_A_1930_367#_c_2004_n 0.00103402f $X=10.655
+ $Y=1.665 $X2=0 $Y2=0
cc_837 N_A_1022_362#_c_1020_n N_A_1930_367#_c_2004_n 0.0301493f $X=9.405 $Y=0.78
+ $X2=0 $Y2=0
cc_838 N_A_1022_362#_c_1013_n N_A_1930_367#_c_2008_n 0.00910951f $X=9.215
+ $Y=1.665 $X2=0 $Y2=0
cc_839 N_A_1022_362#_c_1011_n N_VGND_c_2155_n 7.7537e-19 $X=6.387 $Y=1.185 $X2=0
+ $Y2=0
cc_840 N_A_878_41#_c_1221_n N_B_c_1363_n 0.0128837f $X=7.265 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_841 N_A_878_41#_c_1216_n N_B_c_1363_n 0.00488f $X=7.35 $Y=1.96 $X2=-0.19
+ $Y2=-0.245
cc_842 N_A_878_41#_c_1221_n N_B_c_1356_n 0.00125146f $X=7.265 $Y=2.045 $X2=0
+ $Y2=0
cc_843 N_A_878_41#_c_1216_n N_B_c_1356_n 0.0150931f $X=7.35 $Y=1.96 $X2=0 $Y2=0
cc_844 N_A_878_41#_c_1206_n N_B_M1028_g 0.0211829f $X=8.365 $Y=0.18 $X2=0 $Y2=0
cc_845 N_A_878_41#_c_1216_n N_B_M1028_g 0.0158884f $X=7.35 $Y=1.96 $X2=0 $Y2=0
cc_846 N_A_878_41#_c_1217_n N_B_M1028_g 0.0140642f $X=8.045 $Y=0.975 $X2=0 $Y2=0
cc_847 N_A_878_41#_c_1288_p N_B_M1028_g 8.16773e-19 $X=8.2 $Y=0.555 $X2=0 $Y2=0
cc_848 N_A_878_41#_M1003_g N_B_c_1366_n 0.00737859f $X=9.145 $Y=2.255 $X2=0
+ $Y2=0
cc_849 N_A_878_41#_M1029_g N_B_M1021_g 0.0247445f $X=10.2 $Y=2.255 $X2=0 $Y2=0
cc_850 N_A_878_41#_M1003_g N_B_M1025_g 0.00177801f $X=9.145 $Y=2.255 $X2=0 $Y2=0
cc_851 N_A_878_41#_M1005_g N_B_M1025_g 0.0177412f $X=9.19 $Y=0.945 $X2=0 $Y2=0
cc_852 N_A_878_41#_c_1209_n N_B_M1025_g 0.00737233f $X=10.205 $Y=0.18 $X2=0
+ $Y2=0
cc_853 N_A_878_41#_M1014_g N_B_M1025_g 0.0131606f $X=10.28 $Y=0.915 $X2=0 $Y2=0
cc_854 N_A_878_41#_c_1214_n N_B_M1025_g 0.00448984f $X=10.28 $Y=1.42 $X2=0 $Y2=0
cc_855 N_A_878_41#_M1029_g N_B_c_1368_n 0.00754303f $X=10.2 $Y=2.255 $X2=0 $Y2=0
cc_856 N_A_878_41#_M1029_g N_B_M1009_g 0.03796f $X=10.2 $Y=2.255 $X2=0 $Y2=0
cc_857 N_A_878_41#_M1014_g N_B_M1009_g 0.0287121f $X=10.28 $Y=0.915 $X2=0 $Y2=0
cc_858 N_A_878_41#_c_1217_n N_B_c_1361_n 0.00552968f $X=8.045 $Y=0.975 $X2=0
+ $Y2=0
cc_859 N_A_878_41#_c_1221_n N_B_c_1371_n 0.0032376f $X=7.265 $Y=2.045 $X2=0
+ $Y2=0
cc_860 N_A_878_41#_c_1216_n N_B_c_1371_n 0.00479148f $X=7.35 $Y=1.96 $X2=0 $Y2=0
cc_861 N_A_878_41#_M1003_g N_B_c_1362_n 0.0387123f $X=9.145 $Y=2.255 $X2=0 $Y2=0
cc_862 N_A_878_41#_M1029_g N_B_c_1362_n 0.00448984f $X=10.2 $Y=2.255 $X2=0 $Y2=0
cc_863 N_A_878_41#_c_1221_n N_VPWR_M1022_d 0.00416066f $X=7.265 $Y=2.045 $X2=0
+ $Y2=0
cc_864 N_A_878_41#_c_1216_n N_VPWR_M1022_d 0.00172155f $X=7.35 $Y=1.96 $X2=0
+ $Y2=0
cc_865 N_A_878_41#_c_1221_n N_VPWR_c_1622_n 0.0201549f $X=7.265 $Y=2.045 $X2=0
+ $Y2=0
cc_866 N_A_878_41#_c_1228_n N_VPWR_c_1626_n 0.0110663f $X=6.84 $Y=2.9 $X2=0
+ $Y2=0
cc_867 N_A_878_41#_M1015_d N_VPWR_c_1620_n 0.00633253f $X=6.585 $Y=1.895 $X2=0
+ $Y2=0
cc_868 N_A_878_41#_c_1228_n N_VPWR_c_1620_n 0.006495f $X=6.84 $Y=2.9 $X2=0 $Y2=0
cc_869 N_A_878_41#_c_1215_n N_A_630_100#_c_1833_n 0.0131312f $X=7.265 $Y=0.35
+ $X2=0 $Y2=0
cc_870 N_A_878_41#_M1003_g N_A_1741_367#_c_1926_n 0.0124225f $X=9.145 $Y=2.255
+ $X2=0 $Y2=0
cc_871 N_A_878_41#_M1005_g N_A_1741_367#_c_1922_n 0.00262489f $X=9.19 $Y=0.945
+ $X2=0 $Y2=0
cc_872 N_A_878_41#_c_1212_n N_A_1741_367#_c_1922_n 0.00441866f $X=9.167 $Y=1.525
+ $X2=0 $Y2=0
cc_873 N_A_878_41#_M1003_g N_A_1741_367#_c_1934_n 0.0117087f $X=9.145 $Y=2.255
+ $X2=0 $Y2=0
cc_874 N_A_878_41#_M1029_g N_A_1741_367#_c_1934_n 0.0129916f $X=10.2 $Y=2.255
+ $X2=0 $Y2=0
cc_875 N_A_878_41#_M1029_g N_A_1741_367#_c_1965_n 7.85155e-19 $X=10.2 $Y=2.255
+ $X2=0 $Y2=0
cc_876 N_A_878_41#_M1003_g N_A_1741_367#_c_1924_n 0.00441866f $X=9.145 $Y=2.255
+ $X2=0 $Y2=0
cc_877 N_A_878_41#_M1003_g N_A_1741_367#_c_1929_n 0.00418945f $X=9.145 $Y=2.255
+ $X2=0 $Y2=0
cc_878 N_A_878_41#_M1003_g N_A_1930_367#_c_2000_n 0.00271658f $X=9.145 $Y=2.255
+ $X2=0 $Y2=0
cc_879 N_A_878_41#_M1003_g N_A_1930_367#_c_2011_n 0.00157534f $X=9.145 $Y=2.255
+ $X2=0 $Y2=0
cc_880 N_A_878_41#_M1005_g N_A_1930_367#_c_2001_n 0.00572097f $X=9.19 $Y=0.945
+ $X2=0 $Y2=0
cc_881 N_A_878_41#_c_1217_n N_A_1930_367#_c_2001_n 0.0130075f $X=8.045 $Y=0.975
+ $X2=0 $Y2=0
cc_882 N_A_878_41#_c_1288_p N_A_1930_367#_c_2001_n 0.032567f $X=8.2 $Y=0.555
+ $X2=0 $Y2=0
cc_883 N_A_878_41#_c_1218_n N_A_1930_367#_c_2001_n 0.0140003f $X=8.2 $Y=0.555
+ $X2=0 $Y2=0
cc_884 N_A_878_41#_c_1205_n N_A_1930_367#_c_2002_n 0.00735352f $X=9.115 $Y=0.18
+ $X2=0 $Y2=0
cc_885 N_A_878_41#_M1005_g N_A_1930_367#_c_2002_n 0.017572f $X=9.19 $Y=0.945
+ $X2=0 $Y2=0
cc_886 N_A_878_41#_c_1209_n N_A_1930_367#_c_2002_n 0.00762504f $X=10.205 $Y=0.18
+ $X2=0 $Y2=0
cc_887 N_A_878_41#_c_1205_n N_A_1930_367#_c_2003_n 0.00418768f $X=9.115 $Y=0.18
+ $X2=0 $Y2=0
cc_888 N_A_878_41#_c_1288_p N_A_1930_367#_c_2003_n 0.00362359f $X=8.2 $Y=0.555
+ $X2=0 $Y2=0
cc_889 N_A_878_41#_c_1218_n N_A_1930_367#_c_2003_n 0.00480353f $X=8.2 $Y=0.555
+ $X2=0 $Y2=0
cc_890 N_A_878_41#_M1005_g N_A_1930_367#_c_2004_n 0.00174189f $X=9.19 $Y=0.945
+ $X2=0 $Y2=0
cc_891 N_A_878_41#_M1014_g N_A_1930_367#_c_2004_n 0.0105865f $X=10.28 $Y=0.915
+ $X2=0 $Y2=0
cc_892 N_A_878_41#_M1029_g N_A_1930_367#_c_2013_n 0.00719459f $X=10.2 $Y=2.255
+ $X2=0 $Y2=0
cc_893 N_A_878_41#_M1014_g N_A_1930_367#_c_2005_n 0.0177374f $X=10.28 $Y=0.915
+ $X2=0 $Y2=0
cc_894 N_A_878_41#_c_1217_n N_A_1930_367#_c_2008_n 0.00183871f $X=8.045 $Y=0.975
+ $X2=0 $Y2=0
cc_895 N_A_878_41#_c_1218_n N_A_1930_367#_c_2008_n 3.77083e-19 $X=8.2 $Y=0.555
+ $X2=0 $Y2=0
cc_896 N_A_878_41#_M1029_g N_A_1930_367#_c_2016_n 3.8325e-19 $X=10.2 $Y=2.255
+ $X2=0 $Y2=0
cc_897 N_A_878_41#_c_1209_n N_A_1930_367#_c_2009_n 0.00812903f $X=10.205 $Y=0.18
+ $X2=0 $Y2=0
cc_898 N_A_878_41#_c_1217_n N_VGND_M1028_d 0.00703782f $X=8.045 $Y=0.975 $X2=0
+ $Y2=0
cc_899 N_A_878_41#_c_1206_n N_VGND_c_2149_n 0.00729525f $X=8.365 $Y=0.18 $X2=0
+ $Y2=0
cc_900 N_A_878_41#_c_1217_n N_VGND_c_2149_n 0.0147641f $X=8.045 $Y=0.975 $X2=0
+ $Y2=0
cc_901 N_A_878_41#_c_1288_p N_VGND_c_2149_n 0.0231873f $X=8.2 $Y=0.555 $X2=0
+ $Y2=0
cc_902 N_A_878_41#_c_1215_n N_VGND_c_2155_n 0.174285f $X=7.265 $Y=0.35 $X2=0
+ $Y2=0
cc_903 N_A_878_41#_c_1344_p N_VGND_c_2155_n 0.0111659f $X=7.35 $Y=0.435 $X2=0
+ $Y2=0
cc_904 N_A_878_41#_c_1206_n N_VGND_c_2157_n 0.0540191f $X=8.365 $Y=0.18 $X2=0
+ $Y2=0
cc_905 N_A_878_41#_c_1288_p N_VGND_c_2157_n 0.0111366f $X=8.2 $Y=0.555 $X2=0
+ $Y2=0
cc_906 N_A_878_41#_M1024_s N_VGND_c_2159_n 0.00258405f $X=4.39 $Y=0.205 $X2=0
+ $Y2=0
cc_907 N_A_878_41#_M1028_s N_VGND_c_2159_n 0.0041999f $X=7.205 $Y=0.235 $X2=0
+ $Y2=0
cc_908 N_A_878_41#_c_1205_n N_VGND_c_2159_n 0.0236443f $X=9.115 $Y=0.18 $X2=0
+ $Y2=0
cc_909 N_A_878_41#_c_1206_n N_VGND_c_2159_n 0.0101832f $X=8.365 $Y=0.18 $X2=0
+ $Y2=0
cc_910 N_A_878_41#_c_1209_n N_VGND_c_2159_n 0.028166f $X=10.205 $Y=0.18 $X2=0
+ $Y2=0
cc_911 N_A_878_41#_c_1213_n N_VGND_c_2159_n 0.00371014f $X=9.19 $Y=0.18 $X2=0
+ $Y2=0
cc_912 N_A_878_41#_c_1215_n N_VGND_c_2159_n 0.103927f $X=7.265 $Y=0.35 $X2=0
+ $Y2=0
cc_913 N_A_878_41#_c_1344_p N_VGND_c_2159_n 0.00656694f $X=7.35 $Y=0.435 $X2=0
+ $Y2=0
cc_914 N_A_878_41#_c_1288_p N_VGND_c_2159_n 0.00973671f $X=8.2 $Y=0.555 $X2=0
+ $Y2=0
cc_915 N_B_c_1368_n N_A_2229_269#_M1000_g 0.0271939f $X=10.635 $Y=3.12 $X2=0
+ $Y2=0
cc_916 N_B_M1009_g N_A_2229_269#_c_1483_n 0.0165796f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_917 N_B_M1009_g N_A_2229_269#_c_1484_n 0.0271939f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_918 N_B_c_1363_n N_VPWR_c_1622_n 0.0160637f $X=7.055 $Y=1.725 $X2=0 $Y2=0
cc_919 N_B_c_1356_n N_VPWR_c_1622_n 6.68236e-19 $X=7.49 $Y=1.65 $X2=0 $Y2=0
cc_920 N_B_c_1372_n N_VPWR_c_1622_n 0.00575967f $X=7.87 $Y=2.795 $X2=0 $Y2=0
cc_921 B N_VPWR_c_1622_n 0.0364075f $X=7.835 $Y=2.32 $X2=0 $Y2=0
cc_922 N_B_c_1376_n N_VPWR_c_1622_n 0.00606454f $X=7.87 $Y=2.455 $X2=0 $Y2=0
cc_923 N_B_c_1363_n N_VPWR_c_1626_n 0.00486043f $X=7.055 $Y=1.725 $X2=0 $Y2=0
cc_924 N_B_c_1372_n N_VPWR_c_1630_n 0.066044f $X=7.87 $Y=2.795 $X2=0 $Y2=0
cc_925 B N_VPWR_c_1630_n 0.0125839f $X=7.835 $Y=2.32 $X2=0 $Y2=0
cc_926 N_B_c_1363_n N_VPWR_c_1620_n 0.00847851f $X=7.055 $Y=1.725 $X2=0 $Y2=0
cc_927 N_B_c_1366_n N_VPWR_c_1620_n 0.0446754f $X=9.5 $Y=3.12 $X2=0 $Y2=0
cc_928 N_B_c_1368_n N_VPWR_c_1620_n 0.0291371f $X=10.635 $Y=3.12 $X2=0 $Y2=0
cc_929 N_B_c_1372_n N_VPWR_c_1620_n 0.00568355f $X=7.87 $Y=2.795 $X2=0 $Y2=0
cc_930 N_B_c_1374_n N_VPWR_c_1620_n 0.00375312f $X=9.575 $Y=3.12 $X2=0 $Y2=0
cc_931 B N_VPWR_c_1620_n 0.0110834f $X=7.835 $Y=2.32 $X2=0 $Y2=0
cc_932 N_B_c_1357_n N_A_630_100#_c_1833_n 2.56268e-19 $X=7.13 $Y=1.65 $X2=0
+ $Y2=0
cc_933 N_B_M1021_g N_A_1741_367#_c_1934_n 0.0124424f $X=9.575 $Y=2.255 $X2=0
+ $Y2=0
cc_934 N_B_c_1368_n N_A_1741_367#_c_1934_n 0.00108508f $X=10.635 $Y=3.12 $X2=0
+ $Y2=0
cc_935 N_B_M1009_g N_A_1741_367#_c_1934_n 0.0109139f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_936 N_B_M1009_g N_A_1741_367#_c_1965_n 0.00376316f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_937 N_B_M1009_g N_A_1741_367#_c_1938_n 0.00512748f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_938 N_B_M1009_g N_A_1741_367#_c_1923_n 0.00406775f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_939 N_B_M1009_g N_A_1741_367#_c_1956_n 0.00323552f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_940 N_B_M1009_g N_A_1741_367#_c_1925_n 0.00180295f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_941 N_B_M1028_g N_A_1930_367#_c_2000_n 0.00328363f $X=7.565 $Y=0.655 $X2=0
+ $Y2=0
cc_942 N_B_c_1361_n N_A_1930_367#_c_2000_n 0.0154482f $X=7.78 $Y=1.65 $X2=0
+ $Y2=0
cc_943 B N_A_1930_367#_c_2000_n 0.0287088f $X=7.835 $Y=2.32 $X2=0 $Y2=0
cc_944 N_B_c_1376_n N_A_1930_367#_c_2000_n 0.0119376f $X=7.87 $Y=2.455 $X2=0
+ $Y2=0
cc_945 N_B_c_1366_n N_A_1930_367#_c_2011_n 0.0192625f $X=9.5 $Y=3.12 $X2=0 $Y2=0
cc_946 N_B_M1021_g N_A_1930_367#_c_2011_n 0.0136717f $X=9.575 $Y=2.255 $X2=0
+ $Y2=0
cc_947 N_B_c_1366_n N_A_1930_367#_c_2012_n 0.00432079f $X=9.5 $Y=3.12 $X2=0
+ $Y2=0
cc_948 N_B_c_1372_n N_A_1930_367#_c_2012_n 0.0048782f $X=7.87 $Y=2.795 $X2=0
+ $Y2=0
cc_949 B N_A_1930_367#_c_2012_n 0.00469811f $X=7.835 $Y=2.32 $X2=0 $Y2=0
cc_950 N_B_M1025_g N_A_1930_367#_c_2002_n 0.00331137f $X=9.62 $Y=0.945 $X2=0
+ $Y2=0
cc_951 N_B_M1025_g N_A_1930_367#_c_2004_n 0.00818044f $X=9.62 $Y=0.945 $X2=0
+ $Y2=0
cc_952 N_B_c_1368_n N_A_1930_367#_c_2013_n 0.00786694f $X=10.635 $Y=3.12 $X2=0
+ $Y2=0
cc_953 N_B_M1009_g N_A_1930_367#_c_2013_n 0.0122597f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_954 N_B_M1009_g N_A_1930_367#_c_2005_n 0.00684395f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_955 N_B_M1009_g N_A_1930_367#_c_2066_n 7.51949e-19 $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_956 N_B_M1028_g N_A_1930_367#_c_2008_n 0.00369835f $X=7.565 $Y=0.655 $X2=0
+ $Y2=0
cc_957 N_B_M1021_g N_A_1930_367#_c_2016_n 0.00757667f $X=9.575 $Y=2.255 $X2=0
+ $Y2=0
cc_958 N_B_c_1368_n N_A_1930_367#_c_2016_n 0.00809934f $X=10.635 $Y=3.12 $X2=0
+ $Y2=0
cc_959 N_B_M1009_g N_A_1930_367#_c_2016_n 0.00494646f $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_960 N_B_M1009_g N_A_1930_367#_c_2071_n 8.89287e-19 $X=10.71 $Y=0.915 $X2=0
+ $Y2=0
cc_961 N_B_M1028_g N_VGND_c_2149_n 0.0119537f $X=7.565 $Y=0.655 $X2=0 $Y2=0
cc_962 N_B_M1028_g N_VGND_c_2155_n 0.00486043f $X=7.565 $Y=0.655 $X2=0 $Y2=0
cc_963 N_B_M1028_g N_VGND_c_2159_n 0.00954696f $X=7.565 $Y=0.655 $X2=0 $Y2=0
cc_964 N_A_2229_269#_c_1485_n N_A_M1026_g 0.0162628f $X=12.995 $Y=1.285 $X2=0
+ $Y2=0
cc_965 N_A_2229_269#_c_1486_n N_A_M1026_g 0.00107794f $X=13.16 $Y=0.505 $X2=0
+ $Y2=0
cc_966 N_A_2229_269#_c_1487_n N_A_M1026_g 8.70136e-19 $X=13.16 $Y=2.19 $X2=0
+ $Y2=0
cc_967 N_A_2229_269#_c_1488_n N_A_M1026_g 0.00112688f $X=11.61 $Y=1.285 $X2=0
+ $Y2=0
cc_968 N_A_2229_269#_c_1489_n N_A_M1026_g 0.00404387f $X=11.61 $Y=1.51 $X2=0
+ $Y2=0
cc_969 N_A_2229_269#_c_1485_n N_A_c_1553_n 0.0033869f $X=12.995 $Y=1.285 $X2=0
+ $Y2=0
cc_970 N_A_2229_269#_c_1485_n N_A_M1010_g 0.0149371f $X=12.995 $Y=1.285 $X2=0
+ $Y2=0
cc_971 N_A_2229_269#_c_1486_n N_A_M1010_g 0.0149299f $X=13.16 $Y=0.505 $X2=0
+ $Y2=0
cc_972 N_A_2229_269#_c_1487_n N_A_M1010_g 0.00686217f $X=13.16 $Y=2.19 $X2=0
+ $Y2=0
cc_973 N_A_2229_269#_c_1490_n N_A_M1010_g 0.00383478f $X=13.16 $Y=1.285 $X2=0
+ $Y2=0
cc_974 N_A_2229_269#_c_1487_n N_A_M1016_g 0.0239104f $X=13.16 $Y=2.19 $X2=0
+ $Y2=0
cc_975 N_A_2229_269#_c_1487_n N_A_c_1555_n 0.00674624f $X=13.16 $Y=2.19 $X2=0
+ $Y2=0
cc_976 N_A_2229_269#_c_1485_n N_A_c_1556_n 0.00400978f $X=12.995 $Y=1.285 $X2=0
+ $Y2=0
cc_977 N_A_2229_269#_c_1487_n N_A_c_1556_n 0.00133861f $X=13.16 $Y=2.19 $X2=0
+ $Y2=0
cc_978 N_A_2229_269#_c_1489_n N_A_c_1556_n 0.00268479f $X=11.61 $Y=1.51 $X2=0
+ $Y2=0
cc_979 N_A_2229_269#_c_1485_n N_A_c_1557_n 0.0334708f $X=12.995 $Y=1.285 $X2=0
+ $Y2=0
cc_980 N_A_2229_269#_c_1487_n N_A_c_1557_n 0.0125655f $X=13.16 $Y=2.19 $X2=0
+ $Y2=0
cc_981 N_A_2229_269#_c_1488_n N_A_c_1557_n 0.00591902f $X=11.61 $Y=1.285 $X2=0
+ $Y2=0
cc_982 N_A_2229_269#_c_1489_n N_A_c_1557_n 0.00113556f $X=11.61 $Y=1.51 $X2=0
+ $Y2=0
cc_983 N_A_2229_269#_M1000_g N_VPWR_c_1623_n 0.00979591f $X=11.22 $Y=2.465 $X2=0
+ $Y2=0
cc_984 N_A_2229_269#_c_1487_n N_VPWR_c_1625_n 0.0367071f $X=13.16 $Y=2.19 $X2=0
+ $Y2=0
cc_985 N_A_2229_269#_M1000_g N_VPWR_c_1630_n 0.00401687f $X=11.22 $Y=2.465 $X2=0
+ $Y2=0
cc_986 N_A_2229_269#_c_1487_n N_VPWR_c_1631_n 0.0220321f $X=13.16 $Y=2.19 $X2=0
+ $Y2=0
cc_987 N_A_2229_269#_M1000_g N_VPWR_c_1620_n 0.00754288f $X=11.22 $Y=2.465 $X2=0
+ $Y2=0
cc_988 N_A_2229_269#_c_1487_n N_VPWR_c_1620_n 0.0125808f $X=13.16 $Y=2.19 $X2=0
+ $Y2=0
cc_989 N_A_2229_269#_M1000_g N_A_1741_367#_c_1923_n 0.0158034f $X=11.22 $Y=2.465
+ $X2=0 $Y2=0
cc_990 N_A_2229_269#_c_1484_n N_A_1741_367#_c_1923_n 0.0100028f $X=11.237
+ $Y=1.51 $X2=0 $Y2=0
cc_991 N_A_2229_269#_c_1488_n N_A_1741_367#_c_1923_n 0.0204382f $X=11.61
+ $Y=1.285 $X2=0 $Y2=0
cc_992 N_A_2229_269#_M1000_g N_A_1741_367#_c_1956_n 0.0148063f $X=11.22 $Y=2.465
+ $X2=0 $Y2=0
cc_993 N_A_2229_269#_c_1483_n N_A_1741_367#_c_1925_n 0.00775407f $X=11.255
+ $Y=1.345 $X2=0 $Y2=0
cc_994 N_A_2229_269#_c_1484_n N_A_1741_367#_c_1925_n 0.00187875f $X=11.237
+ $Y=1.51 $X2=0 $Y2=0
cc_995 N_A_2229_269#_c_1488_n N_A_1741_367#_c_1925_n 0.0127624f $X=11.61
+ $Y=1.285 $X2=0 $Y2=0
cc_996 N_A_2229_269#_M1000_g N_A_1930_367#_c_2013_n 0.010424f $X=11.22 $Y=2.465
+ $X2=0 $Y2=0
cc_997 N_A_2229_269#_c_1483_n N_A_1930_367#_c_2005_n 0.0154174f $X=11.255
+ $Y=1.345 $X2=0 $Y2=0
cc_998 N_A_2229_269#_c_1483_n N_A_1930_367#_c_2066_n 0.0135832f $X=11.255
+ $Y=1.345 $X2=0 $Y2=0
cc_999 N_A_2229_269#_M1000_g N_A_1930_367#_c_2014_n 9.20342e-19 $X=11.22
+ $Y=2.465 $X2=0 $Y2=0
cc_1000 N_A_2229_269#_c_1485_n N_A_1930_367#_c_2006_n 0.0522586f $X=12.995
+ $Y=1.285 $X2=0 $Y2=0
cc_1001 N_A_2229_269#_c_1488_n N_A_1930_367#_c_2006_n 0.0226067f $X=11.61
+ $Y=1.285 $X2=0 $Y2=0
cc_1002 N_A_2229_269#_c_1489_n N_A_1930_367#_c_2006_n 0.00146787f $X=11.61
+ $Y=1.51 $X2=0 $Y2=0
cc_1003 N_A_2229_269#_c_1483_n N_A_1930_367#_c_2079_n 0.00715454f $X=11.255
+ $Y=1.345 $X2=0 $Y2=0
cc_1004 N_A_2229_269#_c_1488_n N_A_1930_367#_c_2079_n 0.00243969f $X=11.61
+ $Y=1.285 $X2=0 $Y2=0
cc_1005 N_A_2229_269#_c_1489_n N_A_1930_367#_c_2079_n 0.00334584f $X=11.61
+ $Y=1.51 $X2=0 $Y2=0
cc_1006 N_A_2229_269#_M1000_g N_A_1930_367#_c_2071_n 0.0114358f $X=11.22
+ $Y=2.465 $X2=0 $Y2=0
cc_1007 N_A_2229_269#_c_1485_n N_VGND_M1019_d 0.00129074f $X=12.995 $Y=1.285
+ $X2=0 $Y2=0
cc_1008 N_A_2229_269#_c_1488_n N_VGND_M1019_d 0.00407244f $X=11.61 $Y=1.285
+ $X2=0 $Y2=0
cc_1009 N_A_2229_269#_c_1483_n N_VGND_c_2150_n 0.00209411f $X=11.255 $Y=1.345
+ $X2=0 $Y2=0
cc_1010 N_A_2229_269#_c_1485_n N_VGND_c_2152_n 0.0136256f $X=12.995 $Y=1.285
+ $X2=0 $Y2=0
cc_1011 N_A_2229_269#_c_1486_n N_VGND_c_2152_n 0.0257452f $X=13.16 $Y=0.505
+ $X2=0 $Y2=0
cc_1012 N_A_2229_269#_c_1483_n N_VGND_c_2157_n 0.00336933f $X=11.255 $Y=1.345
+ $X2=0 $Y2=0
cc_1013 N_A_2229_269#_c_1486_n N_VGND_c_2158_n 0.0151738f $X=13.16 $Y=0.505
+ $X2=0 $Y2=0
cc_1014 N_A_2229_269#_c_1483_n N_VGND_c_2159_n 0.00448211f $X=11.255 $Y=1.345
+ $X2=0 $Y2=0
cc_1015 N_A_2229_269#_c_1486_n N_VGND_c_2159_n 0.0120712f $X=13.16 $Y=0.505
+ $X2=0 $Y2=0
cc_1016 N_A_M1030_g N_VPWR_c_1623_n 0.00210814f $X=12.515 $Y=2.545 $X2=0 $Y2=0
cc_1017 N_A_M1030_g N_VPWR_c_1624_n 0.00502664f $X=12.515 $Y=2.545 $X2=0 $Y2=0
cc_1018 N_A_M1030_g N_VPWR_c_1625_n 0.00364626f $X=12.515 $Y=2.545 $X2=0 $Y2=0
cc_1019 N_A_c_1553_n N_VPWR_c_1625_n 0.00335914f $X=12.87 $Y=1.625 $X2=0 $Y2=0
cc_1020 N_A_M1016_g N_VPWR_c_1625_n 0.00364626f $X=12.945 $Y=2.545 $X2=0 $Y2=0
cc_1021 N_A_M1016_g N_VPWR_c_1631_n 0.00502664f $X=12.945 $Y=2.545 $X2=0 $Y2=0
cc_1022 N_A_M1030_g N_VPWR_c_1620_n 0.0103182f $X=12.515 $Y=2.545 $X2=0 $Y2=0
cc_1023 N_A_M1016_g N_VPWR_c_1620_n 0.0100768f $X=12.945 $Y=2.545 $X2=0 $Y2=0
cc_1024 N_A_c_1557_n N_A_1930_367#_c_2014_n 3.03247e-19 $X=12.425 $Y=1.715 $X2=0
+ $Y2=0
cc_1025 N_A_M1026_g N_A_1930_367#_c_2006_n 0.00258257f $X=12.515 $Y=0.68 $X2=0
+ $Y2=0
cc_1026 N_A_M1026_g N_A_1930_367#_c_2007_n 0.00587648f $X=12.515 $Y=0.68 $X2=0
+ $Y2=0
cc_1027 N_A_M1030_g N_A_1930_367#_c_2015_n 0.00678878f $X=12.515 $Y=2.545 $X2=0
+ $Y2=0
cc_1028 N_A_c_1556_n N_A_1930_367#_c_2015_n 0.00399301f $X=12.425 $Y=1.625 $X2=0
+ $Y2=0
cc_1029 N_A_c_1557_n N_A_1930_367#_c_2015_n 0.0239036f $X=12.425 $Y=1.715 $X2=0
+ $Y2=0
cc_1030 N_A_M1030_g N_A_1930_367#_c_2017_n 0.0109048f $X=12.515 $Y=2.545 $X2=0
+ $Y2=0
cc_1031 N_A_M1026_g N_VGND_c_2150_n 0.00312582f $X=12.515 $Y=0.68 $X2=0 $Y2=0
cc_1032 N_A_M1026_g N_VGND_c_2151_n 0.00441827f $X=12.515 $Y=0.68 $X2=0 $Y2=0
cc_1033 N_A_M1026_g N_VGND_c_2152_n 0.00285146f $X=12.515 $Y=0.68 $X2=0 $Y2=0
cc_1034 N_A_M1010_g N_VGND_c_2152_n 0.00285175f $X=12.945 $Y=0.68 $X2=0 $Y2=0
cc_1035 N_A_M1010_g N_VGND_c_2158_n 0.00441827f $X=12.945 $Y=0.68 $X2=0 $Y2=0
cc_1036 N_A_M1026_g N_VGND_c_2159_n 0.0085125f $X=12.515 $Y=0.68 $X2=0 $Y2=0
cc_1037 N_A_M1010_g N_VGND_c_2159_n 0.00847227f $X=12.945 $Y=0.68 $X2=0 $Y2=0
cc_1038 SUM N_VPWR_c_1628_n 0.019758f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_1039 N_SUM_M1018_s N_VPWR_c_1620_n 0.0023218f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_1040 SUM N_VPWR_c_1620_n 0.012508f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_1041 SUM N_COUT_c_1751_n 0.0765593f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_1042 SUM N_COUT_c_1777_n 0.0128808f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_1043 SUM N_COUT_c_1765_n 0.00546985f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_1044 SUM N_COUT_c_1756_n 0.0124395f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_1045 SUM N_VGND_c_2147_n 0.00783164f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_1046 SUM N_VGND_c_2159_n 0.0113167f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_1047 SUM N_VGND_c_2160_n 0.0106618f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_1048 N_VPWR_c_1620_n N_COUT_M1007_s 0.00269239f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1049 N_VPWR_M1018_d N_COUT_c_1751_n 0.00643301f $X=0.57 $Y=1.835 $X2=0 $Y2=0
cc_1050 N_VPWR_M1018_d N_COUT_c_1765_n 0.00774586f $X=0.57 $Y=1.835 $X2=0 $Y2=0
cc_1051 N_VPWR_c_1621_n N_COUT_c_1765_n 0.0358149f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_1052 N_VPWR_c_1629_n N_COUT_c_1755_n 0.0699817f $X=2.845 $Y=3.33 $X2=0 $Y2=0
cc_1053 N_VPWR_c_1620_n N_COUT_c_1755_n 0.0438982f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1054 N_VPWR_M1018_d N_COUT_c_1767_n 0.00253815f $X=0.57 $Y=1.835 $X2=0 $Y2=0
cc_1055 N_VPWR_c_1621_n N_COUT_c_1767_n 0.013252f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_1056 N_VPWR_c_1629_n N_COUT_c_1767_n 0.00932233f $X=2.845 $Y=3.33 $X2=0 $Y2=0
cc_1057 N_VPWR_c_1620_n N_COUT_c_1767_n 0.00646268f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1058 N_VPWR_M1018_d N_COUT_c_1756_n 0.0139143f $X=0.57 $Y=1.835 $X2=0 $Y2=0
cc_1059 N_VPWR_c_1621_n N_COUT_c_1756_n 0.0123597f $X=0.71 $Y=2.545 $X2=0 $Y2=0
cc_1060 N_VPWR_c_1629_n N_COUT_c_1757_n 0.0157238f $X=2.845 $Y=3.33 $X2=0 $Y2=0
cc_1061 N_VPWR_c_1620_n N_COUT_c_1757_n 0.00944948f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1062 N_VPWR_c_1620_n N_A_1741_367#_M1031_d 0.00239376f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1063 N_VPWR_c_1620_n N_A_1741_367#_c_1934_n 0.00346586f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1064 N_VPWR_c_1630_n N_A_1930_367#_c_2011_n 0.0665347f $X=11.62 $Y=3.33 $X2=0
+ $Y2=0
cc_1065 N_VPWR_c_1620_n N_A_1930_367#_c_2011_n 0.0404971f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1066 N_VPWR_c_1630_n N_A_1930_367#_c_2012_n 0.00967019f $X=11.62 $Y=3.33
+ $X2=0 $Y2=0
cc_1067 N_VPWR_c_1620_n N_A_1930_367#_c_2012_n 0.00571933f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1068 N_VPWR_c_1630_n N_A_1930_367#_c_2013_n 0.030286f $X=11.62 $Y=3.33 $X2=0
+ $Y2=0
cc_1069 N_VPWR_c_1620_n N_A_1930_367#_c_2013_n 0.0349729f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1070 N_VPWR_M1000_d N_A_1930_367#_c_2014_n 0.0251232f $X=11.295 $Y=1.835
+ $X2=0 $Y2=0
cc_1071 N_VPWR_c_1623_n N_A_1930_367#_c_2014_n 0.0181122f $X=11.705 $Y=3.025
+ $X2=0 $Y2=0
cc_1072 N_VPWR_c_1624_n N_A_1930_367#_c_2014_n 0.00466398f $X=12.645 $Y=3.33
+ $X2=0 $Y2=0
cc_1073 N_VPWR_c_1630_n N_A_1930_367#_c_2014_n 0.00303264f $X=11.62 $Y=3.33
+ $X2=0 $Y2=0
cc_1074 N_VPWR_c_1620_n N_A_1930_367#_c_2014_n 0.0137511f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1075 N_VPWR_c_1630_n N_A_1930_367#_c_2016_n 0.0178668f $X=11.62 $Y=3.33 $X2=0
+ $Y2=0
cc_1076 N_VPWR_c_1620_n N_A_1930_367#_c_2016_n 0.0108239f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1077 N_VPWR_M1000_d N_A_1930_367#_c_2071_n 0.0118919f $X=11.295 $Y=1.835
+ $X2=0 $Y2=0
cc_1078 N_VPWR_c_1630_n N_A_1930_367#_c_2071_n 0.00380301f $X=11.62 $Y=3.33
+ $X2=0 $Y2=0
cc_1079 N_VPWR_c_1620_n N_A_1930_367#_c_2071_n 0.00542667f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1080 N_VPWR_c_1623_n N_A_1930_367#_c_2017_n 0.0122778f $X=11.705 $Y=3.025
+ $X2=0 $Y2=0
cc_1081 N_VPWR_c_1624_n N_A_1930_367#_c_2017_n 0.0220321f $X=12.645 $Y=3.33
+ $X2=0 $Y2=0
cc_1082 N_VPWR_c_1625_n N_A_1930_367#_c_2017_n 0.0144496f $X=12.73 $Y=2.225
+ $X2=0 $Y2=0
cc_1083 N_VPWR_c_1620_n N_A_1930_367#_c_2017_n 0.0125808f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1084 N_COUT_c_1751_n N_VGND_M1006_d 0.0120312f $X=0.72 $Y=2.03 $X2=-0.19
+ $Y2=-0.245
cc_1085 N_COUT_c_1752_n N_VGND_M1006_d 0.00908711f $X=1.515 $Y=0.825 $X2=-0.19
+ $Y2=-0.245
cc_1086 N_COUT_c_1777_n N_VGND_M1006_d 0.00502249f $X=0.805 $Y=0.825 $X2=-0.19
+ $Y2=-0.245
cc_1087 N_COUT_c_1752_n N_VGND_c_2147_n 0.013723f $X=1.515 $Y=0.825 $X2=0 $Y2=0
cc_1088 N_COUT_c_1777_n N_VGND_c_2147_n 0.0118826f $X=0.805 $Y=0.825 $X2=0 $Y2=0
cc_1089 COUT N_VGND_c_2147_n 0.00477859f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_1090 COUT N_VGND_c_2148_n 0.0154737f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_1091 N_COUT_c_1752_n N_VGND_c_2153_n 0.00647397f $X=1.515 $Y=0.825 $X2=0
+ $Y2=0
cc_1092 COUT N_VGND_c_2153_n 0.0268419f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_1093 N_COUT_c_1752_n N_VGND_c_2159_n 0.012361f $X=1.515 $Y=0.825 $X2=0 $Y2=0
cc_1094 N_COUT_c_1777_n N_VGND_c_2159_n 0.00127336f $X=0.805 $Y=0.825 $X2=0
+ $Y2=0
cc_1095 COUT N_VGND_c_2159_n 0.0197958f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_1096 N_COUT_c_1777_n N_VGND_c_2160_n 3.81535e-19 $X=0.805 $Y=0.825 $X2=0
+ $Y2=0
cc_1097 N_A_1741_367#_c_1934_n N_A_1930_367#_M1021_d 0.00996555f $X=10.76
+ $Y=2.415 $X2=0 $Y2=0
cc_1098 N_A_1741_367#_c_1922_n N_A_1930_367#_c_2000_n 0.00768338f $X=8.975
+ $Y=0.78 $X2=0 $Y2=0
cc_1099 N_A_1741_367#_c_1924_n N_A_1930_367#_c_2000_n 0.0816446f $X=8.872
+ $Y=1.76 $X2=0 $Y2=0
cc_1100 N_A_1741_367#_c_1934_n N_A_1930_367#_c_2011_n 0.0221922f $X=10.76
+ $Y=2.415 $X2=0 $Y2=0
cc_1101 N_A_1741_367#_c_1929_n N_A_1930_367#_c_2011_n 0.0248902f $X=8.85
+ $Y=2.415 $X2=0 $Y2=0
cc_1102 N_A_1741_367#_c_1922_n N_A_1930_367#_c_2001_n 0.0443682f $X=8.975
+ $Y=0.78 $X2=0 $Y2=0
cc_1103 N_A_1741_367#_c_1922_n N_A_1930_367#_c_2002_n 0.0126928f $X=8.975
+ $Y=0.78 $X2=0 $Y2=0
cc_1104 N_A_1741_367#_M1031_d N_A_1930_367#_c_2013_n 0.00483357f $X=10.785
+ $Y=1.835 $X2=0 $Y2=0
cc_1105 N_A_1741_367#_c_1934_n N_A_1930_367#_c_2013_n 0.0617847f $X=10.76
+ $Y=2.415 $X2=0 $Y2=0
cc_1106 N_A_1741_367#_c_1956_n N_A_1930_367#_c_2013_n 0.00308902f $X=11.18
+ $Y=2.045 $X2=0 $Y2=0
cc_1107 N_A_1741_367#_M1009_d N_A_1930_367#_c_2005_n 0.00270919f $X=10.785
+ $Y=0.595 $X2=0 $Y2=0
cc_1108 N_A_1741_367#_c_1938_n N_A_1930_367#_c_2005_n 0.0177591f $X=11.04
+ $Y=0.935 $X2=0 $Y2=0
cc_1109 N_A_1741_367#_c_1922_n N_A_1930_367#_c_2008_n 0.0129484f $X=8.975
+ $Y=0.78 $X2=0 $Y2=0
cc_1110 N_A_1741_367#_c_1924_n N_A_1930_367#_c_2008_n 0.00177249f $X=8.872
+ $Y=1.76 $X2=0 $Y2=0
cc_1111 N_A_1741_367#_c_1934_n N_A_1930_367#_c_2016_n 0.0236666f $X=10.76
+ $Y=2.415 $X2=0 $Y2=0
cc_1112 N_A_1930_367#_c_2005_n N_VGND_M1019_d 8.52337e-19 $X=11.305 $Y=0.35
+ $X2=0 $Y2=0
cc_1113 N_A_1930_367#_c_2066_n N_VGND_M1019_d 0.00610762f $X=11.39 $Y=0.85 $X2=0
+ $Y2=0
cc_1114 N_A_1930_367#_c_2006_n N_VGND_M1019_d 0.0134981f $X=12.135 $Y=0.935
+ $X2=0 $Y2=0
cc_1115 N_A_1930_367#_c_2079_n N_VGND_M1019_d 0.00119004f $X=11.475 $Y=0.935
+ $X2=0 $Y2=0
cc_1116 N_A_1930_367#_c_2003_n N_VGND_c_2149_n 0.00386812f $X=8.71 $Y=0.35 $X2=0
+ $Y2=0
cc_1117 N_A_1930_367#_c_2005_n N_VGND_c_2150_n 0.0139148f $X=11.305 $Y=0.35
+ $X2=0 $Y2=0
cc_1118 N_A_1930_367#_c_2066_n N_VGND_c_2150_n 0.0168102f $X=11.39 $Y=0.85 $X2=0
+ $Y2=0
cc_1119 N_A_1930_367#_c_2006_n N_VGND_c_2150_n 0.0189082f $X=12.135 $Y=0.935
+ $X2=0 $Y2=0
cc_1120 N_A_1930_367#_c_2007_n N_VGND_c_2150_n 0.0217905f $X=12.3 $Y=0.505 $X2=0
+ $Y2=0
cc_1121 N_A_1930_367#_c_2007_n N_VGND_c_2151_n 0.0151738f $X=12.3 $Y=0.505 $X2=0
+ $Y2=0
cc_1122 N_A_1930_367#_c_2006_n N_VGND_c_2152_n 0.00752767f $X=12.135 $Y=0.935
+ $X2=0 $Y2=0
cc_1123 N_A_1930_367#_c_2007_n N_VGND_c_2152_n 0.0189298f $X=12.3 $Y=0.505 $X2=0
+ $Y2=0
cc_1124 N_A_1930_367#_c_2002_n N_VGND_c_2157_n 0.0646808f $X=9.785 $Y=0.35 $X2=0
+ $Y2=0
cc_1125 N_A_1930_367#_c_2003_n N_VGND_c_2157_n 0.0114574f $X=8.71 $Y=0.35 $X2=0
+ $Y2=0
cc_1126 N_A_1930_367#_c_2005_n N_VGND_c_2157_n 0.0826913f $X=11.305 $Y=0.35
+ $X2=0 $Y2=0
cc_1127 N_A_1930_367#_c_2009_n N_VGND_c_2157_n 0.0222408f $X=9.95 $Y=0.35 $X2=0
+ $Y2=0
cc_1128 N_A_1930_367#_c_2002_n N_VGND_c_2159_n 0.0357328f $X=9.785 $Y=0.35 $X2=0
+ $Y2=0
cc_1129 N_A_1930_367#_c_2003_n N_VGND_c_2159_n 0.00589978f $X=8.71 $Y=0.35 $X2=0
+ $Y2=0
cc_1130 N_A_1930_367#_c_2005_n N_VGND_c_2159_n 0.0498801f $X=11.305 $Y=0.35
+ $X2=0 $Y2=0
cc_1131 N_A_1930_367#_c_2006_n N_VGND_c_2159_n 0.0148853f $X=12.135 $Y=0.935
+ $X2=0 $Y2=0
cc_1132 N_A_1930_367#_c_2007_n N_VGND_c_2159_n 0.0120712f $X=12.3 $Y=0.505 $X2=0
+ $Y2=0
cc_1133 N_A_1930_367#_c_2009_n N_VGND_c_2159_n 0.0114525f $X=9.95 $Y=0.35 $X2=0
+ $Y2=0
