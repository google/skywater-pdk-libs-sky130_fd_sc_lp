* File: sky130_fd_sc_lp__or4b_4.pxi.spice
* Created: Fri Aug 28 11:25:59 2020
* 
x_PM_SKY130_FD_SC_LP__OR4B_4%A_83_21# N_A_83_21#_M1006_d N_A_83_21#_M1003_d
+ N_A_83_21#_M1010_d N_A_83_21#_M1000_g N_A_83_21#_M1001_g N_A_83_21#_M1007_g
+ N_A_83_21#_M1005_g N_A_83_21#_M1008_g N_A_83_21#_M1011_g N_A_83_21#_M1012_g
+ N_A_83_21#_M1014_g N_A_83_21#_c_106_n N_A_83_21#_c_107_n N_A_83_21#_c_108_n
+ N_A_83_21#_c_209_p N_A_83_21#_c_215_p N_A_83_21#_c_109_n N_A_83_21#_c_216_p
+ N_A_83_21#_c_117_n N_A_83_21#_c_148_p N_A_83_21#_c_110_n N_A_83_21#_c_111_n
+ N_A_83_21#_c_118_n N_A_83_21#_c_112_n PM_SKY130_FD_SC_LP__OR4B_4%A_83_21#
x_PM_SKY130_FD_SC_LP__OR4B_4%A N_A_M1006_g N_A_M1015_g A N_A_c_227_n N_A_c_228_n
+ PM_SKY130_FD_SC_LP__OR4B_4%A
x_PM_SKY130_FD_SC_LP__OR4B_4%B N_B_M1013_g N_B_M1016_g B B B B N_B_c_265_n
+ N_B_c_266_n PM_SKY130_FD_SC_LP__OR4B_4%B
x_PM_SKY130_FD_SC_LP__OR4B_4%C N_C_c_305_n N_C_M1004_g N_C_c_307_n N_C_M1003_g C
+ C C C N_C_c_308_n PM_SKY130_FD_SC_LP__OR4B_4%C
x_PM_SKY130_FD_SC_LP__OR4B_4%A_737_315# N_A_737_315#_M1017_d
+ N_A_737_315#_M1002_d N_A_737_315#_c_347_n N_A_737_315#_M1010_g
+ N_A_737_315#_c_341_n N_A_737_315#_M1009_g N_A_737_315#_c_342_n
+ N_A_737_315#_c_343_n N_A_737_315#_c_349_n N_A_737_315#_c_350_n
+ N_A_737_315#_c_344_n N_A_737_315#_c_351_n N_A_737_315#_c_345_n
+ N_A_737_315#_c_346_n PM_SKY130_FD_SC_LP__OR4B_4%A_737_315#
x_PM_SKY130_FD_SC_LP__OR4B_4%D_N N_D_N_M1017_g N_D_N_M1002_g N_D_N_c_403_n
+ N_D_N_c_407_n D_N D_N N_D_N_c_409_n PM_SKY130_FD_SC_LP__OR4B_4%D_N
x_PM_SKY130_FD_SC_LP__OR4B_4%VPWR N_VPWR_M1001_d N_VPWR_M1005_d N_VPWR_M1014_d
+ N_VPWR_M1002_s N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n N_VPWR_c_439_n
+ N_VPWR_c_440_n VPWR N_VPWR_c_441_n N_VPWR_c_442_n N_VPWR_c_443_n
+ N_VPWR_c_444_n N_VPWR_c_435_n N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n
+ PM_SKY130_FD_SC_LP__OR4B_4%VPWR
x_PM_SKY130_FD_SC_LP__OR4B_4%X N_X_M1000_d N_X_M1008_d N_X_M1001_s N_X_M1011_s
+ N_X_c_509_n N_X_c_510_n N_X_c_512_n N_X_c_561_p N_X_c_545_n N_X_c_523_n
+ N_X_c_513_n N_X_c_532_n N_X_c_514_n N_X_c_535_n X X N_X_c_516_n X
+ PM_SKY130_FD_SC_LP__OR4B_4%X
x_PM_SKY130_FD_SC_LP__OR4B_4%VGND N_VGND_M1000_s N_VGND_M1007_s N_VGND_M1012_s
+ N_VGND_M1013_d N_VGND_M1009_d N_VGND_c_579_n N_VGND_c_580_n N_VGND_c_581_n
+ N_VGND_c_582_n N_VGND_c_583_n N_VGND_c_584_n N_VGND_c_585_n VGND
+ N_VGND_c_586_n N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n
+ N_VGND_c_591_n N_VGND_c_592_n N_VGND_c_593_n PM_SKY130_FD_SC_LP__OR4B_4%VGND
cc_1 VNB N_A_83_21#_M1000_g 0.0235711f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_2 VNB N_A_83_21#_M1001_g 0.00268533f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_3 VNB N_A_83_21#_M1007_g 0.0205482f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.655
cc_4 VNB N_A_83_21#_M1005_g 0.00249019f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_5 VNB N_A_83_21#_M1008_g 0.0205534f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_6 VNB N_A_83_21#_M1011_g 0.00249134f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_7 VNB N_A_83_21#_M1012_g 0.0202421f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_8 VNB N_A_83_21#_M1014_g 0.00243186f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_9 VNB N_A_83_21#_c_106_n 0.00251486f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.44
cc_10 VNB N_A_83_21#_c_107_n 0.0018086f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.355
cc_11 VNB N_A_83_21#_c_108_n 0.00643342f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=1.085
cc_12 VNB N_A_83_21#_c_109_n 0.00861478f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=1.085
cc_13 VNB N_A_83_21#_c_110_n 0.00491141f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=1.085
cc_14 VNB N_A_83_21#_c_111_n 0.00434787f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=1.085
cc_15 VNB N_A_83_21#_c_112_n 0.0781667f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.44
cc_16 VNB N_A_M1006_g 0.0244732f $X=-0.19 $Y=-0.245 $X2=3.835 $Y2=1.835
cc_17 VNB N_A_c_227_n 0.0260686f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_18 VNB N_A_c_228_n 9.21456e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_M1013_g 0.0267618f $X=-0.19 $Y=-0.245 $X2=3.835 $Y2=1.835
cc_20 VNB N_B_c_265_n 0.0239251f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.275
cc_21 VNB N_B_c_266_n 0.00387868f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.655
cc_22 VNB N_C_c_305_n 0.0403345f $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=0.235
cc_23 VNB N_C_M1004_g 0.00256088f $X=-0.19 $Y=-0.245 $X2=3.835 $Y2=1.835
cc_24 VNB N_C_c_307_n 0.0174266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C_c_308_n 0.00684527f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.275
cc_26 VNB N_A_737_315#_c_341_n 0.018314f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.275
cc_27 VNB N_A_737_315#_c_342_n 9.01663e-19 $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.605
cc_28 VNB N_A_737_315#_c_343_n 0.0164283f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_29 VNB N_A_737_315#_c_344_n 0.0201483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_737_315#_c_345_n 0.00516007f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_31 VNB N_A_737_315#_c_346_n 0.0668661f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.275
cc_32 VNB N_D_N_M1017_g 0.0470129f $X=-0.19 $Y=-0.245 $X2=3.835 $Y2=1.835
cc_33 VNB N_D_N_c_403_n 0.0170344f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_34 VNB D_N 0.0101808f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.605
cc_35 VNB N_VPWR_c_435_n 0.223389f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=0.42
cc_36 VNB N_X_c_509_n 0.00404319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_510_n 0.00886058f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.605
cc_38 VNB X 0.0242612f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.44
cc_39 VNB N_VGND_c_579_n 0.0108441f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_40 VNB N_VGND_c_580_n 0.0261041f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.275
cc_41 VNB N_VGND_c_581_n 3.12649e-19 $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.605
cc_42 VNB N_VGND_c_582_n 3.16188e-19 $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.275
cc_43 VNB N_VGND_c_583_n 0.00174533f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.605
cc_44 VNB N_VGND_c_584_n 0.0133644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_585_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.275
cc_46 VNB N_VGND_c_586_n 0.0122054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_587_n 0.0133881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_588_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.175
cc_49 VNB N_VGND_c_589_n 0.019591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_590_n 0.277368f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=1.085
cc_51 VNB N_VGND_c_591_n 0.00436274f $X=-0.19 $Y=-0.245 $X2=3.945 $Y2=1.175
cc_52 VNB N_VGND_c_592_n 0.010461f $X=-0.19 $Y=-0.245 $X2=3.972 $Y2=1.98
cc_53 VNB N_VGND_c_593_n 0.0354759f $X=-0.19 $Y=-0.245 $X2=3.972 $Y2=1.815
cc_54 VPB N_A_83_21#_M1001_g 0.0226516f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_55 VPB N_A_83_21#_M1005_g 0.0183934f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_56 VPB N_A_83_21#_M1011_g 0.0184118f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_57 VPB N_A_83_21#_M1014_g 0.0206208f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_58 VPB N_A_83_21#_c_117_n 8.51343e-19 $X=-0.19 $Y=1.655 $X2=3.972 $Y2=1.932
cc_59 VPB N_A_83_21#_c_118_n 0.00127423f $X=-0.19 $Y=1.655 $X2=3.972 $Y2=1.815
cc_60 VPB N_A_M1015_g 0.0192297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_c_227_n 0.00647256f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.655
cc_62 VPB N_A_c_228_n 0.00310844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_B_M1016_g 0.0177506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_B_c_265_n 0.00819893f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.275
cc_65 VPB N_B_c_266_n 0.00245768f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.655
cc_66 VPB N_C_M1004_g 0.0206919f $X=-0.19 $Y=1.655 $X2=3.835 $Y2=1.835
cc_67 VPB N_C_c_308_n 0.00274791f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.275
cc_68 VPB N_A_737_315#_c_347_n 0.0203376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_737_315#_c_342_n 0.0146744f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.605
cc_70 VPB N_A_737_315#_c_349_n 0.0168327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_737_315#_c_350_n 0.0074154f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.275
cc_72 VPB N_A_737_315#_c_351_n 0.0231853f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_737_315#_c_346_n 0.0308699f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=1.275
cc_74 VPB N_D_N_M1002_g 0.0471177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_D_N_c_403_n 0.00463815f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.655
cc_76 VPB N_D_N_c_407_n 0.0196212f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB D_N 0.0246006f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.605
cc_78 VPB N_D_N_c_409_n 0.0307752f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.655
cc_79 VPB N_VPWR_c_436_n 0.0108182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_437_n 0.0439112f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_81 VPB N_VPWR_c_438_n 3.18512e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_439_n 0.00493704f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=0.655
cc_83 VPB N_VPWR_c_440_n 0.00830804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_441_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_442_n 0.0151002f $X=-0.19 $Y=1.655 $X2=1.735 $Y2=1.44
cc_86 VPB N_VPWR_c_443_n 0.0599258f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.44
cc_87 VPB N_VPWR_c_444_n 0.015705f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=0.995
cc_88 VPB N_VPWR_c_435_n 0.0560232f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=0.42
cc_89 VPB N_VPWR_c_446_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=0.42
cc_90 VPB N_VPWR_c_447_n 0.00631825f $X=-0.19 $Y=1.655 $X2=3.945 $Y2=1.175
cc_91 VPB N_VPWR_c_448_n 0.00548851f $X=-0.19 $Y=1.655 $X2=3.972 $Y2=1.98
cc_92 VPB N_X_c_512_n 0.00142506f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_93 VPB N_X_c_513_n 0.0049094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_X_c_514_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.44
cc_95 VPB X 0.00198241f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.44
cc_96 VPB N_X_c_516_n 0.00892113f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=0.995
cc_97 N_A_83_21#_M1012_g N_A_M1006_g 0.0200391f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_98 N_A_83_21#_c_107_n N_A_M1006_g 0.00315833f $X=1.82 $Y=1.355 $X2=0 $Y2=0
cc_99 N_A_83_21#_c_108_n N_A_M1006_g 0.0147579f $X=2.35 $Y=1.085 $X2=0 $Y2=0
cc_100 N_A_83_21#_M1014_g N_A_M1015_g 0.0123164f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A_83_21#_c_106_n N_A_c_227_n 0.00106352f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_102 N_A_83_21#_c_108_n N_A_c_227_n 0.00214237f $X=2.35 $Y=1.085 $X2=0 $Y2=0
cc_103 N_A_83_21#_c_110_n N_A_c_227_n 0.00217735f $X=2.455 $Y=1.085 $X2=0 $Y2=0
cc_104 N_A_83_21#_c_112_n N_A_c_227_n 0.0214812f $X=1.78 $Y=1.44 $X2=0 $Y2=0
cc_105 N_A_83_21#_M1014_g N_A_c_228_n 8.92346e-19 $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_83_21#_c_106_n N_A_c_228_n 0.0140311f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_107 N_A_83_21#_c_107_n N_A_c_228_n 6.96048e-19 $X=1.82 $Y=1.355 $X2=0 $Y2=0
cc_108 N_A_83_21#_c_108_n N_A_c_228_n 0.0178143f $X=2.35 $Y=1.085 $X2=0 $Y2=0
cc_109 N_A_83_21#_c_112_n N_A_c_228_n 0.00125866f $X=1.78 $Y=1.44 $X2=0 $Y2=0
cc_110 N_A_83_21#_c_109_n N_B_M1013_g 0.0150872f $X=3.57 $Y=1.085 $X2=0 $Y2=0
cc_111 N_A_83_21#_c_109_n N_B_c_265_n 0.00376228f $X=3.57 $Y=1.085 $X2=0 $Y2=0
cc_112 N_A_83_21#_c_109_n N_B_c_266_n 0.0231932f $X=3.57 $Y=1.085 $X2=0 $Y2=0
cc_113 N_A_83_21#_c_110_n N_B_c_266_n 0.00693362f $X=2.455 $Y=1.085 $X2=0 $Y2=0
cc_114 N_A_83_21#_c_109_n N_C_c_305_n 0.00705389f $X=3.57 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_83_21#_c_118_n N_C_c_305_n 2.71729e-19 $X=3.972 $Y=1.815 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A_83_21#_c_109_n N_C_c_307_n 0.014869f $X=3.57 $Y=1.085 $X2=0 $Y2=0
cc_117 N_A_83_21#_c_118_n N_C_c_307_n 9.89127e-19 $X=3.972 $Y=1.815 $X2=0 $Y2=0
cc_118 N_A_83_21#_c_109_n N_C_c_308_n 0.0440175f $X=3.57 $Y=1.085 $X2=0 $Y2=0
cc_119 N_A_83_21#_c_111_n N_C_c_308_n 0.0106815f $X=3.665 $Y=1.085 $X2=0 $Y2=0
cc_120 N_A_83_21#_c_118_n N_C_c_308_n 0.0397119f $X=3.972 $Y=1.815 $X2=0 $Y2=0
cc_121 N_A_83_21#_c_118_n N_A_737_315#_c_347_n 0.0054879f $X=3.972 $Y=1.815
+ $X2=0 $Y2=0
cc_122 N_A_83_21#_c_111_n N_A_737_315#_c_341_n 0.0142554f $X=3.665 $Y=1.085
+ $X2=0 $Y2=0
cc_123 N_A_83_21#_c_118_n N_A_737_315#_c_341_n 2.82924e-19 $X=3.972 $Y=1.815
+ $X2=0 $Y2=0
cc_124 N_A_83_21#_c_117_n N_A_737_315#_c_342_n 0.0442784f $X=3.972 $Y=1.932
+ $X2=0 $Y2=0
cc_125 N_A_83_21#_c_118_n N_A_737_315#_c_342_n 0.0177305f $X=3.972 $Y=1.815
+ $X2=0 $Y2=0
cc_126 N_A_83_21#_c_148_p N_A_737_315#_c_350_n 0.0144399f $X=3.975 $Y=1.98 $X2=0
+ $Y2=0
cc_127 N_A_83_21#_c_118_n N_A_737_315#_c_345_n 0.0226855f $X=3.972 $Y=1.815
+ $X2=0 $Y2=0
cc_128 N_A_83_21#_c_117_n N_A_737_315#_c_346_n 0.00275985f $X=3.972 $Y=1.932
+ $X2=0 $Y2=0
cc_129 N_A_83_21#_c_111_n N_A_737_315#_c_346_n 0.0043118f $X=3.665 $Y=1.085
+ $X2=0 $Y2=0
cc_130 N_A_83_21#_c_118_n N_A_737_315#_c_346_n 0.0276205f $X=3.972 $Y=1.815
+ $X2=0 $Y2=0
cc_131 N_A_83_21#_c_111_n N_D_N_M1017_g 0.00271582f $X=3.665 $Y=1.085 $X2=0
+ $Y2=0
cc_132 N_A_83_21#_c_117_n N_D_N_M1002_g 5.80193e-19 $X=3.972 $Y=1.932 $X2=0
+ $Y2=0
cc_133 N_A_83_21#_c_148_p N_D_N_M1002_g 0.00424582f $X=3.975 $Y=1.98 $X2=0 $Y2=0
cc_134 N_A_83_21#_M1001_g N_VPWR_c_437_n 0.0169028f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_83_21#_M1005_g N_VPWR_c_437_n 7.44145e-19 $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A_83_21#_M1001_g N_VPWR_c_438_n 7.44145e-19 $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A_83_21#_M1005_g N_VPWR_c_438_n 0.0154271f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A_83_21#_M1011_g N_VPWR_c_438_n 0.0155524f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_83_21#_M1014_g N_VPWR_c_438_n 8.34461e-19 $X=1.78 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_83_21#_M1014_g N_VPWR_c_439_n 0.00269741f $X=1.78 $Y=2.465 $X2=0
+ $Y2=0
cc_141 N_A_83_21#_c_148_p N_VPWR_c_440_n 0.0177095f $X=3.975 $Y=1.98 $X2=0 $Y2=0
cc_142 N_A_83_21#_M1001_g N_VPWR_c_441_n 0.00486043f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_83_21#_M1005_g N_VPWR_c_441_n 0.00486043f $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_83_21#_M1011_g N_VPWR_c_442_n 0.00486043f $X=1.35 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_83_21#_M1014_g N_VPWR_c_442_n 0.00571722f $X=1.78 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_83_21#_c_148_p N_VPWR_c_443_n 0.0151289f $X=3.975 $Y=1.98 $X2=0 $Y2=0
cc_147 N_A_83_21#_M1010_d N_VPWR_c_435_n 0.00323f $X=3.835 $Y=1.835 $X2=0 $Y2=0
cc_148 N_A_83_21#_M1001_g N_VPWR_c_435_n 0.00824727f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_83_21#_M1005_g N_VPWR_c_435_n 0.00824727f $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_83_21#_M1011_g N_VPWR_c_435_n 0.00824727f $X=1.35 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_83_21#_M1014_g N_VPWR_c_435_n 0.0105481f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_83_21#_c_148_p N_VPWR_c_435_n 0.0090585f $X=3.975 $Y=1.98 $X2=0 $Y2=0
cc_153 N_A_83_21#_M1000_g N_X_c_509_n 0.0156099f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_154 N_A_83_21#_M1007_g N_X_c_509_n 0.00311953f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_155 N_A_83_21#_c_106_n N_X_c_509_n 0.0208464f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_156 N_A_83_21#_c_112_n N_X_c_509_n 0.00255521f $X=1.78 $Y=1.44 $X2=0 $Y2=0
cc_157 N_A_83_21#_M1001_g N_X_c_512_n 0.0163482f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_83_21#_c_106_n N_X_c_512_n 0.0072485f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_159 N_A_83_21#_M1007_g N_X_c_523_n 0.0121185f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_160 N_A_83_21#_M1008_g N_X_c_523_n 0.0113554f $X=1.35 $Y=0.655 $X2=0 $Y2=0
cc_161 N_A_83_21#_c_106_n N_X_c_523_n 0.0155221f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_162 N_A_83_21#_c_112_n N_X_c_523_n 0.00186738f $X=1.78 $Y=1.44 $X2=0 $Y2=0
cc_163 N_A_83_21#_M1005_g N_X_c_513_n 0.0139345f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A_83_21#_M1011_g N_X_c_513_n 0.0139345f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_83_21#_M1014_g N_X_c_513_n 0.0049246f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A_83_21#_c_106_n N_X_c_513_n 0.0664507f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_167 N_A_83_21#_c_112_n N_X_c_513_n 0.00503231f $X=1.78 $Y=1.44 $X2=0 $Y2=0
cc_168 N_A_83_21#_M1014_g N_X_c_532_n 0.0131273f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_83_21#_c_106_n N_X_c_514_n 0.0153308f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_170 N_A_83_21#_c_112_n N_X_c_514_n 0.00256759f $X=1.78 $Y=1.44 $X2=0 $Y2=0
cc_171 N_A_83_21#_c_106_n N_X_c_535_n 0.0056637f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_172 N_A_83_21#_c_112_n N_X_c_535_n 0.00193203f $X=1.78 $Y=1.44 $X2=0 $Y2=0
cc_173 N_A_83_21#_M1000_g X 0.02006f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A_83_21#_c_106_n X 0.0137867f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_175 N_A_83_21#_c_108_n N_VGND_M1012_s 0.00219369f $X=2.35 $Y=1.085 $X2=0
+ $Y2=0
cc_176 N_A_83_21#_c_109_n N_VGND_M1013_d 0.00652527f $X=3.57 $Y=1.085 $X2=0
+ $Y2=0
cc_177 N_A_83_21#_c_111_n N_VGND_M1009_d 0.00158361f $X=3.665 $Y=1.085 $X2=0
+ $Y2=0
cc_178 N_A_83_21#_M1000_g N_VGND_c_580_n 0.0112208f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_179 N_A_83_21#_M1007_g N_VGND_c_580_n 6.48667e-19 $X=0.92 $Y=0.655 $X2=0
+ $Y2=0
cc_180 N_A_83_21#_M1000_g N_VGND_c_581_n 5.14991e-19 $X=0.49 $Y=0.655 $X2=0
+ $Y2=0
cc_181 N_A_83_21#_M1007_g N_VGND_c_581_n 0.00663779f $X=0.92 $Y=0.655 $X2=0
+ $Y2=0
cc_182 N_A_83_21#_M1008_g N_VGND_c_581_n 0.00844802f $X=1.35 $Y=0.655 $X2=0
+ $Y2=0
cc_183 N_A_83_21#_M1012_g N_VGND_c_581_n 0.00111219f $X=1.78 $Y=0.655 $X2=0
+ $Y2=0
cc_184 N_A_83_21#_M1008_g N_VGND_c_582_n 0.00111027f $X=1.35 $Y=0.655 $X2=0
+ $Y2=0
cc_185 N_A_83_21#_M1012_g N_VGND_c_582_n 0.0102498f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_186 N_A_83_21#_c_108_n N_VGND_c_582_n 0.0170884f $X=2.35 $Y=1.085 $X2=0 $Y2=0
cc_187 N_A_83_21#_c_209_p N_VGND_c_582_n 2.89978e-19 $X=1.905 $Y=1.085 $X2=0
+ $Y2=0
cc_188 N_A_83_21#_c_109_n N_VGND_c_583_n 0.044913f $X=3.57 $Y=1.085 $X2=0 $Y2=0
cc_189 N_A_83_21#_M1008_g N_VGND_c_584_n 0.00355956f $X=1.35 $Y=0.655 $X2=0
+ $Y2=0
cc_190 N_A_83_21#_M1012_g N_VGND_c_584_n 0.00564095f $X=1.78 $Y=0.655 $X2=0
+ $Y2=0
cc_191 N_A_83_21#_M1000_g N_VGND_c_586_n 0.00486043f $X=0.49 $Y=0.655 $X2=0
+ $Y2=0
cc_192 N_A_83_21#_M1007_g N_VGND_c_586_n 0.00355956f $X=0.92 $Y=0.655 $X2=0
+ $Y2=0
cc_193 N_A_83_21#_c_215_p N_VGND_c_587_n 0.0131621f $X=2.465 $Y=0.42 $X2=0 $Y2=0
cc_194 N_A_83_21#_c_216_p N_VGND_c_588_n 0.0124525f $X=3.665 $Y=0.42 $X2=0 $Y2=0
cc_195 N_A_83_21#_M1006_d N_VGND_c_590_n 0.00467071f $X=2.325 $Y=0.235 $X2=0
+ $Y2=0
cc_196 N_A_83_21#_M1003_d N_VGND_c_590_n 0.00536646f $X=3.525 $Y=0.235 $X2=0
+ $Y2=0
cc_197 N_A_83_21#_M1000_g N_VGND_c_590_n 0.00824727f $X=0.49 $Y=0.655 $X2=0
+ $Y2=0
cc_198 N_A_83_21#_M1007_g N_VGND_c_590_n 0.00415754f $X=0.92 $Y=0.655 $X2=0
+ $Y2=0
cc_199 N_A_83_21#_M1008_g N_VGND_c_590_n 0.00423262f $X=1.35 $Y=0.655 $X2=0
+ $Y2=0
cc_200 N_A_83_21#_M1012_g N_VGND_c_590_n 0.00959071f $X=1.78 $Y=0.655 $X2=0
+ $Y2=0
cc_201 N_A_83_21#_c_215_p N_VGND_c_590_n 0.00808656f $X=2.465 $Y=0.42 $X2=0
+ $Y2=0
cc_202 N_A_83_21#_c_216_p N_VGND_c_590_n 0.00730901f $X=3.665 $Y=0.42 $X2=0
+ $Y2=0
cc_203 N_A_83_21#_c_111_n N_VGND_c_593_n 0.00502853f $X=3.665 $Y=1.085 $X2=0
+ $Y2=0
cc_204 N_A_M1006_g N_B_M1013_g 0.0238189f $X=2.25 $Y=0.655 $X2=0 $Y2=0
cc_205 N_A_M1015_g N_B_M1016_g 0.0594807f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A_M1015_g B 0.00474347f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_M1015_g B 0.0144717f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A_c_227_n N_B_c_265_n 0.0594807f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_209 N_A_c_228_n N_B_c_265_n 3.549e-19 $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_210 N_A_c_227_n N_B_c_266_n 0.00700556f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_211 N_A_c_228_n N_B_c_266_n 0.0315825f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_212 N_A_M1015_g N_VPWR_c_439_n 0.00419107f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A_c_227_n N_VPWR_c_439_n 0.00127919f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_214 N_A_c_228_n N_VPWR_c_439_n 0.0110295f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_215 N_A_M1015_g N_VPWR_c_443_n 0.0057332f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A_M1015_g N_VPWR_c_435_n 0.0104572f $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_M1015_g N_X_c_513_n 4.91772e-19 $X=2.32 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A_c_228_n N_X_c_513_n 0.00256396f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_219 N_A_M1006_g N_VGND_c_582_n 0.00849028f $X=2.25 $Y=0.655 $X2=0 $Y2=0
cc_220 N_A_M1006_g N_VGND_c_583_n 6.33983e-19 $X=2.25 $Y=0.655 $X2=0 $Y2=0
cc_221 N_A_M1006_g N_VGND_c_587_n 0.00564095f $X=2.25 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A_M1006_g N_VGND_c_590_n 0.00950825f $X=2.25 $Y=0.655 $X2=0 $Y2=0
cc_223 N_B_M1013_g N_C_c_305_n 0.00645315f $X=2.68 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_224 N_B_c_265_n N_C_c_305_n 0.0203734f $X=2.77 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_225 N_B_c_266_n N_C_c_305_n 2.88163e-19 $X=2.77 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_226 N_B_M1016_g N_C_M1004_g 0.0466059f $X=2.68 $Y=2.465 $X2=0 $Y2=0
cc_227 N_B_c_266_n N_C_M1004_g 0.00382223f $X=2.77 $Y=1.51 $X2=0 $Y2=0
cc_228 N_B_M1013_g N_C_c_307_n 0.00564364f $X=2.68 $Y=0.655 $X2=0 $Y2=0
cc_229 N_B_M1016_g N_C_c_308_n 0.0042713f $X=2.68 $Y=2.465 $X2=0 $Y2=0
cc_230 N_B_c_265_n N_C_c_308_n 0.00235772f $X=2.77 $Y=1.51 $X2=0 $Y2=0
cc_231 N_B_c_266_n N_C_c_308_n 0.137661f $X=2.77 $Y=1.51 $X2=0 $Y2=0
cc_232 N_B_M1016_g N_VPWR_c_443_n 0.00384307f $X=2.68 $Y=2.465 $X2=0 $Y2=0
cc_233 B N_VPWR_c_443_n 0.014211f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_234 N_B_M1016_g N_VPWR_c_435_n 0.00564664f $X=2.68 $Y=2.465 $X2=0 $Y2=0
cc_235 B N_VPWR_c_435_n 0.0160821f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_236 B A_479_367# 0.00148865f $X=2.555 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_237 B A_479_367# 0.00122477f $X=2.555 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_238 N_B_c_266_n A_479_367# 0.00102518f $X=2.77 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_239 B A_551_367# 0.00212417f $X=2.555 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_240 B A_551_367# 0.00762243f $X=2.555 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_241 N_B_c_266_n A_551_367# 7.53728e-19 $X=2.77 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_242 N_B_M1013_g N_VGND_c_582_n 5.88872e-19 $X=2.68 $Y=0.655 $X2=0 $Y2=0
cc_243 N_B_M1013_g N_VGND_c_583_n 0.0111117f $X=2.68 $Y=0.655 $X2=0 $Y2=0
cc_244 N_B_M1013_g N_VGND_c_587_n 0.00486043f $X=2.68 $Y=0.655 $X2=0 $Y2=0
cc_245 N_B_M1013_g N_VGND_c_590_n 0.0082726f $X=2.68 $Y=0.655 $X2=0 $Y2=0
cc_246 N_C_c_307_n N_A_737_315#_c_341_n 0.011885f $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_247 N_C_c_305_n N_A_737_315#_c_346_n 0.0218832f $X=3.22 $Y=1.595 $X2=0 $Y2=0
cc_248 N_C_M1004_g N_A_737_315#_c_346_n 0.0435676f $X=3.22 $Y=2.465 $X2=0 $Y2=0
cc_249 N_C_c_308_n N_A_737_315#_c_346_n 0.012117f $X=3.31 $Y=1.43 $X2=0 $Y2=0
cc_250 N_C_M1004_g N_VPWR_c_443_n 0.00384307f $X=3.22 $Y=2.465 $X2=0 $Y2=0
cc_251 N_C_c_308_n N_VPWR_c_443_n 0.0213291f $X=3.31 $Y=1.43 $X2=0 $Y2=0
cc_252 N_C_M1004_g N_VPWR_c_435_n 0.00610266f $X=3.22 $Y=2.465 $X2=0 $Y2=0
cc_253 N_C_c_308_n N_VPWR_c_435_n 0.0229718f $X=3.31 $Y=1.43 $X2=0 $Y2=0
cc_254 N_C_c_308_n A_551_367# 0.0108026f $X=3.31 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_255 N_C_c_308_n A_659_367# 0.012879f $X=3.31 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_256 N_C_c_307_n N_VGND_c_583_n 0.0110629f $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_257 N_C_c_307_n N_VGND_c_588_n 0.00486043f $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_258 N_C_c_307_n N_VGND_c_590_n 0.0082726f $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_259 N_C_c_307_n N_VGND_c_593_n 6.29916e-19 $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_260 N_A_737_315#_c_341_n N_D_N_M1017_g 0.00267142f $X=3.88 $Y=1.185 $X2=0
+ $Y2=0
cc_261 N_A_737_315#_c_343_n N_D_N_M1017_g 0.0158016f $X=4.87 $Y=1.27 $X2=0 $Y2=0
cc_262 N_A_737_315#_c_344_n N_D_N_M1017_g 0.00478801f $X=4.965 $Y=0.865 $X2=0
+ $Y2=0
cc_263 N_A_737_315#_c_345_n N_D_N_M1017_g 0.00284733f $X=4.387 $Y=1.27 $X2=0
+ $Y2=0
cc_264 N_A_737_315#_c_346_n N_D_N_M1017_g 0.0310675f $X=3.88 $Y=1.455 $X2=0
+ $Y2=0
cc_265 N_A_737_315#_c_349_n N_D_N_M1002_g 0.0146512f $X=4.925 $Y=2.46 $X2=0
+ $Y2=0
cc_266 N_A_737_315#_c_351_n N_D_N_M1002_g 0.00451176f $X=5.02 $Y=2.835 $X2=0
+ $Y2=0
cc_267 N_A_737_315#_c_342_n N_D_N_c_403_n 0.00267825f $X=4.41 $Y=2.375 $X2=0
+ $Y2=0
cc_268 N_A_737_315#_c_343_n N_D_N_c_403_n 0.00177107f $X=4.87 $Y=1.27 $X2=0
+ $Y2=0
cc_269 N_A_737_315#_c_349_n N_D_N_c_403_n 0.0013374f $X=4.925 $Y=2.46 $X2=0
+ $Y2=0
cc_270 N_A_737_315#_c_349_n N_D_N_c_407_n 0.0013655f $X=4.925 $Y=2.46 $X2=0
+ $Y2=0
cc_271 N_A_737_315#_c_342_n D_N 0.0538981f $X=4.41 $Y=2.375 $X2=0 $Y2=0
cc_272 N_A_737_315#_c_343_n D_N 0.0326583f $X=4.87 $Y=1.27 $X2=0 $Y2=0
cc_273 N_A_737_315#_c_349_n D_N 0.0386651f $X=4.925 $Y=2.46 $X2=0 $Y2=0
cc_274 N_A_737_315#_c_342_n N_D_N_c_409_n 0.0173324f $X=4.41 $Y=2.375 $X2=0
+ $Y2=0
cc_275 N_A_737_315#_c_346_n N_D_N_c_409_n 0.00183821f $X=3.88 $Y=1.455 $X2=0
+ $Y2=0
cc_276 N_A_737_315#_c_347_n N_VPWR_c_440_n 0.0027598f $X=3.76 $Y=1.725 $X2=0
+ $Y2=0
cc_277 N_A_737_315#_c_349_n N_VPWR_c_440_n 0.0128399f $X=4.925 $Y=2.46 $X2=0
+ $Y2=0
cc_278 N_A_737_315#_c_350_n N_VPWR_c_440_n 0.0119971f $X=4.56 $Y=2.46 $X2=0
+ $Y2=0
cc_279 N_A_737_315#_c_351_n N_VPWR_c_440_n 0.0146718f $X=5.02 $Y=2.835 $X2=0
+ $Y2=0
cc_280 N_A_737_315#_c_347_n N_VPWR_c_443_n 0.00585385f $X=3.76 $Y=1.725 $X2=0
+ $Y2=0
cc_281 N_A_737_315#_c_351_n N_VPWR_c_444_n 0.018536f $X=5.02 $Y=2.835 $X2=0
+ $Y2=0
cc_282 N_A_737_315#_c_347_n N_VPWR_c_435_n 0.0124608f $X=3.76 $Y=1.725 $X2=0
+ $Y2=0
cc_283 N_A_737_315#_c_349_n N_VPWR_c_435_n 0.00593841f $X=4.925 $Y=2.46 $X2=0
+ $Y2=0
cc_284 N_A_737_315#_c_350_n N_VPWR_c_435_n 0.00739944f $X=4.56 $Y=2.46 $X2=0
+ $Y2=0
cc_285 N_A_737_315#_c_351_n N_VPWR_c_435_n 0.0100381f $X=5.02 $Y=2.835 $X2=0
+ $Y2=0
cc_286 N_A_737_315#_c_341_n N_VGND_c_583_n 6.2485e-19 $X=3.88 $Y=1.185 $X2=0
+ $Y2=0
cc_287 N_A_737_315#_c_341_n N_VGND_c_588_n 0.00486043f $X=3.88 $Y=1.185 $X2=0
+ $Y2=0
cc_288 N_A_737_315#_c_344_n N_VGND_c_589_n 0.00427512f $X=4.965 $Y=0.865 $X2=0
+ $Y2=0
cc_289 N_A_737_315#_c_341_n N_VGND_c_590_n 0.00822376f $X=3.88 $Y=1.185 $X2=0
+ $Y2=0
cc_290 N_A_737_315#_c_344_n N_VGND_c_590_n 0.00744821f $X=4.965 $Y=0.865 $X2=0
+ $Y2=0
cc_291 N_A_737_315#_c_341_n N_VGND_c_593_n 0.013384f $X=3.88 $Y=1.185 $X2=0
+ $Y2=0
cc_292 N_A_737_315#_c_343_n N_VGND_c_593_n 0.0088133f $X=4.87 $Y=1.27 $X2=0
+ $Y2=0
cc_293 N_A_737_315#_c_345_n N_VGND_c_593_n 0.0302111f $X=4.387 $Y=1.27 $X2=0
+ $Y2=0
cc_294 N_A_737_315#_c_346_n N_VGND_c_593_n 0.00935317f $X=3.88 $Y=1.455 $X2=0
+ $Y2=0
cc_295 N_D_N_M1002_g N_VPWR_c_440_n 0.00983143f $X=4.805 $Y=2.835 $X2=0 $Y2=0
cc_296 N_D_N_M1002_g N_VPWR_c_444_n 0.00445056f $X=4.805 $Y=2.835 $X2=0 $Y2=0
cc_297 N_D_N_M1002_g N_VPWR_c_435_n 0.00489276f $X=4.805 $Y=2.835 $X2=0 $Y2=0
cc_298 N_D_N_M1017_g N_VGND_c_589_n 0.00332367f $X=4.75 $Y=0.865 $X2=0 $Y2=0
cc_299 N_D_N_M1017_g N_VGND_c_590_n 0.0038435f $X=4.75 $Y=0.865 $X2=0 $Y2=0
cc_300 N_D_N_M1017_g N_VGND_c_593_n 0.0164201f $X=4.75 $Y=0.865 $X2=0 $Y2=0
cc_301 N_VPWR_c_435_n N_X_M1001_s 0.00536646f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_302 N_VPWR_c_435_n N_X_M1011_s 0.00380103f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_303 N_VPWR_M1001_d N_X_c_512_n 2.33864e-19 $X=0.15 $Y=1.835 $X2=0 $Y2=0
cc_304 N_VPWR_c_437_n N_X_c_512_n 0.00362085f $X=0.275 $Y=2.12 $X2=0 $Y2=0
cc_305 N_VPWR_c_441_n N_X_c_545_n 0.0124525f $X=0.97 $Y=3.33 $X2=0 $Y2=0
cc_306 N_VPWR_c_435_n N_X_c_545_n 0.00730901f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_307 N_VPWR_M1005_d N_X_c_513_n 0.00176461f $X=0.995 $Y=1.835 $X2=0 $Y2=0
cc_308 N_VPWR_c_438_n N_X_c_513_n 0.0170777f $X=1.135 $Y=2.12 $X2=0 $Y2=0
cc_309 N_VPWR_c_442_n N_X_c_532_n 0.0146655f $X=1.885 $Y=3.33 $X2=0 $Y2=0
cc_310 N_VPWR_c_435_n N_X_c_532_n 0.00933292f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_311 N_VPWR_M1001_d N_X_c_516_n 0.0021884f $X=0.15 $Y=1.835 $X2=0 $Y2=0
cc_312 N_VPWR_c_437_n N_X_c_516_n 0.0203341f $X=0.275 $Y=2.12 $X2=0 $Y2=0
cc_313 N_VPWR_c_435_n A_479_367# 0.00181925f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_314 N_VPWR_c_435_n A_551_367# 0.00926526f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_315 N_VPWR_c_435_n A_659_367# 0.00338003f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_316 N_X_c_509_n N_VGND_M1000_s 2.33864e-19 $X=0.61 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_317 N_X_c_510_n N_VGND_M1000_s 0.00237659f $X=0.335 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_318 N_X_c_523_n N_VGND_M1007_s 0.00446387f $X=1.47 $Y=0.74 $X2=0 $Y2=0
cc_319 N_X_c_509_n N_VGND_c_580_n 0.00362085f $X=0.61 $Y=1.09 $X2=0 $Y2=0
cc_320 N_X_c_510_n N_VGND_c_580_n 0.0203341f $X=0.335 $Y=1.09 $X2=0 $Y2=0
cc_321 N_X_c_523_n N_VGND_c_581_n 0.016098f $X=1.47 $Y=0.74 $X2=0 $Y2=0
cc_322 N_X_c_523_n N_VGND_c_584_n 0.00235176f $X=1.47 $Y=0.74 $X2=0 $Y2=0
cc_323 N_X_c_535_n N_VGND_c_584_n 0.00501641f $X=1.565 $Y=0.65 $X2=0 $Y2=0
cc_324 N_X_c_561_p N_VGND_c_586_n 0.0124525f $X=0.705 $Y=0.42 $X2=0 $Y2=0
cc_325 N_X_c_523_n N_VGND_c_586_n 0.00235807f $X=1.47 $Y=0.74 $X2=0 $Y2=0
cc_326 N_X_M1000_d N_VGND_c_590_n 0.00396356f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_327 N_X_M1008_d N_VGND_c_590_n 0.00365119f $X=1.425 $Y=0.235 $X2=0 $Y2=0
cc_328 N_X_c_561_p N_VGND_c_590_n 0.0073074f $X=0.705 $Y=0.42 $X2=0 $Y2=0
cc_329 N_X_c_523_n N_VGND_c_590_n 0.00972279f $X=1.47 $Y=0.74 $X2=0 $Y2=0
cc_330 N_X_c_535_n N_VGND_c_590_n 0.00684215f $X=1.565 $Y=0.65 $X2=0 $Y2=0
