* File: sky130_fd_sc_lp__o2bb2a_lp.pex.spice
* Created: Wed Sep  2 10:21:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%A_86_22# 1 2 9 13 15 19 21 23 24 25 30 34
+ 41 42 44 48
c99 48 0 1.88541e-19 $X=0.865 $Y=1.025
r100 41 42 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0.962
+ $X2=2.505 $Y2=0.962
r101 38 48 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=0.8 $Y=1.025
+ $X2=0.865 $Y2=1.025
r102 38 45 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=0.8 $Y=1.025
+ $X2=0.505 $Y2=1.025
r103 37 39 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.8 $Y=1.025
+ $X2=0.8 $Y2=1.19
r104 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.8
+ $Y=1.025 $X2=0.8 $Y2=1.025
r105 34 37 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.8 $Y=0.945 $X2=0.8
+ $Y2=1.025
r106 28 44 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.49
+ $X2=2.98 $Y2=2.575
r107 28 30 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.98 $Y=2.49
+ $X2=2.98 $Y2=2.225
r108 27 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0.945
+ $X2=0.8 $Y2=0.945
r109 27 42 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=0.965 $Y=0.945
+ $X2=2.505 $Y2=0.945
r110 24 44 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=2.575
+ $X2=2.98 $Y2=2.575
r111 24 25 131.134 $w=1.68e-07 $l=2.01e-06 $layer=LI1_cond $X=2.815 $Y=2.575
+ $X2=0.805 $Y2=2.575
r112 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=2.49
+ $X2=0.805 $Y2=2.575
r113 23 39 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=0.72 $Y=2.49
+ $X2=0.72 $Y2=1.19
r114 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.865 $Y=0.86
+ $X2=0.865 $Y2=1.025
r115 17 19 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.865 $Y=0.86
+ $X2=0.865 $Y2=0.45
r116 13 21 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.555 $Y=1.555
+ $X2=0.555 $Y2=1.43
r117 13 15 254.665 $w=2.5e-07 $l=1.025e-06 $layer=POLY_cond $X=0.555 $Y=1.555
+ $X2=0.555 $Y2=2.58
r118 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.19
+ $X2=0.505 $Y2=1.025
r119 11 21 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.505 $Y=1.19
+ $X2=0.505 $Y2=1.43
r120 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=0.86
+ $X2=0.505 $Y2=1.025
r121 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.505 $Y=0.86
+ $X2=0.505 $Y2=0.45
r122 2 30 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.84
+ $Y=2.08 $X2=2.98 $Y2=2.225
r123 1 41 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.71 $X2=2.67 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%A1_N 3 7 9 10 18
c44 7 0 1.90762e-19 $X=1.365 $Y=2.58
r45 17 18 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.295 $Y=1.715
+ $X2=1.365 $Y2=1.715
r46 14 17 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.15 $Y=1.715
+ $X2=1.295 $Y2=1.715
r47 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=2.035
r48 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.715 $X2=1.15 $Y2=1.715
r49 5 18 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.88
+ $X2=1.365 $Y2=1.715
r50 5 7 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.365 $Y=1.88 $X2=1.365
+ $Y2=2.58
r51 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.295 $Y=1.55
+ $X2=1.295 $Y2=1.715
r52 1 3 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=1.295 $Y=1.55
+ $X2=1.295 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%A2_N 1 3 8 12 15 16 17 18 19 23
c45 19 0 1.67368e-19 $X=2.16 $Y=1.665
c46 17 0 1.11508e-19 $X=1.895 $Y=1.88
r47 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.895
+ $Y=1.375 $X2=1.895 $Y2=1.375
r48 19 24 4.73076 $w=6.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.895 $Y2=1.545
r49 18 24 3.83816 $w=6.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.545
+ $X2=1.895 $Y2=1.545
r50 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.895 $Y=1.715
+ $X2=1.895 $Y2=1.375
r51 16 17 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.715
+ $X2=1.895 $Y2=1.88
r52 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.21
+ $X2=1.895 $Y2=1.375
r53 10 12 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.685 $Y=0.81
+ $X2=1.805 $Y2=0.81
r54 8 17 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.925 $Y=2.58 $X2=1.925
+ $Y2=1.88
r55 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.805 $Y=0.885
+ $X2=1.805 $Y2=0.81
r56 4 15 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.805 $Y=0.885
+ $X2=1.805 $Y2=1.21
r57 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.685 $Y=0.735
+ $X2=1.685 $Y2=0.81
r58 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.685 $Y=0.735
+ $X2=1.685 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%A_298_416# 1 2 8 11 13 15 16 22 23 26 30
+ 32 39
c75 26 0 1.53316e-19 $X=2.54 $Y=2.06
c76 22 0 3.80012e-20 $X=2.67 $Y=0.43
c77 16 0 2.58786e-19 $X=2.455 $Y=2.185
c78 13 0 1.10062e-19 $X=2.945 $Y=0.595
c79 11 0 1.67368e-19 $X=2.715 $Y=2.58
r80 33 39 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.62 $Y=1.665
+ $X2=2.715 $Y2=1.665
r81 33 36 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=2.62 $Y=1.665
+ $X2=2.375 $Y2=1.665
r82 32 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=1.665
+ $X2=2.62 $Y2=1.83
r83 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.665 $X2=2.62 $Y2=1.665
r84 28 30 5.09823 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=0.472
+ $X2=2.065 $Y2=0.472
r85 26 35 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.54 $Y=2.06
+ $X2=2.54 $Y2=1.83
r86 23 43 47.6799 $w=2.78e-07 $l=2.75e-07 $layer=POLY_cond $X=2.67 $Y=0.43
+ $X2=2.945 $Y2=0.43
r87 22 30 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=2.67 $Y=0.43
+ $X2=2.065 $Y2=0.43
r88 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=0.43 $X2=2.67 $Y2=0.43
r89 16 26 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.455 $Y=2.185
+ $X2=2.54 $Y2=2.06
r90 16 18 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=2.455 $Y=2.185
+ $X2=1.66 $Y2=2.185
r91 13 43 17.1848 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=0.595
+ $X2=2.945 $Y2=0.43
r92 13 15 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.945 $Y=0.595
+ $X2=2.945 $Y2=0.92
r93 9 39 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.83
+ $X2=2.715 $Y2=1.665
r94 9 11 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.715 $Y=1.83
+ $X2=2.715 $Y2=2.58
r95 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.5
+ $X2=2.375 $Y2=1.665
r96 7 23 51.1475 $w=2.78e-07 $l=3.68375e-07 $layer=POLY_cond $X=2.375 $Y=0.595
+ $X2=2.67 $Y2=0.43
r97 7 8 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=2.375 $Y=0.595
+ $X2=2.375 $Y2=1.5
r98 2 18 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=2.08 $X2=1.66 $Y2=2.225
r99 1 28 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=1.76
+ $Y=0.24 $X2=1.9 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%B2 3 9 10 11 12 15 16 17
c47 15 0 4.18084e-20 $X=3.245 $Y=1.715
c48 10 0 3.80012e-20 $X=3.365 $Y=1.205
c49 3 0 6.80235e-20 $X=3.245 $Y=2.58
r50 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.245 $Y=1.715
+ $X2=3.245 $Y2=1.55
r51 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.245
+ $Y=1.715 $X2=3.245 $Y2=1.715
r52 12 16 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.12 $Y=1.715
+ $X2=3.245 $Y2=1.715
r53 11 17 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.335 $Y=1.355
+ $X2=3.335 $Y2=1.55
r54 10 11 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=3.365 $Y=1.205
+ $X2=3.365 $Y2=1.355
r55 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.395 $Y=0.92
+ $X2=3.395 $Y2=1.205
r56 1 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.245 $Y=1.88
+ $X2=3.245 $Y2=1.715
r57 1 3 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.245 $Y=1.88 $X2=3.245
+ $Y2=2.58
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%B1 3 7 9 12
r27 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.715
+ $X2=3.815 $Y2=1.88
r28 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.715
+ $X2=3.815 $Y2=1.55
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.815
+ $Y=1.715 $X2=3.815 $Y2=1.715
r30 9 13 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.08 $Y=1.715
+ $X2=3.815 $Y2=1.715
r31 7 14 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.825 $Y=0.92
+ $X2=3.825 $Y2=1.55
r32 3 15 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.775 $Y=2.58 $X2=3.775
+ $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%X 1 2 7 8 9 10
r17 10 26 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=2.225
r18 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r19 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.925 $X2=0.29
+ $Y2=1.295
r20 7 8 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.29 $Y=0.47 $X2=0.29
+ $Y2=0.925
r21 2 26 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=2.08 $X2=0.29 $Y2=2.225
r22 1 7 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.24 $X2=0.29 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%VPWR 1 2 3 14 18 20 22 26 28 33 42 45 49
r51 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 40 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 34 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.19 $Y2=3.33
r59 34 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 33 48 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.097 $Y2=3.33
r61 33 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.6 $Y2=3.33
r62 32 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 29 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.82 $Y2=3.33
r65 29 31 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 28 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.19 $Y2=3.33
r67 28 31 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 26 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 22 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.04 $Y=2.225
+ $X2=4.04 $Y2=2.935
r72 20 48 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.097 $Y2=3.33
r73 20 25 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=4.04 $Y=3.245
+ $X2=4.04 $Y2=2.935
r74 16 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r75 16 18 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.93
r76 12 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=3.33
r77 12 14 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.93
r78 3 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=2.08 $X2=4.04 $Y2=2.935
r79 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=2.08 $X2=4.04 $Y2=2.225
r80 2 18 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=2.08 $X2=2.19 $Y2=2.93
r81 1 14 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=2.08 $X2=0.82 $Y2=2.93
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
c49 13 0 1.10062e-19 $X=3.61 $Y=0.855
c50 9 0 1.88541e-19 $X=1.08 $Y=0.45
r51 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r52 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r54 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r55 27 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=3.57
+ $Y2=0
r56 27 29 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.695 $Y=0 $X2=4.08
+ $Y2=0
r57 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r58 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r59 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.08
+ $Y2=0
r60 23 25 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=1.245 $Y=0
+ $X2=3.12 $Y2=0
r61 22 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.57
+ $Y2=0
r62 22 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.12
+ $Y2=0
r63 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r64 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.08
+ $Y2=0
r66 17 19 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.72
+ $Y2=0
r67 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r68 15 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r69 11 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0
r70 11 13 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0.855
r71 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=0.085 $X2=1.08
+ $Y2=0
r72 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.08 $Y=0.085
+ $X2=1.08 $Y2=0.45
r73 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.47
+ $Y=0.71 $X2=3.61 $Y2=0.855
r74 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.24 $X2=1.08 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_LP%A_604_142# 1 2 9 11 12 15
r28 13 15 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.04 $Y=1.2 $X2=4.04
+ $Y2=0.96
r29 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.875 $Y=1.285
+ $X2=4.04 $Y2=1.2
r30 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.875 $Y=1.285
+ $X2=3.265 $Y2=1.285
r31 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.14 $Y=1.2
+ $X2=3.265 $Y2=1.285
r32 7 9 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.14 $Y=1.2 $X2=3.14
+ $Y2=0.92
r33 2 15 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.71 $X2=4.04 $Y2=0.96
r34 1 9 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.71 $X2=3.18 $Y2=0.92
.ends

