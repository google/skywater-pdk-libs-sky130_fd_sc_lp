* File: sky130_fd_sc_lp__o21a_1.pxi.spice
* Created: Fri Aug 28 11:03:42 2020
* 
x_PM_SKY130_FD_SC_LP__O21A_1%A_80_21# N_A_80_21#_M1005_s N_A_80_21#_M1007_d
+ N_A_80_21#_c_50_n N_A_80_21#_M1003_g N_A_80_21#_M1002_g N_A_80_21#_c_52_n
+ N_A_80_21#_c_53_n N_A_80_21#_c_62_p N_A_80_21#_c_85_p N_A_80_21#_c_54_n
+ N_A_80_21#_c_73_p N_A_80_21#_c_89_p N_A_80_21#_c_55_n
+ PM_SKY130_FD_SC_LP__O21A_1%A_80_21#
x_PM_SKY130_FD_SC_LP__O21A_1%B1 N_B1_M1005_g N_B1_M1007_g B1 N_B1_c_104_n
+ N_B1_c_105_n PM_SKY130_FD_SC_LP__O21A_1%B1
x_PM_SKY130_FD_SC_LP__O21A_1%A2 N_A2_M1000_g N_A2_M1001_g A2 A2 N_A2_c_139_n
+ PM_SKY130_FD_SC_LP__O21A_1%A2
x_PM_SKY130_FD_SC_LP__O21A_1%A1 N_A1_M1006_g N_A1_M1004_g A1 N_A1_c_173_n
+ N_A1_c_174_n PM_SKY130_FD_SC_LP__O21A_1%A1
x_PM_SKY130_FD_SC_LP__O21A_1%X N_X_M1003_s N_X_M1002_s X X X X X X X N_X_c_196_n
+ X N_X_c_199_n PM_SKY130_FD_SC_LP__O21A_1%X
x_PM_SKY130_FD_SC_LP__O21A_1%VPWR N_VPWR_M1002_d N_VPWR_M1004_d N_VPWR_c_215_n
+ N_VPWR_c_216_n N_VPWR_c_217_n VPWR N_VPWR_c_218_n N_VPWR_c_219_n
+ N_VPWR_c_214_n PM_SKY130_FD_SC_LP__O21A_1%VPWR
x_PM_SKY130_FD_SC_LP__O21A_1%VGND N_VGND_M1003_d N_VGND_M1000_d N_VGND_c_249_n
+ N_VGND_c_250_n VGND N_VGND_c_251_n N_VGND_c_252_n N_VGND_c_253_n
+ N_VGND_c_254_n N_VGND_c_255_n N_VGND_c_256_n PM_SKY130_FD_SC_LP__O21A_1%VGND
x_PM_SKY130_FD_SC_LP__O21A_1%A_300_51# N_A_300_51#_M1005_d N_A_300_51#_M1006_d
+ N_A_300_51#_c_283_n N_A_300_51#_c_284_n N_A_300_51#_c_285_n
+ N_A_300_51#_c_286_n PM_SKY130_FD_SC_LP__O21A_1%A_300_51#
cc_1 VNB N_A_80_21#_c_50_n 0.0222572f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_A_80_21#_M1002_g 0.00764058f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_3 VNB N_A_80_21#_c_52_n 0.0219644f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.515
cc_4 VNB N_A_80_21#_c_53_n 8.38913e-19 $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.93
cc_5 VNB N_A_80_21#_c_54_n 0.0102419f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.42
cc_6 VNB N_A_80_21#_c_55_n 0.0393456f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.35
cc_7 VNB N_B1_M1005_g 0.0283577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_104_n 0.00159725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_105_n 0.0340045f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.515
cc_10 VNB N_A2_M1000_g 0.0245193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A2 0.0062261f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.515
cc_12 VNB N_A2_c_139_n 0.023006f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.515
cc_13 VNB N_A1_M1006_g 0.0285539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_M1004_g 0.00176086f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_15 VNB N_A1_c_173_n 0.0481202f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.515
cc_16 VNB N_A1_c_174_n 0.0117791f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.93
cc_17 VNB N_X_c_196_n 0.0620551f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=2.49
cc_18 VNB N_VPWR_c_214_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.35
cc_19 VNB N_VGND_c_249_n 0.0094015f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_20 VNB N_VGND_c_250_n 0.00621827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_251_n 0.0152818f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.015
cc_22 VNB N_VGND_c_252_n 0.0294847f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=2.1
cc_23 VNB N_VGND_c_253_n 0.0180487f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.385
cc_24 VNB N_VGND_c_254_n 0.185774f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.085
cc_25 VNB N_VGND_c_255_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.35
cc_26 VNB N_VGND_c_256_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.35
cc_27 VNB N_A_300_51#_c_283_n 0.00120843f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_28 VNB N_A_300_51#_c_284_n 0.0140414f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_29 VNB N_A_300_51#_c_285_n 0.00445487f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_30 VNB N_A_300_51#_c_286_n 0.0313482f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.93
cc_31 VPB N_A_80_21#_M1002_g 0.0252113f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_32 VPB N_A_80_21#_c_53_n 0.00169782f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.93
cc_33 VPB N_B1_M1007_g 0.0227192f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_34 VPB N_B1_c_104_n 0.00379563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_B1_c_105_n 0.0109457f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.515
cc_36 VPB N_A2_M1001_g 0.0187037f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_37 VPB A2 0.0108226f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.515
cc_38 VPB N_A2_c_139_n 0.00624595f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.515
cc_39 VPB N_A1_M1004_g 0.0244358f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_40 VPB N_A1_c_174_n 0.00792998f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.93
cc_41 VPB X 0.0163223f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.515
cc_42 VPB N_X_c_196_n 0.00211515f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=2.49
cc_43 VPB N_X_c_199_n 0.0564945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_215_n 0.00220061f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_45 VPB N_VPWR_c_216_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_217_n 0.047982f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=1.93
cc_47 VPB N_VPWR_c_218_n 0.0265791f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_219_n 0.0309373f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.35
cc_49 VPB N_VPWR_c_214_n 0.0461496f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.35
cc_50 N_A_80_21#_c_52_n N_B1_M1005_g 0.00632417f $X=0.82 $Y=1.515 $X2=0 $Y2=0
cc_51 N_A_80_21#_c_55_n N_B1_M1005_g 0.00223708f $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_52 N_A_80_21#_M1002_g N_B1_M1007_g 0.010063f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_53 N_A_80_21#_c_53_n N_B1_M1007_g 0.00288922f $X=0.82 $Y=1.93 $X2=0 $Y2=0
cc_54 N_A_80_21#_c_62_p N_B1_M1007_g 0.0202585f $X=1.605 $Y=2.015 $X2=0 $Y2=0
cc_55 N_A_80_21#_M1002_g N_B1_c_104_n 6.64748e-19 $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_56 N_A_80_21#_c_52_n N_B1_c_104_n 0.0304792f $X=0.82 $Y=1.515 $X2=0 $Y2=0
cc_57 N_A_80_21#_c_53_n N_B1_c_104_n 0.0194299f $X=0.82 $Y=1.93 $X2=0 $Y2=0
cc_58 N_A_80_21#_c_62_p N_B1_c_104_n 0.0243999f $X=1.605 $Y=2.015 $X2=0 $Y2=0
cc_59 N_A_80_21#_c_55_n N_B1_c_104_n 2.384e-19 $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_60 N_A_80_21#_M1002_g N_B1_c_105_n 0.00548941f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_52_n N_B1_c_105_n 0.00901086f $X=0.82 $Y=1.515 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_53_n N_B1_c_105_n 5.17801e-19 $X=0.82 $Y=1.93 $X2=0 $Y2=0
cc_63 N_A_80_21#_c_62_p N_B1_c_105_n 0.00172211f $X=1.605 $Y=2.015 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_55_n N_B1_c_105_n 0.00665127f $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_73_p A2 0.0262157f $X=1.77 $Y=2.1 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_73_p N_A2_c_139_n 9.33109e-19 $X=1.77 $Y=2.1 $X2=0 $Y2=0
cc_67 N_A_80_21#_M1002_g X 0.00616529f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_52_n X 0.00157017f $X=0.82 $Y=1.515 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_53_n X 0.0128764f $X=0.82 $Y=1.93 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_55_n X 0.00613075f $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_50_n N_X_c_196_n 0.0138614f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_72 N_A_80_21#_M1002_g N_X_c_196_n 0.00361291f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_52_n N_X_c_196_n 0.0345708f $X=0.82 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_53_n N_X_c_196_n 0.00731361f $X=0.82 $Y=1.93 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_53_n N_VPWR_M1002_d 0.00145438f $X=0.82 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_76 N_A_80_21#_c_62_p N_VPWR_M1002_d 0.013459f $X=1.605 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_77 N_A_80_21#_c_85_p N_VPWR_M1002_d 0.00118409f $X=0.905 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_78 N_A_80_21#_M1002_g N_VPWR_c_215_n 0.0194707f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_62_p N_VPWR_c_215_n 0.0381982f $X=1.605 $Y=2.015 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_85_p N_VPWR_c_215_n 0.0100733f $X=0.905 $Y=2.015 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_89_p N_VPWR_c_218_n 0.0212513f $X=1.77 $Y=2.49 $X2=0 $Y2=0
cc_82 N_A_80_21#_M1002_g N_VPWR_c_219_n 0.00486043f $X=0.665 $Y=2.465 $X2=0
+ $Y2=0
cc_83 N_A_80_21#_M1007_d N_VPWR_c_214_n 0.00526034f $X=1.56 $Y=1.835 $X2=0 $Y2=0
cc_84 N_A_80_21#_M1002_g N_VPWR_c_214_n 0.00931677f $X=0.665 $Y=2.465 $X2=0
+ $Y2=0
cc_85 N_A_80_21#_c_89_p N_VPWR_c_214_n 0.0127519f $X=1.77 $Y=2.49 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_50_n N_VGND_c_249_n 0.0150697f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_52_n N_VGND_c_249_n 0.0267896f $X=0.82 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_54_n N_VGND_c_249_n 0.0504577f $X=1.21 $Y=0.42 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_55_n N_VGND_c_249_n 0.00123105f $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_50_n N_VGND_c_251_n 0.00486043f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_54_n N_VGND_c_252_n 0.0192303f $X=1.21 $Y=0.42 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_50_n N_VGND_c_254_n 0.00917987f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_54_n N_VGND_c_254_n 0.0115856f $X=1.21 $Y=0.42 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_52_n N_A_300_51#_c_285_n 0.00926935f $X=0.82 $Y=1.515 $X2=0
+ $Y2=0
cc_95 N_B1_M1005_g N_A2_M1000_g 0.0233281f $X=1.425 $Y=0.675 $X2=0 $Y2=0
cc_96 N_B1_M1007_g N_A2_M1001_g 0.0260452f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_97 N_B1_c_104_n A2 0.0280634f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_98 N_B1_c_105_n A2 0.00296801f $X=1.425 $Y=1.51 $X2=0 $Y2=0
cc_99 N_B1_c_105_n N_A2_c_139_n 0.0206549f $X=1.425 $Y=1.51 $X2=0 $Y2=0
cc_100 N_B1_M1007_g N_VPWR_c_215_n 0.0182135f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_101 N_B1_M1007_g N_VPWR_c_218_n 0.00486043f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_102 N_B1_M1007_g N_VPWR_c_214_n 0.00864313f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_103 N_B1_M1005_g N_VGND_c_249_n 0.00320371f $X=1.425 $Y=0.675 $X2=0 $Y2=0
cc_104 N_B1_M1005_g N_VGND_c_252_n 0.00565115f $X=1.425 $Y=0.675 $X2=0 $Y2=0
cc_105 N_B1_M1005_g N_VGND_c_254_n 0.0119838f $X=1.425 $Y=0.675 $X2=0 $Y2=0
cc_106 N_B1_M1005_g N_A_300_51#_c_285_n 8.72721e-19 $X=1.425 $Y=0.675 $X2=0
+ $Y2=0
cc_107 N_B1_c_105_n N_A_300_51#_c_285_n 0.00204132f $X=1.425 $Y=1.51 $X2=0 $Y2=0
cc_108 N_A2_M1000_g N_A1_M1006_g 0.0172084f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_109 N_A2_M1001_g N_A1_M1004_g 0.0565292f $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_110 A2 N_A1_c_173_n 0.00252904f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A2_c_139_n N_A1_c_173_n 0.0565292f $X=1.935 $Y=1.51 $X2=0 $Y2=0
cc_112 A2 N_A1_c_174_n 0.0282277f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A2_c_139_n N_A1_c_174_n 5.39811e-19 $X=1.935 $Y=1.51 $X2=0 $Y2=0
cc_114 N_A2_M1001_g N_VPWR_c_215_n 0.00115983f $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A2_M1001_g N_VPWR_c_217_n 0.00441827f $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A2_M1001_g N_VPWR_c_218_n 0.00585385f $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A2_M1001_g N_VPWR_c_214_n 0.0109726f $X=2.025 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A2_M1000_g N_VGND_c_250_n 0.00317939f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_119 N_A2_M1000_g N_VGND_c_252_n 0.00559232f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_120 N_A2_M1000_g N_VGND_c_254_n 0.0106256f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_121 N_A2_M1000_g N_A_300_51#_c_283_n 0.00988877f $X=1.855 $Y=0.675 $X2=0
+ $Y2=0
cc_122 N_A2_M1000_g N_A_300_51#_c_284_n 0.013442f $X=1.855 $Y=0.675 $X2=0 $Y2=0
cc_123 A2 N_A_300_51#_c_284_n 0.0282762f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A2_c_139_n N_A_300_51#_c_284_n 0.0046292f $X=1.935 $Y=1.51 $X2=0 $Y2=0
cc_125 N_A2_M1000_g N_A_300_51#_c_285_n 0.00113046f $X=1.855 $Y=0.675 $X2=0
+ $Y2=0
cc_126 A2 N_A_300_51#_c_285_n 0.0142361f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A2_c_139_n N_A_300_51#_c_285_n 2.48771e-19 $X=1.935 $Y=1.51 $X2=0 $Y2=0
cc_128 N_A2_M1000_g N_A_300_51#_c_286_n 3.84433e-19 $X=1.855 $Y=0.675 $X2=0
+ $Y2=0
cc_129 N_A1_M1004_g N_VPWR_c_217_n 0.0287066f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A1_c_173_n N_VPWR_c_217_n 0.00154747f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_131 N_A1_c_174_n N_VPWR_c_217_n 0.0261833f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_132 N_A1_M1004_g N_VPWR_c_218_n 0.00486043f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A1_M1004_g N_VPWR_c_214_n 0.00818711f $X=2.385 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A1_M1006_g N_VGND_c_250_n 0.00317939f $X=2.385 $Y=0.675 $X2=0 $Y2=0
cc_135 N_A1_M1006_g N_VGND_c_253_n 0.00559232f $X=2.385 $Y=0.675 $X2=0 $Y2=0
cc_136 N_A1_M1006_g N_VGND_c_254_n 0.0114801f $X=2.385 $Y=0.675 $X2=0 $Y2=0
cc_137 N_A1_M1006_g N_A_300_51#_c_283_n 3.85289e-19 $X=2.385 $Y=0.675 $X2=0
+ $Y2=0
cc_138 N_A1_M1006_g N_A_300_51#_c_284_n 0.0188009f $X=2.385 $Y=0.675 $X2=0 $Y2=0
cc_139 N_A1_c_173_n N_A_300_51#_c_284_n 0.00753227f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_140 N_A1_c_174_n N_A_300_51#_c_284_n 0.0274208f $X=2.59 $Y=1.46 $X2=0 $Y2=0
cc_141 N_A1_M1006_g N_A_300_51#_c_286_n 0.0113432f $X=2.385 $Y=0.675 $X2=0 $Y2=0
cc_142 N_X_c_199_n N_VPWR_c_219_n 0.0321484f $X=0.45 $Y=1.98 $X2=0 $Y2=0
cc_143 N_X_M1002_s N_VPWR_c_214_n 0.00371702f $X=0.325 $Y=1.835 $X2=0 $Y2=0
cc_144 N_X_c_199_n N_VPWR_c_214_n 0.017806f $X=0.45 $Y=1.98 $X2=0 $Y2=0
cc_145 N_X_c_196_n N_VGND_c_251_n 0.018528f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_146 N_X_M1003_s N_VGND_c_254_n 0.00371702f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_147 N_X_c_196_n N_VGND_c_254_n 0.0104192f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_148 N_VPWR_c_214_n A_420_367# 0.00899413f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_149 N_VGND_c_252_n N_A_300_51#_c_283_n 0.015389f $X=1.955 $Y=0 $X2=0 $Y2=0
cc_150 N_VGND_c_254_n N_A_300_51#_c_283_n 0.0103909f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_151 N_VGND_M1000_d N_A_300_51#_c_284_n 0.00290401f $X=1.93 $Y=0.255 $X2=0
+ $Y2=0
cc_152 N_VGND_c_250_n N_A_300_51#_c_284_n 0.0216414f $X=2.12 $Y=0.4 $X2=0 $Y2=0
cc_153 N_VGND_c_253_n N_A_300_51#_c_286_n 0.0196832f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_154 N_VGND_c_254_n N_A_300_51#_c_286_n 0.0119461f $X=2.64 $Y=0 $X2=0 $Y2=0
