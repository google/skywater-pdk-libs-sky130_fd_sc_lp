* File: sky130_fd_sc_lp__or2b_4.pxi.spice
* Created: Fri Aug 28 11:22:34 2020
* 
x_PM_SKY130_FD_SC_LP__OR2B_4%B_N N_B_N_M1008_g N_B_N_c_86_n N_B_N_c_87_n
+ N_B_N_c_88_n N_B_N_M1005_g N_B_N_c_89_n B_N B_N B_N B_N B_N N_B_N_c_91_n
+ PM_SKY130_FD_SC_LP__OR2B_4%B_N
x_PM_SKY130_FD_SC_LP__OR2B_4%A_27_496# N_A_27_496#_M1005_s N_A_27_496#_M1008_s
+ N_A_27_496#_c_120_n N_A_27_496#_c_121_n N_A_27_496#_c_122_n
+ N_A_27_496#_M1013_g N_A_27_496#_M1009_g N_A_27_496#_c_124_n
+ N_A_27_496#_c_128_n N_A_27_496#_c_129_n N_A_27_496#_c_130_n
+ N_A_27_496#_c_125_n N_A_27_496#_c_126_n PM_SKY130_FD_SC_LP__OR2B_4%A_27_496#
x_PM_SKY130_FD_SC_LP__OR2B_4%A N_A_M1001_g N_A_M1000_g A A N_A_c_180_n
+ PM_SKY130_FD_SC_LP__OR2B_4%A
x_PM_SKY130_FD_SC_LP__OR2B_4%A_256_367# N_A_256_367#_M1013_d
+ N_A_256_367#_M1009_s N_A_256_367#_M1002_g N_A_256_367#_M1003_g
+ N_A_256_367#_M1004_g N_A_256_367#_M1006_g N_A_256_367#_M1007_g
+ N_A_256_367#_M1010_g N_A_256_367#_M1012_g N_A_256_367#_M1011_g
+ N_A_256_367#_c_224_n N_A_256_367#_c_214_n N_A_256_367#_c_215_n
+ N_A_256_367#_c_307_p N_A_256_367#_c_216_n N_A_256_367#_c_281_p
+ N_A_256_367#_c_225_n N_A_256_367#_c_217_n N_A_256_367#_c_218_n
+ N_A_256_367#_c_219_n PM_SKY130_FD_SC_LP__OR2B_4%A_256_367#
x_PM_SKY130_FD_SC_LP__OR2B_4%VPWR N_VPWR_M1008_d N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_M1011_d N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n
+ N_VPWR_c_331_n VPWR N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n
+ N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_326_n
+ PM_SKY130_FD_SC_LP__OR2B_4%VPWR
x_PM_SKY130_FD_SC_LP__OR2B_4%X N_X_M1002_s N_X_M1007_s N_X_M1003_s N_X_M1010_s
+ N_X_c_401_n N_X_c_402_n N_X_c_394_n N_X_c_395_n N_X_c_388_n N_X_c_389_n
+ N_X_c_449_p N_X_c_434_n N_X_c_390_n N_X_c_396_n N_X_c_391_n N_X_c_397_n X X
+ N_X_c_392_n X PM_SKY130_FD_SC_LP__OR2B_4%X
x_PM_SKY130_FD_SC_LP__OR2B_4%VGND N_VGND_M1005_d N_VGND_M1000_d N_VGND_M1004_d
+ N_VGND_M1012_d N_VGND_c_456_n N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n
+ N_VGND_c_460_n N_VGND_c_461_n N_VGND_c_462_n N_VGND_c_463_n VGND
+ N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n N_VGND_c_467_n N_VGND_c_468_n
+ PM_SKY130_FD_SC_LP__OR2B_4%VGND
cc_1 VNB N_B_N_M1008_g 0.0135687f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.69
cc_2 VNB N_B_N_c_86_n 0.0428381f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.84
cc_3 VNB N_B_N_c_87_n 0.0190047f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.84
cc_4 VNB N_B_N_c_88_n 0.0210342f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=0.765
cc_5 VNB N_B_N_c_89_n 0.0185695f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.435
cc_6 VNB B_N 0.0648575f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_7 VNB N_B_N_c_91_n 0.030432f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.93
cc_8 VNB N_A_27_496#_c_120_n 0.0275773f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=0.765
cc_9 VNB N_A_27_496#_c_121_n 0.0117531f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=0.445
cc_10 VNB N_A_27_496#_c_122_n 0.0172423f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=0.445
cc_11 VNB N_A_27_496#_M1009_g 0.0160131f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_12 VNB N_A_27_496#_c_124_n 0.00492991f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_13 VNB N_A_27_496#_c_125_n 0.0141557f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.555
cc_14 VNB N_A_27_496#_c_126_n 0.0219686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_M1000_g 0.0238309f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=0.765
cc_16 VNB A 0.00408839f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.915
cc_17 VNB N_A_c_180_n 0.0225315f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_18 VNB N_A_256_367#_M1002_g 0.0227881f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=0.445
cc_19 VNB N_A_256_367#_M1004_g 0.0228084f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_20 VNB N_A_256_367#_M1007_g 0.0221553f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.93
cc_21 VNB N_A_256_367#_M1012_g 0.0270724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_256_367#_c_214_n 0.00311076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_256_367#_c_215_n 0.00127835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_256_367#_c_216_n 0.0111739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_256_367#_c_217_n 0.00502187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_256_367#_c_218_n 0.00190721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_256_367#_c_219_n 0.0699449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_326_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_388_n 0.00124517f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.93
cc_30 VNB N_X_c_389_n 0.00143437f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.555
cc_31 VNB N_X_c_390_n 0.00141276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_391_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_X_c_392_n 0.0106703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.0212534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_456_n 0.00490645f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_36 VNB N_VGND_c_457_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_37 VNB N_VGND_c_458_n 0.00395069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_459_n 3.20903e-19 $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.93
cc_39 VNB N_VGND_c_460_n 0.0114821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_461_n 0.0284267f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.925
cc_41 VNB N_VGND_c_462_n 0.0344047f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.93
cc_42 VNB N_VGND_c_463_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.295
cc_43 VNB N_VGND_c_464_n 0.0148023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_465_n 0.0123119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_466_n 0.00509388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_467_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_468_n 0.236038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_B_N_M1008_g 0.073891f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.69
cc_49 VPB B_N 0.0240169f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.47
cc_50 VPB N_A_27_496#_M1009_g 0.0221505f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_51 VPB N_A_27_496#_c_128_n 0.0194778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_27_496#_c_129_n 0.0167267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_27_496#_c_130_n 0.0101234f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.93
cc_54 VPB N_A_27_496#_c_125_n 0.0110802f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=0.555
cc_55 VPB N_A_27_496#_c_126_n 0.0251934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_M1001_g 0.0186951f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.69
cc_57 VPB A 0.0117617f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.915
cc_58 VPB N_A_c_180_n 0.00624994f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_59 VPB N_A_256_367#_M1003_g 0.0203177f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.47
cc_60 VPB N_A_256_367#_M1006_g 0.0183529f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_256_367#_M1010_g 0.0183339f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=0.925
cc_62 VPB N_A_256_367#_M1011_g 0.0218662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_256_367#_c_224_n 0.0122559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_256_367#_c_225_n 0.00159279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_256_367#_c_217_n 0.00426239f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_256_367#_c_219_n 0.00893359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_327_n 0.0135098f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_68 VPB N_VPWR_c_328_n 0.00495041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_329_n 3.19317e-19 $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.93
cc_70 VPB N_VPWR_c_330_n 0.0114562f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=0.925
cc_71 VPB N_VPWR_c_331_n 0.0399019f $X=-0.19 $Y=1.655 $X2=0.315 $Y2=0.93
cc_72 VPB N_VPWR_c_332_n 0.0170758f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_333_n 0.0357051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_334_n 0.0152106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_335_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_336_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_337_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_338_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_326_n 0.0612066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_X_c_394_n 0.00305125f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.93
cc_81 VPB N_X_c_395_n 0.00181435f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.93
cc_82 VPB N_X_c_396_n 0.0119296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_X_c_397_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB X 0.00517784f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 N_B_N_c_86_n N_A_27_496#_c_121_n 0.0203744f $X=1.02 $Y=0.84 $X2=0 $Y2=0
cc_86 B_N N_A_27_496#_c_121_n 7.228e-19 $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_87 N_B_N_c_91_n N_A_27_496#_c_121_n 0.0170216f $X=0.385 $Y=0.93 $X2=0 $Y2=0
cc_88 N_B_N_c_88_n N_A_27_496#_c_122_n 0.0132213f $X=1.095 $Y=0.765 $X2=0 $Y2=0
cc_89 N_B_N_M1008_g N_A_27_496#_c_128_n 0.00128436f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_90 N_B_N_M1008_g N_A_27_496#_c_129_n 0.0150408f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_91 B_N N_A_27_496#_c_129_n 0.0147321f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_92 B_N N_A_27_496#_c_130_n 0.0241802f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_93 N_B_N_c_86_n N_A_27_496#_c_125_n 0.0196235f $X=1.02 $Y=0.84 $X2=0 $Y2=0
cc_94 N_B_N_c_88_n N_A_27_496#_c_125_n 0.00833452f $X=1.095 $Y=0.765 $X2=0 $Y2=0
cc_95 B_N N_A_27_496#_c_125_n 0.150105f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_96 N_B_N_c_91_n N_A_27_496#_c_125_n 0.0217035f $X=0.385 $Y=0.93 $X2=0 $Y2=0
cc_97 N_B_N_c_89_n N_A_27_496#_c_126_n 0.0170216f $X=0.385 $Y=1.435 $X2=0 $Y2=0
cc_98 N_B_N_M1008_g N_A_256_367#_c_224_n 0.00436065f $X=0.475 $Y=2.69 $X2=0
+ $Y2=0
cc_99 N_B_N_M1008_g N_A_256_367#_c_217_n 5.11241e-19 $X=0.475 $Y=2.69 $X2=0
+ $Y2=0
cc_100 N_B_N_M1008_g N_VPWR_c_327_n 0.011375f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_101 N_B_N_M1008_g N_VPWR_c_332_n 0.00444095f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_102 N_B_N_M1008_g N_VPWR_c_326_n 0.00442501f $X=0.475 $Y=2.69 $X2=0 $Y2=0
cc_103 N_B_N_c_88_n N_VGND_c_456_n 0.00941374f $X=1.095 $Y=0.765 $X2=0 $Y2=0
cc_104 N_B_N_c_86_n N_VGND_c_462_n 6.70861e-19 $X=1.02 $Y=0.84 $X2=0 $Y2=0
cc_105 N_B_N_c_87_n N_VGND_c_462_n 0.00342052f $X=0.55 $Y=0.84 $X2=0 $Y2=0
cc_106 N_B_N_c_88_n N_VGND_c_462_n 0.0054895f $X=1.095 $Y=0.765 $X2=0 $Y2=0
cc_107 B_N N_VGND_c_462_n 0.0261847f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_108 N_B_N_c_87_n N_VGND_c_468_n 0.00368553f $X=0.55 $Y=0.84 $X2=0 $Y2=0
cc_109 N_B_N_c_88_n N_VGND_c_468_n 0.0116582f $X=1.095 $Y=0.765 $X2=0 $Y2=0
cc_110 B_N N_VGND_c_468_n 0.0174527f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_111 N_A_27_496#_c_122_n N_A_M1000_g 0.0235752f $X=1.62 $Y=1.185 $X2=0 $Y2=0
cc_112 N_A_27_496#_M1009_g A 0.0151439f $X=1.62 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_27_496#_M1009_g N_A_c_180_n 0.113303f $X=1.62 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A_27_496#_M1009_g N_A_256_367#_c_224_n 0.0190402f $X=1.62 $Y=2.465
+ $X2=0 $Y2=0
cc_115 N_A_27_496#_c_129_n N_A_256_367#_c_224_n 0.0136484f $X=0.715 $Y=2.385
+ $X2=0 $Y2=0
cc_116 N_A_27_496#_c_120_n N_A_256_367#_c_214_n 0.00622278f $X=1.545 $Y=1.26
+ $X2=0 $Y2=0
cc_117 N_A_27_496#_c_122_n N_A_256_367#_c_214_n 0.0109058f $X=1.62 $Y=1.185
+ $X2=0 $Y2=0
cc_118 N_A_27_496#_c_124_n N_A_256_367#_c_214_n 0.00470611f $X=1.62 $Y=1.26
+ $X2=0 $Y2=0
cc_119 N_A_27_496#_c_120_n N_A_256_367#_c_215_n 0.0050835f $X=1.545 $Y=1.26
+ $X2=0 $Y2=0
cc_120 N_A_27_496#_c_125_n N_A_256_367#_c_215_n 0.0138345f $X=0.88 $Y=0.44 $X2=0
+ $Y2=0
cc_121 N_A_27_496#_c_120_n N_A_256_367#_c_225_n 6.30113e-19 $X=1.545 $Y=1.26
+ $X2=0 $Y2=0
cc_122 N_A_27_496#_M1009_g N_A_256_367#_c_225_n 0.00342165f $X=1.62 $Y=2.465
+ $X2=0 $Y2=0
cc_123 N_A_27_496#_c_120_n N_A_256_367#_c_217_n 0.00800138f $X=1.545 $Y=1.26
+ $X2=0 $Y2=0
cc_124 N_A_27_496#_M1009_g N_A_256_367#_c_217_n 0.00824141f $X=1.62 $Y=2.465
+ $X2=0 $Y2=0
cc_125 N_A_27_496#_c_125_n N_A_256_367#_c_217_n 0.07367f $X=0.88 $Y=0.44 $X2=0
+ $Y2=0
cc_126 N_A_27_496#_c_126_n N_A_256_367#_c_217_n 0.00472456f $X=0.955 $Y=1.35
+ $X2=0 $Y2=0
cc_127 N_A_27_496#_M1009_g N_VPWR_c_327_n 0.00269103f $X=1.62 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_A_27_496#_c_128_n N_VPWR_c_327_n 0.0108805f $X=0.26 $Y=2.69 $X2=0 $Y2=0
cc_129 N_A_27_496#_c_129_n N_VPWR_c_327_n 0.0250281f $X=0.715 $Y=2.385 $X2=0
+ $Y2=0
cc_130 N_A_27_496#_c_128_n N_VPWR_c_332_n 0.00905291f $X=0.26 $Y=2.69 $X2=0
+ $Y2=0
cc_131 N_A_27_496#_M1009_g N_VPWR_c_333_n 0.0054895f $X=1.62 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_A_27_496#_M1009_g N_VPWR_c_326_n 0.0111524f $X=1.62 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_27_496#_c_128_n N_VPWR_c_326_n 0.00911154f $X=0.26 $Y=2.69 $X2=0
+ $Y2=0
cc_134 N_A_27_496#_c_129_n N_VPWR_c_326_n 0.0138391f $X=0.715 $Y=2.385 $X2=0
+ $Y2=0
cc_135 N_A_27_496#_c_120_n N_VGND_c_456_n 0.0017068f $X=1.545 $Y=1.26 $X2=0
+ $Y2=0
cc_136 N_A_27_496#_c_122_n N_VGND_c_456_n 0.01154f $X=1.62 $Y=1.185 $X2=0 $Y2=0
cc_137 N_A_27_496#_c_125_n N_VGND_c_456_n 0.0457501f $X=0.88 $Y=0.44 $X2=0 $Y2=0
cc_138 N_A_27_496#_c_122_n N_VGND_c_457_n 0.00486043f $X=1.62 $Y=1.185 $X2=0
+ $Y2=0
cc_139 N_A_27_496#_c_125_n N_VGND_c_462_n 0.0210467f $X=0.88 $Y=0.44 $X2=0 $Y2=0
cc_140 N_A_27_496#_M1005_s N_VGND_c_468_n 0.00215158f $X=0.755 $Y=0.235 $X2=0
+ $Y2=0
cc_141 N_A_27_496#_c_122_n N_VGND_c_468_n 0.0082726f $X=1.62 $Y=1.185 $X2=0
+ $Y2=0
cc_142 N_A_27_496#_c_125_n N_VGND_c_468_n 0.0125689f $X=0.88 $Y=0.44 $X2=0 $Y2=0
cc_143 N_A_M1000_g N_A_256_367#_M1002_g 0.0215783f $X=2.05 $Y=0.655 $X2=0 $Y2=0
cc_144 N_A_M1001_g N_A_256_367#_M1003_g 0.0249719f $X=1.98 $Y=2.465 $X2=0 $Y2=0
cc_145 A N_A_256_367#_c_214_n 0.0114468f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A_M1000_g N_A_256_367#_c_216_n 0.0163062f $X=2.05 $Y=0.655 $X2=0 $Y2=0
cc_147 A N_A_256_367#_c_216_n 0.0364541f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A_c_180_n N_A_256_367#_c_216_n 0.0037626f $X=2.07 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A_M1001_g N_A_256_367#_c_225_n 0.00320303f $X=1.98 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_M1000_g N_A_256_367#_c_217_n 2.97897e-19 $X=2.05 $Y=0.655 $X2=0 $Y2=0
cc_151 A N_A_256_367#_c_217_n 0.0266975f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_152 A N_A_256_367#_c_218_n 0.0196765f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_153 N_A_c_180_n N_A_256_367#_c_218_n 0.00179872f $X=2.07 $Y=1.51 $X2=0 $Y2=0
cc_154 A N_A_256_367#_c_219_n 0.00592858f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A_c_180_n N_A_256_367#_c_219_n 0.0222569f $X=2.07 $Y=1.51 $X2=0 $Y2=0
cc_156 N_A_M1001_g N_VPWR_c_328_n 0.00417327f $X=1.98 $Y=2.465 $X2=0 $Y2=0
cc_157 A N_VPWR_c_328_n 0.0154451f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A_c_180_n N_VPWR_c_328_n 8.99119e-19 $X=2.07 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A_M1001_g N_VPWR_c_333_n 0.00585385f $X=1.98 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A_M1001_g N_VPWR_c_326_n 0.0107707f $X=1.98 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A_M1001_g N_X_c_395_n 5.50387e-19 $X=1.98 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_M1000_g N_VGND_c_456_n 6.48031e-19 $X=2.05 $Y=0.655 $X2=0 $Y2=0
cc_163 N_A_M1000_g N_VGND_c_457_n 0.00585385f $X=2.05 $Y=0.655 $X2=0 $Y2=0
cc_164 N_A_M1000_g N_VGND_c_458_n 0.00165353f $X=2.05 $Y=0.655 $X2=0 $Y2=0
cc_165 N_A_M1000_g N_VGND_c_468_n 0.0106668f $X=2.05 $Y=0.655 $X2=0 $Y2=0
cc_166 N_A_256_367#_c_224_n N_VPWR_c_327_n 0.0205913f $X=1.405 $Y=2.95 $X2=0
+ $Y2=0
cc_167 N_A_256_367#_M1003_g N_VPWR_c_328_n 0.00849287f $X=2.52 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_256_367#_c_216_n N_VPWR_c_328_n 0.00373213f $X=2.445 $Y=1.165 $X2=0
+ $Y2=0
cc_169 N_A_256_367#_M1003_g N_VPWR_c_329_n 8.13809e-19 $X=2.52 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_256_367#_M1006_g N_VPWR_c_329_n 0.0141531f $X=2.95 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_256_367#_M1010_g N_VPWR_c_329_n 0.0140168f $X=3.38 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_256_367#_M1011_g N_VPWR_c_329_n 7.21513e-19 $X=3.81 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_256_367#_M1010_g N_VPWR_c_331_n 7.21513e-19 $X=3.38 $Y=2.465 $X2=0
+ $Y2=0
cc_174 N_A_256_367#_M1011_g N_VPWR_c_331_n 0.0150803f $X=3.81 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A_256_367#_c_224_n N_VPWR_c_333_n 0.0210467f $X=1.405 $Y=2.95 $X2=0
+ $Y2=0
cc_176 N_A_256_367#_M1003_g N_VPWR_c_334_n 0.00564131f $X=2.52 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_256_367#_M1006_g N_VPWR_c_334_n 0.00486043f $X=2.95 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_256_367#_M1010_g N_VPWR_c_335_n 0.00486043f $X=3.38 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A_256_367#_M1011_g N_VPWR_c_335_n 0.00486043f $X=3.81 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_256_367#_M1009_s N_VPWR_c_326_n 0.00215158f $X=1.28 $Y=1.835 $X2=0
+ $Y2=0
cc_181 N_A_256_367#_M1003_g N_VPWR_c_326_n 0.0105044f $X=2.52 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_256_367#_M1006_g N_VPWR_c_326_n 0.00824727f $X=2.95 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_256_367#_M1010_g N_VPWR_c_326_n 0.00824727f $X=3.38 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_256_367#_M1011_g N_VPWR_c_326_n 0.00824727f $X=3.81 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A_256_367#_c_224_n N_VPWR_c_326_n 0.0125689f $X=1.405 $Y=2.95 $X2=0
+ $Y2=0
cc_186 N_A_256_367#_c_216_n N_X_M1002_s 0.0021281f $X=2.445 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_256_367#_M1002_g N_X_c_401_n 0.00516273f $X=2.52 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A_256_367#_M1003_g N_X_c_402_n 0.0123379f $X=2.52 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_256_367#_M1006_g N_X_c_394_n 0.013815f $X=2.95 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A_256_367#_M1010_g N_X_c_394_n 0.013815f $X=3.38 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_256_367#_c_281_p N_X_c_394_n 0.0471383f $X=3.63 $Y=1.5 $X2=0 $Y2=0
cc_192 N_A_256_367#_c_219_n N_X_c_394_n 0.00247143f $X=3.81 $Y=1.5 $X2=0 $Y2=0
cc_193 N_A_256_367#_M1003_g N_X_c_395_n 0.0048798f $X=2.52 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A_256_367#_c_216_n N_X_c_395_n 0.0181878f $X=2.445 $Y=1.165 $X2=0 $Y2=0
cc_195 N_A_256_367#_c_281_p N_X_c_395_n 0.00322815f $X=3.63 $Y=1.5 $X2=0 $Y2=0
cc_196 N_A_256_367#_c_219_n N_X_c_395_n 0.00256564f $X=3.81 $Y=1.5 $X2=0 $Y2=0
cc_197 N_A_256_367#_M1007_g N_X_c_388_n 0.0208725f $X=3.38 $Y=0.655 $X2=0 $Y2=0
cc_198 N_A_256_367#_c_281_p N_X_c_388_n 0.0215884f $X=3.63 $Y=1.5 $X2=0 $Y2=0
cc_199 N_A_256_367#_M1002_g N_X_c_389_n 0.0028386f $X=2.52 $Y=0.655 $X2=0 $Y2=0
cc_200 N_A_256_367#_M1004_g N_X_c_389_n 0.0209959f $X=2.95 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A_256_367#_c_216_n N_X_c_389_n 0.0308492f $X=2.445 $Y=1.165 $X2=0 $Y2=0
cc_202 N_A_256_367#_c_281_p N_X_c_389_n 0.0238597f $X=3.63 $Y=1.5 $X2=0 $Y2=0
cc_203 N_A_256_367#_c_219_n N_X_c_389_n 0.00298151f $X=3.81 $Y=1.5 $X2=0 $Y2=0
cc_204 N_A_256_367#_M1012_g N_X_c_390_n 0.0171311f $X=3.81 $Y=0.655 $X2=0 $Y2=0
cc_205 N_A_256_367#_c_281_p N_X_c_390_n 0.00728094f $X=3.63 $Y=1.5 $X2=0 $Y2=0
cc_206 N_A_256_367#_M1011_g N_X_c_396_n 0.0164342f $X=3.81 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_256_367#_c_281_p N_X_c_396_n 0.00731186f $X=3.63 $Y=1.5 $X2=0 $Y2=0
cc_208 N_A_256_367#_c_281_p N_X_c_391_n 0.0153308f $X=3.63 $Y=1.5 $X2=0 $Y2=0
cc_209 N_A_256_367#_c_219_n N_X_c_391_n 0.00256759f $X=3.81 $Y=1.5 $X2=0 $Y2=0
cc_210 N_A_256_367#_c_281_p N_X_c_397_n 0.0153308f $X=3.63 $Y=1.5 $X2=0 $Y2=0
cc_211 N_A_256_367#_c_219_n N_X_c_397_n 0.00256759f $X=3.81 $Y=1.5 $X2=0 $Y2=0
cc_212 N_A_256_367#_M1012_g X 0.0198363f $X=3.81 $Y=0.655 $X2=0 $Y2=0
cc_213 N_A_256_367#_c_281_p X 0.0138862f $X=3.63 $Y=1.5 $X2=0 $Y2=0
cc_214 N_A_256_367#_c_215_n N_VGND_M1005_d 0.00149394f $X=1.415 $Y=1.165
+ $X2=-0.19 $Y2=-0.245
cc_215 N_A_256_367#_c_214_n N_VGND_c_456_n 0.00998943f $X=1.74 $Y=1.165 $X2=0
+ $Y2=0
cc_216 N_A_256_367#_c_215_n N_VGND_c_456_n 0.0158256f $X=1.415 $Y=1.165 $X2=0
+ $Y2=0
cc_217 N_A_256_367#_c_307_p N_VGND_c_457_n 0.0136943f $X=1.835 $Y=0.42 $X2=0
+ $Y2=0
cc_218 N_A_256_367#_M1002_g N_VGND_c_458_n 0.00155098f $X=2.52 $Y=0.655 $X2=0
+ $Y2=0
cc_219 N_A_256_367#_c_216_n N_VGND_c_458_n 0.0192759f $X=2.445 $Y=1.165 $X2=0
+ $Y2=0
cc_220 N_A_256_367#_M1002_g N_VGND_c_459_n 4.78045e-19 $X=2.52 $Y=0.655 $X2=0
+ $Y2=0
cc_221 N_A_256_367#_M1004_g N_VGND_c_459_n 0.00779775f $X=2.95 $Y=0.655 $X2=0
+ $Y2=0
cc_222 N_A_256_367#_M1007_g N_VGND_c_459_n 0.00764057f $X=3.38 $Y=0.655 $X2=0
+ $Y2=0
cc_223 N_A_256_367#_M1012_g N_VGND_c_459_n 5.37623e-19 $X=3.81 $Y=0.655 $X2=0
+ $Y2=0
cc_224 N_A_256_367#_M1007_g N_VGND_c_461_n 5.85999e-19 $X=3.38 $Y=0.655 $X2=0
+ $Y2=0
cc_225 N_A_256_367#_M1012_g N_VGND_c_461_n 0.0126465f $X=3.81 $Y=0.655 $X2=0
+ $Y2=0
cc_226 N_A_256_367#_M1002_g N_VGND_c_464_n 0.0054895f $X=2.52 $Y=0.655 $X2=0
+ $Y2=0
cc_227 N_A_256_367#_M1004_g N_VGND_c_464_n 0.00365091f $X=2.95 $Y=0.655 $X2=0
+ $Y2=0
cc_228 N_A_256_367#_M1007_g N_VGND_c_465_n 0.00365202f $X=3.38 $Y=0.655 $X2=0
+ $Y2=0
cc_229 N_A_256_367#_M1012_g N_VGND_c_465_n 0.00486043f $X=3.81 $Y=0.655 $X2=0
+ $Y2=0
cc_230 N_A_256_367#_M1013_d N_VGND_c_468_n 0.0041489f $X=1.695 $Y=0.235 $X2=0
+ $Y2=0
cc_231 N_A_256_367#_M1002_g N_VGND_c_468_n 0.00988472f $X=2.52 $Y=0.655 $X2=0
+ $Y2=0
cc_232 N_A_256_367#_M1004_g N_VGND_c_468_n 0.00432036f $X=2.95 $Y=0.655 $X2=0
+ $Y2=0
cc_233 N_A_256_367#_M1007_g N_VGND_c_468_n 0.00432244f $X=3.38 $Y=0.655 $X2=0
+ $Y2=0
cc_234 N_A_256_367#_M1012_g N_VGND_c_468_n 0.00824727f $X=3.81 $Y=0.655 $X2=0
+ $Y2=0
cc_235 N_A_256_367#_c_307_p N_VGND_c_468_n 0.00866972f $X=1.835 $Y=0.42 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_326_n A_339_367# 0.00899413f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_237 N_VPWR_c_326_n N_X_M1003_s 0.00380103f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_238 N_VPWR_c_326_n N_X_M1010_s 0.00536646f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_c_334_n N_X_c_402_n 0.0150063f $X=3 $Y=3.33 $X2=0 $Y2=0
cc_240 N_VPWR_c_326_n N_X_c_402_n 0.00950443f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_241 N_VPWR_M1006_d N_X_c_394_n 0.00177068f $X=3.025 $Y=1.835 $X2=0 $Y2=0
cc_242 N_VPWR_c_329_n N_X_c_394_n 0.0172078f $X=3.165 $Y=2.2 $X2=0 $Y2=0
cc_243 N_VPWR_c_335_n N_X_c_434_n 0.0124525f $X=3.86 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_326_n N_X_c_434_n 0.00730901f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_M1011_d N_X_c_396_n 0.00314254f $X=3.885 $Y=1.835 $X2=0 $Y2=0
cc_246 N_VPWR_c_331_n N_X_c_396_n 0.0239119f $X=4.025 $Y=2.2 $X2=0 $Y2=0
cc_247 N_X_c_388_n N_VGND_M1004_d 3.43519e-19 $X=3.5 $Y=0.99 $X2=0 $Y2=0
cc_248 N_X_c_389_n N_VGND_M1004_d 0.00142435f $X=3.215 $Y=0.99 $X2=0 $Y2=0
cc_249 N_X_c_390_n N_VGND_M1012_d 2.34277e-19 $X=3.965 $Y=1.155 $X2=0 $Y2=0
cc_250 N_X_c_392_n N_VGND_M1012_d 0.0020943f $X=4.1 $Y=1.245 $X2=0 $Y2=0
cc_251 N_X_c_388_n N_VGND_c_459_n 0.00460669f $X=3.5 $Y=0.99 $X2=0 $Y2=0
cc_252 N_X_c_389_n N_VGND_c_459_n 0.0131604f $X=3.215 $Y=0.99 $X2=0 $Y2=0
cc_253 N_X_c_390_n N_VGND_c_461_n 0.00363499f $X=3.965 $Y=1.155 $X2=0 $Y2=0
cc_254 N_X_c_392_n N_VGND_c_461_n 0.0203341f $X=4.1 $Y=1.245 $X2=0 $Y2=0
cc_255 N_X_c_401_n N_VGND_c_464_n 0.0156443f $X=2.735 $Y=0.42 $X2=0 $Y2=0
cc_256 N_X_c_389_n N_VGND_c_464_n 0.00200795f $X=3.215 $Y=0.99 $X2=0 $Y2=0
cc_257 N_X_c_388_n N_VGND_c_465_n 0.0020876f $X=3.5 $Y=0.99 $X2=0 $Y2=0
cc_258 N_X_c_449_p N_VGND_c_465_n 0.0124525f $X=3.595 $Y=0.42 $X2=0 $Y2=0
cc_259 N_X_M1002_s N_VGND_c_468_n 0.00244952f $X=2.595 $Y=0.235 $X2=0 $Y2=0
cc_260 N_X_M1007_s N_VGND_c_468_n 0.00401561f $X=3.455 $Y=0.235 $X2=0 $Y2=0
cc_261 N_X_c_401_n N_VGND_c_468_n 0.00983564f $X=2.735 $Y=0.42 $X2=0 $Y2=0
cc_262 N_X_c_388_n N_VGND_c_468_n 0.00451994f $X=3.5 $Y=0.99 $X2=0 $Y2=0
cc_263 N_X_c_389_n N_VGND_c_468_n 0.00478653f $X=3.215 $Y=0.99 $X2=0 $Y2=0
cc_264 N_X_c_449_p N_VGND_c_468_n 0.00730901f $X=3.595 $Y=0.42 $X2=0 $Y2=0
