* File: sky130_fd_sc_lp__einvn_1.pxi.spice
* Created: Wed Sep  2 09:51:32 2020
* 
x_PM_SKY130_FD_SC_LP__EINVN_1%A N_A_M1000_g N_A_M1004_g A A N_A_c_46_n
+ N_A_c_47_n PM_SKY130_FD_SC_LP__EINVN_1%A
x_PM_SKY130_FD_SC_LP__EINVN_1%A_214_21# N_A_214_21#_M1002_d N_A_214_21#_M1003_d
+ N_A_214_21#_c_73_n N_A_214_21#_M1001_g N_A_214_21#_c_74_n N_A_214_21#_c_75_n
+ N_A_214_21#_c_76_n N_A_214_21#_c_77_n N_A_214_21#_c_81_n N_A_214_21#_c_78_n
+ N_A_214_21#_c_79_n N_A_214_21#_c_80_n PM_SKY130_FD_SC_LP__EINVN_1%A_214_21#
x_PM_SKY130_FD_SC_LP__EINVN_1%TE_B N_TE_B_c_124_n N_TE_B_M1005_g N_TE_B_c_119_n
+ N_TE_B_c_120_n N_TE_B_M1003_g N_TE_B_M1002_g TE_B TE_B N_TE_B_c_121_n
+ N_TE_B_c_122_n N_TE_B_c_123_n PM_SKY130_FD_SC_LP__EINVN_1%TE_B
x_PM_SKY130_FD_SC_LP__EINVN_1%Z N_Z_M1000_s N_Z_M1004_s N_Z_c_164_n N_Z_c_165_n
+ Z Z Z PM_SKY130_FD_SC_LP__EINVN_1%Z
x_PM_SKY130_FD_SC_LP__EINVN_1%VPWR N_VPWR_M1005_d N_VPWR_c_193_n VPWR
+ N_VPWR_c_194_n N_VPWR_c_195_n N_VPWR_c_192_n N_VPWR_c_197_n
+ PM_SKY130_FD_SC_LP__EINVN_1%VPWR
x_PM_SKY130_FD_SC_LP__EINVN_1%VGND N_VGND_M1001_d N_VGND_c_216_n N_VGND_c_217_n
+ VGND N_VGND_c_218_n N_VGND_c_219_n N_VGND_c_220_n N_VGND_c_221_n
+ PM_SKY130_FD_SC_LP__EINVN_1%VGND
cc_1 VNB N_A_M1004_g 5.05655e-19 $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=2.465
cc_2 VNB A 0.0136979f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_c_46_n 0.0371628f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.48
cc_4 VNB N_A_c_47_n 0.0211217f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.315
cc_5 VNB N_A_214_21#_c_73_n 0.0156157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_214_21#_c_74_n 0.038094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_214_21#_c_75_n 0.012053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_214_21#_c_76_n 0.0222535f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.48
cc_9 VNB N_A_214_21#_c_77_n 0.0185554f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.295
cc_10 VNB N_A_214_21#_c_78_n 0.0187527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_214_21#_c_79_n 0.00869653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_214_21#_c_80_n 0.0551115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_TE_B_c_119_n 0.0164431f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.645
cc_14 VNB N_TE_B_c_120_n 0.00454679f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=2.465
cc_15 VNB N_TE_B_c_121_n 0.0254429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_TE_B_c_122_n 0.00769637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_TE_B_c_123_n 0.0203969f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.48
cc_18 VNB N_Z_c_164_n 0.0256113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Z_c_165_n 0.016666f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_20 VNB Z 0.0329116f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.645
cc_21 VNB N_VPWR_c_192_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.48
cc_22 VNB N_VGND_c_216_n 0.00616313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_217_n 0.00358244f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_24 VNB N_VGND_c_218_n 0.0353989f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.48
cc_25 VNB N_VGND_c_219_n 0.0213186f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.665
cc_26 VNB N_VGND_c_220_n 0.163899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_221_n 0.00552652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A_M1004_g 0.0234701f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=2.465
cc_29 VPB A 0.00390908f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_30 VPB N_A_214_21#_c_81_n 0.040636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_A_214_21#_c_78_n 0.0130082f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_TE_B_c_124_n 0.0181941f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=1.315
cc_33 VPB N_TE_B_c_119_n 0.0147111f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=1.645
cc_34 VPB N_TE_B_c_120_n 0.00192443f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=2.465
cc_35 VPB N_TE_B_M1003_g 0.0268688f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_36 VPB N_TE_B_c_121_n 0.0112211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_TE_B_c_122_n 0.00812009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB Z 0.0814773f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.645
cc_39 VPB N_VPWR_c_193_n 0.0218365f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=2.465
cc_40 VPB N_VPWR_c_194_n 0.0313059f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.48
cc_41 VPB N_VPWR_c_195_n 0.0266462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_192_n 0.0566927f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.48
cc_43 VPB N_VPWR_c_197_n 0.00712807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 A N_A_214_21#_c_73_n 0.00108011f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_45 N_A_c_46_n N_A_214_21#_c_73_n 0.0274771f $X=0.665 $Y=1.48 $X2=0 $Y2=0
cc_46 N_A_c_47_n N_A_214_21#_c_75_n 0.0274771f $X=0.665 $Y=1.315 $X2=0 $Y2=0
cc_47 N_A_M1004_g N_TE_B_c_124_n 0.0437446f $X=0.755 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_48 A N_TE_B_c_120_n 7.09338e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_49 N_A_c_46_n N_TE_B_c_120_n 0.0437446f $X=0.665 $Y=1.48 $X2=0 $Y2=0
cc_50 A N_TE_B_c_122_n 0.0217227f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_51 N_A_c_46_n N_TE_B_c_122_n 5.48234e-19 $X=0.665 $Y=1.48 $X2=0 $Y2=0
cc_52 A N_Z_c_164_n 0.0149154f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_53 N_A_c_46_n N_Z_c_164_n 8.98502e-19 $X=0.665 $Y=1.48 $X2=0 $Y2=0
cc_54 N_A_c_47_n N_Z_c_164_n 0.00727845f $X=0.665 $Y=1.315 $X2=0 $Y2=0
cc_55 N_A_c_47_n N_Z_c_165_n 0.00665995f $X=0.665 $Y=1.315 $X2=0 $Y2=0
cc_56 N_A_M1004_g Z 0.0321466f $X=0.755 $Y=2.465 $X2=0 $Y2=0
cc_57 A Z 0.0694891f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_58 N_A_c_46_n Z 0.00839588f $X=0.665 $Y=1.48 $X2=0 $Y2=0
cc_59 N_A_c_47_n Z 0.00398495f $X=0.665 $Y=1.315 $X2=0 $Y2=0
cc_60 N_A_M1004_g N_VPWR_c_193_n 0.0024397f $X=0.755 $Y=2.465 $X2=0 $Y2=0
cc_61 N_A_M1004_g N_VPWR_c_194_n 0.00357668f $X=0.755 $Y=2.465 $X2=0 $Y2=0
cc_62 N_A_M1004_g N_VPWR_c_192_n 0.00638121f $X=0.755 $Y=2.465 $X2=0 $Y2=0
cc_63 N_A_c_47_n N_VGND_c_216_n 0.00337666f $X=0.665 $Y=1.315 $X2=0 $Y2=0
cc_64 A N_VGND_c_217_n 0.00636008f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_c_47_n N_VGND_c_218_n 0.00437175f $X=0.665 $Y=1.315 $X2=0 $Y2=0
cc_66 N_A_c_47_n N_VGND_c_220_n 0.00833596f $X=0.665 $Y=1.315 $X2=0 $Y2=0
cc_67 N_A_214_21#_c_81_n N_TE_B_c_124_n 4.12285e-19 $X=1.965 $Y=2.05 $X2=-0.19
+ $Y2=-0.245
cc_68 N_A_214_21#_c_73_n N_TE_B_c_120_n 0.00996546f $X=1.145 $Y=0.255 $X2=0
+ $Y2=0
cc_69 N_A_214_21#_c_81_n N_TE_B_M1003_g 0.00798072f $X=1.965 $Y=2.05 $X2=0 $Y2=0
cc_70 N_A_214_21#_c_78_n N_TE_B_M1003_g 0.00362222f $X=2.057 $Y=1.92 $X2=0 $Y2=0
cc_71 N_A_214_21#_c_81_n N_TE_B_c_121_n 8.70296e-19 $X=1.965 $Y=2.05 $X2=0 $Y2=0
cc_72 N_A_214_21#_c_78_n N_TE_B_c_121_n 0.00481961f $X=2.057 $Y=1.92 $X2=0 $Y2=0
cc_73 N_A_214_21#_c_73_n N_TE_B_c_122_n 0.00304635f $X=1.145 $Y=0.255 $X2=0
+ $Y2=0
cc_74 N_A_214_21#_c_81_n N_TE_B_c_122_n 0.0107323f $X=1.965 $Y=2.05 $X2=0 $Y2=0
cc_75 N_A_214_21#_c_78_n N_TE_B_c_122_n 0.0203606f $X=2.057 $Y=1.92 $X2=0 $Y2=0
cc_76 N_A_214_21#_c_73_n N_TE_B_c_123_n 0.004307f $X=1.145 $Y=0.255 $X2=0 $Y2=0
cc_77 N_A_214_21#_c_76_n N_TE_B_c_123_n 0.00392777f $X=2.115 $Y=1.07 $X2=0 $Y2=0
cc_78 N_A_214_21#_c_77_n N_TE_B_c_123_n 0.00319798f $X=1.945 $Y=0.38 $X2=0 $Y2=0
cc_79 N_A_214_21#_c_78_n N_TE_B_c_123_n 0.00301791f $X=2.057 $Y=1.92 $X2=0 $Y2=0
cc_80 N_A_214_21#_c_80_n N_TE_B_c_123_n 0.00825427f $X=1.945 $Y=0.18 $X2=0 $Y2=0
cc_81 N_A_214_21#_c_73_n N_Z_c_164_n 9.39754e-19 $X=1.145 $Y=0.255 $X2=0 $Y2=0
cc_82 N_A_214_21#_c_73_n N_Z_c_165_n 0.00101899f $X=1.145 $Y=0.255 $X2=0 $Y2=0
cc_83 N_A_214_21#_c_81_n N_VPWR_c_193_n 0.0267307f $X=1.965 $Y=2.05 $X2=0 $Y2=0
cc_84 N_A_214_21#_c_81_n N_VPWR_c_192_n 0.0214511f $X=1.965 $Y=2.05 $X2=0 $Y2=0
cc_85 N_A_214_21#_c_73_n N_VGND_c_216_n 0.0141561f $X=1.145 $Y=0.255 $X2=0 $Y2=0
cc_86 N_A_214_21#_c_74_n N_VGND_c_216_n 0.023413f $X=1.78 $Y=0.18 $X2=0 $Y2=0
cc_87 N_A_214_21#_c_75_n N_VGND_c_216_n 0.00363588f $X=1.22 $Y=0.18 $X2=0 $Y2=0
cc_88 N_A_214_21#_c_76_n N_VGND_c_216_n 0.0174849f $X=2.115 $Y=1.07 $X2=0 $Y2=0
cc_89 N_A_214_21#_c_77_n N_VGND_c_216_n 0.0308462f $X=1.945 $Y=0.38 $X2=0 $Y2=0
cc_90 N_A_214_21#_c_80_n N_VGND_c_216_n 0.00305668f $X=1.945 $Y=0.18 $X2=0 $Y2=0
cc_91 N_A_214_21#_c_73_n N_VGND_c_217_n 0.0107449f $X=1.145 $Y=0.255 $X2=0 $Y2=0
cc_92 N_A_214_21#_c_78_n N_VGND_c_217_n 2.35244e-19 $X=2.057 $Y=1.92 $X2=0 $Y2=0
cc_93 N_A_214_21#_c_75_n N_VGND_c_218_n 0.00486043f $X=1.22 $Y=0.18 $X2=0 $Y2=0
cc_94 N_A_214_21#_c_74_n N_VGND_c_219_n 0.0138149f $X=1.78 $Y=0.18 $X2=0 $Y2=0
cc_95 N_A_214_21#_c_77_n N_VGND_c_219_n 0.0344292f $X=1.945 $Y=0.38 $X2=0 $Y2=0
cc_96 N_A_214_21#_c_74_n N_VGND_c_220_n 0.00905438f $X=1.78 $Y=0.18 $X2=0 $Y2=0
cc_97 N_A_214_21#_c_75_n N_VGND_c_220_n 0.00972445f $X=1.22 $Y=0.18 $X2=0 $Y2=0
cc_98 N_A_214_21#_c_77_n N_VGND_c_220_n 0.0190261f $X=1.945 $Y=0.38 $X2=0 $Y2=0
cc_99 N_A_214_21#_c_80_n N_VGND_c_220_n 0.00950499f $X=1.945 $Y=0.18 $X2=0 $Y2=0
cc_100 N_TE_B_c_124_n Z 0.00893316f $X=1.145 $Y=1.725 $X2=0 $Y2=0
cc_101 N_TE_B_c_124_n N_VPWR_c_193_n 0.0351187f $X=1.145 $Y=1.725 $X2=0 $Y2=0
cc_102 N_TE_B_c_119_n N_VPWR_c_193_n 0.00285315f $X=1.63 $Y=1.635 $X2=0 $Y2=0
cc_103 N_TE_B_M1003_g N_VPWR_c_193_n 0.00534125f $X=1.75 $Y=2.225 $X2=0 $Y2=0
cc_104 N_TE_B_c_122_n N_VPWR_c_193_n 0.0336302f $X=1.795 $Y=1.58 $X2=0 $Y2=0
cc_105 N_TE_B_c_124_n N_VPWR_c_194_n 0.00486043f $X=1.145 $Y=1.725 $X2=0 $Y2=0
cc_106 N_TE_B_M1003_g N_VPWR_c_195_n 0.00340167f $X=1.75 $Y=2.225 $X2=0 $Y2=0
cc_107 N_TE_B_c_124_n N_VPWR_c_192_n 0.00827383f $X=1.145 $Y=1.725 $X2=0 $Y2=0
cc_108 N_TE_B_M1003_g N_VPWR_c_192_n 0.00427383f $X=1.75 $Y=2.225 $X2=0 $Y2=0
cc_109 N_TE_B_c_123_n N_VGND_c_216_n 0.00242338f $X=1.795 $Y=1.415 $X2=0 $Y2=0
cc_110 N_TE_B_c_119_n N_VGND_c_217_n 0.00285345f $X=1.63 $Y=1.635 $X2=0 $Y2=0
cc_111 N_TE_B_c_121_n N_VGND_c_217_n 0.00315729f $X=1.795 $Y=1.58 $X2=0 $Y2=0
cc_112 N_TE_B_c_122_n N_VGND_c_217_n 0.0463856f $X=1.795 $Y=1.58 $X2=0 $Y2=0
cc_113 N_TE_B_c_123_n N_VGND_c_217_n 5.7783e-19 $X=1.795 $Y=1.415 $X2=0 $Y2=0
cc_114 N_TE_B_c_123_n N_VGND_c_220_n 4.27605e-19 $X=1.795 $Y=1.415 $X2=0 $Y2=0
cc_115 Z A_166_367# 0.0125693f $X=0.155 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_116 Z N_VPWR_c_193_n 0.0618465f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_117 Z N_VPWR_c_194_n 0.0532917f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_118 N_Z_M1004_s N_VPWR_c_192_n 0.00215158f $X=0.415 $Y=1.835 $X2=0 $Y2=0
cc_119 Z N_VPWR_c_192_n 0.030848f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_120 N_Z_c_164_n N_VGND_c_216_n 0.01131f $X=0.54 $Y=0.705 $X2=0 $Y2=0
cc_121 N_Z_c_165_n N_VGND_c_216_n 0.0116086f $X=0.54 $Y=0.51 $X2=0 $Y2=0
cc_122 N_Z_c_164_n N_VGND_c_218_n 0.00485549f $X=0.54 $Y=0.705 $X2=0 $Y2=0
cc_123 N_Z_c_165_n N_VGND_c_218_n 0.0142054f $X=0.54 $Y=0.51 $X2=0 $Y2=0
cc_124 N_Z_c_164_n N_VGND_c_220_n 0.00813131f $X=0.54 $Y=0.705 $X2=0 $Y2=0
cc_125 N_Z_c_165_n N_VGND_c_220_n 0.0117891f $X=0.54 $Y=0.51 $X2=0 $Y2=0
cc_126 A_166_367# N_VPWR_c_192_n 0.00787867f $X=0.83 $Y=1.835 $X2=0 $Y2=0
