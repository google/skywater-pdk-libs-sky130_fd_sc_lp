* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4_0 A B C D VGND VNB VPB VPWR X
X0 VGND a_54_482# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_137_482# C a_227_482# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_54_482# D a_137_482# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_54_482# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND B a_54_482# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_54_482# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_227_482# B a_317_482# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_317_482# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_54_482# X VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VGND D a_54_482# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
