# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux2_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__mux2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 0.345000 1.905000 1.525000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.200000 2.725000 1.525000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.335000 0.690000 1.695000 ;
        RECT 0.430000 1.695000 3.255000 1.865000 ;
        RECT 2.905000 1.200000 3.255000 1.695000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 0.255000 3.975000 1.065000 ;
        RECT 3.765000 1.065000 5.660000 1.235000 ;
        RECT 3.855000 1.755000 5.660000 1.925000 ;
        RECT 3.855000 1.925000 4.045000 3.075000 ;
        RECT 4.645000 0.255000 4.870000 1.065000 ;
        RECT 4.715000 1.925000 4.895000 3.075000 ;
        RECT 5.435000 0.390000 5.660000 1.065000 ;
        RECT 5.460000 1.235000 5.660000 1.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.760000 0.085000 ;
        RECT 0.870000  0.085000 1.330000 0.815000 ;
        RECT 2.875000  0.085000 3.595000 0.690000 ;
        RECT 4.145000  0.085000 4.475000 0.895000 ;
        RECT 5.040000  0.085000 5.265000 0.895000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 5.760000 3.415000 ;
        RECT 0.595000 2.035000 0.925000 3.245000 ;
        RECT 3.355000 2.445000 3.685000 3.245000 ;
        RECT 4.215000 2.095000 4.545000 3.245000 ;
        RECT 5.075000 2.095000 5.405000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.255000 0.700000 0.985000 ;
      RECT 0.090000 0.985000 1.415000 1.155000 ;
      RECT 0.090000 1.155000 0.260000 2.035000 ;
      RECT 0.090000 2.035000 0.425000 3.075000 ;
      RECT 1.085000 1.155000 1.415000 1.525000 ;
      RECT 1.095000 2.035000 1.355000 2.905000 ;
      RECT 1.095000 2.905000 2.735000 3.075000 ;
      RECT 1.545000 2.035000 1.805000 2.505000 ;
      RECT 1.545000 2.505000 3.185000 2.675000 ;
      RECT 1.545000 2.675000 1.795000 2.735000 ;
      RECT 1.975000 2.035000 3.650000 2.215000 ;
      RECT 1.975000 2.215000 2.305000 2.335000 ;
      RECT 2.085000 0.255000 2.530000 0.860000 ;
      RECT 2.085000 0.860000 3.595000 1.030000 ;
      RECT 2.405000 2.845000 2.735000 2.905000 ;
      RECT 2.925000 2.385000 3.185000 2.505000 ;
      RECT 2.925000 2.675000 3.185000 3.075000 ;
      RECT 3.425000 1.030000 3.595000 1.405000 ;
      RECT 3.425000 1.405000 5.280000 1.585000 ;
      RECT 3.425000 1.585000 3.650000 2.035000 ;
  END
END sky130_fd_sc_lp__mux2_4
