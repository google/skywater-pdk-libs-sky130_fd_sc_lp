# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfxtp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfxtp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.170000 2.755000 1.500000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.400500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.595000 0.440000 10.935000 1.780000 ;
        RECT 10.595000 1.780000 10.925000 3.000000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.175000 0.835000 1.845000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 11.040000 0.085000 ;
        RECT 0.895000  0.085000  1.225000 0.645000 ;
        RECT 2.260000  0.085000  2.590000 0.990000 ;
        RECT 6.320000  0.085000  6.570000 0.685000 ;
        RECT 8.545000  0.085000  8.795000 0.815000 ;
        RECT 9.895000  0.085000 10.145000 0.900000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 11.040000 3.415000 ;
        RECT  0.760000 2.025000  1.090000 3.245000 ;
        RECT  2.540000 2.030000  2.870000 3.245000 ;
        RECT  5.360000 2.075000  5.690000 3.245000 ;
        RECT  8.535000 2.105000  8.865000 3.245000 ;
        RECT 10.065000 1.960000 10.395000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.105000 0.265000  0.435000 0.825000 ;
      RECT  0.105000 0.825000  1.495000 0.995000 ;
      RECT  0.105000 0.995000  0.275000 2.025000 ;
      RECT  0.105000 2.025000  0.560000 3.065000 ;
      RECT  1.165000 0.995000  1.495000 1.495000 ;
      RECT  1.290000 2.025000  1.845000 3.065000 ;
      RECT  1.675000 0.265000  2.015000 0.725000 ;
      RECT  1.675000 0.725000  1.845000 1.680000 ;
      RECT  1.675000 1.680000  3.105000 1.850000 ;
      RECT  1.675000 1.850000  1.845000 2.025000 ;
      RECT  2.935000 1.215000  3.645000 1.545000 ;
      RECT  2.935000 1.545000  3.105000 1.680000 ;
      RECT  3.200000 0.375000  3.530000 0.865000 ;
      RECT  3.200000 0.865000  3.995000 1.035000 ;
      RECT  3.285000 1.725000  3.995000 1.895000 ;
      RECT  3.285000 1.895000  3.615000 2.730000 ;
      RECT  3.710000 0.375000  4.345000 0.685000 ;
      RECT  3.825000 1.035000  3.995000 1.725000 ;
      RECT  4.175000 0.685000  4.345000 1.685000 ;
      RECT  4.175000 1.685000  5.065000 1.855000 ;
      RECT  4.175000 1.855000  4.505000 2.875000 ;
      RECT  4.525000 0.455000  6.140000 0.625000 ;
      RECT  4.525000 0.625000  4.715000 1.485000 ;
      RECT  4.895000 0.805000  5.790000 0.975000 ;
      RECT  4.895000 0.975000  5.065000 1.685000 ;
      RECT  5.245000 1.155000  5.440000 1.725000 ;
      RECT  5.245000 1.725000  8.005000 1.895000 ;
      RECT  5.620000 0.975000  5.790000 1.215000 ;
      RECT  5.620000 1.215000  6.330000 1.545000 ;
      RECT  5.970000 0.625000  6.140000 0.865000 ;
      RECT  5.970000 0.865000  6.680000 1.035000 ;
      RECT  6.510000 1.035000  6.680000 1.215000 ;
      RECT  6.510000 1.215000  7.655000 1.385000 ;
      RECT  6.510000 1.685000  6.840000 1.725000 ;
      RECT  6.510000 1.895000  6.840000 2.935000 ;
      RECT  7.115000 0.605000  7.445000 0.865000 ;
      RECT  7.115000 0.865000  8.005000 1.035000 ;
      RECT  7.120000 2.075000  8.355000 2.245000 ;
      RECT  7.120000 2.245000  7.450000 2.935000 ;
      RECT  7.345000 1.385000  7.655000 1.545000 ;
      RECT  7.675000 0.355000  8.355000 0.685000 ;
      RECT  7.835000 1.035000  8.005000 1.725000 ;
      RECT  8.185000 0.685000  8.355000 0.995000 ;
      RECT  8.185000 0.995000  9.365000 1.165000 ;
      RECT  8.185000 1.165000  8.355000 2.075000 ;
      RECT  8.535000 1.425000  8.845000 1.755000 ;
      RECT  8.535000 1.755000  9.720000 1.925000 ;
      RECT  9.055000 0.905000  9.365000 0.995000 ;
      RECT  9.055000 1.165000  9.365000 1.575000 ;
      RECT  9.255000 0.355000  9.715000 0.725000 ;
      RECT  9.390000 1.925000  9.720000 2.935000 ;
      RECT  9.545000 0.725000  9.715000 1.585000 ;
      RECT  9.545000 1.585000 10.415000 1.755000 ;
      RECT 10.085000 1.085000 10.415000 1.585000 ;
  END
END sky130_fd_sc_lp__dfxtp_lp
