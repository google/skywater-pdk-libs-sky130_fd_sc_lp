* File: sky130_fd_sc_lp__a221oi_lp.pex.spice
* Created: Fri Aug 28 09:53:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221OI_LP%B2 3 7 11 14 15 17 24
c36 24 0 2.42909e-19 $X=0.55 $Y=1.275
c37 11 0 1.66743e-19 $X=0.58 $Y=1.26
r38 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.55
+ $Y=1.275 $X2=0.55 $Y2=1.275
r39 17 25 3.03483 $w=6.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.72 $Y=1.445
+ $X2=0.55 $Y2=1.445
r40 15 25 5.53409 $w=6.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.24 $Y=1.445
+ $X2=0.55 $Y2=1.445
r41 13 24 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.55 $Y=1.63
+ $X2=0.55 $Y2=1.275
r42 13 14 29.7575 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.6 $Y=1.63 $X2=0.6
+ $Y2=1.78
r43 11 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.55 $Y=1.26
+ $X2=0.55 $Y2=1.275
r44 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.58 $Y=1.11
+ $X2=0.58 $Y2=1.26
r45 7 10 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.7 $Y=0.45 $X2=0.7
+ $Y2=1.11
r46 3 14 193.794 $w=2.5e-07 $l=7.8e-07 $layer=POLY_cond $X=0.69 $Y=2.56 $X2=0.69
+ $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_LP%B1 3 7 9 12 15 16 17 18 27
c63 9 0 2.37644e-19 $X=1.565 $Y=1.165
r64 27 30 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.54 $Y=1.735
+ $X2=2.54 $Y2=1.9
r65 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.54
+ $Y=1.735 $X2=2.54 $Y2=1.735
r66 18 28 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.64 $Y=1.735 $X2=2.54
+ $Y2=1.735
r67 17 28 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.16 $Y=1.735
+ $X2=2.54 $Y2=1.735
r68 16 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=1.735
+ $X2=1.735 $Y2=1.735
r69 16 17 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.75 $Y=1.735
+ $X2=2.16 $Y2=1.735
r70 16 31 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.75 $Y=1.735
+ $X2=1.735 $Y2=1.735
r71 15 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=1.57
+ $X2=1.65 $Y2=1.735
r72 14 15 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.65 $Y=1.33
+ $X2=1.65 $Y2=1.57
r73 12 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.165
+ $X2=1.18 $Y2=1
r74 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.165 $X2=1.18 $Y2=1.165
r75 9 14 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.165
+ $X2=1.65 $Y2=1.33
r76 9 11 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.565 $Y=1.165
+ $X2=1.18 $Y2=1.165
r77 7 30 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.57 $Y=2.56 $X2=2.57
+ $Y2=1.9
r78 3 24 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.09 $Y=0.45 $X2=1.09
+ $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_LP%A1 3 7 9 15
c43 9 0 3.24915e-19 $X=1.2 $Y=1.665
c44 3 0 1.7238e-19 $X=1.22 $Y=2.56
r45 12 15 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.22 $Y=1.735
+ $X2=1.63 $Y2=1.735
r46 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.735 $X2=1.22 $Y2=1.735
r47 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.57
+ $X2=1.63 $Y2=1.735
r48 5 7 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.63 $Y=1.57 $X2=1.63
+ $Y2=0.45
r49 1 12 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.9 $X2=1.22
+ $Y2=1.735
r50 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.22 $Y=1.9 $X2=1.22
+ $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_LP%A2 1 3 7 11 12 13 17
c43 17 0 1.3464e-19 $X=2.11 $Y=1.165
c44 1 0 1.52907e-19 $X=2.04 $Y=1.695
r45 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.165
+ $X2=2.11 $Y2=1.33
r46 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.165
+ $X2=2.11 $Y2=1
r47 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.165 $X2=2.11 $Y2=1.165
r48 12 13 14.1839 $w=3.88e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.195
+ $X2=2.64 $Y2=1.195
r49 12 18 1.47749 $w=3.88e-07 $l=5e-08 $layer=LI1_cond $X=2.16 $Y=1.195 $X2=2.11
+ $Y2=1.195
r50 11 20 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.09 $Y=1.57
+ $X2=2.09 $Y2=1.33
r51 7 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.02 $Y=0.45 $X2=2.02
+ $Y2=1
r52 1 11 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.04 $Y=1.695
+ $X2=2.04 $Y2=1.57
r53 1 3 214.912 $w=2.5e-07 $l=8.65e-07 $layer=POLY_cond $X=2.04 $Y=1.695
+ $X2=2.04 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_LP%C1 3 7 11 17 20 21 22 26
c44 21 0 1.3464e-19 $X=3.12 $Y=1.295
c45 7 0 2.54677e-19 $X=3.1 $Y=2.56
r46 21 22 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.11 $Y=1.275
+ $X2=3.11 $Y2=1.665
r47 21 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.11
+ $Y=1.275 $X2=3.11 $Y2=1.275
r48 19 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.11 $Y=1.615
+ $X2=3.11 $Y2=1.275
r49 19 20 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.615
+ $X2=3.11 $Y2=1.78
r50 16 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.11 $Y=1.26
+ $X2=3.11 $Y2=1.275
r51 16 17 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.11 $Y=1.185
+ $X2=3.23 $Y2=1.185
r52 13 16 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.87 $Y=1.185
+ $X2=3.11 $Y2=1.185
r53 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.23 $Y=1.11 $X2=3.23
+ $Y2=1.185
r54 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.23 $Y=1.11 $X2=3.23
+ $Y2=0.45
r55 7 20 193.794 $w=2.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.1 $Y=2.56 $X2=3.1
+ $Y2=1.78
r56 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.87 $Y=1.11 $X2=2.87
+ $Y2=1.185
r57 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.87 $Y=1.11 $X2=2.87
+ $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_LP%A_56_412# 1 2 7 9 11 18
c37 7 0 1.7238e-19 $X=0.425 $Y=2.25
r38 12 16 4.95428 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=0.59 $Y=2.165
+ $X2=0.425 $Y2=2.145
r39 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=2.165
+ $X2=2.835 $Y2=2.165
r40 11 12 135.701 $w=1.68e-07 $l=2.08e-06 $layer=LI1_cond $X=2.67 $Y=2.165
+ $X2=0.59 $Y2=2.165
r41 7 16 2.81189 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=0.425 $Y=2.25
+ $X2=0.425 $Y2=2.145
r42 7 9 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=0.425 $Y=2.25
+ $X2=0.425 $Y2=2.9
r43 2 18 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=2.695
+ $Y=2.06 $X2=2.835 $Y2=2.245
r44 1 16 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.28
+ $Y=2.06 $X2=0.425 $Y2=2.205
r45 1 9 400 $w=1.7e-07 $l=9.09615e-07 $layer=licon1_PDIFF $count=1 $X=0.28
+ $Y=2.06 $X2=0.425 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_LP%A_163_412# 1 2 7 10 11 12
c30 12 0 1.56513e-19 $X=2.305 $Y=2.6
c31 10 0 9.81645e-20 $X=2.14 $Y=2.515
r32 12 14 5.36061 $w=3.3e-07 $l=1.45e-07 $layer=LI1_cond $X=2.305 $Y=2.6
+ $X2=2.305 $Y2=2.745
r33 10 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.14 $Y=2.515
+ $X2=2.305 $Y2=2.6
r34 10 11 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=2.14 $Y=2.515
+ $X2=1.12 $Y2=2.515
r35 7 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.955 $Y=2.6
+ $X2=1.12 $Y2=2.515
r36 7 9 5.36061 $w=3.3e-07 $l=1.45e-07 $layer=LI1_cond $X=0.955 $Y=2.6 $X2=0.955
+ $Y2=2.745
r37 2 14 600 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_PDIFF $count=1 $X=2.165
+ $Y=2.06 $X2=2.305 $Y2=2.745
r38 1 9 600 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_PDIFF $count=1 $X=0.815
+ $Y=2.06 $X2=0.955 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_LP%VPWR 1 6 9 10 11 24 25
r37 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r38 21 24 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r39 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r40 19 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 18 19 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 15 19 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r43 14 18 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 11 25 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.6 $Y2=3.33
r46 11 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 9 18 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.32 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.485 $Y2=3.33
r49 8 21 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.65 $Y=3.33 $X2=1.68
+ $Y2=3.33
r50 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=1.485 $Y2=3.33
r51 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=3.245
+ $X2=1.485 $Y2=3.33
r52 4 6 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.485 $Y=3.245
+ $X2=1.485 $Y2=2.89
r53 1 6 600 $w=1.7e-07 $l=8.97274e-07 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=2.06 $X2=1.485 $Y2=2.89
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_LP%Y 1 2 3 12 15 18 23 24 25 26 30 36
r53 26 36 0.646529 $w=5.53e-07 $l=3e-08 $layer=LI1_cond $X=3.6 $Y=0.542 $X2=3.63
+ $Y2=0.542
r54 26 33 3.3404 $w=5.53e-07 $l=1.55e-07 $layer=LI1_cond $X=3.6 $Y=0.542
+ $X2=3.445 $Y2=0.542
r55 25 33 7.00406 $w=5.53e-07 $l=3.25e-07 $layer=LI1_cond $X=3.12 $Y=0.542
+ $X2=3.445 $Y2=0.542
r56 25 30 8.78658 $w=5.53e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=0.542
+ $X2=3.005 $Y2=0.542
r57 23 24 9.60999 $w=5.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.457 $Y=2.205
+ $X2=3.457 $Y2=2.04
r58 20 36 7.81693 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=3.63 $Y=0.82
+ $X2=3.63 $Y2=0.542
r59 20 24 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=3.63 $Y=0.82
+ $X2=3.63 $Y2=2.04
r60 16 23 2.13668 $w=5.13e-07 $l=9.2e-08 $layer=LI1_cond $X=3.457 $Y=2.297
+ $X2=3.457 $Y2=2.205
r61 16 18 14.0046 $w=5.13e-07 $l=6.03e-07 $layer=LI1_cond $X=3.457 $Y=2.297
+ $X2=3.457 $Y2=2.9
r62 15 30 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=1.58 $Y=0.735
+ $X2=3.005 $Y2=0.735
r63 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.415 $Y=0.65
+ $X2=1.58 $Y2=0.735
r64 10 12 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.415 $Y=0.65
+ $X2=1.415 $Y2=0.47
r65 3 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=2.06 $X2=3.365 $Y2=2.205
r66 3 18 400 $w=1.7e-07 $l=9.07304e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=2.06 $X2=3.365 $Y2=2.9
r67 2 33 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=3.305
+ $Y=0.24 $X2=3.445 $Y2=0.47
r68 1 12 182 $w=1.7e-07 $l=3.4641e-07 $layer=licon1_NDIFF $count=1 $X=1.165
+ $Y=0.24 $X2=1.415 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_LP%VGND 1 2 9 13 16 17 18 24 36 37 40
r45 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r46 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r47 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r48 34 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r49 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r50 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r51 31 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.235
+ $Y2=0
r52 31 33 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r53 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r54 27 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r55 26 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r56 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 24 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.235
+ $Y2=0
r58 24 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.68
+ $Y2=0
r59 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r60 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r61 18 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r62 18 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r63 16 21 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.24
+ $Y2=0
r64 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.485
+ $Y2=0
r65 15 26 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.65 $Y=0 $X2=0.72
+ $Y2=0
r66 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.65 $Y=0 $X2=0.485
+ $Y2=0
r67 11 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0
r68 11 13 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0.385
r69 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.485 $Y=0.085
+ $X2=0.485 $Y2=0
r70 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.485 $Y=0.085
+ $X2=0.485 $Y2=0.45
r71 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.095
+ $Y=0.24 $X2=2.235 $Y2=0.385
r72 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.34
+ $Y=0.24 $X2=0.485 $Y2=0.45
.ends

