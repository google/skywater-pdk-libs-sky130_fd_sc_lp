* File: sky130_fd_sc_lp__mux2i_1.pxi.spice
* Created: Fri Aug 28 10:44:59 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2I_1%A0 N_A0_M1005_g N_A0_M1002_g A0 N_A0_c_66_n
+ N_A0_c_67_n PM_SKY130_FD_SC_LP__MUX2I_1%A0
x_PM_SKY130_FD_SC_LP__MUX2I_1%A1 N_A1_M1000_g N_A1_M1007_g A1 N_A1_c_96_n
+ N_A1_c_99_n PM_SKY130_FD_SC_LP__MUX2I_1%A1
x_PM_SKY130_FD_SC_LP__MUX2I_1%A_304_237# N_A_304_237#_M1003_s
+ N_A_304_237#_M1001_s N_A_304_237#_M1004_g N_A_304_237#_c_131_n
+ N_A_304_237#_M1006_g N_A_304_237#_c_132_n N_A_304_237#_c_133_n
+ N_A_304_237#_c_140_n N_A_304_237#_c_134_n N_A_304_237#_c_135_n
+ N_A_304_237#_c_136_n N_A_304_237#_c_137_n
+ PM_SKY130_FD_SC_LP__MUX2I_1%A_304_237#
x_PM_SKY130_FD_SC_LP__MUX2I_1%S N_S_c_204_n N_S_M1009_g N_S_M1008_g N_S_c_199_n
+ N_S_c_200_n N_S_M1001_g N_S_M1003_g S S N_S_c_202_n N_S_c_203_n N_S_c_209_n
+ PM_SKY130_FD_SC_LP__MUX2I_1%S
x_PM_SKY130_FD_SC_LP__MUX2I_1%A_52_367# N_A_52_367#_M1002_s N_A_52_367#_M1009_d
+ N_A_52_367#_c_253_n N_A_52_367#_c_262_n N_A_52_367#_c_266_n
+ N_A_52_367#_c_254_n N_A_52_367#_c_255_n N_A_52_367#_c_256_n
+ N_A_52_367#_c_257_n N_A_52_367#_c_258_n PM_SKY130_FD_SC_LP__MUX2I_1%A_52_367#
x_PM_SKY130_FD_SC_LP__MUX2I_1%Y N_Y_M1005_d N_Y_M1002_d N_Y_c_305_n N_Y_c_307_n
+ N_Y_c_303_n N_Y_c_312_n Y PM_SKY130_FD_SC_LP__MUX2I_1%Y
x_PM_SKY130_FD_SC_LP__MUX2I_1%VPWR N_VPWR_M1004_d N_VPWR_M1001_d N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n VPWR
+ N_VPWR_c_344_n N_VPWR_c_338_n PM_SKY130_FD_SC_LP__MUX2I_1%VPWR
x_PM_SKY130_FD_SC_LP__MUX2I_1%A_29_73# N_A_29_73#_M1005_s N_A_29_73#_M1006_s
+ N_A_29_73#_c_377_n N_A_29_73#_c_378_n N_A_29_73#_c_379_n N_A_29_73#_c_380_n
+ PM_SKY130_FD_SC_LP__MUX2I_1%A_29_73#
x_PM_SKY130_FD_SC_LP__MUX2I_1%A_212_73# N_A_212_73#_M1000_d N_A_212_73#_M1008_d
+ N_A_212_73#_c_402_n N_A_212_73#_c_403_n N_A_212_73#_c_404_n
+ N_A_212_73#_c_405_n PM_SKY130_FD_SC_LP__MUX2I_1%A_212_73#
x_PM_SKY130_FD_SC_LP__MUX2I_1%VGND N_VGND_M1006_d N_VGND_M1003_d N_VGND_c_433_n
+ N_VGND_c_434_n N_VGND_c_435_n VGND N_VGND_c_436_n N_VGND_c_437_n
+ N_VGND_c_438_n N_VGND_c_439_n PM_SKY130_FD_SC_LP__MUX2I_1%VGND
cc_1 VNB N_A0_M1005_g 0.0247584f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.785
cc_2 VNB N_A0_c_66_n 0.016888f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_3 VNB N_A0_c_67_n 0.0369392f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.51
cc_4 VNB N_A1_M1000_g 0.0214731f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.785
cc_5 VNB N_A1_c_96_n 0.0303988f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_6 VNB N_A_304_237#_c_131_n 0.0196339f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_7 VNB N_A_304_237#_c_132_n 0.0156165f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.51
cc_8 VNB N_A_304_237#_c_133_n 0.0520039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_304_237#_c_134_n 0.00591273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_304_237#_c_135_n 0.0065993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_304_237#_c_136_n 0.00257434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_304_237#_c_137_n 0.00119135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_S_M1008_g 0.0443315f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.465
cc_14 VNB N_S_c_199_n 0.0237604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_S_c_200_n 0.00934934f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB S 0.0201073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_S_c_202_n 0.040007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_S_c_203_n 0.0224069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_303_n 0.00581426f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_20 VNB N_VPWR_c_338_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_29_73#_c_377_n 0.0287893f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_29_73#_c_378_n 0.0118375f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_23 VNB N_A_29_73#_c_379_n 0.00964068f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_24 VNB N_A_29_73#_c_380_n 0.00627997f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.51
cc_25 VNB N_A_212_73#_c_402_n 0.00541478f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_A_212_73#_c_403_n 0.020734f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_27 VNB N_A_212_73#_c_404_n 0.00465651f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_28 VNB N_A_212_73#_c_405_n 0.00830279f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.675
cc_29 VNB N_VGND_c_433_n 0.00494808f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_30 VNB N_VGND_c_434_n 0.0111997f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_31 VNB N_VGND_c_435_n 0.0358916f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_32 VNB N_VGND_c_436_n 0.0510556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_437_n 0.0302975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_438_n 0.00422795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_439_n 0.230443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_A0_M1002_g 0.0238802f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.465
cc_37 VPB N_A0_c_66_n 0.0113903f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_38 VPB N_A0_c_67_n 0.0118054f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.51
cc_39 VPB N_A1_M1007_g 0.0197017f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.465
cc_40 VPB N_A1_c_96_n 0.00856789f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_41 VPB N_A1_c_99_n 0.00311548f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_42 VPB N_A_304_237#_M1004_g 0.0221626f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_43 VPB N_A_304_237#_c_133_n 0.00647369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_304_237#_c_140_n 0.0169342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_S_c_204_n 0.0218864f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.345
cc_46 VPB N_S_c_199_n 0.0314314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_S_c_200_n 0.00651558f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_48 VPB S 0.00842008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_S_c_202_n 0.011931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_S_c_209_n 0.0238302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_52_367#_c_253_n 0.0150427f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_52 VPB N_A_52_367#_c_254_n 0.00370537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_52_367#_c_255_n 0.00100448f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.665
cc_54 VPB N_A_52_367#_c_256_n 0.00435424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_52_367#_c_257_n 0.0128177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_52_367#_c_258_n 0.0314089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_303_n 0.00142808f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_58 VPB N_VPWR_c_339_n 0.00562917f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_59 VPB N_VPWR_c_340_n 0.0116157f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_60 VPB N_VPWR_c_341_n 0.0484529f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.675
cc_61 VPB N_VPWR_c_342_n 0.0561781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_343_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_344_n 0.0334364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_338_n 0.0659178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 N_A0_M1005_g N_A1_M1000_g 0.00948562f $X=0.505 $Y=0.785 $X2=0 $Y2=0
cc_66 N_A0_M1002_g N_A1_M1007_g 0.0442777f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_67 N_A0_c_67_n N_A1_c_96_n 0.0189289f $X=0.505 $Y=1.51 $X2=0 $Y2=0
cc_68 N_A0_M1002_g N_A1_c_99_n 2.10941e-19 $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_69 N_A0_M1002_g N_A_52_367#_c_253_n 0.00430102f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A0_c_66_n N_A_52_367#_c_253_n 0.0238424f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_71 N_A0_c_67_n N_A_52_367#_c_253_n 0.00158197f $X=0.505 $Y=1.51 $X2=0 $Y2=0
cc_72 N_A0_M1002_g N_A_52_367#_c_262_n 0.0148524f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A0_c_67_n N_A_52_367#_c_258_n 0.00124124f $X=0.505 $Y=1.51 $X2=0 $Y2=0
cc_74 N_A0_M1005_g N_Y_c_305_n 0.00304419f $X=0.505 $Y=0.785 $X2=0 $Y2=0
cc_75 N_A0_c_67_n N_Y_c_305_n 0.00125565f $X=0.505 $Y=1.51 $X2=0 $Y2=0
cc_76 N_A0_M1005_g N_Y_c_307_n 0.00462974f $X=0.505 $Y=0.785 $X2=0 $Y2=0
cc_77 N_A0_M1005_g N_Y_c_303_n 0.00552331f $X=0.505 $Y=0.785 $X2=0 $Y2=0
cc_78 N_A0_M1002_g N_Y_c_303_n 0.00962004f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A0_c_66_n N_Y_c_303_n 0.0310007f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_80 N_A0_c_67_n N_Y_c_303_n 0.0050591f $X=0.505 $Y=1.51 $X2=0 $Y2=0
cc_81 N_A0_M1002_g N_Y_c_312_n 0.00356755f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A0_M1002_g N_VPWR_c_342_n 0.00585385f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A0_M1002_g N_VPWR_c_338_n 0.00750563f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_84 N_A0_c_66_n N_A_29_73#_c_377_n 0.0235027f $X=0.385 $Y=1.51 $X2=0 $Y2=0
cc_85 N_A0_c_67_n N_A_29_73#_c_377_n 0.00126468f $X=0.505 $Y=1.51 $X2=0 $Y2=0
cc_86 N_A0_M1005_g N_A_29_73#_c_378_n 0.0134471f $X=0.505 $Y=0.785 $X2=0 $Y2=0
cc_87 N_A0_M1005_g N_VGND_c_436_n 0.0028086f $X=0.505 $Y=0.785 $X2=0 $Y2=0
cc_88 N_A0_M1005_g N_VGND_c_439_n 0.00370953f $X=0.505 $Y=0.785 $X2=0 $Y2=0
cc_89 N_A1_M1007_g N_A_304_237#_M1004_g 0.05621f $X=1.105 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A1_c_99_n N_A_304_237#_M1004_g 0.00172645f $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_91 N_A1_c_96_n N_A_304_237#_c_132_n 6.37767e-19 $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_92 N_A1_c_99_n N_A_304_237#_c_132_n 0.0107083f $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_93 N_A1_M1000_g N_A_304_237#_c_133_n 0.00467083f $X=0.985 $Y=0.785 $X2=0
+ $Y2=0
cc_94 N_A1_c_96_n N_A_304_237#_c_133_n 0.0223826f $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_95 N_A1_c_99_n N_A_304_237#_c_133_n 8.50287e-19 $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_96 N_A1_M1007_g N_A_52_367#_c_262_n 0.015311f $X=1.105 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A1_c_99_n N_A_52_367#_c_262_n 8.15308e-19 $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_98 N_A1_M1007_g N_A_52_367#_c_266_n 0.0035844f $X=1.105 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A1_M1007_g N_A_52_367#_c_255_n 0.00144302f $X=1.105 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A1_M1000_g N_Y_c_303_n 0.00641219f $X=0.985 $Y=0.785 $X2=0 $Y2=0
cc_101 N_A1_M1007_g N_Y_c_303_n 0.00232397f $X=1.105 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A1_c_99_n N_Y_c_303_n 0.0247324f $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_103 N_A1_M1007_g Y 0.0086629f $X=1.105 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A1_c_96_n Y 0.00310929f $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_105 N_A1_c_99_n Y 0.0183035f $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_106 N_A1_M1007_g N_VPWR_c_342_n 0.00585385f $X=1.105 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A1_M1007_g N_VPWR_c_338_n 0.00671188f $X=1.105 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A1_M1000_g N_A_29_73#_c_378_n 0.0158868f $X=0.985 $Y=0.785 $X2=0 $Y2=0
cc_109 N_A1_M1000_g N_A_29_73#_c_380_n 0.00305414f $X=0.985 $Y=0.785 $X2=0 $Y2=0
cc_110 N_A1_M1000_g N_A_212_73#_c_402_n 0.00421736f $X=0.985 $Y=0.785 $X2=0
+ $Y2=0
cc_111 N_A1_M1000_g N_A_212_73#_c_404_n 0.0022996f $X=0.985 $Y=0.785 $X2=0 $Y2=0
cc_112 N_A1_c_96_n N_A_212_73#_c_404_n 0.00689467f $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_113 N_A1_c_99_n N_A_212_73#_c_404_n 0.0204895f $X=1.145 $Y=1.51 $X2=0 $Y2=0
cc_114 N_A1_M1000_g N_VGND_c_436_n 0.0028086f $X=0.985 $Y=0.785 $X2=0 $Y2=0
cc_115 N_A1_M1000_g N_VGND_c_439_n 0.00369932f $X=0.985 $Y=0.785 $X2=0 $Y2=0
cc_116 N_A_304_237#_c_140_n N_S_c_204_n 0.00233396f $X=3.11 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_304_237#_c_131_n N_S_M1008_g 0.0256967f $X=1.965 $Y=1.185 $X2=0 $Y2=0
cc_118 N_A_304_237#_c_132_n N_S_M1008_g 0.0105881f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_119 N_A_304_237#_c_133_n N_S_M1008_g 0.00715251f $X=1.685 $Y=1.5 $X2=0 $Y2=0
cc_120 N_A_304_237#_c_134_n N_S_M1008_g 0.00112869f $X=3.15 $Y=0.525 $X2=0 $Y2=0
cc_121 N_A_304_237#_c_135_n N_S_M1008_g 0.00418195f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_122 N_A_304_237#_c_137_n N_S_M1008_g 6.31488e-19 $X=3.115 $Y=1.095 $X2=0
+ $Y2=0
cc_123 N_A_304_237#_c_132_n N_S_c_199_n 0.0217933f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_124 N_A_304_237#_c_140_n N_S_c_199_n 0.0169281f $X=3.11 $Y=2.045 $X2=0 $Y2=0
cc_125 N_A_304_237#_c_136_n N_S_c_199_n 0.00530855f $X=3.075 $Y=1.5 $X2=0 $Y2=0
cc_126 N_A_304_237#_M1004_g N_S_c_200_n 0.0223989f $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_304_237#_c_132_n N_S_c_200_n 0.00832163f $X=2.945 $Y=1.5 $X2=0 $Y2=0
cc_128 N_A_304_237#_c_133_n N_S_c_200_n 0.00621888f $X=1.685 $Y=1.5 $X2=0 $Y2=0
cc_129 N_A_304_237#_c_140_n S 0.0123198f $X=3.11 $Y=2.045 $X2=0 $Y2=0
cc_130 N_A_304_237#_c_135_n S 0.0158037f $X=3.095 $Y=1.415 $X2=0 $Y2=0
cc_131 N_A_304_237#_c_136_n S 0.0144294f $X=3.075 $Y=1.5 $X2=0 $Y2=0
cc_132 N_A_304_237#_c_135_n N_S_c_202_n 0.00325694f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_133 N_A_304_237#_c_136_n N_S_c_202_n 0.00449979f $X=3.075 $Y=1.5 $X2=0 $Y2=0
cc_134 N_A_304_237#_c_135_n N_S_c_203_n 0.00566865f $X=3.095 $Y=1.415 $X2=0
+ $Y2=0
cc_135 N_A_304_237#_c_140_n N_S_c_209_n 0.00596708f $X=3.11 $Y=2.045 $X2=0 $Y2=0
cc_136 N_A_304_237#_M1004_g N_A_52_367#_c_262_n 0.00976877f $X=1.595 $Y=2.465
+ $X2=0 $Y2=0
cc_137 N_A_304_237#_M1004_g N_A_52_367#_c_266_n 0.00886513f $X=1.595 $Y=2.465
+ $X2=0 $Y2=0
cc_138 N_A_304_237#_M1004_g N_A_52_367#_c_254_n 0.00619663f $X=1.595 $Y=2.465
+ $X2=0 $Y2=0
cc_139 N_A_304_237#_c_132_n N_A_52_367#_c_254_n 0.0383672f $X=2.945 $Y=1.5 $X2=0
+ $Y2=0
cc_140 N_A_304_237#_c_133_n N_A_52_367#_c_254_n 0.005892f $X=1.685 $Y=1.5 $X2=0
+ $Y2=0
cc_141 N_A_304_237#_M1004_g N_A_52_367#_c_255_n 0.00454058f $X=1.595 $Y=2.465
+ $X2=0 $Y2=0
cc_142 N_A_304_237#_c_132_n N_A_52_367#_c_255_n 0.00627388f $X=2.945 $Y=1.5
+ $X2=0 $Y2=0
cc_143 N_A_304_237#_c_132_n N_A_52_367#_c_256_n 0.0192945f $X=2.945 $Y=1.5 $X2=0
+ $Y2=0
cc_144 N_A_304_237#_c_140_n N_A_52_367#_c_256_n 0.00895415f $X=3.11 $Y=2.045
+ $X2=0 $Y2=0
cc_145 N_A_304_237#_c_140_n N_A_52_367#_c_257_n 0.0536892f $X=3.11 $Y=2.045
+ $X2=0 $Y2=0
cc_146 N_A_304_237#_M1004_g Y 7.34957e-19 $X=1.595 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_304_237#_M1004_g N_VPWR_c_339_n 0.0206386f $X=1.595 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_304_237#_M1004_g N_VPWR_c_342_n 0.00585385f $X=1.595 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_304_237#_c_140_n N_VPWR_c_344_n 0.0178111f $X=3.11 $Y=2.045 $X2=0
+ $Y2=0
cc_150 N_A_304_237#_M1001_s N_VPWR_c_338_n 0.00371702f $X=2.985 $Y=1.835 $X2=0
+ $Y2=0
cc_151 N_A_304_237#_M1004_g N_VPWR_c_338_n 0.00838452f $X=1.595 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_304_237#_c_140_n N_VPWR_c_338_n 0.0100304f $X=3.11 $Y=2.045 $X2=0
+ $Y2=0
cc_153 N_A_304_237#_c_131_n N_A_29_73#_c_380_n 0.00810964f $X=1.965 $Y=1.185
+ $X2=0 $Y2=0
cc_154 N_A_304_237#_c_133_n N_A_29_73#_c_380_n 0.00166511f $X=1.685 $Y=1.5 $X2=0
+ $Y2=0
cc_155 N_A_304_237#_c_131_n N_A_212_73#_c_402_n 0.00368285f $X=1.965 $Y=1.185
+ $X2=0 $Y2=0
cc_156 N_A_304_237#_c_131_n N_A_212_73#_c_403_n 0.0112877f $X=1.965 $Y=1.185
+ $X2=0 $Y2=0
cc_157 N_A_304_237#_c_132_n N_A_212_73#_c_403_n 0.0925578f $X=2.945 $Y=1.5 $X2=0
+ $Y2=0
cc_158 N_A_304_237#_c_133_n N_A_212_73#_c_403_n 0.0169444f $X=1.685 $Y=1.5 $X2=0
+ $Y2=0
cc_159 N_A_304_237#_c_137_n N_A_212_73#_c_403_n 0.0125761f $X=3.115 $Y=1.095
+ $X2=0 $Y2=0
cc_160 N_A_304_237#_c_134_n N_A_212_73#_c_405_n 0.0497997f $X=3.15 $Y=0.525
+ $X2=0 $Y2=0
cc_161 N_A_304_237#_c_131_n N_VGND_c_433_n 0.00284552f $X=1.965 $Y=1.185 $X2=0
+ $Y2=0
cc_162 N_A_304_237#_c_131_n N_VGND_c_436_n 0.00547432f $X=1.965 $Y=1.185 $X2=0
+ $Y2=0
cc_163 N_A_304_237#_c_134_n N_VGND_c_437_n 0.0105928f $X=3.15 $Y=0.525 $X2=0
+ $Y2=0
cc_164 N_A_304_237#_c_131_n N_VGND_c_439_n 0.0110536f $X=1.965 $Y=1.185 $X2=0
+ $Y2=0
cc_165 N_A_304_237#_c_134_n N_VGND_c_439_n 0.00947127f $X=3.15 $Y=0.525 $X2=0
+ $Y2=0
cc_166 N_S_c_204_n N_A_52_367#_c_266_n 3.28686e-19 $X=2.215 $Y=1.725 $X2=0 $Y2=0
cc_167 N_S_c_204_n N_A_52_367#_c_254_n 0.0145701f $X=2.215 $Y=1.725 $X2=0 $Y2=0
cc_168 N_S_c_200_n N_A_52_367#_c_256_n 0.0063861f $X=2.47 $Y=1.65 $X2=0 $Y2=0
cc_169 N_S_c_204_n N_VPWR_c_339_n 0.00342995f $X=2.215 $Y=1.725 $X2=0 $Y2=0
cc_170 S N_VPWR_c_341_n 0.0269148f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_171 N_S_c_202_n N_VPWR_c_341_n 0.00163524f $X=3.48 $Y=1.46 $X2=0 $Y2=0
cc_172 N_S_c_209_n N_VPWR_c_341_n 0.0224724f $X=3.447 $Y=1.725 $X2=0 $Y2=0
cc_173 N_S_c_204_n N_VPWR_c_344_n 0.00585385f $X=2.215 $Y=1.725 $X2=0 $Y2=0
cc_174 N_S_c_209_n N_VPWR_c_344_n 0.00486043f $X=3.447 $Y=1.725 $X2=0 $Y2=0
cc_175 N_S_c_204_n N_VPWR_c_338_n 0.0122513f $X=2.215 $Y=1.725 $X2=0 $Y2=0
cc_176 N_S_c_209_n N_VPWR_c_338_n 0.00954696f $X=3.447 $Y=1.725 $X2=0 $Y2=0
cc_177 N_S_M1008_g N_A_212_73#_c_403_n 0.0164148f $X=2.395 $Y=0.655 $X2=0 $Y2=0
cc_178 N_S_c_199_n N_A_212_73#_c_403_n 0.00117872f $X=3.25 $Y=1.65 $X2=0 $Y2=0
cc_179 N_S_c_200_n N_A_212_73#_c_403_n 8.50214e-19 $X=2.47 $Y=1.65 $X2=0 $Y2=0
cc_180 N_S_c_203_n N_A_212_73#_c_405_n 0.00264824f $X=3.447 $Y=1.295 $X2=0 $Y2=0
cc_181 N_S_M1008_g N_VGND_c_433_n 0.00301542f $X=2.395 $Y=0.655 $X2=0 $Y2=0
cc_182 S N_VGND_c_435_n 0.0269149f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_183 N_S_c_202_n N_VGND_c_435_n 0.00115333f $X=3.48 $Y=1.46 $X2=0 $Y2=0
cc_184 N_S_c_203_n N_VGND_c_435_n 0.0155587f $X=3.447 $Y=1.295 $X2=0 $Y2=0
cc_185 N_S_M1008_g N_VGND_c_437_n 0.00585385f $X=2.395 $Y=0.655 $X2=0 $Y2=0
cc_186 N_S_c_203_n N_VGND_c_437_n 0.00400407f $X=3.447 $Y=1.295 $X2=0 $Y2=0
cc_187 N_S_M1008_g N_VGND_c_439_n 0.0118611f $X=2.395 $Y=0.655 $X2=0 $Y2=0
cc_188 N_S_c_203_n N_VGND_c_439_n 0.00804497f $X=3.447 $Y=1.295 $X2=0 $Y2=0
cc_189 N_A_52_367#_c_262_n N_Y_M1002_d 0.0065545f $X=1.455 $Y=2.43 $X2=0 $Y2=0
cc_190 N_A_52_367#_c_255_n N_Y_c_303_n 0.00334559f $X=1.625 $Y=1.9 $X2=0 $Y2=0
cc_191 N_A_52_367#_c_253_n N_Y_c_312_n 0.0169848f $X=0.385 $Y=2.095 $X2=0 $Y2=0
cc_192 N_A_52_367#_c_262_n N_Y_c_312_n 0.00896709f $X=1.455 $Y=2.43 $X2=0 $Y2=0
cc_193 N_A_52_367#_c_262_n Y 0.0265177f $X=1.455 $Y=2.43 $X2=0 $Y2=0
cc_194 N_A_52_367#_c_266_n Y 0.0124385f $X=1.54 $Y=2.31 $X2=0 $Y2=0
cc_195 N_A_52_367#_c_255_n Y 0.00484964f $X=1.625 $Y=1.9 $X2=0 $Y2=0
cc_196 N_A_52_367#_c_262_n A_236_367# 0.0111476f $X=1.455 $Y=2.43 $X2=-0.19
+ $Y2=1.655
cc_197 N_A_52_367#_c_266_n A_236_367# 0.00346838f $X=1.54 $Y=2.31 $X2=-0.19
+ $Y2=1.655
cc_198 N_A_52_367#_c_255_n A_236_367# 0.00209931f $X=1.625 $Y=1.9 $X2=-0.19
+ $Y2=1.655
cc_199 N_A_52_367#_c_254_n N_VPWR_M1004_d 0.00659079f $X=2.295 $Y=1.9 $X2=-0.19
+ $Y2=1.655
cc_200 N_A_52_367#_c_262_n N_VPWR_c_339_n 0.0197769f $X=1.455 $Y=2.43 $X2=0
+ $Y2=0
cc_201 N_A_52_367#_c_266_n N_VPWR_c_339_n 0.011435f $X=1.54 $Y=2.31 $X2=0 $Y2=0
cc_202 N_A_52_367#_c_254_n N_VPWR_c_339_n 0.0233499f $X=2.295 $Y=1.9 $X2=0 $Y2=0
cc_203 N_A_52_367#_c_258_n N_VPWR_c_342_n 0.0218897f $X=0.41 $Y=2.49 $X2=0 $Y2=0
cc_204 N_A_52_367#_c_257_n N_VPWR_c_344_n 0.0192303f $X=2.43 $Y=2.91 $X2=0 $Y2=0
cc_205 N_A_52_367#_M1002_s N_VPWR_c_338_n 0.00246193f $X=0.26 $Y=1.835 $X2=0
+ $Y2=0
cc_206 N_A_52_367#_M1009_d N_VPWR_c_338_n 0.00232552f $X=2.29 $Y=1.835 $X2=0
+ $Y2=0
cc_207 N_A_52_367#_c_262_n N_VPWR_c_338_n 0.0386732f $X=1.455 $Y=2.43 $X2=0
+ $Y2=0
cc_208 N_A_52_367#_c_257_n N_VPWR_c_338_n 0.0115856f $X=2.43 $Y=2.91 $X2=0 $Y2=0
cc_209 N_A_52_367#_c_258_n N_VPWR_c_338_n 0.0127519f $X=0.41 $Y=2.49 $X2=0 $Y2=0
cc_210 N_A_52_367#_c_255_n N_A_212_73#_c_403_n 0.0021965f $X=1.625 $Y=1.9 $X2=0
+ $Y2=0
cc_211 Y A_236_367# 0.002792f $X=1.115 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_212 N_Y_M1002_d N_VPWR_c_338_n 0.0045459f $X=0.7 $Y=1.835 $X2=0 $Y2=0
cc_213 N_Y_M1005_d N_A_29_73#_c_378_n 0.00229612f $X=0.58 $Y=0.365 $X2=0 $Y2=0
cc_214 N_Y_c_307_n N_A_29_73#_c_378_n 0.018046f $X=0.72 $Y=0.68 $X2=0 $Y2=0
cc_215 N_Y_c_305_n N_A_212_73#_c_404_n 6.11933e-19 $X=0.72 $Y=1 $X2=0 $Y2=0
cc_216 N_Y_c_303_n N_A_212_73#_c_404_n 0.00417432f $X=0.725 $Y=1.93 $X2=0 $Y2=0
cc_217 A_236_367# N_VPWR_c_338_n 0.00468268f $X=1.18 $Y=1.835 $X2=0 $Y2=0
cc_218 N_A_29_73#_c_378_n N_A_212_73#_M1000_d 0.00290554f $X=1.585 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_219 N_A_29_73#_c_378_n N_A_212_73#_c_402_n 0.0205822f $X=1.585 $Y=0.34 $X2=0
+ $Y2=0
cc_220 N_A_29_73#_c_380_n N_A_212_73#_c_402_n 0.0230301f $X=1.75 $Y=0.38 $X2=0
+ $Y2=0
cc_221 N_A_29_73#_c_378_n N_A_212_73#_c_403_n 0.00587992f $X=1.585 $Y=0.34 $X2=0
+ $Y2=0
cc_222 N_A_29_73#_c_380_n N_A_212_73#_c_403_n 0.0243529f $X=1.75 $Y=0.38 $X2=0
+ $Y2=0
cc_223 N_A_29_73#_c_378_n N_VGND_c_436_n 0.0763704f $X=1.585 $Y=0.34 $X2=0 $Y2=0
cc_224 N_A_29_73#_c_379_n N_VGND_c_436_n 0.0200723f $X=0.385 $Y=0.34 $X2=0 $Y2=0
cc_225 N_A_29_73#_c_380_n N_VGND_c_436_n 0.0211235f $X=1.75 $Y=0.38 $X2=0 $Y2=0
cc_226 N_A_29_73#_M1006_s N_VGND_c_439_n 0.00215158f $X=1.625 $Y=0.235 $X2=0
+ $Y2=0
cc_227 N_A_29_73#_c_378_n N_VGND_c_439_n 0.0437442f $X=1.585 $Y=0.34 $X2=0 $Y2=0
cc_228 N_A_29_73#_c_379_n N_VGND_c_439_n 0.0108858f $X=0.385 $Y=0.34 $X2=0 $Y2=0
cc_229 N_A_29_73#_c_380_n N_VGND_c_439_n 0.012627f $X=1.75 $Y=0.38 $X2=0 $Y2=0
cc_230 N_A_212_73#_c_403_n N_VGND_c_433_n 0.0156925f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A_212_73#_c_405_n N_VGND_c_435_n 0.00300084f $X=2.61 $Y=0.42 $X2=0
+ $Y2=0
cc_232 N_A_212_73#_c_405_n N_VGND_c_437_n 0.0186981f $X=2.61 $Y=0.42 $X2=0 $Y2=0
cc_233 N_A_212_73#_M1008_d N_VGND_c_439_n 0.00284733f $X=2.47 $Y=0.235 $X2=0
+ $Y2=0
cc_234 N_A_212_73#_c_405_n N_VGND_c_439_n 0.0110024f $X=2.61 $Y=0.42 $X2=0 $Y2=0
