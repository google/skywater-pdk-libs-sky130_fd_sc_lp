* File: sky130_fd_sc_lp__o221ai_lp.pex.spice
* Created: Wed Sep  2 10:19:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221AI_LP%C1 1 3 7 9
r35 9 12 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=1.215 $X2=0.71 $Y2=1.215
r36 5 12 42.9487 $w=5.39e-07 $l=2.52357e-07 $layer=POLY_cond $X=1.005 $Y=1.05
+ $X2=0.822 $Y2=1.215
r37 5 7 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.005 $Y=1.05
+ $X2=1.005 $Y2=0.485
r38 1 12 59.131 $w=5.39e-07 $l=5.76446e-07 $layer=POLY_cond $X=0.975 $Y=1.72
+ $X2=0.822 $Y2=1.215
r39 1 3 217.397 $w=2.5e-07 $l=8.75e-07 $layer=POLY_cond $X=0.975 $Y=1.72
+ $X2=0.975 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_LP%B1 3 6 9 11 12 13 17
r47 17 19 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.547 $Y=1.345
+ $X2=1.547 $Y2=1.18
r48 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.57
+ $Y=1.345 $X2=1.57 $Y2=1.345
r49 13 18 9.45594 $w=3.88e-07 $l=3.2e-07 $layer=LI1_cond $X=1.6 $Y=1.665 $X2=1.6
+ $Y2=1.345
r50 12 18 1.47749 $w=3.88e-07 $l=5e-08 $layer=LI1_cond $X=1.6 $Y=1.295 $X2=1.6
+ $Y2=1.345
r51 9 11 185.098 $w=2.5e-07 $l=7.45e-07 $layer=POLY_cond $X=1.61 $Y=2.595
+ $X2=1.61 $Y2=1.85
r52 6 11 33.9275 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=1.547 $Y=1.663
+ $X2=1.547 $Y2=1.85
r53 5 17 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=1.547 $Y=1.367
+ $X2=1.547 $Y2=1.345
r54 5 6 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=1.547 $Y=1.367
+ $X2=1.547 $Y2=1.663
r55 3 19 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.435 $Y=0.485
+ $X2=1.435 $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_LP%B2 3 7 11 14 15 20 21 25 26
c62 7 0 1.79821e-20 $X=3.58 $Y=0.485
r63 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.67
+ $Y=1.06 $X2=3.67 $Y2=1.06
r64 20 21 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.66 $Y=1.295
+ $X2=3.66 $Y2=1.665
r65 20 26 7.73783 $w=3.48e-07 $l=2.35e-07 $layer=LI1_cond $X=3.66 $Y=1.295
+ $X2=3.66 $Y2=1.06
r66 19 21 3.29269 $w=3.48e-07 $l=1e-07 $layer=LI1_cond $X=3.66 $Y=1.765 $X2=3.66
+ $Y2=1.665
r67 15 30 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.77
+ $X2=2.14 $Y2=1.935
r68 14 17 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.14 $Y=1.77 $X2=2.14
+ $Y2=1.85
r69 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.77 $X2=2.14 $Y2=1.77
r70 12 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=1.85
+ $X2=2.14 $Y2=1.85
r71 11 19 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=3.485 $Y=1.85
+ $X2=3.66 $Y2=1.765
r72 11 12 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=3.485 $Y=1.85
+ $X2=2.305 $Y2=1.85
r73 10 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=0.895
+ $X2=3.67 $Y2=1.06
r74 7 10 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.58 $Y=0.485
+ $X2=3.58 $Y2=0.895
r75 3 30 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.1 $Y=2.595 $X2=2.1
+ $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_LP%A2 3 4 5 8 10 13 14 16 17 18 22
c62 22 0 1.32013e-19 $X=2.185 $Y=1.2
c63 13 0 1.17138e-19 $X=2.11 $Y=0.79
r64 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.185
+ $Y=1.2 $X2=2.185 $Y2=1.2
r65 18 23 13.983 $w=3.73e-07 $l=4.55e-07 $layer=LI1_cond $X=2.64 $Y=1.222
+ $X2=2.185 $Y2=1.222
r66 17 23 0.768295 $w=3.73e-07 $l=2.5e-08 $layer=LI1_cond $X=2.16 $Y=1.222
+ $X2=2.185 $Y2=1.222
r67 15 22 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.185 $Y=1.215
+ $X2=2.185 $Y2=1.2
r68 14 22 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=2.185 $Y=0.94
+ $X2=2.185 $Y2=1.2
r69 13 14 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.11 $Y=0.79
+ $X2=2.11 $Y2=0.94
r70 8 16 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.67 $Y=1.95
+ $X2=2.67 $Y2=1.825
r71 8 10 160.253 $w=2.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.67 $Y=1.95
+ $X2=2.67 $Y2=2.595
r72 6 16 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.62 $Y=1.365
+ $X2=2.62 $Y2=1.825
r73 5 15 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.35 $Y=1.29
+ $X2=2.185 $Y2=1.215
r74 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.545 $Y=1.29
+ $X2=2.62 $Y2=1.365
r75 4 5 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.545 $Y=1.29
+ $X2=2.35 $Y2=1.29
r76 3 13 98.0067 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.945 $Y=0.485
+ $X2=1.945 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_LP%A1 3 5 9 13 14 15 16 19 20
c48 20 0 1.32013e-19 $X=3.1 $Y=1.08
r49 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.1 $Y=1.08
+ $X2=3.1 $Y2=1.08
r50 16 20 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.1 $Y=1.295
+ $X2=3.1 $Y2=1.08
r51 14 15 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.11 $Y=1.585
+ $X2=3.11 $Y2=1.805
r52 13 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.1 $Y=1.42 $X2=3.1
+ $Y2=1.08
r53 13 14 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.42 $X2=3.1
+ $Y2=1.585
r54 12 19 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=0.915
+ $X2=3.1 $Y2=1.08
r55 9 12 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.15 $Y=0.485
+ $X2=3.15 $Y2=0.915
r56 3 15 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=3.16 $Y=1.93
+ $X2=3.16 $Y2=1.805
r57 3 5 165.222 $w=2.5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.16 $Y=1.93 $X2=3.16
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_LP%Y 1 2 3 12 14 16 20 22 23 31
r44 23 39 2.31242 $w=7.48e-07 $l=1.45e-07 $layer=LI1_cond $X=0.5 $Y=2.405
+ $X2=0.5 $Y2=2.55
r45 23 35 2.63137 $w=7.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.5 $Y=2.405
+ $X2=0.5 $Y2=2.24
r46 22 35 3.26928 $w=7.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.5 $Y=2.035
+ $X2=0.5 $Y2=2.24
r47 22 31 10.3256 $w=7.48e-07 $l=1.15e-07 $layer=LI1_cond $X=0.5 $Y=2.035
+ $X2=0.5 $Y2=1.92
r48 18 20 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.365 $Y=2.635
+ $X2=2.365 $Y2=2.765
r49 17 39 9.77808 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=0.875 $Y=2.55
+ $X2=0.5 $Y2=2.55
r50 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.2 $Y=2.55
+ $X2=2.365 $Y2=2.635
r51 16 17 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=2.2 $Y=2.55
+ $X2=0.875 $Y2=2.55
r52 12 14 13.1569 $w=4.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.295 $Y=0.49
+ $X2=0.79 $Y2=0.49
r53 10 12 8.80477 $w=4.5e-07 $l=2.64102e-07 $layer=LI1_cond $X=0.21 $Y=0.715
+ $X2=0.295 $Y2=0.49
r54 10 31 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=0.21 $Y=0.715
+ $X2=0.21 $Y2=1.92
r55 3 20 600 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=2.095 $X2=2.365 $Y2=2.765
r56 2 35 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.565
+ $Y=2.095 $X2=0.71 $Y2=2.24
r57 1 14 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.645
+ $Y=0.275 $X2=0.79 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_LP%VPWR 1 2 9 13 16 17 18 20 33 34 37
r42 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r44 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=3.33
+ $X2=1.24 $Y2=3.33
r50 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.405 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=1.24 $Y2=3.33
r54 20 22 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.075 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 18 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 16 30 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.425 $Y2=3.33
r59 15 33 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.59 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=3.33
+ $X2=3.425 $Y2=3.33
r61 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.425 $Y2=3.33
r62 11 13 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.425 $Y2=2.79
r63 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=3.245 $X2=1.24
+ $Y2=3.33
r64 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.24 $Y=3.245 $X2=1.24
+ $Y2=2.925
r65 2 13 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=2.095 $X2=3.425 $Y2=2.79
r66 1 9 600 $w=1.7e-07 $l=8.97274e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=2.095 $X2=1.24 $Y2=2.925
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_LP%A_216_55# 1 2 9 12 13 14 16 17 21
c58 9 0 1.17138e-19 $X=1.22 $Y=0.49
r59 19 21 5.98039 $w=4.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.875 $Y=0.49
+ $X2=4.1 $Y2=0.49
r60 15 21 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=4.1 $Y=0.715 $X2=4.1
+ $Y2=0.49
r61 15 16 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=4.1 $Y=0.715 $X2=4.1
+ $Y2=2.115
r62 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=2.2
+ $X2=4.1 $Y2=2.115
r63 13 14 182.021 $w=1.68e-07 $l=2.79e-06 $layer=LI1_cond $X=4.015 $Y=2.2
+ $X2=1.225 $Y2=2.2
r64 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.14 $Y=2.115
+ $X2=1.225 $Y2=2.2
r65 12 17 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=1.14 $Y=2.115
+ $X2=1.14 $Y2=0.895
r66 7 17 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=0.73
+ $X2=1.22 $Y2=0.895
r67 7 9 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.22 $Y=0.73 $X2=1.22
+ $Y2=0.49
r68 2 19 182 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_NDIFF $count=1 $X=3.655
+ $Y=0.275 $X2=3.875 $Y2=0.49
r69 1 9 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.275 $X2=1.22 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_LP%A_302_55# 1 2 9 11 12 13 15 20
c49 13 0 1.79821e-20 $X=3.2 $Y=0.63
r50 20 22 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.365 $Y=0.49
+ $X2=3.365 $Y2=0.63
r51 15 17 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.67 $Y=0.63
+ $X2=2.67 $Y2=0.77
r52 14 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.63
+ $X2=2.67 $Y2=0.63
r53 13 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=0.63
+ $X2=3.365 $Y2=0.63
r54 13 14 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.2 $Y=0.63
+ $X2=2.755 $Y2=0.63
r55 11 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.77
+ $X2=2.67 $Y2=0.77
r56 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.585 $Y=0.77
+ $X2=1.895 $Y2=0.77
r57 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.73 $Y=0.685
+ $X2=1.895 $Y2=0.77
r58 7 9 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.73 $Y=0.685
+ $X2=1.73 $Y2=0.49
r59 2 20 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.275 $X2=3.365 $Y2=0.49
r60 1 9 182 $w=1.7e-07 $l=3.09354e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.275 $X2=1.73 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_LP%VGND 1 6 8 10 23 24 27
r42 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r43 21 24 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r44 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r45 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 18 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.24
+ $Y2=0
r47 18 20 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.64
+ $Y2=0
r48 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r49 13 17 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r50 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r51 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 10 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.24
+ $Y2=0
r53 10 16 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=1.68
+ $Y2=0
r54 8 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r55 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r56 8 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r57 4 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=0.085 $X2=2.24
+ $Y2=0
r58 4 6 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.24 $Y=0.085 $X2=2.24
+ $Y2=0.42
r59 1 6 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.275 $X2=2.24 $Y2=0.42
.ends

