* File: sky130_fd_sc_lp__sdfrbp_1.pxi.spice
* Created: Fri Aug 28 11:27:38 2020
* 
x_PM_SKY130_FD_SC_LP__SDFRBP_1%SCE N_SCE_M1042_g N_SCE_c_293_n N_SCE_c_294_n
+ N_SCE_c_304_n N_SCE_c_305_n N_SCE_M1000_g N_SCE_c_306_n N_SCE_c_307_n
+ N_SCE_M1020_g N_SCE_M1038_g N_SCE_c_308_n N_SCE_c_296_n N_SCE_c_309_n
+ N_SCE_c_297_n N_SCE_c_298_n SCE SCE N_SCE_c_299_n N_SCE_c_300_n N_SCE_c_317_p
+ SCE N_SCE_c_301_n PM_SKY130_FD_SC_LP__SDFRBP_1%SCE
x_PM_SKY130_FD_SC_LP__SDFRBP_1%A_27_75# N_A_27_75#_M1042_s N_A_27_75#_M1000_s
+ N_A_27_75#_c_396_n N_A_27_75#_M1029_g N_A_27_75#_M1009_g N_A_27_75#_c_397_n
+ N_A_27_75#_c_398_n N_A_27_75#_c_404_n N_A_27_75#_c_405_n N_A_27_75#_c_399_n
+ N_A_27_75#_c_400_n N_A_27_75#_c_406_n N_A_27_75#_c_407_n N_A_27_75#_c_408_n
+ N_A_27_75#_c_401_n N_A_27_75#_c_409_n PM_SKY130_FD_SC_LP__SDFRBP_1%A_27_75#
x_PM_SKY130_FD_SC_LP__SDFRBP_1%D N_D_c_478_n N_D_M1028_g N_D_M1011_g D D
+ PM_SKY130_FD_SC_LP__SDFRBP_1%D
x_PM_SKY130_FD_SC_LP__SDFRBP_1%SCD N_SCD_M1017_g N_SCD_M1030_g N_SCD_c_522_n
+ N_SCD_c_527_n SCD SCD SCD N_SCD_c_524_n PM_SKY130_FD_SC_LP__SDFRBP_1%SCD
x_PM_SKY130_FD_SC_LP__SDFRBP_1%CLK N_CLK_M1015_g N_CLK_M1023_g N_CLK_M1001_g CLK
+ CLK CLK N_CLK_c_571_n PM_SKY130_FD_SC_LP__SDFRBP_1%CLK
x_PM_SKY130_FD_SC_LP__SDFRBP_1%A_1024_367# N_A_1024_367#_M1013_d
+ N_A_1024_367#_M1006_d N_A_1024_367#_M1022_g N_A_1024_367#_c_613_n
+ N_A_1024_367#_M1033_g N_A_1024_367#_M1043_g N_A_1024_367#_M1003_g
+ N_A_1024_367#_c_615_n N_A_1024_367#_c_616_n N_A_1024_367#_c_617_n
+ N_A_1024_367#_c_618_n N_A_1024_367#_c_619_n N_A_1024_367#_c_634_p
+ N_A_1024_367#_c_639_p N_A_1024_367#_c_620_n N_A_1024_367#_c_621_n
+ N_A_1024_367#_c_622_n N_A_1024_367#_c_623_n N_A_1024_367#_c_624_n
+ N_A_1024_367#_c_631_n N_A_1024_367#_c_632_n N_A_1024_367#_c_625_n
+ N_A_1024_367#_c_626_n PM_SKY130_FD_SC_LP__SDFRBP_1%A_1024_367#
x_PM_SKY130_FD_SC_LP__SDFRBP_1%A_1374_362# N_A_1374_362#_M1004_d
+ N_A_1374_362#_M1012_d N_A_1374_362#_M1037_g N_A_1374_362#_M1026_g
+ N_A_1374_362#_c_779_n N_A_1374_362#_c_787_n N_A_1374_362#_c_780_n
+ N_A_1374_362#_c_781_n N_A_1374_362#_c_788_n N_A_1374_362#_c_789_n
+ N_A_1374_362#_c_782_n N_A_1374_362#_c_783_n
+ PM_SKY130_FD_SC_LP__SDFRBP_1%A_1374_362#
x_PM_SKY130_FD_SC_LP__SDFRBP_1%RESET_B N_RESET_B_M1021_g N_RESET_B_M1040_g
+ N_RESET_B_c_864_n N_RESET_B_c_865_n N_RESET_B_c_874_n N_RESET_B_M1010_g
+ N_RESET_B_M1014_g N_RESET_B_M1027_g N_RESET_B_c_868_n N_RESET_B_M1002_g
+ N_RESET_B_c_869_n N_RESET_B_c_870_n N_RESET_B_c_877_n N_RESET_B_c_878_n
+ N_RESET_B_c_879_n N_RESET_B_c_937_p RESET_B N_RESET_B_c_880_n
+ N_RESET_B_c_881_n N_RESET_B_c_882_n N_RESET_B_c_883_n N_RESET_B_c_884_n
+ N_RESET_B_c_885_n N_RESET_B_c_871_n PM_SKY130_FD_SC_LP__SDFRBP_1%RESET_B
x_PM_SKY130_FD_SC_LP__SDFRBP_1%A_1246_463# N_A_1246_463#_M1031_d
+ N_A_1246_463#_M1022_d N_A_1246_463#_M1010_d N_A_1246_463#_M1004_g
+ N_A_1246_463#_M1012_g N_A_1246_463#_c_1079_n N_A_1246_463#_c_1074_n
+ N_A_1246_463#_c_1103_n N_A_1246_463#_c_1081_n N_A_1246_463#_c_1075_n
+ N_A_1246_463#_c_1076_n N_A_1246_463#_c_1077_n N_A_1246_463#_c_1083_n
+ N_A_1246_463#_c_1094_n N_A_1246_463#_c_1084_n N_A_1246_463#_c_1118_n
+ PM_SKY130_FD_SC_LP__SDFRBP_1%A_1246_463#
x_PM_SKY130_FD_SC_LP__SDFRBP_1%A_840_119# N_A_840_119#_M1015_s
+ N_A_840_119#_M1001_s N_A_840_119#_M1006_g N_A_840_119#_M1013_g
+ N_A_840_119#_c_1190_n N_A_840_119#_M1018_g N_A_840_119#_c_1202_n
+ N_A_840_119#_c_1191_n N_A_840_119#_c_1192_n N_A_840_119#_c_1204_n
+ N_A_840_119#_c_1205_n N_A_840_119#_M1007_g N_A_840_119#_c_1193_n
+ N_A_840_119#_M1031_g N_A_840_119#_c_1207_n N_A_840_119#_M1041_g
+ N_A_840_119#_c_1194_n N_A_840_119#_c_1195_n N_A_840_119#_M1024_g
+ N_A_840_119#_c_1211_n N_A_840_119#_c_1212_n N_A_840_119#_c_1197_n
+ N_A_840_119#_c_1198_n N_A_840_119#_c_1199_n N_A_840_119#_c_1214_n
+ N_A_840_119#_c_1200_n PM_SKY130_FD_SC_LP__SDFRBP_1%A_840_119#
x_PM_SKY130_FD_SC_LP__SDFRBP_1%A_2002_42# N_A_2002_42#_M1005_d
+ N_A_2002_42#_M1002_d N_A_2002_42#_M1019_g N_A_2002_42#_M1032_g
+ N_A_2002_42#_c_1366_n N_A_2002_42#_c_1372_n N_A_2002_42#_c_1392_n
+ N_A_2002_42#_c_1373_n N_A_2002_42#_c_1374_n N_A_2002_42#_c_1367_n
+ N_A_2002_42#_c_1368_n N_A_2002_42#_c_1369_n N_A_2002_42#_c_1370_n
+ N_A_2002_42#_c_1376_n PM_SKY130_FD_SC_LP__SDFRBP_1%A_2002_42#
x_PM_SKY130_FD_SC_LP__SDFRBP_1%A_1812_379# N_A_1812_379#_M1043_d
+ N_A_1812_379#_M1041_d N_A_1812_379#_M1005_g N_A_1812_379#_c_1478_n
+ N_A_1812_379#_M1025_g N_A_1812_379#_c_1500_n N_A_1812_379#_c_1501_n
+ N_A_1812_379#_c_1480_n N_A_1812_379#_c_1481_n N_A_1812_379#_M1035_g
+ N_A_1812_379#_c_1483_n N_A_1812_379#_M1036_g N_A_1812_379#_M1016_g
+ N_A_1812_379#_M1034_g N_A_1812_379#_c_1485_n N_A_1812_379#_c_1486_n
+ N_A_1812_379#_c_1487_n N_A_1812_379#_c_1488_n N_A_1812_379#_c_1504_n
+ N_A_1812_379#_c_1489_n N_A_1812_379#_c_1505_n N_A_1812_379#_c_1490_n
+ N_A_1812_379#_c_1491_n N_A_1812_379#_c_1507_n N_A_1812_379#_c_1508_n
+ N_A_1812_379#_c_1492_n N_A_1812_379#_c_1493_n N_A_1812_379#_c_1494_n
+ N_A_1812_379#_c_1495_n N_A_1812_379#_c_1511_n N_A_1812_379#_c_1512_n
+ N_A_1812_379#_c_1496_n N_A_1812_379#_c_1497_n N_A_1812_379#_c_1498_n
+ PM_SKY130_FD_SC_LP__SDFRBP_1%A_1812_379#
x_PM_SKY130_FD_SC_LP__SDFRBP_1%A_2352_327# N_A_2352_327#_M1036_d
+ N_A_2352_327#_M1035_d N_A_2352_327#_c_1692_n N_A_2352_327#_M1039_g
+ N_A_2352_327#_c_1694_n N_A_2352_327#_M1008_g N_A_2352_327#_c_1695_n
+ N_A_2352_327#_c_1696_n N_A_2352_327#_c_1697_n N_A_2352_327#_c_1698_n
+ PM_SKY130_FD_SC_LP__SDFRBP_1%A_2352_327#
x_PM_SKY130_FD_SC_LP__SDFRBP_1%VPWR N_VPWR_M1000_d N_VPWR_M1017_d N_VPWR_M1001_d
+ N_VPWR_M1037_d N_VPWR_M1012_s N_VPWR_M1032_d N_VPWR_M1025_d N_VPWR_M1035_s
+ N_VPWR_M1039_d N_VPWR_c_1744_n N_VPWR_c_1745_n N_VPWR_c_1746_n N_VPWR_c_1747_n
+ N_VPWR_c_1748_n N_VPWR_c_1749_n N_VPWR_c_1750_n N_VPWR_c_1751_n
+ N_VPWR_c_1752_n N_VPWR_c_1753_n N_VPWR_c_1754_n N_VPWR_c_1755_n
+ N_VPWR_c_1756_n N_VPWR_c_1757_n N_VPWR_c_1758_n N_VPWR_c_1759_n
+ N_VPWR_c_1760_n N_VPWR_c_1761_n N_VPWR_c_1762_n N_VPWR_c_1763_n VPWR
+ N_VPWR_c_1764_n N_VPWR_c_1765_n N_VPWR_c_1766_n N_VPWR_c_1743_n
+ N_VPWR_c_1768_n N_VPWR_c_1769_n PM_SKY130_FD_SC_LP__SDFRBP_1%VPWR
x_PM_SKY130_FD_SC_LP__SDFRBP_1%A_367_491# N_A_367_491#_M1011_d
+ N_A_367_491#_M1031_s N_A_367_491#_M1028_d N_A_367_491#_M1040_d
+ N_A_367_491#_M1022_s N_A_367_491#_c_1928_n N_A_367_491#_c_1924_n
+ N_A_367_491#_c_1925_n N_A_367_491#_c_1930_n N_A_367_491#_c_1931_n
+ N_A_367_491#_c_1932_n N_A_367_491#_c_1926_n N_A_367_491#_c_1934_n
+ N_A_367_491#_c_1927_n N_A_367_491#_c_1935_n N_A_367_491#_c_1936_n
+ PM_SKY130_FD_SC_LP__SDFRBP_1%A_367_491#
x_PM_SKY130_FD_SC_LP__SDFRBP_1%Q N_Q_M1008_s N_Q_M1039_s Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__SDFRBP_1%Q
x_PM_SKY130_FD_SC_LP__SDFRBP_1%Q_N N_Q_N_M1034_d N_Q_N_M1016_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_2078_n Q_N Q_N PM_SKY130_FD_SC_LP__SDFRBP_1%Q_N
x_PM_SKY130_FD_SC_LP__SDFRBP_1%VGND N_VGND_M1042_d N_VGND_M1021_d N_VGND_M1023_d
+ N_VGND_M1018_s N_VGND_M1014_d N_VGND_M1019_d N_VGND_M1036_s N_VGND_M1008_d
+ N_VGND_c_2096_n N_VGND_c_2097_n N_VGND_c_2098_n N_VGND_c_2099_n
+ N_VGND_c_2100_n N_VGND_c_2101_n N_VGND_c_2102_n N_VGND_c_2103_n
+ N_VGND_c_2104_n N_VGND_c_2105_n N_VGND_c_2106_n N_VGND_c_2107_n
+ N_VGND_c_2108_n N_VGND_c_2109_n N_VGND_c_2110_n N_VGND_c_2111_n VGND
+ N_VGND_c_2112_n N_VGND_c_2113_n N_VGND_c_2114_n N_VGND_c_2115_n
+ N_VGND_c_2116_n N_VGND_c_2117_n N_VGND_c_2118_n N_VGND_c_2119_n
+ N_VGND_c_2120_n N_VGND_c_2121_n PM_SKY130_FD_SC_LP__SDFRBP_1%VGND
x_PM_SKY130_FD_SC_LP__SDFRBP_1%noxref_25 N_noxref_25_M1029_s N_noxref_25_M1030_d
+ N_noxref_25_c_2236_n N_noxref_25_c_2237_n N_noxref_25_c_2238_n
+ N_noxref_25_c_2239_n PM_SKY130_FD_SC_LP__SDFRBP_1%noxref_25
cc_1 VNB N_SCE_M1042_g 0.070491f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.585
cc_2 VNB N_SCE_c_293_n 0.0134183f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.7
cc_3 VNB N_SCE_c_294_n 0.00492231f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.7
cc_4 VNB N_SCE_M1038_g 0.0194437f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=0.615
cc_5 VNB N_SCE_c_296_n 0.0116412f $X=-0.19 $Y=-0.245 $X2=2.345 $Y2=1.21
cc_6 VNB N_SCE_c_297_n 0.00240003f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=1.56
cc_7 VNB N_SCE_c_298_n 0.0230204f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=1.56
cc_8 VNB N_SCE_c_299_n 0.0131662f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.7
cc_9 VNB N_SCE_c_300_n 0.0103648f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=1.395
cc_10 VNB N_SCE_c_301_n 0.00244357f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.7
cc_11 VNB N_A_27_75#_c_396_n 0.0221648f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.865
cc_12 VNB N_A_27_75#_c_397_n 0.00510363f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.775
cc_13 VNB N_A_27_75#_c_398_n 0.0198135f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=1.06
cc_14 VNB N_A_27_75#_c_399_n 0.0144004f $X=-0.19 $Y=-0.245 $X2=2.345 $Y2=1.06
cc_15 VNB N_A_27_75#_c_400_n 0.0560468f $X=-0.19 $Y=-0.245 $X2=2.345 $Y2=1.21
cc_16 VNB N_A_27_75#_c_401_n 0.0158625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_D_c_478_n 0.0731859f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.535
cc_18 VNB N_D_M1028_g 0.00341434f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.585
cc_19 VNB N_D_M1011_g 0.0193357f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.865
cc_20 VNB D 0.00355081f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.345
cc_21 VNB N_SCD_M1030_g 0.0383246f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.865
cc_22 VNB N_SCD_c_522_n 0.00240776f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.775
cc_23 VNB SCD 0.00738129f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=2.27
cc_24 VNB N_SCD_c_524_n 0.0156115f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=0.615
cc_25 VNB N_CLK_M1015_g 0.0258266f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.585
cc_26 VNB N_CLK_M1023_g 0.0204922f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.865
cc_27 VNB N_CLK_M1001_g 0.00692573f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.775
cc_28 VNB CLK 0.0359398f $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=1.21
cc_29 VNB N_CLK_c_571_n 0.0561109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_1024_367#_c_613_n 0.0547127f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.775
cc_31 VNB N_A_1024_367#_M1033_g 0.0295774f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.775
cc_32 VNB N_A_1024_367#_c_615_n 0.014546f $X=-0.19 $Y=-0.245 $X2=2.345 $Y2=1.06
cc_33 VNB N_A_1024_367#_c_616_n 6.27072e-19 $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=1.78
cc_34 VNB N_A_1024_367#_c_617_n 0.0344038f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=1.56
cc_35 VNB N_A_1024_367#_c_618_n 0.00260871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1024_367#_c_619_n 0.00253915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1024_367#_c_620_n 0.00480485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1024_367#_c_621_n 0.00434663f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.7
cc_39 VNB N_A_1024_367#_c_622_n 0.0350462f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.7
cc_40 VNB N_A_1024_367#_c_623_n 0.00583458f $X=-0.19 $Y=-0.245 $X2=2.235
+ $Y2=1.56
cc_41 VNB N_A_1024_367#_c_624_n 0.00215342f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.7
cc_42 VNB N_A_1024_367#_c_625_n 0.0168712f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.665
cc_43 VNB N_A_1024_367#_c_626_n 0.019479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1374_362#_M1026_g 0.0360929f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=2.27
cc_45 VNB N_A_1374_362#_c_779_n 0.00321052f $X=-0.19 $Y=-0.245 $X2=2.325
+ $Y2=1.21
cc_46 VNB N_A_1374_362#_c_780_n 0.0215524f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=0.615
cc_47 VNB N_A_1374_362#_c_781_n 0.0016026f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=0.615
cc_48 VNB N_A_1374_362#_c_782_n 0.00154381f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=1.78
cc_49 VNB N_A_1374_362#_c_783_n 0.00634396f $X=-0.19 $Y=-0.245 $X2=2.227
+ $Y2=1.56
cc_50 VNB N_RESET_B_M1021_g 0.0601426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_RESET_B_c_864_n 0.341702f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.345
cc_52 VNB N_RESET_B_c_865_n 0.0126405f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.775
cc_53 VNB N_RESET_B_M1014_g 0.0529632f $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=1.21
cc_54 VNB N_RESET_B_M1027_g 0.0218057f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=0.615
cc_55 VNB N_RESET_B_c_868_n 0.00422336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_RESET_B_c_869_n 0.00309655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_c_870_n 0.0211515f $X=-0.19 $Y=-0.245 $X2=2.227 $Y2=1.78
cc_58 VNB N_RESET_B_c_871_n 0.00271421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1246_463#_M1004_g 0.0397436f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=2.27
cc_60 VNB N_A_1246_463#_c_1074_n 0.00846753f $X=-0.19 $Y=-0.245 $X2=0.97
+ $Y2=2.27
cc_61 VNB N_A_1246_463#_c_1075_n 8.92097e-19 $X=-0.19 $Y=-0.245 $X2=2.227
+ $Y2=1.56
cc_62 VNB N_A_1246_463#_c_1076_n 0.00838559f $X=-0.19 $Y=-0.245 $X2=2.235
+ $Y2=1.56
cc_63 VNB N_A_1246_463#_c_1077_n 0.0277172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_840_119#_M1013_g 0.0233645f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=2.27
cc_65 VNB N_A_840_119#_c_1190_n 0.013666f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.775
cc_66 VNB N_A_840_119#_c_1191_n 0.0632462f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=0.615
cc_67 VNB N_A_840_119#_c_1192_n 0.0513917f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=0.615
cc_68 VNB N_A_840_119#_c_1193_n 0.0146382f $X=-0.19 $Y=-0.245 $X2=2.227 $Y2=1.56
cc_69 VNB N_A_840_119#_c_1194_n 0.0143881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_840_119#_c_1195_n 0.00880019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_840_119#_M1024_g 0.0510636f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.7
cc_72 VNB N_A_840_119#_c_1197_n 0.00583251f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.7
cc_73 VNB N_A_840_119#_c_1198_n 0.00428462f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.7
cc_74 VNB N_A_840_119#_c_1199_n 0.0018853f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.7
cc_75 VNB N_A_840_119#_c_1200_n 0.00140294f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.7
cc_76 VNB N_A_2002_42#_M1019_g 0.0278377f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.345
cc_77 VNB N_A_2002_42#_M1032_g 0.0114276f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=2.27
cc_78 VNB N_A_2002_42#_c_1366_n 0.00678376f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.775
cc_79 VNB N_A_2002_42#_c_1367_n 0.00373208f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=1.78
cc_80 VNB N_A_2002_42#_c_1368_n 0.00506697f $X=-0.19 $Y=-0.245 $X2=1.305
+ $Y2=1.78
cc_81 VNB N_A_2002_42#_c_1369_n 0.0299462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_2002_42#_c_1370_n 0.0137325f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_83 VNB N_A_1812_379#_c_1478_n 0.0131117f $X=-0.19 $Y=-0.245 $X2=0.97
+ $Y2=2.775
cc_84 VNB N_A_1812_379#_M1025_g 0.00460903f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.775
cc_85 VNB N_A_1812_379#_c_1480_n 0.0199409f $X=-0.19 $Y=-0.245 $X2=2.325
+ $Y2=1.395
cc_86 VNB N_A_1812_379#_c_1481_n 0.0149749f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=0.615
cc_87 VNB N_A_1812_379#_M1035_g 0.00841505f $X=-0.19 $Y=-0.245 $X2=2.345
+ $Y2=1.06
cc_88 VNB N_A_1812_379#_c_1483_n 0.02203f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=1.78
cc_89 VNB N_A_1812_379#_M1034_g 0.0229092f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_90 VNB N_A_1812_379#_c_1485_n 0.0162845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1812_379#_c_1486_n 0.00365984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1812_379#_c_1487_n 0.0299653f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.7
cc_93 VNB N_A_1812_379#_c_1488_n 0.00762525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1812_379#_c_1489_n 0.00873124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1812_379#_c_1490_n 0.00307798f $X=-0.19 $Y=-0.245 $X2=1.2
+ $Y2=1.665
cc_96 VNB N_A_1812_379#_c_1491_n 0.00855604f $X=-0.19 $Y=-0.245 $X2=1.305
+ $Y2=1.7
cc_97 VNB N_A_1812_379#_c_1492_n 0.00415648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1812_379#_c_1493_n 0.00798731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1812_379#_c_1494_n 0.00226815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1812_379#_c_1495_n 0.00135953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1812_379#_c_1496_n 0.00314557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1812_379#_c_1497_n 0.0264999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1812_379#_c_1498_n 0.0274139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2352_327#_c_1692_n 0.0383268f $X=-0.19 $Y=-0.245 $X2=0.97
+ $Y2=1.865
cc_105 VNB N_A_2352_327#_M1039_g 0.0110845f $X=-0.19 $Y=-0.245 $X2=0.97
+ $Y2=2.775
cc_106 VNB N_A_2352_327#_c_1694_n 0.0198814f $X=-0.19 $Y=-0.245 $X2=1.045
+ $Y2=2.27
cc_107 VNB N_A_2352_327#_c_1695_n 0.00796065f $X=-0.19 $Y=-0.245 $X2=1.4
+ $Y2=2.775
cc_108 VNB N_A_2352_327#_c_1696_n 0.0158086f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=1.06
cc_109 VNB N_A_2352_327#_c_1697_n 0.0357499f $X=-0.19 $Y=-0.245 $X2=0.97
+ $Y2=2.27
cc_110 VNB N_A_2352_327#_c_1698_n 2.87661e-19 $X=-0.19 $Y=-0.245 $X2=2.345
+ $Y2=1.21
cc_111 VNB N_VPWR_c_1743_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_367_491#_c_1924_n 0.00958349f $X=-0.19 $Y=-0.245 $X2=2.365
+ $Y2=0.615
cc_113 VNB N_A_367_491#_c_1925_n 0.00479741f $X=-0.19 $Y=-0.245 $X2=0.97
+ $Y2=2.27
cc_114 VNB N_A_367_491#_c_1926_n 0.00553676f $X=-0.19 $Y=-0.245 $X2=2.227
+ $Y2=1.78
cc_115 VNB N_A_367_491#_c_1927_n 0.00434751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB Q 0.0136359f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.865
cc_117 VNB Q_N 0.00777199f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.195
cc_118 VNB Q_N 0.0227731f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.345
cc_119 VNB N_Q_N_c_2078_n 0.0301157f $X=-0.19 $Y=-0.245 $X2=2.345 $Y2=1.21
cc_120 VNB N_VGND_c_2096_n 0.00863513f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.78
cc_121 VNB N_VGND_c_2097_n 0.00607943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2098_n 0.0142784f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_123 VNB N_VGND_c_2099_n 0.00882909f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.7
cc_124 VNB N_VGND_c_2100_n 0.0086398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2101_n 0.00574937f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.7
cc_126 VNB N_VGND_c_2102_n 0.00774686f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.7
cc_127 VNB N_VGND_c_2103_n 0.00879948f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.7
cc_128 VNB N_VGND_c_2104_n 0.0308765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2105_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2106_n 0.0176323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2107_n 0.00239704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2108_n 0.048766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2109_n 0.00631594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2110_n 0.0294063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2111_n 0.00452017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2112_n 0.019513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2113_n 0.0583104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2114_n 0.0516825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2115_n 0.0302681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2116_n 0.0214128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2117_n 0.716116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2118_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2119_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2120_n 0.00590529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2121_n 0.00510637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_noxref_25_c_2236_n 0.00346516f $X=-0.19 $Y=-0.245 $X2=0.97
+ $Y2=2.345
cc_147 VNB N_noxref_25_c_2237_n 0.00943229f $X=-0.19 $Y=-0.245 $X2=0.97
+ $Y2=2.775
cc_148 VNB N_noxref_25_c_2238_n 0.00391027f $X=-0.19 $Y=-0.245 $X2=1.325
+ $Y2=2.27
cc_149 VNB N_noxref_25_c_2239_n 0.00393383f $X=-0.19 $Y=-0.245 $X2=1.045
+ $Y2=2.27
cc_150 VPB N_SCE_c_293_n 0.0159295f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=1.7
cc_151 VPB N_SCE_c_294_n 0.0125399f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.7
cc_152 VPB N_SCE_c_304_n 0.0192523f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.195
cc_153 VPB N_SCE_c_305_n 0.0200329f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.345
cc_154 VPB N_SCE_c_306_n 0.021084f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=2.27
cc_155 VPB N_SCE_c_307_n 0.0154392f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=2.345
cc_156 VPB N_SCE_c_308_n 0.00664226f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.27
cc_157 VPB N_SCE_c_309_n 0.0139144f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=1.78
cc_158 VPB N_SCE_c_297_n 0.0030934f $X=-0.19 $Y=1.655 $X2=2.235 $Y2=1.56
cc_159 VPB N_SCE_c_298_n 0.00903814f $X=-0.19 $Y=1.655 $X2=2.235 $Y2=1.56
cc_160 VPB N_SCE_c_299_n 0.0151669f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.7
cc_161 VPB N_SCE_c_301_n 0.00100706f $X=-0.19 $Y=1.655 $X2=1.305 $Y2=1.7
cc_162 VPB N_A_27_75#_M1009_g 0.0192434f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=2.27
cc_163 VPB N_A_27_75#_c_398_n 0.0190153f $X=-0.19 $Y=1.655 $X2=2.365 $Y2=1.06
cc_164 VPB N_A_27_75#_c_404_n 0.0150297f $X=-0.19 $Y=1.655 $X2=2.365 $Y2=0.615
cc_165 VPB N_A_27_75#_c_405_n 0.0153049f $X=-0.19 $Y=1.655 $X2=2.365 $Y2=0.615
cc_166 VPB N_A_27_75#_c_406_n 0.0342881f $X=-0.19 $Y=1.655 $X2=2.235 $Y2=1.56
cc_167 VPB N_A_27_75#_c_407_n 0.0170194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_27_75#_c_408_n 0.030857f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_169 VPB N_A_27_75#_c_409_n 0.00266323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_D_M1028_g 0.0589909f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.585
cc_171 VPB N_SCD_M1017_g 0.0290546f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.585
cc_172 VPB N_SCD_c_522_n 0.0225815f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.775
cc_173 VPB N_SCD_c_527_n 0.015621f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=2.27
cc_174 VPB SCD 0.00929358f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=2.27
cc_175 VPB N_CLK_M1001_g 0.0255172f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.775
cc_176 VPB CLK 0.0143454f $X=-0.19 $Y=1.655 $X2=2.325 $Y2=1.21
cc_177 VPB N_A_1024_367#_M1022_g 0.0297976f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.345
cc_178 VPB N_A_1024_367#_M1003_g 0.0231454f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_1024_367#_c_621_n 0.00323267f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.7
cc_180 VPB N_A_1024_367#_c_623_n 0.0051484f $X=-0.19 $Y=1.655 $X2=2.235 $Y2=1.56
cc_181 VPB N_A_1024_367#_c_631_n 0.00564878f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_1024_367#_c_632_n 0.0332902f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.7
cc_183 VPB N_A_1024_367#_c_625_n 0.0327067f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.665
cc_184 VPB N_A_1374_362#_M1037_g 0.0185311f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.345
cc_185 VPB N_A_1374_362#_M1026_g 0.00186457f $X=-0.19 $Y=1.655 $X2=1.045
+ $Y2=2.27
cc_186 VPB N_A_1374_362#_c_779_n 0.00399028f $X=-0.19 $Y=1.655 $X2=2.325
+ $Y2=1.21
cc_187 VPB N_A_1374_362#_c_787_n 0.0626506f $X=-0.19 $Y=1.655 $X2=2.325
+ $Y2=1.395
cc_188 VPB N_A_1374_362#_c_788_n 0.00132561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1374_362#_c_789_n 0.00355404f $X=-0.19 $Y=1.655 $X2=2.345
+ $Y2=1.06
cc_190 VPB N_A_1374_362#_c_783_n 0.00205353f $X=-0.19 $Y=1.655 $X2=2.227
+ $Y2=1.56
cc_191 VPB N_RESET_B_M1021_g 0.0141715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_RESET_B_M1040_g 0.0275614f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=1.865
cc_193 VPB N_RESET_B_c_874_n 0.0166756f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.775
cc_194 VPB N_RESET_B_M1014_g 0.00964634f $X=-0.19 $Y=1.655 $X2=2.325 $Y2=1.21
cc_195 VPB N_RESET_B_M1002_g 0.0305593f $X=-0.19 $Y=1.655 $X2=2.227 $Y2=1.56
cc_196 VPB N_RESET_B_c_877_n 0.0220153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_RESET_B_c_878_n 0.00344624f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_198 VPB N_RESET_B_c_879_n 0.0128147f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_199 VPB N_RESET_B_c_880_n 0.0522016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_RESET_B_c_881_n 0.00675524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_RESET_B_c_882_n 0.0554078f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.665
cc_202 VPB N_RESET_B_c_883_n 0.00498243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_RESET_B_c_884_n 0.0311625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_RESET_B_c_885_n 0.00539788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_RESET_B_c_871_n 0.0117946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1246_463#_M1012_g 0.0205283f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=2.775
cc_207 VPB N_A_1246_463#_c_1079_n 0.00326366f $X=-0.19 $Y=1.655 $X2=2.325
+ $Y2=1.395
cc_208 VPB N_A_1246_463#_c_1074_n 0.00542445f $X=-0.19 $Y=1.655 $X2=0.97
+ $Y2=2.27
cc_209 VPB N_A_1246_463#_c_1081_n 0.00532687f $X=-0.19 $Y=1.655 $X2=1.305
+ $Y2=1.78
cc_210 VPB N_A_1246_463#_c_1077_n 0.0112995f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_1246_463#_c_1083_n 0.00410744f $X=-0.19 $Y=1.655 $X2=1.115
+ $Y2=1.58
cc_212 VPB N_A_1246_463#_c_1084_n 0.00122638f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.7
cc_213 VPB N_A_840_119#_M1006_g 0.0183579f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.345
cc_214 VPB N_A_840_119#_c_1202_n 0.0764725f $X=-0.19 $Y=1.655 $X2=2.365 $Y2=1.06
cc_215 VPB N_A_840_119#_c_1192_n 0.00797095f $X=-0.19 $Y=1.655 $X2=2.365
+ $Y2=0.615
cc_216 VPB N_A_840_119#_c_1204_n 0.0626892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_840_119#_c_1205_n 0.00989679f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.27
cc_218 VPB N_A_840_119#_M1007_g 0.0352706f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=1.78
cc_219 VPB N_A_840_119#_c_1207_n 0.178445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_840_119#_M1041_g 0.0286603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_840_119#_c_1194_n 0.0286127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_840_119#_c_1195_n 0.00365263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_840_119#_c_1211_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_840_119#_c_1212_n 0.00350191f $X=-0.19 $Y=1.655 $X2=2.235
+ $Y2=1.56
cc_225 VPB N_A_840_119#_c_1199_n 0.00105539f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.7
cc_226 VPB N_A_840_119#_c_1214_n 9.04689e-19 $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.665
cc_227 VPB N_A_2002_42#_M1032_g 0.0553269f $X=-0.19 $Y=1.655 $X2=1.045 $Y2=2.27
cc_228 VPB N_A_2002_42#_c_1372_n 0.00474457f $X=-0.19 $Y=1.655 $X2=2.325
+ $Y2=1.21
cc_229 VPB N_A_2002_42#_c_1373_n 0.00338593f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.27
cc_230 VPB N_A_2002_42#_c_1374_n 0.00274155f $X=-0.19 $Y=1.655 $X2=2.345
+ $Y2=1.06
cc_231 VPB N_A_2002_42#_c_1367_n 0.00407966f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=1.78
cc_232 VPB N_A_2002_42#_c_1376_n 0.00358816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_1812_379#_M1025_g 0.0558408f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=2.775
cc_234 VPB N_A_1812_379#_c_1500_n 0.0732492f $X=-0.19 $Y=1.655 $X2=1.4 $Y2=2.775
cc_235 VPB N_A_1812_379#_c_1501_n 0.012251f $X=-0.19 $Y=1.655 $X2=2.325 $Y2=1.21
cc_236 VPB N_A_1812_379#_M1035_g 0.0252092f $X=-0.19 $Y=1.655 $X2=2.345 $Y2=1.06
cc_237 VPB N_A_1812_379#_M1016_g 0.0221586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_1812_379#_c_1504_n 0.00731894f $X=-0.19 $Y=1.655 $X2=2.235
+ $Y2=1.395
cc_239 VPB N_A_1812_379#_c_1505_n 0.015365f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.7
cc_240 VPB N_A_1812_379#_c_1490_n 0.00297532f $X=-0.19 $Y=1.655 $X2=1.2
+ $Y2=1.665
cc_241 VPB N_A_1812_379#_c_1507_n 0.00928278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_1812_379#_c_1508_n 0.0013757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1812_379#_c_1493_n 0.00196228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_1812_379#_c_1494_n 3.17313e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_1812_379#_c_1511_n 0.00209091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_1812_379#_c_1512_n 0.0641552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_1812_379#_c_1496_n 4.76632e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_1812_379#_c_1497_n 0.00728842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_1812_379#_c_1498_n 0.00155927f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_2352_327#_M1039_g 0.022701f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.775
cc_251 VPB N_A_2352_327#_c_1696_n 0.00127343f $X=-0.19 $Y=1.655 $X2=2.365
+ $Y2=1.06
cc_252 VPB N_A_2352_327#_c_1697_n 0.00654255f $X=-0.19 $Y=1.655 $X2=0.97
+ $Y2=2.27
cc_253 VPB N_A_2352_327#_c_1698_n 0.0237644f $X=-0.19 $Y=1.655 $X2=2.345
+ $Y2=1.21
cc_254 VPB N_VPWR_c_1744_n 0.00448053f $X=-0.19 $Y=1.655 $X2=2.235 $Y2=1.56
cc_255 VPB N_VPWR_c_1745_n 0.0055721f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_256 VPB N_VPWR_c_1746_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1747_n 0.0136159f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.7
cc_258 VPB N_VPWR_c_1748_n 0.0161695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1749_n 0.0113045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1750_n 0.0121427f $X=-0.19 $Y=1.655 $X2=1.212 $Y2=1.7
cc_261 VPB N_VPWR_c_1751_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1752_n 0.0384826f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1753_n 0.00631541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1754_n 0.0405967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1755_n 0.00436584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1756_n 0.0562589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1757_n 0.00437061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1758_n 0.050608f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1759_n 0.0049622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1760_n 0.0186006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1761_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1762_n 0.0324517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1763_n 0.00436557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1764_n 0.0336194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1765_n 0.0229598f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1766_n 0.0196387f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1743_n 0.107687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1768_n 0.00375865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1769_n 0.00303699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_A_367_491#_c_1928_n 0.0121852f $X=-0.19 $Y=1.655 $X2=2.325
+ $Y2=1.395
cc_281 VPB N_A_367_491#_c_1925_n 0.00514565f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.27
cc_282 VPB N_A_367_491#_c_1930_n 0.0263059f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=1.78
cc_283 VPB N_A_367_491#_c_1931_n 0.002387f $X=-0.19 $Y=1.655 $X2=1.305 $Y2=1.78
cc_284 VPB N_A_367_491#_c_1932_n 0.0012266f $X=-0.19 $Y=1.655 $X2=2.227 $Y2=1.56
cc_285 VPB N_A_367_491#_c_1926_n 0.00884133f $X=-0.19 $Y=1.655 $X2=2.227
+ $Y2=1.78
cc_286 VPB N_A_367_491#_c_1934_n 0.00238405f $X=-0.19 $Y=1.655 $X2=1.115
+ $Y2=1.58
cc_287 VPB N_A_367_491#_c_1935_n 0.0178583f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_A_367_491#_c_1936_n 0.00382435f $X=-0.19 $Y=1.655 $X2=2.235
+ $Y2=1.56
cc_289 VPB Q 0.00753462f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=1.865
cc_290 VPB Q_N 0.0095607f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.345
cc_291 VPB Q_N 0.0535353f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=2.775
cc_292 N_SCE_M1042_g N_A_27_75#_c_397_n 0.00443261f $X=0.475 $Y=0.585 $X2=0
+ $Y2=0
cc_293 N_SCE_M1042_g N_A_27_75#_c_398_n 0.0213798f $X=0.475 $Y=0.585 $X2=0 $Y2=0
cc_294 N_SCE_c_304_n N_A_27_75#_c_398_n 0.00424163f $X=0.97 $Y=2.195 $X2=0 $Y2=0
cc_295 N_SCE_c_317_p N_A_27_75#_c_398_n 0.0208533f $X=1.14 $Y=1.7 $X2=0 $Y2=0
cc_296 N_SCE_c_294_n N_A_27_75#_c_404_n 0.00721273f $X=0.55 $Y=1.7 $X2=0 $Y2=0
cc_297 N_SCE_c_317_p N_A_27_75#_c_404_n 0.00260402f $X=1.14 $Y=1.7 $X2=0 $Y2=0
cc_298 N_SCE_M1042_g N_A_27_75#_c_399_n 0.0293433f $X=0.475 $Y=0.585 $X2=0 $Y2=0
cc_299 N_SCE_c_293_n N_A_27_75#_c_399_n 0.00750542f $X=0.895 $Y=1.7 $X2=0 $Y2=0
cc_300 N_SCE_c_299_n N_A_27_75#_c_399_n 0.00140075f $X=1.07 $Y=1.7 $X2=0 $Y2=0
cc_301 N_SCE_c_317_p N_A_27_75#_c_399_n 0.033836f $X=1.14 $Y=1.7 $X2=0 $Y2=0
cc_302 N_SCE_M1042_g N_A_27_75#_c_400_n 0.0109334f $X=0.475 $Y=0.585 $X2=0 $Y2=0
cc_303 N_SCE_c_309_n N_A_27_75#_c_400_n 0.00413039f $X=2.07 $Y=1.78 $X2=0 $Y2=0
cc_304 N_SCE_c_299_n N_A_27_75#_c_400_n 0.0133313f $X=1.07 $Y=1.7 $X2=0 $Y2=0
cc_305 N_SCE_c_317_p N_A_27_75#_c_400_n 0.00130943f $X=1.14 $Y=1.7 $X2=0 $Y2=0
cc_306 N_SCE_c_301_n N_A_27_75#_c_400_n 0.0018749f $X=1.305 $Y=1.7 $X2=0 $Y2=0
cc_307 N_SCE_c_305_n N_A_27_75#_c_406_n 0.0104806f $X=0.97 $Y=2.345 $X2=0 $Y2=0
cc_308 N_SCE_c_307_n N_A_27_75#_c_406_n 6.2413e-19 $X=1.4 $Y=2.345 $X2=0 $Y2=0
cc_309 N_SCE_c_308_n N_A_27_75#_c_406_n 0.00875086f $X=0.97 $Y=2.27 $X2=0 $Y2=0
cc_310 N_SCE_c_304_n N_A_27_75#_c_407_n 0.00491923f $X=0.97 $Y=2.195 $X2=0 $Y2=0
cc_311 N_SCE_c_306_n N_A_27_75#_c_407_n 0.0178533f $X=1.325 $Y=2.27 $X2=0 $Y2=0
cc_312 N_SCE_c_308_n N_A_27_75#_c_407_n 0.00574277f $X=0.97 $Y=2.27 $X2=0 $Y2=0
cc_313 N_SCE_c_297_n N_A_27_75#_c_407_n 0.0238511f $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_314 N_SCE_c_298_n N_A_27_75#_c_407_n 2.67229e-19 $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_315 N_SCE_c_299_n N_A_27_75#_c_407_n 0.00130086f $X=1.07 $Y=1.7 $X2=0 $Y2=0
cc_316 N_SCE_c_317_p N_A_27_75#_c_407_n 0.0853974f $X=1.14 $Y=1.7 $X2=0 $Y2=0
cc_317 N_SCE_c_309_n N_A_27_75#_c_408_n 6.08855e-19 $X=2.07 $Y=1.78 $X2=0 $Y2=0
cc_318 N_SCE_c_297_n N_A_27_75#_c_408_n 0.00230542f $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_319 N_SCE_c_298_n N_A_27_75#_c_408_n 0.0164111f $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_320 N_SCE_c_293_n N_A_27_75#_c_409_n 0.00708493f $X=0.895 $Y=1.7 $X2=0 $Y2=0
cc_321 N_SCE_c_304_n N_A_27_75#_c_409_n 0.00466026f $X=0.97 $Y=2.195 $X2=0 $Y2=0
cc_322 N_SCE_c_308_n N_A_27_75#_c_409_n 5.46893e-19 $X=0.97 $Y=2.27 $X2=0 $Y2=0
cc_323 N_SCE_c_317_p N_A_27_75#_c_409_n 0.0276796f $X=1.14 $Y=1.7 $X2=0 $Y2=0
cc_324 N_SCE_c_296_n N_D_c_478_n 0.0125751f $X=2.345 $Y=1.21 $X2=-0.19
+ $Y2=-0.245
cc_325 N_SCE_c_309_n N_D_c_478_n 0.0104488f $X=2.07 $Y=1.78 $X2=-0.19 $Y2=-0.245
cc_326 N_SCE_c_297_n N_D_c_478_n 9.92476e-19 $X=2.235 $Y=1.56 $X2=-0.19
+ $Y2=-0.245
cc_327 N_SCE_c_298_n N_D_c_478_n 0.0128787f $X=2.235 $Y=1.56 $X2=-0.19
+ $Y2=-0.245
cc_328 N_SCE_c_299_n N_D_c_478_n 0.00322691f $X=1.07 $Y=1.7 $X2=-0.19 $Y2=-0.245
cc_329 N_SCE_c_301_n N_D_c_478_n 0.00164041f $X=1.305 $Y=1.7 $X2=-0.19
+ $Y2=-0.245
cc_330 N_SCE_c_304_n N_D_M1028_g 0.002734f $X=0.97 $Y=2.195 $X2=0 $Y2=0
cc_331 N_SCE_c_306_n N_D_M1028_g 0.0630552f $X=1.325 $Y=2.27 $X2=0 $Y2=0
cc_332 N_SCE_c_309_n N_D_M1028_g 0.0131306f $X=2.07 $Y=1.78 $X2=0 $Y2=0
cc_333 N_SCE_c_297_n N_D_M1028_g 0.00124251f $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_334 N_SCE_c_298_n N_D_M1028_g 0.00737535f $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_335 N_SCE_c_299_n N_D_M1028_g 0.00613667f $X=1.07 $Y=1.7 $X2=0 $Y2=0
cc_336 N_SCE_c_301_n N_D_M1028_g 0.00227739f $X=1.305 $Y=1.7 $X2=0 $Y2=0
cc_337 N_SCE_M1038_g N_D_M1011_g 0.0216104f $X=2.365 $Y=0.615 $X2=0 $Y2=0
cc_338 N_SCE_M1038_g D 2.30294e-19 $X=2.365 $Y=0.615 $X2=0 $Y2=0
cc_339 N_SCE_c_296_n D 0.00167288f $X=2.345 $Y=1.21 $X2=0 $Y2=0
cc_340 N_SCE_c_309_n D 0.0257659f $X=2.07 $Y=1.78 $X2=0 $Y2=0
cc_341 N_SCE_c_297_n D 0.00681824f $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_342 N_SCE_c_298_n D 4.17052e-19 $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_343 N_SCE_M1038_g N_SCD_M1030_g 0.0584175f $X=2.365 $Y=0.615 $X2=0 $Y2=0
cc_344 N_SCE_c_300_n N_SCD_M1030_g 0.0113519f $X=2.235 $Y=1.395 $X2=0 $Y2=0
cc_345 N_SCE_c_297_n N_SCD_c_522_n 8.92637e-19 $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_346 N_SCE_c_296_n SCD 0.00132488f $X=2.345 $Y=1.21 $X2=0 $Y2=0
cc_347 N_SCE_c_297_n SCD 0.037411f $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_348 N_SCE_c_300_n SCD 0.00622877f $X=2.235 $Y=1.395 $X2=0 $Y2=0
cc_349 N_SCE_c_297_n N_SCD_c_524_n 2.99474e-19 $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_350 N_SCE_c_298_n N_SCD_c_524_n 0.0171212f $X=2.235 $Y=1.56 $X2=0 $Y2=0
cc_351 N_SCE_c_305_n N_VPWR_c_1744_n 0.00304035f $X=0.97 $Y=2.345 $X2=0 $Y2=0
cc_352 N_SCE_c_306_n N_VPWR_c_1744_n 0.0022993f $X=1.325 $Y=2.27 $X2=0 $Y2=0
cc_353 N_SCE_c_307_n N_VPWR_c_1744_n 0.0155746f $X=1.4 $Y=2.345 $X2=0 $Y2=0
cc_354 N_SCE_c_307_n N_VPWR_c_1752_n 0.00486043f $X=1.4 $Y=2.345 $X2=0 $Y2=0
cc_355 N_SCE_c_305_n N_VPWR_c_1764_n 0.0054895f $X=0.97 $Y=2.345 $X2=0 $Y2=0
cc_356 N_SCE_c_305_n N_VPWR_c_1743_n 0.0110654f $X=0.97 $Y=2.345 $X2=0 $Y2=0
cc_357 N_SCE_c_307_n N_VPWR_c_1743_n 0.00818711f $X=1.4 $Y=2.345 $X2=0 $Y2=0
cc_358 N_SCE_c_297_n N_A_367_491#_c_1928_n 3.46948e-19 $X=2.235 $Y=1.56 $X2=0
+ $Y2=0
cc_359 N_SCE_c_298_n N_A_367_491#_c_1928_n 4.53601e-19 $X=2.235 $Y=1.56 $X2=0
+ $Y2=0
cc_360 N_SCE_M1038_g N_A_367_491#_c_1924_n 0.0104572f $X=2.365 $Y=0.615 $X2=0
+ $Y2=0
cc_361 N_SCE_c_297_n N_A_367_491#_c_1924_n 0.00249918f $X=2.235 $Y=1.56 $X2=0
+ $Y2=0
cc_362 N_SCE_c_307_n N_A_367_491#_c_1934_n 0.00198712f $X=1.4 $Y=2.345 $X2=0
+ $Y2=0
cc_363 N_SCE_M1038_g N_A_367_491#_c_1927_n 0.00736162f $X=2.365 $Y=0.615 $X2=0
+ $Y2=0
cc_364 N_SCE_c_296_n N_A_367_491#_c_1927_n 0.00133331f $X=2.345 $Y=1.21 $X2=0
+ $Y2=0
cc_365 N_SCE_c_297_n N_A_367_491#_c_1927_n 0.0103131f $X=2.235 $Y=1.56 $X2=0
+ $Y2=0
cc_366 N_SCE_c_298_n N_A_367_491#_c_1927_n 0.00115418f $X=2.235 $Y=1.56 $X2=0
+ $Y2=0
cc_367 N_SCE_M1042_g N_VGND_c_2096_n 0.00526731f $X=0.475 $Y=0.585 $X2=0 $Y2=0
cc_368 N_SCE_M1042_g N_VGND_c_2112_n 0.00457417f $X=0.475 $Y=0.585 $X2=0 $Y2=0
cc_369 N_SCE_M1038_g N_VGND_c_2113_n 9.15902e-19 $X=2.365 $Y=0.615 $X2=0 $Y2=0
cc_370 N_SCE_M1042_g N_VGND_c_2117_n 0.00544287f $X=0.475 $Y=0.585 $X2=0 $Y2=0
cc_371 N_SCE_M1042_g N_noxref_25_c_2236_n 0.00141203f $X=0.475 $Y=0.585 $X2=0
+ $Y2=0
cc_372 N_SCE_M1038_g N_noxref_25_c_2237_n 0.0103366f $X=2.365 $Y=0.615 $X2=0
+ $Y2=0
cc_373 N_SCE_M1038_g N_noxref_25_c_2239_n 0.00105726f $X=2.365 $Y=0.615 $X2=0
+ $Y2=0
cc_374 N_A_27_75#_c_400_n N_D_c_478_n 0.00870429f $X=1.07 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_375 N_A_27_75#_M1009_g N_D_M1028_g 0.0142398f $X=2.19 $Y=2.775 $X2=0 $Y2=0
cc_376 N_A_27_75#_c_407_n N_D_M1028_g 0.0157855f $X=2.21 $Y=2.13 $X2=0 $Y2=0
cc_377 N_A_27_75#_c_408_n N_D_M1028_g 0.022163f $X=2.21 $Y=2.13 $X2=0 $Y2=0
cc_378 N_A_27_75#_c_396_n N_D_M1011_g 0.0231395f $X=1.425 $Y=0.905 $X2=0 $Y2=0
cc_379 N_A_27_75#_c_396_n D 0.00741535f $X=1.425 $Y=0.905 $X2=0 $Y2=0
cc_380 N_A_27_75#_c_399_n D 0.0206055f $X=1.07 $Y=1.07 $X2=0 $Y2=0
cc_381 N_A_27_75#_c_400_n D 0.00550757f $X=1.07 $Y=1.07 $X2=0 $Y2=0
cc_382 N_A_27_75#_M1009_g N_SCD_M1017_g 0.033131f $X=2.19 $Y=2.775 $X2=0 $Y2=0
cc_383 N_A_27_75#_c_407_n N_SCD_c_527_n 2.02046e-19 $X=2.21 $Y=2.13 $X2=0 $Y2=0
cc_384 N_A_27_75#_c_408_n N_SCD_c_527_n 0.0187608f $X=2.21 $Y=2.13 $X2=0 $Y2=0
cc_385 N_A_27_75#_c_407_n SCD 0.0142186f $X=2.21 $Y=2.13 $X2=0 $Y2=0
cc_386 N_A_27_75#_c_408_n SCD 0.00223032f $X=2.21 $Y=2.13 $X2=0 $Y2=0
cc_387 N_A_27_75#_c_406_n N_VPWR_c_1744_n 0.0247768f $X=0.755 $Y=2.6 $X2=0 $Y2=0
cc_388 N_A_27_75#_c_407_n N_VPWR_c_1744_n 0.0170992f $X=2.21 $Y=2.13 $X2=0 $Y2=0
cc_389 N_A_27_75#_M1009_g N_VPWR_c_1752_n 0.00424295f $X=2.19 $Y=2.775 $X2=0
+ $Y2=0
cc_390 N_A_27_75#_c_406_n N_VPWR_c_1764_n 0.0210467f $X=0.755 $Y=2.6 $X2=0 $Y2=0
cc_391 N_A_27_75#_M1000_s N_VPWR_c_1743_n 0.00215158f $X=0.63 $Y=2.455 $X2=0
+ $Y2=0
cc_392 N_A_27_75#_M1009_g N_VPWR_c_1743_n 0.00621075f $X=2.19 $Y=2.775 $X2=0
+ $Y2=0
cc_393 N_A_27_75#_c_406_n N_VPWR_c_1743_n 0.0125689f $X=0.755 $Y=2.6 $X2=0 $Y2=0
cc_394 N_A_27_75#_M1009_g N_A_367_491#_c_1928_n 0.0106995f $X=2.19 $Y=2.775
+ $X2=0 $Y2=0
cc_395 N_A_27_75#_c_407_n N_A_367_491#_c_1928_n 0.016799f $X=2.21 $Y=2.13 $X2=0
+ $Y2=0
cc_396 N_A_27_75#_c_408_n N_A_367_491#_c_1928_n 0.00273319f $X=2.21 $Y=2.13
+ $X2=0 $Y2=0
cc_397 N_A_27_75#_M1009_g N_A_367_491#_c_1934_n 0.0106681f $X=2.19 $Y=2.775
+ $X2=0 $Y2=0
cc_398 N_A_27_75#_c_407_n N_A_367_491#_c_1934_n 0.0273313f $X=2.21 $Y=2.13 $X2=0
+ $Y2=0
cc_399 N_A_27_75#_c_408_n N_A_367_491#_c_1934_n 0.00179489f $X=2.21 $Y=2.13
+ $X2=0 $Y2=0
cc_400 N_A_27_75#_c_396_n N_A_367_491#_c_1927_n 0.00101333f $X=1.425 $Y=0.905
+ $X2=0 $Y2=0
cc_401 N_A_27_75#_c_396_n N_VGND_c_2096_n 7.73277e-19 $X=1.425 $Y=0.905 $X2=0
+ $Y2=0
cc_402 N_A_27_75#_c_399_n N_VGND_c_2096_n 0.0141832f $X=1.07 $Y=1.07 $X2=0 $Y2=0
cc_403 N_A_27_75#_c_397_n N_VGND_c_2112_n 0.00549742f $X=0.26 $Y=0.65 $X2=0
+ $Y2=0
cc_404 N_A_27_75#_c_396_n N_VGND_c_2113_n 0.00275707f $X=1.425 $Y=0.905 $X2=0
+ $Y2=0
cc_405 N_A_27_75#_c_396_n N_VGND_c_2117_n 0.00544287f $X=1.425 $Y=0.905 $X2=0
+ $Y2=0
cc_406 N_A_27_75#_c_397_n N_VGND_c_2117_n 0.00703216f $X=0.26 $Y=0.65 $X2=0
+ $Y2=0
cc_407 N_A_27_75#_c_399_n N_noxref_25_c_2236_n 0.0152444f $X=1.07 $Y=1.07 $X2=0
+ $Y2=0
cc_408 N_A_27_75#_c_400_n N_noxref_25_c_2236_n 0.00679837f $X=1.07 $Y=1.07 $X2=0
+ $Y2=0
cc_409 N_A_27_75#_c_396_n N_noxref_25_c_2237_n 0.0138742f $X=1.425 $Y=0.905
+ $X2=0 $Y2=0
cc_410 N_D_M1028_g N_VPWR_c_1744_n 0.00295574f $X=1.76 $Y=2.775 $X2=0 $Y2=0
cc_411 N_D_M1028_g N_VPWR_c_1752_n 0.0054895f $X=1.76 $Y=2.775 $X2=0 $Y2=0
cc_412 N_D_M1028_g N_VPWR_c_1743_n 0.00987805f $X=1.76 $Y=2.775 $X2=0 $Y2=0
cc_413 N_D_M1028_g N_A_367_491#_c_1934_n 0.0124738f $X=1.76 $Y=2.775 $X2=0 $Y2=0
cc_414 N_D_M1011_g N_A_367_491#_c_1927_n 0.00894524f $X=1.935 $Y=0.615 $X2=0
+ $Y2=0
cc_415 D N_A_367_491#_c_1927_n 0.013701f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_416 N_D_M1011_g N_VGND_c_2113_n 9.15902e-19 $X=1.935 $Y=0.615 $X2=0 $Y2=0
cc_417 N_D_c_478_n N_noxref_25_c_2237_n 3.74292e-19 $X=1.76 $Y=1.595 $X2=0 $Y2=0
cc_418 N_D_M1011_g N_noxref_25_c_2237_n 0.0139954f $X=1.935 $Y=0.615 $X2=0 $Y2=0
cc_419 D N_noxref_25_c_2237_n 0.010806f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_420 D noxref_26 0.00405852f $X=1.595 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_421 N_SCD_M1030_g N_RESET_B_M1021_g 0.0330012f $X=2.725 $Y=0.615 $X2=0 $Y2=0
cc_422 SCD N_RESET_B_M1021_g 0.00144841f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_423 N_SCD_c_524_n N_RESET_B_M1021_g 0.0206795f $X=2.775 $Y=1.615 $X2=0 $Y2=0
cc_424 N_SCD_M1017_g N_RESET_B_c_880_n 0.0261242f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_425 N_SCD_c_522_n N_RESET_B_c_880_n 0.0206795f $X=2.775 $Y=1.955 $X2=0 $Y2=0
cc_426 SCD N_RESET_B_c_880_n 2.77759e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_427 N_SCD_M1017_g N_VPWR_c_1745_n 0.00334233f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_428 N_SCD_M1017_g N_VPWR_c_1752_n 0.00435799f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_429 N_SCD_M1017_g N_VPWR_c_1743_n 0.00639962f $X=2.685 $Y=2.775 $X2=0 $Y2=0
cc_430 N_SCD_M1017_g N_A_367_491#_c_1928_n 0.0158218f $X=2.685 $Y=2.775 $X2=0
+ $Y2=0
cc_431 N_SCD_c_527_n N_A_367_491#_c_1928_n 0.00365836f $X=2.775 $Y=2.12 $X2=0
+ $Y2=0
cc_432 SCD N_A_367_491#_c_1928_n 0.0249002f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_433 N_SCD_M1030_g N_A_367_491#_c_1924_n 0.0112462f $X=2.725 $Y=0.615 $X2=0
+ $Y2=0
cc_434 SCD N_A_367_491#_c_1924_n 0.0242725f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_435 N_SCD_c_524_n N_A_367_491#_c_1924_n 0.00280204f $X=2.775 $Y=1.615 $X2=0
+ $Y2=0
cc_436 N_SCD_M1017_g N_A_367_491#_c_1925_n 0.00348269f $X=2.685 $Y=2.775 $X2=0
+ $Y2=0
cc_437 N_SCD_M1030_g N_A_367_491#_c_1925_n 0.00418665f $X=2.725 $Y=0.615 $X2=0
+ $Y2=0
cc_438 SCD N_A_367_491#_c_1925_n 0.0768936f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_439 N_SCD_c_524_n N_A_367_491#_c_1925_n 0.00415403f $X=2.775 $Y=1.615 $X2=0
+ $Y2=0
cc_440 N_SCD_M1017_g N_A_367_491#_c_1934_n 0.00168777f $X=2.685 $Y=2.775 $X2=0
+ $Y2=0
cc_441 N_SCD_M1030_g N_A_367_491#_c_1927_n 0.00106536f $X=2.725 $Y=0.615 $X2=0
+ $Y2=0
cc_442 N_SCD_M1017_g N_A_367_491#_c_1935_n 6.29265e-19 $X=2.685 $Y=2.775 $X2=0
+ $Y2=0
cc_443 N_SCD_M1030_g N_VGND_c_2113_n 9.09582e-19 $X=2.725 $Y=0.615 $X2=0 $Y2=0
cc_444 N_SCD_M1030_g N_noxref_25_c_2237_n 0.00801173f $X=2.725 $Y=0.615 $X2=0
+ $Y2=0
cc_445 N_SCD_M1030_g N_noxref_25_c_2239_n 0.00674782f $X=2.725 $Y=0.615 $X2=0
+ $Y2=0
cc_446 CLK N_RESET_B_M1021_g 0.0127448f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_447 N_CLK_M1015_g N_RESET_B_c_864_n 0.0104164f $X=4.125 $Y=0.805 $X2=0 $Y2=0
cc_448 N_CLK_M1023_g N_RESET_B_c_864_n 0.0100709f $X=4.555 $Y=0.805 $X2=0 $Y2=0
cc_449 CLK N_RESET_B_c_877_n 0.0197286f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_450 CLK N_RESET_B_c_878_n 0.00848611f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_451 CLK N_RESET_B_c_880_n 0.00432175f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_452 CLK N_RESET_B_c_881_n 0.0244549f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_453 N_CLK_M1001_g N_A_840_119#_M1006_g 0.052748f $X=4.615 $Y=2.465 $X2=0
+ $Y2=0
cc_454 N_CLK_M1023_g N_A_840_119#_M1013_g 0.0171343f $X=4.555 $Y=0.805 $X2=0
+ $Y2=0
cc_455 N_CLK_c_571_n N_A_840_119#_M1013_g 0.00148f $X=4.615 $Y=1.375 $X2=0 $Y2=0
cc_456 CLK N_A_840_119#_c_1192_n 4.10738e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_457 N_CLK_c_571_n N_A_840_119#_c_1192_n 0.0263228f $X=4.615 $Y=1.375 $X2=0
+ $Y2=0
cc_458 N_CLK_M1001_g N_A_840_119#_c_1212_n 0.0127748f $X=4.615 $Y=2.465 $X2=0
+ $Y2=0
cc_459 CLK N_A_840_119#_c_1212_n 0.0282526f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_460 N_CLK_c_571_n N_A_840_119#_c_1212_n 0.00119299f $X=4.615 $Y=1.375 $X2=0
+ $Y2=0
cc_461 N_CLK_M1023_g N_A_840_119#_c_1197_n 0.00836466f $X=4.555 $Y=0.805 $X2=0
+ $Y2=0
cc_462 CLK N_A_840_119#_c_1197_n 0.0170276f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_463 N_CLK_c_571_n N_A_840_119#_c_1197_n 0.00194922f $X=4.615 $Y=1.375 $X2=0
+ $Y2=0
cc_464 N_CLK_M1023_g N_A_840_119#_c_1198_n 0.0036424f $X=4.555 $Y=0.805 $X2=0
+ $Y2=0
cc_465 CLK N_A_840_119#_c_1198_n 0.0110224f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_466 N_CLK_c_571_n N_A_840_119#_c_1198_n 9.52696e-19 $X=4.615 $Y=1.375 $X2=0
+ $Y2=0
cc_467 CLK N_A_840_119#_c_1199_n 0.0300243f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_468 N_CLK_c_571_n N_A_840_119#_c_1199_n 0.00234761f $X=4.615 $Y=1.375 $X2=0
+ $Y2=0
cc_469 N_CLK_M1001_g N_A_840_119#_c_1214_n 0.00405806f $X=4.615 $Y=2.465 $X2=0
+ $Y2=0
cc_470 CLK N_A_840_119#_c_1214_n 0.00486037f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_471 N_CLK_M1015_g N_A_840_119#_c_1200_n 3.38323e-19 $X=4.125 $Y=0.805 $X2=0
+ $Y2=0
cc_472 CLK N_A_840_119#_c_1200_n 0.0147697f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_473 N_CLK_c_571_n N_A_840_119#_c_1200_n 7.27255e-19 $X=4.615 $Y=1.375 $X2=0
+ $Y2=0
cc_474 N_CLK_M1001_g N_VPWR_c_1746_n 0.0181451f $X=4.615 $Y=2.465 $X2=0 $Y2=0
cc_475 N_CLK_M1001_g N_VPWR_c_1754_n 0.00362386f $X=4.615 $Y=2.465 $X2=0 $Y2=0
cc_476 N_CLK_M1001_g N_VPWR_c_1743_n 0.00574617f $X=4.615 $Y=2.465 $X2=0 $Y2=0
cc_477 CLK N_A_367_491#_c_1925_n 0.0412895f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_478 N_CLK_M1001_g N_A_367_491#_c_1930_n 0.01421f $X=4.615 $Y=2.465 $X2=0
+ $Y2=0
cc_479 CLK N_A_367_491#_c_1930_n 0.00590486f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_480 N_CLK_M1015_g N_VGND_c_2097_n 0.00527445f $X=4.125 $Y=0.805 $X2=0 $Y2=0
cc_481 CLK N_VGND_c_2097_n 0.00757882f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_482 N_CLK_M1023_g N_VGND_c_2098_n 0.00435905f $X=4.555 $Y=0.805 $X2=0 $Y2=0
cc_483 N_CLK_M1015_g N_VGND_c_2117_n 9.39239e-19 $X=4.125 $Y=0.805 $X2=0 $Y2=0
cc_484 N_CLK_M1023_g N_VGND_c_2117_n 9.39239e-19 $X=4.555 $Y=0.805 $X2=0 $Y2=0
cc_485 N_A_1024_367#_c_634_p N_A_1374_362#_M1004_d 0.018976f $X=9.085 $Y=0.805
+ $X2=-0.19 $Y2=-0.245
cc_486 N_A_1024_367#_M1022_g N_A_1374_362#_M1037_g 0.00236682f $X=6.155 $Y=2.525
+ $X2=0 $Y2=0
cc_487 N_A_1024_367#_M1033_g N_A_1374_362#_M1026_g 0.0692272f $X=7.075 $Y=0.805
+ $X2=0 $Y2=0
cc_488 N_A_1024_367#_c_617_n N_A_1374_362#_M1026_g 0.00202915f $X=7.61 $Y=0.34
+ $X2=0 $Y2=0
cc_489 N_A_1024_367#_c_619_n N_A_1374_362#_M1026_g 0.00477256f $X=7.695 $Y=0.72
+ $X2=0 $Y2=0
cc_490 N_A_1024_367#_c_639_p N_A_1374_362#_M1026_g 0.00241473f $X=7.78 $Y=0.805
+ $X2=0 $Y2=0
cc_491 N_A_1024_367#_c_613_n N_A_1374_362#_c_779_n 0.00464197f $X=7 $Y=1.525
+ $X2=0 $Y2=0
cc_492 N_A_1024_367#_M1033_g N_A_1374_362#_c_779_n 0.00289511f $X=7.075 $Y=0.805
+ $X2=0 $Y2=0
cc_493 N_A_1024_367#_c_613_n N_A_1374_362#_c_787_n 0.0200287f $X=7 $Y=1.525
+ $X2=0 $Y2=0
cc_494 N_A_1024_367#_c_625_n N_A_1374_362#_c_787_n 0.00236682f $X=6.025 $Y=1.525
+ $X2=0 $Y2=0
cc_495 N_A_1024_367#_c_617_n N_A_1374_362#_c_780_n 0.0105928f $X=7.61 $Y=0.34
+ $X2=0 $Y2=0
cc_496 N_A_1024_367#_c_634_p N_A_1374_362#_c_780_n 0.0652026f $X=9.085 $Y=0.805
+ $X2=0 $Y2=0
cc_497 N_A_1024_367#_c_639_p N_A_1374_362#_c_780_n 0.0113273f $X=7.78 $Y=0.805
+ $X2=0 $Y2=0
cc_498 N_A_1024_367#_M1033_g N_A_1374_362#_c_781_n 0.00856162f $X=7.075 $Y=0.805
+ $X2=0 $Y2=0
cc_499 N_A_1024_367#_c_617_n N_A_1374_362#_c_781_n 0.00448945f $X=7.61 $Y=0.34
+ $X2=0 $Y2=0
cc_500 N_A_1024_367#_c_631_n N_A_1374_362#_c_788_n 0.013305f $X=9.217 $Y=2.135
+ $X2=0 $Y2=0
cc_501 N_A_1024_367#_c_631_n N_A_1374_362#_c_789_n 0.00143309f $X=9.217 $Y=2.135
+ $X2=0 $Y2=0
cc_502 N_A_1024_367#_c_632_n N_A_1374_362#_c_789_n 2.08435e-19 $X=9.635 $Y=2.155
+ $X2=0 $Y2=0
cc_503 N_A_1024_367#_c_634_p N_A_1374_362#_c_782_n 0.013831f $X=9.085 $Y=0.805
+ $X2=0 $Y2=0
cc_504 N_A_1024_367#_c_624_n N_A_1374_362#_c_782_n 0.01992f $X=9.217 $Y=1.09
+ $X2=0 $Y2=0
cc_505 N_A_1024_367#_c_626_n N_A_1374_362#_c_782_n 0.00109f $X=9.265 $Y=1.09
+ $X2=0 $Y2=0
cc_506 N_A_1024_367#_c_621_n N_A_1374_362#_c_783_n 0.0470361f $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_507 N_A_1024_367#_c_622_n N_A_1374_362#_c_783_n 4.63584e-19 $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_508 N_A_1024_367#_M1033_g N_RESET_B_c_864_n 0.00882199f $X=7.075 $Y=0.805
+ $X2=0 $Y2=0
cc_509 N_A_1024_367#_c_616_n N_RESET_B_c_864_n 0.00450293f $X=5.32 $Y=0.845
+ $X2=0 $Y2=0
cc_510 N_A_1024_367#_c_617_n N_RESET_B_c_864_n 0.0280956f $X=7.61 $Y=0.34 $X2=0
+ $Y2=0
cc_511 N_A_1024_367#_c_618_n N_RESET_B_c_864_n 0.00420304f $X=6.175 $Y=0.34
+ $X2=0 $Y2=0
cc_512 N_A_1024_367#_c_617_n N_RESET_B_M1014_g 0.0062523f $X=7.61 $Y=0.34 $X2=0
+ $Y2=0
cc_513 N_A_1024_367#_c_619_n N_RESET_B_M1014_g 0.00728364f $X=7.695 $Y=0.72
+ $X2=0 $Y2=0
cc_514 N_A_1024_367#_c_634_p N_RESET_B_M1014_g 0.00785328f $X=9.085 $Y=0.805
+ $X2=0 $Y2=0
cc_515 N_A_1024_367#_c_639_p N_RESET_B_M1014_g 0.00261366f $X=7.78 $Y=0.805
+ $X2=0 $Y2=0
cc_516 N_A_1024_367#_M1006_d N_RESET_B_c_877_n 8.11436e-19 $X=5.12 $Y=1.835
+ $X2=0 $Y2=0
cc_517 N_A_1024_367#_M1022_g N_RESET_B_c_877_n 0.00421651f $X=6.155 $Y=2.525
+ $X2=0 $Y2=0
cc_518 N_A_1024_367#_c_613_n N_RESET_B_c_877_n 0.0060198f $X=7 $Y=1.525 $X2=0
+ $Y2=0
cc_519 N_A_1024_367#_c_623_n N_RESET_B_c_877_n 0.0679201f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_520 N_A_1024_367#_c_625_n N_RESET_B_c_877_n 0.00479087f $X=6.025 $Y=1.525
+ $X2=0 $Y2=0
cc_521 N_A_1024_367#_c_631_n N_RESET_B_c_879_n 0.0382376f $X=9.217 $Y=2.135
+ $X2=0 $Y2=0
cc_522 N_A_1024_367#_c_632_n N_RESET_B_c_879_n 0.00179783f $X=9.635 $Y=2.155
+ $X2=0 $Y2=0
cc_523 N_A_1024_367#_c_619_n N_A_1246_463#_M1004_g 8.05761e-19 $X=7.695 $Y=0.72
+ $X2=0 $Y2=0
cc_524 N_A_1024_367#_c_634_p N_A_1246_463#_M1004_g 0.0142408f $X=9.085 $Y=0.805
+ $X2=0 $Y2=0
cc_525 N_A_1024_367#_c_624_n N_A_1246_463#_M1004_g 0.00186588f $X=9.217 $Y=1.09
+ $X2=0 $Y2=0
cc_526 N_A_1024_367#_c_626_n N_A_1246_463#_M1004_g 0.0233604f $X=9.265 $Y=1.09
+ $X2=0 $Y2=0
cc_527 N_A_1024_367#_M1022_g N_A_1246_463#_c_1079_n 0.00509651f $X=6.155
+ $Y=2.525 $X2=0 $Y2=0
cc_528 N_A_1024_367#_M1022_g N_A_1246_463#_c_1074_n 8.55642e-19 $X=6.155
+ $Y=2.525 $X2=0 $Y2=0
cc_529 N_A_1024_367#_c_613_n N_A_1246_463#_c_1074_n 0.0143424f $X=7 $Y=1.525
+ $X2=0 $Y2=0
cc_530 N_A_1024_367#_M1033_g N_A_1246_463#_c_1074_n 0.00713341f $X=7.075
+ $Y=0.805 $X2=0 $Y2=0
cc_531 N_A_1024_367#_c_622_n N_A_1246_463#_c_1077_n 6.03145e-19 $X=9.265
+ $Y=1.255 $X2=0 $Y2=0
cc_532 N_A_1024_367#_c_613_n N_A_1246_463#_c_1094_n 0.00131347f $X=7 $Y=1.525
+ $X2=0 $Y2=0
cc_533 N_A_1024_367#_c_617_n N_A_1246_463#_c_1094_n 0.0116303f $X=7.61 $Y=0.34
+ $X2=0 $Y2=0
cc_534 N_A_1024_367#_c_623_n N_A_840_119#_M1006_g 0.00156669f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_535 N_A_1024_367#_c_616_n N_A_840_119#_M1013_g 5.92176e-19 $X=5.32 $Y=0.845
+ $X2=0 $Y2=0
cc_536 N_A_1024_367#_c_623_n N_A_840_119#_M1013_g 0.00161174f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_537 N_A_1024_367#_c_615_n N_A_840_119#_c_1190_n 0.00253392f $X=5.335 $Y=1.085
+ $X2=0 $Y2=0
cc_538 N_A_1024_367#_c_616_n N_A_840_119#_c_1190_n 0.00645513f $X=5.32 $Y=0.845
+ $X2=0 $Y2=0
cc_539 N_A_1024_367#_c_623_n N_A_840_119#_c_1190_n 0.00251185f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_540 N_A_1024_367#_M1022_g N_A_840_119#_c_1202_n 0.016423f $X=6.155 $Y=2.525
+ $X2=0 $Y2=0
cc_541 N_A_1024_367#_c_623_n N_A_840_119#_c_1202_n 0.019527f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_542 N_A_1024_367#_c_615_n N_A_840_119#_c_1191_n 0.00609584f $X=5.335 $Y=1.085
+ $X2=0 $Y2=0
cc_543 N_A_1024_367#_c_617_n N_A_840_119#_c_1191_n 0.00393175f $X=7.61 $Y=0.34
+ $X2=0 $Y2=0
cc_544 N_A_1024_367#_c_623_n N_A_840_119#_c_1191_n 0.0269711f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_545 N_A_1024_367#_c_625_n N_A_840_119#_c_1191_n 0.0609309f $X=6.025 $Y=1.525
+ $X2=0 $Y2=0
cc_546 N_A_1024_367#_c_623_n N_A_840_119#_c_1192_n 0.0388674f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_547 N_A_1024_367#_c_625_n N_A_840_119#_c_1192_n 0.0337552f $X=6.025 $Y=1.525
+ $X2=0 $Y2=0
cc_548 N_A_1024_367#_M1022_g N_A_840_119#_c_1204_n 0.0102906f $X=6.155 $Y=2.525
+ $X2=0 $Y2=0
cc_549 N_A_1024_367#_M1022_g N_A_840_119#_M1007_g 0.0158227f $X=6.155 $Y=2.525
+ $X2=0 $Y2=0
cc_550 N_A_1024_367#_c_613_n N_A_840_119#_M1007_g 0.00299189f $X=7 $Y=1.525
+ $X2=0 $Y2=0
cc_551 N_A_1024_367#_M1033_g N_A_840_119#_c_1193_n 0.0166217f $X=7.075 $Y=0.805
+ $X2=0 $Y2=0
cc_552 N_A_1024_367#_c_615_n N_A_840_119#_c_1193_n 0.00602089f $X=5.335 $Y=1.085
+ $X2=0 $Y2=0
cc_553 N_A_1024_367#_c_617_n N_A_840_119#_c_1193_n 0.0037178f $X=7.61 $Y=0.34
+ $X2=0 $Y2=0
cc_554 N_A_1024_367#_M1003_g N_A_840_119#_M1041_g 0.0137491f $X=9.69 $Y=2.69
+ $X2=0 $Y2=0
cc_555 N_A_1024_367#_c_621_n N_A_840_119#_M1041_g 0.00372022f $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_556 N_A_1024_367#_c_631_n N_A_840_119#_M1041_g 0.00270465f $X=9.217 $Y=2.135
+ $X2=0 $Y2=0
cc_557 N_A_1024_367#_c_632_n N_A_840_119#_M1041_g 0.00895892f $X=9.635 $Y=2.155
+ $X2=0 $Y2=0
cc_558 N_A_1024_367#_c_621_n N_A_840_119#_c_1194_n 0.0168231f $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_559 N_A_1024_367#_c_622_n N_A_840_119#_c_1194_n 0.0215454f $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_560 N_A_1024_367#_c_631_n N_A_840_119#_c_1194_n 0.00718236f $X=9.217 $Y=2.135
+ $X2=0 $Y2=0
cc_561 N_A_1024_367#_c_632_n N_A_840_119#_c_1194_n 0.0219548f $X=9.635 $Y=2.155
+ $X2=0 $Y2=0
cc_562 N_A_1024_367#_c_620_n N_A_840_119#_M1024_g 3.10126e-19 $X=9.217 $Y=1.222
+ $X2=0 $Y2=0
cc_563 N_A_1024_367#_c_621_n N_A_840_119#_M1024_g 0.00117797f $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_564 N_A_1024_367#_c_622_n N_A_840_119#_M1024_g 0.0192237f $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_565 N_A_1024_367#_c_624_n N_A_840_119#_M1024_g 3.87935e-19 $X=9.217 $Y=1.09
+ $X2=0 $Y2=0
cc_566 N_A_1024_367#_c_626_n N_A_840_119#_M1024_g 0.0186916f $X=9.265 $Y=1.09
+ $X2=0 $Y2=0
cc_567 N_A_1024_367#_c_623_n N_A_840_119#_c_1212_n 0.0124972f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_568 N_A_1024_367#_c_616_n N_A_840_119#_c_1197_n 0.00112126f $X=5.32 $Y=0.845
+ $X2=0 $Y2=0
cc_569 N_A_1024_367#_c_616_n N_A_840_119#_c_1198_n 0.00392578f $X=5.32 $Y=0.845
+ $X2=0 $Y2=0
cc_570 N_A_1024_367#_c_623_n N_A_840_119#_c_1198_n 0.0149127f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_571 N_A_1024_367#_c_623_n N_A_840_119#_c_1199_n 0.0311072f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_572 N_A_1024_367#_c_623_n N_A_840_119#_c_1214_n 0.00818288f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_573 N_A_1024_367#_M1003_g N_A_2002_42#_M1032_g 0.0171673f $X=9.69 $Y=2.69
+ $X2=0 $Y2=0
cc_574 N_A_1024_367#_c_632_n N_A_2002_42#_M1032_g 0.0096407f $X=9.635 $Y=2.155
+ $X2=0 $Y2=0
cc_575 N_A_1024_367#_c_631_n N_A_1812_379#_M1041_d 0.00753743f $X=9.217 $Y=2.135
+ $X2=0 $Y2=0
cc_576 N_A_1024_367#_M1003_g N_A_1812_379#_c_1504_n 0.0227395f $X=9.69 $Y=2.69
+ $X2=0 $Y2=0
cc_577 N_A_1024_367#_c_631_n N_A_1812_379#_c_1504_n 0.0319565f $X=9.217 $Y=2.135
+ $X2=0 $Y2=0
cc_578 N_A_1024_367#_c_632_n N_A_1812_379#_c_1504_n 0.0023049f $X=9.635 $Y=2.155
+ $X2=0 $Y2=0
cc_579 N_A_1024_367#_c_620_n N_A_1812_379#_c_1489_n 0.0292831f $X=9.217 $Y=1.222
+ $X2=0 $Y2=0
cc_580 N_A_1024_367#_c_622_n N_A_1812_379#_c_1489_n 0.0022145f $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_581 N_A_1024_367#_c_624_n N_A_1812_379#_c_1489_n 0.00696723f $X=9.217 $Y=1.09
+ $X2=0 $Y2=0
cc_582 N_A_1024_367#_c_626_n N_A_1812_379#_c_1489_n 6.17791e-19 $X=9.265 $Y=1.09
+ $X2=0 $Y2=0
cc_583 N_A_1024_367#_M1003_g N_A_1812_379#_c_1505_n 0.00404275f $X=9.69 $Y=2.69
+ $X2=0 $Y2=0
cc_584 N_A_1024_367#_c_621_n N_A_1812_379#_c_1505_n 0.0076211f $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_585 N_A_1024_367#_c_631_n N_A_1812_379#_c_1505_n 0.0273878f $X=9.217 $Y=2.135
+ $X2=0 $Y2=0
cc_586 N_A_1024_367#_c_632_n N_A_1812_379#_c_1505_n 0.00262369f $X=9.635
+ $Y=2.155 $X2=0 $Y2=0
cc_587 N_A_1024_367#_c_626_n N_A_1812_379#_c_1492_n 0.0108267f $X=9.265 $Y=1.09
+ $X2=0 $Y2=0
cc_588 N_A_1024_367#_c_621_n N_A_1812_379#_c_1493_n 0.0152705f $X=9.265 $Y=1.255
+ $X2=0 $Y2=0
cc_589 N_A_1024_367#_c_631_n N_A_1812_379#_c_1493_n 0.00949859f $X=9.217
+ $Y=2.135 $X2=0 $Y2=0
cc_590 N_A_1024_367#_c_632_n N_A_1812_379#_c_1493_n 6.29304e-19 $X=9.635
+ $Y=2.155 $X2=0 $Y2=0
cc_591 N_A_1024_367#_M1003_g N_VPWR_c_1758_n 0.00386641f $X=9.69 $Y=2.69 $X2=0
+ $Y2=0
cc_592 N_A_1024_367#_M1006_d N_VPWR_c_1743_n 0.00337311f $X=5.12 $Y=1.835 $X2=0
+ $Y2=0
cc_593 N_A_1024_367#_M1022_g N_VPWR_c_1743_n 9.39239e-19 $X=6.155 $Y=2.525 $X2=0
+ $Y2=0
cc_594 N_A_1024_367#_M1003_g N_VPWR_c_1743_n 0.00526787f $X=9.69 $Y=2.69 $X2=0
+ $Y2=0
cc_595 N_A_1024_367#_M1006_d N_A_367_491#_c_1930_n 0.00633816f $X=5.12 $Y=1.835
+ $X2=0 $Y2=0
cc_596 N_A_1024_367#_c_623_n N_A_367_491#_c_1930_n 0.0227337f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_597 N_A_1024_367#_M1022_g N_A_367_491#_c_1932_n 0.0134931f $X=6.155 $Y=2.525
+ $X2=0 $Y2=0
cc_598 N_A_1024_367#_c_613_n N_A_367_491#_c_1932_n 0.00261237f $X=7 $Y=1.525
+ $X2=0 $Y2=0
cc_599 N_A_1024_367#_c_623_n N_A_367_491#_c_1932_n 0.00768066f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_600 N_A_1024_367#_c_625_n N_A_367_491#_c_1932_n 3.09106e-19 $X=6.025 $Y=1.525
+ $X2=0 $Y2=0
cc_601 N_A_1024_367#_c_613_n N_A_367_491#_c_1926_n 0.0121695f $X=7 $Y=1.525
+ $X2=0 $Y2=0
cc_602 N_A_1024_367#_c_615_n N_A_367_491#_c_1926_n 0.0316237f $X=5.335 $Y=1.085
+ $X2=0 $Y2=0
cc_603 N_A_1024_367#_c_617_n N_A_367_491#_c_1926_n 0.00867491f $X=7.61 $Y=0.34
+ $X2=0 $Y2=0
cc_604 N_A_1024_367#_c_623_n N_A_367_491#_c_1926_n 0.0670522f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_605 N_A_1024_367#_c_625_n N_A_367_491#_c_1926_n 0.0112359f $X=6.025 $Y=1.525
+ $X2=0 $Y2=0
cc_606 N_A_1024_367#_M1022_g N_A_367_491#_c_1936_n 5.70334e-19 $X=6.155 $Y=2.525
+ $X2=0 $Y2=0
cc_607 N_A_1024_367#_c_623_n N_A_367_491#_c_1936_n 0.0193153f $X=5.985 $Y=1.805
+ $X2=0 $Y2=0
cc_608 N_A_1024_367#_c_625_n N_A_367_491#_c_1936_n 0.00161809f $X=6.025 $Y=1.525
+ $X2=0 $Y2=0
cc_609 N_A_1024_367#_c_634_p N_VGND_M1014_d 0.0101789f $X=9.085 $Y=0.805 $X2=0
+ $Y2=0
cc_610 N_A_1024_367#_c_615_n N_VGND_c_2099_n 0.0399305f $X=5.335 $Y=1.085 $X2=0
+ $Y2=0
cc_611 N_A_1024_367#_c_618_n N_VGND_c_2099_n 0.0144144f $X=6.175 $Y=0.34 $X2=0
+ $Y2=0
cc_612 N_A_1024_367#_c_623_n N_VGND_c_2099_n 0.0150621f $X=5.985 $Y=1.805 $X2=0
+ $Y2=0
cc_613 N_A_1024_367#_c_617_n N_VGND_c_2100_n 0.0140942f $X=7.61 $Y=0.34 $X2=0
+ $Y2=0
cc_614 N_A_1024_367#_c_619_n N_VGND_c_2100_n 0.00921517f $X=7.695 $Y=0.72 $X2=0
+ $Y2=0
cc_615 N_A_1024_367#_c_634_p N_VGND_c_2100_n 0.0256243f $X=9.085 $Y=0.805 $X2=0
+ $Y2=0
cc_616 N_A_1024_367#_c_616_n N_VGND_c_2106_n 0.0041894f $X=5.32 $Y=0.845 $X2=0
+ $Y2=0
cc_617 N_A_1024_367#_c_617_n N_VGND_c_2108_n 0.10385f $X=7.61 $Y=0.34 $X2=0
+ $Y2=0
cc_618 N_A_1024_367#_c_618_n N_VGND_c_2108_n 0.0115893f $X=6.175 $Y=0.34 $X2=0
+ $Y2=0
cc_619 N_A_1024_367#_c_634_p N_VGND_c_2108_n 0.00198542f $X=9.085 $Y=0.805 $X2=0
+ $Y2=0
cc_620 N_A_1024_367#_c_634_p N_VGND_c_2114_n 0.012915f $X=9.085 $Y=0.805 $X2=0
+ $Y2=0
cc_621 N_A_1024_367#_c_626_n N_VGND_c_2114_n 0.00355214f $X=9.265 $Y=1.09 $X2=0
+ $Y2=0
cc_622 N_A_1024_367#_c_616_n N_VGND_c_2117_n 0.00747125f $X=5.32 $Y=0.845 $X2=0
+ $Y2=0
cc_623 N_A_1024_367#_c_617_n N_VGND_c_2117_n 0.054012f $X=7.61 $Y=0.34 $X2=0
+ $Y2=0
cc_624 N_A_1024_367#_c_618_n N_VGND_c_2117_n 0.00583135f $X=6.175 $Y=0.34 $X2=0
+ $Y2=0
cc_625 N_A_1024_367#_c_634_p N_VGND_c_2117_n 0.0302863f $X=9.085 $Y=0.805 $X2=0
+ $Y2=0
cc_626 N_A_1024_367#_c_626_n N_VGND_c_2117_n 0.00511725f $X=9.265 $Y=1.09 $X2=0
+ $Y2=0
cc_627 N_A_1024_367#_c_619_n A_1502_119# 0.00160545f $X=7.695 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_628 N_A_1024_367#_c_639_p A_1502_119# 0.00314214f $X=7.78 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_629 N_A_1374_362#_M1026_g N_RESET_B_c_864_n 0.00882199f $X=7.435 $Y=0.805
+ $X2=0 $Y2=0
cc_630 N_A_1374_362#_M1026_g N_RESET_B_M1014_g 0.0441382f $X=7.435 $Y=0.805
+ $X2=0 $Y2=0
cc_631 N_A_1374_362#_c_780_n N_RESET_B_M1014_g 0.0136243f $X=8.745 $Y=1.177
+ $X2=0 $Y2=0
cc_632 N_A_1374_362#_c_779_n N_RESET_B_c_877_n 0.0147994f $X=7.15 $Y=1.99 $X2=0
+ $Y2=0
cc_633 N_A_1374_362#_c_787_n N_RESET_B_c_877_n 0.0127689f $X=7.15 $Y=1.99 $X2=0
+ $Y2=0
cc_634 N_A_1374_362#_M1012_d N_RESET_B_c_879_n 0.00212996f $X=8.63 $Y=1.895
+ $X2=0 $Y2=0
cc_635 N_A_1374_362#_c_788_n N_RESET_B_c_879_n 0.0144689f $X=8.787 $Y=2.002
+ $X2=0 $Y2=0
cc_636 N_A_1374_362#_c_789_n N_RESET_B_c_879_n 0.0184507f $X=8.77 $Y=2.04 $X2=0
+ $Y2=0
cc_637 N_A_1374_362#_M1037_g N_RESET_B_c_882_n 0.0124836f $X=6.945 $Y=2.525
+ $X2=0 $Y2=0
cc_638 N_A_1374_362#_c_787_n N_RESET_B_c_882_n 0.0548485f $X=7.15 $Y=1.99 $X2=0
+ $Y2=0
cc_639 N_A_1374_362#_c_783_n N_RESET_B_c_883_n 0.00163775f $X=8.787 $Y=1.875
+ $X2=0 $Y2=0
cc_640 N_A_1374_362#_c_780_n N_A_1246_463#_M1004_g 0.0154659f $X=8.745 $Y=1.177
+ $X2=0 $Y2=0
cc_641 N_A_1374_362#_c_783_n N_A_1246_463#_M1004_g 0.00208113f $X=8.787 $Y=1.875
+ $X2=0 $Y2=0
cc_642 N_A_1374_362#_c_788_n N_A_1246_463#_M1012_g 0.00207119f $X=8.787 $Y=2.002
+ $X2=0 $Y2=0
cc_643 N_A_1374_362#_M1037_g N_A_1246_463#_c_1074_n 0.00449837f $X=6.945
+ $Y=2.525 $X2=0 $Y2=0
cc_644 N_A_1374_362#_c_779_n N_A_1246_463#_c_1074_n 0.0602009f $X=7.15 $Y=1.99
+ $X2=0 $Y2=0
cc_645 N_A_1374_362#_c_787_n N_A_1246_463#_c_1074_n 0.00946436f $X=7.15 $Y=1.99
+ $X2=0 $Y2=0
cc_646 N_A_1374_362#_c_781_n N_A_1246_463#_c_1074_n 0.0181875f $X=7.245 $Y=1.177
+ $X2=0 $Y2=0
cc_647 N_A_1374_362#_M1037_g N_A_1246_463#_c_1103_n 0.00826835f $X=6.945
+ $Y=2.525 $X2=0 $Y2=0
cc_648 N_A_1374_362#_c_779_n N_A_1246_463#_c_1103_n 0.0120197f $X=7.15 $Y=1.99
+ $X2=0 $Y2=0
cc_649 N_A_1374_362#_c_787_n N_A_1246_463#_c_1103_n 0.00731357f $X=7.15 $Y=1.99
+ $X2=0 $Y2=0
cc_650 N_A_1374_362#_M1037_g N_A_1246_463#_c_1081_n 0.00136387f $X=6.945
+ $Y=2.525 $X2=0 $Y2=0
cc_651 N_A_1374_362#_M1026_g N_A_1246_463#_c_1081_n 8.08062e-19 $X=7.435
+ $Y=0.805 $X2=0 $Y2=0
cc_652 N_A_1374_362#_c_779_n N_A_1246_463#_c_1081_n 0.0334443f $X=7.15 $Y=1.99
+ $X2=0 $Y2=0
cc_653 N_A_1374_362#_c_787_n N_A_1246_463#_c_1081_n 0.00892453f $X=7.15 $Y=1.99
+ $X2=0 $Y2=0
cc_654 N_A_1374_362#_M1026_g N_A_1246_463#_c_1075_n 0.0055818f $X=7.435 $Y=0.805
+ $X2=0 $Y2=0
cc_655 N_A_1374_362#_c_779_n N_A_1246_463#_c_1075_n 0.0142126f $X=7.15 $Y=1.99
+ $X2=0 $Y2=0
cc_656 N_A_1374_362#_c_780_n N_A_1246_463#_c_1075_n 0.0148274f $X=8.745 $Y=1.177
+ $X2=0 $Y2=0
cc_657 N_A_1374_362#_c_780_n N_A_1246_463#_c_1076_n 0.0723085f $X=8.745 $Y=1.177
+ $X2=0 $Y2=0
cc_658 N_A_1374_362#_c_783_n N_A_1246_463#_c_1076_n 0.0146236f $X=8.787 $Y=1.875
+ $X2=0 $Y2=0
cc_659 N_A_1374_362#_c_780_n N_A_1246_463#_c_1077_n 0.00719495f $X=8.745
+ $Y=1.177 $X2=0 $Y2=0
cc_660 N_A_1374_362#_c_783_n N_A_1246_463#_c_1077_n 0.0112907f $X=8.787 $Y=1.875
+ $X2=0 $Y2=0
cc_661 N_A_1374_362#_M1037_g N_A_1246_463#_c_1084_n 0.00922727f $X=6.945
+ $Y=2.525 $X2=0 $Y2=0
cc_662 N_A_1374_362#_M1037_g N_A_1246_463#_c_1118_n 5.55128e-19 $X=6.945
+ $Y=2.525 $X2=0 $Y2=0
cc_663 N_A_1374_362#_M1037_g N_A_840_119#_M1007_g 0.0416539f $X=6.945 $Y=2.525
+ $X2=0 $Y2=0
cc_664 N_A_1374_362#_M1037_g N_A_840_119#_c_1207_n 0.00992967f $X=6.945 $Y=2.525
+ $X2=0 $Y2=0
cc_665 N_A_1374_362#_c_789_n N_A_840_119#_c_1207_n 0.00363004f $X=8.77 $Y=2.04
+ $X2=0 $Y2=0
cc_666 N_A_1374_362#_c_788_n N_A_840_119#_M1041_g 0.00122481f $X=8.787 $Y=2.002
+ $X2=0 $Y2=0
cc_667 N_A_1374_362#_c_789_n N_A_840_119#_M1041_g 0.0190811f $X=8.77 $Y=2.04
+ $X2=0 $Y2=0
cc_668 N_A_1374_362#_c_783_n N_A_840_119#_M1041_g 0.00159221f $X=8.787 $Y=1.875
+ $X2=0 $Y2=0
cc_669 N_A_1374_362#_c_783_n N_A_840_119#_c_1195_n 0.00327346f $X=8.787 $Y=1.875
+ $X2=0 $Y2=0
cc_670 N_A_1374_362#_c_789_n N_A_1812_379#_c_1504_n 0.023752f $X=8.77 $Y=2.04
+ $X2=0 $Y2=0
cc_671 N_A_1374_362#_M1037_g N_VPWR_c_1747_n 0.00337028f $X=6.945 $Y=2.525 $X2=0
+ $Y2=0
cc_672 N_A_1374_362#_c_788_n N_VPWR_c_1748_n 0.0429672f $X=8.787 $Y=2.002 $X2=0
+ $Y2=0
cc_673 N_A_1374_362#_c_789_n N_VPWR_c_1758_n 0.00907063f $X=8.77 $Y=2.04 $X2=0
+ $Y2=0
cc_674 N_A_1374_362#_M1037_g N_VPWR_c_1743_n 9.39239e-19 $X=6.945 $Y=2.525 $X2=0
+ $Y2=0
cc_675 N_A_1374_362#_c_789_n N_VPWR_c_1743_n 0.00795555f $X=8.77 $Y=2.04 $X2=0
+ $Y2=0
cc_676 N_A_1374_362#_M1037_g N_A_367_491#_c_1932_n 2.13429e-19 $X=6.945 $Y=2.525
+ $X2=0 $Y2=0
cc_677 N_A_1374_362#_c_787_n N_A_367_491#_c_1926_n 9.19997e-19 $X=7.15 $Y=1.99
+ $X2=0 $Y2=0
cc_678 N_RESET_B_c_864_n N_A_1246_463#_M1004_g 0.0246579f $X=7.72 $Y=0.18 $X2=0
+ $Y2=0
cc_679 N_RESET_B_M1014_g N_A_1246_463#_M1012_g 0.00245662f $X=7.795 $Y=0.805
+ $X2=0 $Y2=0
cc_680 N_RESET_B_c_879_n N_A_1246_463#_M1012_g 0.00929882f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_681 N_RESET_B_c_882_n N_A_1246_463#_M1012_g 0.00612174f $X=7.795 $Y=2.03
+ $X2=0 $Y2=0
cc_682 N_RESET_B_c_883_n N_A_1246_463#_M1012_g 8.59057e-19 $X=7.89 $Y=1.99 $X2=0
+ $Y2=0
cc_683 N_RESET_B_c_877_n N_A_1246_463#_c_1079_n 0.00868662f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_684 N_RESET_B_c_877_n N_A_1246_463#_c_1074_n 0.0191659f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_685 N_RESET_B_c_877_n N_A_1246_463#_c_1103_n 0.0146739f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_686 N_RESET_B_c_874_n N_A_1246_463#_c_1081_n 0.00334082f $X=7.605 $Y=2.24
+ $X2=0 $Y2=0
cc_687 N_RESET_B_M1014_g N_A_1246_463#_c_1081_n 0.00539843f $X=7.795 $Y=0.805
+ $X2=0 $Y2=0
cc_688 N_RESET_B_c_877_n N_A_1246_463#_c_1081_n 0.0193344f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_689 N_RESET_B_c_937_p N_A_1246_463#_c_1081_n 0.00220786f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_690 N_RESET_B_c_882_n N_A_1246_463#_c_1081_n 0.00665424f $X=7.795 $Y=2.03
+ $X2=0 $Y2=0
cc_691 N_RESET_B_c_883_n N_A_1246_463#_c_1081_n 0.0236069f $X=7.89 $Y=1.99 $X2=0
+ $Y2=0
cc_692 N_RESET_B_M1014_g N_A_1246_463#_c_1076_n 0.0111361f $X=7.795 $Y=0.805
+ $X2=0 $Y2=0
cc_693 N_RESET_B_c_877_n N_A_1246_463#_c_1076_n 0.00631543f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_694 N_RESET_B_c_879_n N_A_1246_463#_c_1076_n 0.0112508f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_695 N_RESET_B_c_937_p N_A_1246_463#_c_1076_n 0.00167348f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_696 N_RESET_B_c_882_n N_A_1246_463#_c_1076_n 0.00391783f $X=7.795 $Y=2.03
+ $X2=0 $Y2=0
cc_697 N_RESET_B_c_883_n N_A_1246_463#_c_1076_n 0.0212037f $X=7.89 $Y=1.99 $X2=0
+ $Y2=0
cc_698 N_RESET_B_M1014_g N_A_1246_463#_c_1077_n 0.0114317f $X=7.795 $Y=0.805
+ $X2=0 $Y2=0
cc_699 N_RESET_B_c_874_n N_A_1246_463#_c_1083_n 0.00473864f $X=7.605 $Y=2.24
+ $X2=0 $Y2=0
cc_700 N_RESET_B_c_877_n N_A_1246_463#_c_1083_n 0.00683731f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_701 N_RESET_B_c_937_p N_A_1246_463#_c_1083_n 0.00165837f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_702 N_RESET_B_c_882_n N_A_1246_463#_c_1083_n 0.00895701f $X=7.795 $Y=2.03
+ $X2=0 $Y2=0
cc_703 N_RESET_B_c_883_n N_A_1246_463#_c_1083_n 0.0153013f $X=7.89 $Y=1.99 $X2=0
+ $Y2=0
cc_704 N_RESET_B_c_874_n N_A_1246_463#_c_1084_n 5.56839e-19 $X=7.605 $Y=2.24
+ $X2=0 $Y2=0
cc_705 N_RESET_B_c_877_n N_A_1246_463#_c_1084_n 3.96873e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_706 N_RESET_B_c_874_n N_A_1246_463#_c_1118_n 0.0085993f $X=7.605 $Y=2.24
+ $X2=0 $Y2=0
cc_707 N_RESET_B_c_877_n N_A_840_119#_M1006_g 0.00258239f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_708 N_RESET_B_c_864_n N_A_840_119#_M1013_g 0.0104164f $X=7.72 $Y=0.18 $X2=0
+ $Y2=0
cc_709 N_RESET_B_c_864_n N_A_840_119#_c_1190_n 0.0103256f $X=7.72 $Y=0.18 $X2=0
+ $Y2=0
cc_710 N_RESET_B_c_877_n N_A_840_119#_c_1202_n 0.00273949f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_877_n N_A_840_119#_M1007_g 0.00266744f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_712 N_RESET_B_c_864_n N_A_840_119#_c_1193_n 0.00882199f $X=7.72 $Y=0.18 $X2=0
+ $Y2=0
cc_713 N_RESET_B_c_874_n N_A_840_119#_c_1207_n 0.00987666f $X=7.605 $Y=2.24
+ $X2=0 $Y2=0
cc_714 N_RESET_B_c_879_n N_A_840_119#_M1041_g 0.0127134f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_715 N_RESET_B_c_879_n N_A_840_119#_c_1194_n 0.00156333f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_716 N_RESET_B_c_877_n N_A_840_119#_c_1212_n 0.0457809f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_878_n N_A_840_119#_c_1212_n 4.62217e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_718 N_RESET_B_c_880_n N_A_840_119#_c_1212_n 0.0012151f $X=3.475 $Y=2.115
+ $X2=0 $Y2=0
cc_719 N_RESET_B_c_881_n N_A_840_119#_c_1212_n 0.00817049f $X=3.475 $Y=2.115
+ $X2=0 $Y2=0
cc_720 N_RESET_B_c_864_n N_A_840_119#_c_1197_n 0.00144731f $X=7.72 $Y=0.18 $X2=0
+ $Y2=0
cc_721 N_RESET_B_c_877_n N_A_840_119#_c_1199_n 0.00692644f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_722 N_RESET_B_c_864_n N_A_840_119#_c_1200_n 0.0030155f $X=7.72 $Y=0.18 $X2=0
+ $Y2=0
cc_723 N_RESET_B_M1027_g N_A_2002_42#_M1019_g 0.0190089f $X=10.615 $Y=0.55 $X2=0
+ $Y2=0
cc_724 N_RESET_B_c_870_n N_A_2002_42#_M1019_g 0.00183827f $X=10.62 $Y=1.52 $X2=0
+ $Y2=0
cc_725 N_RESET_B_c_868_n N_A_2002_42#_M1032_g 0.0206622f $X=10.62 $Y=1.6 $X2=0
+ $Y2=0
cc_726 N_RESET_B_M1002_g N_A_2002_42#_M1032_g 0.0154226f $X=10.72 $Y=2.755 $X2=0
+ $Y2=0
cc_727 N_RESET_B_c_870_n N_A_2002_42#_M1032_g 0.00548914f $X=10.62 $Y=1.52 $X2=0
+ $Y2=0
cc_728 N_RESET_B_c_879_n N_A_2002_42#_M1032_g 0.00130748f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_729 RESET_B N_A_2002_42#_M1032_g 0.00361565f $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_730 N_RESET_B_c_884_n N_A_2002_42#_M1032_g 0.020719f $X=10.7 $Y=2.035 $X2=0
+ $Y2=0
cc_731 N_RESET_B_c_885_n N_A_2002_42#_M1032_g 0.0126124f $X=10.7 $Y=2.035 $X2=0
+ $Y2=0
cc_732 N_RESET_B_c_869_n N_A_2002_42#_c_1366_n 0.00474034f $X=10.62 $Y=1.02
+ $X2=0 $Y2=0
cc_733 N_RESET_B_c_870_n N_A_2002_42#_c_1366_n 0.0037282f $X=10.62 $Y=1.52 $X2=0
+ $Y2=0
cc_734 N_RESET_B_M1002_g N_A_2002_42#_c_1372_n 0.00503951f $X=10.72 $Y=2.755
+ $X2=0 $Y2=0
cc_735 N_RESET_B_c_884_n N_A_2002_42#_c_1372_n 0.00300997f $X=10.7 $Y=2.035
+ $X2=0 $Y2=0
cc_736 N_RESET_B_M1002_g N_A_2002_42#_c_1392_n 0.00357671f $X=10.72 $Y=2.755
+ $X2=0 $Y2=0
cc_737 N_RESET_B_c_871_n N_A_2002_42#_c_1374_n 0.00422048f $X=10.7 $Y=1.87 $X2=0
+ $Y2=0
cc_738 N_RESET_B_c_870_n N_A_2002_42#_c_1368_n 8.50731e-19 $X=10.62 $Y=1.52
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_870_n N_A_2002_42#_c_1369_n 0.020653f $X=10.62 $Y=1.52 $X2=0
+ $Y2=0
cc_740 N_RESET_B_M1027_g N_A_2002_42#_c_1370_n 0.0100326f $X=10.615 $Y=0.55
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_869_n N_A_2002_42#_c_1370_n 0.00131805f $X=10.62 $Y=1.02
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_870_n N_A_2002_42#_c_1370_n 0.00246325f $X=10.62 $Y=1.52
+ $X2=0 $Y2=0
cc_743 N_RESET_B_M1002_g N_A_2002_42#_c_1376_n 0.00349481f $X=10.72 $Y=2.755
+ $X2=0 $Y2=0
cc_744 RESET_B N_A_2002_42#_c_1376_n 8.53555e-19 $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_745 N_RESET_B_c_884_n N_A_2002_42#_c_1376_n 0.00203249f $X=10.7 $Y=2.035
+ $X2=0 $Y2=0
cc_746 N_RESET_B_c_885_n N_A_2002_42#_c_1376_n 0.0252204f $X=10.7 $Y=2.035 $X2=0
+ $Y2=0
cc_747 N_RESET_B_c_871_n N_A_2002_42#_c_1376_n 2.7054e-19 $X=10.7 $Y=1.87 $X2=0
+ $Y2=0
cc_748 N_RESET_B_c_879_n N_A_1812_379#_M1041_d 0.00129571f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_749 N_RESET_B_M1027_g N_A_1812_379#_c_1478_n 0.00388812f $X=10.615 $Y=0.55
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_869_n N_A_1812_379#_c_1478_n 0.0159777f $X=10.62 $Y=1.02
+ $X2=0 $Y2=0
cc_751 N_RESET_B_M1002_g N_A_1812_379#_M1025_g 0.0216529f $X=10.72 $Y=2.755
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_870_n N_A_1812_379#_M1025_g 0.0112444f $X=10.62 $Y=1.52 $X2=0
+ $Y2=0
cc_753 N_RESET_B_c_884_n N_A_1812_379#_M1025_g 0.0203599f $X=10.7 $Y=2.035 $X2=0
+ $Y2=0
cc_754 N_RESET_B_c_885_n N_A_1812_379#_M1025_g 2.97558e-19 $X=10.7 $Y=2.035
+ $X2=0 $Y2=0
cc_755 N_RESET_B_M1027_g N_A_1812_379#_c_1485_n 0.0429647f $X=10.615 $Y=0.55
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_879_n N_A_1812_379#_c_1504_n 0.00933414f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_879_n N_A_1812_379#_c_1505_n 0.0165161f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_758 RESET_B N_A_1812_379#_c_1505_n 0.00238569f $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_759 N_RESET_B_c_885_n N_A_1812_379#_c_1505_n 0.0229718f $X=10.7 $Y=2.035
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_868_n N_A_1812_379#_c_1490_n 3.59463e-19 $X=10.62 $Y=1.6
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_879_n N_A_1812_379#_c_1490_n 0.00460976f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_762 RESET_B N_A_1812_379#_c_1490_n 0.00355947f $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_763 N_RESET_B_c_885_n N_A_1812_379#_c_1490_n 0.0186871f $X=10.7 $Y=2.035
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_870_n N_A_1812_379#_c_1491_n 0.00313352f $X=10.62 $Y=1.52
+ $X2=0 $Y2=0
cc_765 N_RESET_B_c_884_n N_A_1812_379#_c_1491_n 0.00433242f $X=10.7 $Y=2.035
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_885_n N_A_1812_379#_c_1491_n 0.00491336f $X=10.7 $Y=2.035
+ $X2=0 $Y2=0
cc_767 N_RESET_B_c_879_n N_A_1812_379#_c_1493_n 0.0089057f $X=10.175 $Y=2.035
+ $X2=0 $Y2=0
cc_768 N_RESET_B_c_868_n N_A_1812_379#_c_1494_n 0.00249728f $X=10.62 $Y=1.6
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_870_n N_A_1812_379#_c_1494_n 0.00495741f $X=10.62 $Y=1.52
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_885_n N_A_1812_379#_c_1494_n 0.0120861f $X=10.7 $Y=2.035
+ $X2=0 $Y2=0
cc_771 N_RESET_B_c_871_n N_A_1812_379#_c_1494_n 0.00453566f $X=10.7 $Y=1.87
+ $X2=0 $Y2=0
cc_772 N_RESET_B_c_870_n N_A_1812_379#_c_1495_n 7.39192e-19 $X=10.62 $Y=1.52
+ $X2=0 $Y2=0
cc_773 N_RESET_B_c_870_n N_A_1812_379#_c_1498_n 0.0159777f $X=10.62 $Y=1.52
+ $X2=0 $Y2=0
cc_774 N_RESET_B_c_879_n N_VPWR_M1012_s 0.00170757f $X=10.175 $Y=2.035 $X2=0
+ $Y2=0
cc_775 N_RESET_B_M1040_g N_VPWR_c_1745_n 0.00486065f $X=3.225 $Y=2.775 $X2=0
+ $Y2=0
cc_776 N_RESET_B_c_874_n N_VPWR_c_1747_n 0.00463903f $X=7.605 $Y=2.24 $X2=0
+ $Y2=0
cc_777 N_RESET_B_c_874_n N_VPWR_c_1748_n 0.00519476f $X=7.605 $Y=2.24 $X2=0
+ $Y2=0
cc_778 N_RESET_B_c_879_n N_VPWR_c_1748_n 0.0215432f $X=10.175 $Y=2.035 $X2=0
+ $Y2=0
cc_779 N_RESET_B_c_937_p N_VPWR_c_1748_n 6.69218e-19 $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_780 N_RESET_B_c_882_n N_VPWR_c_1748_n 0.00192009f $X=7.795 $Y=2.03 $X2=0
+ $Y2=0
cc_781 N_RESET_B_c_883_n N_VPWR_c_1748_n 0.0211499f $X=7.89 $Y=1.99 $X2=0 $Y2=0
cc_782 N_RESET_B_M1002_g N_VPWR_c_1749_n 0.00469162f $X=10.72 $Y=2.755 $X2=0
+ $Y2=0
cc_783 RESET_B N_VPWR_c_1749_n 8.57425e-19 $X=10.235 $Y=1.95 $X2=0 $Y2=0
cc_784 N_RESET_B_c_884_n N_VPWR_c_1749_n 0.00168792f $X=10.7 $Y=2.035 $X2=0
+ $Y2=0
cc_785 N_RESET_B_c_885_n N_VPWR_c_1749_n 0.0111193f $X=10.7 $Y=2.035 $X2=0 $Y2=0
cc_786 N_RESET_B_M1040_g N_VPWR_c_1754_n 0.0042418f $X=3.225 $Y=2.775 $X2=0
+ $Y2=0
cc_787 N_RESET_B_M1002_g N_VPWR_c_1760_n 0.00461195f $X=10.72 $Y=2.755 $X2=0
+ $Y2=0
cc_788 N_RESET_B_M1040_g N_VPWR_c_1743_n 0.00743583f $X=3.225 $Y=2.775 $X2=0
+ $Y2=0
cc_789 N_RESET_B_c_874_n N_VPWR_c_1743_n 9.39239e-19 $X=7.605 $Y=2.24 $X2=0
+ $Y2=0
cc_790 N_RESET_B_M1002_g N_VPWR_c_1743_n 0.00907238f $X=10.72 $Y=2.755 $X2=0
+ $Y2=0
cc_791 N_RESET_B_M1021_g N_A_367_491#_c_1924_n 0.0125196f $X=3.225 $Y=0.615
+ $X2=0 $Y2=0
cc_792 N_RESET_B_M1021_g N_A_367_491#_c_1925_n 0.0303891f $X=3.225 $Y=0.615
+ $X2=0 $Y2=0
cc_793 N_RESET_B_M1040_g N_A_367_491#_c_1925_n 0.00534244f $X=3.225 $Y=2.775
+ $X2=0 $Y2=0
cc_794 N_RESET_B_c_878_n N_A_367_491#_c_1925_n 0.00236242f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_795 N_RESET_B_c_880_n N_A_367_491#_c_1925_n 0.00840091f $X=3.475 $Y=2.115
+ $X2=0 $Y2=0
cc_796 N_RESET_B_c_881_n N_A_367_491#_c_1925_n 0.0226939f $X=3.475 $Y=2.115
+ $X2=0 $Y2=0
cc_797 N_RESET_B_c_877_n N_A_367_491#_c_1930_n 0.0308685f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_878_n N_A_367_491#_c_1930_n 7.71213e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_799 N_RESET_B_c_880_n N_A_367_491#_c_1930_n 7.82525e-19 $X=3.475 $Y=2.115
+ $X2=0 $Y2=0
cc_800 N_RESET_B_c_881_n N_A_367_491#_c_1930_n 0.0105736f $X=3.475 $Y=2.115
+ $X2=0 $Y2=0
cc_801 N_RESET_B_M1040_g N_A_367_491#_c_1931_n 0.0166122f $X=3.225 $Y=2.775
+ $X2=0 $Y2=0
cc_802 N_RESET_B_c_878_n N_A_367_491#_c_1931_n 9.28705e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_803 N_RESET_B_c_880_n N_A_367_491#_c_1931_n 0.00871367f $X=3.475 $Y=2.115
+ $X2=0 $Y2=0
cc_804 N_RESET_B_c_881_n N_A_367_491#_c_1931_n 0.0179037f $X=3.475 $Y=2.115
+ $X2=0 $Y2=0
cc_805 N_RESET_B_c_877_n N_A_367_491#_c_1932_n 0.011966f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_806 N_RESET_B_c_877_n N_A_367_491#_c_1926_n 0.0159774f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_807 N_RESET_B_M1040_g N_A_367_491#_c_1935_n 0.00648897f $X=3.225 $Y=2.775
+ $X2=0 $Y2=0
cc_808 N_RESET_B_c_877_n N_A_367_491#_c_1936_n 0.00779817f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_809 N_RESET_B_M1021_g N_VGND_c_2097_n 0.00657535f $X=3.225 $Y=0.615 $X2=0
+ $Y2=0
cc_810 N_RESET_B_c_864_n N_VGND_c_2097_n 0.0182194f $X=7.72 $Y=0.18 $X2=0 $Y2=0
cc_811 N_RESET_B_c_865_n N_VGND_c_2097_n 0.00388727f $X=3.3 $Y=0.18 $X2=0 $Y2=0
cc_812 N_RESET_B_c_864_n N_VGND_c_2098_n 0.0246905f $X=7.72 $Y=0.18 $X2=0 $Y2=0
cc_813 N_RESET_B_c_864_n N_VGND_c_2099_n 0.016885f $X=7.72 $Y=0.18 $X2=0 $Y2=0
cc_814 N_RESET_B_c_864_n N_VGND_c_2100_n 0.0078465f $X=7.72 $Y=0.18 $X2=0 $Y2=0
cc_815 N_RESET_B_M1027_g N_VGND_c_2101_n 0.00948771f $X=10.615 $Y=0.55 $X2=0
+ $Y2=0
cc_816 N_RESET_B_c_864_n N_VGND_c_2104_n 0.0356412f $X=7.72 $Y=0.18 $X2=0 $Y2=0
cc_817 N_RESET_B_c_864_n N_VGND_c_2106_n 0.0202037f $X=7.72 $Y=0.18 $X2=0 $Y2=0
cc_818 N_RESET_B_c_864_n N_VGND_c_2108_n 0.0448727f $X=7.72 $Y=0.18 $X2=0 $Y2=0
cc_819 N_RESET_B_c_865_n N_VGND_c_2113_n 0.00486043f $X=3.3 $Y=0.18 $X2=0 $Y2=0
cc_820 N_RESET_B_M1027_g N_VGND_c_2115_n 0.00438567f $X=10.615 $Y=0.55 $X2=0
+ $Y2=0
cc_821 N_RESET_B_c_864_n N_VGND_c_2117_n 0.120257f $X=7.72 $Y=0.18 $X2=0 $Y2=0
cc_822 N_RESET_B_c_865_n N_VGND_c_2117_n 0.00803016f $X=3.3 $Y=0.18 $X2=0 $Y2=0
cc_823 N_RESET_B_M1027_g N_VGND_c_2117_n 0.00788543f $X=10.615 $Y=0.55 $X2=0
+ $Y2=0
cc_824 N_RESET_B_M1021_g N_noxref_25_c_2239_n 0.00310474f $X=3.225 $Y=0.615
+ $X2=0 $Y2=0
cc_825 N_A_1246_463#_c_1079_n N_A_840_119#_c_1202_n 4.04116e-19 $X=6.725
+ $Y=2.635 $X2=0 $Y2=0
cc_826 N_A_1246_463#_c_1079_n N_A_840_119#_c_1204_n 0.00377074f $X=6.725
+ $Y=2.635 $X2=0 $Y2=0
cc_827 N_A_1246_463#_c_1079_n N_A_840_119#_M1007_g 0.0126499f $X=6.725 $Y=2.635
+ $X2=0 $Y2=0
cc_828 N_A_1246_463#_c_1074_n N_A_840_119#_M1007_g 0.00111222f $X=6.81 $Y=2.335
+ $X2=0 $Y2=0
cc_829 N_A_1246_463#_c_1084_n N_A_840_119#_M1007_g 0.00485082f $X=6.815 $Y=2.555
+ $X2=0 $Y2=0
cc_830 N_A_1246_463#_c_1074_n N_A_840_119#_c_1193_n 0.0022109f $X=6.81 $Y=2.335
+ $X2=0 $Y2=0
cc_831 N_A_1246_463#_M1012_g N_A_840_119#_c_1207_n 0.0104164f $X=8.555 $Y=2.315
+ $X2=0 $Y2=0
cc_832 N_A_1246_463#_c_1103_n N_A_840_119#_c_1207_n 0.00193378f $X=7.425 $Y=2.43
+ $X2=0 $Y2=0
cc_833 N_A_1246_463#_c_1083_n N_A_840_119#_c_1207_n 0.00558975f $X=7.82 $Y=2.52
+ $X2=0 $Y2=0
cc_834 N_A_1246_463#_c_1084_n N_A_840_119#_c_1207_n 0.00257797f $X=6.815
+ $Y=2.555 $X2=0 $Y2=0
cc_835 N_A_1246_463#_c_1118_n N_A_840_119#_c_1207_n 0.0021936f $X=7.425 $Y=2.335
+ $X2=0 $Y2=0
cc_836 N_A_1246_463#_M1012_g N_A_840_119#_M1041_g 0.0112486f $X=8.555 $Y=2.315
+ $X2=0 $Y2=0
cc_837 N_A_1246_463#_c_1077_n N_A_840_119#_c_1195_n 0.0112486f $X=8.41 $Y=1.555
+ $X2=0 $Y2=0
cc_838 N_A_1246_463#_c_1103_n N_VPWR_M1037_d 0.00697033f $X=7.425 $Y=2.43 $X2=0
+ $Y2=0
cc_839 N_A_1246_463#_c_1081_n N_VPWR_M1037_d 2.64675e-19 $X=7.515 $Y=2.335 $X2=0
+ $Y2=0
cc_840 N_A_1246_463#_c_1118_n N_VPWR_M1037_d 4.55983e-19 $X=7.425 $Y=2.335 $X2=0
+ $Y2=0
cc_841 N_A_1246_463#_c_1103_n N_VPWR_c_1747_n 0.0255129f $X=7.425 $Y=2.43 $X2=0
+ $Y2=0
cc_842 N_A_1246_463#_c_1084_n N_VPWR_c_1747_n 0.00501406f $X=6.815 $Y=2.555
+ $X2=0 $Y2=0
cc_843 N_A_1246_463#_M1012_g N_VPWR_c_1748_n 0.00646507f $X=8.555 $Y=2.315 $X2=0
+ $Y2=0
cc_844 N_A_1246_463#_c_1081_n N_VPWR_c_1748_n 0.0042563f $X=7.515 $Y=2.335 $X2=0
+ $Y2=0
cc_845 N_A_1246_463#_c_1076_n N_VPWR_c_1748_n 0.0136664f $X=8.41 $Y=1.555 $X2=0
+ $Y2=0
cc_846 N_A_1246_463#_c_1077_n N_VPWR_c_1748_n 0.00601524f $X=8.41 $Y=1.555 $X2=0
+ $Y2=0
cc_847 N_A_1246_463#_c_1083_n N_VPWR_c_1748_n 0.0213452f $X=7.82 $Y=2.52 $X2=0
+ $Y2=0
cc_848 N_A_1246_463#_c_1079_n N_VPWR_c_1756_n 0.0113548f $X=6.725 $Y=2.635 $X2=0
+ $Y2=0
cc_849 N_A_1246_463#_c_1084_n N_VPWR_c_1756_n 0.00423883f $X=6.815 $Y=2.555
+ $X2=0 $Y2=0
cc_850 N_A_1246_463#_c_1083_n N_VPWR_c_1765_n 0.00635792f $X=7.82 $Y=2.52 $X2=0
+ $Y2=0
cc_851 N_A_1246_463#_c_1118_n N_VPWR_c_1765_n 3.42346e-19 $X=7.425 $Y=2.335
+ $X2=0 $Y2=0
cc_852 N_A_1246_463#_M1012_g N_VPWR_c_1743_n 9.39239e-19 $X=8.555 $Y=2.315 $X2=0
+ $Y2=0
cc_853 N_A_1246_463#_c_1079_n N_VPWR_c_1743_n 0.0138069f $X=6.725 $Y=2.635 $X2=0
+ $Y2=0
cc_854 N_A_1246_463#_c_1103_n N_VPWR_c_1743_n 0.00686979f $X=7.425 $Y=2.43 $X2=0
+ $Y2=0
cc_855 N_A_1246_463#_c_1083_n N_VPWR_c_1743_n 0.00962807f $X=7.82 $Y=2.52 $X2=0
+ $Y2=0
cc_856 N_A_1246_463#_c_1084_n N_VPWR_c_1743_n 0.00502303f $X=6.815 $Y=2.555
+ $X2=0 $Y2=0
cc_857 N_A_1246_463#_c_1118_n N_VPWR_c_1743_n 0.00615122f $X=7.425 $Y=2.335
+ $X2=0 $Y2=0
cc_858 N_A_1246_463#_M1022_d N_A_367_491#_c_1932_n 0.00180549f $X=6.23 $Y=2.315
+ $X2=0 $Y2=0
cc_859 N_A_1246_463#_c_1079_n N_A_367_491#_c_1932_n 0.0147392f $X=6.725 $Y=2.635
+ $X2=0 $Y2=0
cc_860 N_A_1246_463#_c_1074_n N_A_367_491#_c_1932_n 0.0113861f $X=6.81 $Y=2.335
+ $X2=0 $Y2=0
cc_861 N_A_1246_463#_c_1074_n N_A_367_491#_c_1926_n 0.0711159f $X=6.81 $Y=2.335
+ $X2=0 $Y2=0
cc_862 N_A_1246_463#_c_1084_n A_1332_463# 0.00208311f $X=6.815 $Y=2.555
+ $X2=-0.19 $Y2=-0.245
cc_863 N_A_1246_463#_M1004_g N_VGND_c_2100_n 0.00936599f $X=8.455 $Y=0.66 $X2=0
+ $Y2=0
cc_864 N_A_1246_463#_M1004_g N_VGND_c_2114_n 0.00355322f $X=8.455 $Y=0.66 $X2=0
+ $Y2=0
cc_865 N_A_1246_463#_M1004_g N_VGND_c_2117_n 0.00517216f $X=8.455 $Y=0.66 $X2=0
+ $Y2=0
cc_866 N_A_840_119#_M1024_g N_A_2002_42#_M1019_g 0.0737658f $X=9.725 $Y=0.55
+ $X2=0 $Y2=0
cc_867 N_A_840_119#_M1024_g N_A_2002_42#_M1032_g 0.010723f $X=9.725 $Y=0.55
+ $X2=0 $Y2=0
cc_868 N_A_840_119#_M1024_g N_A_2002_42#_c_1368_n 0.00108253f $X=9.725 $Y=0.55
+ $X2=0 $Y2=0
cc_869 N_A_840_119#_M1041_g N_A_1812_379#_c_1504_n 0.00489308f $X=8.985 $Y=2.315
+ $X2=0 $Y2=0
cc_870 N_A_840_119#_c_1194_n N_A_1812_379#_c_1489_n 6.09738e-19 $X=9.65 $Y=1.705
+ $X2=0 $Y2=0
cc_871 N_A_840_119#_M1024_g N_A_1812_379#_c_1489_n 0.0150317f $X=9.725 $Y=0.55
+ $X2=0 $Y2=0
cc_872 N_A_840_119#_c_1194_n N_A_1812_379#_c_1505_n 7.77711e-19 $X=9.65 $Y=1.705
+ $X2=0 $Y2=0
cc_873 N_A_840_119#_c_1194_n N_A_1812_379#_c_1492_n 0.00286811f $X=9.65 $Y=1.705
+ $X2=0 $Y2=0
cc_874 N_A_840_119#_M1024_g N_A_1812_379#_c_1492_n 0.0136999f $X=9.725 $Y=0.55
+ $X2=0 $Y2=0
cc_875 N_A_840_119#_c_1194_n N_A_1812_379#_c_1493_n 0.00812139f $X=9.65 $Y=1.705
+ $X2=0 $Y2=0
cc_876 N_A_840_119#_M1024_g N_A_1812_379#_c_1493_n 0.00554251f $X=9.725 $Y=0.55
+ $X2=0 $Y2=0
cc_877 N_A_840_119#_c_1212_n N_VPWR_M1001_d 0.00517466f $X=4.825 $Y=2.082 $X2=0
+ $Y2=0
cc_878 N_A_840_119#_c_1214_n N_VPWR_M1001_d 0.00129419f $X=4.91 $Y=1.95 $X2=0
+ $Y2=0
cc_879 N_A_840_119#_M1006_g N_VPWR_c_1746_n 0.0110094f $X=5.045 $Y=2.465 $X2=0
+ $Y2=0
cc_880 N_A_840_119#_c_1202_n N_VPWR_c_1746_n 0.00253831f $X=5.535 $Y=3.075 $X2=0
+ $Y2=0
cc_881 N_A_840_119#_M1007_g N_VPWR_c_1747_n 0.00614754f $X=6.585 $Y=2.525 $X2=0
+ $Y2=0
cc_882 N_A_840_119#_c_1207_n N_VPWR_c_1747_n 0.0252266f $X=8.91 $Y=3.15 $X2=0
+ $Y2=0
cc_883 N_A_840_119#_c_1207_n N_VPWR_c_1748_n 0.0203716f $X=8.91 $Y=3.15 $X2=0
+ $Y2=0
cc_884 N_A_840_119#_M1041_g N_VPWR_c_1748_n 0.00452821f $X=8.985 $Y=2.315 $X2=0
+ $Y2=0
cc_885 N_A_840_119#_M1006_g N_VPWR_c_1756_n 0.00362386f $X=5.045 $Y=2.465 $X2=0
+ $Y2=0
cc_886 N_A_840_119#_c_1205_n N_VPWR_c_1756_n 0.0451203f $X=5.61 $Y=3.15 $X2=0
+ $Y2=0
cc_887 N_A_840_119#_c_1207_n N_VPWR_c_1758_n 0.0179991f $X=8.91 $Y=3.15 $X2=0
+ $Y2=0
cc_888 N_A_840_119#_c_1207_n N_VPWR_c_1765_n 0.0255036f $X=8.91 $Y=3.15 $X2=0
+ $Y2=0
cc_889 N_A_840_119#_M1001_s N_VPWR_c_1743_n 0.00340169f $X=4.275 $Y=1.835 $X2=0
+ $Y2=0
cc_890 N_A_840_119#_M1006_g N_VPWR_c_1743_n 0.00450596f $X=5.045 $Y=2.465 $X2=0
+ $Y2=0
cc_891 N_A_840_119#_c_1204_n N_VPWR_c_1743_n 0.0262432f $X=6.51 $Y=3.15 $X2=0
+ $Y2=0
cc_892 N_A_840_119#_c_1205_n N_VPWR_c_1743_n 0.00551146f $X=5.61 $Y=3.15 $X2=0
+ $Y2=0
cc_893 N_A_840_119#_c_1207_n N_VPWR_c_1743_n 0.0647516f $X=8.91 $Y=3.15 $X2=0
+ $Y2=0
cc_894 N_A_840_119#_c_1211_n N_VPWR_c_1743_n 0.00412439f $X=6.585 $Y=3.15 $X2=0
+ $Y2=0
cc_895 N_A_840_119#_M1001_s N_A_367_491#_c_1930_n 0.00713304f $X=4.275 $Y=1.835
+ $X2=0 $Y2=0
cc_896 N_A_840_119#_M1006_g N_A_367_491#_c_1930_n 0.0128009f $X=5.045 $Y=2.465
+ $X2=0 $Y2=0
cc_897 N_A_840_119#_c_1202_n N_A_367_491#_c_1930_n 0.0137053f $X=5.535 $Y=3.075
+ $X2=0 $Y2=0
cc_898 N_A_840_119#_c_1204_n N_A_367_491#_c_1930_n 0.00124696f $X=6.51 $Y=3.15
+ $X2=0 $Y2=0
cc_899 N_A_840_119#_c_1212_n N_A_367_491#_c_1930_n 0.030975f $X=4.825 $Y=2.082
+ $X2=0 $Y2=0
cc_900 N_A_840_119#_M1007_g N_A_367_491#_c_1932_n 0.00313167f $X=6.585 $Y=2.525
+ $X2=0 $Y2=0
cc_901 N_A_840_119#_c_1191_n N_A_367_491#_c_1926_n 0.010413f $X=6.57 $Y=1.165
+ $X2=0 $Y2=0
cc_902 N_A_840_119#_c_1193_n N_A_367_491#_c_1926_n 0.00166658f $X=6.645 $Y=1.09
+ $X2=0 $Y2=0
cc_903 N_A_840_119#_c_1202_n N_A_367_491#_c_1936_n 0.00822086f $X=5.535 $Y=3.075
+ $X2=0 $Y2=0
cc_904 N_A_840_119#_c_1204_n N_A_367_491#_c_1936_n 0.0048013f $X=6.51 $Y=3.15
+ $X2=0 $Y2=0
cc_905 N_A_840_119#_c_1197_n N_VGND_M1023_d 0.00418757f $X=4.825 $Y=0.945 $X2=0
+ $Y2=0
cc_906 N_A_840_119#_M1013_g N_VGND_c_2098_n 0.00270145f $X=5.105 $Y=0.805 $X2=0
+ $Y2=0
cc_907 N_A_840_119#_c_1192_n N_VGND_c_2098_n 2.95613e-19 $X=5.61 $Y=1.165 $X2=0
+ $Y2=0
cc_908 N_A_840_119#_c_1197_n N_VGND_c_2098_n 0.0240111f $X=4.825 $Y=0.945 $X2=0
+ $Y2=0
cc_909 N_A_840_119#_c_1190_n N_VGND_c_2099_n 0.00377681f $X=5.535 $Y=1.09 $X2=0
+ $Y2=0
cc_910 N_A_840_119#_c_1191_n N_VGND_c_2099_n 0.0028073f $X=6.57 $Y=1.165 $X2=0
+ $Y2=0
cc_911 N_A_840_119#_M1024_g N_VGND_c_2101_n 0.00100535f $X=9.725 $Y=0.55 $X2=0
+ $Y2=0
cc_912 N_A_840_119#_c_1200_n N_VGND_c_2104_n 0.00285367f $X=4.34 $Y=0.865 $X2=0
+ $Y2=0
cc_913 N_A_840_119#_M1024_g N_VGND_c_2114_n 0.00305546f $X=9.725 $Y=0.55 $X2=0
+ $Y2=0
cc_914 N_A_840_119#_M1013_g N_VGND_c_2117_n 9.39239e-19 $X=5.105 $Y=0.805 $X2=0
+ $Y2=0
cc_915 N_A_840_119#_c_1190_n N_VGND_c_2117_n 9.39239e-19 $X=5.535 $Y=1.09 $X2=0
+ $Y2=0
cc_916 N_A_840_119#_M1024_g N_VGND_c_2117_n 0.00414861f $X=9.725 $Y=0.55 $X2=0
+ $Y2=0
cc_917 N_A_840_119#_c_1197_n N_VGND_c_2117_n 0.00782023f $X=4.825 $Y=0.945 $X2=0
+ $Y2=0
cc_918 N_A_840_119#_c_1200_n N_VGND_c_2117_n 0.0041548f $X=4.34 $Y=0.865 $X2=0
+ $Y2=0
cc_919 N_A_2002_42#_c_1367_n N_A_1812_379#_c_1478_n 0.00161746f $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_920 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1478_n 0.00773714f $X=11.19
+ $Y=0.615 $X2=0 $Y2=0
cc_921 N_A_2002_42#_c_1372_n N_A_1812_379#_M1025_g 0.00424803f $X=10.962
+ $Y=2.542 $X2=0 $Y2=0
cc_922 N_A_2002_42#_c_1392_n N_A_1812_379#_M1025_g 0.00596055f $X=10.935
+ $Y=2.755 $X2=0 $Y2=0
cc_923 N_A_2002_42#_c_1373_n N_A_1812_379#_M1025_g 0.00986239f $X=11.36 $Y=1.77
+ $X2=0 $Y2=0
cc_924 N_A_2002_42#_c_1374_n N_A_1812_379#_M1025_g 0.00325489f $X=11.135 $Y=1.77
+ $X2=0 $Y2=0
cc_925 N_A_2002_42#_c_1367_n N_A_1812_379#_M1025_g 0.00435137f $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_926 N_A_2002_42#_c_1376_n N_A_1812_379#_M1025_g 0.0108963f $X=10.962 $Y=2.37
+ $X2=0 $Y2=0
cc_927 N_A_2002_42#_c_1373_n N_A_1812_379#_c_1480_n 0.00268461f $X=11.36 $Y=1.77
+ $X2=0 $Y2=0
cc_928 N_A_2002_42#_c_1367_n N_A_1812_379#_c_1480_n 0.0120394f $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_929 N_A_2002_42#_c_1367_n N_A_1812_379#_c_1481_n 0.00534197f $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_930 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1481_n 0.00219113f $X=11.19
+ $Y=0.615 $X2=0 $Y2=0
cc_931 N_A_2002_42#_c_1367_n N_A_1812_379#_M1035_g 0.00471601f $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_932 N_A_2002_42#_c_1376_n N_A_1812_379#_M1035_g 4.97487e-19 $X=10.962 $Y=2.37
+ $X2=0 $Y2=0
cc_933 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1483_n 0.00437605f $X=11.19
+ $Y=0.615 $X2=0 $Y2=0
cc_934 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1485_n 0.011022f $X=11.19 $Y=0.615
+ $X2=0 $Y2=0
cc_935 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1486_n 0.00310261f $X=11.19
+ $Y=0.615 $X2=0 $Y2=0
cc_936 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1487_n 0.00655754f $X=11.19
+ $Y=0.615 $X2=0 $Y2=0
cc_937 N_A_2002_42#_c_1367_n N_A_1812_379#_c_1488_n 0.00312905f $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_938 N_A_2002_42#_M1032_g N_A_1812_379#_c_1504_n 0.00558743f $X=10.245 $Y=2.69
+ $X2=0 $Y2=0
cc_939 N_A_2002_42#_M1019_g N_A_1812_379#_c_1489_n 0.0010935f $X=10.085 $Y=0.55
+ $X2=0 $Y2=0
cc_940 N_A_2002_42#_M1032_g N_A_1812_379#_c_1489_n 0.00193135f $X=10.245 $Y=2.69
+ $X2=0 $Y2=0
cc_941 N_A_2002_42#_c_1368_n N_A_1812_379#_c_1489_n 0.0288416f $X=10.17 $Y=1.08
+ $X2=0 $Y2=0
cc_942 N_A_2002_42#_c_1369_n N_A_1812_379#_c_1489_n 0.00155827f $X=10.175
+ $Y=1.25 $X2=0 $Y2=0
cc_943 N_A_2002_42#_M1032_g N_A_1812_379#_c_1505_n 0.0152759f $X=10.245 $Y=2.69
+ $X2=0 $Y2=0
cc_944 N_A_2002_42#_M1032_g N_A_1812_379#_c_1490_n 0.0102306f $X=10.245 $Y=2.69
+ $X2=0 $Y2=0
cc_945 N_A_2002_42#_c_1366_n N_A_1812_379#_c_1490_n 0.0077694f $X=10.635 $Y=1.08
+ $X2=0 $Y2=0
cc_946 N_A_2002_42#_c_1369_n N_A_1812_379#_c_1490_n 5.03006e-19 $X=10.175
+ $Y=1.25 $X2=0 $Y2=0
cc_947 N_A_2002_42#_c_1374_n N_A_1812_379#_c_1491_n 8.44452e-19 $X=11.135
+ $Y=1.77 $X2=0 $Y2=0
cc_948 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1491_n 0.0145576f $X=11.19 $Y=0.615
+ $X2=0 $Y2=0
cc_949 N_A_2002_42#_M1019_g N_A_1812_379#_c_1492_n 0.00649664f $X=10.085 $Y=0.55
+ $X2=0 $Y2=0
cc_950 N_A_2002_42#_M1032_g N_A_1812_379#_c_1493_n 0.00111826f $X=10.245 $Y=2.69
+ $X2=0 $Y2=0
cc_951 N_A_2002_42#_c_1368_n N_A_1812_379#_c_1493_n 0.0245256f $X=10.17 $Y=1.08
+ $X2=0 $Y2=0
cc_952 N_A_2002_42#_c_1369_n N_A_1812_379#_c_1493_n 0.00453595f $X=10.175
+ $Y=1.25 $X2=0 $Y2=0
cc_953 N_A_2002_42#_M1032_g N_A_1812_379#_c_1494_n 0.00210697f $X=10.245 $Y=2.69
+ $X2=0 $Y2=0
cc_954 N_A_2002_42#_c_1366_n N_A_1812_379#_c_1494_n 0.00879841f $X=10.635
+ $Y=1.08 $X2=0 $Y2=0
cc_955 N_A_2002_42#_c_1369_n N_A_1812_379#_c_1494_n 0.00142933f $X=10.175
+ $Y=1.25 $X2=0 $Y2=0
cc_956 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1494_n 0.00326387f $X=11.19
+ $Y=0.615 $X2=0 $Y2=0
cc_957 N_A_2002_42#_c_1373_n N_A_1812_379#_c_1495_n 0.00387821f $X=11.36 $Y=1.77
+ $X2=0 $Y2=0
cc_958 N_A_2002_42#_c_1374_n N_A_1812_379#_c_1495_n 0.0137234f $X=11.135 $Y=1.77
+ $X2=0 $Y2=0
cc_959 N_A_2002_42#_c_1367_n N_A_1812_379#_c_1495_n 0.0269578f $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_960 N_A_2002_42#_c_1368_n N_A_1812_379#_c_1495_n 0.00438017f $X=10.17 $Y=1.08
+ $X2=0 $Y2=0
cc_961 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1495_n 0.0186935f $X=11.19 $Y=0.615
+ $X2=0 $Y2=0
cc_962 N_A_2002_42#_c_1373_n N_A_1812_379#_c_1498_n 0.00125939f $X=11.36 $Y=1.77
+ $X2=0 $Y2=0
cc_963 N_A_2002_42#_c_1374_n N_A_1812_379#_c_1498_n 7.6518e-19 $X=11.135 $Y=1.77
+ $X2=0 $Y2=0
cc_964 N_A_2002_42#_c_1367_n N_A_1812_379#_c_1498_n 0.00150664f $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_965 N_A_2002_42#_c_1370_n N_A_1812_379#_c_1498_n 0.00539052f $X=11.19
+ $Y=0.615 $X2=0 $Y2=0
cc_966 N_A_2002_42#_c_1367_n N_A_2352_327#_c_1696_n 0.023053f $X=11.475 $Y=1.685
+ $X2=0 $Y2=0
cc_967 N_A_2002_42#_c_1370_n N_A_2352_327#_c_1696_n 0.0099481f $X=11.19 $Y=0.615
+ $X2=0 $Y2=0
cc_968 N_A_2002_42#_c_1367_n N_A_2352_327#_c_1697_n 4.34377e-19 $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_969 N_A_2002_42#_c_1367_n N_A_2352_327#_c_1698_n 0.00134837f $X=11.475
+ $Y=1.685 $X2=0 $Y2=0
cc_970 N_A_2002_42#_c_1373_n N_VPWR_M1035_s 0.00506527f $X=11.36 $Y=1.77 $X2=0
+ $Y2=0
cc_971 N_A_2002_42#_c_1367_n N_VPWR_M1035_s 9.78397e-19 $X=11.475 $Y=1.685 $X2=0
+ $Y2=0
cc_972 N_A_2002_42#_M1032_g N_VPWR_c_1749_n 0.00320586f $X=10.245 $Y=2.69 $X2=0
+ $Y2=0
cc_973 N_A_2002_42#_c_1373_n N_VPWR_c_1750_n 0.021713f $X=11.36 $Y=1.77 $X2=0
+ $Y2=0
cc_974 N_A_2002_42#_c_1376_n N_VPWR_c_1750_n 0.0686967f $X=10.962 $Y=2.37 $X2=0
+ $Y2=0
cc_975 N_A_2002_42#_M1032_g N_VPWR_c_1758_n 0.00534427f $X=10.245 $Y=2.69 $X2=0
+ $Y2=0
cc_976 N_A_2002_42#_c_1392_n N_VPWR_c_1760_n 0.00990475f $X=10.935 $Y=2.755
+ $X2=0 $Y2=0
cc_977 N_A_2002_42#_M1032_g N_VPWR_c_1743_n 0.00526787f $X=10.245 $Y=2.69 $X2=0
+ $Y2=0
cc_978 N_A_2002_42#_c_1392_n N_VPWR_c_1743_n 0.0118144f $X=10.935 $Y=2.755 $X2=0
+ $Y2=0
cc_979 N_A_2002_42#_M1019_g N_VGND_c_2101_n 0.00848513f $X=10.085 $Y=0.55 $X2=0
+ $Y2=0
cc_980 N_A_2002_42#_c_1366_n N_VGND_c_2101_n 0.00571153f $X=10.635 $Y=1.08 $X2=0
+ $Y2=0
cc_981 N_A_2002_42#_c_1368_n N_VGND_c_2101_n 0.00827931f $X=10.17 $Y=1.08 $X2=0
+ $Y2=0
cc_982 N_A_2002_42#_c_1369_n N_VGND_c_2101_n 8.62589e-19 $X=10.175 $Y=1.25 $X2=0
+ $Y2=0
cc_983 N_A_2002_42#_c_1370_n N_VGND_c_2101_n 0.00305228f $X=11.19 $Y=0.615 $X2=0
+ $Y2=0
cc_984 N_A_2002_42#_c_1370_n N_VGND_c_2102_n 0.00742183f $X=11.19 $Y=0.615 $X2=0
+ $Y2=0
cc_985 N_A_2002_42#_M1019_g N_VGND_c_2114_n 0.0040395f $X=10.085 $Y=0.55 $X2=0
+ $Y2=0
cc_986 N_A_2002_42#_c_1370_n N_VGND_c_2115_n 0.0158229f $X=11.19 $Y=0.615 $X2=0
+ $Y2=0
cc_987 N_A_2002_42#_M1019_g N_VGND_c_2117_n 0.00773564f $X=10.085 $Y=0.55 $X2=0
+ $Y2=0
cc_988 N_A_2002_42#_c_1370_n N_VGND_c_2117_n 0.0261483f $X=11.19 $Y=0.615 $X2=0
+ $Y2=0
cc_989 N_A_2002_42#_c_1370_n A_2138_68# 0.00191422f $X=11.19 $Y=0.615 $X2=-0.19
+ $Y2=-0.245
cc_990 N_A_1812_379#_M1016_g N_A_2352_327#_M1039_g 0.0494897f $X=13.28 $Y=2.465
+ $X2=0 $Y2=0
cc_991 N_A_1812_379#_c_1507_n N_A_2352_327#_M1039_g 0.0159132f $X=13.04 $Y=2.54
+ $X2=0 $Y2=0
cc_992 N_A_1812_379#_c_1508_n N_A_2352_327#_M1039_g 0.00803727f $X=13.135
+ $Y=2.455 $X2=0 $Y2=0
cc_993 N_A_1812_379#_c_1511_n N_A_2352_327#_M1039_g 0.00198581f $X=12.135 $Y=2.6
+ $X2=0 $Y2=0
cc_994 N_A_1812_379#_c_1512_n N_A_2352_327#_M1039_g 0.0193448f $X=12.135 $Y=2.6
+ $X2=0 $Y2=0
cc_995 N_A_1812_379#_c_1496_n N_A_2352_327#_M1039_g 0.00138323f $X=13.33 $Y=1.51
+ $X2=0 $Y2=0
cc_996 N_A_1812_379#_c_1497_n N_A_2352_327#_M1039_g 0.00988188f $X=13.33 $Y=1.51
+ $X2=0 $Y2=0
cc_997 N_A_1812_379#_M1034_g N_A_2352_327#_c_1694_n 0.0147918f $X=13.31 $Y=0.795
+ $X2=0 $Y2=0
cc_998 N_A_1812_379#_c_1496_n N_A_2352_327#_c_1695_n 0.0010747f $X=13.33 $Y=1.51
+ $X2=0 $Y2=0
cc_999 N_A_1812_379#_c_1497_n N_A_2352_327#_c_1695_n 0.00853212f $X=13.33
+ $Y=1.51 $X2=0 $Y2=0
cc_1000 N_A_1812_379#_c_1481_n N_A_2352_327#_c_1696_n 0.0046899f $X=11.662
+ $Y=1.145 $X2=0 $Y2=0
cc_1001 N_A_1812_379#_M1035_g N_A_2352_327#_c_1696_n 0.00274066f $X=11.685
+ $Y=1.955 $X2=0 $Y2=0
cc_1002 N_A_1812_379#_c_1483_n N_A_2352_327#_c_1696_n 0.00901422f $X=11.925
+ $Y=0.765 $X2=0 $Y2=0
cc_1003 N_A_1812_379#_c_1488_n N_A_2352_327#_c_1696_n 0.00122237f $X=11.662
+ $Y=1.22 $X2=0 $Y2=0
cc_1004 N_A_1812_379#_c_1487_n N_A_2352_327#_c_1697_n 3.50304e-19 $X=11.925
+ $Y=0.84 $X2=0 $Y2=0
cc_1005 N_A_1812_379#_c_1488_n N_A_2352_327#_c_1697_n 0.0188202f $X=11.662
+ $Y=1.22 $X2=0 $Y2=0
cc_1006 N_A_1812_379#_M1035_g N_A_2352_327#_c_1698_n 6.99232e-19 $X=11.685
+ $Y=1.955 $X2=0 $Y2=0
cc_1007 N_A_1812_379#_c_1487_n N_A_2352_327#_c_1698_n 0.00508415f $X=11.925
+ $Y=0.84 $X2=0 $Y2=0
cc_1008 N_A_1812_379#_c_1511_n N_A_2352_327#_c_1698_n 0.0292186f $X=12.135
+ $Y=2.6 $X2=0 $Y2=0
cc_1009 N_A_1812_379#_c_1512_n N_A_2352_327#_c_1698_n 0.00919545f $X=12.135
+ $Y=2.6 $X2=0 $Y2=0
cc_1010 N_A_1812_379#_c_1507_n N_VPWR_M1039_d 0.00391543f $X=13.04 $Y=2.54 $X2=0
+ $Y2=0
cc_1011 N_A_1812_379#_c_1508_n N_VPWR_M1039_d 0.00603397f $X=13.135 $Y=2.455
+ $X2=0 $Y2=0
cc_1012 N_A_1812_379#_M1025_g N_VPWR_c_1749_n 0.00265776f $X=11.15 $Y=2.755
+ $X2=0 $Y2=0
cc_1013 N_A_1812_379#_c_1504_n N_VPWR_c_1749_n 0.0119002f $X=9.89 $Y=2.707 $X2=0
+ $Y2=0
cc_1014 N_A_1812_379#_M1025_g N_VPWR_c_1750_n 0.0139606f $X=11.15 $Y=2.755 $X2=0
+ $Y2=0
cc_1015 N_A_1812_379#_c_1500_n N_VPWR_c_1750_n 0.0250557f $X=11.97 $Y=3.15 $X2=0
+ $Y2=0
cc_1016 N_A_1812_379#_M1035_g N_VPWR_c_1750_n 0.011313f $X=11.685 $Y=1.955 $X2=0
+ $Y2=0
cc_1017 N_A_1812_379#_c_1511_n N_VPWR_c_1750_n 0.0300503f $X=12.135 $Y=2.6 $X2=0
+ $Y2=0
cc_1018 N_A_1812_379#_c_1512_n N_VPWR_c_1750_n 0.0109717f $X=12.135 $Y=2.6 $X2=0
+ $Y2=0
cc_1019 N_A_1812_379#_M1016_g N_VPWR_c_1751_n 0.00870422f $X=13.28 $Y=2.465
+ $X2=0 $Y2=0
cc_1020 N_A_1812_379#_c_1507_n N_VPWR_c_1751_n 0.0173237f $X=13.04 $Y=2.54 $X2=0
+ $Y2=0
cc_1021 N_A_1812_379#_c_1511_n N_VPWR_c_1751_n 0.00738921f $X=12.135 $Y=2.6
+ $X2=0 $Y2=0
cc_1022 N_A_1812_379#_c_1512_n N_VPWR_c_1751_n 0.00191217f $X=12.135 $Y=2.6
+ $X2=0 $Y2=0
cc_1023 N_A_1812_379#_c_1504_n N_VPWR_c_1758_n 0.0299387f $X=9.89 $Y=2.707 $X2=0
+ $Y2=0
cc_1024 N_A_1812_379#_c_1501_n N_VPWR_c_1760_n 0.00816041f $X=11.225 $Y=3.15
+ $X2=0 $Y2=0
cc_1025 N_A_1812_379#_c_1500_n N_VPWR_c_1762_n 0.0200205f $X=11.97 $Y=3.15 $X2=0
+ $Y2=0
cc_1026 N_A_1812_379#_c_1507_n N_VPWR_c_1762_n 0.00864277f $X=13.04 $Y=2.54
+ $X2=0 $Y2=0
cc_1027 N_A_1812_379#_c_1511_n N_VPWR_c_1762_n 0.0222109f $X=12.135 $Y=2.6 $X2=0
+ $Y2=0
cc_1028 N_A_1812_379#_M1016_g N_VPWR_c_1766_n 0.00486043f $X=13.28 $Y=2.465
+ $X2=0 $Y2=0
cc_1029 N_A_1812_379#_c_1500_n N_VPWR_c_1743_n 0.0328256f $X=11.97 $Y=3.15 $X2=0
+ $Y2=0
cc_1030 N_A_1812_379#_c_1501_n N_VPWR_c_1743_n 0.00931549f $X=11.225 $Y=3.15
+ $X2=0 $Y2=0
cc_1031 N_A_1812_379#_M1016_g N_VPWR_c_1743_n 0.00930295f $X=13.28 $Y=2.465
+ $X2=0 $Y2=0
cc_1032 N_A_1812_379#_c_1504_n N_VPWR_c_1743_n 0.0303562f $X=9.89 $Y=2.707 $X2=0
+ $Y2=0
cc_1033 N_A_1812_379#_c_1507_n N_VPWR_c_1743_n 0.0170176f $X=13.04 $Y=2.54 $X2=0
+ $Y2=0
cc_1034 N_A_1812_379#_c_1511_n N_VPWR_c_1743_n 0.0112205f $X=12.135 $Y=2.6 $X2=0
+ $Y2=0
cc_1035 N_A_1812_379#_c_1504_n A_1953_496# 0.00825055f $X=9.89 $Y=2.707
+ $X2=-0.19 $Y2=-0.245
cc_1036 N_A_1812_379#_c_1505_n A_1953_496# 4.0332e-19 $X=9.975 $Y=2.495
+ $X2=-0.19 $Y2=-0.245
cc_1037 N_A_1812_379#_c_1507_n N_Q_M1039_s 0.00691017f $X=13.04 $Y=2.54 $X2=0
+ $Y2=0
cc_1038 N_A_1812_379#_M1016_g Q 5.23259e-19 $X=13.28 $Y=2.465 $X2=0 $Y2=0
cc_1039 N_A_1812_379#_M1034_g Q 9.70295e-19 $X=13.31 $Y=0.795 $X2=0 $Y2=0
cc_1040 N_A_1812_379#_c_1507_n Q 0.0231038f $X=13.04 $Y=2.54 $X2=0 $Y2=0
cc_1041 N_A_1812_379#_c_1508_n Q 0.0375943f $X=13.135 $Y=2.455 $X2=0 $Y2=0
cc_1042 N_A_1812_379#_c_1496_n Q 0.0217474f $X=13.33 $Y=1.51 $X2=0 $Y2=0
cc_1043 N_A_1812_379#_c_1497_n Q 2.813e-19 $X=13.33 $Y=1.51 $X2=0 $Y2=0
cc_1044 N_A_1812_379#_c_1497_n Q_N 0.00253611f $X=13.33 $Y=1.51 $X2=0 $Y2=0
cc_1045 N_A_1812_379#_M1016_g Q_N 0.00254244f $X=13.28 $Y=2.465 $X2=0 $Y2=0
cc_1046 N_A_1812_379#_M1034_g Q_N 0.00398808f $X=13.31 $Y=0.795 $X2=0 $Y2=0
cc_1047 N_A_1812_379#_c_1508_n Q_N 0.00542448f $X=13.135 $Y=2.455 $X2=0 $Y2=0
cc_1048 N_A_1812_379#_c_1496_n Q_N 0.0251217f $X=13.33 $Y=1.51 $X2=0 $Y2=0
cc_1049 N_A_1812_379#_c_1497_n Q_N 0.00817336f $X=13.33 $Y=1.51 $X2=0 $Y2=0
cc_1050 N_A_1812_379#_c_1496_n Q_N 6.33027e-19 $X=13.33 $Y=1.51 $X2=0 $Y2=0
cc_1051 N_A_1812_379#_c_1497_n Q_N 0.0026802f $X=13.33 $Y=1.51 $X2=0 $Y2=0
cc_1052 N_A_1812_379#_M1034_g N_Q_N_c_2078_n 0.00248525f $X=13.31 $Y=0.795 $X2=0
+ $Y2=0
cc_1053 N_A_1812_379#_c_1492_n N_VGND_c_2101_n 0.0068398f $X=9.51 $Y=0.535 $X2=0
+ $Y2=0
cc_1054 N_A_1812_379#_c_1483_n N_VGND_c_2102_n 0.0118122f $X=11.925 $Y=0.765
+ $X2=0 $Y2=0
cc_1055 N_A_1812_379#_c_1485_n N_VGND_c_2102_n 0.00646705f $X=10.98 $Y=0.835
+ $X2=0 $Y2=0
cc_1056 N_A_1812_379#_c_1487_n N_VGND_c_2102_n 0.01012f $X=11.925 $Y=0.84 $X2=0
+ $Y2=0
cc_1057 N_A_1812_379#_M1034_g N_VGND_c_2103_n 0.00366731f $X=13.31 $Y=0.795
+ $X2=0 $Y2=0
cc_1058 N_A_1812_379#_c_1496_n N_VGND_c_2103_n 0.0136441f $X=13.33 $Y=1.51 $X2=0
+ $Y2=0
cc_1059 N_A_1812_379#_c_1497_n N_VGND_c_2103_n 0.00130922f $X=13.33 $Y=1.51
+ $X2=0 $Y2=0
cc_1060 N_A_1812_379#_c_1483_n N_VGND_c_2110_n 0.00486043f $X=11.925 $Y=0.765
+ $X2=0 $Y2=0
cc_1061 N_A_1812_379#_c_1492_n N_VGND_c_2114_n 0.0190328f $X=9.51 $Y=0.535 $X2=0
+ $Y2=0
cc_1062 N_A_1812_379#_c_1485_n N_VGND_c_2115_n 0.00351444f $X=10.98 $Y=0.835
+ $X2=0 $Y2=0
cc_1063 N_A_1812_379#_M1034_g N_VGND_c_2116_n 0.00457417f $X=13.31 $Y=0.795
+ $X2=0 $Y2=0
cc_1064 N_A_1812_379#_c_1483_n N_VGND_c_2117_n 0.00975473f $X=11.925 $Y=0.765
+ $X2=0 $Y2=0
cc_1065 N_A_1812_379#_M1034_g N_VGND_c_2117_n 0.00544287f $X=13.31 $Y=0.795
+ $X2=0 $Y2=0
cc_1066 N_A_1812_379#_c_1485_n N_VGND_c_2117_n 0.00512192f $X=10.98 $Y=0.835
+ $X2=0 $Y2=0
cc_1067 N_A_1812_379#_c_1492_n N_VGND_c_2117_n 0.0143264f $X=9.51 $Y=0.535 $X2=0
+ $Y2=0
cc_1068 N_A_2352_327#_c_1698_n N_VPWR_c_1750_n 0.0101545f $X=11.9 $Y=1.78 $X2=0
+ $Y2=0
cc_1069 N_A_2352_327#_M1039_g N_VPWR_c_1751_n 0.0109651f $X=12.85 $Y=2.465 $X2=0
+ $Y2=0
cc_1070 N_A_2352_327#_M1039_g N_VPWR_c_1762_n 0.00361815f $X=12.85 $Y=2.465
+ $X2=0 $Y2=0
cc_1071 N_A_2352_327#_M1039_g N_VPWR_c_1743_n 0.00479281f $X=12.85 $Y=2.465
+ $X2=0 $Y2=0
cc_1072 N_A_2352_327#_c_1692_n Q 0.0206843f $X=12.775 $Y=1.4 $X2=0 $Y2=0
cc_1073 N_A_2352_327#_M1039_g Q 0.0198674f $X=12.85 $Y=2.465 $X2=0 $Y2=0
cc_1074 N_A_2352_327#_c_1694_n Q 0.0157777f $X=12.88 $Y=1.325 $X2=0 $Y2=0
cc_1075 N_A_2352_327#_c_1695_n Q 0.00288526f $X=12.865 $Y=1.4 $X2=0 $Y2=0
cc_1076 N_A_2352_327#_c_1696_n Q 0.159221f $X=12.14 $Y=0.445 $X2=0 $Y2=0
cc_1077 N_A_2352_327#_c_1697_n Q 0.00167269f $X=12.16 $Y=1.31 $X2=0 $Y2=0
cc_1078 N_A_2352_327#_c_1694_n N_VGND_c_2103_n 0.00353791f $X=12.88 $Y=1.325
+ $X2=0 $Y2=0
cc_1079 N_A_2352_327#_c_1694_n N_VGND_c_2110_n 0.0044174f $X=12.88 $Y=1.325
+ $X2=0 $Y2=0
cc_1080 N_A_2352_327#_c_1696_n N_VGND_c_2110_n 0.0153489f $X=12.14 $Y=0.445
+ $X2=0 $Y2=0
cc_1081 N_A_2352_327#_M1036_d N_VGND_c_2117_n 0.00376753f $X=12 $Y=0.235 $X2=0
+ $Y2=0
cc_1082 N_A_2352_327#_c_1694_n N_VGND_c_2117_n 0.00544287f $X=12.88 $Y=1.325
+ $X2=0 $Y2=0
cc_1083 N_A_2352_327#_c_1696_n N_VGND_c_2117_n 0.00990863f $X=12.14 $Y=0.445
+ $X2=0 $Y2=0
cc_1084 N_VPWR_c_1743_n A_295_491# 0.00899413f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1085 N_VPWR_c_1743_n N_A_367_491#_M1028_d 0.00223559f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1086 N_VPWR_c_1743_n N_A_367_491#_M1040_d 0.00215158f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1087 N_VPWR_M1017_d N_A_367_491#_c_1928_n 0.00259179f $X=2.76 $Y=2.455 $X2=0
+ $Y2=0
cc_1088 N_VPWR_c_1745_n N_A_367_491#_c_1928_n 0.0177127f $X=2.94 $Y=2.895 $X2=0
+ $Y2=0
cc_1089 N_VPWR_c_1752_n N_A_367_491#_c_1928_n 0.00842033f $X=2.775 $Y=3.33 $X2=0
+ $Y2=0
cc_1090 N_VPWR_c_1743_n N_A_367_491#_c_1928_n 0.0169822f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1091 N_VPWR_M1001_d N_A_367_491#_c_1930_n 0.00363026f $X=4.69 $Y=1.835 $X2=0
+ $Y2=0
cc_1092 N_VPWR_c_1746_n N_A_367_491#_c_1930_n 0.0163525f $X=4.83 $Y=2.895 $X2=0
+ $Y2=0
cc_1093 N_VPWR_c_1754_n N_A_367_491#_c_1930_n 0.0157544f $X=4.665 $Y=3.33 $X2=0
+ $Y2=0
cc_1094 N_VPWR_c_1756_n N_A_367_491#_c_1930_n 0.0110698f $X=7.075 $Y=3.33 $X2=0
+ $Y2=0
cc_1095 N_VPWR_c_1743_n N_A_367_491#_c_1930_n 0.0482728f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1096 N_VPWR_M1017_d N_A_367_491#_c_1931_n 5.70704e-19 $X=2.76 $Y=2.455 $X2=0
+ $Y2=0
cc_1097 N_VPWR_c_1745_n N_A_367_491#_c_1931_n 0.00456214f $X=2.94 $Y=2.895 $X2=0
+ $Y2=0
cc_1098 N_VPWR_c_1754_n N_A_367_491#_c_1931_n 0.00217767f $X=4.665 $Y=3.33 $X2=0
+ $Y2=0
cc_1099 N_VPWR_c_1743_n N_A_367_491#_c_1931_n 0.00443319f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1100 N_VPWR_c_1744_n N_A_367_491#_c_1934_n 0.0213871f $X=1.185 $Y=2.6 $X2=0
+ $Y2=0
cc_1101 N_VPWR_c_1752_n N_A_367_491#_c_1934_n 0.0189395f $X=2.775 $Y=3.33 $X2=0
+ $Y2=0
cc_1102 N_VPWR_c_1743_n N_A_367_491#_c_1934_n 0.0123908f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1103 N_VPWR_c_1754_n N_A_367_491#_c_1935_n 0.0209292f $X=4.665 $Y=3.33 $X2=0
+ $Y2=0
cc_1104 N_VPWR_c_1743_n N_A_367_491#_c_1935_n 0.0125409f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1105 N_VPWR_c_1756_n N_A_367_491#_c_1936_n 0.00467875f $X=7.075 $Y=3.33 $X2=0
+ $Y2=0
cc_1106 N_VPWR_c_1743_n N_A_367_491#_c_1936_n 0.00666895f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_1107 N_VPWR_c_1743_n A_453_491# 0.00439141f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1108 N_VPWR_c_1743_n N_Q_M1039_s 0.003382f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1109 N_VPWR_c_1743_n N_Q_N_M1016_d 0.00371702f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1110 N_VPWR_c_1766_n Q_N 0.0253382f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1111 N_VPWR_c_1743_n Q_N 0.0141126f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1112 N_A_367_491#_c_1928_n A_453_491# 0.00441364f $X=3.04 $Y=2.502 $X2=-0.19
+ $Y2=-0.245
cc_1113 N_A_367_491#_c_1924_n N_VGND_c_2117_n 0.00560423f $X=3.04 $Y=0.9 $X2=0
+ $Y2=0
cc_1114 N_A_367_491#_c_1924_n N_noxref_25_M1030_d 0.00248206f $X=3.04 $Y=0.9
+ $X2=0 $Y2=0
cc_1115 N_A_367_491#_M1011_d N_noxref_25_c_2237_n 0.00176461f $X=2.01 $Y=0.405
+ $X2=0 $Y2=0
cc_1116 N_A_367_491#_c_1924_n N_noxref_25_c_2237_n 0.0107288f $X=3.04 $Y=0.9
+ $X2=0 $Y2=0
cc_1117 N_A_367_491#_c_1927_n N_noxref_25_c_2237_n 0.0153209f $X=2.15 $Y=0.7
+ $X2=0 $Y2=0
cc_1118 N_A_367_491#_c_1924_n N_noxref_25_c_2239_n 0.0199717f $X=3.04 $Y=0.9
+ $X2=0 $Y2=0
cc_1119 N_A_367_491#_c_1927_n N_noxref_25_c_2239_n 0.00167287f $X=2.15 $Y=0.7
+ $X2=0 $Y2=0
cc_1120 N_A_367_491#_c_1924_n noxref_27 0.00147531f $X=3.04 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_1121 Q N_VGND_c_2103_n 0.0317293f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_1122 Q N_VGND_c_2110_n 0.0149624f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_1123 Q N_VGND_c_2117_n 0.0125623f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_1124 N_Q_N_c_2078_n N_VGND_c_2103_n 0.00155513f $X=13.525 $Y=0.52 $X2=0 $Y2=0
cc_1125 N_Q_N_c_2078_n N_VGND_c_2116_n 0.0160975f $X=13.525 $Y=0.52 $X2=0 $Y2=0
cc_1126 N_Q_N_c_2078_n N_VGND_c_2117_n 0.0135505f $X=13.525 $Y=0.52 $X2=0 $Y2=0
cc_1127 N_VGND_c_2096_n N_noxref_25_c_2236_n 0.015285f $X=0.69 $Y=0.52 $X2=0
+ $Y2=0
cc_1128 N_VGND_c_2113_n N_noxref_25_c_2237_n 0.0942291f $X=3.275 $Y=0 $X2=0
+ $Y2=0
cc_1129 N_VGND_c_2117_n N_noxref_25_c_2237_n 0.0545822f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1130 N_VGND_c_2096_n N_noxref_25_c_2238_n 0.0110442f $X=0.69 $Y=0.52 $X2=0
+ $Y2=0
cc_1131 N_VGND_c_2113_n N_noxref_25_c_2238_n 0.018162f $X=3.275 $Y=0 $X2=0 $Y2=0
cc_1132 N_VGND_c_2117_n N_noxref_25_c_2238_n 0.0100189f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1133 N_VGND_c_2097_n N_noxref_25_c_2239_n 0.0207954f $X=3.44 $Y=0.56 $X2=0
+ $Y2=0
cc_1134 N_VGND_c_2113_n N_noxref_25_c_2239_n 0.022561f $X=3.275 $Y=0 $X2=0 $Y2=0
cc_1135 N_VGND_c_2117_n N_noxref_25_c_2239_n 0.0125743f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_1136 N_noxref_25_c_2237_n noxref_26 0.00354478f $X=2.775 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1137 N_noxref_25_c_2237_n noxref_27 0.00151984f $X=2.775 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
