* File: sky130_fd_sc_lp__a211oi_1.spice
* Created: Wed Sep  2 09:18:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a211oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a211oi_1  VNB VPB A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1002 A_110_49# N_A2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1007 N_Y_M1007_d N_A1_M1007_g A_110_49# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=11.424 NRS=7.14 M=1 R=5.6 SA=75000.6 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_B1_M1001_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=13.56 NRS=4.284 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_C1_M1005_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=2.136 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_A2_M1006_g N_A_27_367#_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.3339 PD=1.65 PS=3.05 NRD=8.5892 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1000 N_A_27_367#_M1000_d N_A1_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=9.3772 NRS=8.5892 M=1 R=8.4 SA=75000.7
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 A_326_367# N_B1_M1003_g N_A_27_367#_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.2457 PD=1.47 PS=1.65 NRD=7.8012 NRS=7.8012 M=1 R=8.4 SA=75001.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_C1_M1004_g A_326_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.3339
+ AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.6 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__a211oi_1.pxi.spice"
*
.ends
*
*
