# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__srsdfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__srsdfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.24000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.180000 1.805000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.585900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.795000 0.265000 18.135000 3.075000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.598000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.605000 0.255000 7.070000 0.425000 ;
        RECT 6.900000 0.425000 7.070000 1.610000 ;
        RECT 6.900000 1.610000 8.140000 1.780000 ;
        RECT 7.805000 1.215000 8.140000 1.610000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.605000 2.870000 2.275000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 1.095000 0.915000 1.780000 ;
    END
  END SCE
  PIN SLEEP_B
    ANTENNAGATEAREA  0.598000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.195000 1.295000 11.560000 1.780000 ;
    END
  END SLEEP_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 10.205000 1.555000 10.685000 1.840000 ;
    END
  END CLK_N
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT  0.070000 2.675000 18.170000 2.945000 ;
        RECT  7.775000 2.660000  8.065000 2.675000 ;
        RECT  8.255000 2.660000  8.545000 2.675000 ;
        RECT 11.615000 2.660000 11.905000 2.675000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 18.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 18.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.240000 0.085000 ;
      RECT  0.000000  3.245000 18.240000 3.415000 ;
      RECT  0.105000  0.255000  0.355000 1.950000 ;
      RECT  0.105000  1.950000  2.305000 2.120000 ;
      RECT  0.105000  2.120000  0.610000 3.075000 ;
      RECT  0.535000  0.085000  0.865000 0.715000 ;
      RECT  0.780000  2.435000  1.110000 3.245000 ;
      RECT  1.070000  0.255000  3.080000 0.425000 ;
      RECT  1.070000  0.425000  1.320000 0.925000 ;
      RECT  1.500000  0.595000  2.145000 0.925000 ;
      RECT  1.600000  2.445000  3.260000 2.615000 ;
      RECT  1.600000  2.615000  1.930000 3.075000 ;
      RECT  1.975000  0.925000  2.145000 1.265000 ;
      RECT  1.975000  1.265000  3.210000 1.435000 ;
      RECT  1.975000  1.945000  2.305000 1.950000 ;
      RECT  1.975000  2.120000  2.305000 2.275000 ;
      RECT  2.400000  0.595000  2.570000 0.925000 ;
      RECT  2.400000  0.925000  4.700000 1.095000 ;
      RECT  2.670000  2.785000  2.920000 3.245000 ;
      RECT  2.750000  0.425000  3.080000 0.755000 ;
      RECT  3.040000  1.435000  3.210000 2.445000 ;
      RECT  3.090000  2.615000  3.260000 2.905000 ;
      RECT  3.090000  2.905000  4.115000 3.075000 ;
      RECT  3.380000  1.265000  3.735000 1.595000 ;
      RECT  3.485000  1.595000  3.735000 2.735000 ;
      RECT  3.835000  0.085000  4.165000 0.755000 ;
      RECT  3.945000  1.735000  4.805000 1.905000 ;
      RECT  3.945000  1.905000  4.115000 2.905000 ;
      RECT  4.285000  2.075000  4.455000 3.245000 ;
      RECT  4.370000  0.595000  4.700000 0.925000 ;
      RECT  4.635000  1.265000  5.380000 1.435000 ;
      RECT  4.635000  1.435000  4.805000 1.735000 ;
      RECT  4.635000  1.905000  4.805000 2.105000 ;
      RECT  4.635000  2.105000  4.965000 2.755000 ;
      RECT  5.015000  0.595000  6.730000 0.765000 ;
      RECT  5.050000  1.605000  5.380000 1.935000 ;
      RECT  5.210000  0.935000  6.670000 1.105000 ;
      RECT  5.210000  1.105000  5.380000 1.265000 ;
      RECT  5.210000  1.935000  5.380000 2.905000 ;
      RECT  5.210000  2.905000  7.245000 3.075000 ;
      RECT  5.550000  1.275000  5.985000 2.320000 ;
      RECT  5.550000  2.320000  6.905000 2.490000 ;
      RECT  5.550000  2.490000  5.985000 2.735000 ;
      RECT  6.155000  1.605000  6.565000 2.150000 ;
      RECT  6.340000  1.105000  6.670000 1.435000 ;
      RECT  6.735000  1.950000  8.185000 2.010000 ;
      RECT  6.735000  2.010000 10.335000 2.180000 ;
      RECT  6.735000  2.180000  6.905000 2.320000 ;
      RECT  7.075000  2.350000  9.580000 2.520000 ;
      RECT  7.075000  2.520000  7.245000 2.905000 ;
      RECT  7.240000  0.365000  7.570000 0.535000 ;
      RECT  7.240000  0.535000  8.645000 0.705000 ;
      RECT  7.240000  0.875000  9.865000 1.045000 ;
      RECT  7.240000  1.045000  7.570000 1.440000 ;
      RECT  7.415000  2.690000  8.035000 3.075000 ;
      RECT  7.780000  0.085000  8.110000 0.365000 ;
      RECT  8.285000  2.690000  9.240000 3.020000 ;
      RECT  8.315000  0.255000  8.645000 0.535000 ;
      RECT  8.355000  1.045000  8.525000 1.670000 ;
      RECT  8.355000  1.670000  9.960000 1.840000 ;
      RECT  8.695000  1.215000 10.205000 1.385000 ;
      RECT  8.695000  1.385000  9.025000 1.500000 ;
      RECT  8.825000  0.085000  9.075000 0.675000 ;
      RECT  9.410000  2.520000  9.580000 2.725000 ;
      RECT  9.410000  2.725000 10.675000 2.895000 ;
      RECT  9.535000  0.255000 11.705000 0.425000 ;
      RECT  9.535000  0.425000  9.865000 0.875000 ;
      RECT  9.630000  1.590000  9.960000 1.670000 ;
      RECT 10.035000  0.595000 11.365000 0.765000 ;
      RECT 10.035000  0.765000 10.205000 1.215000 ;
      RECT 10.080000  2.180000 10.335000 2.555000 ;
      RECT 10.420000  0.935000 11.025000 1.265000 ;
      RECT 10.505000  2.010000 12.080000 2.120000 ;
      RECT 10.505000  2.120000 11.445000 2.180000 ;
      RECT 10.505000  2.180000 10.675000 2.725000 ;
      RECT 10.845000  2.350000 11.015000 2.905000 ;
      RECT 10.845000  2.905000 12.050000 3.075000 ;
      RECT 10.855000  1.265000 11.025000 2.010000 ;
      RECT 11.195000  0.765000 11.365000 0.955000 ;
      RECT 11.195000  0.955000 13.485000 1.125000 ;
      RECT 11.195000  1.950000 12.080000 2.010000 ;
      RECT 11.195000  2.180000 11.445000 2.735000 ;
      RECT 11.535000  0.425000 11.705000 0.615000 ;
      RECT 11.535000  0.615000 12.595000 0.785000 ;
      RECT 11.645000  2.290000 12.050000 2.905000 ;
      RECT 11.910000  0.085000 12.160000 0.445000 ;
      RECT 11.910000  1.375000 13.145000 1.545000 ;
      RECT 11.910000  1.545000 12.080000 1.950000 ;
      RECT 12.250000  1.715000 12.580000 1.905000 ;
      RECT 12.250000  1.905000 13.485000 2.075000 ;
      RECT 12.250000  2.075000 12.580000 2.755000 ;
      RECT 12.425000  0.255000 14.700000 0.425000 ;
      RECT 12.425000  0.425000 12.595000 0.615000 ;
      RECT 12.750000  1.545000 13.145000 1.735000 ;
      RECT 12.765000  0.595000 13.095000 0.955000 ;
      RECT 12.770000  2.245000 13.100000 2.905000 ;
      RECT 12.770000  2.905000 15.265000 3.075000 ;
      RECT 13.315000  1.125000 13.485000 1.905000 ;
      RECT 13.325000  0.425000 13.655000 0.615000 ;
      RECT 13.655000  0.785000 14.155000 0.955000 ;
      RECT 13.655000  0.955000 13.905000 2.565000 ;
      RECT 13.655000  2.565000 14.925000 2.735000 ;
      RECT 13.825000  0.595000 14.155000 0.785000 ;
      RECT 14.075000  1.125000 14.360000 1.455000 ;
      RECT 14.075000  1.455000 14.245000 2.150000 ;
      RECT 14.415000  1.625000 14.700000 1.795000 ;
      RECT 14.415000  1.795000 14.585000 2.395000 ;
      RECT 14.530000  0.425000 14.700000 1.625000 ;
      RECT 14.755000  1.965000 15.040000 2.135000 ;
      RECT 14.755000  2.135000 14.925000 2.565000 ;
      RECT 14.870000  1.105000 15.790000 1.275000 ;
      RECT 14.870000  1.275000 15.040000 1.965000 ;
      RECT 15.095000  2.305000 15.265000 2.905000 ;
      RECT 15.120000  0.085000 15.450000 0.935000 ;
      RECT 15.210000  1.805000 16.205000 2.135000 ;
      RECT 15.445000  2.305000 15.695000 3.245000 ;
      RECT 15.620000  0.255000 16.650000 0.425000 ;
      RECT 15.620000  0.425000 15.790000 1.105000 ;
      RECT 15.875000  2.135000 16.205000 2.755000 ;
      RECT 16.035000  0.595000 16.305000 0.935000 ;
      RECT 16.035000  0.935000 16.205000 1.805000 ;
      RECT 16.385000  2.295000 16.635000 3.245000 ;
      RECT 16.480000  0.425000 16.650000 0.895000 ;
      RECT 16.480000  0.895000 16.810000 1.565000 ;
      RECT 16.820000  0.265000 17.150000 0.725000 ;
      RECT 16.840000  2.435000 17.170000 3.075000 ;
      RECT 16.980000  0.725000 17.150000 1.315000 ;
      RECT 16.980000  1.315000 17.625000 1.645000 ;
      RECT 16.980000  1.645000 17.170000 2.435000 ;
      RECT 17.365000  0.085000 17.615000 1.145000 ;
      RECT 17.375000  1.815000 17.625000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  1.950000  3.685000 2.120000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.950000  6.565000 2.120000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  2.690000  8.005000 2.860000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  2.690000  8.485000 2.860000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  2.690000 11.845000 2.860000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  1.950000 14.245000 2.120000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.245000 18.085000 3.415000 ;
    LAYER met1 ;
      RECT  3.455000 1.920000  3.745000 1.965000 ;
      RECT  3.455000 1.965000 14.305000 2.105000 ;
      RECT  3.455000 2.105000  3.745000 2.150000 ;
      RECT  6.335000 1.920000  6.625000 1.965000 ;
      RECT  6.335000 2.105000  6.625000 2.150000 ;
      RECT 14.015000 1.920000 14.305000 1.965000 ;
      RECT 14.015000 2.105000 14.305000 2.150000 ;
  END
END sky130_fd_sc_lp__srsdfrtn_1
END LIBRARY
