* File: sky130_fd_sc_lp__a22o_m.pxi.spice
* Created: Wed Sep  2 09:22:52 2020
* 
x_PM_SKY130_FD_SC_LP__A22O_M%A_85_317# N_A_85_317#_M1004_d N_A_85_317#_M1000_d
+ N_A_85_317#_M1002_g N_A_85_317#_M1001_g N_A_85_317#_c_66_n N_A_85_317#_c_72_n
+ N_A_85_317#_c_67_n N_A_85_317#_c_73_n N_A_85_317#_c_68_n N_A_85_317#_c_75_n
+ N_A_85_317#_c_69_n N_A_85_317#_c_76_n N_A_85_317#_c_93_p N_A_85_317#_c_77_n
+ PM_SKY130_FD_SC_LP__A22O_M%A_85_317#
x_PM_SKY130_FD_SC_LP__A22O_M%A2 N_A2_M1007_g N_A2_M1005_g A2 A2 N_A2_c_147_n
+ N_A2_c_148_n PM_SKY130_FD_SC_LP__A22O_M%A2
x_PM_SKY130_FD_SC_LP__A22O_M%A1 N_A1_M1004_g N_A1_M1003_g N_A1_c_191_n
+ N_A1_c_183_n N_A1_c_184_n A1 A1 A1 A1 N_A1_c_187_n N_A1_c_188_n N_A1_c_189_n
+ PM_SKY130_FD_SC_LP__A22O_M%A1
x_PM_SKY130_FD_SC_LP__A22O_M%B1 N_B1_M1000_g N_B1_c_242_n N_B1_M1009_g B1 B1
+ N_B1_c_244_n PM_SKY130_FD_SC_LP__A22O_M%B1
x_PM_SKY130_FD_SC_LP__A22O_M%B2 N_B2_c_282_n N_B2_M1006_g N_B2_M1008_g B2 B2 B2
+ N_B2_c_285_n PM_SKY130_FD_SC_LP__A22O_M%B2
x_PM_SKY130_FD_SC_LP__A22O_M%X N_X_M1001_s N_X_M1002_s N_X_c_325_n N_X_c_326_n X
+ X X X X N_X_c_329_n PM_SKY130_FD_SC_LP__A22O_M%X
x_PM_SKY130_FD_SC_LP__A22O_M%VPWR N_VPWR_M1002_d N_VPWR_M1003_d N_VPWR_c_348_n
+ N_VPWR_c_349_n N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n VPWR
+ N_VPWR_c_353_n N_VPWR_c_347_n PM_SKY130_FD_SC_LP__A22O_M%VPWR
x_PM_SKY130_FD_SC_LP__A22O_M%A_265_501# N_A_265_501#_M1005_d
+ N_A_265_501#_M1006_d N_A_265_501#_c_384_n N_A_265_501#_c_385_n
+ N_A_265_501#_c_386_n PM_SKY130_FD_SC_LP__A22O_M%A_265_501#
x_PM_SKY130_FD_SC_LP__A22O_M%VGND N_VGND_M1001_d N_VGND_M1008_d N_VGND_c_409_n
+ N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n
+ VGND N_VGND_c_415_n N_VGND_c_416_n PM_SKY130_FD_SC_LP__A22O_M%VGND
cc_1 VNB N_A_85_317#_M1001_g 0.0473901f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.835
cc_2 VNB N_A_85_317#_c_66_n 0.012021f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.735
cc_3 VNB N_A_85_317#_c_67_n 0.00352803f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.755
cc_4 VNB N_A_85_317#_c_68_n 0.0102964f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.67
cc_5 VNB N_A_85_317#_c_69_n 0.00484425f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.585
cc_6 VNB N_A2_M1005_g 0.00899688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB A2 0.0093938f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.715
cc_8 VNB N_A2_c_147_n 0.0325535f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.835
cc_9 VNB N_A2_c_148_n 0.0177931f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.735
cc_10 VNB N_A1_c_183_n 0.0255818f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.585
cc_11 VNB N_A1_c_184_n 0.0466824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A1 0.0293543f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.09
cc_13 VNB A1 0.0138756f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.255
cc_14 VNB N_A1_c_187_n 0.012711f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.67
cc_15 VNB N_A1_c_188_n 0.015532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_189_n 0.0081723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_M1000_g 0.00479172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_242_n 0.0167827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB B1 0.00893891f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.715
cc_20 VNB N_B1_c_244_n 0.0569578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B2_M1008_g 0.0485369f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.255
cc_22 VNB N_X_c_325_n 0.0127826f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.255
cc_23 VNB N_X_c_326_n 0.00143848f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.715
cc_24 VNB X 0.0324271f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.835
cc_25 VNB N_VPWR_c_347_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_409_n 0.0250375f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.715
cc_27 VNB N_VGND_c_410_n 0.0247208f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.835
cc_28 VNB N_VGND_c_411_n 0.0282373f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.585
cc_29 VNB N_VGND_c_412_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.735
cc_30 VNB N_VGND_c_413_n 0.0423326f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.255
cc_31 VNB N_VGND_c_414_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.755
cc_32 VNB N_VGND_c_415_n 0.0140765f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=0.81
cc_33 VNB N_VGND_c_416_n 0.237659f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=0.81
cc_34 VPB N_A_85_317#_M1002_g 0.0302376f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.715
cc_35 VPB N_A_85_317#_c_66_n 0.00717895f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.735
cc_36 VPB N_A_85_317#_c_72_n 0.01771f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.255
cc_37 VPB N_A_85_317#_c_73_n 0.0117645f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.04
cc_38 VPB N_A_85_317#_c_68_n 0.00703312f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=1.67
cc_39 VPB N_A_85_317#_c_75_n 0.0140606f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=2.41
cc_40 VPB N_A_85_317#_c_76_n 0.0269798f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.75
cc_41 VPB N_A_85_317#_c_77_n 0.00696766f $X=-0.19 $Y=1.655 $X2=2.01 $Y2=2.41
cc_42 VPB N_A2_M1005_g 0.0558835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A1_M1003_g 0.029703f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A1_c_191_n 0.0239163f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB A1 0.046397f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.255
cc_46 VPB N_A1_c_187_n 0.0367122f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.67
cc_47 VPB N_B1_M1000_g 0.0565567f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB B1 0.00360114f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.715
cc_49 VPB N_B2_c_282_n 0.064314f $X=-0.19 $Y=1.655 $X2=1.685 $Y2=0.625
cc_50 VPB N_B2_M1006_g 0.0333515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B2_M1008_g 0.00239931f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.255
cc_52 VPB N_B2_c_285_n 0.0155089f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.735
cc_53 VPB X 0.0417284f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.835
cc_54 VPB N_X_c_329_n 0.0166666f $X=-0.19 $Y=1.655 $X2=1.825 $Y2=0.81
cc_55 VPB N_VPWR_c_348_n 0.00867537f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.715
cc_56 VPB N_VPWR_c_349_n 0.014379f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.585
cc_57 VPB N_VPWR_c_350_n 0.0200055f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.835
cc_58 VPB N_VPWR_c_351_n 0.022934f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.585
cc_59 VPB N_VPWR_c_352_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.735
cc_60 VPB N_VPWR_c_353_n 0.0438678f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=2.41
cc_61 VPB N_VPWR_c_347_n 0.0701993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_265_501#_c_384_n 0.005626f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.255
cc_63 VPB N_A_265_501#_c_385_n 0.00253418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_265_501#_c_386_n 0.00252845f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.735
cc_65 N_A_85_317#_M1002_g N_A2_M1005_g 0.0136593f $X=0.66 $Y=2.715 $X2=0 $Y2=0
cc_66 N_A_85_317#_M1001_g N_A2_M1005_g 0.00805859f $X=0.71 $Y=0.835 $X2=0 $Y2=0
cc_67 N_A_85_317#_c_73_n N_A2_M1005_g 0.0100087f $X=0.72 $Y=2.04 $X2=0 $Y2=0
cc_68 N_A_85_317#_c_68_n N_A2_M1005_g 0.0111471f $X=1.625 $Y=1.67 $X2=0 $Y2=0
cc_69 N_A_85_317#_c_75_n N_A2_M1005_g 0.0123531f $X=1.845 $Y=2.41 $X2=0 $Y2=0
cc_70 N_A_85_317#_c_76_n N_A2_M1005_g 0.0125496f $X=0.59 $Y=1.75 $X2=0 $Y2=0
cc_71 N_A_85_317#_M1001_g A2 0.0137423f $X=0.71 $Y=0.835 $X2=0 $Y2=0
cc_72 N_A_85_317#_c_67_n A2 0.0232842f $X=0.72 $Y=1.755 $X2=0 $Y2=0
cc_73 N_A_85_317#_c_68_n A2 0.0266206f $X=1.625 $Y=1.67 $X2=0 $Y2=0
cc_74 N_A_85_317#_c_69_n A2 0.0100716f $X=1.71 $Y=1.585 $X2=0 $Y2=0
cc_75 N_A_85_317#_M1001_g N_A2_c_147_n 0.0217873f $X=0.71 $Y=0.835 $X2=0 $Y2=0
cc_76 N_A_85_317#_c_68_n N_A2_c_147_n 0.00440824f $X=1.625 $Y=1.67 $X2=0 $Y2=0
cc_77 N_A_85_317#_c_69_n N_A2_c_147_n 0.00280434f $X=1.71 $Y=1.585 $X2=0 $Y2=0
cc_78 N_A_85_317#_M1001_g N_A2_c_148_n 0.014051f $X=0.71 $Y=0.835 $X2=0 $Y2=0
cc_79 N_A_85_317#_c_69_n N_A2_c_148_n 0.00109697f $X=1.71 $Y=1.585 $X2=0 $Y2=0
cc_80 N_A_85_317#_c_93_p N_A2_c_148_n 0.00121678f $X=1.825 $Y=0.81 $X2=0 $Y2=0
cc_81 N_A_85_317#_c_93_p N_A1_c_183_n 0.016009f $X=1.825 $Y=0.81 $X2=0 $Y2=0
cc_82 N_A_85_317#_c_93_p N_A1_c_184_n 0.00421546f $X=1.825 $Y=0.81 $X2=0 $Y2=0
cc_83 N_A_85_317#_c_77_n A1 0.00740644f $X=2.01 $Y=2.41 $X2=0 $Y2=0
cc_84 N_A_85_317#_c_68_n N_A1_c_188_n 0.0023592f $X=1.625 $Y=1.67 $X2=0 $Y2=0
cc_85 N_A_85_317#_c_69_n N_A1_c_188_n 0.00597906f $X=1.71 $Y=1.585 $X2=0 $Y2=0
cc_86 N_A_85_317#_c_93_p N_A1_c_188_n 0.00731983f $X=1.825 $Y=0.81 $X2=0 $Y2=0
cc_87 N_A_85_317#_c_69_n N_A1_c_189_n 0.00451908f $X=1.71 $Y=1.585 $X2=0 $Y2=0
cc_88 N_A_85_317#_c_93_p N_A1_c_189_n 0.0102015f $X=1.825 $Y=0.81 $X2=0 $Y2=0
cc_89 N_A_85_317#_c_68_n N_B1_M1000_g 0.00863234f $X=1.625 $Y=1.67 $X2=0 $Y2=0
cc_90 N_A_85_317#_c_75_n N_B1_M1000_g 0.0112858f $X=1.845 $Y=2.41 $X2=0 $Y2=0
cc_91 N_A_85_317#_c_69_n N_B1_M1000_g 6.46889e-19 $X=1.71 $Y=1.585 $X2=0 $Y2=0
cc_92 N_A_85_317#_c_77_n N_B1_M1000_g 0.00599338f $X=2.01 $Y=2.41 $X2=0 $Y2=0
cc_93 N_A_85_317#_c_69_n N_B1_c_242_n 0.00167867f $X=1.71 $Y=1.585 $X2=0 $Y2=0
cc_94 N_A_85_317#_c_93_p N_B1_c_242_n 0.00382187f $X=1.825 $Y=0.81 $X2=0 $Y2=0
cc_95 N_A_85_317#_c_68_n B1 0.0138158f $X=1.625 $Y=1.67 $X2=0 $Y2=0
cc_96 N_A_85_317#_c_69_n B1 0.0299646f $X=1.71 $Y=1.585 $X2=0 $Y2=0
cc_97 N_A_85_317#_c_69_n N_B1_c_244_n 0.0128691f $X=1.71 $Y=1.585 $X2=0 $Y2=0
cc_98 N_A_85_317#_c_93_p N_B1_c_244_n 0.0045498f $X=1.825 $Y=0.81 $X2=0 $Y2=0
cc_99 N_A_85_317#_c_68_n N_B2_c_282_n 2.0352e-19 $X=1.625 $Y=1.67 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_85_317#_c_77_n N_B2_c_282_n 0.00170484f $X=2.01 $Y=2.41 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_85_317#_c_77_n N_B2_M1006_g 0.00794051f $X=2.01 $Y=2.41 $X2=0 $Y2=0
cc_102 N_A_85_317#_c_73_n N_B2_c_285_n 0.0145313f $X=0.72 $Y=2.04 $X2=0 $Y2=0
cc_103 N_A_85_317#_c_68_n N_B2_c_285_n 0.045438f $X=1.625 $Y=1.67 $X2=0 $Y2=0
cc_104 N_A_85_317#_c_75_n N_B2_c_285_n 0.0459007f $X=1.845 $Y=2.41 $X2=0 $Y2=0
cc_105 N_A_85_317#_c_76_n N_B2_c_285_n 4.99486e-19 $X=0.59 $Y=1.75 $X2=0 $Y2=0
cc_106 N_A_85_317#_c_77_n N_B2_c_285_n 0.0229334f $X=2.01 $Y=2.41 $X2=0 $Y2=0
cc_107 N_A_85_317#_M1001_g N_X_c_326_n 0.0032215f $X=0.71 $Y=0.835 $X2=0 $Y2=0
cc_108 N_A_85_317#_c_66_n N_X_c_326_n 0.00268795f $X=0.605 $Y=1.735 $X2=0 $Y2=0
cc_109 N_A_85_317#_c_67_n N_X_c_326_n 0.00307643f $X=0.72 $Y=1.755 $X2=0 $Y2=0
cc_110 N_A_85_317#_M1002_g X 0.0054029f $X=0.66 $Y=2.715 $X2=0 $Y2=0
cc_111 N_A_85_317#_M1001_g X 0.0120094f $X=0.71 $Y=0.835 $X2=0 $Y2=0
cc_112 N_A_85_317#_c_66_n X 0.0164252f $X=0.605 $Y=1.735 $X2=0 $Y2=0
cc_113 N_A_85_317#_c_67_n X 0.0129659f $X=0.72 $Y=1.755 $X2=0 $Y2=0
cc_114 N_A_85_317#_c_73_n X 0.0467967f $X=0.72 $Y=2.04 $X2=0 $Y2=0
cc_115 N_A_85_317#_c_72_n N_X_c_329_n 0.00337708f $X=0.59 $Y=2.255 $X2=0 $Y2=0
cc_116 N_A_85_317#_c_73_n N_X_c_329_n 0.00193458f $X=0.72 $Y=2.04 $X2=0 $Y2=0
cc_117 N_A_85_317#_M1002_g N_VPWR_c_348_n 0.0117381f $X=0.66 $Y=2.715 $X2=0
+ $Y2=0
cc_118 N_A_85_317#_c_73_n N_VPWR_c_348_n 0.0141725f $X=0.72 $Y=2.04 $X2=0 $Y2=0
cc_119 N_A_85_317#_c_75_n N_VPWR_c_348_n 0.00953553f $X=1.845 $Y=2.41 $X2=0
+ $Y2=0
cc_120 N_A_85_317#_M1002_g N_VPWR_c_351_n 0.00532616f $X=0.66 $Y=2.715 $X2=0
+ $Y2=0
cc_121 N_A_85_317#_M1002_g N_VPWR_c_347_n 0.00520409f $X=0.66 $Y=2.715 $X2=0
+ $Y2=0
cc_122 N_A_85_317#_c_73_n N_VPWR_c_347_n 6.40905e-19 $X=0.72 $Y=2.04 $X2=0 $Y2=0
cc_123 N_A_85_317#_c_75_n N_VPWR_c_347_n 0.00947399f $X=1.845 $Y=2.41 $X2=0
+ $Y2=0
cc_124 N_A_85_317#_M1000_d N_A_265_501#_c_384_n 0.0052373f $X=1.755 $Y=2.505
+ $X2=0 $Y2=0
cc_125 N_A_85_317#_c_75_n N_A_265_501#_c_384_n 0.00564952f $X=1.845 $Y=2.41
+ $X2=0 $Y2=0
cc_126 N_A_85_317#_c_77_n N_A_265_501#_c_384_n 0.0228434f $X=2.01 $Y=2.41 $X2=0
+ $Y2=0
cc_127 N_A_85_317#_c_75_n N_A_265_501#_c_385_n 0.0193109f $X=1.845 $Y=2.41 $X2=0
+ $Y2=0
cc_128 N_A_85_317#_c_77_n N_A_265_501#_c_385_n 0.00259213f $X=2.01 $Y=2.41 $X2=0
+ $Y2=0
cc_129 N_A_85_317#_M1001_g N_VGND_c_409_n 0.00523461f $X=0.71 $Y=0.835 $X2=0
+ $Y2=0
cc_130 N_A_85_317#_M1001_g N_VGND_c_411_n 0.00415323f $X=0.71 $Y=0.835 $X2=0
+ $Y2=0
cc_131 N_A_85_317#_M1001_g N_VGND_c_416_n 0.00469432f $X=0.71 $Y=0.835 $X2=0
+ $Y2=0
cc_132 N_A2_c_148_n N_A1_c_184_n 0.0203471f $X=1.16 $Y=1.155 $X2=0 $Y2=0
cc_133 N_A2_c_147_n N_A1_c_188_n 0.0203471f $X=1.16 $Y=1.32 $X2=0 $Y2=0
cc_134 N_A2_M1005_g N_B1_M1000_g 0.0303253f $X=1.25 $Y=2.715 $X2=0 $Y2=0
cc_135 N_A2_c_147_n N_B1_c_244_n 0.0337193f $X=1.16 $Y=1.32 $X2=0 $Y2=0
cc_136 N_A2_M1005_g N_B2_c_285_n 0.010104f $X=1.25 $Y=2.715 $X2=0 $Y2=0
cc_137 A2 N_X_c_326_n 2.69546e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_138 N_A2_c_148_n N_X_c_326_n 3.82584e-19 $X=1.16 $Y=1.155 $X2=0 $Y2=0
cc_139 A2 X 0.00982706f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A2_M1005_g N_VPWR_c_348_n 0.00357217f $X=1.25 $Y=2.715 $X2=0 $Y2=0
cc_141 N_A2_M1005_g N_VPWR_c_353_n 0.00478816f $X=1.25 $Y=2.715 $X2=0 $Y2=0
cc_142 N_A2_M1005_g N_VPWR_c_347_n 0.0044912f $X=1.25 $Y=2.715 $X2=0 $Y2=0
cc_143 N_A2_M1005_g N_A_265_501#_c_385_n 0.00675732f $X=1.25 $Y=2.715 $X2=0
+ $Y2=0
cc_144 A2 N_VGND_c_409_n 0.014802f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_145 N_A2_c_147_n N_VGND_c_409_n 0.00333381f $X=1.16 $Y=1.32 $X2=0 $Y2=0
cc_146 N_A2_c_148_n N_VGND_c_409_n 0.00382662f $X=1.16 $Y=1.155 $X2=0 $Y2=0
cc_147 N_A2_c_148_n N_VGND_c_413_n 0.00415323f $X=1.16 $Y=1.155 $X2=0 $Y2=0
cc_148 N_A2_c_148_n N_VGND_c_416_n 0.00469432f $X=1.16 $Y=1.155 $X2=0 $Y2=0
cc_149 N_A1_c_183_n N_B1_c_242_n 0.00701919f $X=2.445 $Y=0.35 $X2=0 $Y2=0
cc_150 N_A1_c_184_n N_B1_c_242_n 0.00134682f $X=1.7 $Y=0.35 $X2=0 $Y2=0
cc_151 N_A1_c_188_n N_B1_c_242_n 0.0124073f $X=1.7 $Y=0.515 $X2=0 $Y2=0
cc_152 N_A1_c_189_n N_B1_c_242_n 0.00292194f $X=2.825 $Y=1.21 $X2=0 $Y2=0
cc_153 A1 B1 0.0184535f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_154 N_A1_c_189_n B1 0.0159679f $X=2.825 $Y=1.21 $X2=0 $Y2=0
cc_155 N_A1_c_188_n N_B1_c_244_n 0.00594549f $X=1.7 $Y=0.515 $X2=0 $Y2=0
cc_156 N_A1_c_189_n N_B1_c_244_n 2.66291e-19 $X=2.825 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A1_c_191_n N_B2_c_282_n 0.00333459f $X=2.91 $Y=2.28 $X2=-0.19
+ $Y2=-0.245
cc_158 A1 N_B2_c_282_n 0.00577546f $X=3.035 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_159 N_A1_c_187_n N_B2_c_282_n 0.00896733f $X=2.96 $Y=1.775 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A1_c_191_n N_B2_M1006_g 0.0244587f $X=2.91 $Y=2.28 $X2=0 $Y2=0
cc_161 A1 N_B2_M1006_g 0.0047598f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A1_c_183_n N_B2_M1008_g 4.48397e-19 $X=2.445 $Y=0.35 $X2=0 $Y2=0
cc_163 A1 N_B2_M1008_g 0.0138342f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_164 A1 N_B2_M1008_g 0.0108263f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A1_c_187_n N_B2_M1008_g 0.0141231f $X=2.96 $Y=1.775 $X2=0 $Y2=0
cc_166 N_A1_c_189_n N_B2_M1008_g 0.0306054f $X=2.825 $Y=1.21 $X2=0 $Y2=0
cc_167 A1 N_B2_c_285_n 0.0141182f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A1_M1003_g N_VPWR_c_350_n 0.00631532f $X=2.77 $Y=2.755 $X2=0 $Y2=0
cc_169 N_A1_c_191_n N_VPWR_c_350_n 0.00123833f $X=2.91 $Y=2.28 $X2=0 $Y2=0
cc_170 A1 N_VPWR_c_350_n 0.0212931f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_171 N_A1_M1003_g N_VPWR_c_353_n 0.00448616f $X=2.77 $Y=2.755 $X2=0 $Y2=0
cc_172 N_A1_M1003_g N_VPWR_c_347_n 0.0044931f $X=2.77 $Y=2.755 $X2=0 $Y2=0
cc_173 A1 N_VPWR_c_347_n 0.00889181f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_174 N_A1_M1003_g N_A_265_501#_c_386_n 7.56271e-19 $X=2.77 $Y=2.755 $X2=0
+ $Y2=0
cc_175 A1 N_A_265_501#_c_386_n 0.00263682f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A1_c_183_n N_VGND_c_409_n 0.0076368f $X=2.445 $Y=0.35 $X2=0 $Y2=0
cc_177 N_A1_c_184_n N_VGND_c_409_n 0.00558812f $X=1.7 $Y=0.35 $X2=0 $Y2=0
cc_178 N_A1_c_183_n N_VGND_c_410_n 0.0138932f $X=2.445 $Y=0.35 $X2=0 $Y2=0
cc_179 A1 N_VGND_c_410_n 0.0122128f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A1_c_187_n N_VGND_c_410_n 6.81723e-19 $X=2.96 $Y=1.775 $X2=0 $Y2=0
cc_181 N_A1_c_189_n N_VGND_c_410_n 0.0247562f $X=2.825 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A1_c_183_n N_VGND_c_413_n 0.0656671f $X=2.445 $Y=0.35 $X2=0 $Y2=0
cc_183 N_A1_c_184_n N_VGND_c_413_n 0.00651318f $X=1.7 $Y=0.35 $X2=0 $Y2=0
cc_184 N_A1_c_183_n N_VGND_c_416_n 0.0390724f $X=2.445 $Y=0.35 $X2=0 $Y2=0
cc_185 N_A1_c_184_n N_VGND_c_416_n 0.0101042f $X=1.7 $Y=0.35 $X2=0 $Y2=0
cc_186 N_B1_M1000_g N_B2_c_282_n 0.0171755f $X=1.68 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_187 B1 N_B2_c_282_n 0.00245171f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_188 N_B1_c_244_n N_B2_c_282_n 0.00328311f $X=2.06 $Y=1.32 $X2=-0.19
+ $Y2=-0.245
cc_189 N_B1_M1000_g N_B2_M1006_g 0.0161355f $X=1.68 $Y=2.715 $X2=0 $Y2=0
cc_190 N_B1_M1000_g N_B2_M1008_g 0.0012487f $X=1.68 $Y=2.715 $X2=0 $Y2=0
cc_191 N_B1_c_242_n N_B2_M1008_g 0.0578572f $X=2.15 $Y=1.155 $X2=0 $Y2=0
cc_192 B1 N_B2_M1008_g 0.00412677f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_193 N_B1_c_244_n N_B2_M1008_g 0.00205965f $X=2.06 $Y=1.32 $X2=0 $Y2=0
cc_194 N_B1_M1000_g N_B2_c_285_n 0.0110766f $X=1.68 $Y=2.715 $X2=0 $Y2=0
cc_195 B1 N_B2_c_285_n 0.0194221f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_196 N_B1_c_244_n N_B2_c_285_n 0.00604328f $X=2.06 $Y=1.32 $X2=0 $Y2=0
cc_197 N_B1_M1000_g N_VPWR_c_353_n 9.22791e-19 $X=1.68 $Y=2.715 $X2=0 $Y2=0
cc_198 N_B1_M1000_g N_A_265_501#_c_384_n 0.00964875f $X=1.68 $Y=2.715 $X2=0
+ $Y2=0
cc_199 N_B1_M1000_g N_A_265_501#_c_385_n 0.00737326f $X=1.68 $Y=2.715 $X2=0
+ $Y2=0
cc_200 N_B2_M1006_g N_VPWR_c_353_n 0.00282336f $X=2.34 $Y=2.755 $X2=0 $Y2=0
cc_201 N_B2_M1006_g N_VPWR_c_347_n 0.00372843f $X=2.34 $Y=2.755 $X2=0 $Y2=0
cc_202 N_B2_c_282_n N_A_265_501#_c_384_n 0.00147946f $X=2.34 $Y=2.2 $X2=0 $Y2=0
cc_203 N_B2_M1006_g N_A_265_501#_c_384_n 0.013244f $X=2.34 $Y=2.755 $X2=0 $Y2=0
cc_204 N_B2_M1006_g N_A_265_501#_c_385_n 8.82209e-19 $X=2.34 $Y=2.755 $X2=0
+ $Y2=0
cc_205 N_B2_M1006_g N_A_265_501#_c_386_n 2.46537e-19 $X=2.34 $Y=2.755 $X2=0
+ $Y2=0
cc_206 N_B2_M1008_g N_VGND_c_410_n 0.00288905f $X=2.51 $Y=0.835 $X2=0 $Y2=0
cc_207 N_B2_M1008_g N_VGND_c_413_n 5.31375e-19 $X=2.51 $Y=0.835 $X2=0 $Y2=0
cc_208 N_X_c_329_n N_VPWR_c_351_n 0.0107262f $X=0.445 $Y=2.695 $X2=0 $Y2=0
cc_209 N_X_c_329_n N_VPWR_c_347_n 0.0131021f $X=0.445 $Y=2.695 $X2=0 $Y2=0
cc_210 N_X_c_325_n N_VGND_c_416_n 0.00697456f $X=0.325 $Y=0.9 $X2=0 $Y2=0
cc_211 N_X_c_326_n N_VGND_c_416_n 0.0114768f $X=0.475 $Y=0.9 $X2=0 $Y2=0
cc_212 N_VPWR_c_353_n N_A_265_501#_c_384_n 0.0492907f $X=2.84 $Y=3.33 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_347_n N_A_265_501#_c_384_n 0.0299592f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_348_n N_A_265_501#_c_385_n 0.0235017f $X=0.895 $Y=2.78 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_353_n N_A_265_501#_c_385_n 0.021223f $X=2.84 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_347_n N_A_265_501#_c_385_n 0.0125082f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_350_n N_A_265_501#_c_386_n 0.0162385f $X=3.005 $Y=2.82 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_353_n N_A_265_501#_c_386_n 0.0134585f $X=2.84 $Y=3.33 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_347_n N_A_265_501#_c_386_n 0.00793202f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
