* File: sky130_fd_sc_lp__o22ai_0.pxi.spice
* Created: Wed Sep  2 10:20:28 2020
* 
x_PM_SKY130_FD_SC_LP__O22AI_0%B1 N_B1_M1004_g N_B1_c_53_n N_B1_M1001_g
+ N_B1_c_59_n B1 B1 B1 B1 N_B1_c_55_n N_B1_c_56_n PM_SKY130_FD_SC_LP__O22AI_0%B1
x_PM_SKY130_FD_SC_LP__O22AI_0%B2 N_B2_M1007_g N_B2_M1002_g N_B2_c_91_n
+ N_B2_c_96_n B2 B2 B2 N_B2_c_93_n PM_SKY130_FD_SC_LP__O22AI_0%B2
x_PM_SKY130_FD_SC_LP__O22AI_0%A2 N_A2_M1005_g N_A2_M1000_g A2 A2 A2 N_A2_c_136_n
+ PM_SKY130_FD_SC_LP__O22AI_0%A2
x_PM_SKY130_FD_SC_LP__O22AI_0%A1 N_A1_M1003_g N_A1_c_173_n N_A1_M1006_g
+ N_A1_c_174_n N_A1_c_175_n N_A1_c_179_n A1 A1 A1 PM_SKY130_FD_SC_LP__O22AI_0%A1
x_PM_SKY130_FD_SC_LP__O22AI_0%VPWR N_VPWR_M1001_s N_VPWR_M1003_d N_VPWR_c_206_n
+ N_VPWR_c_207_n N_VPWR_c_208_n N_VPWR_c_209_n VPWR N_VPWR_c_210_n
+ N_VPWR_c_205_n PM_SKY130_FD_SC_LP__O22AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O22AI_0%Y N_Y_M1004_d N_Y_M1002_d N_Y_c_237_n N_Y_c_238_n
+ Y Y N_Y_c_240_n PM_SKY130_FD_SC_LP__O22AI_0%Y
x_PM_SKY130_FD_SC_LP__O22AI_0%A_27_85# N_A_27_85#_M1004_s N_A_27_85#_M1007_d
+ N_A_27_85#_M1006_d N_A_27_85#_c_277_n N_A_27_85#_c_278_n N_A_27_85#_c_279_n
+ N_A_27_85#_c_280_n N_A_27_85#_c_281_n N_A_27_85#_c_282_n
+ PM_SKY130_FD_SC_LP__O22AI_0%A_27_85#
x_PM_SKY130_FD_SC_LP__O22AI_0%VGND N_VGND_M1005_d N_VGND_c_314_n VGND
+ N_VGND_c_315_n N_VGND_c_316_n N_VGND_c_317_n N_VGND_c_318_n
+ PM_SKY130_FD_SC_LP__O22AI_0%VGND
cc_1 VNB N_B1_c_53_n 0.00141401f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.12
cc_2 VNB B1 0.0316126f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_3 VNB N_B1_c_55_n 0.0794771f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_4 VNB N_B1_c_56_n 0.017889f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.955
cc_5 VNB N_B2_M1007_g 0.0302778f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.635
cc_6 VNB N_B2_c_91_n 0.0179584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB B2 0.00670532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B2_c_93_n 0.0155944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A2_M1005_g 0.0365198f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.635
cc_10 VNB A2 0.00543059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_c_136_n 0.0252393f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_A1_c_173_n 0.0203548f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.12
cc_13 VNB N_A1_c_174_n 0.0693579f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.735
cc_14 VNB N_A1_c_175_n 0.00710449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A1 0.0186375f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_16 VNB N_VPWR_c_205_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.235 $Y2=1.12
cc_17 VNB N_Y_c_237_n 0.00455734f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.735
cc_18 VNB N_Y_c_238_n 0.00454382f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.735
cc_19 VNB N_A_27_85#_c_277_n 0.0136039f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.195
cc_20 VNB N_A_27_85#_c_278_n 3.9412e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_21 VNB N_A_27_85#_c_279_n 0.0167972f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_27_85#_c_280_n 0.00545059f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_23 VNB N_A_27_85#_c_281_n 0.0156484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_85#_c_282_n 0.0190513f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.12
cc_25 VNB N_VGND_c_314_n 0.00705229f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.27
cc_26 VNB N_VGND_c_315_n 0.039025f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.195
cc_27 VNB N_VGND_c_316_n 0.0177708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_317_n 0.167905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_318_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.12
cc_30 VPB N_B1_c_53_n 0.0239027f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.12
cc_31 VPB N_B1_M1001_g 0.0204367f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.735
cc_32 VPB N_B1_c_59_n 0.0221674f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.195
cc_33 VPB B1 0.0277238f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_34 VPB N_B2_M1002_g 0.0359602f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.735
cc_35 VPB N_B2_c_91_n 0.00379765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_B2_c_96_n 0.015961f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.195
cc_37 VPB B2 0.00670832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A2_M1000_g 0.0467077f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.735
cc_39 VPB A2 0.00415405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A2_c_136_n 0.00644233f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_41 VPB N_A1_M1003_g 0.0365366f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.635
cc_42 VPB N_A1_c_175_n 0.0175532f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A1_c_179_n 0.025715f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.195
cc_44 VPB A1 0.0275258f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_45 VPB N_VPWR_c_206_n 0.022551f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.735
cc_46 VPB N_VPWR_c_207_n 0.026517f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.735
cc_47 VPB N_VPWR_c_208_n 0.0132721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_209_n 0.0357365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_210_n 0.0356524f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_50 VPB N_VPWR_c_205_n 0.0552099f $X=-0.19 $Y=1.655 $X2=0.235 $Y2=1.12
cc_51 VPB N_Y_c_238_n 0.00947777f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=2.735
cc_52 VPB N_Y_c_240_n 0.0169154f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 N_B1_c_56_n N_B2_M1007_g 0.0226497f $X=0.345 $Y=0.955 $X2=0 $Y2=0
cc_54 N_B1_c_53_n N_B2_M1002_g 0.0071316f $X=0.5 $Y=2.12 $X2=0 $Y2=0
cc_55 N_B1_c_59_n N_B2_M1002_g 0.0546071f $X=0.64 $Y=2.195 $X2=0 $Y2=0
cc_56 N_B1_c_53_n N_B2_c_91_n 0.0174084f $X=0.5 $Y=2.12 $X2=0 $Y2=0
cc_57 N_B1_c_53_n B2 6.61775e-19 $X=0.5 $Y=2.12 $X2=0 $Y2=0
cc_58 N_B1_c_55_n B2 5.69816e-19 $X=0.28 $Y=1.12 $X2=0 $Y2=0
cc_59 N_B1_c_55_n N_B2_c_93_n 0.0174084f $X=0.28 $Y=1.12 $X2=0 $Y2=0
cc_60 N_B1_M1001_g N_VPWR_c_206_n 0.0121823f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_61 N_B1_c_59_n N_VPWR_c_206_n 0.00410048f $X=0.64 $Y=2.195 $X2=0 $Y2=0
cc_62 B1 N_VPWR_c_206_n 0.0173159f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_63 N_B1_M1001_g N_VPWR_c_207_n 0.00866029f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_64 N_B1_M1001_g N_VPWR_c_210_n 0.00452967f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_65 N_B1_M1001_g N_VPWR_c_205_n 0.00435436f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_66 B1 N_Y_c_237_n 0.0127189f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_67 N_B1_c_55_n N_Y_c_237_n 0.00151868f $X=0.28 $Y=1.12 $X2=0 $Y2=0
cc_68 N_B1_c_56_n N_Y_c_237_n 0.00355263f $X=0.345 $Y=0.955 $X2=0 $Y2=0
cc_69 N_B1_c_53_n N_Y_c_238_n 0.00903197f $X=0.5 $Y=2.12 $X2=0 $Y2=0
cc_70 N_B1_M1001_g N_Y_c_238_n 0.011996f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_71 N_B1_c_59_n N_Y_c_238_n 0.0119845f $X=0.64 $Y=2.195 $X2=0 $Y2=0
cc_72 B1 N_Y_c_238_n 0.0809122f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_73 N_B1_c_55_n N_Y_c_238_n 0.0140853f $X=0.28 $Y=1.12 $X2=0 $Y2=0
cc_74 N_B1_M1001_g N_Y_c_240_n 0.00206334f $X=0.64 $Y=2.735 $X2=0 $Y2=0
cc_75 B1 N_A_27_85#_M1004_s 0.00254342f $X=0.155 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_76 N_B1_c_56_n N_A_27_85#_c_277_n 0.0110264f $X=0.345 $Y=0.955 $X2=0 $Y2=0
cc_77 B1 N_A_27_85#_c_282_n 0.0214331f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_78 N_B1_c_55_n N_A_27_85#_c_282_n 0.00146666f $X=0.28 $Y=1.12 $X2=0 $Y2=0
cc_79 N_B1_c_56_n N_A_27_85#_c_282_n 0.00841007f $X=0.345 $Y=0.955 $X2=0 $Y2=0
cc_80 N_B1_c_56_n N_VGND_c_315_n 8.57629e-19 $X=0.345 $Y=0.955 $X2=0 $Y2=0
cc_81 B1 N_VGND_c_317_n 0.00167468f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_82 N_B2_M1007_g N_A2_M1005_g 0.0197676f $X=1.005 $Y=0.635 $X2=0 $Y2=0
cc_83 B2 N_A2_M1005_g 0.00630223f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_84 N_B2_c_93_n N_A2_M1005_g 0.0112906f $X=0.98 $Y=1.375 $X2=0 $Y2=0
cc_85 N_B2_M1002_g N_A2_M1000_g 0.0298177f $X=1.03 $Y=2.735 $X2=0 $Y2=0
cc_86 N_B2_c_96_n N_A2_M1000_g 0.0112906f $X=0.98 $Y=1.88 $X2=0 $Y2=0
cc_87 N_B2_M1002_g A2 2.52679e-19 $X=1.03 $Y=2.735 $X2=0 $Y2=0
cc_88 B2 A2 0.0735812f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_89 N_B2_c_93_n A2 5.69077e-19 $X=0.98 $Y=1.375 $X2=0 $Y2=0
cc_90 N_B2_c_91_n N_A2_c_136_n 0.0112906f $X=0.98 $Y=1.715 $X2=0 $Y2=0
cc_91 N_B2_M1002_g N_VPWR_c_206_n 6.56073e-19 $X=1.03 $Y=2.735 $X2=0 $Y2=0
cc_92 N_B2_M1002_g N_VPWR_c_207_n 0.00142016f $X=1.03 $Y=2.735 $X2=0 $Y2=0
cc_93 N_B2_M1002_g N_VPWR_c_210_n 0.00511657f $X=1.03 $Y=2.735 $X2=0 $Y2=0
cc_94 N_B2_M1002_g N_VPWR_c_205_n 0.00585924f $X=1.03 $Y=2.735 $X2=0 $Y2=0
cc_95 N_B2_M1007_g N_Y_c_237_n 0.00724024f $X=1.005 $Y=0.635 $X2=0 $Y2=0
cc_96 B2 N_Y_c_237_n 0.00428008f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_97 N_B2_c_93_n N_Y_c_237_n 0.00376241f $X=0.98 $Y=1.375 $X2=0 $Y2=0
cc_98 N_B2_M1007_g N_Y_c_238_n 0.00377641f $X=1.005 $Y=0.635 $X2=0 $Y2=0
cc_99 N_B2_M1002_g N_Y_c_238_n 0.00408641f $X=1.03 $Y=2.735 $X2=0 $Y2=0
cc_100 B2 N_Y_c_238_n 0.0703431f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B2_c_93_n N_Y_c_238_n 0.00445899f $X=0.98 $Y=1.375 $X2=0 $Y2=0
cc_102 N_B2_M1002_g N_Y_c_240_n 0.0224248f $X=1.03 $Y=2.735 $X2=0 $Y2=0
cc_103 N_B2_c_96_n N_Y_c_240_n 0.00282493f $X=0.98 $Y=1.88 $X2=0 $Y2=0
cc_104 B2 N_Y_c_240_n 0.0329251f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B2_M1007_g N_A_27_85#_c_277_n 0.0130821f $X=1.005 $Y=0.635 $X2=0 $Y2=0
cc_106 N_B2_M1007_g N_A_27_85#_c_278_n 3.20578e-19 $X=1.005 $Y=0.635 $X2=0 $Y2=0
cc_107 N_B2_M1007_g N_A_27_85#_c_280_n 0.00161237f $X=1.005 $Y=0.635 $X2=0 $Y2=0
cc_108 B2 N_A_27_85#_c_280_n 0.0148525f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B2_M1007_g N_A_27_85#_c_282_n 6.48565e-19 $X=1.005 $Y=0.635 $X2=0 $Y2=0
cc_110 N_B2_M1007_g N_VGND_c_315_n 8.63546e-19 $X=1.005 $Y=0.635 $X2=0 $Y2=0
cc_111 A2 N_A1_M1003_g 0.00427264f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_112 N_A2_M1005_g N_A1_c_173_n 0.0177787f $X=1.46 $Y=0.635 $X2=0 $Y2=0
cc_113 N_A2_M1005_g N_A1_c_174_n 0.00670095f $X=1.46 $Y=0.635 $X2=0 $Y2=0
cc_114 A2 N_A1_c_174_n 0.00524314f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A2_c_136_n N_A1_c_174_n 0.0160199f $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_116 N_A2_M1000_g N_A1_c_175_n 0.00520106f $X=1.46 $Y=2.735 $X2=0 $Y2=0
cc_117 N_A2_M1000_g N_A1_c_179_n 0.0658128f $X=1.46 $Y=2.735 $X2=0 $Y2=0
cc_118 A2 N_A1_c_179_n 0.00571804f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_119 N_A2_M1000_g A1 2.81256e-19 $X=1.46 $Y=2.735 $X2=0 $Y2=0
cc_120 A2 A1 0.0724075f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_121 N_A2_c_136_n A1 3.20566e-19 $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_122 N_A2_M1000_g N_VPWR_c_210_n 0.00333733f $X=1.46 $Y=2.735 $X2=0 $Y2=0
cc_123 N_A2_M1000_g N_VPWR_c_205_n 0.00494322f $X=1.46 $Y=2.735 $X2=0 $Y2=0
cc_124 N_A2_M1000_g N_Y_c_240_n 0.0248306f $X=1.46 $Y=2.735 $X2=0 $Y2=0
cc_125 A2 N_Y_c_240_n 0.0272976f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_126 N_A2_c_136_n N_Y_c_240_n 5.74484e-19 $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_127 N_A2_M1005_g N_A_27_85#_c_277_n 0.00114761f $X=1.46 $Y=0.635 $X2=0 $Y2=0
cc_128 N_A2_M1005_g N_A_27_85#_c_278_n 4.88584e-19 $X=1.46 $Y=0.635 $X2=0 $Y2=0
cc_129 N_A2_M1005_g N_A_27_85#_c_279_n 0.0168434f $X=1.46 $Y=0.635 $X2=0 $Y2=0
cc_130 A2 N_A_27_85#_c_279_n 0.0300865f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_131 N_A2_c_136_n N_A_27_85#_c_279_n 9.06402e-19 $X=1.55 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A2_M1005_g N_VGND_c_314_n 0.00565659f $X=1.46 $Y=0.635 $X2=0 $Y2=0
cc_133 N_A2_M1005_g N_VGND_c_315_n 0.00500822f $X=1.46 $Y=0.635 $X2=0 $Y2=0
cc_134 N_A2_M1005_g N_VGND_c_317_n 0.00496652f $X=1.46 $Y=0.635 $X2=0 $Y2=0
cc_135 N_A1_M1003_g N_VPWR_c_209_n 0.0052935f $X=1.85 $Y=2.735 $X2=0 $Y2=0
cc_136 N_A1_c_179_n N_VPWR_c_209_n 0.00311141f $X=2.04 $Y=1.99 $X2=0 $Y2=0
cc_137 A1 N_VPWR_c_209_n 0.0197361f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_138 N_A1_M1003_g N_VPWR_c_210_n 0.00545548f $X=1.85 $Y=2.735 $X2=0 $Y2=0
cc_139 N_A1_M1003_g N_VPWR_c_205_n 0.0110042f $X=1.85 $Y=2.735 $X2=0 $Y2=0
cc_140 N_A1_M1003_g N_Y_c_240_n 0.00590786f $X=1.85 $Y=2.735 $X2=0 $Y2=0
cc_141 N_A1_c_173_n N_A_27_85#_c_279_n 0.0100915f $X=1.925 $Y=0.955 $X2=0 $Y2=0
cc_142 N_A1_c_174_n N_A_27_85#_c_279_n 0.0159767f $X=2.04 $Y=1.54 $X2=0 $Y2=0
cc_143 A1 N_A_27_85#_c_279_n 0.026066f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A1_c_173_n N_A_27_85#_c_281_n 0.001033f $X=1.925 $Y=0.955 $X2=0 $Y2=0
cc_145 N_A1_c_173_n N_VGND_c_314_n 0.011101f $X=1.925 $Y=0.955 $X2=0 $Y2=0
cc_146 N_A1_c_173_n N_VGND_c_316_n 0.00518754f $X=1.925 $Y=0.955 $X2=0 $Y2=0
cc_147 N_A1_c_173_n N_VGND_c_317_n 0.00514264f $X=1.925 $Y=0.955 $X2=0 $Y2=0
cc_148 N_VPWR_c_206_n N_Y_c_238_n 0.00666363f $X=0.357 $Y=2.892 $X2=0 $Y2=0
cc_149 N_VPWR_c_205_n N_Y_c_238_n 0.00449208f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_150 N_VPWR_c_206_n N_Y_c_240_n 0.00799855f $X=0.357 $Y=2.892 $X2=0 $Y2=0
cc_151 N_VPWR_c_207_n N_Y_c_240_n 0.00593525f $X=0.357 $Y=3.245 $X2=0 $Y2=0
cc_152 N_VPWR_c_209_n N_Y_c_240_n 0.00244605f $X=2.065 $Y=2.56 $X2=0 $Y2=0
cc_153 N_VPWR_c_210_n N_Y_c_240_n 0.0454483f $X=1.935 $Y=3.33 $X2=0 $Y2=0
cc_154 N_VPWR_c_205_n N_Y_c_240_n 0.0370982f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_155 A_143_483# N_Y_c_240_n 0.00256757f $X=0.715 $Y=2.415 $X2=1.08 $Y2=2.395
cc_156 N_Y_c_237_n N_A_27_85#_c_277_n 0.0239923f $X=0.64 $Y=1.005 $X2=0 $Y2=0
cc_157 N_Y_c_237_n N_A_27_85#_c_278_n 0.0108148f $X=0.64 $Y=1.005 $X2=0 $Y2=0
cc_158 N_Y_c_237_n N_A_27_85#_c_280_n 0.0110989f $X=0.64 $Y=1.005 $X2=0 $Y2=0
cc_159 N_Y_c_238_n N_A_27_85#_c_280_n 0.00157669f $X=0.64 $Y=2.3 $X2=0 $Y2=0
cc_160 N_A_27_85#_c_277_n N_VGND_c_314_n 0.0144534f $X=1.135 $Y=0.34 $X2=0 $Y2=0
cc_161 N_A_27_85#_c_279_n N_VGND_c_314_n 0.0218367f $X=2.025 $Y=0.955 $X2=0
+ $Y2=0
cc_162 N_A_27_85#_c_277_n N_VGND_c_315_n 0.0601906f $X=1.135 $Y=0.34 $X2=0 $Y2=0
cc_163 N_A_27_85#_c_282_n N_VGND_c_315_n 0.0226635f $X=0.28 $Y=0.34 $X2=0 $Y2=0
cc_164 N_A_27_85#_c_281_n N_VGND_c_316_n 0.00757938f $X=2.14 $Y=0.635 $X2=0
+ $Y2=0
cc_165 N_A_27_85#_c_277_n N_VGND_c_317_n 0.0344916f $X=1.135 $Y=0.34 $X2=0 $Y2=0
cc_166 N_A_27_85#_c_281_n N_VGND_c_317_n 0.00942937f $X=2.14 $Y=0.635 $X2=0
+ $Y2=0
cc_167 N_A_27_85#_c_282_n N_VGND_c_317_n 0.0125932f $X=0.28 $Y=0.34 $X2=0 $Y2=0
