* File: sky130_fd_sc_lp__invlp_4.pxi.spice
* Created: Wed Sep  2 09:57:14 2020
* 
x_PM_SKY130_FD_SC_LP__INVLP_4%A N_A_M1000_g N_A_M1002_g N_A_M1009_g N_A_M1004_g
+ N_A_M1005_g N_A_M1011_g N_A_M1001_g N_A_M1003_g N_A_M1008_g N_A_M1006_g
+ N_A_M1007_g N_A_M1010_g N_A_M1014_g N_A_M1013_g N_A_M1012_g N_A_M1015_g
+ N_A_c_65_n N_A_c_66_n A A A N_A_c_78_n N_A_c_67_n N_A_c_80_n
+ PM_SKY130_FD_SC_LP__INVLP_4%A
x_PM_SKY130_FD_SC_LP__INVLP_4%VPWR N_VPWR_M1002_d N_VPWR_M1004_d N_VPWR_M1012_d
+ N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n N_VPWR_c_230_n N_VPWR_c_231_n
+ VPWR N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_226_n
+ PM_SKY130_FD_SC_LP__INVLP_4%VPWR
x_PM_SKY130_FD_SC_LP__INVLP_4%A_118_367# N_A_118_367#_M1002_s
+ N_A_118_367#_M1005_s N_A_118_367#_M1008_d N_A_118_367#_M1013_d
+ N_A_118_367#_c_283_n N_A_118_367#_c_287_n N_A_118_367#_c_290_n
+ N_A_118_367#_c_292_n N_A_118_367#_c_296_n N_A_118_367#_c_298_n
+ N_A_118_367#_c_300_n N_A_118_367#_c_302_n N_A_118_367#_c_304_n
+ N_A_118_367#_c_305_n N_A_118_367#_c_308_n N_A_118_367#_c_309_n
+ PM_SKY130_FD_SC_LP__INVLP_4%A_118_367#
x_PM_SKY130_FD_SC_LP__INVLP_4%Y N_Y_M1003_s N_Y_M1007_s N_Y_M1001_s N_Y_M1010_s
+ N_Y_c_346_n N_Y_c_341_n N_Y_c_356_n N_Y_c_396_n N_Y_c_419_p N_Y_c_342_n
+ N_Y_c_367_n N_Y_c_372_n N_Y_c_373_n N_Y_c_376_n N_Y_c_343_n N_Y_c_344_n
+ N_Y_c_385_n N_Y_c_345_n Y PM_SKY130_FD_SC_LP__INVLP_4%Y
x_PM_SKY130_FD_SC_LP__INVLP_4%VGND N_VGND_M1000_d N_VGND_M1009_d N_VGND_M1015_d
+ N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n
+ VGND N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n
+ PM_SKY130_FD_SC_LP__INVLP_4%VGND
x_PM_SKY130_FD_SC_LP__INVLP_4%A_114_53# N_A_114_53#_M1000_s N_A_114_53#_M1011_s
+ N_A_114_53#_M1006_d N_A_114_53#_M1014_d N_A_114_53#_c_480_n
+ N_A_114_53#_c_489_n N_A_114_53#_c_493_n N_A_114_53#_c_497_n
+ N_A_114_53#_c_481_n N_A_114_53#_c_482_n N_A_114_53#_c_483_n
+ N_A_114_53#_c_484_n N_A_114_53#_c_485_n PM_SKY130_FD_SC_LP__INVLP_4%A_114_53#
cc_1 VNB N_A_M1000_g 0.0317431f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.685
cc_2 VNB N_A_M1009_g 0.0233467f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.685
cc_3 VNB N_A_M1011_g 0.0240921f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.685
cc_4 VNB N_A_M1003_g 0.0222343f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.685
cc_5 VNB N_A_M1006_g 0.0222372f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.685
cc_6 VNB N_A_M1007_g 0.0232397f $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=0.685
cc_7 VNB N_A_M1014_g 0.0245555f $X=-0.19 $Y=-0.245 $X2=3.285 $Y2=0.685
cc_8 VNB N_A_M1015_g 0.0327026f $X=-0.19 $Y=-0.245 $X2=3.785 $Y2=0.685
cc_9 VNB N_A_c_65_n 0.0125848f $X=-0.19 $Y=-0.245 $X2=3.93 $Y2=1.51
cc_10 VNB N_A_c_66_n 0.179787f $X=-0.19 $Y=-0.245 $X2=3.93 $Y2=1.51
cc_11 VNB N_A_c_67_n 9.31901e-19 $X=-0.19 $Y=-0.245 $X2=2 $Y2=1.562
cc_12 VNB N_VPWR_c_226_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=2.465
cc_13 VNB N_Y_c_341_n 0.00625221f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.465
cc_14 VNB N_Y_c_342_n 0.00545048f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.675
cc_15 VNB N_Y_c_343_n 0.00288027f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.345
cc_16 VNB N_Y_c_344_n 0.00482817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_345_n 0.00124913f $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=0.685
cc_18 VNB N_VGND_c_426_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.685
cc_19 VNB N_VGND_c_427_n 0.0486288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_428_n 0.00645394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_429_n 0.0119539f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=2.465
cc_22 VNB N_VGND_c_430_n 0.0424868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_431_n 0.0175438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_432_n 0.0586603f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.345
cc_25 VNB N_VGND_c_433_n 0.00630919f $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=1.345
cc_26 VNB N_VGND_c_434_n 0.248702f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=1.675
cc_27 VNB N_A_114_53#_c_480_n 0.00203831f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.465
cc_28 VNB N_A_114_53#_c_481_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.685
cc_29 VNB N_A_114_53#_c_482_n 0.00203277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_114_53#_c_483_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.465
cc_31 VNB N_A_114_53#_c_484_n 0.00203277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_114_53#_c_485_n 0.0049581f $X=-0.19 $Y=-0.245 $X2=2.305 $Y2=2.465
cc_33 VPB N_A_M1002_g 0.0254819f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.465
cc_34 VPB N_A_M1004_g 0.0184913f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_35 VPB N_A_M1005_g 0.0186707f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=2.465
cc_36 VPB N_A_M1001_g 0.01866f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.465
cc_37 VPB N_A_M1008_g 0.0194537f $X=-0.19 $Y=1.655 $X2=2.305 $Y2=2.465
cc_38 VPB N_A_M1010_g 0.0198938f $X=-0.19 $Y=1.655 $X2=2.805 $Y2=2.465
cc_39 VPB N_A_M1013_g 0.0195323f $X=-0.19 $Y=1.655 $X2=3.305 $Y2=2.465
cc_40 VPB N_A_M1012_g 0.0261051f $X=-0.19 $Y=1.655 $X2=3.735 $Y2=2.465
cc_41 VPB N_A_c_65_n 7.73822e-19 $X=-0.19 $Y=1.655 $X2=3.93 $Y2=1.51
cc_42 VPB N_A_c_66_n 0.0431164f $X=-0.19 $Y=1.655 $X2=3.93 $Y2=1.51
cc_43 VPB N_A_c_78_n 0.00359974f $X=-0.19 $Y=1.655 $X2=2.538 $Y2=1.562
cc_44 VPB N_A_c_67_n 0.00374338f $X=-0.19 $Y=1.655 $X2=2 $Y2=1.562
cc_45 VPB N_A_c_80_n 0.00179264f $X=-0.19 $Y=1.655 $X2=2.755 $Y2=1.562
cc_46 VPB N_VPWR_c_227_n 0.0112901f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.685
cc_47 VPB N_VPWR_c_228_n 0.0617459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_229_n 0.00231123f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=2.465
cc_49 VPB N_VPWR_c_230_n 0.0128252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_231_n 0.0535687f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=0.685
cc_51 VPB N_VPWR_c_232_n 0.0158404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_233_n 0.0609301f $X=-0.19 $Y=1.655 $X2=2.305 $Y2=1.675
cc_53 VPB N_VPWR_c_234_n 0.00356964f $X=-0.19 $Y=1.655 $X2=2.785 $Y2=0.685
cc_54 VPB N_VPWR_c_226_n 0.0469265f $X=-0.19 $Y=1.655 $X2=2.805 $Y2=2.465
cc_55 VPB N_A_118_367#_c_283_n 0.00305603f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_56 VPB N_Y_c_346_n 0.00267097f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_57 N_A_M1002_g N_VPWR_c_228_n 0.00721235f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_58 N_A_M1002_g N_VPWR_c_229_n 6.42741e-19 $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A_M1004_g N_VPWR_c_229_n 0.00943178f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_60 N_A_M1005_g N_VPWR_c_229_n 0.00313805f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_61 N_A_M1012_g N_VPWR_c_231_n 0.0288467f $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_62 N_A_c_65_n N_VPWR_c_231_n 0.0192431f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_63 N_A_c_66_n N_VPWR_c_231_n 0.00554992f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_64 N_A_M1002_g N_VPWR_c_232_n 0.0054895f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_65 N_A_M1004_g N_VPWR_c_232_n 0.00486043f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_M1005_g N_VPWR_c_233_n 0.00547432f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_VPWR_c_233_n 0.00357842f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A_M1008_g N_VPWR_c_233_n 0.00357877f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_69 N_A_M1010_g N_VPWR_c_233_n 0.00357842f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_M1013_g N_VPWR_c_233_n 0.00357877f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_71 N_A_M1012_g N_VPWR_c_233_n 0.00547432f $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_72 N_A_M1002_g N_VPWR_c_226_n 0.0107613f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_VPWR_c_226_n 0.00824727f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_74 N_A_M1005_g N_VPWR_c_226_n 0.0098633f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_75 N_A_M1001_g N_VPWR_c_226_n 0.00553547f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_76 N_A_M1008_g N_VPWR_c_226_n 0.0057905f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A_M1010_g N_VPWR_c_226_n 0.00570659f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_M1013_g N_VPWR_c_226_n 0.00553549f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A_M1012_g N_VPWR_c_226_n 0.0109358f $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A_M1002_g N_A_118_367#_c_283_n 0.00727789f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_81 N_A_M1004_g N_A_118_367#_c_283_n 4.75665e-19 $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A_c_66_n N_A_118_367#_c_283_n 0.00287442f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_83 N_A_M1004_g N_A_118_367#_c_287_n 0.0168101f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_84 N_A_M1005_g N_A_118_367#_c_287_n 0.01115f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_c_66_n N_A_118_367#_c_287_n 2.86047e-19 $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_86 N_A_M1005_g N_A_118_367#_c_290_n 7.32094e-19 $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_M1001_g N_A_118_367#_c_290_n 0.00209265f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_88 N_A_M1004_g N_A_118_367#_c_292_n 6.18158e-19 $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_M1005_g N_A_118_367#_c_292_n 0.00677393f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A_M1001_g N_A_118_367#_c_292_n 0.00695801f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_91 N_A_M1008_g N_A_118_367#_c_292_n 4.62714e-19 $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A_M1001_g N_A_118_367#_c_296_n 0.0109138f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_93 N_A_M1008_g N_A_118_367#_c_296_n 0.0143648f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_M1005_g N_A_118_367#_c_298_n 0.00197018f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A_M1001_g N_A_118_367#_c_298_n 5.89773e-19 $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A_M1010_g N_A_118_367#_c_300_n 0.00892877f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A_M1013_g N_A_118_367#_c_300_n 8.75074e-19 $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_M1010_g N_A_118_367#_c_302_n 0.0109138f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_M1013_g N_A_118_367#_c_302_n 0.0118963f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_M1012_g N_A_118_367#_c_304_n 0.00202381f $X=3.735 $Y=2.465 $X2=0
+ $Y2=0
cc_101 N_A_M1012_g N_A_118_367#_c_305_n 0.0127124f $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_c_65_n N_A_118_367#_c_305_n 0.0177688f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_103 N_A_c_66_n N_A_118_367#_c_305_n 0.00232957f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_104 N_A_M1002_g N_A_118_367#_c_308_n 0.00944473f $X=0.515 $Y=2.465 $X2=0
+ $Y2=0
cc_105 N_A_M1010_g N_A_118_367#_c_309_n 5.89773e-19 $X=2.805 $Y=2.465 $X2=0
+ $Y2=0
cc_106 N_A_M1004_g N_Y_c_346_n 0.00414614f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_M1005_g N_Y_c_346_n 0.00481775f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_c_66_n N_Y_c_346_n 0.0212306f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A_c_67_n N_Y_c_346_n 0.00535098f $X=2 $Y=1.562 $X2=0 $Y2=0
cc_110 N_A_M1011_g N_Y_c_341_n 0.0104123f $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_111 N_A_M1003_g N_Y_c_341_n 0.0114627f $X=1.925 $Y=0.685 $X2=0 $Y2=0
cc_112 N_A_c_66_n N_Y_c_341_n 0.00546875f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_113 N_A_c_78_n N_Y_c_341_n 0.0041468f $X=2.538 $Y=1.562 $X2=0 $Y2=0
cc_114 N_A_c_67_n N_Y_c_341_n 0.0460352f $X=2 $Y=1.562 $X2=0 $Y2=0
cc_115 N_A_M1005_g N_Y_c_356_n 0.0129088f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_M1001_g N_Y_c_356_n 0.0146497f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_c_66_n N_Y_c_356_n 5.55909e-19 $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A_c_67_n N_Y_c_356_n 0.0317143f $X=2 $Y=1.562 $X2=0 $Y2=0
cc_119 N_A_M1006_g N_Y_c_342_n 0.0115018f $X=2.355 $Y=0.685 $X2=0 $Y2=0
cc_120 N_A_M1007_g N_Y_c_342_n 0.0125117f $X=2.785 $Y=0.685 $X2=0 $Y2=0
cc_121 N_A_M1014_g N_Y_c_342_n 0.00434728f $X=3.285 $Y=0.685 $X2=0 $Y2=0
cc_122 N_A_M1015_g N_Y_c_342_n 2.71338e-19 $X=3.785 $Y=0.685 $X2=0 $Y2=0
cc_123 N_A_c_65_n N_Y_c_342_n 0.0273607f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_124 N_A_c_66_n N_Y_c_342_n 0.00625627f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_125 N_A_c_78_n N_Y_c_342_n 0.0506943f $X=2.538 $Y=1.562 $X2=0 $Y2=0
cc_126 N_A_M1008_g N_Y_c_367_n 0.0115433f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_M1010_g N_Y_c_367_n 0.0155875f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_c_65_n N_Y_c_367_n 0.00720235f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A_c_66_n N_Y_c_367_n 9.26083e-19 $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A_c_78_n N_Y_c_367_n 0.0346418f $X=2.538 $Y=1.562 $X2=0 $Y2=0
cc_131 N_A_M1014_g N_Y_c_372_n 0.00536639f $X=3.285 $Y=0.685 $X2=0 $Y2=0
cc_132 N_A_M1013_g N_Y_c_373_n 0.00314442f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A_c_65_n N_Y_c_373_n 0.024044f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A_c_66_n N_Y_c_373_n 0.00403915f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A_M1013_g N_Y_c_376_n 0.0087304f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_M1012_g N_Y_c_376_n 2.37719e-19 $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_M1009_g N_Y_c_343_n 0.00306462f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_138 N_A_M1011_g N_Y_c_343_n 0.00381768f $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_139 N_A_c_66_n N_Y_c_343_n 0.00477392f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_140 N_A_c_67_n N_Y_c_343_n 0.0251038f $X=2 $Y=1.562 $X2=0 $Y2=0
cc_141 N_A_M1000_g N_Y_c_344_n 0.00482622f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_142 N_A_M1009_g N_Y_c_344_n 0.00792459f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_143 N_A_c_66_n N_Y_c_344_n 0.0221477f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A_M1008_g N_Y_c_385_n 0.00976964f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1010_g N_Y_c_385_n 5.97816e-19 $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_c_66_n N_Y_c_385_n 0.00104552f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_147 N_A_c_78_n N_Y_c_385_n 0.0197412f $X=2.538 $Y=1.562 $X2=0 $Y2=0
cc_148 N_A_c_67_n N_Y_c_385_n 0.00612547f $X=2 $Y=1.562 $X2=0 $Y2=0
cc_149 N_A_c_66_n N_Y_c_345_n 0.00251211f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A_c_78_n N_Y_c_345_n 0.0144295f $X=2.538 $Y=1.562 $X2=0 $Y2=0
cc_151 N_A_M1000_g N_VGND_c_427_n 0.00822358f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_152 N_A_M1009_g N_VGND_c_428_n 0.0043892f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_153 N_A_M1011_g N_VGND_c_428_n 0.00438904f $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_154 N_A_M1015_g N_VGND_c_430_n 0.00787605f $X=3.785 $Y=0.685 $X2=0 $Y2=0
cc_155 N_A_c_65_n N_VGND_c_430_n 0.0124468f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_156 N_A_c_66_n N_VGND_c_430_n 0.00406184f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A_M1000_g N_VGND_c_431_n 0.00520505f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_158 N_A_M1009_g N_VGND_c_431_n 0.00395047f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_159 N_A_M1011_g N_VGND_c_432_n 0.003936f $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_160 N_A_M1003_g N_VGND_c_432_n 0.0033828f $X=1.925 $Y=0.685 $X2=0 $Y2=0
cc_161 N_A_M1006_g N_VGND_c_432_n 0.0033828f $X=2.355 $Y=0.685 $X2=0 $Y2=0
cc_162 N_A_M1007_g N_VGND_c_432_n 0.0033828f $X=2.785 $Y=0.685 $X2=0 $Y2=0
cc_163 N_A_M1014_g N_VGND_c_432_n 0.00338313f $X=3.285 $Y=0.685 $X2=0 $Y2=0
cc_164 N_A_M1015_g N_VGND_c_432_n 0.00519058f $X=3.785 $Y=0.685 $X2=0 $Y2=0
cc_165 N_A_M1000_g N_VGND_c_434_n 0.0104451f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_166 N_A_M1009_g N_VGND_c_434_n 0.00576893f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_167 N_A_M1011_g N_VGND_c_434_n 0.00577802f $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_168 N_A_M1003_g N_VGND_c_434_n 0.00509122f $X=1.925 $Y=0.685 $X2=0 $Y2=0
cc_169 N_A_M1006_g N_VGND_c_434_n 0.00509122f $X=2.355 $Y=0.685 $X2=0 $Y2=0
cc_170 N_A_M1007_g N_VGND_c_434_n 0.00523601f $X=2.785 $Y=0.685 $X2=0 $Y2=0
cc_171 N_A_M1014_g N_VGND_c_434_n 0.00538083f $X=3.285 $Y=0.685 $X2=0 $Y2=0
cc_172 N_A_M1015_g N_VGND_c_434_n 0.0105813f $X=3.785 $Y=0.685 $X2=0 $Y2=0
cc_173 N_A_M1000_g N_A_114_53#_c_480_n 0.00518099f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_174 N_A_M1009_g N_A_114_53#_c_480_n 0.00663493f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_175 N_A_M1011_g N_A_114_53#_c_480_n 5.79146e-19 $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_176 N_A_M1009_g N_A_114_53#_c_489_n 0.0100974f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_177 N_A_M1011_g N_A_114_53#_c_489_n 0.011185f $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_178 N_A_M1003_g N_A_114_53#_c_489_n 0.00326815f $X=1.925 $Y=0.685 $X2=0 $Y2=0
cc_179 N_A_c_66_n N_A_114_53#_c_489_n 5.8517e-19 $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A_M1000_g N_A_114_53#_c_493_n 0.00502503f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_181 N_A_M1009_g N_A_114_53#_c_493_n 0.00421868f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_182 N_A_M1011_g N_A_114_53#_c_493_n 7.79642e-19 $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_183 N_A_c_66_n N_A_114_53#_c_493_n 5.35171e-19 $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_184 N_A_M1009_g N_A_114_53#_c_497_n 5.45135e-19 $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_185 N_A_M1011_g N_A_114_53#_c_497_n 0.00415295f $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_186 N_A_M1003_g N_A_114_53#_c_497_n 0.0036618f $X=1.925 $Y=0.685 $X2=0 $Y2=0
cc_187 N_A_M1006_g N_A_114_53#_c_497_n 5.20259e-19 $X=2.355 $Y=0.685 $X2=0 $Y2=0
cc_188 N_A_M1003_g N_A_114_53#_c_481_n 0.00827312f $X=1.925 $Y=0.685 $X2=0 $Y2=0
cc_189 N_A_M1006_g N_A_114_53#_c_481_n 0.00827312f $X=2.355 $Y=0.685 $X2=0 $Y2=0
cc_190 N_A_M1011_g N_A_114_53#_c_482_n 0.00310094f $X=1.495 $Y=0.685 $X2=0 $Y2=0
cc_191 N_A_M1003_g N_A_114_53#_c_482_n 0.00172424f $X=1.925 $Y=0.685 $X2=0 $Y2=0
cc_192 N_A_M1007_g N_A_114_53#_c_483_n 0.00866637f $X=2.785 $Y=0.685 $X2=0 $Y2=0
cc_193 N_A_M1014_g N_A_114_53#_c_483_n 0.0142587f $X=3.285 $Y=0.685 $X2=0 $Y2=0
cc_194 N_A_M1003_g N_A_114_53#_c_484_n 5.71288e-19 $X=1.925 $Y=0.685 $X2=0 $Y2=0
cc_195 N_A_M1006_g N_A_114_53#_c_484_n 0.00644132f $X=2.355 $Y=0.685 $X2=0 $Y2=0
cc_196 N_A_M1007_g N_A_114_53#_c_484_n 0.00684043f $X=2.785 $Y=0.685 $X2=0 $Y2=0
cc_197 N_A_M1014_g N_A_114_53#_c_484_n 6.22096e-19 $X=3.285 $Y=0.685 $X2=0 $Y2=0
cc_198 N_A_M1014_g N_A_114_53#_c_485_n 0.00371159f $X=3.285 $Y=0.685 $X2=0 $Y2=0
cc_199 N_A_M1015_g N_A_114_53#_c_485_n 0.0122586f $X=3.785 $Y=0.685 $X2=0 $Y2=0
cc_200 N_A_c_65_n N_A_114_53#_c_485_n 0.022699f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_201 N_A_c_66_n N_A_114_53#_c_485_n 0.00411924f $X=3.93 $Y=1.51 $X2=0 $Y2=0
cc_202 N_VPWR_c_226_n N_A_118_367#_M1002_s 0.0041489f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_203 N_VPWR_c_226_n N_A_118_367#_M1005_s 0.00223559f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_226_n N_A_118_367#_M1008_d 0.00280658f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_226_n N_A_118_367#_M1013_d 0.00223562f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_228_n N_A_118_367#_c_283_n 0.0170091f $X=0.3 $Y=1.98 $X2=0 $Y2=0
cc_207 N_VPWR_M1004_d N_A_118_367#_c_287_n 0.00338954f $X=1.02 $Y=1.835 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_229_n N_A_118_367#_c_287_n 0.0153337f $X=1.16 $Y=2.87 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_233_n N_A_118_367#_c_296_n 0.0374555f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_226_n N_A_118_367#_c_296_n 0.0239316f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_233_n N_A_118_367#_c_298_n 0.01906f $X=3.855 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_226_n N_A_118_367#_c_298_n 0.0124545f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_233_n N_A_118_367#_c_302_n 0.037782f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_226_n N_A_118_367#_c_302_n 0.024237f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_215 N_VPWR_c_233_n N_A_118_367#_c_304_n 0.0154369f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_216 N_VPWR_c_226_n N_A_118_367#_c_304_n 0.00952129f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_232_n N_A_118_367#_c_308_n 0.0153332f $X=0.995 $Y=3.33 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_226_n N_A_118_367#_c_308_n 0.00945339f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_233_n N_A_118_367#_c_309_n 0.0207136f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_226_n N_A_118_367#_c_309_n 0.0126421f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_226_n N_Y_M1001_s 0.00281482f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_226_n N_Y_M1010_s 0.00281482f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_M1004_d N_Y_c_346_n 0.0014879f $X=1.02 $Y=1.835 $X2=0 $Y2=0
cc_224 N_VPWR_M1004_d N_Y_c_356_n 0.00131791f $X=1.02 $Y=1.835 $X2=0 $Y2=0
cc_225 N_VPWR_M1004_d N_Y_c_396_n 0.001903f $X=1.02 $Y=1.835 $X2=0 $Y2=0
cc_226 N_A_118_367#_c_296_n N_Y_M1001_s 0.00472489f $X=2.425 $Y=2.99 $X2=0 $Y2=0
cc_227 N_A_118_367#_c_302_n N_Y_M1010_s 0.00472489f $X=3.435 $Y=2.99 $X2=0 $Y2=0
cc_228 N_A_118_367#_c_283_n N_Y_c_346_n 0.0011916f $X=0.73 $Y=1.98 $X2=0 $Y2=0
cc_229 N_A_118_367#_M1005_s N_Y_c_356_n 0.00346799f $X=1.45 $Y=1.835 $X2=0 $Y2=0
cc_230 N_A_118_367#_c_287_n N_Y_c_356_n 0.0104361f $X=1.425 $Y=2.375 $X2=0 $Y2=0
cc_231 N_A_118_367#_c_290_n N_Y_c_356_n 0.01723f $X=1.59 $Y=2.46 $X2=0 $Y2=0
cc_232 N_A_118_367#_c_287_n N_Y_c_396_n 0.0111826f $X=1.425 $Y=2.375 $X2=0 $Y2=0
cc_233 N_A_118_367#_M1008_d N_Y_c_367_n 0.00469238f $X=2.38 $Y=1.835 $X2=0 $Y2=0
cc_234 N_A_118_367#_c_300_n N_Y_c_367_n 0.0209867f $X=2.59 $Y=2.455 $X2=0 $Y2=0
cc_235 N_A_118_367#_c_302_n N_Y_c_376_n 0.0196355f $X=3.435 $Y=2.99 $X2=0 $Y2=0
cc_236 N_A_118_367#_c_283_n N_Y_c_344_n 0.00902076f $X=0.73 $Y=1.98 $X2=0 $Y2=0
cc_237 N_A_118_367#_c_296_n N_Y_c_385_n 0.0196355f $X=2.425 $Y=2.99 $X2=0 $Y2=0
cc_238 N_Y_c_341_n N_VGND_M1009_d 0.00194702f $X=2.055 $Y=1.09 $X2=0 $Y2=0
cc_239 N_Y_c_343_n N_VGND_M1009_d 0.00217186f $X=1.13 $Y=1.09 $X2=0 $Y2=0
cc_240 N_Y_c_341_n N_A_114_53#_M1011_s 0.00176461f $X=2.055 $Y=1.09 $X2=0 $Y2=0
cc_241 N_Y_c_342_n N_A_114_53#_M1006_d 0.00176461f $X=2.905 $Y=1.09 $X2=0 $Y2=0
cc_242 N_Y_c_341_n N_A_114_53#_c_489_n 0.0362786f $X=2.055 $Y=1.09 $X2=0 $Y2=0
cc_243 N_Y_c_343_n N_A_114_53#_c_489_n 0.0127733f $X=1.13 $Y=1.09 $X2=0 $Y2=0
cc_244 N_Y_c_344_n N_A_114_53#_c_489_n 0.00598592f $X=1.045 $Y=1.295 $X2=0 $Y2=0
cc_245 N_Y_c_344_n N_A_114_53#_c_493_n 0.0190512f $X=1.045 $Y=1.295 $X2=0 $Y2=0
cc_246 N_Y_M1003_s N_A_114_53#_c_481_n 0.00176461f $X=2 $Y=0.265 $X2=0 $Y2=0
cc_247 N_Y_c_341_n N_A_114_53#_c_481_n 0.00305513f $X=2.055 $Y=1.09 $X2=0 $Y2=0
cc_248 N_Y_c_419_p N_A_114_53#_c_481_n 0.0124813f $X=2.14 $Y=0.86 $X2=0 $Y2=0
cc_249 N_Y_c_342_n N_A_114_53#_c_481_n 0.00305513f $X=2.905 $Y=1.09 $X2=0 $Y2=0
cc_250 N_Y_M1007_s N_A_114_53#_c_483_n 0.00250873f $X=2.86 $Y=0.265 $X2=0 $Y2=0
cc_251 N_Y_c_342_n N_A_114_53#_c_483_n 0.00306745f $X=2.905 $Y=1.09 $X2=0 $Y2=0
cc_252 N_Y_c_372_n N_A_114_53#_c_483_n 0.0194333f $X=3.07 $Y=0.86 $X2=0 $Y2=0
cc_253 N_Y_c_342_n N_A_114_53#_c_484_n 0.0168576f $X=2.905 $Y=1.09 $X2=0 $Y2=0
cc_254 N_Y_c_342_n N_A_114_53#_c_485_n 0.00584871f $X=2.905 $Y=1.09 $X2=0 $Y2=0
cc_255 N_VGND_c_427_n N_A_114_53#_c_480_n 0.0150039f $X=0.28 $Y=0.41 $X2=0 $Y2=0
cc_256 N_VGND_c_428_n N_A_114_53#_c_480_n 0.00937982f $X=1.21 $Y=0.41 $X2=0
+ $Y2=0
cc_257 N_VGND_c_431_n N_A_114_53#_c_480_n 0.0233446f $X=1.045 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_434_n N_A_114_53#_c_480_n 0.0125323f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_259 N_VGND_M1009_d N_A_114_53#_c_489_n 0.00667164f $X=1 $Y=0.265 $X2=0 $Y2=0
cc_260 N_VGND_c_428_n N_A_114_53#_c_489_n 0.0235432f $X=1.21 $Y=0.41 $X2=0 $Y2=0
cc_261 N_VGND_c_431_n N_A_114_53#_c_489_n 0.00229766f $X=1.045 $Y=0 $X2=0 $Y2=0
cc_262 N_VGND_c_432_n N_A_114_53#_c_489_n 0.00229766f $X=3.915 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_434_n N_A_114_53#_c_489_n 0.00970368f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_264 N_VGND_c_432_n N_A_114_53#_c_481_n 0.0333615f $X=3.915 $Y=0 $X2=0 $Y2=0
cc_265 N_VGND_c_434_n N_A_114_53#_c_481_n 0.0187823f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_c_428_n N_A_114_53#_c_482_n 0.00753712f $X=1.21 $Y=0.41 $X2=0
+ $Y2=0
cc_267 N_VGND_c_432_n N_A_114_53#_c_482_n 0.0232022f $X=3.915 $Y=0 $X2=0 $Y2=0
cc_268 N_VGND_c_434_n N_A_114_53#_c_482_n 0.0125478f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_c_432_n N_A_114_53#_c_483_n 0.0423044f $X=3.915 $Y=0 $X2=0 $Y2=0
cc_270 N_VGND_c_434_n N_A_114_53#_c_483_n 0.0239316f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_271 N_VGND_c_432_n N_A_114_53#_c_484_n 0.0232038f $X=3.915 $Y=0 $X2=0 $Y2=0
cc_272 N_VGND_c_434_n N_A_114_53#_c_484_n 0.0125481f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_273 N_VGND_c_430_n N_A_114_53#_c_485_n 0.0329656f $X=4 $Y=0.41 $X2=0 $Y2=0
cc_274 N_VGND_c_432_n N_A_114_53#_c_485_n 0.0235688f $X=3.915 $Y=0 $X2=0 $Y2=0
cc_275 N_VGND_c_434_n N_A_114_53#_c_485_n 0.0127152f $X=4.08 $Y=0 $X2=0 $Y2=0
