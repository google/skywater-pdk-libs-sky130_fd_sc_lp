# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a2bb2oi_0
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a2bb2oi_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.455000 1.840000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.780000 1.365000 1.435000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 0.780000 3.275000 1.475000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055000 0.780000 2.550000 1.475000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.287200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.570000 0.780000 1.885000 1.915000 ;
        RECT 1.570000 1.915000 1.935000 2.950000 ;
        RECT 1.715000 0.275000 2.280000 0.610000 ;
        RECT 1.715000 0.610000 1.885000 0.780000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.095000  0.085000 0.385000 0.610000 ;
      RECT 0.095000  2.115000 0.425000 3.245000 ;
      RECT 0.555000  0.280000 0.830000 0.610000 ;
      RECT 0.625000  0.610000 0.830000 1.645000 ;
      RECT 0.625000  1.645000 1.400000 2.155000 ;
      RECT 0.885000  2.155000 1.215000 2.795000 ;
      RECT 1.000000  0.085000 1.545000 0.610000 ;
      RECT 2.105000  1.645000 3.265000 1.815000 ;
      RECT 2.105000  1.815000 2.335000 2.595000 ;
      RECT 2.505000  1.985000 2.835000 3.245000 ;
      RECT 2.910000  0.085000 3.240000 0.610000 ;
      RECT 3.015000  1.815000 3.265000 2.595000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__a2bb2oi_0
END LIBRARY
