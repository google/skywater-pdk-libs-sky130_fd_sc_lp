* File: sky130_fd_sc_lp__and2_2.pex.spice
* Created: Wed Sep  2 09:30:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2_2%A 1 3 4 6 10 11 12 16 17
r34 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r35 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.665
r36 11 17 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.12
r37 10 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.27 $Y2=1.12
r38 4 16 68.5308 $w=2.11e-07 $l=4.82208e-07 $layer=POLY_cond $X=0.57 $Y=0.765
+ $X2=0.27 $Y2=1.12
r39 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.57 $Y=0.765 $X2=0.57
+ $Y2=0.445
r40 1 10 73.5404 $w=2.72e-07 $l=5.17373e-07 $layer=POLY_cond $X=0.5 $Y=1.875
+ $X2=0.27 $Y2=1.46
r41 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.5 $Y=1.875 $X2=0.5
+ $Y2=2.195
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_2%B 3 7 9 12 13
c38 13 0 1.49631e-19 $X=0.84 $Y=1.32
c39 12 0 1.94859e-19 $X=0.84 $Y=1.32
r40 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.32
+ $X2=0.84 $Y2=1.485
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.32
+ $X2=0.84 $Y2=1.155
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.84
+ $Y=1.32 $X2=0.84 $Y2=1.32
r43 9 13 4.5342 $w=3.03e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.277 $X2=0.84
+ $Y2=1.277
r44 7 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.93 $Y=2.195
+ $X2=0.93 $Y2=1.485
r45 3 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.93 $Y=0.445
+ $X2=0.93 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_2%A_46_47# 1 2 9 13 15 19 23 25 28 30 31 34 36
+ 37 40 43 45 46
c86 40 0 1.94859e-19 $X=1.35 $Y=1.385
c87 9 0 1.49631e-19 $X=1.455 $Y=0.655
r88 46 47 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.38 $Y=1.345
+ $X2=1.38 $Y2=1.27
r89 44 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.435
+ $X2=1.38 $Y2=1.6
r90 44 46 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.38 $Y=1.435 $X2=1.38
+ $Y2=1.345
r91 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.38
+ $Y=1.435 $X2=1.38 $Y2=1.435
r92 41 43 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=1.6
+ $X2=1.35 $Y2=1.435
r93 40 45 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.35 $Y=1.385
+ $X2=1.35 $Y2=1.27
r94 40 43 2.50531 $w=2.28e-07 $l=5e-08 $layer=LI1_cond $X=1.35 $Y=1.385 $X2=1.35
+ $Y2=1.435
r95 38 45 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.32 $Y=0.865
+ $X2=1.32 $Y2=1.27
r96 36 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.235 $Y=1.685
+ $X2=1.35 $Y2=1.6
r97 36 37 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.235 $Y=1.685
+ $X2=0.845 $Y2=1.685
r98 32 37 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.732 $Y=1.77
+ $X2=0.845 $Y2=1.685
r99 32 34 21.7684 $w=2.23e-07 $l=4.25e-07 $layer=LI1_cond $X=0.732 $Y=1.77
+ $X2=0.732 $Y2=2.195
r100 30 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.235 $Y=0.78
+ $X2=1.32 $Y2=0.865
r101 30 31 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.235 $Y=0.78
+ $X2=0.52 $Y2=0.78
r102 26 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.355 $Y=0.695
+ $X2=0.52 $Y2=0.78
r103 26 28 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.355 $Y=0.695
+ $X2=0.355 $Y2=0.445
r104 21 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=1.42
+ $X2=1.885 $Y2=1.345
r105 21 23 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=1.885 $Y=1.42
+ $X2=1.885 $Y2=2.465
r106 17 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=1.27
+ $X2=1.885 $Y2=1.345
r107 17 19 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.885 $Y=1.27
+ $X2=1.885 $Y2=0.655
r108 16 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.545 $Y=1.345
+ $X2=1.38 $Y2=1.345
r109 15 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.81 $Y=1.345
+ $X2=1.885 $Y2=1.345
r110 15 16 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=1.81 $Y=1.345
+ $X2=1.545 $Y2=1.345
r111 13 49 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=1.455 $Y=2.465
+ $X2=1.455 $Y2=1.6
r112 9 47 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.455 $Y=0.655
+ $X2=1.455 $Y2=1.27
r113 2 34 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.985 $X2=0.715 $Y2=2.195
r114 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.23
+ $Y=0.235 $X2=0.355 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_2%VPWR 1 2 3 10 12 16 20 22 26 28 33 42 46
r30 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 37 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 34 42 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.36 $Y=3.33
+ $X2=1.187 $Y2=3.33
r35 34 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.36 $Y=3.33 $X2=1.68
+ $Y2=3.33
r36 33 45 4.24382 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.192 $Y2=3.33
r37 33 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 32 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r39 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 29 39 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.225 $Y2=3.33
r41 29 31 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=3.33 $X2=0.72
+ $Y2=3.33
r42 28 42 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.187 $Y2=3.33
r43 28 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 26 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 22 25 39.9239 $w=2.78e-07 $l=9.7e-07 $layer=LI1_cond $X=2.125 $Y=1.98
+ $X2=2.125 $Y2=2.95
r48 20 45 3.11623 $w=2.8e-07 $l=1.13666e-07 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.192 $Y2=3.33
r49 20 25 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=2.95
r50 16 19 14.5308 $w=3.43e-07 $l=4.35e-07 $layer=LI1_cond $X=1.187 $Y=2.11
+ $X2=1.187 $Y2=2.545
r51 14 42 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.187 $Y=3.245
+ $X2=1.187 $Y2=3.33
r52 14 19 23.3829 $w=3.43e-07 $l=7e-07 $layer=LI1_cond $X=1.187 $Y=3.245
+ $X2=1.187 $Y2=2.545
r53 10 39 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.225 $Y2=3.33
r54 10 12 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.285 $Y2=2.195
r55 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.835 $X2=2.1 $Y2=2.95
r56 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.835 $X2=2.1 $Y2=1.98
r57 2 19 300 $w=1.7e-07 $l=6.67233e-07 $layer=licon1_PDIFF $count=2 $X=1.005
+ $Y=1.985 $X2=1.24 $Y2=2.545
r58 2 16 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.985 $X2=1.145 $Y2=2.11
r59 1 12 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.985 $X2=0.285 $Y2=2.195
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_2%X 1 2 9 13 14 15 16 32 34
r28 21 34 1.90052 $w=2.83e-07 $l=4.7e-08 $layer=LI1_cond $X=1.672 $Y=2.082
+ $X2=1.672 $Y2=2.035
r29 16 29 5.45894 $w=2.83e-07 $l=1.35e-07 $layer=LI1_cond $X=1.672 $Y=2.775
+ $X2=1.672 $Y2=2.91
r30 15 16 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.672 $Y=2.405
+ $X2=1.672 $Y2=2.775
r31 14 34 0.768295 $w=2.83e-07 $l=1.9e-08 $layer=LI1_cond $X=1.672 $Y=2.016
+ $X2=1.672 $Y2=2.035
r32 14 32 4.6303 $w=2.83e-07 $l=7.6e-08 $layer=LI1_cond $X=1.672 $Y=2.016
+ $X2=1.672 $Y2=1.94
r33 14 15 12.2927 $w=2.83e-07 $l=3.04e-07 $layer=LI1_cond $X=1.672 $Y=2.101
+ $X2=1.672 $Y2=2.405
r34 14 21 0.768295 $w=2.83e-07 $l=1.9e-08 $layer=LI1_cond $X=1.672 $Y=2.101
+ $X2=1.672 $Y2=2.082
r35 13 32 52.3737 $w=1.78e-07 $l=8.5e-07 $layer=LI1_cond $X=1.725 $Y=1.09
+ $X2=1.725 $Y2=1.94
r36 7 13 6.50835 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=1.695 $Y=0.97
+ $X2=1.695 $Y2=1.09
r37 7 9 26.4102 $w=2.38e-07 $l=5.5e-07 $layer=LI1_cond $X=1.695 $Y=0.97
+ $X2=1.695 $Y2=0.42
r38 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.835 $X2=1.67 $Y2=2.91
r39 2 14 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.835 $X2=1.67 $Y2=2.105
r40 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.53
+ $Y=0.235 $X2=1.67 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_2%VGND 1 2 9 11 13 15 17 22 28 32
r33 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r35 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r36 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=0 $X2=1.195
+ $Y2=0
r37 23 25 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.36 $Y=0 $X2=1.68
+ $Y2=0
r38 22 31 4.24382 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.192
+ $Y2=0
r39 22 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=1.68
+ $Y2=0
r40 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.195
+ $Y2=0
r42 17 19 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r43 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r44 15 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r45 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 11 31 3.11623 $w=2.8e-07 $l=1.13666e-07 $layer=LI1_cond $X=2.125 $Y=0.085
+ $X2=2.192 $Y2=0
r47 11 13 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.125 $Y=0.085
+ $X2=2.125 $Y2=0.38
r48 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0
r49 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0.4
r50 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.96
+ $Y=0.235 $X2=2.1 $Y2=0.38
r51 1 9 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.195 $Y2=0.4
.ends

