# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__xnor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 1.425000 1.825000 1.750000 ;
        RECT 1.655000 1.005000 2.635000 1.175000 ;
        RECT 1.655000 1.175000 1.825000 1.425000 ;
        RECT 2.465000 1.175000 2.635000 1.405000 ;
        RECT 2.465000 1.405000 3.135000 1.575000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.345000 2.285000 1.675000 ;
        RECT 2.115000 1.675000 2.285000 1.745000 ;
        RECT 2.115000 1.745000 4.500000 1.750000 ;
        RECT 2.115000 1.750000 3.475000 1.915000 ;
        RECT 3.305000 1.405000 4.500000 1.745000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.255800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.095000 2.260000 5.215000 2.430000 ;
        RECT 4.095000 2.430000 4.355000 2.635000 ;
        RECT 5.025000 1.775000 6.155000 1.945000 ;
        RECT 5.025000 1.945000 5.215000 2.260000 ;
        RECT 5.025000 2.430000 5.215000 3.075000 ;
        RECT 5.315000 0.595000 5.645000 1.065000 ;
        RECT 5.315000 1.065000 6.155000 1.235000 ;
        RECT 5.885000 1.235000 6.155000 1.775000 ;
        RECT 5.885000 1.945000 6.155000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.095000  0.255000 0.415000 0.735000 ;
      RECT 0.095000  0.735000 1.145000 0.905000 ;
      RECT 0.095000  0.905000 0.425000 1.095000 ;
      RECT 0.300000  1.815000 0.510000 2.270000 ;
      RECT 0.300000  2.270000 0.645000 3.245000 ;
      RECT 0.585000  0.085000 0.805000 0.565000 ;
      RECT 0.680000  1.075000 1.485000 1.245000 ;
      RECT 0.680000  1.245000 0.850000 1.920000 ;
      RECT 0.680000  1.920000 1.945000 2.085000 ;
      RECT 0.680000  2.085000 4.855000 2.090000 ;
      RECT 0.680000  2.090000 1.065000 2.100000 ;
      RECT 0.815000  2.100000 1.065000 3.075000 ;
      RECT 0.975000  0.255000 2.515000 0.445000 ;
      RECT 0.975000  0.445000 1.145000 0.735000 ;
      RECT 1.235000  2.260000 1.565000 3.245000 ;
      RECT 1.315000  0.615000 2.015000 0.815000 ;
      RECT 1.315000  0.815000 1.485000 1.075000 ;
      RECT 1.745000  2.090000 3.855000 2.255000 ;
      RECT 1.745000  2.255000 2.015000 3.075000 ;
      RECT 2.185000  0.445000 2.515000 0.835000 ;
      RECT 2.195000  2.435000 2.525000 3.245000 ;
      RECT 2.700000  2.435000 3.855000 2.605000 ;
      RECT 2.700000  2.605000 3.030000 3.075000 ;
      RECT 2.805000  0.300000 2.995000 1.065000 ;
      RECT 2.805000  1.065000 5.145000 1.235000 ;
      RECT 3.165000  0.085000 3.495000 0.895000 ;
      RECT 3.200000  2.775000 3.460000 3.245000 ;
      RECT 3.630000  2.605000 3.855000 2.895000 ;
      RECT 3.630000  2.895000 4.855000 3.065000 ;
      RECT 3.645000  1.920000 4.855000 2.085000 ;
      RECT 3.665000  0.300000 3.855000 1.065000 ;
      RECT 4.025000  0.085000 4.785000 0.895000 ;
      RECT 4.525000  2.600000 4.855000 2.895000 ;
      RECT 4.685000  1.405000 5.715000 1.605000 ;
      RECT 4.685000  1.605000 4.855000 1.920000 ;
      RECT 4.955000  0.255000 6.145000 0.425000 ;
      RECT 4.955000  0.425000 5.145000 1.065000 ;
      RECT 5.385000  2.115000 5.715000 3.245000 ;
      RECT 5.815000  0.425000 6.145000 0.895000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__xnor2_2
END LIBRARY
