* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
X0 a_52_367# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_304_237# S VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_304_237# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_29_73# a_304_237# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND S a_212_73# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_29_73# A0 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Y A1 a_236_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VPWR S a_52_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Y A1 a_212_73# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_236_367# a_304_237# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
