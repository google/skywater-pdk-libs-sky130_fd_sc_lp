* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4b_lp A B C D_N VGND VNB VPB VPWR Y
X0 a_31_409# D_N a_144_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_799_57# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Y C a_466_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_144_57# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_31_409# a_302_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y a_31_409# a_537_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VGND B a_641_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_537_409# C a_635_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_641_57# B Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_31_409# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_635_409# B a_733_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 Y A a_799_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_733_409# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_466_57# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_302_57# a_31_409# Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
