* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_781_51# a_823_25# a_432_109# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_823_25# a_1109_21# a_1204_459# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_1204_459# a_1246_339# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 VPWR GATE a_1109_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VGND a_432_109# a_1067_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_432_109# a_981_503# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR D a_1246_339# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VGND a_80_21# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_432_109# a_823_25# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_981_503# a_1023_405# a_823_25# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VGND a_432_109# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 Q_N a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VPWR RESET_B a_432_109# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 Q a_432_109# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VPWR a_80_21# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND RESET_B a_781_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_1023_405# a_1109_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_432_109# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VGND GATE a_1109_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_80_21# a_432_109# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_1225_119# a_1246_339# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1023_405# a_1109_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 Q a_432_109# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_823_25# a_1023_405# a_1225_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_80_21# a_432_109# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND D a_1246_339# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 Q_N a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_1067_119# a_1109_21# a_823_25# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
