* File: sky130_fd_sc_lp__dfsbp_lp.pxi.spice
* Created: Wed Sep  2 09:44:14 2020
* 
x_PM_SKY130_FD_SC_LP__DFSBP_LP%D N_D_c_280_n N_D_M1019_g N_D_M1002_g N_D_c_281_n
+ N_D_M1010_g N_D_c_282_n D D N_D_c_283_n N_D_c_284_n N_D_c_285_n
+ PM_SKY130_FD_SC_LP__DFSBP_LP%D
x_PM_SKY130_FD_SC_LP__DFSBP_LP%CLK N_CLK_M1001_g N_CLK_c_315_n N_CLK_M1036_g
+ N_CLK_c_316_n N_CLK_c_317_n N_CLK_M1024_g N_CLK_c_318_n CLK N_CLK_c_320_n
+ N_CLK_c_321_n PM_SKY130_FD_SC_LP__DFSBP_LP%CLK
x_PM_SKY130_FD_SC_LP__DFSBP_LP%A_476_409# N_A_476_409#_M1021_d
+ N_A_476_409#_M1026_d N_A_476_409#_M1005_g N_A_476_409#_M1017_g
+ N_A_476_409#_M1009_g N_A_476_409#_M1015_g N_A_476_409#_c_386_n
+ N_A_476_409#_c_387_n N_A_476_409#_c_388_n N_A_476_409#_c_374_n
+ N_A_476_409#_c_389_n N_A_476_409#_c_375_n N_A_476_409#_c_376_n
+ N_A_476_409#_c_377_n N_A_476_409#_c_402_p N_A_476_409#_c_403_p
+ N_A_476_409#_c_397_p N_A_476_409#_c_420_p N_A_476_409#_c_378_n
+ N_A_476_409#_c_379_n N_A_476_409#_c_394_n N_A_476_409#_c_380_n
+ N_A_476_409#_c_381_n N_A_476_409#_c_409_p N_A_476_409#_c_382_n
+ N_A_476_409#_c_383_n PM_SKY130_FD_SC_LP__DFSBP_LP%A_476_409#
x_PM_SKY130_FD_SC_LP__DFSBP_LP%A_946_99# N_A_946_99#_M1034_s N_A_946_99#_M1003_d
+ N_A_946_99#_M1008_g N_A_946_99#_c_582_n N_A_946_99#_M1032_g
+ N_A_946_99#_c_583_n N_A_946_99#_c_589_n N_A_946_99#_c_584_n
+ N_A_946_99#_c_590_n N_A_946_99#_c_591_n N_A_946_99#_c_585_n
+ N_A_946_99#_c_586_n PM_SKY130_FD_SC_LP__DFSBP_LP%A_946_99#
x_PM_SKY130_FD_SC_LP__DFSBP_LP%A_712_419# N_A_712_419#_M1020_d
+ N_A_712_419#_M1005_d N_A_712_419#_M1003_g N_A_712_419#_M1034_g
+ N_A_712_419#_M1018_g N_A_712_419#_M1029_g N_A_712_419#_c_661_n
+ N_A_712_419#_c_662_n N_A_712_419#_c_683_n N_A_712_419#_c_699_n
+ N_A_712_419#_c_663_n N_A_712_419#_c_684_n N_A_712_419#_c_685_n
+ N_A_712_419#_c_664_n N_A_712_419#_c_665_n N_A_712_419#_c_666_n
+ N_A_712_419#_c_667_n N_A_712_419#_c_668_n N_A_712_419#_c_669_n
+ N_A_712_419#_c_670_n N_A_712_419#_c_671_n N_A_712_419#_c_672_n
+ N_A_712_419#_c_673_n N_A_712_419#_c_674_n N_A_712_419#_c_675_n
+ N_A_712_419#_c_676_n N_A_712_419#_c_767_n N_A_712_419#_c_677_n
+ N_A_712_419#_c_678_n N_A_712_419#_c_679_n
+ PM_SKY130_FD_SC_LP__DFSBP_LP%A_712_419#
x_PM_SKY130_FD_SC_LP__DFSBP_LP%SET_B N_SET_B_M1027_g N_SET_B_M1022_g
+ N_SET_B_c_849_n N_SET_B_M1037_g N_SET_B_c_850_n N_SET_B_c_851_n
+ N_SET_B_M1013_g N_SET_B_c_852_n N_SET_B_c_853_n N_SET_B_c_861_n
+ N_SET_B_c_862_n N_SET_B_c_875_n SET_B N_SET_B_c_854_n N_SET_B_c_855_n
+ N_SET_B_c_856_n N_SET_B_c_857_n PM_SKY130_FD_SC_LP__DFSBP_LP%SET_B
x_PM_SKY130_FD_SC_LP__DFSBP_LP%A_263_409# N_A_263_409#_M1036_s
+ N_A_263_409#_M1001_s N_A_263_409#_M1026_g N_A_263_409#_c_987_n
+ N_A_263_409#_M1028_g N_A_263_409#_c_988_n N_A_263_409#_c_989_n
+ N_A_263_409#_c_990_n N_A_263_409#_M1021_g N_A_263_409#_c_991_n
+ N_A_263_409#_c_992_n N_A_263_409#_c_993_n N_A_263_409#_M1020_g
+ N_A_263_409#_c_1006_n N_A_263_409#_c_1007_n N_A_263_409#_c_995_n
+ N_A_263_409#_c_996_n N_A_263_409#_c_1008_n N_A_263_409#_M1016_g
+ N_A_263_409#_c_1009_n N_A_263_409#_M1038_g N_A_263_409#_c_1010_n
+ N_A_263_409#_c_1011_n N_A_263_409#_M1000_g N_A_263_409#_c_998_n
+ N_A_263_409#_c_999_n N_A_263_409#_c_1000_n N_A_263_409#_c_1001_n
+ N_A_263_409#_c_1014_n N_A_263_409#_c_1015_n N_A_263_409#_c_1002_n
+ N_A_263_409#_c_1017_n N_A_263_409#_c_1003_n
+ PM_SKY130_FD_SC_LP__DFSBP_LP%A_263_409#
x_PM_SKY130_FD_SC_LP__DFSBP_LP%A_1686_40# N_A_1686_40#_M1006_s
+ N_A_1686_40#_M1007_s N_A_1686_40#_M1039_g N_A_1686_40#_c_1191_n
+ N_A_1686_40#_c_1192_n N_A_1686_40#_M1033_g N_A_1686_40#_c_1193_n
+ N_A_1686_40#_c_1194_n N_A_1686_40#_c_1195_n N_A_1686_40#_c_1196_n
+ N_A_1686_40#_c_1197_n N_A_1686_40#_c_1198_n N_A_1686_40#_c_1199_n
+ N_A_1686_40#_c_1200_n N_A_1686_40#_c_1201_n
+ PM_SKY130_FD_SC_LP__DFSBP_LP%A_1686_40#
x_PM_SKY130_FD_SC_LP__DFSBP_LP%A_1519_125# N_A_1519_125#_M1009_d
+ N_A_1519_125#_M1038_d N_A_1519_125#_M1013_d N_A_1519_125#_c_1287_n
+ N_A_1519_125#_M1006_g N_A_1519_125#_c_1288_n N_A_1519_125#_c_1289_n
+ N_A_1519_125#_c_1290_n N_A_1519_125#_M1035_g N_A_1519_125#_c_1291_n
+ N_A_1519_125#_M1007_g N_A_1519_125#_c_1292_n N_A_1519_125#_M1011_g
+ N_A_1519_125#_c_1293_n N_A_1519_125#_c_1294_n N_A_1519_125#_c_1295_n
+ N_A_1519_125#_c_1296_n N_A_1519_125#_M1012_g N_A_1519_125#_M1014_g
+ N_A_1519_125#_c_1298_n N_A_1519_125#_c_1299_n N_A_1519_125#_c_1300_n
+ N_A_1519_125#_c_1301_n N_A_1519_125#_M1023_g N_A_1519_125#_M1004_g
+ N_A_1519_125#_c_1303_n N_A_1519_125#_M1025_g N_A_1519_125#_c_1304_n
+ N_A_1519_125#_c_1305_n N_A_1519_125#_c_1306_n N_A_1519_125#_c_1324_n
+ N_A_1519_125#_c_1307_n N_A_1519_125#_c_1308_n N_A_1519_125#_c_1331_n
+ N_A_1519_125#_c_1309_n N_A_1519_125#_c_1351_n N_A_1519_125#_c_1316_n
+ N_A_1519_125#_c_1317_n N_A_1519_125#_c_1318_n N_A_1519_125#_c_1319_n
+ N_A_1519_125#_c_1310_n N_A_1519_125#_c_1320_n N_A_1519_125#_c_1321_n
+ N_A_1519_125#_c_1401_n N_A_1519_125#_c_1322_n N_A_1519_125#_c_1311_n
+ PM_SKY130_FD_SC_LP__DFSBP_LP%A_1519_125#
x_PM_SKY130_FD_SC_LP__DFSBP_LP%A_2383_57# N_A_2383_57#_M1023_s
+ N_A_2383_57#_M1004_s N_A_2383_57#_M1040_g N_A_2383_57#_M1030_g
+ N_A_2383_57#_M1031_g N_A_2383_57#_c_1509_n N_A_2383_57#_c_1510_n
+ N_A_2383_57#_c_1511_n N_A_2383_57#_c_1519_n N_A_2383_57#_c_1512_n
+ N_A_2383_57#_c_1513_n N_A_2383_57#_c_1514_n N_A_2383_57#_c_1515_n
+ N_A_2383_57#_c_1516_n PM_SKY130_FD_SC_LP__DFSBP_LP%A_2383_57#
x_PM_SKY130_FD_SC_LP__DFSBP_LP%VPWR N_VPWR_M1002_s N_VPWR_M1001_d N_VPWR_M1032_d
+ N_VPWR_M1027_d N_VPWR_M1033_d N_VPWR_M1007_d N_VPWR_M1004_d N_VPWR_c_1575_n
+ N_VPWR_c_1576_n N_VPWR_c_1577_n N_VPWR_c_1578_n N_VPWR_c_1579_n
+ N_VPWR_c_1580_n N_VPWR_c_1581_n N_VPWR_c_1582_n N_VPWR_c_1583_n
+ N_VPWR_c_1584_n N_VPWR_c_1585_n N_VPWR_c_1586_n VPWR N_VPWR_c_1587_n
+ N_VPWR_c_1588_n N_VPWR_c_1589_n N_VPWR_c_1590_n N_VPWR_c_1591_n
+ N_VPWR_c_1574_n N_VPWR_c_1593_n N_VPWR_c_1594_n N_VPWR_c_1595_n
+ N_VPWR_c_1596_n PM_SKY130_FD_SC_LP__DFSBP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DFSBP_LP%A_145_409# N_A_145_409#_M1010_d
+ N_A_145_409#_M1020_s N_A_145_409#_M1002_d N_A_145_409#_M1005_s
+ N_A_145_409#_c_1727_n N_A_145_409#_c_1728_n N_A_145_409#_c_1715_n
+ N_A_145_409#_c_1716_n N_A_145_409#_c_1717_n N_A_145_409#_c_1718_n
+ N_A_145_409#_c_1719_n N_A_145_409#_c_1720_n N_A_145_409#_c_1721_n
+ N_A_145_409#_c_1722_n N_A_145_409#_c_1730_n N_A_145_409#_c_1731_n
+ N_A_145_409#_c_1732_n N_A_145_409#_c_1723_n N_A_145_409#_c_1724_n
+ N_A_145_409#_c_1725_n N_A_145_409#_c_1726_n
+ PM_SKY130_FD_SC_LP__DFSBP_LP%A_145_409#
x_PM_SKY130_FD_SC_LP__DFSBP_LP%Q_N N_Q_N_M1012_d N_Q_N_M1014_d N_Q_N_c_1847_n
+ N_Q_N_c_1844_n Q_N Q_N N_Q_N_c_1846_n PM_SKY130_FD_SC_LP__DFSBP_LP%Q_N
x_PM_SKY130_FD_SC_LP__DFSBP_LP%Q N_Q_M1031_d N_Q_M1030_d N_Q_c_1883_n Q Q Q
+ N_Q_c_1886_n N_Q_c_1884_n PM_SKY130_FD_SC_LP__DFSBP_LP%Q
x_PM_SKY130_FD_SC_LP__DFSBP_LP%VGND N_VGND_M1019_s N_VGND_M1024_d N_VGND_M1008_d
+ N_VGND_M1022_d N_VGND_M1037_d N_VGND_M1035_d N_VGND_M1025_d N_VGND_c_1906_n
+ N_VGND_c_1907_n N_VGND_c_1908_n N_VGND_c_1909_n N_VGND_c_1910_n
+ N_VGND_c_1911_n N_VGND_c_1912_n N_VGND_c_1913_n N_VGND_c_1914_n
+ N_VGND_c_1915_n N_VGND_c_1916_n N_VGND_c_1917_n N_VGND_c_1918_n VGND
+ N_VGND_c_1919_n N_VGND_c_1920_n N_VGND_c_1921_n N_VGND_c_1922_n
+ N_VGND_c_1923_n N_VGND_c_1924_n N_VGND_c_1925_n N_VGND_c_1926_n
+ N_VGND_c_1927_n PM_SKY130_FD_SC_LP__DFSBP_LP%VGND
cc_1 VNB N_D_c_280_n 0.0175114f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.78
cc_2 VNB N_D_c_281_n 0.0174678f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.78
cc_3 VNB N_D_c_282_n 0.0304469f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.855
cc_4 VNB N_D_c_283_n 0.0634179f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_5 VNB N_D_c_284_n 0.0245402f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_6 VNB N_D_c_285_n 0.0194264f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.11
cc_7 VNB N_CLK_c_315_n 0.0156366f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.11
cc_8 VNB N_CLK_c_316_n 0.0182382f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.78
cc_9 VNB N_CLK_c_317_n 0.0135295f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.495
cc_10 VNB N_CLK_c_318_n 0.00702308f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=0.855
cc_11 VNB CLK 0.00222853f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.855
cc_12 VNB N_CLK_c_320_n 0.0218013f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_CLK_c_321_n 0.0168058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_476_409#_M1017_g 0.0255674f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.855
cc_15 VNB N_A_476_409#_M1009_g 0.0240529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_476_409#_c_374_n 0.00843919f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.665
cc_17 VNB N_A_476_409#_c_375_n 0.00690406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_476_409#_c_376_n 0.00952385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_476_409#_c_377_n 0.0234764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_476_409#_c_378_n 4.47893e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_476_409#_c_379_n 0.0129681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_476_409#_c_380_n 0.00950533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_476_409#_c_381_n 0.0178381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_476_409#_c_382_n 0.0303001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_476_409#_c_383_n 0.00388401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_946_99#_M1008_g 0.0220347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_946_99#_c_582_n 0.0582162f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.495
cc_28 VNB N_A_946_99#_c_583_n 0.00315929f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=0.855
cc_29 VNB N_A_946_99#_c_584_n 0.0170838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_946_99#_c_585_n 0.00688544f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_31 VNB N_A_946_99#_c_586_n 0.0116299f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_32 VNB N_A_712_419#_M1034_g 0.0204585f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=0.855
cc_33 VNB N_A_712_419#_M1029_g 0.0205744f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_34 VNB N_A_712_419#_c_661_n 0.025845f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.275
cc_35 VNB N_A_712_419#_c_662_n 0.0169648f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_36 VNB N_A_712_419#_c_663_n 0.00436449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_712_419#_c_664_n 0.00652238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_712_419#_c_665_n 0.00252665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_712_419#_c_666_n 0.00454688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_712_419#_c_667_n 0.00704227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_712_419#_c_668_n 0.012364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_712_419#_c_669_n 0.025229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_712_419#_c_670_n 0.00348498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_712_419#_c_671_n 0.0018543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_712_419#_c_672_n 0.0102377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_712_419#_c_673_n 0.00314283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_712_419#_c_674_n 0.00967025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_712_419#_c_675_n 0.00934316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_712_419#_c_676_n 0.00513594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_712_419#_c_677_n 0.00309778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_712_419#_c_678_n 0.0145769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_712_419#_c_679_n 0.0129404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_SET_B_M1022_g 0.0399696f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.545
cc_54 VNB N_SET_B_c_849_n 0.0187067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_SET_B_c_850_n 0.0519874f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.495
cc_56 VNB N_SET_B_c_851_n 0.00674719f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.855
cc_57 VNB N_SET_B_c_852_n 0.0194997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_SET_B_c_853_n 0.0161115f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.275
cc_59 VNB N_SET_B_c_854_n 0.0165464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_SET_B_c_855_n 0.00583734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_SET_B_c_856_n 0.0011472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_SET_B_c_857_n 0.0121328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_263_409#_c_987_n 0.0135295f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.495
cc_64 VNB N_A_263_409#_c_988_n 0.0243533f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=0.855
cc_65 VNB N_A_263_409#_c_989_n 0.00901312f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.855
cc_66 VNB N_A_263_409#_c_990_n 0.0156237f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_67 VNB N_A_263_409#_c_991_n 0.0483904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_263_409#_c_992_n 0.0152186f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_69 VNB N_A_263_409#_c_993_n 0.0228024f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_70 VNB N_A_263_409#_M1020_g 0.0218556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_263_409#_c_995_n 0.305402f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_72 VNB N_A_263_409#_c_996_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_263_409#_M1000_g 0.0576265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_263_409#_c_998_n 0.0046367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_263_409#_c_999_n 0.0100371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_263_409#_c_1000_n 0.0175557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_263_409#_c_1001_n 0.012491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_263_409#_c_1002_n 0.0034243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_263_409#_c_1003_n 0.0189167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1686_40#_M1039_g 0.0373462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1686_40#_c_1191_n 0.0373289f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.495
cc_82 VNB N_A_1686_40#_c_1192_n 0.00835867f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.495
cc_83 VNB N_A_1686_40#_c_1193_n 0.00120563f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_84 VNB N_A_1686_40#_c_1194_n 0.00234083f $X=-0.19 $Y=-0.245 $X2=0.472
+ $Y2=1.275
cc_85 VNB N_A_1686_40#_c_1195_n 0.0260001f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.275
cc_86 VNB N_A_1686_40#_c_1196_n 0.007392f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.11
cc_87 VNB N_A_1686_40#_c_1197_n 8.22949e-19 $X=-0.19 $Y=-0.245 $X2=0.472
+ $Y2=1.78
cc_88 VNB N_A_1686_40#_c_1198_n 0.0127228f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.295
cc_89 VNB N_A_1686_40#_c_1199_n 0.0164805f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.665
cc_90 VNB N_A_1686_40#_c_1200_n 0.00942875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1686_40#_c_1201_n 0.00664779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1519_125#_c_1287_n 0.0175304f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.78
cc_93 VNB N_A_1519_125#_c_1288_n 0.0101801f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=0.855
cc_94 VNB N_A_1519_125#_c_1289_n 0.00937291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1519_125#_c_1290_n 0.0136552f $X=-0.19 $Y=-0.245 $X2=0.562
+ $Y2=0.855
cc_96 VNB N_A_1519_125#_c_1291_n 0.0160628f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_97 VNB N_A_1519_125#_c_1292_n 0.0136573f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.275
cc_98 VNB N_A_1519_125#_c_1293_n 0.00747072f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.275
cc_99 VNB N_A_1519_125#_c_1294_n 0.007351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1519_125#_c_1295_n 0.00977986f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.295
cc_101 VNB N_A_1519_125#_c_1296_n 0.0171659f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.665
cc_102 VNB N_A_1519_125#_M1014_g 0.0237112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1519_125#_c_1298_n 0.0134123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1519_125#_c_1299_n 0.0386698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1519_125#_c_1300_n 0.0186068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1519_125#_c_1301_n 0.0174911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1519_125#_M1004_g 0.0501546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1519_125#_c_1303_n 0.0137559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1519_125#_c_1304_n 0.00494546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1519_125#_c_1305_n 0.00838945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1519_125#_c_1306_n 0.0176414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1519_125#_c_1307_n 0.0174792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1519_125#_c_1308_n 0.00718231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1519_125#_c_1309_n 0.00507043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1519_125#_c_1310_n 0.00396923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_1519_125#_c_1311_n 0.0607429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2383_57#_M1040_g 0.0241564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2383_57#_M1031_g 0.0293965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2383_57#_c_1509_n 0.0256228f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.275
cc_120 VNB N_A_2383_57#_c_1510_n 0.0123107f $X=-0.19 $Y=-0.245 $X2=0.472
+ $Y2=1.78
cc_121 VNB N_A_2383_57#_c_1511_n 0.0132686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2383_57#_c_1512_n 0.0114987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_2383_57#_c_1513_n 0.00121962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2383_57#_c_1514_n 0.0285181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2383_57#_c_1515_n 0.00849853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_2383_57#_c_1516_n 0.0074766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VPWR_c_1574_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_145_409#_c_1715_n 0.0213108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_145_409#_c_1716_n 0.00159743f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.275
cc_130 VNB N_A_145_409#_c_1717_n 0.00975871f $X=-0.19 $Y=-0.245 $X2=0.472
+ $Y2=1.11
cc_131 VNB N_A_145_409#_c_1718_n 0.00746485f $X=-0.19 $Y=-0.245 $X2=0.472
+ $Y2=1.78
cc_132 VNB N_A_145_409#_c_1719_n 0.00159816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_145_409#_c_1720_n 0.0030969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_145_409#_c_1721_n 0.0204674f $X=-0.19 $Y=-0.245 $X2=0.337
+ $Y2=1.665
cc_135 VNB N_A_145_409#_c_1722_n 0.00291864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_145_409#_c_1723_n 0.00787639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_145_409#_c_1724_n 0.0167037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_145_409#_c_1725_n 0.0140178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_145_409#_c_1726_n 5.74534e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_Q_N_c_1844_n 0.00976104f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.855
cc_141 VNB Q_N 0.010094f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_142 VNB N_Q_N_c_1846_n 0.00445616f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_143 VNB N_Q_c_1883_n 0.0251105f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.78
cc_144 VNB N_Q_c_1884_n 0.0449413f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_145 VNB N_VGND_c_1906_n 0.0107448f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.275
cc_146 VNB N_VGND_c_1907_n 0.0265531f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_147 VNB N_VGND_c_1908_n 0.0132052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_1909_n 0.0105502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_1910_n 0.016709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_1911_n 0.0125499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_1912_n 0.00656177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_1913_n 0.0495856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_1914_n 0.0131801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_1915_n 0.0469158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_1916_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_1917_n 0.0557136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_1918_n 0.00585462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_1919_n 0.0645969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_1920_n 0.0379159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_1921_n 0.0366067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_1922_n 0.0271986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_1923_n 0.741253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_1924_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_1925_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_1926_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_1927_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VPB N_D_M1002_g 0.0458742f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.545
cc_168 VPB N_D_c_283_n 0.0206452f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_169 VPB N_D_c_284_n 0.00989638f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_170 VPB N_CLK_M1001_g 0.0367128f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.495
cc_171 VPB CLK 7.36937e-19 $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.855
cc_172 VPB N_CLK_c_320_n 0.0118764f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_173 VPB N_A_476_409#_M1005_g 0.0414125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_476_409#_M1015_g 0.0266119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_476_409#_c_386_n 0.00725725f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.11
cc_176 VPB N_A_476_409#_c_387_n 0.0157333f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.275
cc_177 VPB N_A_476_409#_c_388_n 0.00246318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_476_409#_c_389_n 0.00336316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_476_409#_c_375_n 0.00375693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_476_409#_c_376_n 0.00972083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_476_409#_c_377_n 0.00548403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_476_409#_c_378_n 0.00836007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_476_409#_c_394_n 2.8107e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_476_409#_c_380_n 0.0217105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_476_409#_c_381_n 0.0104571f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_946_99#_c_582_n 0.0364222f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.495
cc_187 VPB N_A_946_99#_M1032_g 0.0316319f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.855
cc_188 VPB N_A_946_99#_c_589_n 0.00332961f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.855
cc_189 VPB N_A_946_99#_c_590_n 3.51419e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_190 VPB N_A_946_99#_c_591_n 0.0114334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_712_419#_M1003_g 0.0316395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_712_419#_M1018_g 0.0273769f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_193 VPB N_A_712_419#_c_662_n 0.00718046f $X=-0.19 $Y=1.655 $X2=0.337
+ $Y2=1.665
cc_194 VPB N_A_712_419#_c_683_n 0.0145467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_712_419#_c_684_n 0.00697694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_712_419#_c_685_n 0.00238935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_712_419#_c_666_n 0.00640603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_712_419#_c_671_n 0.00397103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_712_419#_c_672_n 0.0160659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_712_419#_c_677_n 9.02542e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_SET_B_M1027_g 0.026945f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.495
cc_202 VPB N_SET_B_M1013_g 0.0308779f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.855
cc_203 VPB N_SET_B_c_853_n 0.00819959f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.275
cc_204 VPB N_SET_B_c_861_n 0.0153854f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_205 VPB N_SET_B_c_862_n 0.0242791f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_206 VPB SET_B 0.00290381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_SET_B_c_855_n 0.00411011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_SET_B_c_856_n 0.00200631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_SET_B_c_857_n 0.0288497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_263_409#_M1026_g 0.0293306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_263_409#_c_993_n 0.0140979f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_212 VPB N_A_263_409#_c_1006_n 0.0244652f $X=-0.19 $Y=1.655 $X2=0.337
+ $Y2=1.295
cc_213 VPB N_A_263_409#_c_1007_n 0.0108148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_263_409#_c_1008_n 0.0224979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_263_409#_c_1009_n 0.0212961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_263_409#_c_1010_n 0.0283612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_263_409#_c_1011_n 0.00935016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_263_409#_M1000_g 0.0101541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_263_409#_c_1001_n 0.00616039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_263_409#_c_1014_n 0.0134196f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_263_409#_c_1015_n 0.00929625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_263_409#_c_1002_n 7.01084e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_263_409#_c_1017_n 0.00986418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_263_409#_c_1003_n 0.0305389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1686_40#_M1033_g 0.0289122f $X=-0.19 $Y=1.655 $X2=0.562 $Y2=0.855
cc_226 VPB N_A_1686_40#_c_1193_n 0.0253082f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_227 VPB N_A_1686_40#_c_1194_n 0.0024701f $X=-0.19 $Y=1.655 $X2=0.472
+ $Y2=1.275
cc_228 VPB N_A_1686_40#_c_1200_n 0.0117268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_1519_125#_M1007_g 0.0296186f $X=-0.19 $Y=1.655 $X2=0.472
+ $Y2=1.275
cc_230 VPB N_A_1519_125#_M1014_g 0.0451827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_1519_125#_M1004_g 0.0316849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_1519_125#_c_1309_n 0.00354889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_1519_125#_c_1316_n 0.00256112f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_1519_125#_c_1317_n 0.00404091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_1519_125#_c_1318_n 0.014292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_1519_125#_c_1319_n 3.42419e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_1519_125#_c_1320_n 0.00175974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_1519_125#_c_1321_n 0.0029268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_1519_125#_c_1322_n 0.006464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_1519_125#_c_1311_n 0.0349895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_2383_57#_M1030_g 0.0343439f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.855
cc_242 VPB N_A_2383_57#_c_1510_n 0.00266792f $X=-0.19 $Y=1.655 $X2=0.472
+ $Y2=1.78
cc_243 VPB N_A_2383_57#_c_1519_n 0.0165762f $X=-0.19 $Y=1.655 $X2=0.337
+ $Y2=1.665
cc_244 VPB N_A_2383_57#_c_1512_n 0.00348674f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1575_n 0.0131113f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.275
cc_246 VPB N_VPWR_c_1576_n 0.0465021f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_247 VPB N_VPWR_c_1577_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1578_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1579_n 0.00487982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1580_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1581_n 0.00452326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1582_n 0.0139381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1583_n 0.0338291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1584_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1585_n 0.0324567f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1586_n 0.00631504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1587_n 0.066177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1588_n 0.0653177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1589_n 0.043549f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1590_n 0.0353069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1591_n 0.0270929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1574_n 0.106202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1593_n 0.00510188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1594_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1595_n 0.00428995f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1596_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_145_409#_c_1727_n 0.00694835f $X=-0.19 $Y=1.655 $X2=0.562
+ $Y2=0.855
cc_268 VPB N_A_145_409#_c_1728_n 0.00960744f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_145_409#_c_1720_n 0.003636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_145_409#_c_1730_n 0.0173148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_145_409#_c_1731_n 0.00617618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_145_409#_c_1732_n 0.00723729f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_145_409#_c_1724_n 0.00796123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_Q_N_c_1847_n 0.0148801f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.495
cc_275 VPB Q_N 0.00151544f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_276 VPB Q 0.043146f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_Q_c_1886_n 0.0282671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_Q_c_1884_n 0.00985254f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.295
cc_279 N_D_c_281_n N_A_263_409#_c_1000_n 0.00119574f $X=0.835 $Y=0.78 $X2=0
+ $Y2=0
cc_280 N_D_M1002_g N_A_263_409#_c_1014_n 0.00152794f $X=0.6 $Y=2.545 $X2=0 $Y2=0
cc_281 N_D_M1002_g N_A_263_409#_c_1017_n 2.35528e-19 $X=0.6 $Y=2.545 $X2=0 $Y2=0
cc_282 N_D_M1002_g N_VPWR_c_1576_n 0.0250417f $X=0.6 $Y=2.545 $X2=0 $Y2=0
cc_283 N_D_c_283_n N_VPWR_c_1576_n 0.00191238f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_284 N_D_c_284_n N_VPWR_c_1576_n 0.0223028f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_285 N_D_M1002_g N_VPWR_c_1583_n 0.00769046f $X=0.6 $Y=2.545 $X2=0 $Y2=0
cc_286 N_D_M1002_g N_VPWR_c_1574_n 0.0143431f $X=0.6 $Y=2.545 $X2=0 $Y2=0
cc_287 N_D_M1002_g N_A_145_409#_c_1727_n 0.00451956f $X=0.6 $Y=2.545 $X2=0 $Y2=0
cc_288 N_D_M1002_g N_A_145_409#_c_1728_n 0.015872f $X=0.6 $Y=2.545 $X2=0 $Y2=0
cc_289 N_D_c_281_n N_A_145_409#_c_1724_n 0.00184816f $X=0.835 $Y=0.78 $X2=0
+ $Y2=0
cc_290 N_D_c_282_n N_A_145_409#_c_1724_n 0.0106456f $X=0.835 $Y=0.855 $X2=0
+ $Y2=0
cc_291 N_D_c_284_n N_A_145_409#_c_1724_n 0.0327571f $X=0.385 $Y=1.275 $X2=0
+ $Y2=0
cc_292 N_D_c_285_n N_A_145_409#_c_1724_n 0.0343919f $X=0.472 $Y=1.11 $X2=0 $Y2=0
cc_293 N_D_c_280_n N_A_145_409#_c_1725_n 0.00158738f $X=0.475 $Y=0.78 $X2=0
+ $Y2=0
cc_294 N_D_c_281_n N_A_145_409#_c_1725_n 0.00967975f $X=0.835 $Y=0.78 $X2=0
+ $Y2=0
cc_295 N_D_c_280_n N_VGND_c_1907_n 0.0140511f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_296 N_D_c_281_n N_VGND_c_1907_n 0.00209399f $X=0.835 $Y=0.78 $X2=0 $Y2=0
cc_297 N_D_c_283_n N_VGND_c_1907_n 0.0012686f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_298 N_D_c_284_n N_VGND_c_1907_n 0.014708f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_299 N_D_c_280_n N_VGND_c_1915_n 0.00445056f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_300 N_D_c_281_n N_VGND_c_1915_n 0.00467918f $X=0.835 $Y=0.78 $X2=0 $Y2=0
cc_301 N_D_c_282_n N_VGND_c_1915_n 5.84996e-19 $X=0.835 $Y=0.855 $X2=0 $Y2=0
cc_302 N_D_c_280_n N_VGND_c_1923_n 0.00796275f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_303 N_D_c_281_n N_VGND_c_1923_n 0.00937674f $X=0.835 $Y=0.78 $X2=0 $Y2=0
cc_304 N_D_c_282_n N_VGND_c_1923_n 7.94744e-19 $X=0.835 $Y=0.855 $X2=0 $Y2=0
cc_305 N_CLK_c_317_n N_A_263_409#_c_987_n 0.00851747f $X=2.15 $Y=1.06 $X2=0
+ $Y2=0
cc_306 CLK N_A_263_409#_c_988_n 5.14737e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_307 N_CLK_c_320_n N_A_263_409#_c_988_n 0.00222567f $X=1.725 $Y=1.615 $X2=0
+ $Y2=0
cc_308 N_CLK_c_321_n N_A_263_409#_c_988_n 0.00488548f $X=1.725 $Y=1.45 $X2=0
+ $Y2=0
cc_309 N_CLK_c_316_n N_A_263_409#_c_998_n 0.00851747f $X=2.075 $Y=1.135 $X2=0
+ $Y2=0
cc_310 N_CLK_c_315_n N_A_263_409#_c_1000_n 0.00644031f $X=1.79 $Y=1.06 $X2=0
+ $Y2=0
cc_311 N_CLK_c_317_n N_A_263_409#_c_1000_n 3.49297e-19 $X=2.15 $Y=1.06 $X2=0
+ $Y2=0
cc_312 N_CLK_c_318_n N_A_263_409#_c_1000_n 0.00114563f $X=1.79 $Y=1.135 $X2=0
+ $Y2=0
cc_313 CLK N_A_263_409#_c_1000_n 0.0080165f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_314 N_CLK_c_320_n N_A_263_409#_c_1000_n 0.00102834f $X=1.725 $Y=1.615 $X2=0
+ $Y2=0
cc_315 N_CLK_M1001_g N_A_263_409#_c_1001_n 0.00445693f $X=1.725 $Y=2.545 $X2=0
+ $Y2=0
cc_316 N_CLK_c_318_n N_A_263_409#_c_1001_n 0.0082313f $X=1.79 $Y=1.135 $X2=0
+ $Y2=0
cc_317 CLK N_A_263_409#_c_1001_n 0.0237562f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_318 N_CLK_c_320_n N_A_263_409#_c_1001_n 0.00735127f $X=1.725 $Y=1.615 $X2=0
+ $Y2=0
cc_319 N_CLK_M1001_g N_A_263_409#_c_1014_n 0.017065f $X=1.725 $Y=2.545 $X2=0
+ $Y2=0
cc_320 N_CLK_M1001_g N_A_263_409#_c_1015_n 0.0178513f $X=1.725 $Y=2.545 $X2=0
+ $Y2=0
cc_321 CLK N_A_263_409#_c_1015_n 0.0182122f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_322 N_CLK_c_320_n N_A_263_409#_c_1015_n 2.70163e-19 $X=1.725 $Y=1.615 $X2=0
+ $Y2=0
cc_323 N_CLK_M1001_g N_A_263_409#_c_1002_n 0.00117819f $X=1.725 $Y=2.545 $X2=0
+ $Y2=0
cc_324 CLK N_A_263_409#_c_1002_n 0.0128184f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_325 N_CLK_c_320_n N_A_263_409#_c_1002_n 8.28332e-19 $X=1.725 $Y=1.615 $X2=0
+ $Y2=0
cc_326 N_CLK_M1001_g N_A_263_409#_c_1017_n 0.00255958f $X=1.725 $Y=2.545 $X2=0
+ $Y2=0
cc_327 CLK N_A_263_409#_c_1017_n 0.00508007f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_328 N_CLK_c_320_n N_A_263_409#_c_1017_n 3.06379e-19 $X=1.725 $Y=1.615 $X2=0
+ $Y2=0
cc_329 N_CLK_M1001_g N_A_263_409#_c_1003_n 0.031641f $X=1.725 $Y=2.545 $X2=0
+ $Y2=0
cc_330 N_CLK_c_316_n N_A_263_409#_c_1003_n 0.00331226f $X=2.075 $Y=1.135 $X2=0
+ $Y2=0
cc_331 CLK N_A_263_409#_c_1003_n 9.04713e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_332 N_CLK_c_320_n N_A_263_409#_c_1003_n 0.012071f $X=1.725 $Y=1.615 $X2=0
+ $Y2=0
cc_333 N_CLK_M1001_g N_VPWR_c_1577_n 0.0189165f $X=1.725 $Y=2.545 $X2=0 $Y2=0
cc_334 N_CLK_M1001_g N_VPWR_c_1583_n 0.00769046f $X=1.725 $Y=2.545 $X2=0 $Y2=0
cc_335 N_CLK_M1001_g N_VPWR_c_1574_n 0.0143431f $X=1.725 $Y=2.545 $X2=0 $Y2=0
cc_336 N_CLK_c_315_n N_A_145_409#_c_1715_n 0.00705993f $X=1.79 $Y=1.06 $X2=0
+ $Y2=0
cc_337 N_CLK_c_317_n N_A_145_409#_c_1715_n 2.48962e-19 $X=2.15 $Y=1.06 $X2=0
+ $Y2=0
cc_338 N_CLK_c_315_n N_A_145_409#_c_1716_n 0.004761f $X=1.79 $Y=1.06 $X2=0 $Y2=0
cc_339 N_CLK_c_316_n N_A_145_409#_c_1716_n 0.00310288f $X=2.075 $Y=1.135 $X2=0
+ $Y2=0
cc_340 N_CLK_c_317_n N_A_145_409#_c_1716_n 0.0108002f $X=2.15 $Y=1.06 $X2=0
+ $Y2=0
cc_341 N_CLK_c_316_n N_A_145_409#_c_1717_n 0.00960072f $X=2.075 $Y=1.135 $X2=0
+ $Y2=0
cc_342 N_CLK_c_316_n N_A_145_409#_c_1718_n 0.00711534f $X=2.075 $Y=1.135 $X2=0
+ $Y2=0
cc_343 N_CLK_c_321_n N_A_145_409#_c_1718_n 0.00111729f $X=1.725 $Y=1.45 $X2=0
+ $Y2=0
cc_344 N_CLK_c_317_n N_A_145_409#_c_1719_n 6.89573e-19 $X=2.15 $Y=1.06 $X2=0
+ $Y2=0
cc_345 N_CLK_M1001_g N_A_145_409#_c_1724_n 0.00246486f $X=1.725 $Y=2.545 $X2=0
+ $Y2=0
cc_346 N_CLK_c_315_n N_A_145_409#_c_1724_n 6.39523e-19 $X=1.79 $Y=1.06 $X2=0
+ $Y2=0
cc_347 N_CLK_c_318_n N_A_145_409#_c_1724_n 0.00100521f $X=1.79 $Y=1.135 $X2=0
+ $Y2=0
cc_348 N_CLK_c_315_n N_A_145_409#_c_1725_n 0.00475564f $X=1.79 $Y=1.06 $X2=0
+ $Y2=0
cc_349 N_CLK_c_317_n N_VGND_c_1908_n 9.43806e-19 $X=2.15 $Y=1.06 $X2=0 $Y2=0
cc_350 N_CLK_c_317_n N_VGND_c_1915_n 0.00409299f $X=2.15 $Y=1.06 $X2=0 $Y2=0
cc_351 N_CLK_c_317_n N_VGND_c_1923_n 0.00437698f $X=2.15 $Y=1.06 $X2=0 $Y2=0
cc_352 N_A_476_409#_c_397_p N_A_946_99#_M1003_d 0.0047688f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_353 N_A_476_409#_M1017_g N_A_946_99#_M1008_g 0.0264501f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_354 N_A_476_409#_c_376_n N_A_946_99#_c_582_n 0.00116447f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_355 N_A_476_409#_c_377_n N_A_946_99#_c_582_n 0.042729f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_356 N_A_476_409#_c_397_p N_A_946_99#_c_582_n 9.21303e-19 $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_357 N_A_476_409#_c_402_p N_A_946_99#_M1032_g 0.00180461f $X=4.375 $Y=2.98
+ $X2=0 $Y2=0
cc_358 N_A_476_409#_c_403_p N_A_946_99#_M1032_g 0.00403868f $X=4.46 $Y=2.895
+ $X2=0 $Y2=0
cc_359 N_A_476_409#_c_397_p N_A_946_99#_M1032_g 0.0233251f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_360 N_A_476_409#_c_397_p N_A_946_99#_c_590_n 0.0243994f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_361 N_A_476_409#_c_397_p N_A_946_99#_c_591_n 0.0461265f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_362 N_A_476_409#_c_389_n N_A_712_419#_M1005_d 0.0086935f $X=3.6 $Y=2.895
+ $X2=0 $Y2=0
cc_363 N_A_476_409#_c_402_p N_A_712_419#_M1005_d 0.0159428f $X=4.375 $Y=2.98
+ $X2=0 $Y2=0
cc_364 N_A_476_409#_c_409_p N_A_712_419#_M1005_d 6.69812e-19 $X=3.6 $Y=2.98
+ $X2=0 $Y2=0
cc_365 N_A_476_409#_c_397_p N_A_712_419#_M1003_g 0.0187081f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_366 N_A_476_409#_c_397_p N_A_712_419#_M1018_g 0.020982f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_367 N_A_476_409#_M1009_g N_A_712_419#_M1029_g 0.0417634f $X=7.52 $Y=0.835
+ $X2=0 $Y2=0
cc_368 N_A_476_409#_c_378_n N_A_712_419#_c_662_n 0.00968448f $X=7.5 $Y=2.505
+ $X2=0 $Y2=0
cc_369 N_A_476_409#_c_383_n N_A_712_419#_c_662_n 7.44355e-19 $X=7.745 $Y=1.465
+ $X2=0 $Y2=0
cc_370 N_A_476_409#_c_397_p N_A_712_419#_c_683_n 2.21279e-19 $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_371 N_A_476_409#_M1005_g N_A_712_419#_c_699_n 0.00152258f $X=3.435 $Y=2.595
+ $X2=0 $Y2=0
cc_372 N_A_476_409#_c_389_n N_A_712_419#_c_699_n 0.0343853f $X=3.6 $Y=2.895
+ $X2=0 $Y2=0
cc_373 N_A_476_409#_c_402_p N_A_712_419#_c_699_n 0.0194739f $X=4.375 $Y=2.98
+ $X2=0 $Y2=0
cc_374 N_A_476_409#_c_403_p N_A_712_419#_c_699_n 0.00269616f $X=4.46 $Y=2.895
+ $X2=0 $Y2=0
cc_375 N_A_476_409#_c_420_p N_A_712_419#_c_699_n 0.0129587f $X=4.545 $Y=2.59
+ $X2=0 $Y2=0
cc_376 N_A_476_409#_M1017_g N_A_712_419#_c_663_n 0.00338635f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_377 N_A_476_409#_c_376_n N_A_712_419#_c_684_n 0.0171133f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_378 N_A_476_409#_c_377_n N_A_712_419#_c_684_n 6.69682e-19 $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_379 N_A_476_409#_c_402_p N_A_712_419#_c_684_n 0.00396791f $X=4.375 $Y=2.98
+ $X2=0 $Y2=0
cc_380 N_A_476_409#_c_397_p N_A_712_419#_c_684_n 0.0142858f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_381 N_A_476_409#_c_420_p N_A_712_419#_c_684_n 0.00637416f $X=4.545 $Y=2.59
+ $X2=0 $Y2=0
cc_382 N_A_476_409#_M1005_g N_A_712_419#_c_685_n 6.20042e-19 $X=3.435 $Y=2.595
+ $X2=0 $Y2=0
cc_383 N_A_476_409#_c_389_n N_A_712_419#_c_685_n 0.0133149f $X=3.6 $Y=2.895
+ $X2=0 $Y2=0
cc_384 N_A_476_409#_c_376_n N_A_712_419#_c_685_n 0.0196999f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_385 N_A_476_409#_M1017_g N_A_712_419#_c_664_n 0.0126144f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_386 N_A_476_409#_c_376_n N_A_712_419#_c_664_n 0.00972422f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_387 N_A_476_409#_c_377_n N_A_712_419#_c_664_n 7.36044e-19 $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_388 N_A_476_409#_c_376_n N_A_712_419#_c_665_n 0.0158582f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_389 N_A_476_409#_c_377_n N_A_712_419#_c_665_n 0.00318967f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_390 N_A_476_409#_M1017_g N_A_712_419#_c_666_n 0.00521452f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_391 N_A_476_409#_c_376_n N_A_712_419#_c_666_n 0.0348234f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_392 N_A_476_409#_c_377_n N_A_712_419#_c_666_n 0.00100293f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_393 N_A_476_409#_M1009_g N_A_712_419#_c_677_n 3.5045e-19 $X=7.52 $Y=0.835
+ $X2=0 $Y2=0
cc_394 N_A_476_409#_c_397_p N_A_712_419#_c_677_n 0.00337217f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_395 N_A_476_409#_c_378_n N_A_712_419#_c_677_n 0.0182476f $X=7.5 $Y=2.505
+ $X2=0 $Y2=0
cc_396 N_A_476_409#_c_382_n N_A_712_419#_c_677_n 2.69668e-19 $X=7.58 $Y=1.465
+ $X2=0 $Y2=0
cc_397 N_A_476_409#_c_383_n N_A_712_419#_c_677_n 0.0218887f $X=7.745 $Y=1.465
+ $X2=0 $Y2=0
cc_398 N_A_476_409#_c_382_n N_A_712_419#_c_678_n 0.0209697f $X=7.58 $Y=1.465
+ $X2=0 $Y2=0
cc_399 N_A_476_409#_c_397_p N_SET_B_M1027_g 0.0225097f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_400 N_A_476_409#_M1015_g N_SET_B_c_862_n 0.00812824f $X=8.47 $Y=2.595 $X2=0
+ $Y2=0
cc_401 N_A_476_409#_c_397_p N_SET_B_c_862_n 0.0221796f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_402 N_A_476_409#_c_378_n N_SET_B_c_862_n 0.0220497f $X=7.5 $Y=2.505 $X2=0
+ $Y2=0
cc_403 N_A_476_409#_c_394_n N_SET_B_c_862_n 0.00818755f $X=8.48 $Y=1.77 $X2=0
+ $Y2=0
cc_404 N_A_476_409#_c_380_n N_SET_B_c_862_n 0.00133741f $X=8.48 $Y=1.77 $X2=0
+ $Y2=0
cc_405 N_A_476_409#_c_382_n N_SET_B_c_862_n 8.24116e-19 $X=7.58 $Y=1.465 $X2=0
+ $Y2=0
cc_406 N_A_476_409#_c_383_n N_SET_B_c_862_n 0.0217434f $X=7.745 $Y=1.465 $X2=0
+ $Y2=0
cc_407 N_A_476_409#_c_397_p N_SET_B_c_875_n 0.00353311f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_408 N_A_476_409#_c_397_p N_SET_B_c_856_n 0.00697942f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_409 N_A_476_409#_c_397_p N_SET_B_c_857_n 7.95656e-19 $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_410 N_A_476_409#_c_386_n N_A_263_409#_M1026_g 0.0108317f $X=2.52 $Y=2.475
+ $X2=0 $Y2=0
cc_411 N_A_476_409#_c_388_n N_A_263_409#_M1026_g 0.00359736f $X=2.685 $Y=2.98
+ $X2=0 $Y2=0
cc_412 N_A_476_409#_c_374_n N_A_263_409#_c_987_n 3.49778e-19 $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_413 N_A_476_409#_c_374_n N_A_263_409#_c_988_n 6.26784e-19 $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_414 N_A_476_409#_c_375_n N_A_263_409#_c_988_n 0.00176338f $X=3.685 $Y=1.555
+ $X2=0 $Y2=0
cc_415 N_A_476_409#_c_381_n N_A_263_409#_c_988_n 0.00491746f $X=3.395 $Y=1.615
+ $X2=0 $Y2=0
cc_416 N_A_476_409#_c_374_n N_A_263_409#_c_990_n 0.00623642f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_417 N_A_476_409#_c_374_n N_A_263_409#_c_991_n 0.021909f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_418 N_A_476_409#_c_375_n N_A_263_409#_c_991_n 0.00924413f $X=3.685 $Y=1.555
+ $X2=0 $Y2=0
cc_419 N_A_476_409#_c_381_n N_A_263_409#_c_991_n 0.0168615f $X=3.395 $Y=1.615
+ $X2=0 $Y2=0
cc_420 N_A_476_409#_M1017_g N_A_263_409#_c_992_n 0.00897248f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_421 N_A_476_409#_c_374_n N_A_263_409#_c_992_n 0.00324629f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_422 N_A_476_409#_c_376_n N_A_263_409#_c_992_n 6.37995e-19 $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_423 N_A_476_409#_c_374_n N_A_263_409#_c_993_n 0.00320191f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_424 N_A_476_409#_c_389_n N_A_263_409#_c_993_n 0.00537872f $X=3.6 $Y=2.895
+ $X2=0 $Y2=0
cc_425 N_A_476_409#_c_376_n N_A_263_409#_c_993_n 0.029096f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_426 N_A_476_409#_c_377_n N_A_263_409#_c_993_n 0.0180853f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_427 N_A_476_409#_c_381_n N_A_263_409#_c_993_n 0.0153399f $X=3.395 $Y=1.615
+ $X2=0 $Y2=0
cc_428 N_A_476_409#_M1017_g N_A_263_409#_M1020_g 0.0133216f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_429 N_A_476_409#_c_374_n N_A_263_409#_M1020_g 0.00194081f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_430 N_A_476_409#_c_376_n N_A_263_409#_c_1006_n 0.00802552f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_431 N_A_476_409#_c_377_n N_A_263_409#_c_1006_n 0.015098f $X=4.355 $Y=1.495
+ $X2=0 $Y2=0
cc_432 N_A_476_409#_M1005_g N_A_263_409#_c_1007_n 0.0153399f $X=3.435 $Y=2.595
+ $X2=0 $Y2=0
cc_433 N_A_476_409#_M1017_g N_A_263_409#_c_995_n 0.00865213f $X=4.445 $Y=0.835
+ $X2=0 $Y2=0
cc_434 N_A_476_409#_M1009_g N_A_263_409#_c_995_n 0.00907339f $X=7.52 $Y=0.835
+ $X2=0 $Y2=0
cc_435 N_A_476_409#_M1005_g N_A_263_409#_c_1008_n 0.0145942f $X=3.435 $Y=2.595
+ $X2=0 $Y2=0
cc_436 N_A_476_409#_c_389_n N_A_263_409#_c_1008_n 0.00490093f $X=3.6 $Y=2.895
+ $X2=0 $Y2=0
cc_437 N_A_476_409#_c_402_p N_A_263_409#_c_1008_n 0.0163067f $X=4.375 $Y=2.98
+ $X2=0 $Y2=0
cc_438 N_A_476_409#_c_403_p N_A_263_409#_c_1008_n 0.0102029f $X=4.46 $Y=2.895
+ $X2=0 $Y2=0
cc_439 N_A_476_409#_c_420_p N_A_263_409#_c_1008_n 0.00640761f $X=4.545 $Y=2.59
+ $X2=0 $Y2=0
cc_440 N_A_476_409#_M1015_g N_A_263_409#_c_1009_n 0.0144374f $X=8.47 $Y=2.595
+ $X2=0 $Y2=0
cc_441 N_A_476_409#_c_397_p N_A_263_409#_c_1009_n 0.00882806f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_442 N_A_476_409#_c_378_n N_A_263_409#_c_1009_n 0.0126461f $X=7.5 $Y=2.505
+ $X2=0 $Y2=0
cc_443 N_A_476_409#_M1015_g N_A_263_409#_c_1010_n 0.00529911f $X=8.47 $Y=2.595
+ $X2=0 $Y2=0
cc_444 N_A_476_409#_c_379_n N_A_263_409#_c_1010_n 0.00491141f $X=8.315 $Y=1.545
+ $X2=0 $Y2=0
cc_445 N_A_476_409#_c_378_n N_A_263_409#_c_1011_n 0.00909518f $X=7.5 $Y=2.505
+ $X2=0 $Y2=0
cc_446 N_A_476_409#_c_382_n N_A_263_409#_c_1011_n 0.0171208f $X=7.58 $Y=1.465
+ $X2=0 $Y2=0
cc_447 N_A_476_409#_c_383_n N_A_263_409#_c_1011_n 0.00124929f $X=7.745 $Y=1.465
+ $X2=0 $Y2=0
cc_448 N_A_476_409#_M1009_g N_A_263_409#_M1000_g 0.0204057f $X=7.52 $Y=0.835
+ $X2=0 $Y2=0
cc_449 N_A_476_409#_c_378_n N_A_263_409#_M1000_g 0.00415307f $X=7.5 $Y=2.505
+ $X2=0 $Y2=0
cc_450 N_A_476_409#_c_379_n N_A_263_409#_M1000_g 0.0133649f $X=8.315 $Y=1.545
+ $X2=0 $Y2=0
cc_451 N_A_476_409#_c_394_n N_A_263_409#_M1000_g 0.00218718f $X=8.48 $Y=1.77
+ $X2=0 $Y2=0
cc_452 N_A_476_409#_c_380_n N_A_263_409#_M1000_g 0.0222538f $X=8.48 $Y=1.77
+ $X2=0 $Y2=0
cc_453 N_A_476_409#_c_382_n N_A_263_409#_M1000_g 0.0205198f $X=7.58 $Y=1.465
+ $X2=0 $Y2=0
cc_454 N_A_476_409#_c_383_n N_A_263_409#_M1000_g 0.00106267f $X=7.745 $Y=1.465
+ $X2=0 $Y2=0
cc_455 N_A_476_409#_c_374_n N_A_263_409#_c_999_n 0.0028974f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_456 N_A_476_409#_c_375_n N_A_263_409#_c_999_n 0.00153296f $X=3.685 $Y=1.555
+ $X2=0 $Y2=0
cc_457 N_A_476_409#_M1026_d N_A_263_409#_c_1015_n 0.00121183f $X=2.38 $Y=2.045
+ $X2=0 $Y2=0
cc_458 N_A_476_409#_c_386_n N_A_263_409#_c_1015_n 0.00383775f $X=2.52 $Y=2.475
+ $X2=0 $Y2=0
cc_459 N_A_476_409#_M1005_g N_A_263_409#_c_1003_n 0.00128846f $X=3.435 $Y=2.595
+ $X2=0 $Y2=0
cc_460 N_A_476_409#_c_386_n N_A_263_409#_c_1003_n 0.0068691f $X=2.52 $Y=2.475
+ $X2=0 $Y2=0
cc_461 N_A_476_409#_c_379_n N_A_1686_40#_c_1192_n 0.00170606f $X=8.315 $Y=1.545
+ $X2=0 $Y2=0
cc_462 N_A_476_409#_c_380_n N_A_1686_40#_c_1192_n 0.0120516f $X=8.48 $Y=1.77
+ $X2=0 $Y2=0
cc_463 N_A_476_409#_M1015_g N_A_1686_40#_M1033_g 0.0601746f $X=8.47 $Y=2.595
+ $X2=0 $Y2=0
cc_464 N_A_476_409#_c_379_n N_A_1686_40#_c_1195_n 8.64347e-19 $X=8.315 $Y=1.545
+ $X2=0 $Y2=0
cc_465 N_A_476_409#_c_394_n N_A_1686_40#_c_1195_n 2.76776e-19 $X=8.48 $Y=1.77
+ $X2=0 $Y2=0
cc_466 N_A_476_409#_c_380_n N_A_1686_40#_c_1195_n 0.017217f $X=8.48 $Y=1.77
+ $X2=0 $Y2=0
cc_467 N_A_476_409#_c_397_p N_A_1519_125#_c_1324_n 0.0114736f $X=7.415 $Y=2.59
+ $X2=0 $Y2=0
cc_468 N_A_476_409#_c_379_n N_A_1519_125#_c_1307_n 0.0214314f $X=8.315 $Y=1.545
+ $X2=0 $Y2=0
cc_469 N_A_476_409#_c_380_n N_A_1519_125#_c_1307_n 6.31835e-19 $X=8.48 $Y=1.77
+ $X2=0 $Y2=0
cc_470 N_A_476_409#_M1009_g N_A_1519_125#_c_1308_n 0.003274f $X=7.52 $Y=0.835
+ $X2=0 $Y2=0
cc_471 N_A_476_409#_c_379_n N_A_1519_125#_c_1308_n 0.0150765f $X=8.315 $Y=1.545
+ $X2=0 $Y2=0
cc_472 N_A_476_409#_c_382_n N_A_1519_125#_c_1308_n 0.00210396f $X=7.58 $Y=1.465
+ $X2=0 $Y2=0
cc_473 N_A_476_409#_c_383_n N_A_1519_125#_c_1308_n 0.00608888f $X=7.745 $Y=1.465
+ $X2=0 $Y2=0
cc_474 N_A_476_409#_M1015_g N_A_1519_125#_c_1331_n 0.0194756f $X=8.47 $Y=2.595
+ $X2=0 $Y2=0
cc_475 N_A_476_409#_c_394_n N_A_1519_125#_c_1331_n 0.00470629f $X=8.48 $Y=1.77
+ $X2=0 $Y2=0
cc_476 N_A_476_409#_M1015_g N_A_1519_125#_c_1309_n 0.00513213f $X=8.47 $Y=2.595
+ $X2=0 $Y2=0
cc_477 N_A_476_409#_c_379_n N_A_1519_125#_c_1309_n 0.0136719f $X=8.315 $Y=1.545
+ $X2=0 $Y2=0
cc_478 N_A_476_409#_c_394_n N_A_1519_125#_c_1309_n 0.0215584f $X=8.48 $Y=1.77
+ $X2=0 $Y2=0
cc_479 N_A_476_409#_c_380_n N_A_1519_125#_c_1309_n 0.0021337f $X=8.48 $Y=1.77
+ $X2=0 $Y2=0
cc_480 N_A_476_409#_M1015_g N_A_1519_125#_c_1321_n 0.0187883f $X=8.47 $Y=2.595
+ $X2=0 $Y2=0
cc_481 N_A_476_409#_c_378_n N_A_1519_125#_c_1321_n 0.0257837f $X=7.5 $Y=2.505
+ $X2=0 $Y2=0
cc_482 N_A_476_409#_c_379_n N_A_1519_125#_c_1321_n 0.00766198f $X=8.315 $Y=1.545
+ $X2=0 $Y2=0
cc_483 N_A_476_409#_c_397_p N_VPWR_M1032_d 0.0159709f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_484 N_A_476_409#_c_397_p N_VPWR_M1027_d 0.0121213f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_485 N_A_476_409#_c_386_n N_VPWR_c_1577_n 0.0385131f $X=2.52 $Y=2.475 $X2=0
+ $Y2=0
cc_486 N_A_476_409#_c_388_n N_VPWR_c_1577_n 0.0119061f $X=2.685 $Y=2.98 $X2=0
+ $Y2=0
cc_487 N_A_476_409#_c_402_p N_VPWR_c_1578_n 0.0067281f $X=4.375 $Y=2.98 $X2=0
+ $Y2=0
cc_488 N_A_476_409#_c_403_p N_VPWR_c_1578_n 0.00139649f $X=4.46 $Y=2.895 $X2=0
+ $Y2=0
cc_489 N_A_476_409#_c_397_p N_VPWR_c_1578_n 0.0196062f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_490 N_A_476_409#_c_397_p N_VPWR_c_1579_n 0.0238466f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_491 N_A_476_409#_M1015_g N_VPWR_c_1580_n 0.00263095f $X=8.47 $Y=2.595 $X2=0
+ $Y2=0
cc_492 N_A_476_409#_c_397_p N_VPWR_c_1585_n 0.0174681f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_493 N_A_476_409#_M1005_g N_VPWR_c_1587_n 0.00599878f $X=3.435 $Y=2.595 $X2=0
+ $Y2=0
cc_494 N_A_476_409#_c_387_n N_VPWR_c_1587_n 0.0478968f $X=3.515 $Y=2.98 $X2=0
+ $Y2=0
cc_495 N_A_476_409#_c_388_n N_VPWR_c_1587_n 0.0221635f $X=2.685 $Y=2.98 $X2=0
+ $Y2=0
cc_496 N_A_476_409#_c_402_p N_VPWR_c_1587_n 0.0483813f $X=4.375 $Y=2.98 $X2=0
+ $Y2=0
cc_497 N_A_476_409#_c_397_p N_VPWR_c_1587_n 0.00666313f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_498 N_A_476_409#_c_409_p N_VPWR_c_1587_n 0.00921724f $X=3.6 $Y=2.98 $X2=0
+ $Y2=0
cc_499 N_A_476_409#_M1015_g N_VPWR_c_1588_n 0.00975641f $X=8.47 $Y=2.595 $X2=0
+ $Y2=0
cc_500 N_A_476_409#_c_397_p N_VPWR_c_1588_n 0.0111957f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_501 N_A_476_409#_M1005_g N_VPWR_c_1574_n 0.0100086f $X=3.435 $Y=2.595 $X2=0
+ $Y2=0
cc_502 N_A_476_409#_M1015_g N_VPWR_c_1574_n 0.0105056f $X=8.47 $Y=2.595 $X2=0
+ $Y2=0
cc_503 N_A_476_409#_c_387_n N_VPWR_c_1574_n 0.0300734f $X=3.515 $Y=2.98 $X2=0
+ $Y2=0
cc_504 N_A_476_409#_c_388_n N_VPWR_c_1574_n 0.0126536f $X=2.685 $Y=2.98 $X2=0
+ $Y2=0
cc_505 N_A_476_409#_c_402_p N_VPWR_c_1574_n 0.0311775f $X=4.375 $Y=2.98 $X2=0
+ $Y2=0
cc_506 N_A_476_409#_c_397_p N_VPWR_c_1574_n 0.0646345f $X=7.415 $Y=2.59 $X2=0
+ $Y2=0
cc_507 N_A_476_409#_c_409_p N_VPWR_c_1574_n 0.00636028f $X=3.6 $Y=2.98 $X2=0
+ $Y2=0
cc_508 N_A_476_409#_c_387_n N_A_145_409#_M1005_s 0.00564752f $X=3.515 $Y=2.98
+ $X2=0 $Y2=0
cc_509 N_A_476_409#_c_374_n N_A_145_409#_c_1719_n 0.0212837f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_510 N_A_476_409#_M1005_g N_A_145_409#_c_1720_n 0.00365402f $X=3.435 $Y=2.595
+ $X2=0 $Y2=0
cc_511 N_A_476_409#_c_374_n N_A_145_409#_c_1720_n 0.00453283f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_512 N_A_476_409#_c_375_n N_A_145_409#_c_1720_n 0.036332f $X=3.685 $Y=1.555
+ $X2=0 $Y2=0
cc_513 N_A_476_409#_c_381_n N_A_145_409#_c_1720_n 7.37948e-19 $X=3.395 $Y=1.615
+ $X2=0 $Y2=0
cc_514 N_A_476_409#_c_374_n N_A_145_409#_c_1721_n 0.0221619f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_515 N_A_476_409#_M1005_g N_A_145_409#_c_1730_n 0.00728752f $X=3.435 $Y=2.595
+ $X2=0 $Y2=0
cc_516 N_A_476_409#_c_389_n N_A_145_409#_c_1730_n 0.012389f $X=3.6 $Y=2.895
+ $X2=0 $Y2=0
cc_517 N_A_476_409#_c_375_n N_A_145_409#_c_1730_n 0.0292335f $X=3.685 $Y=1.555
+ $X2=0 $Y2=0
cc_518 N_A_476_409#_c_381_n N_A_145_409#_c_1730_n 0.00185447f $X=3.395 $Y=1.615
+ $X2=0 $Y2=0
cc_519 N_A_476_409#_M1026_d N_A_145_409#_c_1731_n 0.00115503f $X=2.38 $Y=2.045
+ $X2=0 $Y2=0
cc_520 N_A_476_409#_c_386_n N_A_145_409#_c_1731_n 0.00386824f $X=2.52 $Y=2.475
+ $X2=0 $Y2=0
cc_521 N_A_476_409#_M1005_g N_A_145_409#_c_1732_n 0.0140272f $X=3.435 $Y=2.595
+ $X2=0 $Y2=0
cc_522 N_A_476_409#_c_386_n N_A_145_409#_c_1732_n 0.0217627f $X=2.52 $Y=2.475
+ $X2=0 $Y2=0
cc_523 N_A_476_409#_c_387_n N_A_145_409#_c_1732_n 0.0196206f $X=3.515 $Y=2.98
+ $X2=0 $Y2=0
cc_524 N_A_476_409#_c_389_n N_A_145_409#_c_1732_n 0.0398689f $X=3.6 $Y=2.895
+ $X2=0 $Y2=0
cc_525 N_A_476_409#_c_374_n N_A_145_409#_c_1723_n 0.0207906f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_526 N_A_476_409#_c_375_n N_A_145_409#_c_1723_n 0.0147418f $X=3.685 $Y=1.555
+ $X2=0 $Y2=0
cc_527 N_A_476_409#_c_374_n N_A_145_409#_c_1726_n 0.0134816f $X=3.155 $Y=0.81
+ $X2=0 $Y2=0
cc_528 N_A_476_409#_c_402_p A_884_419# 0.00293005f $X=4.375 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_529 N_A_476_409#_c_403_p A_884_419# 0.00263862f $X=4.46 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_530 N_A_476_409#_c_397_p A_884_419# 0.00478283f $X=7.415 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_531 N_A_476_409#_c_420_p A_884_419# 9.0912e-19 $X=4.545 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_532 N_A_476_409#_c_397_p A_1441_419# 0.00434279f $X=7.415 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_533 N_A_476_409#_M1009_g N_VGND_c_1910_n 0.00189704f $X=7.52 $Y=0.835 $X2=0
+ $Y2=0
cc_534 N_A_476_409#_M1017_g N_VGND_c_1923_n 9.49986e-19 $X=4.445 $Y=0.835 $X2=0
+ $Y2=0
cc_535 N_A_476_409#_M1009_g N_VGND_c_1923_n 9.49986e-19 $X=7.52 $Y=0.835 $X2=0
+ $Y2=0
cc_536 N_A_946_99#_M1032_g N_A_712_419#_M1003_g 0.0176391f $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_537 N_A_946_99#_c_589_n N_A_712_419#_M1003_g 0.00433088f $X=5.215 $Y=2.075
+ $X2=0 $Y2=0
cc_538 N_A_946_99#_c_591_n N_A_712_419#_M1003_g 0.0180572f $X=6.05 $Y=2.24 $X2=0
+ $Y2=0
cc_539 N_A_946_99#_c_585_n N_A_712_419#_M1034_g 0.00303189f $X=5.78 $Y=1.215
+ $X2=0 $Y2=0
cc_540 N_A_946_99#_c_586_n N_A_712_419#_M1034_g 0.00643264f $X=5.955 $Y=0.84
+ $X2=0 $Y2=0
cc_541 N_A_946_99#_c_582_n N_A_712_419#_c_661_n 0.00946257f $X=4.885 $Y=1.885
+ $X2=0 $Y2=0
cc_542 N_A_946_99#_c_584_n N_A_712_419#_c_661_n 0.00672112f $X=5.695 $Y=1.3
+ $X2=0 $Y2=0
cc_543 N_A_946_99#_c_586_n N_A_712_419#_c_661_n 0.00639222f $X=5.955 $Y=0.84
+ $X2=0 $Y2=0
cc_544 N_A_946_99#_M1032_g N_A_712_419#_c_699_n 0.00120947f $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_545 N_A_946_99#_M1032_g N_A_712_419#_c_684_n 0.00762113f $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_546 N_A_946_99#_c_590_n N_A_712_419#_c_684_n 0.00772304f $X=5.38 $Y=2.2 $X2=0
+ $Y2=0
cc_547 N_A_946_99#_M1008_g N_A_712_419#_c_666_n 0.00766293f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_548 N_A_946_99#_c_582_n N_A_712_419#_c_666_n 0.0222544f $X=4.885 $Y=1.885
+ $X2=0 $Y2=0
cc_549 N_A_946_99#_M1032_g N_A_712_419#_c_666_n 0.00480674f $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_550 N_A_946_99#_c_583_n N_A_712_419#_c_666_n 0.0123662f $X=5.215 $Y=1.385
+ $X2=0 $Y2=0
cc_551 N_A_946_99#_c_589_n N_A_712_419#_c_666_n 0.0477088f $X=5.215 $Y=2.075
+ $X2=0 $Y2=0
cc_552 N_A_946_99#_M1008_g N_A_712_419#_c_667_n 0.00465503f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_553 N_A_946_99#_c_582_n N_A_712_419#_c_667_n 0.00828624f $X=4.885 $Y=1.885
+ $X2=0 $Y2=0
cc_554 N_A_946_99#_c_583_n N_A_712_419#_c_667_n 0.0252887f $X=5.215 $Y=1.385
+ $X2=0 $Y2=0
cc_555 N_A_946_99#_c_584_n N_A_712_419#_c_667_n 0.0109129f $X=5.695 $Y=1.3 $X2=0
+ $Y2=0
cc_556 N_A_946_99#_c_586_n N_A_712_419#_c_667_n 0.0147702f $X=5.955 $Y=0.84
+ $X2=0 $Y2=0
cc_557 N_A_946_99#_M1008_g N_A_712_419#_c_668_n 0.00475951f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_558 N_A_946_99#_c_586_n N_A_712_419#_c_668_n 0.0193977f $X=5.955 $Y=0.84
+ $X2=0 $Y2=0
cc_559 N_A_946_99#_c_586_n N_A_712_419#_c_669_n 0.0308596f $X=5.955 $Y=0.84
+ $X2=0 $Y2=0
cc_560 N_A_946_99#_c_582_n N_A_712_419#_c_671_n 0.0013234f $X=4.885 $Y=1.885
+ $X2=0 $Y2=0
cc_561 N_A_946_99#_c_589_n N_A_712_419#_c_671_n 0.019676f $X=5.215 $Y=2.075
+ $X2=0 $Y2=0
cc_562 N_A_946_99#_c_584_n N_A_712_419#_c_671_n 0.0180217f $X=5.695 $Y=1.3 $X2=0
+ $Y2=0
cc_563 N_A_946_99#_c_591_n N_A_712_419#_c_671_n 0.0444498f $X=6.05 $Y=2.24 $X2=0
+ $Y2=0
cc_564 N_A_946_99#_c_586_n N_A_712_419#_c_671_n 0.00690068f $X=5.955 $Y=0.84
+ $X2=0 $Y2=0
cc_565 N_A_946_99#_c_582_n N_A_712_419#_c_672_n 0.0179213f $X=4.885 $Y=1.885
+ $X2=0 $Y2=0
cc_566 N_A_946_99#_c_589_n N_A_712_419#_c_672_n 4.48216e-19 $X=5.215 $Y=2.075
+ $X2=0 $Y2=0
cc_567 N_A_946_99#_c_584_n N_A_712_419#_c_672_n 0.00459325f $X=5.695 $Y=1.3
+ $X2=0 $Y2=0
cc_568 N_A_946_99#_c_591_n N_A_712_419#_c_672_n 0.00194249f $X=6.05 $Y=2.24
+ $X2=0 $Y2=0
cc_569 N_A_946_99#_c_589_n N_A_712_419#_c_673_n 0.00392036f $X=5.215 $Y=2.075
+ $X2=0 $Y2=0
cc_570 N_A_946_99#_c_584_n N_A_712_419#_c_674_n 0.00117634f $X=5.695 $Y=1.3
+ $X2=0 $Y2=0
cc_571 N_A_946_99#_c_585_n N_A_712_419#_c_674_n 0.00584978f $X=5.78 $Y=1.215
+ $X2=0 $Y2=0
cc_572 N_A_946_99#_c_586_n N_A_712_419#_c_674_n 0.0177205f $X=5.955 $Y=0.84
+ $X2=0 $Y2=0
cc_573 N_A_946_99#_c_589_n N_A_712_419#_c_676_n 8.46358e-19 $X=5.215 $Y=2.075
+ $X2=0 $Y2=0
cc_574 N_A_946_99#_c_584_n N_A_712_419#_c_676_n 0.0112835f $X=5.695 $Y=1.3 $X2=0
+ $Y2=0
cc_575 N_A_946_99#_c_586_n N_A_712_419#_c_676_n 0.00546182f $X=5.955 $Y=0.84
+ $X2=0 $Y2=0
cc_576 N_A_946_99#_M1008_g N_A_712_419#_c_767_n 0.00744392f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_577 N_A_946_99#_c_589_n N_A_712_419#_c_679_n 7.05606e-19 $X=5.215 $Y=2.075
+ $X2=0 $Y2=0
cc_578 N_A_946_99#_c_584_n N_A_712_419#_c_679_n 0.00148137f $X=5.695 $Y=1.3
+ $X2=0 $Y2=0
cc_579 N_A_946_99#_c_591_n N_SET_B_M1027_g 0.0105502f $X=6.05 $Y=2.24 $X2=0
+ $Y2=0
cc_580 N_A_946_99#_c_591_n N_SET_B_c_875_n 0.00213762f $X=6.05 $Y=2.24 $X2=0
+ $Y2=0
cc_581 N_A_946_99#_c_591_n N_SET_B_c_856_n 0.00458741f $X=6.05 $Y=2.24 $X2=0
+ $Y2=0
cc_582 N_A_946_99#_c_582_n N_A_263_409#_c_1006_n 0.0243832f $X=4.885 $Y=1.885
+ $X2=0 $Y2=0
cc_583 N_A_946_99#_M1008_g N_A_263_409#_c_995_n 0.00865112f $X=4.805 $Y=0.835
+ $X2=0 $Y2=0
cc_584 N_A_946_99#_M1032_g N_A_263_409#_c_1008_n 0.0243832f $X=4.885 $Y=2.595
+ $X2=0 $Y2=0
cc_585 N_A_946_99#_c_590_n N_VPWR_M1032_d 0.00754175f $X=5.38 $Y=2.2 $X2=0 $Y2=0
cc_586 N_A_946_99#_c_591_n N_VPWR_M1032_d 0.00370683f $X=6.05 $Y=2.24 $X2=0
+ $Y2=0
cc_587 N_A_946_99#_M1032_g N_VPWR_c_1578_n 0.0104296f $X=4.885 $Y=2.595 $X2=0
+ $Y2=0
cc_588 N_A_946_99#_M1032_g N_VPWR_c_1587_n 0.00641304f $X=4.885 $Y=2.595 $X2=0
+ $Y2=0
cc_589 N_A_946_99#_M1003_d N_VPWR_c_1574_n 0.00333718f $X=5.91 $Y=2.095 $X2=0
+ $Y2=0
cc_590 N_A_946_99#_M1032_g N_VPWR_c_1574_n 0.00732096f $X=4.885 $Y=2.595 $X2=0
+ $Y2=0
cc_591 N_A_946_99#_M1008_g N_VGND_c_1909_n 0.00488157f $X=4.805 $Y=0.835 $X2=0
+ $Y2=0
cc_592 N_A_946_99#_M1008_g N_VGND_c_1923_n 9.49986e-19 $X=4.805 $Y=0.835 $X2=0
+ $Y2=0
cc_593 N_A_712_419#_M1018_g N_SET_B_M1027_g 0.0311542f $X=7.08 $Y=2.595 $X2=0
+ $Y2=0
cc_594 N_A_712_419#_M1034_g N_SET_B_M1022_g 0.0391773f $X=6.17 $Y=0.835 $X2=0
+ $Y2=0
cc_595 N_A_712_419#_M1029_g N_SET_B_M1022_g 0.0132779f $X=7.13 $Y=0.835 $X2=0
+ $Y2=0
cc_596 N_A_712_419#_c_671_n N_SET_B_M1022_g 5.0341e-19 $X=6.045 $Y=1.73 $X2=0
+ $Y2=0
cc_597 N_A_712_419#_c_673_n N_SET_B_M1022_g 0.00160166f $X=6.13 $Y=1.565 $X2=0
+ $Y2=0
cc_598 N_A_712_419#_c_674_n N_SET_B_M1022_g 0.00739191f $X=6.385 $Y=1.245 $X2=0
+ $Y2=0
cc_599 N_A_712_419#_c_675_n N_SET_B_M1022_g 0.0149115f $X=6.875 $Y=1.33 $X2=0
+ $Y2=0
cc_600 N_A_712_419#_c_677_n N_SET_B_M1022_g 7.66983e-19 $X=7.04 $Y=1.41 $X2=0
+ $Y2=0
cc_601 N_A_712_419#_c_678_n N_SET_B_M1022_g 0.0193547f $X=7.04 $Y=1.41 $X2=0
+ $Y2=0
cc_602 N_A_712_419#_c_679_n N_SET_B_M1022_g 0.00342877f $X=5.785 $Y=1.565 $X2=0
+ $Y2=0
cc_603 N_A_712_419#_M1018_g N_SET_B_c_862_n 0.00872782f $X=7.08 $Y=2.595 $X2=0
+ $Y2=0
cc_604 N_A_712_419#_c_675_n N_SET_B_c_862_n 0.00680665f $X=6.875 $Y=1.33 $X2=0
+ $Y2=0
cc_605 N_A_712_419#_c_677_n N_SET_B_c_862_n 0.0114042f $X=7.04 $Y=1.41 $X2=0
+ $Y2=0
cc_606 N_A_712_419#_M1003_g N_SET_B_c_875_n 7.4775e-19 $X=5.785 $Y=2.595 $X2=0
+ $Y2=0
cc_607 N_A_712_419#_c_676_n N_SET_B_c_875_n 0.00274858f $X=6.47 $Y=1.33 $X2=0
+ $Y2=0
cc_608 N_A_712_419#_M1003_g N_SET_B_c_856_n 0.00132031f $X=5.785 $Y=2.595 $X2=0
+ $Y2=0
cc_609 N_A_712_419#_M1018_g N_SET_B_c_856_n 0.00391297f $X=7.08 $Y=2.595 $X2=0
+ $Y2=0
cc_610 N_A_712_419#_c_662_n N_SET_B_c_856_n 0.00107785f $X=7.04 $Y=1.75 $X2=0
+ $Y2=0
cc_611 N_A_712_419#_c_671_n N_SET_B_c_856_n 0.0215561f $X=6.045 $Y=1.73 $X2=0
+ $Y2=0
cc_612 N_A_712_419#_c_676_n N_SET_B_c_856_n 0.0179594f $X=6.47 $Y=1.33 $X2=0
+ $Y2=0
cc_613 N_A_712_419#_c_677_n N_SET_B_c_856_n 0.0193167f $X=7.04 $Y=1.41 $X2=0
+ $Y2=0
cc_614 N_A_712_419#_M1003_g N_SET_B_c_857_n 0.0503031f $X=5.785 $Y=2.595 $X2=0
+ $Y2=0
cc_615 N_A_712_419#_M1018_g N_SET_B_c_857_n 9.59604e-19 $X=7.08 $Y=2.595 $X2=0
+ $Y2=0
cc_616 N_A_712_419#_c_661_n N_SET_B_c_857_n 0.00307435f $X=6.17 $Y=1.29 $X2=0
+ $Y2=0
cc_617 N_A_712_419#_c_662_n N_SET_B_c_857_n 0.0193959f $X=7.04 $Y=1.75 $X2=0
+ $Y2=0
cc_618 N_A_712_419#_c_671_n N_SET_B_c_857_n 0.00839444f $X=6.045 $Y=1.73 $X2=0
+ $Y2=0
cc_619 N_A_712_419#_c_672_n N_SET_B_c_857_n 0.0159864f $X=5.785 $Y=1.73 $X2=0
+ $Y2=0
cc_620 N_A_712_419#_c_676_n N_SET_B_c_857_n 0.00739497f $X=6.47 $Y=1.33 $X2=0
+ $Y2=0
cc_621 N_A_712_419#_c_677_n N_SET_B_c_857_n 0.00115553f $X=7.04 $Y=1.41 $X2=0
+ $Y2=0
cc_622 N_A_712_419#_c_663_n N_A_263_409#_M1020_g 0.00474949f $X=4.21 $Y=0.865
+ $X2=0 $Y2=0
cc_623 N_A_712_419#_c_665_n N_A_263_409#_M1020_g 0.00572819f $X=4.335 $Y=0.965
+ $X2=0 $Y2=0
cc_624 N_A_712_419#_c_666_n N_A_263_409#_c_1006_n 0.00400794f $X=4.785 $Y=2.075
+ $X2=0 $Y2=0
cc_625 N_A_712_419#_c_685_n N_A_263_409#_c_1007_n 0.00839223f $X=4.195 $Y=2.16
+ $X2=0 $Y2=0
cc_626 N_A_712_419#_M1034_g N_A_263_409#_c_995_n 0.00737233f $X=6.17 $Y=0.835
+ $X2=0 $Y2=0
cc_627 N_A_712_419#_M1029_g N_A_263_409#_c_995_n 0.00894529f $X=7.13 $Y=0.835
+ $X2=0 $Y2=0
cc_628 N_A_712_419#_c_663_n N_A_263_409#_c_995_n 0.00557013f $X=4.21 $Y=0.865
+ $X2=0 $Y2=0
cc_629 N_A_712_419#_c_664_n N_A_263_409#_c_995_n 0.00350913f $X=4.7 $Y=0.965
+ $X2=0 $Y2=0
cc_630 N_A_712_419#_c_667_n N_A_263_409#_c_995_n 0.00466247f $X=5.345 $Y=0.95
+ $X2=0 $Y2=0
cc_631 N_A_712_419#_c_669_n N_A_263_409#_c_995_n 0.0201004f $X=6.3 $Y=0.35 $X2=0
+ $Y2=0
cc_632 N_A_712_419#_c_670_n N_A_263_409#_c_995_n 0.00418768f $X=5.515 $Y=0.35
+ $X2=0 $Y2=0
cc_633 N_A_712_419#_c_767_n N_A_263_409#_c_995_n 4.4656e-19 $X=4.785 $Y=0.965
+ $X2=0 $Y2=0
cc_634 N_A_712_419#_c_699_n N_A_263_409#_c_1008_n 0.0112107f $X=4.03 $Y=2.395
+ $X2=0 $Y2=0
cc_635 N_A_712_419#_c_684_n N_A_263_409#_c_1008_n 0.0145132f $X=4.7 $Y=2.16
+ $X2=0 $Y2=0
cc_636 N_A_712_419#_c_685_n N_A_263_409#_c_1008_n 0.00267092f $X=4.195 $Y=2.16
+ $X2=0 $Y2=0
cc_637 N_A_712_419#_M1018_g N_A_263_409#_c_1009_n 0.0378072f $X=7.08 $Y=2.595
+ $X2=0 $Y2=0
cc_638 N_A_712_419#_c_683_n N_A_263_409#_c_1011_n 0.0378072f $X=7.04 $Y=1.915
+ $X2=0 $Y2=0
cc_639 N_A_712_419#_M1003_g N_VPWR_c_1578_n 0.00718354f $X=5.785 $Y=2.595 $X2=0
+ $Y2=0
cc_640 N_A_712_419#_M1018_g N_VPWR_c_1579_n 0.00938575f $X=7.08 $Y=2.595 $X2=0
+ $Y2=0
cc_641 N_A_712_419#_M1003_g N_VPWR_c_1585_n 0.00713369f $X=5.785 $Y=2.595 $X2=0
+ $Y2=0
cc_642 N_A_712_419#_M1018_g N_VPWR_c_1588_n 0.00713369f $X=7.08 $Y=2.595 $X2=0
+ $Y2=0
cc_643 N_A_712_419#_M1005_d N_VPWR_c_1574_n 0.00499582f $X=3.56 $Y=2.095 $X2=0
+ $Y2=0
cc_644 N_A_712_419#_M1003_g N_VPWR_c_1574_n 0.00975378f $X=5.785 $Y=2.595 $X2=0
+ $Y2=0
cc_645 N_A_712_419#_M1018_g N_VPWR_c_1574_n 0.00943869f $X=7.08 $Y=2.595 $X2=0
+ $Y2=0
cc_646 N_A_712_419#_c_663_n N_A_145_409#_c_1721_n 6.23999e-19 $X=4.21 $Y=0.865
+ $X2=0 $Y2=0
cc_647 N_A_712_419#_c_663_n N_A_145_409#_c_1723_n 0.0246404f $X=4.21 $Y=0.865
+ $X2=0 $Y2=0
cc_648 N_A_712_419#_c_665_n N_A_145_409#_c_1723_n 0.00124673f $X=4.335 $Y=0.965
+ $X2=0 $Y2=0
cc_649 N_A_712_419#_c_684_n A_884_419# 0.00286141f $X=4.7 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_650 N_A_712_419#_c_667_n N_VGND_M1008_d 0.00764644f $X=5.345 $Y=0.95 $X2=0
+ $Y2=0
cc_651 N_A_712_419#_c_663_n N_VGND_c_1909_n 0.00670855f $X=4.21 $Y=0.865 $X2=0
+ $Y2=0
cc_652 N_A_712_419#_c_667_n N_VGND_c_1909_n 0.0176954f $X=5.345 $Y=0.95 $X2=0
+ $Y2=0
cc_653 N_A_712_419#_c_668_n N_VGND_c_1909_n 0.0182235f $X=5.43 $Y=0.865 $X2=0
+ $Y2=0
cc_654 N_A_712_419#_c_670_n N_VGND_c_1909_n 0.0140721f $X=5.515 $Y=0.35 $X2=0
+ $Y2=0
cc_655 N_A_712_419#_M1029_g N_VGND_c_1910_n 0.0131814f $X=7.13 $Y=0.835 $X2=0
+ $Y2=0
cc_656 N_A_712_419#_c_669_n N_VGND_c_1910_n 0.0106161f $X=6.3 $Y=0.35 $X2=0
+ $Y2=0
cc_657 N_A_712_419#_c_674_n N_VGND_c_1910_n 0.0233392f $X=6.385 $Y=1.245 $X2=0
+ $Y2=0
cc_658 N_A_712_419#_c_675_n N_VGND_c_1910_n 0.0100207f $X=6.875 $Y=1.33 $X2=0
+ $Y2=0
cc_659 N_A_712_419#_c_677_n N_VGND_c_1910_n 0.0172864f $X=7.04 $Y=1.41 $X2=0
+ $Y2=0
cc_660 N_A_712_419#_c_678_n N_VGND_c_1910_n 0.00139828f $X=7.04 $Y=1.41 $X2=0
+ $Y2=0
cc_661 N_A_712_419#_c_663_n N_VGND_c_1919_n 0.00844359f $X=4.21 $Y=0.865 $X2=0
+ $Y2=0
cc_662 N_A_712_419#_c_669_n N_VGND_c_1920_n 0.0589829f $X=6.3 $Y=0.35 $X2=0
+ $Y2=0
cc_663 N_A_712_419#_c_670_n N_VGND_c_1920_n 0.0114574f $X=5.515 $Y=0.35 $X2=0
+ $Y2=0
cc_664 N_A_712_419#_M1029_g N_VGND_c_1923_n 7.97988e-19 $X=7.13 $Y=0.835 $X2=0
+ $Y2=0
cc_665 N_A_712_419#_c_663_n N_VGND_c_1923_n 0.00771942f $X=4.21 $Y=0.865 $X2=0
+ $Y2=0
cc_666 N_A_712_419#_c_669_n N_VGND_c_1923_n 0.032098f $X=6.3 $Y=0.35 $X2=0 $Y2=0
cc_667 N_A_712_419#_c_670_n N_VGND_c_1923_n 0.00589978f $X=5.515 $Y=0.35 $X2=0
+ $Y2=0
cc_668 N_A_712_419#_c_767_n N_VGND_c_1923_n 0.00537264f $X=4.785 $Y=0.965 $X2=0
+ $Y2=0
cc_669 N_A_712_419#_c_664_n A_904_125# 0.00165482f $X=4.7 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_670 N_A_712_419#_c_674_n A_1249_125# 0.00292914f $X=6.385 $Y=1.245 $X2=-0.19
+ $Y2=-0.245
cc_671 N_SET_B_M1022_g N_A_263_409#_c_995_n 0.00907339f $X=6.56 $Y=0.835 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_862_n N_A_263_409#_c_1009_n 0.00556136f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_862_n N_A_263_409#_c_1010_n 0.00845492f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_862_n N_A_263_409#_c_1011_n 0.00107753f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_849_n N_A_1686_40#_M1039_g 0.0433565f $X=8.895 $Y=0.825 $X2=0
+ $Y2=0
cc_676 N_SET_B_c_851_n N_A_1686_40#_c_1191_n 0.0320355f $X=8.97 $Y=0.9 $X2=0
+ $Y2=0
cc_677 N_SET_B_c_852_n N_A_1686_40#_c_1191_n 0.00297689f $X=9.75 $Y=1.265 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_862_n N_A_1686_40#_c_1191_n 0.00201561f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_854_n N_A_1686_40#_c_1191_n 0.013005f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_680 N_SET_B_c_855_n N_A_1686_40#_c_1191_n 0.00234594f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_681 N_SET_B_c_861_n N_A_1686_40#_M1033_g 0.0299651f $X=9.75 $Y=1.935 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_862_n N_A_1686_40#_M1033_g 0.0115655f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_855_n N_A_1686_40#_M1033_g 0.00109739f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_684 N_SET_B_c_861_n N_A_1686_40#_c_1193_n 0.013005f $X=9.75 $Y=1.935 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_852_n N_A_1686_40#_c_1194_n 0.00465821f $X=9.75 $Y=1.265 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_862_n N_A_1686_40#_c_1194_n 0.00880383f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_854_n N_A_1686_40#_c_1194_n 0.00215461f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_688 N_SET_B_c_855_n N_A_1686_40#_c_1194_n 0.0388635f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_853_n N_A_1686_40#_c_1195_n 0.013005f $X=9.75 $Y=1.77 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_850_n N_A_1686_40#_c_1196_n 0.0199151f $X=9.615 $Y=0.9 $X2=0
+ $Y2=0
cc_691 N_SET_B_c_852_n N_A_1686_40#_c_1196_n 0.00580443f $X=9.75 $Y=1.265 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_855_n N_A_1686_40#_c_1196_n 0.0123704f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_693 N_SET_B_c_850_n N_A_1686_40#_c_1197_n 0.0107799f $X=9.615 $Y=0.9 $X2=0
+ $Y2=0
cc_694 N_SET_B_c_850_n N_A_1686_40#_c_1198_n 0.00564421f $X=9.615 $Y=0.9 $X2=0
+ $Y2=0
cc_695 N_SET_B_M1013_g N_A_1686_40#_c_1200_n 0.00600933f $X=9.71 $Y=2.595 $X2=0
+ $Y2=0
cc_696 N_SET_B_c_852_n N_A_1686_40#_c_1200_n 0.00275969f $X=9.75 $Y=1.265 $X2=0
+ $Y2=0
cc_697 SET_B N_A_1686_40#_c_1200_n 0.0064453f $X=9.755 $Y=1.95 $X2=0 $Y2=0
cc_698 N_SET_B_c_854_n N_A_1686_40#_c_1200_n 0.00274297f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_699 N_SET_B_c_855_n N_A_1686_40#_c_1200_n 0.0356517f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_850_n N_A_1686_40#_c_1201_n 0.00117215f $X=9.615 $Y=0.9 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_852_n N_A_1686_40#_c_1201_n 0.0024422f $X=9.75 $Y=1.265 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_854_n N_A_1686_40#_c_1201_n 0.00116535f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_703 N_SET_B_c_855_n N_A_1686_40#_c_1201_n 0.0171207f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_704 N_SET_B_c_862_n N_A_1519_125#_M1038_d 0.00598621f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_705 SET_B N_A_1519_125#_M1013_d 0.00138519f $X=9.755 $Y=1.95 $X2=0 $Y2=0
cc_706 N_SET_B_c_855_n N_A_1519_125#_M1013_d 8.58146e-19 $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_707 N_SET_B_c_850_n N_A_1519_125#_c_1289_n 0.00450356f $X=9.615 $Y=0.9 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_850_n N_A_1519_125#_c_1291_n 0.00196892f $X=9.615 $Y=0.9 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_851_n N_A_1519_125#_c_1307_n 0.00899895f $X=8.97 $Y=0.9 $X2=0
+ $Y2=0
cc_710 N_SET_B_c_852_n N_A_1519_125#_c_1307_n 3.25903e-19 $X=9.75 $Y=1.265 $X2=0
+ $Y2=0
cc_711 N_SET_B_c_862_n N_A_1519_125#_c_1331_n 0.0213707f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_712 N_SET_B_c_861_n N_A_1519_125#_c_1309_n 0.00158509f $X=9.75 $Y=1.935 $X2=0
+ $Y2=0
cc_713 N_SET_B_c_862_n N_A_1519_125#_c_1309_n 0.0244076f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_855_n N_A_1519_125#_c_1309_n 0.00413203f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_715 N_SET_B_M1013_g N_A_1519_125#_c_1351_n 0.0146858f $X=9.71 $Y=2.595 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_862_n N_A_1519_125#_c_1351_n 0.0232406f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_717 SET_B N_A_1519_125#_c_1351_n 8.13195e-19 $X=9.755 $Y=1.95 $X2=0 $Y2=0
cc_718 N_SET_B_c_855_n N_A_1519_125#_c_1351_n 0.0138025f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_719 N_SET_B_M1013_g N_A_1519_125#_c_1316_n 7.27872e-19 $X=9.71 $Y=2.595 $X2=0
+ $Y2=0
cc_720 N_SET_B_c_861_n N_A_1519_125#_c_1316_n 2.66149e-19 $X=9.75 $Y=1.935 $X2=0
+ $Y2=0
cc_721 SET_B N_A_1519_125#_c_1316_n 0.00289373f $X=9.755 $Y=1.95 $X2=0 $Y2=0
cc_722 N_SET_B_c_855_n N_A_1519_125#_c_1316_n 0.00678617f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_723 N_SET_B_M1013_g N_A_1519_125#_c_1317_n 0.00812382f $X=9.71 $Y=2.595 $X2=0
+ $Y2=0
cc_724 N_SET_B_M1013_g N_A_1519_125#_c_1319_n 0.00317906f $X=9.71 $Y=2.595 $X2=0
+ $Y2=0
cc_725 N_SET_B_c_862_n N_A_1519_125#_c_1321_n 0.0235822f $X=9.695 $Y=2.035 $X2=0
+ $Y2=0
cc_726 N_SET_B_c_852_n N_A_1519_125#_c_1311_n 0.00196892f $X=9.75 $Y=1.265 $X2=0
+ $Y2=0
cc_727 N_SET_B_c_854_n N_A_1519_125#_c_1311_n 0.0109681f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_728 N_SET_B_c_855_n N_A_1519_125#_c_1311_n 0.00230701f $X=9.75 $Y=1.43 $X2=0
+ $Y2=0
cc_729 N_SET_B_c_862_n N_VPWR_M1027_d 0.00304251f $X=9.695 $Y=2.035 $X2=0 $Y2=0
cc_730 N_SET_B_c_875_n N_VPWR_M1027_d 0.00132627f $X=6.625 $Y=2.035 $X2=0 $Y2=0
cc_731 N_SET_B_c_856_n N_VPWR_M1027_d 0.00262643f $X=6.5 $Y=1.77 $X2=0 $Y2=0
cc_732 N_SET_B_c_862_n N_VPWR_M1033_d 0.00382981f $X=9.695 $Y=2.035 $X2=0 $Y2=0
cc_733 N_SET_B_M1027_g N_VPWR_c_1579_n 0.00515373f $X=6.315 $Y=2.595 $X2=0 $Y2=0
cc_734 N_SET_B_M1013_g N_VPWR_c_1580_n 0.007692f $X=9.71 $Y=2.595 $X2=0 $Y2=0
cc_735 N_SET_B_M1027_g N_VPWR_c_1585_n 0.00713369f $X=6.315 $Y=2.595 $X2=0 $Y2=0
cc_736 N_SET_B_M1013_g N_VPWR_c_1589_n 0.00938036f $X=9.71 $Y=2.595 $X2=0 $Y2=0
cc_737 N_SET_B_M1027_g N_VPWR_c_1574_n 0.00942759f $X=6.315 $Y=2.595 $X2=0 $Y2=0
cc_738 N_SET_B_M1013_g N_VPWR_c_1574_n 0.0111949f $X=9.71 $Y=2.595 $X2=0 $Y2=0
cc_739 N_SET_B_c_862_n A_1441_419# 0.00218517f $X=9.695 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_740 N_SET_B_c_862_n A_1719_419# 0.00138626f $X=9.695 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_741 N_SET_B_M1022_g N_VGND_c_1910_n 0.00556619f $X=6.56 $Y=0.835 $X2=0 $Y2=0
cc_742 N_SET_B_c_849_n N_VGND_c_1911_n 0.0136022f $X=8.895 $Y=0.825 $X2=0 $Y2=0
cc_743 N_SET_B_c_850_n N_VGND_c_1911_n 0.00839872f $X=9.615 $Y=0.9 $X2=0 $Y2=0
cc_744 N_SET_B_c_849_n N_VGND_c_1917_n 0.00411131f $X=8.895 $Y=0.825 $X2=0 $Y2=0
cc_745 N_SET_B_M1022_g N_VGND_c_1923_n 9.49986e-19 $X=6.56 $Y=0.835 $X2=0 $Y2=0
cc_746 N_SET_B_c_849_n N_VGND_c_1923_n 0.00781653f $X=8.895 $Y=0.825 $X2=0 $Y2=0
cc_747 N_SET_B_c_850_n N_VGND_c_1923_n 0.0106417f $X=9.615 $Y=0.9 $X2=0 $Y2=0
cc_748 N_A_263_409#_c_995_n N_A_1686_40#_M1039_g 0.0243333f $X=7.955 $Y=0.18
+ $X2=0 $Y2=0
cc_749 N_A_263_409#_M1000_g N_A_1686_40#_c_1192_n 0.0243333f $X=8.03 $Y=0.835
+ $X2=0 $Y2=0
cc_750 N_A_263_409#_M1000_g N_A_1519_125#_c_1307_n 0.00294207f $X=8.03 $Y=0.835
+ $X2=0 $Y2=0
cc_751 N_A_263_409#_c_995_n N_A_1519_125#_c_1308_n 0.00414475f $X=7.955 $Y=0.18
+ $X2=0 $Y2=0
cc_752 N_A_263_409#_M1000_g N_A_1519_125#_c_1308_n 0.0180849f $X=8.03 $Y=0.835
+ $X2=0 $Y2=0
cc_753 N_A_263_409#_M1000_g N_A_1519_125#_c_1309_n 0.00290079f $X=8.03 $Y=0.835
+ $X2=0 $Y2=0
cc_754 N_A_263_409#_c_1009_n N_A_1519_125#_c_1321_n 0.018917f $X=7.57 $Y=2.02
+ $X2=0 $Y2=0
cc_755 N_A_263_409#_c_1010_n N_A_1519_125#_c_1321_n 0.0074013f $X=7.955 $Y=1.945
+ $X2=0 $Y2=0
cc_756 N_A_263_409#_c_1015_n N_VPWR_M1001_d 0.00180746f $X=2.13 $Y=2.045 $X2=0
+ $Y2=0
cc_757 N_A_263_409#_M1026_g N_VPWR_c_1577_n 0.0189086f $X=2.255 $Y=2.545 $X2=0
+ $Y2=0
cc_758 N_A_263_409#_c_1014_n N_VPWR_c_1577_n 0.0506352f $X=1.46 $Y=2.19 $X2=0
+ $Y2=0
cc_759 N_A_263_409#_c_1015_n N_VPWR_c_1577_n 0.0164812f $X=2.13 $Y=2.045 $X2=0
+ $Y2=0
cc_760 N_A_263_409#_c_1008_n N_VPWR_c_1578_n 0.00109287f $X=4.295 $Y=2.02 $X2=0
+ $Y2=0
cc_761 N_A_263_409#_c_1014_n N_VPWR_c_1583_n 0.0277632f $X=1.46 $Y=2.19 $X2=0
+ $Y2=0
cc_762 N_A_263_409#_M1026_g N_VPWR_c_1587_n 0.00767656f $X=2.255 $Y=2.545 $X2=0
+ $Y2=0
cc_763 N_A_263_409#_c_1008_n N_VPWR_c_1587_n 0.00599878f $X=4.295 $Y=2.02 $X2=0
+ $Y2=0
cc_764 N_A_263_409#_c_1009_n N_VPWR_c_1588_n 0.00828633f $X=7.57 $Y=2.02 $X2=0
+ $Y2=0
cc_765 N_A_263_409#_M1026_g N_VPWR_c_1574_n 0.014306f $X=2.255 $Y=2.545 $X2=0
+ $Y2=0
cc_766 N_A_263_409#_c_1008_n N_VPWR_c_1574_n 0.00876498f $X=4.295 $Y=2.02 $X2=0
+ $Y2=0
cc_767 N_A_263_409#_c_1009_n N_VPWR_c_1574_n 0.0132413f $X=7.57 $Y=2.02 $X2=0
+ $Y2=0
cc_768 N_A_263_409#_c_1014_n N_VPWR_c_1574_n 0.0158697f $X=1.46 $Y=2.19 $X2=0
+ $Y2=0
cc_769 N_A_263_409#_c_1014_n N_A_145_409#_c_1727_n 0.0760189f $X=1.46 $Y=2.19
+ $X2=0 $Y2=0
cc_770 N_A_263_409#_c_1000_n N_A_145_409#_c_1715_n 0.0296483f $X=1.295 $Y=1.075
+ $X2=0 $Y2=0
cc_771 N_A_263_409#_c_987_n N_A_145_409#_c_1716_n 6.98761e-19 $X=2.58 $Y=1.06
+ $X2=0 $Y2=0
cc_772 N_A_263_409#_c_1000_n N_A_145_409#_c_1716_n 0.0201676f $X=1.295 $Y=1.075
+ $X2=0 $Y2=0
cc_773 N_A_263_409#_c_988_n N_A_145_409#_c_1717_n 0.00755896f $X=2.58 $Y=1.555
+ $X2=0 $Y2=0
cc_774 N_A_263_409#_c_998_n N_A_145_409#_c_1717_n 0.00842211f $X=2.58 $Y=1.135
+ $X2=0 $Y2=0
cc_775 N_A_263_409#_c_1002_n N_A_145_409#_c_1717_n 0.0175365f $X=2.295 $Y=1.72
+ $X2=0 $Y2=0
cc_776 N_A_263_409#_c_1003_n N_A_145_409#_c_1717_n 0.00333091f $X=2.58 $Y=1.72
+ $X2=0 $Y2=0
cc_777 N_A_263_409#_c_1001_n N_A_145_409#_c_1718_n 0.00506527f $X=1.295 $Y=1.96
+ $X2=0 $Y2=0
cc_778 N_A_263_409#_c_987_n N_A_145_409#_c_1719_n 0.0108002f $X=2.58 $Y=1.06
+ $X2=0 $Y2=0
cc_779 N_A_263_409#_c_989_n N_A_145_409#_c_1719_n 0.00183437f $X=2.865 $Y=1.135
+ $X2=0 $Y2=0
cc_780 N_A_263_409#_c_990_n N_A_145_409#_c_1719_n 0.0047621f $X=2.94 $Y=1.06
+ $X2=0 $Y2=0
cc_781 N_A_263_409#_c_998_n N_A_145_409#_c_1719_n 6.70354e-19 $X=2.58 $Y=1.135
+ $X2=0 $Y2=0
cc_782 N_A_263_409#_M1026_g N_A_145_409#_c_1720_n 4.35785e-19 $X=2.255 $Y=2.545
+ $X2=0 $Y2=0
cc_783 N_A_263_409#_c_988_n N_A_145_409#_c_1720_n 0.0156171f $X=2.58 $Y=1.555
+ $X2=0 $Y2=0
cc_784 N_A_263_409#_c_1002_n N_A_145_409#_c_1720_n 0.0281451f $X=2.295 $Y=1.72
+ $X2=0 $Y2=0
cc_785 N_A_263_409#_c_1003_n N_A_145_409#_c_1720_n 0.00963292f $X=2.58 $Y=1.72
+ $X2=0 $Y2=0
cc_786 N_A_263_409#_c_990_n N_A_145_409#_c_1721_n 0.00707754f $X=2.94 $Y=1.06
+ $X2=0 $Y2=0
cc_787 N_A_263_409#_c_991_n N_A_145_409#_c_1721_n 0.00495317f $X=3.8 $Y=1.135
+ $X2=0 $Y2=0
cc_788 N_A_263_409#_M1020_g N_A_145_409#_c_1721_n 0.0119864f $X=3.89 $Y=0.655
+ $X2=0 $Y2=0
cc_789 N_A_263_409#_c_987_n N_A_145_409#_c_1722_n 2.48962e-19 $X=2.58 $Y=1.06
+ $X2=0 $Y2=0
cc_790 N_A_263_409#_M1026_g N_A_145_409#_c_1731_n 0.0010942f $X=2.255 $Y=2.545
+ $X2=0 $Y2=0
cc_791 N_A_263_409#_c_1015_n N_A_145_409#_c_1731_n 0.0150105f $X=2.13 $Y=2.045
+ $X2=0 $Y2=0
cc_792 N_A_263_409#_M1026_g N_A_145_409#_c_1732_n 0.00492177f $X=2.255 $Y=2.545
+ $X2=0 $Y2=0
cc_793 N_A_263_409#_c_990_n N_A_145_409#_c_1723_n 0.00472179f $X=2.94 $Y=1.06
+ $X2=0 $Y2=0
cc_794 N_A_263_409#_c_991_n N_A_145_409#_c_1723_n 0.00747149f $X=3.8 $Y=1.135
+ $X2=0 $Y2=0
cc_795 N_A_263_409#_c_992_n N_A_145_409#_c_1723_n 5.41301e-19 $X=3.875 $Y=1.21
+ $X2=0 $Y2=0
cc_796 N_A_263_409#_M1020_g N_A_145_409#_c_1723_n 0.00723319f $X=3.89 $Y=0.655
+ $X2=0 $Y2=0
cc_797 N_A_263_409#_c_1000_n N_A_145_409#_c_1724_n 0.0216895f $X=1.295 $Y=1.075
+ $X2=0 $Y2=0
cc_798 N_A_263_409#_c_1001_n N_A_145_409#_c_1724_n 0.0647658f $X=1.295 $Y=1.96
+ $X2=0 $Y2=0
cc_799 N_A_263_409#_c_1017_n N_A_145_409#_c_1724_n 0.0141548f $X=1.417 $Y=2.045
+ $X2=0 $Y2=0
cc_800 N_A_263_409#_c_1000_n N_A_145_409#_c_1725_n 0.00839784f $X=1.295 $Y=1.075
+ $X2=0 $Y2=0
cc_801 N_A_263_409#_c_988_n N_A_145_409#_c_1726_n 0.00111403f $X=2.58 $Y=1.555
+ $X2=0 $Y2=0
cc_802 N_A_263_409#_c_989_n N_A_145_409#_c_1726_n 0.00484021f $X=2.865 $Y=1.135
+ $X2=0 $Y2=0
cc_803 N_A_263_409#_c_987_n N_VGND_c_1908_n 9.43806e-19 $X=2.58 $Y=1.06 $X2=0
+ $Y2=0
cc_804 N_A_263_409#_c_995_n N_VGND_c_1909_n 0.0210695f $X=7.955 $Y=0.18 $X2=0
+ $Y2=0
cc_805 N_A_263_409#_c_995_n N_VGND_c_1910_n 0.0258253f $X=7.955 $Y=0.18 $X2=0
+ $Y2=0
cc_806 N_A_263_409#_c_995_n N_VGND_c_1917_n 0.0321435f $X=7.955 $Y=0.18 $X2=0
+ $Y2=0
cc_807 N_A_263_409#_c_987_n N_VGND_c_1919_n 0.00409299f $X=2.58 $Y=1.06 $X2=0
+ $Y2=0
cc_808 N_A_263_409#_c_996_n N_VGND_c_1919_n 0.036089f $X=3.965 $Y=0.18 $X2=0
+ $Y2=0
cc_809 N_A_263_409#_c_995_n N_VGND_c_1920_n 0.0390017f $X=7.955 $Y=0.18 $X2=0
+ $Y2=0
cc_810 N_A_263_409#_c_987_n N_VGND_c_1923_n 0.00437698f $X=2.58 $Y=1.06 $X2=0
+ $Y2=0
cc_811 N_A_263_409#_c_995_n N_VGND_c_1923_n 0.124122f $X=7.955 $Y=0.18 $X2=0
+ $Y2=0
cc_812 N_A_263_409#_c_996_n N_VGND_c_1923_n 0.0106778f $X=3.965 $Y=0.18 $X2=0
+ $Y2=0
cc_813 N_A_1686_40#_c_1198_n N_A_1519_125#_c_1287_n 0.0109596f $X=9.92 $Y=0.495
+ $X2=0 $Y2=0
cc_814 N_A_1686_40#_c_1199_n N_A_1519_125#_c_1288_n 0.0136954f $X=10.365 $Y=1
+ $X2=0 $Y2=0
cc_815 N_A_1686_40#_c_1198_n N_A_1519_125#_c_1289_n 0.00832939f $X=9.92 $Y=0.495
+ $X2=0 $Y2=0
cc_816 N_A_1686_40#_c_1199_n N_A_1519_125#_c_1289_n 0.0078115f $X=10.365 $Y=1
+ $X2=0 $Y2=0
cc_817 N_A_1686_40#_c_1201_n N_A_1519_125#_c_1289_n 6.58392e-19 $X=9.92 $Y=1
+ $X2=0 $Y2=0
cc_818 N_A_1686_40#_c_1198_n N_A_1519_125#_c_1290_n 0.00152289f $X=9.92 $Y=0.495
+ $X2=0 $Y2=0
cc_819 N_A_1686_40#_c_1199_n N_A_1519_125#_c_1291_n 0.00756497f $X=10.365 $Y=1
+ $X2=0 $Y2=0
cc_820 N_A_1686_40#_c_1200_n N_A_1519_125#_c_1291_n 0.00331326f $X=10.53
+ $Y=2.145 $X2=0 $Y2=0
cc_821 N_A_1686_40#_c_1200_n N_A_1519_125#_M1007_g 0.00425362f $X=10.53 $Y=2.145
+ $X2=0 $Y2=0
cc_822 N_A_1686_40#_c_1199_n N_A_1519_125#_c_1294_n 4.0175e-19 $X=10.365 $Y=1
+ $X2=0 $Y2=0
cc_823 N_A_1686_40#_c_1199_n N_A_1519_125#_c_1304_n 0.00718699f $X=10.365 $Y=1
+ $X2=0 $Y2=0
cc_824 N_A_1686_40#_M1039_g N_A_1519_125#_c_1307_n 0.0164657f $X=8.505 $Y=0.54
+ $X2=0 $Y2=0
cc_825 N_A_1686_40#_c_1191_n N_A_1519_125#_c_1307_n 0.00639996f $X=8.885 $Y=1.29
+ $X2=0 $Y2=0
cc_826 N_A_1686_40#_c_1197_n N_A_1519_125#_c_1307_n 0.0147435f $X=9.375 $Y=1
+ $X2=0 $Y2=0
cc_827 N_A_1686_40#_M1039_g N_A_1519_125#_c_1308_n 0.00183671f $X=8.505 $Y=0.54
+ $X2=0 $Y2=0
cc_828 N_A_1686_40#_M1039_g N_A_1519_125#_c_1309_n 0.00436911f $X=8.505 $Y=0.54
+ $X2=0 $Y2=0
cc_829 N_A_1686_40#_c_1191_n N_A_1519_125#_c_1309_n 0.0125962f $X=8.885 $Y=1.29
+ $X2=0 $Y2=0
cc_830 N_A_1686_40#_M1033_g N_A_1519_125#_c_1309_n 0.0127223f $X=9.01 $Y=2.595
+ $X2=0 $Y2=0
cc_831 N_A_1686_40#_c_1193_n N_A_1519_125#_c_1309_n 0.0057925f $X=9.13 $Y=1.885
+ $X2=0 $Y2=0
cc_832 N_A_1686_40#_c_1194_n N_A_1519_125#_c_1309_n 0.0544305f $X=9.21 $Y=1.38
+ $X2=0 $Y2=0
cc_833 N_A_1686_40#_c_1195_n N_A_1519_125#_c_1309_n 0.00908532f $X=9.21 $Y=1.38
+ $X2=0 $Y2=0
cc_834 N_A_1686_40#_M1033_g N_A_1519_125#_c_1351_n 0.0141446f $X=9.01 $Y=2.595
+ $X2=0 $Y2=0
cc_835 N_A_1686_40#_c_1193_n N_A_1519_125#_c_1351_n 0.00116124f $X=9.13 $Y=1.885
+ $X2=0 $Y2=0
cc_836 N_A_1686_40#_c_1194_n N_A_1519_125#_c_1351_n 0.00406247f $X=9.21 $Y=1.38
+ $X2=0 $Y2=0
cc_837 N_A_1686_40#_c_1200_n N_A_1519_125#_c_1316_n 0.0121086f $X=10.53 $Y=2.145
+ $X2=0 $Y2=0
cc_838 N_A_1686_40#_M1033_g N_A_1519_125#_c_1317_n 8.08161e-19 $X=9.01 $Y=2.595
+ $X2=0 $Y2=0
cc_839 N_A_1686_40#_c_1200_n N_A_1519_125#_c_1317_n 0.0143799f $X=10.53 $Y=2.145
+ $X2=0 $Y2=0
cc_840 N_A_1686_40#_M1007_s N_A_1519_125#_c_1318_n 0.00308696f $X=10.385 $Y=2
+ $X2=0 $Y2=0
cc_841 N_A_1686_40#_c_1200_n N_A_1519_125#_c_1318_n 0.0179944f $X=10.53 $Y=2.145
+ $X2=0 $Y2=0
cc_842 N_A_1686_40#_c_1200_n N_A_1519_125#_c_1310_n 0.0813762f $X=10.53 $Y=2.145
+ $X2=0 $Y2=0
cc_843 N_A_1686_40#_M1033_g N_A_1519_125#_c_1401_n 0.00401057f $X=9.01 $Y=2.595
+ $X2=0 $Y2=0
cc_844 N_A_1686_40#_c_1200_n N_A_1519_125#_c_1311_n 0.0329024f $X=10.53 $Y=2.145
+ $X2=0 $Y2=0
cc_845 N_A_1686_40#_M1033_g N_VPWR_c_1580_n 0.0144332f $X=9.01 $Y=2.595 $X2=0
+ $Y2=0
cc_846 N_A_1686_40#_M1033_g N_VPWR_c_1588_n 0.008763f $X=9.01 $Y=2.595 $X2=0
+ $Y2=0
cc_847 N_A_1686_40#_M1033_g N_VPWR_c_1574_n 0.0078527f $X=9.01 $Y=2.595 $X2=0
+ $Y2=0
cc_848 N_A_1686_40#_M1039_g N_VGND_c_1911_n 0.00279447f $X=8.505 $Y=0.54 $X2=0
+ $Y2=0
cc_849 N_A_1686_40#_c_1197_n N_VGND_c_1911_n 0.0137416f $X=9.375 $Y=1 $X2=0
+ $Y2=0
cc_850 N_A_1686_40#_c_1198_n N_VGND_c_1911_n 0.0190942f $X=9.92 $Y=0.495 $X2=0
+ $Y2=0
cc_851 N_A_1686_40#_c_1198_n N_VGND_c_1912_n 0.0153904f $X=9.92 $Y=0.495 $X2=0
+ $Y2=0
cc_852 N_A_1686_40#_c_1199_n N_VGND_c_1912_n 0.00575192f $X=10.365 $Y=1 $X2=0
+ $Y2=0
cc_853 N_A_1686_40#_M1039_g N_VGND_c_1917_n 0.00495161f $X=8.505 $Y=0.54 $X2=0
+ $Y2=0
cc_854 N_A_1686_40#_c_1198_n N_VGND_c_1921_n 0.0220321f $X=9.92 $Y=0.495 $X2=0
+ $Y2=0
cc_855 N_A_1686_40#_M1039_g N_VGND_c_1923_n 0.00983461f $X=8.505 $Y=0.54 $X2=0
+ $Y2=0
cc_856 N_A_1686_40#_c_1198_n N_VGND_c_1923_n 0.0125808f $X=9.92 $Y=0.495 $X2=0
+ $Y2=0
cc_857 N_A_1519_125#_c_1303_n N_A_2383_57#_M1040_g 0.0238263f $X=12.635 $Y=0.78
+ $X2=0 $Y2=0
cc_858 N_A_1519_125#_c_1306_n N_A_2383_57#_c_1509_n 0.0238263f $X=12.635
+ $Y=0.855 $X2=0 $Y2=0
cc_859 N_A_1519_125#_M1004_g N_A_2383_57#_c_1510_n 0.0238263f $X=12.585 $Y=2.37
+ $X2=0 $Y2=0
cc_860 N_A_1519_125#_c_1298_n N_A_2383_57#_c_1511_n 0.00243501f $X=11.545
+ $Y=1.17 $X2=0 $Y2=0
cc_861 N_A_1519_125#_c_1299_n N_A_2383_57#_c_1511_n 0.00701321f $X=12.2 $Y=0.855
+ $X2=0 $Y2=0
cc_862 N_A_1519_125#_c_1301_n N_A_2383_57#_c_1511_n 0.00192082f $X=12.275
+ $Y=0.78 $X2=0 $Y2=0
cc_863 N_A_1519_125#_M1004_g N_A_2383_57#_c_1511_n 0.0199796f $X=12.585 $Y=2.37
+ $X2=0 $Y2=0
cc_864 N_A_1519_125#_c_1306_n N_A_2383_57#_c_1511_n 0.00909497f $X=12.635
+ $Y=0.855 $X2=0 $Y2=0
cc_865 N_A_1519_125#_M1014_g N_A_2383_57#_c_1519_n 0.00272198f $X=11.495 $Y=2.5
+ $X2=0 $Y2=0
cc_866 N_A_1519_125#_M1004_g N_A_2383_57#_c_1519_n 0.0264529f $X=12.585 $Y=2.37
+ $X2=0 $Y2=0
cc_867 N_A_1519_125#_M1004_g N_A_2383_57#_c_1512_n 0.0245727f $X=12.585 $Y=2.37
+ $X2=0 $Y2=0
cc_868 N_A_1519_125#_M1004_g N_A_2383_57#_c_1513_n 0.00329386f $X=12.585 $Y=2.37
+ $X2=0 $Y2=0
cc_869 N_A_1519_125#_c_1296_n N_A_2383_57#_c_1515_n 9.77935e-19 $X=11.285
+ $Y=0.78 $X2=0 $Y2=0
cc_870 N_A_1519_125#_c_1299_n N_A_2383_57#_c_1515_n 0.00871991f $X=12.2 $Y=0.855
+ $X2=0 $Y2=0
cc_871 N_A_1519_125#_c_1301_n N_A_2383_57#_c_1515_n 0.0104516f $X=12.275 $Y=0.78
+ $X2=0 $Y2=0
cc_872 N_A_1519_125#_c_1303_n N_A_2383_57#_c_1515_n 0.00165639f $X=12.635
+ $Y=0.78 $X2=0 $Y2=0
cc_873 N_A_1519_125#_M1014_g N_A_2383_57#_c_1516_n 7.06177e-19 $X=11.495 $Y=2.5
+ $X2=0 $Y2=0
cc_874 N_A_1519_125#_M1004_g N_A_2383_57#_c_1516_n 0.00525478f $X=12.585 $Y=2.37
+ $X2=0 $Y2=0
cc_875 N_A_1519_125#_c_1306_n N_A_2383_57#_c_1516_n 0.00306103f $X=12.635
+ $Y=0.855 $X2=0 $Y2=0
cc_876 N_A_1519_125#_c_1351_n N_VPWR_M1033_d 0.00962408f $X=9.81 $Y=2.415 $X2=0
+ $Y2=0
cc_877 N_A_1519_125#_c_1351_n N_VPWR_c_1580_n 0.0197154f $X=9.81 $Y=2.415 $X2=0
+ $Y2=0
cc_878 N_A_1519_125#_c_1317_n N_VPWR_c_1580_n 0.0091605f $X=9.975 $Y=2.895 $X2=0
+ $Y2=0
cc_879 N_A_1519_125#_c_1319_n N_VPWR_c_1580_n 0.00767604f $X=10.14 $Y=2.98 $X2=0
+ $Y2=0
cc_880 N_A_1519_125#_M1007_g N_VPWR_c_1581_n 0.00481654f $X=10.795 $Y=2.5 $X2=0
+ $Y2=0
cc_881 N_A_1519_125#_c_1295_n N_VPWR_c_1581_n 0.00155013f $X=11.37 $Y=1.245
+ $X2=0 $Y2=0
cc_882 N_A_1519_125#_M1014_g N_VPWR_c_1581_n 0.0279424f $X=11.495 $Y=2.5 $X2=0
+ $Y2=0
cc_883 N_A_1519_125#_c_1318_n N_VPWR_c_1581_n 0.0092562f $X=10.795 $Y=2.98 $X2=0
+ $Y2=0
cc_884 N_A_1519_125#_M1004_g N_VPWR_c_1582_n 0.0257488f $X=12.585 $Y=2.37 $X2=0
+ $Y2=0
cc_885 N_A_1519_125#_c_1324_n N_VPWR_c_1588_n 0.0216692f $X=7.97 $Y=2.9 $X2=0
+ $Y2=0
cc_886 N_A_1519_125#_M1007_g N_VPWR_c_1589_n 0.00502067f $X=10.795 $Y=2.5 $X2=0
+ $Y2=0
cc_887 N_A_1519_125#_c_1318_n N_VPWR_c_1589_n 0.0503047f $X=10.795 $Y=2.98 $X2=0
+ $Y2=0
cc_888 N_A_1519_125#_c_1319_n N_VPWR_c_1589_n 0.0198962f $X=10.14 $Y=2.98 $X2=0
+ $Y2=0
cc_889 N_A_1519_125#_M1014_g N_VPWR_c_1590_n 0.00711337f $X=11.495 $Y=2.5 $X2=0
+ $Y2=0
cc_890 N_A_1519_125#_M1004_g N_VPWR_c_1590_n 0.00747382f $X=12.585 $Y=2.37 $X2=0
+ $Y2=0
cc_891 N_A_1519_125#_M1038_d N_VPWR_c_1574_n 0.0105425f $X=7.695 $Y=2.095 $X2=0
+ $Y2=0
cc_892 N_A_1519_125#_M1013_d N_VPWR_c_1574_n 0.00227987f $X=9.835 $Y=2.095 $X2=0
+ $Y2=0
cc_893 N_A_1519_125#_M1007_g N_VPWR_c_1574_n 0.00731936f $X=10.795 $Y=2.5 $X2=0
+ $Y2=0
cc_894 N_A_1519_125#_M1014_g N_VPWR_c_1574_n 0.0135914f $X=11.495 $Y=2.5 $X2=0
+ $Y2=0
cc_895 N_A_1519_125#_M1004_g N_VPWR_c_1574_n 0.00779694f $X=12.585 $Y=2.37 $X2=0
+ $Y2=0
cc_896 N_A_1519_125#_c_1324_n N_VPWR_c_1574_n 0.0126914f $X=7.97 $Y=2.9 $X2=0
+ $Y2=0
cc_897 N_A_1519_125#_c_1331_n N_VPWR_c_1574_n 0.0199763f $X=8.76 $Y=2.415 $X2=0
+ $Y2=0
cc_898 N_A_1519_125#_c_1351_n N_VPWR_c_1574_n 0.017375f $X=9.81 $Y=2.415 $X2=0
+ $Y2=0
cc_899 N_A_1519_125#_c_1318_n N_VPWR_c_1574_n 0.0298966f $X=10.795 $Y=2.98 $X2=0
+ $Y2=0
cc_900 N_A_1519_125#_c_1319_n N_VPWR_c_1574_n 0.0125808f $X=10.14 $Y=2.98 $X2=0
+ $Y2=0
cc_901 N_A_1519_125#_c_1401_n N_VPWR_c_1574_n 0.00637762f $X=8.845 $Y=2.415
+ $X2=0 $Y2=0
cc_902 N_A_1519_125#_c_1331_n A_1719_419# 0.00360016f $X=8.76 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_903 N_A_1519_125#_c_1309_n A_1719_419# 0.00316122f $X=8.845 $Y=2.33 $X2=-0.19
+ $Y2=-0.245
cc_904 N_A_1519_125#_c_1401_n A_1719_419# 0.00157762f $X=8.845 $Y=2.415
+ $X2=-0.19 $Y2=-0.245
cc_905 N_A_1519_125#_M1007_g N_Q_N_c_1847_n 3.25651e-19 $X=10.795 $Y=2.5 $X2=0
+ $Y2=0
cc_906 N_A_1519_125#_M1014_g N_Q_N_c_1847_n 0.0272278f $X=11.495 $Y=2.5 $X2=0
+ $Y2=0
cc_907 N_A_1519_125#_M1004_g N_Q_N_c_1847_n 0.00294351f $X=12.585 $Y=2.37 $X2=0
+ $Y2=0
cc_908 N_A_1519_125#_c_1320_n N_Q_N_c_1847_n 0.00465284f $X=10.88 $Y=2.895 $X2=0
+ $Y2=0
cc_909 N_A_1519_125#_c_1322_n N_Q_N_c_1847_n 0.00195406f $X=10.96 $Y=1.84 $X2=0
+ $Y2=0
cc_910 N_A_1519_125#_c_1292_n N_Q_N_c_1844_n 0.00125204f $X=10.925 $Y=0.78 $X2=0
+ $Y2=0
cc_911 N_A_1519_125#_c_1295_n N_Q_N_c_1844_n 4.94579e-19 $X=11.37 $Y=1.245 $X2=0
+ $Y2=0
cc_912 N_A_1519_125#_c_1296_n N_Q_N_c_1844_n 0.0093567f $X=11.285 $Y=0.78 $X2=0
+ $Y2=0
cc_913 N_A_1519_125#_c_1300_n N_Q_N_c_1844_n 0.00218345f $X=11.62 $Y=0.855 $X2=0
+ $Y2=0
cc_914 N_A_1519_125#_c_1301_n N_Q_N_c_1844_n 0.00122373f $X=12.275 $Y=0.78 $X2=0
+ $Y2=0
cc_915 N_A_1519_125#_M1014_g Q_N 0.0253748f $X=11.495 $Y=2.5 $X2=0 $Y2=0
cc_916 N_A_1519_125#_c_1299_n Q_N 0.00762733f $X=12.2 $Y=0.855 $X2=0 $Y2=0
cc_917 N_A_1519_125#_M1004_g Q_N 0.00283114f $X=12.585 $Y=2.37 $X2=0 $Y2=0
cc_918 N_A_1519_125#_c_1305_n Q_N 0.00751862f $X=11.495 $Y=1.245 $X2=0 $Y2=0
cc_919 N_A_1519_125#_c_1322_n Q_N 0.0124621f $X=10.96 $Y=1.84 $X2=0 $Y2=0
cc_920 N_A_1519_125#_c_1311_n Q_N 0.0016202f $X=11.125 $Y=1.505 $X2=0 $Y2=0
cc_921 N_A_1519_125#_c_1296_n N_Q_N_c_1846_n 0.00192025f $X=11.285 $Y=0.78 $X2=0
+ $Y2=0
cc_922 N_A_1519_125#_c_1298_n N_Q_N_c_1846_n 0.0163993f $X=11.545 $Y=1.17 $X2=0
+ $Y2=0
cc_923 N_A_1519_125#_c_1299_n N_Q_N_c_1846_n 0.00504367f $X=12.2 $Y=0.855 $X2=0
+ $Y2=0
cc_924 N_A_1519_125#_c_1300_n N_Q_N_c_1846_n 0.0109715f $X=11.62 $Y=0.855 $X2=0
+ $Y2=0
cc_925 N_A_1519_125#_c_1305_n N_Q_N_c_1846_n 4.27513e-19 $X=11.495 $Y=1.245
+ $X2=0 $Y2=0
cc_926 N_A_1519_125#_c_1310_n N_Q_N_c_1846_n 0.0124621f $X=10.96 $Y=1.335 $X2=0
+ $Y2=0
cc_927 N_A_1519_125#_M1004_g N_Q_c_1886_n 2.74877e-19 $X=12.585 $Y=2.37 $X2=0
+ $Y2=0
cc_928 N_A_1519_125#_c_1308_n N_VGND_c_1910_n 0.00710794f $X=8.095 $Y=1 $X2=0
+ $Y2=0
cc_929 N_A_1519_125#_c_1287_n N_VGND_c_1912_n 0.002112f $X=10.135 $Y=0.78 $X2=0
+ $Y2=0
cc_930 N_A_1519_125#_c_1290_n N_VGND_c_1912_n 0.0125929f $X=10.495 $Y=0.78 $X2=0
+ $Y2=0
cc_931 N_A_1519_125#_c_1292_n N_VGND_c_1912_n 0.012598f $X=10.925 $Y=0.78 $X2=0
+ $Y2=0
cc_932 N_A_1519_125#_c_1296_n N_VGND_c_1912_n 0.002112f $X=11.285 $Y=0.78 $X2=0
+ $Y2=0
cc_933 N_A_1519_125#_c_1310_n N_VGND_c_1912_n 0.00326237f $X=10.96 $Y=1.335
+ $X2=0 $Y2=0
cc_934 N_A_1519_125#_c_1311_n N_VGND_c_1912_n 0.00531303f $X=11.125 $Y=1.505
+ $X2=0 $Y2=0
cc_935 N_A_1519_125#_c_1292_n N_VGND_c_1913_n 0.00445056f $X=10.925 $Y=0.78
+ $X2=0 $Y2=0
cc_936 N_A_1519_125#_c_1293_n N_VGND_c_1913_n 4.57848e-19 $X=11.21 $Y=0.855
+ $X2=0 $Y2=0
cc_937 N_A_1519_125#_c_1296_n N_VGND_c_1913_n 0.00502664f $X=11.285 $Y=0.78
+ $X2=0 $Y2=0
cc_938 N_A_1519_125#_c_1299_n N_VGND_c_1913_n 0.00384753f $X=12.2 $Y=0.855 $X2=0
+ $Y2=0
cc_939 N_A_1519_125#_c_1300_n N_VGND_c_1913_n 3.90485e-19 $X=11.62 $Y=0.855
+ $X2=0 $Y2=0
cc_940 N_A_1519_125#_c_1301_n N_VGND_c_1913_n 0.00433172f $X=12.275 $Y=0.78
+ $X2=0 $Y2=0
cc_941 N_A_1519_125#_c_1303_n N_VGND_c_1913_n 0.00445056f $X=12.635 $Y=0.78
+ $X2=0 $Y2=0
cc_942 N_A_1519_125#_c_1306_n N_VGND_c_1913_n 5.84996e-19 $X=12.635 $Y=0.855
+ $X2=0 $Y2=0
cc_943 N_A_1519_125#_c_1301_n N_VGND_c_1914_n 0.00207566f $X=12.275 $Y=0.78
+ $X2=0 $Y2=0
cc_944 N_A_1519_125#_c_1303_n N_VGND_c_1914_n 0.0130071f $X=12.635 $Y=0.78 $X2=0
+ $Y2=0
cc_945 N_A_1519_125#_c_1308_n N_VGND_c_1917_n 0.0090144f $X=8.095 $Y=1 $X2=0
+ $Y2=0
cc_946 N_A_1519_125#_c_1287_n N_VGND_c_1921_n 0.00502664f $X=10.135 $Y=0.78
+ $X2=0 $Y2=0
cc_947 N_A_1519_125#_c_1288_n N_VGND_c_1921_n 4.57848e-19 $X=10.42 $Y=0.855
+ $X2=0 $Y2=0
cc_948 N_A_1519_125#_c_1290_n N_VGND_c_1921_n 0.00445056f $X=10.495 $Y=0.78
+ $X2=0 $Y2=0
cc_949 N_A_1519_125#_c_1287_n N_VGND_c_1923_n 0.010303f $X=10.135 $Y=0.78 $X2=0
+ $Y2=0
cc_950 N_A_1519_125#_c_1288_n N_VGND_c_1923_n 6.33118e-19 $X=10.42 $Y=0.855
+ $X2=0 $Y2=0
cc_951 N_A_1519_125#_c_1290_n N_VGND_c_1923_n 0.00796275f $X=10.495 $Y=0.78
+ $X2=0 $Y2=0
cc_952 N_A_1519_125#_c_1292_n N_VGND_c_1923_n 0.00796275f $X=10.925 $Y=0.78
+ $X2=0 $Y2=0
cc_953 N_A_1519_125#_c_1293_n N_VGND_c_1923_n 6.33118e-19 $X=11.21 $Y=0.855
+ $X2=0 $Y2=0
cc_954 N_A_1519_125#_c_1296_n N_VGND_c_1923_n 0.010303f $X=11.285 $Y=0.78 $X2=0
+ $Y2=0
cc_955 N_A_1519_125#_c_1300_n N_VGND_c_1923_n 0.00516662f $X=11.62 $Y=0.855
+ $X2=0 $Y2=0
cc_956 N_A_1519_125#_c_1301_n N_VGND_c_1923_n 0.0084505f $X=12.275 $Y=0.78 $X2=0
+ $Y2=0
cc_957 N_A_1519_125#_c_1303_n N_VGND_c_1923_n 0.00796275f $X=12.635 $Y=0.78
+ $X2=0 $Y2=0
cc_958 N_A_1519_125#_c_1306_n N_VGND_c_1923_n 7.94744e-19 $X=12.635 $Y=0.855
+ $X2=0 $Y2=0
cc_959 N_A_1519_125#_c_1308_n N_VGND_c_1923_n 0.011636f $X=8.095 $Y=1 $X2=0
+ $Y2=0
cc_960 N_A_1519_125#_c_1307_n A_1621_125# 0.00736402f $X=8.76 $Y=1 $X2=-0.19
+ $Y2=-0.245
cc_961 N_A_2383_57#_M1030_g N_VPWR_c_1582_n 0.0257478f $X=13.115 $Y=2.37 $X2=0
+ $Y2=0
cc_962 N_A_2383_57#_c_1519_n N_VPWR_c_1582_n 0.0692741f $X=12.32 $Y=2.015 $X2=0
+ $Y2=0
cc_963 N_A_2383_57#_c_1512_n N_VPWR_c_1582_n 0.0253501f $X=12.99 $Y=1.575 $X2=0
+ $Y2=0
cc_964 N_A_2383_57#_c_1519_n N_VPWR_c_1590_n 0.0122968f $X=12.32 $Y=2.015 $X2=0
+ $Y2=0
cc_965 N_A_2383_57#_M1030_g N_VPWR_c_1591_n 0.00747382f $X=13.115 $Y=2.37 $X2=0
+ $Y2=0
cc_966 N_A_2383_57#_M1030_g N_VPWR_c_1574_n 0.00779694f $X=13.115 $Y=2.37 $X2=0
+ $Y2=0
cc_967 N_A_2383_57#_c_1519_n N_VPWR_c_1574_n 0.0131561f $X=12.32 $Y=2.015 $X2=0
+ $Y2=0
cc_968 N_A_2383_57#_c_1515_n N_Q_N_c_1844_n 0.0313468f $X=12.06 $Y=0.495 $X2=0
+ $Y2=0
cc_969 N_A_2383_57#_c_1511_n Q_N 0.0240775f $X=12.19 $Y=1.49 $X2=0 $Y2=0
cc_970 N_A_2383_57#_c_1519_n Q_N 0.0995518f $X=12.32 $Y=2.015 $X2=0 $Y2=0
cc_971 N_A_2383_57#_c_1515_n Q_N 0.00127638f $X=12.06 $Y=0.495 $X2=0 $Y2=0
cc_972 N_A_2383_57#_c_1516_n Q_N 0.0147194f $X=12.295 $Y=1.575 $X2=0 $Y2=0
cc_973 N_A_2383_57#_c_1511_n N_Q_N_c_1846_n 0.0165535f $X=12.19 $Y=1.49 $X2=0
+ $Y2=0
cc_974 N_A_2383_57#_M1040_g N_Q_c_1883_n 0.00125204f $X=13.065 $Y=0.495 $X2=0
+ $Y2=0
cc_975 N_A_2383_57#_M1031_g N_Q_c_1883_n 0.0100348f $X=13.425 $Y=0.495 $X2=0
+ $Y2=0
cc_976 N_A_2383_57#_M1030_g Q 0.0134647f $X=13.115 $Y=2.37 $X2=0 $Y2=0
cc_977 N_A_2383_57#_M1030_g N_Q_c_1886_n 0.00585731f $X=13.115 $Y=2.37 $X2=0
+ $Y2=0
cc_978 N_A_2383_57#_c_1510_n N_Q_c_1886_n 6.17296e-19 $X=13.155 $Y=1.66 $X2=0
+ $Y2=0
cc_979 N_A_2383_57#_c_1512_n N_Q_c_1886_n 0.00840259f $X=12.99 $Y=1.575 $X2=0
+ $Y2=0
cc_980 N_A_2383_57#_M1030_g N_Q_c_1884_n 0.00399218f $X=13.115 $Y=2.37 $X2=0
+ $Y2=0
cc_981 N_A_2383_57#_M1031_g N_Q_c_1884_n 0.0117228f $X=13.425 $Y=0.495 $X2=0
+ $Y2=0
cc_982 N_A_2383_57#_c_1512_n N_Q_c_1884_n 0.00851731f $X=12.99 $Y=1.575 $X2=0
+ $Y2=0
cc_983 N_A_2383_57#_c_1513_n N_Q_c_1884_n 0.0236709f $X=13.155 $Y=1.155 $X2=0
+ $Y2=0
cc_984 N_A_2383_57#_c_1514_n N_Q_c_1884_n 0.00811515f $X=13.155 $Y=1.155 $X2=0
+ $Y2=0
cc_985 N_A_2383_57#_c_1515_n N_VGND_c_1913_n 0.0248255f $X=12.06 $Y=0.495 $X2=0
+ $Y2=0
cc_986 N_A_2383_57#_M1040_g N_VGND_c_1914_n 0.0125983f $X=13.065 $Y=0.495 $X2=0
+ $Y2=0
cc_987 N_A_2383_57#_M1031_g N_VGND_c_1914_n 0.002112f $X=13.425 $Y=0.495 $X2=0
+ $Y2=0
cc_988 N_A_2383_57#_c_1513_n N_VGND_c_1914_n 0.00135938f $X=13.155 $Y=1.155
+ $X2=0 $Y2=0
cc_989 N_A_2383_57#_c_1515_n N_VGND_c_1914_n 0.0171525f $X=12.06 $Y=0.495 $X2=0
+ $Y2=0
cc_990 N_A_2383_57#_M1040_g N_VGND_c_1922_n 0.00445056f $X=13.065 $Y=0.495 $X2=0
+ $Y2=0
cc_991 N_A_2383_57#_M1031_g N_VGND_c_1922_n 0.00502664f $X=13.425 $Y=0.495 $X2=0
+ $Y2=0
cc_992 N_A_2383_57#_M1040_g N_VGND_c_1923_n 0.00796275f $X=13.065 $Y=0.495 $X2=0
+ $Y2=0
cc_993 N_A_2383_57#_M1031_g N_VGND_c_1923_n 0.0100616f $X=13.425 $Y=0.495 $X2=0
+ $Y2=0
cc_994 N_A_2383_57#_c_1515_n N_VGND_c_1923_n 0.0142018f $X=12.06 $Y=0.495 $X2=0
+ $Y2=0
cc_995 N_VPWR_c_1574_n N_A_145_409#_M1005_s 0.00233022f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_996 N_VPWR_c_1576_n N_A_145_409#_c_1727_n 0.0684934f $X=0.335 $Y=2.19 $X2=0
+ $Y2=0
cc_997 N_VPWR_c_1583_n N_A_145_409#_c_1728_n 0.0220321f $X=1.825 $Y=3.33 $X2=0
+ $Y2=0
cc_998 N_VPWR_c_1574_n N_A_145_409#_c_1728_n 0.0125808f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_999 N_VPWR_c_1574_n A_884_419# 0.00356886f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1000 N_VPWR_c_1574_n A_1441_419# 0.00286f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1001 N_VPWR_c_1574_n A_1719_419# 0.00421038f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1002 N_VPWR_c_1581_n N_Q_N_c_1847_n 0.0645184f $X=11.23 $Y=2.185 $X2=0 $Y2=0
cc_1003 N_VPWR_c_1590_n N_Q_N_c_1847_n 0.0173442f $X=12.685 $Y=3.33 $X2=0 $Y2=0
cc_1004 N_VPWR_c_1574_n N_Q_N_c_1847_n 0.0122839f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1005 N_VPWR_c_1591_n Q 0.0191637f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1006 N_VPWR_c_1574_n Q 0.0204781f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_1007 N_VPWR_c_1582_n N_Q_c_1886_n 0.071673f $X=12.85 $Y=2.015 $X2=0 $Y2=0
cc_1008 N_A_145_409#_c_1725_n N_VGND_c_1907_n 0.0162324f $X=1.037 $Y=0.35 $X2=0
+ $Y2=0
cc_1009 N_A_145_409#_c_1715_n N_VGND_c_1908_n 0.0132716f $X=1.92 $Y=0.35 $X2=0
+ $Y2=0
cc_1010 N_A_145_409#_c_1716_n N_VGND_c_1908_n 0.0194919f $X=2.005 $Y=1.1 $X2=0
+ $Y2=0
cc_1011 N_A_145_409#_c_1717_n N_VGND_c_1908_n 0.013238f $X=2.64 $Y=1.185 $X2=0
+ $Y2=0
cc_1012 N_A_145_409#_c_1719_n N_VGND_c_1908_n 0.0194919f $X=2.725 $Y=1.1 $X2=0
+ $Y2=0
cc_1013 N_A_145_409#_c_1722_n N_VGND_c_1908_n 0.0132716f $X=2.81 $Y=0.35 $X2=0
+ $Y2=0
cc_1014 N_A_145_409#_c_1715_n N_VGND_c_1915_n 0.0541822f $X=1.92 $Y=0.35 $X2=0
+ $Y2=0
cc_1015 N_A_145_409#_c_1725_n N_VGND_c_1915_n 0.0232749f $X=1.037 $Y=0.35 $X2=0
+ $Y2=0
cc_1016 N_A_145_409#_c_1721_n N_VGND_c_1919_n 0.0644006f $X=3.51 $Y=0.35 $X2=0
+ $Y2=0
cc_1017 N_A_145_409#_c_1722_n N_VGND_c_1919_n 0.0114622f $X=2.81 $Y=0.35 $X2=0
+ $Y2=0
cc_1018 N_A_145_409#_c_1715_n N_VGND_c_1923_n 0.0329217f $X=1.92 $Y=0.35 $X2=0
+ $Y2=0
cc_1019 N_A_145_409#_c_1721_n N_VGND_c_1923_n 0.0387747f $X=3.51 $Y=0.35 $X2=0
+ $Y2=0
cc_1020 N_A_145_409#_c_1722_n N_VGND_c_1923_n 0.00657784f $X=2.81 $Y=0.35 $X2=0
+ $Y2=0
cc_1021 N_A_145_409#_c_1725_n N_VGND_c_1923_n 0.0133596f $X=1.037 $Y=0.35 $X2=0
+ $Y2=0
cc_1022 N_Q_N_c_1844_n N_VGND_c_1912_n 0.0153904f $X=11.5 $Y=0.495 $X2=0 $Y2=0
cc_1023 N_Q_N_c_1844_n N_VGND_c_1913_n 0.0217285f $X=11.5 $Y=0.495 $X2=0 $Y2=0
cc_1024 N_Q_N_c_1844_n N_VGND_c_1923_n 0.0125175f $X=11.5 $Y=0.495 $X2=0 $Y2=0
cc_1025 N_Q_c_1883_n N_VGND_c_1914_n 0.0153904f $X=13.64 $Y=0.495 $X2=0 $Y2=0
cc_1026 N_Q_c_1883_n N_VGND_c_1922_n 0.0217285f $X=13.64 $Y=0.495 $X2=0 $Y2=0
cc_1027 N_Q_c_1883_n N_VGND_c_1923_n 0.0125175f $X=13.64 $Y=0.495 $X2=0 $Y2=0
