* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or3b_lp A B C_N VGND VNB VPB VPWR X
X0 a_114_47# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_47# C_N a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_27_47# a_272_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_350_47# A a_640_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_640_101# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_27_47# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_804_101# a_350_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_263_373# B a_628_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_466_185# B a_350_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_350_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VGND a_350_47# a_804_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_628_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_272_47# a_27_47# a_350_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_263_373# a_27_47# a_350_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VGND B a_466_185# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
