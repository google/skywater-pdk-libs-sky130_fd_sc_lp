* File: sky130_fd_sc_lp__maj3_0.spice
* Created: Wed Sep  2 09:59:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__maj3_0.pex.spice"
.subckt sky130_fd_sc_lp__maj3_0  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 A_149_57# N_C_M1000_g N_A_28_431#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g A_149_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1001 A_313_57# N_A_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_28_431#_M1002_d N_B_M1002_g A_313_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1007 A_477_57# N_B_M1007_g N_A_28_431#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_C_M1011_g A_477_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_28_431#_M1003_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1013 A_115_431# N_C_M1013_g N_A_28_431#_M1013_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g A_115_431# VPB PHIGHVT L=0.15 W=0.42 AD=0.1071
+ AS=0.0441 PD=0.93 PS=0.63 NRD=53.9386 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1008 A_319_431# N_A_M1008_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.1071 PD=0.63 PS=0.93 NRD=23.443 NRS=53.9386 M=1 R=2.8 SA=75001.2 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_28_431#_M1006_d N_B_M1006_g A_319_431# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.6
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1004 A_477_431# N_B_M1004_g N_A_28_431#_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75002
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_C_M1005_g A_477_431# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0914094 AS=0.0441 PD=0.824151 PS=0.63 NRD=56.2829 NRS=23.443 M=1 R=2.8
+ SA=75002.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_28_431#_M1009_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.256 AS=0.139291 PD=2.08 PS=1.25585 NRD=35.3812 NRS=0 M=1 R=4.26667
+ SA=75002 SB=75000.3 A=0.096 P=1.58 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__maj3_0.pxi.spice"
*
.ends
*
*
