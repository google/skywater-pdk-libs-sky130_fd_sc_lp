* File: sky130_fd_sc_lp__dlrbp_lp.pxi.spice
* Created: Fri Aug 28 10:26:18 2020
* 
x_PM_SKY130_FD_SC_LP__DLRBP_LP%D N_D_M1014_g N_D_M1027_g N_D_M1006_g N_D_c_196_n
+ N_D_c_197_n D D N_D_c_199_n PM_SKY130_FD_SC_LP__DLRBP_LP%D
x_PM_SKY130_FD_SC_LP__DLRBP_LP%GATE N_GATE_M1013_g N_GATE_M1008_g N_GATE_M1000_g
+ N_GATE_c_236_n N_GATE_c_241_n GATE GATE N_GATE_c_238_n
+ PM_SKY130_FD_SC_LP__DLRBP_LP%GATE
x_PM_SKY130_FD_SC_LP__DLRBP_LP%A_272_419# N_A_272_419#_M1000_d
+ N_A_272_419#_M1013_d N_A_272_419#_M1016_g N_A_272_419#_M1011_g
+ N_A_272_419#_M1010_g N_A_272_419#_M1007_g N_A_272_419#_M1019_g
+ N_A_272_419#_c_297_n N_A_272_419#_c_285_n N_A_272_419#_c_299_n
+ N_A_272_419#_c_286_n N_A_272_419#_c_322_p N_A_272_419#_c_287_n
+ N_A_272_419#_c_288_n N_A_272_419#_c_302_n N_A_272_419#_c_303_n
+ N_A_272_419#_c_304_n N_A_272_419#_c_289_n N_A_272_419#_c_306_n
+ N_A_272_419#_c_290_n N_A_272_419#_c_307_n N_A_272_419#_c_291_n
+ N_A_272_419#_c_292_n N_A_272_419#_c_293_n N_A_272_419#_c_294_n
+ PM_SKY130_FD_SC_LP__DLRBP_LP%A_272_419#
x_PM_SKY130_FD_SC_LP__DLRBP_LP%A_27_112# N_A_27_112#_M1014_s N_A_27_112#_M1027_s
+ N_A_27_112#_c_447_n N_A_27_112#_c_448_n N_A_27_112#_M1025_g
+ N_A_27_112#_M1018_g N_A_27_112#_c_443_n N_A_27_112#_c_444_n
+ N_A_27_112#_c_451_n N_A_27_112#_c_452_n N_A_27_112#_c_453_n
+ N_A_27_112#_c_445_n N_A_27_112#_c_454_n N_A_27_112#_c_446_n
+ PM_SKY130_FD_SC_LP__DLRBP_LP%A_27_112#
x_PM_SKY130_FD_SC_LP__DLRBP_LP%A_455_49# N_A_455_49#_M1016_s N_A_455_49#_M1011_s
+ N_A_455_49#_M1026_g N_A_455_49#_c_527_n N_A_455_49#_c_528_n
+ N_A_455_49#_c_529_n N_A_455_49#_c_530_n N_A_455_49#_M1009_g
+ N_A_455_49#_c_531_n N_A_455_49#_c_532_n N_A_455_49#_c_533_n
+ N_A_455_49#_c_542_n N_A_455_49#_c_534_n N_A_455_49#_c_535_n
+ N_A_455_49#_c_536_n N_A_455_49#_c_537_n PM_SKY130_FD_SC_LP__DLRBP_LP%A_455_49#
x_PM_SKY130_FD_SC_LP__DLRBP_LP%A_1028_23# N_A_1028_23#_M1020_s
+ N_A_1028_23#_M1021_d N_A_1028_23#_M1028_g N_A_1028_23#_M1002_g
+ N_A_1028_23#_M1003_g N_A_1028_23#_M1005_g N_A_1028_23#_M1024_g
+ N_A_1028_23#_c_624_n N_A_1028_23#_c_625_n N_A_1028_23#_c_626_n
+ N_A_1028_23#_M1029_g N_A_1028_23#_M1004_g N_A_1028_23#_c_628_n
+ N_A_1028_23#_M1001_g N_A_1028_23#_c_629_n N_A_1028_23#_c_630_n
+ N_A_1028_23#_c_631_n N_A_1028_23#_c_632_n N_A_1028_23#_c_645_n
+ N_A_1028_23#_c_646_n N_A_1028_23#_c_647_n N_A_1028_23#_c_633_n
+ N_A_1028_23#_c_648_n N_A_1028_23#_c_634_n N_A_1028_23#_c_635_n
+ N_A_1028_23#_c_636_n N_A_1028_23#_c_637_n N_A_1028_23#_c_650_n
+ N_A_1028_23#_c_638_n PM_SKY130_FD_SC_LP__DLRBP_LP%A_1028_23#
x_PM_SKY130_FD_SC_LP__DLRBP_LP%A_778_49# N_A_778_49#_M1026_d N_A_778_49#_M1007_d
+ N_A_778_49#_M1021_g N_A_778_49#_c_790_n N_A_778_49#_c_791_n
+ N_A_778_49#_M1020_g N_A_778_49#_c_793_n N_A_778_49#_c_804_n
+ N_A_778_49#_c_794_n N_A_778_49#_c_795_n N_A_778_49#_c_796_n
+ N_A_778_49#_c_797_n N_A_778_49#_c_798_n N_A_778_49#_c_799_n
+ N_A_778_49#_c_800_n N_A_778_49#_c_801_n PM_SKY130_FD_SC_LP__DLRBP_LP%A_778_49#
x_PM_SKY130_FD_SC_LP__DLRBP_LP%RESET_B N_RESET_B_M1015_g N_RESET_B_M1023_g
+ N_RESET_B_c_893_n N_RESET_B_c_894_n N_RESET_B_c_895_n N_RESET_B_c_891_n
+ N_RESET_B_c_897_n RESET_B RESET_B RESET_B N_RESET_B_c_899_n
+ PM_SKY130_FD_SC_LP__DLRBP_LP%RESET_B
x_PM_SKY130_FD_SC_LP__DLRBP_LP%A_1614_74# N_A_1614_74#_M1029_s
+ N_A_1614_74#_M1004_s N_A_1614_74#_M1017_g N_A_1614_74#_M1022_g
+ N_A_1614_74#_M1012_g N_A_1614_74#_c_943_n N_A_1614_74#_c_944_n
+ N_A_1614_74#_c_945_n N_A_1614_74#_c_946_n N_A_1614_74#_c_947_n
+ N_A_1614_74#_c_948_n N_A_1614_74#_c_949_n N_A_1614_74#_c_950_n
+ PM_SKY130_FD_SC_LP__DLRBP_LP%A_1614_74#
x_PM_SKY130_FD_SC_LP__DLRBP_LP%VPWR N_VPWR_M1027_d N_VPWR_M1011_d N_VPWR_M1002_d
+ N_VPWR_M1015_d N_VPWR_M1004_d N_VPWR_c_1005_n N_VPWR_c_1006_n N_VPWR_c_1007_n
+ N_VPWR_c_1008_n N_VPWR_c_1009_n N_VPWR_c_1010_n N_VPWR_c_1011_n
+ N_VPWR_c_1012_n N_VPWR_c_1013_n VPWR N_VPWR_c_1014_n N_VPWR_c_1015_n
+ N_VPWR_c_1016_n N_VPWR_c_1017_n N_VPWR_c_1004_n N_VPWR_c_1019_n
+ N_VPWR_c_1020_n N_VPWR_c_1021_n PM_SKY130_FD_SC_LP__DLRBP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DLRBP_LP%Q N_Q_M1024_d N_Q_M1003_d N_Q_c_1114_n
+ N_Q_c_1112_n N_Q_c_1113_n Q Q Q PM_SKY130_FD_SC_LP__DLRBP_LP%Q
x_PM_SKY130_FD_SC_LP__DLRBP_LP%Q_N N_Q_N_M1012_d N_Q_N_M1022_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1151_n PM_SKY130_FD_SC_LP__DLRBP_LP%Q_N
x_PM_SKY130_FD_SC_LP__DLRBP_LP%VGND N_VGND_M1006_d N_VGND_M1010_d N_VGND_M1028_d
+ N_VGND_M1023_d N_VGND_M1001_d N_VGND_c_1169_n N_VGND_c_1170_n N_VGND_c_1171_n
+ N_VGND_c_1172_n N_VGND_c_1173_n N_VGND_c_1174_n N_VGND_c_1175_n VGND
+ N_VGND_c_1176_n N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n
+ N_VGND_c_1180_n N_VGND_c_1181_n N_VGND_c_1182_n N_VGND_c_1183_n
+ N_VGND_c_1184_n N_VGND_c_1185_n PM_SKY130_FD_SC_LP__DLRBP_LP%VGND
cc_1 VNB N_D_M1014_g 0.0258512f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.77
cc_2 VNB N_D_M1006_g 0.0197639f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.77
cc_3 VNB N_D_c_196_n 0.0209367f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.33
cc_4 VNB N_D_c_197_n 8.47018e-19 $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.85
cc_5 VNB D 0.00372538f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_D_c_199_n 0.0265117f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.345
cc_7 VNB N_GATE_M1008_g 0.019763f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.595
cc_8 VNB N_GATE_M1000_g 0.0225937f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.33
cc_9 VNB N_GATE_c_236_n 0.0209917f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.33
cc_10 VNB GATE 0.00580494f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.85
cc_11 VNB N_GATE_c_238_n 0.0247575f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.345
cc_12 VNB N_A_272_419#_M1016_g 0.0385512f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.18
cc_13 VNB N_A_272_419#_M1011_g 0.00201031f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.33
cc_14 VNB N_A_272_419#_M1010_g 0.0311821f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.85
cc_15 VNB N_A_272_419#_M1019_g 0.0259676f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.295
cc_16 VNB N_A_272_419#_c_285_n 0.0136059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_272_419#_c_286_n 2.86674e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_272_419#_c_287_n 0.00566592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_272_419#_c_288_n 0.00361034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_272_419#_c_289_n 0.00458574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_272_419#_c_290_n 0.0129885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_272_419#_c_291_n 0.0128062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_272_419#_c_292_n 0.00338023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_272_419#_c_293_n 0.0348968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_272_419#_c_294_n 0.0394172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_112#_M1018_g 0.0232695f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.85
cc_27 VNB N_A_27_112#_c_443_n 0.0251144f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_28 VNB N_A_27_112#_c_444_n 0.0102048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_112#_c_445_n 0.0263877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_112#_c_446_n 0.0307989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_455_49#_c_527_n 0.0269744f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.77
cc_32 VNB N_A_455_49#_c_528_n 0.0256726f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.33
cc_33 VNB N_A_455_49#_c_529_n 0.0166722f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.18
cc_34 VNB N_A_455_49#_c_530_n 0.00196635f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.33
cc_35 VNB N_A_455_49#_c_531_n 0.0106837f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.345
cc_36 VNB N_A_455_49#_c_532_n 0.0114273f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.295
cc_37 VNB N_A_455_49#_c_533_n 0.00769386f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.665
cc_38 VNB N_A_455_49#_c_534_n 0.00304656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_455_49#_c_535_n 0.0321157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_455_49#_c_536_n 0.0171242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_455_49#_c_537_n 0.01889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1028_23#_M1028_g 0.0559366f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.18
cc_43 VNB N_A_1028_23#_M1005_g 0.019756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1028_23#_M1024_g 0.024576f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.295
cc_45 VNB N_A_1028_23#_c_624_n 0.0647644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1028_23#_c_625_n 0.0200864f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.665
cc_47 VNB N_A_1028_23#_c_626_n 0.0174644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1028_23#_M1004_g 0.0466586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1028_23#_c_628_n 0.01411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1028_23#_c_629_n 0.00922328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1028_23#_c_630_n 0.0170774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1028_23#_c_631_n 0.00211689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1028_23#_c_632_n 0.0166613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1028_23#_c_633_n 0.00800005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1028_23#_c_634_n 0.0146979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1028_23#_c_635_n 0.00102481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1028_23#_c_636_n 0.0266809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1028_23#_c_637_n 0.00660298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1028_23#_c_638_n 8.15863e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_778_49#_c_790_n 0.0203806f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.77
cc_61 VNB N_A_778_49#_c_791_n 0.0173699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_778_49#_M1020_g 0.0271258f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.33
cc_63 VNB N_A_778_49#_c_793_n 0.0094023f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_64 VNB N_A_778_49#_c_794_n 0.00797567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_778_49#_c_795_n 0.00200591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_778_49#_c_796_n 0.0182288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_778_49#_c_797_n 0.00343203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_778_49#_c_798_n 0.00975234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_778_49#_c_799_n 0.00691179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_778_49#_c_800_n 0.00546617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_778_49#_c_801_n 0.0300992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_RESET_B_M1023_g 0.0484191f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.595
cc_73 VNB N_RESET_B_c_891_n 0.0123096f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.18
cc_74 VNB N_A_1614_74#_M1017_g 0.0202979f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.18
cc_75 VNB N_A_1614_74#_M1012_g 0.0250777f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.85
cc_76 VNB N_A_1614_74#_c_943_n 0.0245507f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.345
cc_77 VNB N_A_1614_74#_c_944_n 0.0128053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1614_74#_c_945_n 0.00752635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1614_74#_c_946_n 0.021225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1614_74#_c_947_n 0.0121926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1614_74#_c_948_n 0.0118388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1614_74#_c_949_n 0.00142556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1614_74#_c_950_n 0.028193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VPWR_c_1004_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_Q_c_1112_n 0.0207239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_Q_c_1113_n 0.00668943f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.18
cc_87 VNB Q_N 0.0229441f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.595
cc_88 VNB Q_N 0.0430852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1169_n 0.0272649f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_90 VNB N_VGND_c_1170_n 0.0517644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1171_n 7.46595e-19 $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.345
cc_92 VNB N_VGND_c_1172_n 0.0123624f $X=-0.19 $Y=-0.245 $X2=0.667 $Y2=1.665
cc_93 VNB N_VGND_c_1173_n 0.00977238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1174_n 0.0503917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1175_n 0.00664583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1176_n 0.0291794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1177_n 0.0573607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1178_n 0.0273224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1179_n 0.028381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1180_n 0.542804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1181_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1182_n 0.00449123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1183_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1184_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1185_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VPB N_D_M1027_g 0.0365954f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.595
cc_107 VPB N_D_c_197_n 0.0204226f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.85
cc_108 VPB D 0.00225823f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_109 VPB N_GATE_M1013_g 0.0349256f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.77
cc_110 VPB N_GATE_c_236_n 0.0041927f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.33
cc_111 VPB N_GATE_c_241_n 0.0286408f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.645
cc_112 VPB GATE 0.00510958f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.85
cc_113 VPB N_A_272_419#_M1011_g 0.0268374f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.33
cc_114 VPB N_A_272_419#_M1007_g 0.0242948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_272_419#_c_297_n 0.00801535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_272_419#_c_285_n 0.0128498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_272_419#_c_299_n 0.0165963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_272_419#_c_287_n 0.0175976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_272_419#_c_288_n 0.00133768f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_272_419#_c_302_n 0.00427271f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_272_419#_c_303_n 0.0197426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_272_419#_c_304_n 0.00393773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_272_419#_c_289_n 0.00288813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_272_419#_c_306_n 0.00314224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_272_419#_c_307_n 0.00225528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_272_419#_c_291_n 0.0132055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_27_112#_c_447_n 0.0983434f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.595
cc_128 VPB N_A_27_112#_c_448_n 0.0107704f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.18
cc_129 VPB N_A_27_112#_M1025_g 0.0157983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_27_112#_c_443_n 0.00982688f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_131 VPB N_A_27_112#_c_451_n 0.0102056f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.345
cc_132 VPB N_A_27_112#_c_452_n 0.00130908f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.665
cc_133 VPB N_A_27_112#_c_453_n 0.0620527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_27_112#_c_454_n 0.0536844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_27_112#_c_446_n 0.02041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_455_49#_c_529_n 0.00968557f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.18
cc_137 VPB N_A_455_49#_c_530_n 0.00718554f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.33
cc_138 VPB N_A_455_49#_M1009_g 0.0333518f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_139 VPB N_A_455_49#_c_532_n 0.0040104f $X=-0.19 $Y=1.655 $X2=0.667 $Y2=1.295
cc_140 VPB N_A_455_49#_c_542_n 0.010301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_1028_23#_M1002_g 0.0246358f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.33
cc_142 VPB N_A_1028_23#_M1003_g 0.0260756f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.85
cc_143 VPB N_A_1028_23#_M1004_g 0.0317243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_1028_23#_c_629_n 0.00525472f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_1028_23#_c_631_n 4.28226e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_1028_23#_c_632_n 0.015829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_1028_23#_c_645_n 0.00854148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_1028_23#_c_646_n 9.08934e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_1028_23#_c_647_n 0.0053507f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_1028_23#_c_648_n 0.00343771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_1028_23#_c_634_n 0.00410174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_1028_23#_c_650_n 0.00369126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_1028_23#_c_638_n 2.51035e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_778_49#_M1021_g 0.0359489f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.18
cc_155 VPB N_A_778_49#_c_793_n 0.00525575f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_156 VPB N_A_778_49#_c_804_n 0.00320365f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.345
cc_157 VPB N_A_778_49#_c_798_n 0.00357502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_778_49#_c_800_n 7.55834e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_RESET_B_M1015_g 0.042217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_c_893_n 0.0915238f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.18
cc_161 VPB N_RESET_B_c_894_n 0.0176343f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.77
cc_162 VPB N_RESET_B_c_895_n 0.0183783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_RESET_B_c_891_n 0.00396925f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.18
cc_164 VPB N_RESET_B_c_897_n 0.0198149f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.645
cc_165 VPB RESET_B 0.0211467f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.85
cc_166 VPB N_RESET_B_c_899_n 0.054623f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.345
cc_167 VPB N_A_1614_74#_M1022_g 0.0329914f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.33
cc_168 VPB N_A_1614_74#_c_944_n 0.00265483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_1614_74#_c_946_n 0.0217623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_1614_74#_c_949_n 7.69351e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1005_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_172 VPB N_VPWR_c_1006_n 0.0117269f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.345
cc_173 VPB N_VPWR_c_1007_n 0.0145629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1008_n 0.0101157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1009_n 0.0226092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1010_n 0.0213315f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1011_n 0.00436154f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1012_n 0.0262049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1013_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1014_n 0.0483255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1015_n 0.0555299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1016_n 0.0516141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1017_n 0.027252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1004_n 0.118553f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1019_n 0.00473485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1020_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1021_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_Q_c_1114_n 0.0152261f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.77
cc_189 VPB N_Q_c_1112_n 0.010972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB Q 0.0155221f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.85
cc_191 VPB Q_N 0.0107983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB Q_N 0.043146f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_Q_N_c_1151_n 0.0256541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 N_D_M1027_g N_GATE_M1013_g 0.0285821f $X=0.705 $Y=2.595 $X2=0 $Y2=0
cc_195 N_D_M1006_g N_GATE_M1008_g 0.0119294f $X=0.855 $Y=0.77 $X2=0 $Y2=0
cc_196 N_D_c_197_n N_GATE_c_236_n 0.00555375f $X=0.625 $Y=1.85 $X2=0 $Y2=0
cc_197 N_D_c_197_n N_GATE_c_241_n 0.0285821f $X=0.625 $Y=1.85 $X2=0 $Y2=0
cc_198 D N_GATE_c_241_n 5.43316e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_199 N_D_c_196_n GATE 0.00132304f $X=0.675 $Y=1.33 $X2=0 $Y2=0
cc_200 D GATE 0.0439882f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_201 N_D_c_199_n GATE 0.00227004f $X=0.665 $Y=1.345 $X2=0 $Y2=0
cc_202 N_D_c_196_n N_GATE_c_238_n 0.0119294f $X=0.675 $Y=1.33 $X2=0 $Y2=0
cc_203 D N_GATE_c_238_n 0.00128705f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_204 N_D_c_199_n N_GATE_c_238_n 0.00555375f $X=0.665 $Y=1.345 $X2=0 $Y2=0
cc_205 N_D_M1027_g N_A_272_419#_c_306_n 0.00110445f $X=0.705 $Y=2.595 $X2=0
+ $Y2=0
cc_206 N_D_M1027_g N_A_27_112#_c_451_n 0.0174967f $X=0.705 $Y=2.595 $X2=0 $Y2=0
cc_207 D N_A_27_112#_c_451_n 0.00553203f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_208 N_D_M1014_g N_A_27_112#_c_445_n 0.0102796f $X=0.495 $Y=0.77 $X2=0 $Y2=0
cc_209 N_D_M1006_g N_A_27_112#_c_445_n 0.00125204f $X=0.855 $Y=0.77 $X2=0 $Y2=0
cc_210 N_D_M1027_g N_A_27_112#_c_454_n 0.024464f $X=0.705 $Y=2.595 $X2=0 $Y2=0
cc_211 N_D_c_197_n N_A_27_112#_c_454_n 0.00429185f $X=0.625 $Y=1.85 $X2=0 $Y2=0
cc_212 D N_A_27_112#_c_454_n 0.00731237f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_213 N_D_M1014_g N_A_27_112#_c_446_n 0.0214749f $X=0.495 $Y=0.77 $X2=0 $Y2=0
cc_214 N_D_M1027_g N_A_27_112#_c_446_n 0.0055452f $X=0.705 $Y=2.595 $X2=0 $Y2=0
cc_215 D N_A_27_112#_c_446_n 0.042203f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_216 N_D_M1027_g N_VPWR_c_1005_n 0.00990743f $X=0.705 $Y=2.595 $X2=0 $Y2=0
cc_217 N_D_M1027_g N_VPWR_c_1010_n 0.00629498f $X=0.705 $Y=2.595 $X2=0 $Y2=0
cc_218 N_D_M1027_g N_VPWR_c_1004_n 0.00798245f $X=0.705 $Y=2.595 $X2=0 $Y2=0
cc_219 N_D_M1014_g N_VGND_c_1169_n 0.00180376f $X=0.495 $Y=0.77 $X2=0 $Y2=0
cc_220 N_D_M1006_g N_VGND_c_1169_n 0.0130197f $X=0.855 $Y=0.77 $X2=0 $Y2=0
cc_221 N_D_M1014_g N_VGND_c_1176_n 0.0043356f $X=0.495 $Y=0.77 $X2=0 $Y2=0
cc_222 N_D_M1006_g N_VGND_c_1176_n 0.00375057f $X=0.855 $Y=0.77 $X2=0 $Y2=0
cc_223 N_D_M1014_g N_VGND_c_1180_n 0.00487769f $X=0.495 $Y=0.77 $X2=0 $Y2=0
cc_224 N_D_M1006_g N_VGND_c_1180_n 0.00409726f $X=0.855 $Y=0.77 $X2=0 $Y2=0
cc_225 N_GATE_c_241_n N_A_272_419#_c_297_n 0.00168779f $X=1.415 $Y=1.85 $X2=0
+ $Y2=0
cc_226 GATE N_A_272_419#_c_297_n 4.2716e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_227 N_GATE_M1013_g N_A_272_419#_c_285_n 0.00598512f $X=1.235 $Y=2.595 $X2=0
+ $Y2=0
cc_228 N_GATE_M1000_g N_A_272_419#_c_285_n 0.0236714f $X=1.645 $Y=0.77 $X2=0
+ $Y2=0
cc_229 GATE N_A_272_419#_c_285_n 0.0503813f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_230 N_GATE_M1013_g N_A_272_419#_c_306_n 0.00663217f $X=1.235 $Y=2.595 $X2=0
+ $Y2=0
cc_231 N_GATE_c_241_n N_A_272_419#_c_306_n 0.00208181f $X=1.415 $Y=1.85 $X2=0
+ $Y2=0
cc_232 GATE N_A_272_419#_c_306_n 0.0218921f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_233 N_GATE_M1008_g N_A_272_419#_c_290_n 0.00125204f $X=1.285 $Y=0.77 $X2=0
+ $Y2=0
cc_234 N_GATE_M1000_g N_A_272_419#_c_290_n 0.0102796f $X=1.645 $Y=0.77 $X2=0
+ $Y2=0
cc_235 N_GATE_M1013_g N_A_27_112#_c_451_n 0.0223973f $X=1.235 $Y=2.595 $X2=0
+ $Y2=0
cc_236 GATE N_A_27_112#_c_451_n 0.00589011f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_237 N_GATE_M1013_g N_A_27_112#_c_452_n 0.00335737f $X=1.235 $Y=2.595 $X2=0
+ $Y2=0
cc_238 N_GATE_M1013_g N_A_27_112#_c_453_n 0.0124741f $X=1.235 $Y=2.595 $X2=0
+ $Y2=0
cc_239 N_GATE_M1013_g N_A_27_112#_c_454_n 0.00249613f $X=1.235 $Y=2.595 $X2=0
+ $Y2=0
cc_240 N_GATE_M1000_g N_A_455_49#_c_531_n 0.00328677f $X=1.645 $Y=0.77 $X2=0
+ $Y2=0
cc_241 N_GATE_M1013_g N_VPWR_c_1005_n 0.0106066f $X=1.235 $Y=2.595 $X2=0 $Y2=0
cc_242 N_GATE_M1013_g N_VPWR_c_1014_n 0.00639129f $X=1.235 $Y=2.595 $X2=0 $Y2=0
cc_243 N_GATE_M1013_g N_VPWR_c_1004_n 0.00775836f $X=1.235 $Y=2.595 $X2=0 $Y2=0
cc_244 N_GATE_M1008_g N_VGND_c_1169_n 0.0122426f $X=1.285 $Y=0.77 $X2=0 $Y2=0
cc_245 N_GATE_M1000_g N_VGND_c_1169_n 0.00180376f $X=1.645 $Y=0.77 $X2=0 $Y2=0
cc_246 N_GATE_c_241_n N_VGND_c_1169_n 2.87206e-19 $X=1.415 $Y=1.85 $X2=0 $Y2=0
cc_247 GATE N_VGND_c_1169_n 0.0130791f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_248 N_GATE_M1008_g N_VGND_c_1170_n 0.00375057f $X=1.285 $Y=0.77 $X2=0 $Y2=0
cc_249 N_GATE_M1000_g N_VGND_c_1170_n 0.0043356f $X=1.645 $Y=0.77 $X2=0 $Y2=0
cc_250 N_GATE_M1008_g N_VGND_c_1180_n 0.00409726f $X=1.285 $Y=0.77 $X2=0 $Y2=0
cc_251 N_GATE_M1000_g N_VGND_c_1180_n 0.00487769f $X=1.645 $Y=0.77 $X2=0 $Y2=0
cc_252 N_A_272_419#_M1011_g N_A_27_112#_c_447_n 0.0152142f $X=2.725 $Y=2.175
+ $X2=0 $Y2=0
cc_253 N_A_272_419#_M1011_g N_A_27_112#_c_448_n 0.030133f $X=2.725 $Y=2.175
+ $X2=0 $Y2=0
cc_254 N_A_272_419#_c_322_p N_A_27_112#_c_448_n 0.00932134f $X=2.89 $Y=2.165
+ $X2=0 $Y2=0
cc_255 N_A_272_419#_c_287_n N_A_27_112#_c_448_n 0.00516995f $X=3.67 $Y=1.51
+ $X2=0 $Y2=0
cc_256 N_A_272_419#_c_299_n N_A_27_112#_M1025_g 0.00454006f $X=2.805 $Y=2.25
+ $X2=0 $Y2=0
cc_257 N_A_272_419#_c_304_n N_A_27_112#_M1025_g 0.00322161f $X=4 $Y=2.98 $X2=0
+ $Y2=0
cc_258 N_A_272_419#_M1010_g N_A_27_112#_M1018_g 0.0223531f $X=2.995 $Y=0.455
+ $X2=0 $Y2=0
cc_259 N_A_272_419#_M1011_g N_A_27_112#_c_443_n 0.00527654f $X=2.725 $Y=2.175
+ $X2=0 $Y2=0
cc_260 N_A_272_419#_M1007_g N_A_27_112#_c_443_n 0.0668746f $X=3.825 $Y=2.335
+ $X2=0 $Y2=0
cc_261 N_A_272_419#_c_286_n N_A_27_112#_c_443_n 0.00110736f $X=2.89 $Y=1.675
+ $X2=0 $Y2=0
cc_262 N_A_272_419#_c_322_p N_A_27_112#_c_443_n 5.3184e-19 $X=2.89 $Y=2.165
+ $X2=0 $Y2=0
cc_263 N_A_272_419#_c_287_n N_A_27_112#_c_443_n 0.0226472f $X=3.67 $Y=1.51 $X2=0
+ $Y2=0
cc_264 N_A_272_419#_c_302_n N_A_27_112#_c_443_n 0.00704244f $X=3.835 $Y=2.895
+ $X2=0 $Y2=0
cc_265 N_A_272_419#_c_291_n N_A_27_112#_c_443_n 0.0213276f $X=3.835 $Y=1.51
+ $X2=0 $Y2=0
cc_266 N_A_272_419#_c_294_n N_A_27_112#_c_443_n 0.0146132f $X=2.995 $Y=1.3 $X2=0
+ $Y2=0
cc_267 N_A_272_419#_M1010_g N_A_27_112#_c_444_n 0.0146132f $X=2.995 $Y=0.455
+ $X2=0 $Y2=0
cc_268 N_A_272_419#_c_287_n N_A_27_112#_c_444_n 0.0010845f $X=3.67 $Y=1.51 $X2=0
+ $Y2=0
cc_269 N_A_272_419#_M1013_d N_A_27_112#_c_451_n 0.00729992f $X=1.36 $Y=2.095
+ $X2=0 $Y2=0
cc_270 N_A_272_419#_M1011_g N_A_27_112#_c_451_n 0.00549535f $X=2.725 $Y=2.175
+ $X2=0 $Y2=0
cc_271 N_A_272_419#_c_297_n N_A_27_112#_c_451_n 0.002356f $X=1.855 $Y=2.25 $X2=0
+ $Y2=0
cc_272 N_A_272_419#_c_299_n N_A_27_112#_c_451_n 0.0103256f $X=2.805 $Y=2.25
+ $X2=0 $Y2=0
cc_273 N_A_272_419#_c_306_n N_A_27_112#_c_451_n 0.0310262f $X=1.665 $Y=2.205
+ $X2=0 $Y2=0
cc_274 N_A_272_419#_c_307_n N_A_27_112#_c_451_n 0.0149615f $X=1.94 $Y=2.25 $X2=0
+ $Y2=0
cc_275 N_A_272_419#_M1011_g N_A_27_112#_c_452_n 0.00186695f $X=2.725 $Y=2.175
+ $X2=0 $Y2=0
cc_276 N_A_272_419#_M1011_g N_A_27_112#_c_453_n 0.00213425f $X=2.725 $Y=2.175
+ $X2=0 $Y2=0
cc_277 N_A_272_419#_c_299_n N_A_27_112#_c_453_n 5.41696e-19 $X=2.805 $Y=2.25
+ $X2=0 $Y2=0
cc_278 N_A_272_419#_c_307_n N_A_27_112#_c_453_n 8.11211e-19 $X=1.94 $Y=2.25
+ $X2=0 $Y2=0
cc_279 N_A_272_419#_c_299_n N_A_455_49#_M1011_s 0.0121642f $X=2.805 $Y=2.25
+ $X2=0 $Y2=0
cc_280 N_A_272_419#_c_292_n N_A_455_49#_c_527_n 2.8257e-19 $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_281 N_A_272_419#_c_293_n N_A_455_49#_c_527_n 0.0150044f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_282 N_A_272_419#_c_288_n N_A_455_49#_c_528_n 8.51879e-19 $X=3.835 $Y=1.675
+ $X2=0 $Y2=0
cc_283 N_A_272_419#_c_289_n N_A_455_49#_c_528_n 0.00138519f $X=4.815 $Y=2.895
+ $X2=0 $Y2=0
cc_284 N_A_272_419#_c_291_n N_A_455_49#_c_528_n 0.0151486f $X=3.835 $Y=1.51
+ $X2=0 $Y2=0
cc_285 N_A_272_419#_c_289_n N_A_455_49#_c_529_n 0.00536378f $X=4.815 $Y=2.895
+ $X2=0 $Y2=0
cc_286 N_A_272_419#_c_292_n N_A_455_49#_c_529_n 0.00120658f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_287 N_A_272_419#_c_293_n N_A_455_49#_c_529_n 0.0116031f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_288 N_A_272_419#_M1007_g N_A_455_49#_M1009_g 0.0134653f $X=3.825 $Y=2.335
+ $X2=0 $Y2=0
cc_289 N_A_272_419#_c_302_n N_A_455_49#_M1009_g 0.00163057f $X=3.835 $Y=2.895
+ $X2=0 $Y2=0
cc_290 N_A_272_419#_c_303_n N_A_455_49#_M1009_g 0.0166036f $X=4.73 $Y=2.98 $X2=0
+ $Y2=0
cc_291 N_A_272_419#_c_289_n N_A_455_49#_M1009_g 0.0374806f $X=4.815 $Y=2.895
+ $X2=0 $Y2=0
cc_292 N_A_272_419#_c_291_n N_A_455_49#_M1009_g 0.00145282f $X=3.835 $Y=1.51
+ $X2=0 $Y2=0
cc_293 N_A_272_419#_M1016_g N_A_455_49#_c_531_n 0.0114161f $X=2.635 $Y=0.455
+ $X2=0 $Y2=0
cc_294 N_A_272_419#_M1010_g N_A_455_49#_c_531_n 0.0018251f $X=2.995 $Y=0.455
+ $X2=0 $Y2=0
cc_295 N_A_272_419#_c_290_n N_A_455_49#_c_531_n 0.0164838f $X=1.86 $Y=0.77 $X2=0
+ $Y2=0
cc_296 N_A_272_419#_M1016_g N_A_455_49#_c_532_n 0.0150008f $X=2.635 $Y=0.455
+ $X2=0 $Y2=0
cc_297 N_A_272_419#_M1011_g N_A_455_49#_c_532_n 0.0044138f $X=2.725 $Y=2.175
+ $X2=0 $Y2=0
cc_298 N_A_272_419#_c_286_n N_A_455_49#_c_532_n 0.0292025f $X=2.89 $Y=1.675
+ $X2=0 $Y2=0
cc_299 N_A_272_419#_c_290_n N_A_455_49#_c_532_n 0.0427608f $X=1.86 $Y=0.77 $X2=0
+ $Y2=0
cc_300 N_A_272_419#_M1016_g N_A_455_49#_c_533_n 0.00501003f $X=2.635 $Y=0.455
+ $X2=0 $Y2=0
cc_301 N_A_272_419#_c_290_n N_A_455_49#_c_533_n 0.0121616f $X=1.86 $Y=0.77 $X2=0
+ $Y2=0
cc_302 N_A_272_419#_M1011_g N_A_455_49#_c_542_n 0.00725407f $X=2.725 $Y=2.175
+ $X2=0 $Y2=0
cc_303 N_A_272_419#_c_285_n N_A_455_49#_c_542_n 0.0213217f $X=1.94 $Y=2.165
+ $X2=0 $Y2=0
cc_304 N_A_272_419#_c_299_n N_A_455_49#_c_542_n 0.0228981f $X=2.805 $Y=2.25
+ $X2=0 $Y2=0
cc_305 N_A_272_419#_c_286_n N_A_455_49#_c_542_n 0.00146755f $X=2.89 $Y=1.675
+ $X2=0 $Y2=0
cc_306 N_A_272_419#_c_322_p N_A_455_49#_c_542_n 0.0213455f $X=2.89 $Y=2.165
+ $X2=0 $Y2=0
cc_307 N_A_272_419#_c_294_n N_A_455_49#_c_542_n 0.00173673f $X=2.995 $Y=1.3
+ $X2=0 $Y2=0
cc_308 N_A_272_419#_c_288_n N_A_455_49#_c_534_n 0.0175491f $X=3.835 $Y=1.675
+ $X2=0 $Y2=0
cc_309 N_A_272_419#_c_291_n N_A_455_49#_c_534_n 3.67923e-19 $X=3.835 $Y=1.51
+ $X2=0 $Y2=0
cc_310 N_A_272_419#_M1019_g N_A_455_49#_c_535_n 0.00288312f $X=4.645 $Y=0.455
+ $X2=0 $Y2=0
cc_311 N_A_272_419#_c_288_n N_A_455_49#_c_535_n 0.00115457f $X=3.835 $Y=1.675
+ $X2=0 $Y2=0
cc_312 N_A_272_419#_c_291_n N_A_455_49#_c_535_n 0.0160177f $X=3.835 $Y=1.51
+ $X2=0 $Y2=0
cc_313 N_A_272_419#_M1016_g N_A_455_49#_c_536_n 0.00974192f $X=2.635 $Y=0.455
+ $X2=0 $Y2=0
cc_314 N_A_272_419#_M1010_g N_A_455_49#_c_536_n 0.0117997f $X=2.995 $Y=0.455
+ $X2=0 $Y2=0
cc_315 N_A_272_419#_c_286_n N_A_455_49#_c_536_n 0.0241297f $X=2.89 $Y=1.675
+ $X2=0 $Y2=0
cc_316 N_A_272_419#_c_287_n N_A_455_49#_c_536_n 0.0290215f $X=3.67 $Y=1.51 $X2=0
+ $Y2=0
cc_317 N_A_272_419#_c_288_n N_A_455_49#_c_536_n 0.00168948f $X=3.835 $Y=1.675
+ $X2=0 $Y2=0
cc_318 N_A_272_419#_c_291_n N_A_455_49#_c_536_n 2.31103e-19 $X=3.835 $Y=1.51
+ $X2=0 $Y2=0
cc_319 N_A_272_419#_c_294_n N_A_455_49#_c_536_n 2.06137e-19 $X=2.995 $Y=1.3
+ $X2=0 $Y2=0
cc_320 N_A_272_419#_M1019_g N_A_455_49#_c_537_n 0.00564444f $X=4.645 $Y=0.455
+ $X2=0 $Y2=0
cc_321 N_A_272_419#_M1019_g N_A_1028_23#_M1028_g 0.0211033f $X=4.645 $Y=0.455
+ $X2=0 $Y2=0
cc_322 N_A_272_419#_c_289_n N_A_1028_23#_M1028_g 0.00861415f $X=4.815 $Y=2.895
+ $X2=0 $Y2=0
cc_323 N_A_272_419#_c_292_n N_A_1028_23#_M1028_g 0.00123098f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_324 N_A_272_419#_c_293_n N_A_1028_23#_M1028_g 0.0178736f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_325 N_A_272_419#_c_303_n N_A_1028_23#_M1002_g 7.47481e-19 $X=4.73 $Y=2.98
+ $X2=0 $Y2=0
cc_326 N_A_272_419#_c_289_n N_A_1028_23#_M1002_g 0.011568f $X=4.815 $Y=2.895
+ $X2=0 $Y2=0
cc_327 N_A_272_419#_c_289_n N_A_1028_23#_c_631_n 0.0214281f $X=4.815 $Y=2.895
+ $X2=0 $Y2=0
cc_328 N_A_272_419#_c_289_n N_A_1028_23#_c_646_n 0.0104011f $X=4.815 $Y=2.895
+ $X2=0 $Y2=0
cc_329 N_A_272_419#_M1007_g N_A_778_49#_c_804_n 0.00342901f $X=3.825 $Y=2.335
+ $X2=0 $Y2=0
cc_330 N_A_272_419#_c_302_n N_A_778_49#_c_804_n 0.0353442f $X=3.835 $Y=2.895
+ $X2=0 $Y2=0
cc_331 N_A_272_419#_c_303_n N_A_778_49#_c_804_n 0.0227215f $X=4.73 $Y=2.98 $X2=0
+ $Y2=0
cc_332 N_A_272_419#_c_289_n N_A_778_49#_c_804_n 0.0254791f $X=4.815 $Y=2.895
+ $X2=0 $Y2=0
cc_333 N_A_272_419#_M1019_g N_A_778_49#_c_794_n 0.0102393f $X=4.645 $Y=0.455
+ $X2=0 $Y2=0
cc_334 N_A_272_419#_c_292_n N_A_778_49#_c_794_n 0.0232055f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_335 N_A_272_419#_c_293_n N_A_778_49#_c_794_n 0.00124625f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_336 N_A_272_419#_M1019_g N_A_778_49#_c_795_n 0.00312316f $X=4.645 $Y=0.455
+ $X2=0 $Y2=0
cc_337 N_A_272_419#_c_292_n N_A_778_49#_c_797_n 0.0137327f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_338 N_A_272_419#_c_293_n N_A_778_49#_c_797_n 0.00111656f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_339 N_A_272_419#_M1007_g N_A_778_49#_c_798_n 4.90769e-19 $X=3.825 $Y=2.335
+ $X2=0 $Y2=0
cc_340 N_A_272_419#_M1019_g N_A_778_49#_c_798_n 0.00629113f $X=4.645 $Y=0.455
+ $X2=0 $Y2=0
cc_341 N_A_272_419#_c_288_n N_A_778_49#_c_798_n 0.0207504f $X=3.835 $Y=1.675
+ $X2=0 $Y2=0
cc_342 N_A_272_419#_c_302_n N_A_778_49#_c_798_n 0.00920001f $X=3.835 $Y=2.895
+ $X2=0 $Y2=0
cc_343 N_A_272_419#_c_289_n N_A_778_49#_c_798_n 0.0267693f $X=4.815 $Y=2.895
+ $X2=0 $Y2=0
cc_344 N_A_272_419#_c_291_n N_A_778_49#_c_798_n 6.4808e-19 $X=3.835 $Y=1.51
+ $X2=0 $Y2=0
cc_345 N_A_272_419#_c_292_n N_A_778_49#_c_798_n 0.0237562f $X=4.735 $Y=1.03
+ $X2=0 $Y2=0
cc_346 N_A_272_419#_c_299_n N_VPWR_M1011_d 0.0032149f $X=2.805 $Y=2.25 $X2=0
+ $Y2=0
cc_347 N_A_272_419#_c_322_p N_VPWR_M1011_d 0.0059706f $X=2.89 $Y=2.165 $X2=0
+ $Y2=0
cc_348 N_A_272_419#_M1011_g N_VPWR_c_1006_n 0.00465843f $X=2.725 $Y=2.175 $X2=0
+ $Y2=0
cc_349 N_A_272_419#_M1007_g N_VPWR_c_1006_n 4.06898e-19 $X=3.825 $Y=2.335 $X2=0
+ $Y2=0
cc_350 N_A_272_419#_c_299_n N_VPWR_c_1006_n 0.00587285f $X=2.805 $Y=2.25 $X2=0
+ $Y2=0
cc_351 N_A_272_419#_c_302_n N_VPWR_c_1006_n 0.007925f $X=3.835 $Y=2.895 $X2=0
+ $Y2=0
cc_352 N_A_272_419#_c_304_n N_VPWR_c_1006_n 0.00708746f $X=4 $Y=2.98 $X2=0 $Y2=0
cc_353 N_A_272_419#_c_303_n N_VPWR_c_1007_n 0.00718123f $X=4.73 $Y=2.98 $X2=0
+ $Y2=0
cc_354 N_A_272_419#_c_289_n N_VPWR_c_1007_n 0.0281395f $X=4.815 $Y=2.895 $X2=0
+ $Y2=0
cc_355 N_A_272_419#_M1007_g N_VPWR_c_1015_n 0.00121131f $X=3.825 $Y=2.335 $X2=0
+ $Y2=0
cc_356 N_A_272_419#_c_303_n N_VPWR_c_1015_n 0.0556369f $X=4.73 $Y=2.98 $X2=0
+ $Y2=0
cc_357 N_A_272_419#_c_304_n N_VPWR_c_1015_n 0.0222501f $X=4 $Y=2.98 $X2=0 $Y2=0
cc_358 N_A_272_419#_M1013_d N_VPWR_c_1004_n 0.00339068f $X=1.36 $Y=2.095 $X2=0
+ $Y2=0
cc_359 N_A_272_419#_M1011_g N_VPWR_c_1004_n 0.00152501f $X=2.725 $Y=2.175 $X2=0
+ $Y2=0
cc_360 N_A_272_419#_c_303_n N_VPWR_c_1004_n 0.0338465f $X=4.73 $Y=2.98 $X2=0
+ $Y2=0
cc_361 N_A_272_419#_c_304_n N_VPWR_c_1004_n 0.0127687f $X=4 $Y=2.98 $X2=0 $Y2=0
cc_362 N_A_272_419#_c_289_n A_955_367# 0.0127974f $X=4.815 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_363 N_A_272_419#_c_290_n N_VGND_c_1169_n 0.0153904f $X=1.86 $Y=0.77 $X2=0
+ $Y2=0
cc_364 N_A_272_419#_M1016_g N_VGND_c_1170_n 0.00539624f $X=2.635 $Y=0.455 $X2=0
+ $Y2=0
cc_365 N_A_272_419#_M1010_g N_VGND_c_1170_n 0.00477554f $X=2.995 $Y=0.455 $X2=0
+ $Y2=0
cc_366 N_A_272_419#_c_290_n N_VGND_c_1170_n 0.0080399f $X=1.86 $Y=0.77 $X2=0
+ $Y2=0
cc_367 N_A_272_419#_M1016_g N_VGND_c_1171_n 0.00212301f $X=2.635 $Y=0.455 $X2=0
+ $Y2=0
cc_368 N_A_272_419#_M1010_g N_VGND_c_1171_n 0.0108492f $X=2.995 $Y=0.455 $X2=0
+ $Y2=0
cc_369 N_A_272_419#_M1019_g N_VGND_c_1177_n 0.00398459f $X=4.645 $Y=0.455 $X2=0
+ $Y2=0
cc_370 N_A_272_419#_M1016_g N_VGND_c_1180_n 0.00721898f $X=2.635 $Y=0.455 $X2=0
+ $Y2=0
cc_371 N_A_272_419#_M1010_g N_VGND_c_1180_n 0.00425739f $X=2.995 $Y=0.455 $X2=0
+ $Y2=0
cc_372 N_A_272_419#_M1019_g N_VGND_c_1180_n 0.00667084f $X=4.645 $Y=0.455 $X2=0
+ $Y2=0
cc_373 N_A_272_419#_c_290_n N_VGND_c_1180_n 0.0105548f $X=1.86 $Y=0.77 $X2=0
+ $Y2=0
cc_374 N_A_27_112#_c_444_n N_A_455_49#_c_534_n 0.00101551f $X=3.405 $Y=1.105
+ $X2=0 $Y2=0
cc_375 N_A_27_112#_M1018_g N_A_455_49#_c_535_n 0.0206784f $X=3.425 $Y=0.455
+ $X2=0 $Y2=0
cc_376 N_A_27_112#_M1018_g N_A_455_49#_c_536_n 0.0119386f $X=3.425 $Y=0.455
+ $X2=0 $Y2=0
cc_377 N_A_27_112#_c_444_n N_A_455_49#_c_536_n 0.00142275f $X=3.405 $Y=1.105
+ $X2=0 $Y2=0
cc_378 N_A_27_112#_M1018_g N_A_455_49#_c_537_n 0.0368884f $X=3.425 $Y=0.455
+ $X2=0 $Y2=0
cc_379 N_A_27_112#_c_451_n N_VPWR_M1027_d 0.00807251f $X=1.825 $Y=2.6 $X2=-0.19
+ $Y2=-0.245
cc_380 N_A_27_112#_c_451_n N_VPWR_c_1005_n 0.0152435f $X=1.825 $Y=2.6 $X2=0
+ $Y2=0
cc_381 N_A_27_112#_c_453_n N_VPWR_c_1005_n 0.00152277f $X=1.99 $Y=2.9 $X2=0
+ $Y2=0
cc_382 N_A_27_112#_c_454_n N_VPWR_c_1005_n 0.0135888f $X=0.44 $Y=2.24 $X2=0
+ $Y2=0
cc_383 N_A_27_112#_c_447_n N_VPWR_c_1006_n 0.02365f $X=3.21 $Y=3.12 $X2=0 $Y2=0
cc_384 N_A_27_112#_M1025_g N_VPWR_c_1006_n 0.015064f $X=3.335 $Y=2.335 $X2=0
+ $Y2=0
cc_385 N_A_27_112#_c_451_n N_VPWR_c_1010_n 0.00318192f $X=1.825 $Y=2.6 $X2=0
+ $Y2=0
cc_386 N_A_27_112#_c_454_n N_VPWR_c_1010_n 0.0305459f $X=0.44 $Y=2.24 $X2=0
+ $Y2=0
cc_387 N_A_27_112#_c_451_n N_VPWR_c_1014_n 0.0112247f $X=1.825 $Y=2.6 $X2=0
+ $Y2=0
cc_388 N_A_27_112#_c_452_n N_VPWR_c_1014_n 0.0206619f $X=1.99 $Y=2.9 $X2=0 $Y2=0
cc_389 N_A_27_112#_c_453_n N_VPWR_c_1014_n 0.0325454f $X=1.99 $Y=2.9 $X2=0 $Y2=0
cc_390 N_A_27_112#_c_447_n N_VPWR_c_1015_n 0.00831182f $X=3.21 $Y=3.12 $X2=0
+ $Y2=0
cc_391 N_A_27_112#_M1027_s N_VPWR_c_1004_n 0.0023218f $X=0.295 $Y=2.095 $X2=0
+ $Y2=0
cc_392 N_A_27_112#_c_447_n N_VPWR_c_1004_n 0.0517126f $X=3.21 $Y=3.12 $X2=0
+ $Y2=0
cc_393 N_A_27_112#_c_451_n N_VPWR_c_1004_n 0.0246264f $X=1.825 $Y=2.6 $X2=0
+ $Y2=0
cc_394 N_A_27_112#_c_452_n N_VPWR_c_1004_n 0.0111091f $X=1.99 $Y=2.9 $X2=0 $Y2=0
cc_395 N_A_27_112#_c_453_n N_VPWR_c_1004_n 0.00890056f $X=1.99 $Y=2.9 $X2=0
+ $Y2=0
cc_396 N_A_27_112#_c_454_n N_VPWR_c_1004_n 0.0186989f $X=0.44 $Y=2.24 $X2=0
+ $Y2=0
cc_397 N_A_27_112#_c_445_n N_VGND_c_1169_n 0.0153904f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_398 N_A_27_112#_M1018_g N_VGND_c_1171_n 0.0114632f $X=3.425 $Y=0.455 $X2=0
+ $Y2=0
cc_399 N_A_27_112#_c_445_n N_VGND_c_1176_n 0.0080399f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_400 N_A_27_112#_M1018_g N_VGND_c_1177_n 0.00477554f $X=3.425 $Y=0.455 $X2=0
+ $Y2=0
cc_401 N_A_27_112#_M1018_g N_VGND_c_1180_n 0.00437771f $X=3.425 $Y=0.455 $X2=0
+ $Y2=0
cc_402 N_A_27_112#_c_445_n N_VGND_c_1180_n 0.0105548f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_403 N_A_455_49#_M1009_g N_A_1028_23#_M1002_g 0.0229405f $X=4.65 $Y=2.335
+ $X2=0 $Y2=0
cc_404 N_A_455_49#_c_529_n N_A_1028_23#_c_631_n 2.96074e-19 $X=4.525 $Y=1.51
+ $X2=0 $Y2=0
cc_405 N_A_455_49#_c_529_n N_A_1028_23#_c_632_n 0.0229405f $X=4.525 $Y=1.51
+ $X2=0 $Y2=0
cc_406 N_A_455_49#_c_529_n N_A_778_49#_c_804_n 0.00458624f $X=4.525 $Y=1.51
+ $X2=0 $Y2=0
cc_407 N_A_455_49#_c_530_n N_A_778_49#_c_804_n 4.46821e-19 $X=4.36 $Y=1.51 $X2=0
+ $Y2=0
cc_408 N_A_455_49#_M1009_g N_A_778_49#_c_804_n 0.00194315f $X=4.65 $Y=2.335
+ $X2=0 $Y2=0
cc_409 N_A_455_49#_c_527_n N_A_778_49#_c_798_n 0.00710526f $X=4.21 $Y=1.03 $X2=0
+ $Y2=0
cc_410 N_A_455_49#_c_528_n N_A_778_49#_c_798_n 0.0171883f $X=4.285 $Y=1.435
+ $X2=0 $Y2=0
cc_411 N_A_455_49#_c_529_n N_A_778_49#_c_798_n 0.00474087f $X=4.525 $Y=1.51
+ $X2=0 $Y2=0
cc_412 N_A_455_49#_c_530_n N_A_778_49#_c_798_n 0.00629218f $X=4.36 $Y=1.51 $X2=0
+ $Y2=0
cc_413 N_A_455_49#_M1009_g N_A_778_49#_c_798_n 0.00264528f $X=4.65 $Y=2.335
+ $X2=0 $Y2=0
cc_414 N_A_455_49#_c_534_n N_A_778_49#_c_798_n 0.0238727f $X=3.875 $Y=0.94 $X2=0
+ $Y2=0
cc_415 N_A_455_49#_c_535_n N_A_778_49#_c_798_n 6.88674e-19 $X=3.875 $Y=0.94
+ $X2=0 $Y2=0
cc_416 N_A_455_49#_c_537_n N_A_778_49#_c_798_n 0.00178552f $X=3.875 $Y=0.775
+ $X2=0 $Y2=0
cc_417 N_A_455_49#_c_527_n N_A_778_49#_c_799_n 5.00678e-19 $X=4.21 $Y=1.03 $X2=0
+ $Y2=0
cc_418 N_A_455_49#_c_537_n N_A_778_49#_c_799_n 0.00990824f $X=3.875 $Y=0.775
+ $X2=0 $Y2=0
cc_419 N_A_455_49#_M1009_g N_VPWR_c_1007_n 7.33128e-19 $X=4.65 $Y=2.335 $X2=0
+ $Y2=0
cc_420 N_A_455_49#_M1009_g N_VPWR_c_1015_n 0.00123074f $X=4.65 $Y=2.335 $X2=0
+ $Y2=0
cc_421 N_A_455_49#_c_531_n N_VGND_c_1170_n 0.0197956f $X=2.42 $Y=0.475 $X2=0
+ $Y2=0
cc_422 N_A_455_49#_c_531_n N_VGND_c_1171_n 0.0113755f $X=2.42 $Y=0.475 $X2=0
+ $Y2=0
cc_423 N_A_455_49#_c_536_n N_VGND_c_1171_n 0.0199112f $X=3.71 $Y=0.94 $X2=0
+ $Y2=0
cc_424 N_A_455_49#_c_537_n N_VGND_c_1171_n 0.00284061f $X=3.875 $Y=0.775 $X2=0
+ $Y2=0
cc_425 N_A_455_49#_c_535_n N_VGND_c_1177_n 0.00311545f $X=3.875 $Y=0.94 $X2=0
+ $Y2=0
cc_426 N_A_455_49#_c_537_n N_VGND_c_1177_n 0.00575161f $X=3.875 $Y=0.775 $X2=0
+ $Y2=0
cc_427 N_A_455_49#_M1016_s N_VGND_c_1180_n 0.00229455f $X=2.275 $Y=0.245 $X2=0
+ $Y2=0
cc_428 N_A_455_49#_c_531_n N_VGND_c_1180_n 0.0125833f $X=2.42 $Y=0.475 $X2=0
+ $Y2=0
cc_429 N_A_455_49#_c_534_n N_VGND_c_1180_n 0.0110376f $X=3.875 $Y=0.94 $X2=0
+ $Y2=0
cc_430 N_A_455_49#_c_535_n N_VGND_c_1180_n 0.00423998f $X=3.875 $Y=0.94 $X2=0
+ $Y2=0
cc_431 N_A_455_49#_c_536_n N_VGND_c_1180_n 0.0272995f $X=3.71 $Y=0.94 $X2=0
+ $Y2=0
cc_432 N_A_455_49#_c_537_n N_VGND_c_1180_n 0.00690128f $X=3.875 $Y=0.775 $X2=0
+ $Y2=0
cc_433 N_A_1028_23#_M1002_g N_A_778_49#_M1021_g 0.0214851f $X=5.265 $Y=2.335
+ $X2=0 $Y2=0
cc_434 N_A_1028_23#_c_631_n N_A_778_49#_M1021_g 8.78527e-19 $X=5.305 $Y=1.51
+ $X2=0 $Y2=0
cc_435 N_A_1028_23#_c_645_n N_A_778_49#_M1021_g 0.0232926f $X=6.015 $Y=1.8 $X2=0
+ $Y2=0
cc_436 N_A_1028_23#_c_647_n N_A_778_49#_M1021_g 0.00685128f $X=6.18 $Y=2.69
+ $X2=0 $Y2=0
cc_437 N_A_1028_23#_c_648_n N_A_778_49#_M1021_g 0.00364325f $X=6.305 $Y=1.715
+ $X2=0 $Y2=0
cc_438 N_A_1028_23#_c_633_n N_A_778_49#_c_790_n 0.0080528f $X=6.305 $Y=1.365
+ $X2=0 $Y2=0
cc_439 N_A_1028_23#_c_637_n N_A_778_49#_c_790_n 0.00650364f $X=6.305 $Y=0.495
+ $X2=0 $Y2=0
cc_440 N_A_1028_23#_c_650_n N_A_778_49#_c_790_n 0.00429414f $X=6.18 $Y=1.88
+ $X2=0 $Y2=0
cc_441 N_A_1028_23#_M1028_g N_A_778_49#_c_791_n 0.0141198f $X=5.215 $Y=0.455
+ $X2=0 $Y2=0
cc_442 N_A_1028_23#_c_637_n N_A_778_49#_c_791_n 9.53509e-19 $X=6.305 $Y=0.495
+ $X2=0 $Y2=0
cc_443 N_A_1028_23#_c_633_n N_A_778_49#_M1020_g 0.0101949f $X=6.305 $Y=1.365
+ $X2=0 $Y2=0
cc_444 N_A_1028_23#_c_637_n N_A_778_49#_M1020_g 0.0090435f $X=6.305 $Y=0.495
+ $X2=0 $Y2=0
cc_445 N_A_1028_23#_c_645_n N_A_778_49#_c_793_n 3.7612e-19 $X=6.015 $Y=1.8 $X2=0
+ $Y2=0
cc_446 N_A_1028_23#_M1028_g N_A_778_49#_c_794_n 0.00758478f $X=5.215 $Y=0.455
+ $X2=0 $Y2=0
cc_447 N_A_1028_23#_M1028_g N_A_778_49#_c_795_n 0.00978509f $X=5.215 $Y=0.455
+ $X2=0 $Y2=0
cc_448 N_A_1028_23#_M1028_g N_A_778_49#_c_796_n 0.00573508f $X=5.215 $Y=0.455
+ $X2=0 $Y2=0
cc_449 N_A_1028_23#_c_631_n N_A_778_49#_c_796_n 0.0107668f $X=5.305 $Y=1.51
+ $X2=0 $Y2=0
cc_450 N_A_1028_23#_c_632_n N_A_778_49#_c_796_n 0.00110453f $X=5.305 $Y=1.51
+ $X2=0 $Y2=0
cc_451 N_A_1028_23#_M1028_g N_A_778_49#_c_797_n 0.004593f $X=5.215 $Y=0.455
+ $X2=0 $Y2=0
cc_452 N_A_1028_23#_c_631_n N_A_778_49#_c_797_n 0.00546986f $X=5.305 $Y=1.51
+ $X2=0 $Y2=0
cc_453 N_A_1028_23#_M1028_g N_A_778_49#_c_800_n 0.00174987f $X=5.215 $Y=0.455
+ $X2=0 $Y2=0
cc_454 N_A_1028_23#_c_631_n N_A_778_49#_c_800_n 0.0107959f $X=5.305 $Y=1.51
+ $X2=0 $Y2=0
cc_455 N_A_1028_23#_c_632_n N_A_778_49#_c_800_n 6.98837e-19 $X=5.305 $Y=1.51
+ $X2=0 $Y2=0
cc_456 N_A_1028_23#_c_645_n N_A_778_49#_c_800_n 0.0222574f $X=6.015 $Y=1.8 $X2=0
+ $Y2=0
cc_457 N_A_1028_23#_c_633_n N_A_778_49#_c_800_n 0.0360857f $X=6.305 $Y=1.365
+ $X2=0 $Y2=0
cc_458 N_A_1028_23#_c_637_n N_A_778_49#_c_800_n 0.0102709f $X=6.305 $Y=0.495
+ $X2=0 $Y2=0
cc_459 N_A_1028_23#_c_650_n N_A_778_49#_c_800_n 0.00204652f $X=6.18 $Y=1.88
+ $X2=0 $Y2=0
cc_460 N_A_1028_23#_c_638_n N_A_778_49#_c_800_n 0.0136967f $X=6.305 $Y=1.45
+ $X2=0 $Y2=0
cc_461 N_A_1028_23#_c_631_n N_A_778_49#_c_801_n 0.00164466f $X=5.305 $Y=1.51
+ $X2=0 $Y2=0
cc_462 N_A_1028_23#_c_632_n N_A_778_49#_c_801_n 0.0178661f $X=5.305 $Y=1.51
+ $X2=0 $Y2=0
cc_463 N_A_1028_23#_c_633_n N_A_778_49#_c_801_n 0.00307165f $X=6.305 $Y=1.365
+ $X2=0 $Y2=0
cc_464 N_A_1028_23#_c_638_n N_A_778_49#_c_801_n 0.00138125f $X=6.305 $Y=1.45
+ $X2=0 $Y2=0
cc_465 N_A_1028_23#_c_629_n N_RESET_B_M1015_g 0.0159863f $X=7.1 $Y=1.535 $X2=0
+ $Y2=0
cc_466 N_A_1028_23#_c_647_n N_RESET_B_M1015_g 0.00796692f $X=6.18 $Y=2.69 $X2=0
+ $Y2=0
cc_467 N_A_1028_23#_c_648_n N_RESET_B_M1015_g 0.00504707f $X=6.305 $Y=1.715
+ $X2=0 $Y2=0
cc_468 N_A_1028_23#_c_634_n N_RESET_B_M1015_g 0.0106959f $X=6.935 $Y=1.45 $X2=0
+ $Y2=0
cc_469 N_A_1028_23#_c_650_n N_RESET_B_M1015_g 0.00140473f $X=6.18 $Y=1.88 $X2=0
+ $Y2=0
cc_470 N_A_1028_23#_M1005_g N_RESET_B_M1023_g 0.016618f $X=7.08 $Y=0.455 $X2=0
+ $Y2=0
cc_471 N_A_1028_23#_c_625_n N_RESET_B_M1023_g 0.0207394f $X=7.515 $Y=0.94 $X2=0
+ $Y2=0
cc_472 N_A_1028_23#_c_633_n N_RESET_B_M1023_g 0.00881247f $X=6.305 $Y=1.365
+ $X2=0 $Y2=0
cc_473 N_A_1028_23#_c_634_n N_RESET_B_M1023_g 0.00694572f $X=6.935 $Y=1.45 $X2=0
+ $Y2=0
cc_474 N_A_1028_23#_c_635_n N_RESET_B_M1023_g 0.00191323f $X=7.1 $Y=1.03 $X2=0
+ $Y2=0
cc_475 N_A_1028_23#_c_637_n N_RESET_B_M1023_g 0.00102965f $X=6.305 $Y=0.495
+ $X2=0 $Y2=0
cc_476 N_A_1028_23#_M1003_g N_RESET_B_c_893_n 0.0170394f $X=7.06 $Y=2.235 $X2=0
+ $Y2=0
cc_477 N_A_1028_23#_M1004_g N_RESET_B_c_895_n 0.00258039f $X=8.74 $Y=2.37 $X2=0
+ $Y2=0
cc_478 N_A_1028_23#_c_634_n N_RESET_B_c_891_n 0.0109187f $X=6.935 $Y=1.45 $X2=0
+ $Y2=0
cc_479 N_A_1028_23#_c_636_n N_RESET_B_c_891_n 0.0207394f $X=7.1 $Y=1.03 $X2=0
+ $Y2=0
cc_480 N_A_1028_23#_M1003_g N_RESET_B_c_899_n 0.0047934f $X=7.06 $Y=2.235 $X2=0
+ $Y2=0
cc_481 N_A_1028_23#_M1004_g N_RESET_B_c_899_n 0.00609841f $X=8.74 $Y=2.37 $X2=0
+ $Y2=0
cc_482 N_A_1028_23#_c_628_n N_A_1614_74#_M1017_g 0.0214027f $X=8.79 $Y=0.865
+ $X2=0 $Y2=0
cc_483 N_A_1028_23#_c_630_n N_A_1614_74#_c_943_n 0.0214027f $X=8.79 $Y=0.94
+ $X2=0 $Y2=0
cc_484 N_A_1028_23#_M1004_g N_A_1614_74#_c_944_n 0.0214027f $X=8.74 $Y=2.37
+ $X2=0 $Y2=0
cc_485 N_A_1028_23#_M1024_g N_A_1614_74#_c_945_n 0.001582f $X=7.44 $Y=0.455
+ $X2=0 $Y2=0
cc_486 N_A_1028_23#_c_624_n N_A_1614_74#_c_945_n 0.0123233f $X=8.355 $Y=0.94
+ $X2=0 $Y2=0
cc_487 N_A_1028_23#_c_626_n N_A_1614_74#_c_945_n 0.011008f $X=8.43 $Y=0.865
+ $X2=0 $Y2=0
cc_488 N_A_1028_23#_c_628_n N_A_1614_74#_c_945_n 0.00152289f $X=8.79 $Y=0.865
+ $X2=0 $Y2=0
cc_489 N_A_1028_23#_c_630_n N_A_1614_74#_c_945_n 0.00596677f $X=8.79 $Y=0.94
+ $X2=0 $Y2=0
cc_490 N_A_1028_23#_c_624_n N_A_1614_74#_c_946_n 0.00112211f $X=8.355 $Y=0.94
+ $X2=0 $Y2=0
cc_491 N_A_1028_23#_M1004_g N_A_1614_74#_c_946_n 0.0460456f $X=8.74 $Y=2.37
+ $X2=0 $Y2=0
cc_492 N_A_1028_23#_M1004_g N_A_1614_74#_c_947_n 0.0146055f $X=8.74 $Y=2.37
+ $X2=0 $Y2=0
cc_493 N_A_1028_23#_c_630_n N_A_1614_74#_c_947_n 0.00997648f $X=8.79 $Y=0.94
+ $X2=0 $Y2=0
cc_494 N_A_1028_23#_c_624_n N_A_1614_74#_c_948_n 0.00746669f $X=8.355 $Y=0.94
+ $X2=0 $Y2=0
cc_495 N_A_1028_23#_M1004_g N_A_1614_74#_c_948_n 0.00370646f $X=8.74 $Y=2.37
+ $X2=0 $Y2=0
cc_496 N_A_1028_23#_c_630_n N_A_1614_74#_c_948_n 0.0150096f $X=8.79 $Y=0.94
+ $X2=0 $Y2=0
cc_497 N_A_1028_23#_M1004_g N_A_1614_74#_c_949_n 0.00205744f $X=8.74 $Y=2.37
+ $X2=0 $Y2=0
cc_498 N_A_1028_23#_c_645_n N_VPWR_M1002_d 0.00198167f $X=6.015 $Y=1.8 $X2=0
+ $Y2=0
cc_499 N_A_1028_23#_c_646_n N_VPWR_M1002_d 2.47671e-19 $X=5.47 $Y=1.8 $X2=0
+ $Y2=0
cc_500 N_A_1028_23#_M1002_g N_VPWR_c_1007_n 0.0203193f $X=5.265 $Y=2.335 $X2=0
+ $Y2=0
cc_501 N_A_1028_23#_c_632_n N_VPWR_c_1007_n 2.67792e-19 $X=5.305 $Y=1.51 $X2=0
+ $Y2=0
cc_502 N_A_1028_23#_c_645_n N_VPWR_c_1007_n 0.0142305f $X=6.015 $Y=1.8 $X2=0
+ $Y2=0
cc_503 N_A_1028_23#_c_646_n N_VPWR_c_1007_n 0.00382016f $X=5.47 $Y=1.8 $X2=0
+ $Y2=0
cc_504 N_A_1028_23#_c_647_n N_VPWR_c_1007_n 0.00102756f $X=6.18 $Y=2.69 $X2=0
+ $Y2=0
cc_505 N_A_1028_23#_M1003_g N_VPWR_c_1008_n 0.0220602f $X=7.06 $Y=2.235 $X2=0
+ $Y2=0
cc_506 N_A_1028_23#_c_647_n N_VPWR_c_1008_n 0.0321224f $X=6.18 $Y=2.69 $X2=0
+ $Y2=0
cc_507 N_A_1028_23#_c_634_n N_VPWR_c_1008_n 0.0263569f $X=6.935 $Y=1.45 $X2=0
+ $Y2=0
cc_508 N_A_1028_23#_c_650_n N_VPWR_c_1008_n 0.00564652f $X=6.18 $Y=1.88 $X2=0
+ $Y2=0
cc_509 N_A_1028_23#_M1004_g N_VPWR_c_1009_n 0.0266261f $X=8.74 $Y=2.37 $X2=0
+ $Y2=0
cc_510 N_A_1028_23#_c_647_n N_VPWR_c_1012_n 0.0110296f $X=6.18 $Y=2.69 $X2=0
+ $Y2=0
cc_511 N_A_1028_23#_M1002_g N_VPWR_c_1015_n 0.00735144f $X=5.265 $Y=2.335 $X2=0
+ $Y2=0
cc_512 N_A_1028_23#_M1004_g N_VPWR_c_1016_n 0.00747382f $X=8.74 $Y=2.37 $X2=0
+ $Y2=0
cc_513 N_A_1028_23#_M1002_g N_VPWR_c_1004_n 0.00763694f $X=5.265 $Y=2.335 $X2=0
+ $Y2=0
cc_514 N_A_1028_23#_M1003_g N_VPWR_c_1004_n 0.00129615f $X=7.06 $Y=2.235 $X2=0
+ $Y2=0
cc_515 N_A_1028_23#_M1004_g N_VPWR_c_1004_n 0.00779694f $X=8.74 $Y=2.37 $X2=0
+ $Y2=0
cc_516 N_A_1028_23#_c_647_n N_VPWR_c_1004_n 0.0126983f $X=6.18 $Y=2.69 $X2=0
+ $Y2=0
cc_517 N_A_1028_23#_M1003_g N_Q_c_1114_n 0.00466735f $X=7.06 $Y=2.235 $X2=0
+ $Y2=0
cc_518 N_A_1028_23#_c_625_n N_Q_c_1114_n 0.00252629f $X=7.515 $Y=0.94 $X2=0
+ $Y2=0
cc_519 N_A_1028_23#_c_629_n N_Q_c_1114_n 6.21329e-19 $X=7.1 $Y=1.535 $X2=0 $Y2=0
cc_520 N_A_1028_23#_c_634_n N_Q_c_1114_n 0.00875918f $X=6.935 $Y=1.45 $X2=0
+ $Y2=0
cc_521 N_A_1028_23#_M1003_g N_Q_c_1112_n 0.00590404f $X=7.06 $Y=2.235 $X2=0
+ $Y2=0
cc_522 N_A_1028_23#_M1024_g N_Q_c_1112_n 0.00640238f $X=7.44 $Y=0.455 $X2=0
+ $Y2=0
cc_523 N_A_1028_23#_c_624_n N_Q_c_1112_n 0.00746452f $X=8.355 $Y=0.94 $X2=0
+ $Y2=0
cc_524 N_A_1028_23#_c_625_n N_Q_c_1112_n 0.00482365f $X=7.515 $Y=0.94 $X2=0
+ $Y2=0
cc_525 N_A_1028_23#_c_634_n N_Q_c_1112_n 0.0129674f $X=6.935 $Y=1.45 $X2=0 $Y2=0
cc_526 N_A_1028_23#_c_635_n N_Q_c_1112_n 0.0353562f $X=7.1 $Y=1.03 $X2=0 $Y2=0
cc_527 N_A_1028_23#_c_636_n N_Q_c_1112_n 0.00895567f $X=7.1 $Y=1.03 $X2=0 $Y2=0
cc_528 N_A_1028_23#_M1005_g N_Q_c_1113_n 0.0022222f $X=7.08 $Y=0.455 $X2=0 $Y2=0
cc_529 N_A_1028_23#_M1024_g N_Q_c_1113_n 0.00891319f $X=7.44 $Y=0.455 $X2=0
+ $Y2=0
cc_530 N_A_1028_23#_c_624_n N_Q_c_1113_n 0.00773111f $X=8.355 $Y=0.94 $X2=0
+ $Y2=0
cc_531 N_A_1028_23#_c_626_n N_Q_c_1113_n 0.00286361f $X=8.43 $Y=0.865 $X2=0
+ $Y2=0
cc_532 N_A_1028_23#_M1003_g Q 0.0181517f $X=7.06 $Y=2.235 $X2=0 $Y2=0
cc_533 N_A_1028_23#_M1004_g N_Q_N_c_1151_n 2.74877e-19 $X=8.74 $Y=2.37 $X2=0
+ $Y2=0
cc_534 N_A_1028_23#_M1028_g N_VGND_c_1172_n 0.0172259f $X=5.215 $Y=0.455 $X2=0
+ $Y2=0
cc_535 N_A_1028_23#_c_637_n N_VGND_c_1172_n 0.0257883f $X=6.305 $Y=0.495 $X2=0
+ $Y2=0
cc_536 N_A_1028_23#_M1005_g N_VGND_c_1173_n 0.0123852f $X=7.08 $Y=0.455 $X2=0
+ $Y2=0
cc_537 N_A_1028_23#_M1024_g N_VGND_c_1173_n 0.00231094f $X=7.44 $Y=0.455 $X2=0
+ $Y2=0
cc_538 N_A_1028_23#_c_625_n N_VGND_c_1173_n 5.35752e-19 $X=7.515 $Y=0.94 $X2=0
+ $Y2=0
cc_539 N_A_1028_23#_c_635_n N_VGND_c_1173_n 0.00762588f $X=7.1 $Y=1.03 $X2=0
+ $Y2=0
cc_540 N_A_1028_23#_c_637_n N_VGND_c_1173_n 0.00931701f $X=6.305 $Y=0.495 $X2=0
+ $Y2=0
cc_541 N_A_1028_23#_M1005_g N_VGND_c_1174_n 0.00477554f $X=7.08 $Y=0.455 $X2=0
+ $Y2=0
cc_542 N_A_1028_23#_M1024_g N_VGND_c_1174_n 0.00472992f $X=7.44 $Y=0.455 $X2=0
+ $Y2=0
cc_543 N_A_1028_23#_c_626_n N_VGND_c_1174_n 0.00434272f $X=8.43 $Y=0.865 $X2=0
+ $Y2=0
cc_544 N_A_1028_23#_c_628_n N_VGND_c_1174_n 0.00383152f $X=8.79 $Y=0.865 $X2=0
+ $Y2=0
cc_545 N_A_1028_23#_c_626_n N_VGND_c_1175_n 0.00182089f $X=8.43 $Y=0.865 $X2=0
+ $Y2=0
cc_546 N_A_1028_23#_c_628_n N_VGND_c_1175_n 0.0122129f $X=8.79 $Y=0.865 $X2=0
+ $Y2=0
cc_547 N_A_1028_23#_M1028_g N_VGND_c_1177_n 0.00445461f $X=5.215 $Y=0.455 $X2=0
+ $Y2=0
cc_548 N_A_1028_23#_c_637_n N_VGND_c_1178_n 0.0221634f $X=6.305 $Y=0.495 $X2=0
+ $Y2=0
cc_549 N_A_1028_23#_M1020_s N_VGND_c_1180_n 0.00232384f $X=5.93 $Y=0.245 $X2=0
+ $Y2=0
cc_550 N_A_1028_23#_M1028_g N_VGND_c_1180_n 0.00865943f $X=5.215 $Y=0.455 $X2=0
+ $Y2=0
cc_551 N_A_1028_23#_M1005_g N_VGND_c_1180_n 0.00442294f $X=7.08 $Y=0.455 $X2=0
+ $Y2=0
cc_552 N_A_1028_23#_M1024_g N_VGND_c_1180_n 0.00941849f $X=7.44 $Y=0.455 $X2=0
+ $Y2=0
cc_553 N_A_1028_23#_c_624_n N_VGND_c_1180_n 0.00466911f $X=8.355 $Y=0.94 $X2=0
+ $Y2=0
cc_554 N_A_1028_23#_c_625_n N_VGND_c_1180_n 2.77112e-19 $X=7.515 $Y=0.94 $X2=0
+ $Y2=0
cc_555 N_A_1028_23#_c_626_n N_VGND_c_1180_n 0.00825516f $X=8.43 $Y=0.865 $X2=0
+ $Y2=0
cc_556 N_A_1028_23#_c_628_n N_VGND_c_1180_n 0.00756787f $X=8.79 $Y=0.865 $X2=0
+ $Y2=0
cc_557 N_A_1028_23#_c_630_n N_VGND_c_1180_n 7.5656e-19 $X=8.79 $Y=0.94 $X2=0
+ $Y2=0
cc_558 N_A_1028_23#_c_635_n N_VGND_c_1180_n 0.00796506f $X=7.1 $Y=1.03 $X2=0
+ $Y2=0
cc_559 N_A_1028_23#_c_637_n N_VGND_c_1180_n 0.0171542f $X=6.305 $Y=0.495 $X2=0
+ $Y2=0
cc_560 N_A_778_49#_M1021_g N_RESET_B_M1015_g 0.029173f $X=5.835 $Y=2.335 $X2=0
+ $Y2=0
cc_561 N_A_778_49#_M1020_g N_RESET_B_M1023_g 0.0546129f $X=6.29 $Y=0.455 $X2=0
+ $Y2=0
cc_562 N_A_778_49#_c_801_n N_RESET_B_M1023_g 0.00519515f $X=5.875 $Y=1.03 $X2=0
+ $Y2=0
cc_563 N_A_778_49#_c_793_n N_RESET_B_c_891_n 0.00485955f $X=5.875 $Y=1.535 $X2=0
+ $Y2=0
cc_564 N_A_778_49#_M1021_g N_VPWR_c_1007_n 0.00390445f $X=5.835 $Y=2.335 $X2=0
+ $Y2=0
cc_565 N_A_778_49#_M1021_g N_VPWR_c_1008_n 7.49999e-19 $X=5.835 $Y=2.335 $X2=0
+ $Y2=0
cc_566 N_A_778_49#_M1021_g N_VPWR_c_1012_n 0.00818076f $X=5.835 $Y=2.335 $X2=0
+ $Y2=0
cc_567 N_A_778_49#_M1021_g N_VPWR_c_1004_n 0.00844794f $X=5.835 $Y=2.335 $X2=0
+ $Y2=0
cc_568 N_A_778_49#_M1020_g N_VGND_c_1172_n 0.00354768f $X=6.29 $Y=0.455 $X2=0
+ $Y2=0
cc_569 N_A_778_49#_c_794_n N_VGND_c_1172_n 0.0131617f $X=5.08 $Y=0.6 $X2=0 $Y2=0
cc_570 N_A_778_49#_c_796_n N_VGND_c_1172_n 0.0201141f $X=5.71 $Y=0.95 $X2=0
+ $Y2=0
cc_571 N_A_778_49#_M1020_g N_VGND_c_1173_n 0.0017887f $X=6.29 $Y=0.455 $X2=0
+ $Y2=0
cc_572 N_A_778_49#_c_794_n N_VGND_c_1177_n 0.0148453f $X=5.08 $Y=0.6 $X2=0 $Y2=0
cc_573 N_A_778_49#_c_799_n N_VGND_c_1177_n 0.0198132f $X=4.55 $Y=0.475 $X2=0
+ $Y2=0
cc_574 N_A_778_49#_M1020_g N_VGND_c_1178_n 0.00361198f $X=6.29 $Y=0.455 $X2=0
+ $Y2=0
cc_575 N_A_778_49#_M1026_d N_VGND_c_1180_n 0.0126135f $X=3.89 $Y=0.245 $X2=0
+ $Y2=0
cc_576 N_A_778_49#_M1020_g N_VGND_c_1180_n 0.0064746f $X=6.29 $Y=0.455 $X2=0
+ $Y2=0
cc_577 N_A_778_49#_c_794_n N_VGND_c_1180_n 0.0208527f $X=5.08 $Y=0.6 $X2=0 $Y2=0
cc_578 N_A_778_49#_c_799_n N_VGND_c_1180_n 0.0125997f $X=4.55 $Y=0.475 $X2=0
+ $Y2=0
cc_579 N_A_778_49#_c_800_n N_VGND_c_1180_n 0.00712208f $X=5.875 $Y=1.03 $X2=0
+ $Y2=0
cc_580 N_A_778_49#_c_794_n A_944_49# 0.00499687f $X=5.08 $Y=0.6 $X2=-0.19
+ $Y2=-0.245
cc_581 RESET_B N_A_1614_74#_c_946_n 0.0732652f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_582 N_RESET_B_c_899_n N_A_1614_74#_c_946_n 0.00600415f $X=7.96 $Y=2.385 $X2=0
+ $Y2=0
cc_583 N_RESET_B_M1015_g N_VPWR_c_1008_n 0.029939f $X=6.525 $Y=2.235 $X2=0 $Y2=0
cc_584 N_RESET_B_c_893_n N_VPWR_c_1008_n 0.0184879f $X=7.795 $Y=3.15 $X2=0 $Y2=0
cc_585 N_RESET_B_c_894_n N_VPWR_c_1008_n 0.0041055f $X=6.65 $Y=3.15 $X2=0 $Y2=0
cc_586 N_RESET_B_c_891_n N_VPWR_c_1008_n 5.6787e-19 $X=6.562 $Y=1.525 $X2=0
+ $Y2=0
cc_587 N_RESET_B_c_894_n N_VPWR_c_1012_n 0.008763f $X=6.65 $Y=3.15 $X2=0 $Y2=0
cc_588 N_RESET_B_c_893_n N_VPWR_c_1016_n 0.0280947f $X=7.795 $Y=3.15 $X2=0 $Y2=0
cc_589 N_RESET_B_c_897_n N_VPWR_c_1016_n 9.00552e-19 $X=7.96 $Y=2.89 $X2=0 $Y2=0
cc_590 RESET_B N_VPWR_c_1016_n 0.00985655f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_591 N_RESET_B_c_893_n N_VPWR_c_1004_n 0.0341933f $X=7.795 $Y=3.15 $X2=0 $Y2=0
cc_592 N_RESET_B_c_894_n N_VPWR_c_1004_n 0.0160133f $X=6.65 $Y=3.15 $X2=0 $Y2=0
cc_593 RESET_B N_VPWR_c_1004_n 0.010519f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_594 N_RESET_B_M1015_g N_Q_c_1114_n 3.46043e-19 $X=6.525 $Y=2.235 $X2=0 $Y2=0
cc_595 RESET_B N_Q_c_1114_n 0.076641f $X=7.835 $Y=1.95 $X2=0 $Y2=0
cc_596 N_RESET_B_c_893_n Q 0.00980269f $X=7.795 $Y=3.15 $X2=0 $Y2=0
cc_597 N_RESET_B_c_899_n Q 0.00727818f $X=7.96 $Y=2.385 $X2=0 $Y2=0
cc_598 N_RESET_B_M1023_g N_VGND_c_1173_n 0.0125728f $X=6.65 $Y=0.455 $X2=0 $Y2=0
cc_599 N_RESET_B_M1023_g N_VGND_c_1178_n 0.00477554f $X=6.65 $Y=0.455 $X2=0
+ $Y2=0
cc_600 N_RESET_B_M1023_g N_VGND_c_1180_n 0.00814835f $X=6.65 $Y=0.455 $X2=0
+ $Y2=0
cc_601 N_A_1614_74#_M1022_g N_VPWR_c_1009_n 0.0257325f $X=9.27 $Y=2.37 $X2=0
+ $Y2=0
cc_602 N_A_1614_74#_c_946_n N_VPWR_c_1009_n 0.0685263f $X=8.475 $Y=2.015 $X2=0
+ $Y2=0
cc_603 N_A_1614_74#_c_949_n N_VPWR_c_1009_n 0.00177713f $X=9.31 $Y=1.155 $X2=0
+ $Y2=0
cc_604 N_A_1614_74#_c_946_n N_VPWR_c_1016_n 0.0106618f $X=8.475 $Y=2.015 $X2=0
+ $Y2=0
cc_605 N_A_1614_74#_M1022_g N_VPWR_c_1017_n 0.00747382f $X=9.27 $Y=2.37 $X2=0
+ $Y2=0
cc_606 N_A_1614_74#_M1022_g N_VPWR_c_1004_n 0.00779694f $X=9.27 $Y=2.37 $X2=0
+ $Y2=0
cc_607 N_A_1614_74#_c_946_n N_VPWR_c_1004_n 0.0114128f $X=8.475 $Y=2.015 $X2=0
+ $Y2=0
cc_608 N_A_1614_74#_c_945_n N_Q_c_1112_n 0.0116112f $X=8.215 $Y=0.58 $X2=0 $Y2=0
cc_609 N_A_1614_74#_c_948_n N_Q_c_1112_n 0.00719162f $X=8.64 $Y=1.075 $X2=0
+ $Y2=0
cc_610 N_A_1614_74#_c_945_n N_Q_c_1113_n 0.0228056f $X=8.215 $Y=0.58 $X2=0 $Y2=0
cc_611 N_A_1614_74#_M1017_g Q_N 0.00125204f $X=9.22 $Y=0.58 $X2=0 $Y2=0
cc_612 N_A_1614_74#_M1012_g Q_N 0.0100639f $X=9.58 $Y=0.58 $X2=0 $Y2=0
cc_613 N_A_1614_74#_M1022_g Q_N 0.00600337f $X=9.27 $Y=2.37 $X2=0 $Y2=0
cc_614 N_A_1614_74#_M1012_g Q_N 0.0114523f $X=9.58 $Y=0.58 $X2=0 $Y2=0
cc_615 N_A_1614_74#_c_949_n Q_N 0.039205f $X=9.31 $Y=1.155 $X2=0 $Y2=0
cc_616 N_A_1614_74#_c_950_n Q_N 0.0108326f $X=9.31 $Y=1.155 $X2=0 $Y2=0
cc_617 N_A_1614_74#_M1022_g Q_N 0.0134647f $X=9.27 $Y=2.37 $X2=0 $Y2=0
cc_618 N_A_1614_74#_M1022_g N_Q_N_c_1151_n 0.00585731f $X=9.27 $Y=2.37 $X2=0
+ $Y2=0
cc_619 N_A_1614_74#_c_944_n N_Q_N_c_1151_n 6.09582e-19 $X=9.31 $Y=1.66 $X2=0
+ $Y2=0
cc_620 N_A_1614_74#_c_949_n N_Q_N_c_1151_n 0.00832065f $X=9.31 $Y=1.155 $X2=0
+ $Y2=0
cc_621 N_A_1614_74#_c_945_n N_VGND_c_1174_n 0.0144999f $X=8.215 $Y=0.58 $X2=0
+ $Y2=0
cc_622 N_A_1614_74#_M1017_g N_VGND_c_1175_n 0.0122119f $X=9.22 $Y=0.58 $X2=0
+ $Y2=0
cc_623 N_A_1614_74#_M1012_g N_VGND_c_1175_n 0.00182089f $X=9.58 $Y=0.58 $X2=0
+ $Y2=0
cc_624 N_A_1614_74#_c_945_n N_VGND_c_1175_n 0.0153904f $X=8.215 $Y=0.58 $X2=0
+ $Y2=0
cc_625 N_A_1614_74#_c_947_n N_VGND_c_1175_n 0.024419f $X=9.145 $Y=1.075 $X2=0
+ $Y2=0
cc_626 N_A_1614_74#_c_949_n N_VGND_c_1175_n 0.00193744f $X=9.31 $Y=1.155 $X2=0
+ $Y2=0
cc_627 N_A_1614_74#_M1017_g N_VGND_c_1179_n 0.00383152f $X=9.22 $Y=0.58 $X2=0
+ $Y2=0
cc_628 N_A_1614_74#_M1012_g N_VGND_c_1179_n 0.00434272f $X=9.58 $Y=0.58 $X2=0
+ $Y2=0
cc_629 N_A_1614_74#_M1017_g N_VGND_c_1180_n 0.00756787f $X=9.22 $Y=0.58 $X2=0
+ $Y2=0
cc_630 N_A_1614_74#_M1012_g N_VGND_c_1180_n 0.00824192f $X=9.58 $Y=0.58 $X2=0
+ $Y2=0
cc_631 N_A_1614_74#_c_945_n N_VGND_c_1180_n 0.0119734f $X=8.215 $Y=0.58 $X2=0
+ $Y2=0
cc_632 N_VPWR_c_1008_n N_Q_c_1114_n 0.0780031f $X=6.79 $Y=1.88 $X2=0 $Y2=0
cc_633 N_VPWR_c_1016_n Q 0.0147934f $X=8.84 $Y=3.33 $X2=0 $Y2=0
cc_634 N_VPWR_c_1004_n Q 0.0139796f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_635 N_VPWR_c_1017_n Q_N 0.0191637f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_636 N_VPWR_c_1004_n Q_N 0.0204781f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_637 N_VPWR_c_1009_n N_Q_N_c_1151_n 0.071673f $X=9.005 $Y=2.015 $X2=0 $Y2=0
cc_638 N_Q_c_1113_n N_VGND_c_1173_n 0.0154867f $X=7.655 $Y=0.475 $X2=0 $Y2=0
cc_639 N_Q_c_1113_n N_VGND_c_1174_n 0.0222062f $X=7.655 $Y=0.475 $X2=0 $Y2=0
cc_640 N_Q_M1024_d N_VGND_c_1180_n 0.00229455f $X=7.515 $Y=0.245 $X2=0 $Y2=0
cc_641 N_Q_c_1113_n N_VGND_c_1180_n 0.0140153f $X=7.655 $Y=0.475 $X2=0 $Y2=0
cc_642 Q_N N_VGND_c_1175_n 0.0153904f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_643 Q_N N_VGND_c_1179_n 0.0144513f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_644 Q_N N_VGND_c_1180_n 0.0119539f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_645 N_VGND_c_1180_n A_542_49# 0.00290859f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_646 N_VGND_c_1180_n A_700_49# 0.00331961f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_647 N_VGND_c_1180_n A_944_49# 0.00418818f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_648 N_VGND_c_1180_n A_1273_49# 0.00811909f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_649 N_VGND_c_1180_n A_1431_49# 0.00571915f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
