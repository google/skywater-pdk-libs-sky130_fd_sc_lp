* File: sky130_fd_sc_lp__mux2_2.pxi.spice
* Created: Fri Aug 28 10:43:55 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2_2%A_86_21# N_A_86_21#_M1013_d N_A_86_21#_M1010_d
+ N_A_86_21#_M1007_g N_A_86_21#_M1006_g N_A_86_21#_M1008_g N_A_86_21#_M1011_g
+ N_A_86_21#_c_82_n N_A_86_21#_c_83_n N_A_86_21#_c_161_p N_A_86_21#_c_97_p
+ N_A_86_21#_c_131_p N_A_86_21#_c_91_p N_A_86_21#_c_92_p N_A_86_21#_c_84_n
+ N_A_86_21#_c_85_n N_A_86_21#_c_98_p PM_SKY130_FD_SC_LP__MUX2_2%A_86_21#
x_PM_SKY130_FD_SC_LP__MUX2_2%A_284_279# N_A_284_279#_M1009_d
+ N_A_284_279#_M1012_d N_A_284_279#_M1001_g N_A_284_279#_M1000_g
+ N_A_284_279#_c_181_n N_A_284_279#_c_187_n N_A_284_279#_c_182_n
+ N_A_284_279#_c_183_n N_A_284_279#_c_189_n N_A_284_279#_c_190_n
+ N_A_284_279#_c_184_n N_A_284_279#_c_192_n N_A_284_279#_c_193_n
+ PM_SKY130_FD_SC_LP__MUX2_2%A_284_279#
x_PM_SKY130_FD_SC_LP__MUX2_2%A0 N_A0_M1013_g N_A0_M1004_g N_A0_c_260_n
+ N_A0_c_261_n N_A0_c_262_n A0 N_A0_c_266_n N_A0_c_263_n A0
+ PM_SKY130_FD_SC_LP__MUX2_2%A0
x_PM_SKY130_FD_SC_LP__MUX2_2%A1 N_A1_M1010_g N_A1_c_312_n N_A1_c_313_n
+ N_A1_M1005_g A1 A1 A1 N_A1_c_316_n PM_SKY130_FD_SC_LP__MUX2_2%A1
x_PM_SKY130_FD_SC_LP__MUX2_2%S N_S_c_367_n N_S_M1003_g N_S_M1002_g N_S_c_368_n
+ N_S_M1009_g N_S_c_370_n N_S_M1012_g N_S_c_371_n N_S_c_372_n S S S N_S_c_374_n
+ PM_SKY130_FD_SC_LP__MUX2_2%S
x_PM_SKY130_FD_SC_LP__MUX2_2%VPWR N_VPWR_M1006_s N_VPWR_M1011_s N_VPWR_M1002_d
+ N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n VPWR
+ N_VPWR_c_427_n N_VPWR_c_428_n N_VPWR_c_429_n N_VPWR_c_422_n N_VPWR_c_431_n
+ N_VPWR_c_432_n PM_SKY130_FD_SC_LP__MUX2_2%VPWR
x_PM_SKY130_FD_SC_LP__MUX2_2%X N_X_M1007_d N_X_M1006_d N_X_c_494_p N_X_c_475_n X
+ X X X N_X_c_476_n PM_SKY130_FD_SC_LP__MUX2_2%X
x_PM_SKY130_FD_SC_LP__MUX2_2%VGND N_VGND_M1007_s N_VGND_M1008_s N_VGND_M1003_d
+ N_VGND_c_501_n N_VGND_c_502_n N_VGND_c_503_n N_VGND_c_504_n VGND
+ N_VGND_c_505_n N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n N_VGND_c_509_n
+ N_VGND_c_510_n PM_SKY130_FD_SC_LP__MUX2_2%VGND
cc_1 VNB N_A_86_21#_M1007_g 0.0287234f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_2 VNB N_A_86_21#_M1006_g 0.00392723f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_3 VNB N_A_86_21#_M1008_g 0.0217491f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.655
cc_4 VNB N_A_86_21#_M1011_g 0.00249837f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_5 VNB N_A_86_21#_c_82_n 3.43945e-19 $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=2.515
cc_6 VNB N_A_86_21#_c_83_n 0.00986879f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.68
cc_7 VNB N_A_86_21#_c_84_n 0.0660186f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.44
cc_8 VNB N_A_86_21#_c_85_n 0.00204977f $X=-0.19 $Y=-0.245 $X2=1.052 $Y2=1.275
cc_9 VNB N_A_284_279#_M1001_g 0.0523986f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_10 VNB N_A_284_279#_c_181_n 0.00683053f $X=-0.19 $Y=-0.245 $X2=0.935
+ $Y2=0.655
cc_11 VNB N_A_284_279#_c_182_n 0.00299044f $X=-0.19 $Y=-0.245 $X2=0.935
+ $Y2=2.465
cc_12 VNB N_A_284_279#_c_183_n 0.0165438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_284_279#_c_184_n 0.0692716f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.68
cc_14 VNB N_A0_M1013_g 0.0203078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A0_c_260_n 0.00382383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A0_c_261_n 0.00560455f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_17 VNB N_A0_c_262_n 0.0329139f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_18 VNB N_A0_c_263_n 0.00498967f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=1.275
cc_19 VNB N_A1_M1010_g 0.00648344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_312_n 0.0178438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_313_n 0.00646789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_M1005_g 0.033597f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_23 VNB A1 0.00482463f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.605
cc_24 VNB N_A1_c_316_n 0.0387618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_S_c_367_n 0.0161327f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=0.24
cc_26 VNB N_S_c_368_n 0.0126523f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_27 VNB N_S_M1009_g 0.0213469f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_28 VNB N_S_c_370_n 0.0125172f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.275
cc_29 VNB N_S_c_371_n 0.0235772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_S_c_372_n 0.0101476f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=1.605
cc_31 VNB S 0.00352274f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=2.515
cc_32 VNB N_S_c_374_n 0.0502869f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=0.46
cc_33 VNB N_VPWR_c_422_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=2.68
cc_34 VNB N_X_c_475_n 0.00323438f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_35 VNB N_X_c_476_n 0.00359679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_501_n 0.0116702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_502_n 0.0491101f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_38 VNB N_VGND_c_503_n 0.00457869f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.655
cc_39 VNB N_VGND_c_504_n 0.00580583f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_40 VNB N_VGND_c_505_n 0.0175624f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=1.275
cc_41 VNB N_VGND_c_506_n 0.0410896f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.6
cc_42 VNB N_VGND_c_507_n 0.0186996f $X=-0.19 $Y=-0.245 $X2=1.052 $Y2=1.605
cc_43 VNB N_VGND_c_508_n 0.209368f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=2.6
cc_44 VNB N_VGND_c_509_n 0.00631189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_510_n 0.00632255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_A_86_21#_M1006_g 0.0272005f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_47 VPB N_A_86_21#_M1011_g 0.0216025f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_48 VPB N_A_86_21#_c_82_n 0.00126347f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=2.515
cc_49 VPB N_A_284_279#_M1000_g 0.0211451f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_50 VPB N_A_284_279#_c_181_n 0.018415f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.655
cc_51 VPB N_A_284_279#_c_187_n 0.0175692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_284_279#_c_182_n 8.50772e-19 $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_53 VPB N_A_284_279#_c_189_n 0.0203314f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=1.275
cc_54 VPB N_A_284_279#_c_190_n 5.52508e-19 $X=-0.19 $Y=1.655 $X2=1.09 $Y2=1.605
cc_55 VPB N_A_284_279#_c_184_n 0.0278589f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=0.68
cc_56 VPB N_A_284_279#_c_192_n 0.023344f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.46
cc_57 VPB N_A_284_279#_c_193_n 0.00739525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A0_M1004_g 0.0193151f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.275
cc_59 VPB N_A0_c_260_n 2.34762e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A0_c_266_n 0.0274626f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=0.765
cc_61 VPB N_A0_c_263_n 0.00502101f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=1.275
cc_62 VPB N_A1_M1010_g 0.0386534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_S_M1002_g 0.0300532f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_S_M1012_g 0.0353594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB S 0.00121317f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=2.515
cc_66 VPB N_S_c_374_n 0.0258511f $X=-0.19 $Y=1.655 $X2=2.105 $Y2=0.46
cc_67 VPB N_VPWR_c_423_n 0.0116443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_424_n 0.0650173f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_69 VPB N_VPWR_c_425_n 0.00713258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_426_n 0.00990545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_427_n 0.0150765f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=2.515
cc_72 VPB N_VPWR_c_428_n 0.0477519f $X=-0.19 $Y=1.655 $X2=2.06 $Y2=0.595
cc_73 VPB N_VPWR_c_429_n 0.0171442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_422_n 0.081029f $X=-0.19 $Y=1.655 $X2=2.25 $Y2=2.68
cc_75 VPB N_VPWR_c_431_n 0.00510188f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.44
cc_76 VPB N_VPWR_c_432_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_X_c_476_n 0.00306489f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 N_A_86_21#_M1008_g N_A_284_279#_M1001_g 0.0277005f $X=0.935 $Y=0.655 $X2=0
+ $Y2=0
cc_79 N_A_86_21#_c_83_n N_A_284_279#_M1001_g 0.0140291f $X=1.93 $Y=0.68 $X2=0
+ $Y2=0
cc_80 N_A_86_21#_c_91_p N_A_284_279#_M1001_g 0.00134074f $X=2.105 $Y=0.46 $X2=0
+ $Y2=0
cc_81 N_A_86_21#_c_92_p N_A_284_279#_M1001_g 7.53375e-19 $X=1.015 $Y=1.44 $X2=0
+ $Y2=0
cc_82 N_A_86_21#_c_84_n N_A_284_279#_M1001_g 0.00648763f $X=1.015 $Y=1.44 $X2=0
+ $Y2=0
cc_83 N_A_86_21#_c_85_n N_A_284_279#_M1001_g 0.00751047f $X=1.052 $Y=1.275 $X2=0
+ $Y2=0
cc_84 N_A_86_21#_M1011_g N_A_284_279#_M1000_g 0.0130061f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_85 N_A_86_21#_c_82_n N_A_284_279#_M1000_g 0.0036861f $X=1.09 $Y=2.515 $X2=0
+ $Y2=0
cc_86 N_A_86_21#_c_97_p N_A_284_279#_M1000_g 0.0122451f $X=2.085 $Y=2.6 $X2=0
+ $Y2=0
cc_87 N_A_86_21#_c_98_p N_A_284_279#_M1000_g 8.79113e-19 $X=2.25 $Y=2.6 $X2=0
+ $Y2=0
cc_88 N_A_86_21#_M1011_g N_A_284_279#_c_181_n 0.011665f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_89 N_A_86_21#_c_82_n N_A_284_279#_c_181_n 0.00343859f $X=1.09 $Y=2.515 $X2=0
+ $Y2=0
cc_90 N_A_86_21#_c_97_p N_A_284_279#_c_187_n 5.95576e-19 $X=2.085 $Y=2.6 $X2=0
+ $Y2=0
cc_91 N_A_86_21#_M1011_g N_A_284_279#_c_182_n 8.12315e-19 $X=0.935 $Y=2.465
+ $X2=0 $Y2=0
cc_92 N_A_86_21#_c_83_n N_A_284_279#_c_182_n 0.00904474f $X=1.93 $Y=0.68 $X2=0
+ $Y2=0
cc_93 N_A_86_21#_c_92_p N_A_284_279#_c_182_n 0.0439656f $X=1.015 $Y=1.44 $X2=0
+ $Y2=0
cc_94 N_A_86_21#_c_84_n N_A_284_279#_c_182_n 8.99284e-19 $X=1.015 $Y=1.44 $X2=0
+ $Y2=0
cc_95 N_A_86_21#_c_83_n N_A_284_279#_c_183_n 8.76872e-19 $X=1.93 $Y=0.68 $X2=0
+ $Y2=0
cc_96 N_A_86_21#_c_92_p N_A_284_279#_c_183_n 7.65238e-19 $X=1.015 $Y=1.44 $X2=0
+ $Y2=0
cc_97 N_A_86_21#_c_84_n N_A_284_279#_c_183_n 0.011537f $X=1.015 $Y=1.44 $X2=0
+ $Y2=0
cc_98 N_A_86_21#_M1010_d N_A_284_279#_c_189_n 0.00176461f $X=2.11 $Y=2.245 $X2=0
+ $Y2=0
cc_99 N_A_86_21#_c_97_p N_A_284_279#_c_189_n 0.0154453f $X=2.085 $Y=2.6 $X2=0
+ $Y2=0
cc_100 N_A_86_21#_c_98_p N_A_284_279#_c_189_n 0.0161182f $X=2.25 $Y=2.6 $X2=0
+ $Y2=0
cc_101 N_A_86_21#_M1011_g N_A_284_279#_c_190_n 6.09603e-19 $X=0.935 $Y=2.465
+ $X2=0 $Y2=0
cc_102 N_A_86_21#_c_82_n N_A_284_279#_c_190_n 0.0106803f $X=1.09 $Y=2.515 $X2=0
+ $Y2=0
cc_103 N_A_86_21#_c_97_p N_A_284_279#_c_190_n 0.0213572f $X=2.085 $Y=2.6 $X2=0
+ $Y2=0
cc_104 N_A_86_21#_c_83_n N_A0_M1013_g 0.00983426f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_105 N_A_86_21#_c_91_p N_A0_M1013_g 0.00614095f $X=2.105 $Y=0.46 $X2=0 $Y2=0
cc_106 N_A_86_21#_c_98_p N_A0_M1004_g 0.00669579f $X=2.25 $Y=2.6 $X2=0 $Y2=0
cc_107 N_A_86_21#_c_83_n N_A0_c_261_n 0.0261396f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_108 N_A_86_21#_c_85_n N_A0_c_261_n 0.00668939f $X=1.052 $Y=1.275 $X2=0 $Y2=0
cc_109 N_A_86_21#_c_83_n N_A0_c_262_n 0.00459069f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_110 N_A_86_21#_c_97_p N_A1_M1010_g 0.00829071f $X=2.085 $Y=2.6 $X2=0 $Y2=0
cc_111 N_A_86_21#_c_98_p N_A1_M1010_g 0.00430644f $X=2.25 $Y=2.6 $X2=0 $Y2=0
cc_112 N_A_86_21#_c_83_n N_A1_c_312_n 0.00134423f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_113 N_A_86_21#_c_83_n N_A1_M1005_g 0.00131627f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_114 N_A_86_21#_c_91_p N_A1_M1005_g 0.00604962f $X=2.105 $Y=0.46 $X2=0 $Y2=0
cc_115 N_A_86_21#_c_83_n A1 0.0143491f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_116 N_A_86_21#_c_91_p A1 0.00958184f $X=2.105 $Y=0.46 $X2=0 $Y2=0
cc_117 N_A_86_21#_c_98_p N_S_M1002_g 9.98726e-19 $X=2.25 $Y=2.6 $X2=0 $Y2=0
cc_118 N_A_86_21#_c_82_n N_VPWR_M1011_s 0.0077229f $X=1.09 $Y=2.515 $X2=0 $Y2=0
cc_119 N_A_86_21#_c_97_p N_VPWR_M1011_s 0.0180111f $X=2.085 $Y=2.6 $X2=0 $Y2=0
cc_120 N_A_86_21#_c_131_p N_VPWR_M1011_s 0.00114013f $X=1.175 $Y=2.6 $X2=0 $Y2=0
cc_121 N_A_86_21#_M1006_g N_VPWR_c_424_n 0.00757458f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_122 N_A_86_21#_M1006_g N_VPWR_c_425_n 5.33797e-19 $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_86_21#_M1011_g N_VPWR_c_425_n 0.00838765f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_124 N_A_86_21#_c_97_p N_VPWR_c_425_n 0.0105971f $X=2.085 $Y=2.6 $X2=0 $Y2=0
cc_125 N_A_86_21#_c_131_p N_VPWR_c_425_n 0.00939871f $X=1.175 $Y=2.6 $X2=0 $Y2=0
cc_126 N_A_86_21#_c_98_p N_VPWR_c_426_n 0.00914141f $X=2.25 $Y=2.6 $X2=0 $Y2=0
cc_127 N_A_86_21#_M1006_g N_VPWR_c_427_n 0.00585385f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_A_86_21#_M1011_g N_VPWR_c_427_n 0.00486043f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_A_86_21#_c_97_p N_VPWR_c_428_n 0.0115379f $X=2.085 $Y=2.6 $X2=0 $Y2=0
cc_130 N_A_86_21#_c_98_p N_VPWR_c_428_n 0.00725597f $X=2.25 $Y=2.6 $X2=0 $Y2=0
cc_131 N_A_86_21#_M1006_g N_VPWR_c_422_n 0.0115095f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_A_86_21#_M1011_g N_VPWR_c_422_n 0.00824727f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_86_21#_c_97_p N_VPWR_c_422_n 0.0221806f $X=2.085 $Y=2.6 $X2=0 $Y2=0
cc_134 N_A_86_21#_c_131_p N_VPWR_c_422_n 8.42036e-19 $X=1.175 $Y=2.6 $X2=0 $Y2=0
cc_135 N_A_86_21#_c_98_p N_VPWR_c_422_n 0.0107066f $X=2.25 $Y=2.6 $X2=0 $Y2=0
cc_136 N_A_86_21#_M1007_g N_X_c_475_n 0.00530663f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_137 N_A_86_21#_M1008_g N_X_c_475_n 6.89086e-19 $X=0.935 $Y=0.655 $X2=0 $Y2=0
cc_138 N_A_86_21#_c_84_n N_X_c_475_n 8.7928e-19 $X=1.015 $Y=1.44 $X2=0 $Y2=0
cc_139 N_A_86_21#_c_85_n N_X_c_475_n 0.0119101f $X=1.052 $Y=1.275 $X2=0 $Y2=0
cc_140 N_A_86_21#_c_84_n X 8.2005e-19 $X=1.015 $Y=1.44 $X2=0 $Y2=0
cc_141 N_A_86_21#_M1006_g N_X_c_476_n 0.00606647f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_86_21#_M1008_g N_X_c_476_n 0.00131346f $X=0.935 $Y=0.655 $X2=0 $Y2=0
cc_143 N_A_86_21#_M1011_g N_X_c_476_n 0.00173399f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_86_21#_c_82_n N_X_c_476_n 0.0128777f $X=1.09 $Y=2.515 $X2=0 $Y2=0
cc_145 N_A_86_21#_c_92_p N_X_c_476_n 0.0219826f $X=1.015 $Y=1.44 $X2=0 $Y2=0
cc_146 N_A_86_21#_c_84_n N_X_c_476_n 0.0263205f $X=1.015 $Y=1.44 $X2=0 $Y2=0
cc_147 N_A_86_21#_c_85_n N_X_c_476_n 0.00946172f $X=1.052 $Y=1.275 $X2=0 $Y2=0
cc_148 N_A_86_21#_c_97_p A_350_449# 0.00271391f $X=2.085 $Y=2.6 $X2=-0.19
+ $Y2=-0.245
cc_149 N_A_86_21#_c_83_n N_VGND_M1008_s 0.00883365f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_150 N_A_86_21#_c_161_p N_VGND_M1008_s 0.00113918f $X=1.175 $Y=0.68 $X2=0
+ $Y2=0
cc_151 N_A_86_21#_c_85_n N_VGND_M1008_s 0.00423273f $X=1.052 $Y=1.275 $X2=0
+ $Y2=0
cc_152 N_A_86_21#_M1007_g N_VGND_c_502_n 0.00705785f $X=0.505 $Y=0.655 $X2=0
+ $Y2=0
cc_153 N_A_86_21#_M1008_g N_VGND_c_503_n 0.00309232f $X=0.935 $Y=0.655 $X2=0
+ $Y2=0
cc_154 N_A_86_21#_c_83_n N_VGND_c_503_n 0.0149394f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_155 N_A_86_21#_c_161_p N_VGND_c_503_n 0.00897221f $X=1.175 $Y=0.68 $X2=0
+ $Y2=0
cc_156 N_A_86_21#_c_91_p N_VGND_c_503_n 0.00513201f $X=2.105 $Y=0.46 $X2=0 $Y2=0
cc_157 N_A_86_21#_M1007_g N_VGND_c_505_n 0.00585385f $X=0.505 $Y=0.655 $X2=0
+ $Y2=0
cc_158 N_A_86_21#_M1008_g N_VGND_c_505_n 0.00579836f $X=0.935 $Y=0.655 $X2=0
+ $Y2=0
cc_159 N_A_86_21#_c_161_p N_VGND_c_505_n 4.69325e-19 $X=1.175 $Y=0.68 $X2=0
+ $Y2=0
cc_160 N_A_86_21#_c_83_n N_VGND_c_506_n 0.00886543f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_161 N_A_86_21#_c_91_p N_VGND_c_506_n 0.0158128f $X=2.105 $Y=0.46 $X2=0 $Y2=0
cc_162 N_A_86_21#_M1013_d N_VGND_c_508_n 0.00856311f $X=1.955 $Y=0.24 $X2=0
+ $Y2=0
cc_163 N_A_86_21#_M1007_g N_VGND_c_508_n 0.0115095f $X=0.505 $Y=0.655 $X2=0
+ $Y2=0
cc_164 N_A_86_21#_M1008_g N_VGND_c_508_n 0.0109466f $X=0.935 $Y=0.655 $X2=0
+ $Y2=0
cc_165 N_A_86_21#_c_83_n N_VGND_c_508_n 0.0159798f $X=1.93 $Y=0.68 $X2=0 $Y2=0
cc_166 N_A_86_21#_c_161_p N_VGND_c_508_n 0.00193263f $X=1.175 $Y=0.68 $X2=0
+ $Y2=0
cc_167 N_A_86_21#_c_91_p N_VGND_c_508_n 0.00984655f $X=2.105 $Y=0.46 $X2=0 $Y2=0
cc_168 N_A_86_21#_c_83_n A_319_48# 0.00159304f $X=1.93 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_284_279#_M1001_g N_A0_M1013_g 0.0676921f $X=1.52 $Y=0.45 $X2=0 $Y2=0
cc_170 N_A_284_279#_c_189_n N_A0_M1004_g 0.0142611f $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_171 N_A_284_279#_M1001_g N_A0_c_260_n 0.00578662f $X=1.52 $Y=0.45 $X2=0 $Y2=0
cc_172 N_A_284_279#_c_182_n N_A0_c_260_n 0.0391432f $X=1.585 $Y=1.56 $X2=0 $Y2=0
cc_173 N_A_284_279#_c_183_n N_A0_c_260_n 0.00210058f $X=1.585 $Y=1.56 $X2=0
+ $Y2=0
cc_174 N_A_284_279#_c_189_n N_A0_c_260_n 0.0131148f $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_175 N_A_284_279#_M1001_g N_A0_c_261_n 0.00100222f $X=1.52 $Y=0.45 $X2=0 $Y2=0
cc_176 N_A_284_279#_c_189_n N_A0_c_266_n 0.0044365f $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_177 N_A_284_279#_c_189_n N_A0_c_263_n 0.0398695f $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_178 N_A_284_279#_c_187_n N_A1_M1010_g 0.0500949f $X=1.585 $Y=2.065 $X2=0
+ $Y2=0
cc_179 N_A_284_279#_c_189_n N_A1_M1010_g 0.0100627f $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_180 N_A_284_279#_c_189_n N_A1_c_312_n 2.5505e-19 $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_181 N_A_284_279#_c_182_n N_A1_c_313_n 0.0031015f $X=1.585 $Y=1.56 $X2=0 $Y2=0
cc_182 N_A_284_279#_c_183_n N_A1_c_313_n 0.0500949f $X=1.585 $Y=1.56 $X2=0 $Y2=0
cc_183 N_A_284_279#_c_189_n N_S_M1002_g 0.0174862f $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_184 N_A_284_279#_c_184_n N_S_M1009_g 0.00587194f $X=3.55 $Y=0.44 $X2=0 $Y2=0
cc_185 N_A_284_279#_c_189_n N_S_M1012_g 0.0180672f $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_186 N_A_284_279#_c_192_n N_S_M1012_g 2.21843e-19 $X=3.58 $Y=2.39 $X2=0 $Y2=0
cc_187 N_A_284_279#_c_184_n N_S_c_372_n 0.0441825f $X=3.55 $Y=0.44 $X2=0 $Y2=0
cc_188 N_A_284_279#_c_189_n S 0.0154051f $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_189 N_A_284_279#_c_184_n S 0.0843856f $X=3.55 $Y=0.44 $X2=0 $Y2=0
cc_190 N_A_284_279#_c_189_n N_S_c_374_n 6.08118e-19 $X=3.445 $Y=2.26 $X2=0 $Y2=0
cc_191 N_A_284_279#_c_190_n N_VPWR_M1011_s 0.00247564f $X=1.75 $Y=2.26 $X2=0
+ $Y2=0
cc_192 N_A_284_279#_c_189_n N_VPWR_M1002_d 0.00176461f $X=3.445 $Y=2.26 $X2=0
+ $Y2=0
cc_193 N_A_284_279#_M1000_g N_VPWR_c_425_n 0.00367301f $X=1.675 $Y=2.565 $X2=0
+ $Y2=0
cc_194 N_A_284_279#_c_189_n N_VPWR_c_426_n 0.0170777f $X=3.445 $Y=2.26 $X2=0
+ $Y2=0
cc_195 N_A_284_279#_c_192_n N_VPWR_c_426_n 0.0146197f $X=3.58 $Y=2.39 $X2=0
+ $Y2=0
cc_196 N_A_284_279#_M1000_g N_VPWR_c_428_n 0.00402706f $X=1.675 $Y=2.565 $X2=0
+ $Y2=0
cc_197 N_A_284_279#_c_192_n N_VPWR_c_429_n 0.00856503f $X=3.58 $Y=2.39 $X2=0
+ $Y2=0
cc_198 N_A_284_279#_M1000_g N_VPWR_c_422_n 0.0052212f $X=1.675 $Y=2.565 $X2=0
+ $Y2=0
cc_199 N_A_284_279#_c_192_n N_VPWR_c_422_n 0.00902581f $X=3.58 $Y=2.39 $X2=0
+ $Y2=0
cc_200 N_A_284_279#_c_189_n A_350_449# 0.00102299f $X=3.445 $Y=2.26 $X2=-0.19
+ $Y2=-0.245
cc_201 N_A_284_279#_c_189_n A_508_449# 0.00786004f $X=3.445 $Y=2.26 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A_284_279#_M1001_g N_VGND_c_503_n 0.00583713f $X=1.52 $Y=0.45 $X2=0
+ $Y2=0
cc_203 N_A_284_279#_M1001_g N_VGND_c_506_n 0.00414956f $X=1.52 $Y=0.45 $X2=0
+ $Y2=0
cc_204 N_A_284_279#_c_184_n N_VGND_c_507_n 0.0180131f $X=3.55 $Y=0.44 $X2=0
+ $Y2=0
cc_205 N_A_284_279#_M1009_d N_VGND_c_508_n 0.00269748f $X=3.41 $Y=0.24 $X2=0
+ $Y2=0
cc_206 N_A_284_279#_M1001_g N_VGND_c_508_n 0.00600042f $X=1.52 $Y=0.45 $X2=0
+ $Y2=0
cc_207 N_A_284_279#_c_184_n N_VGND_c_508_n 0.0114738f $X=3.55 $Y=0.44 $X2=0
+ $Y2=0
cc_208 N_A0_M1004_g N_A1_M1010_g 0.0261519f $X=2.465 $Y=2.565 $X2=0 $Y2=0
cc_209 N_A0_c_260_n N_A1_M1010_g 0.0176509f $X=2.05 $Y=1.55 $X2=0 $Y2=0
cc_210 N_A0_c_266_n N_A1_M1010_g 0.0215387f $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_211 N_A0_c_260_n N_A1_c_312_n 0.00723334f $X=2.05 $Y=1.55 $X2=0 $Y2=0
cc_212 N_A0_c_266_n N_A1_c_312_n 0.0112535f $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_213 N_A0_c_263_n N_A1_c_312_n 0.0109858f $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_214 N_A0_c_260_n N_A1_c_313_n 0.00416632f $X=2.05 $Y=1.55 $X2=0 $Y2=0
cc_215 N_A0_c_262_n N_A1_c_313_n 0.0113732f $X=1.97 $Y=1.02 $X2=0 $Y2=0
cc_216 N_A0_M1013_g N_A1_M1005_g 0.0152182f $X=1.88 $Y=0.45 $X2=0 $Y2=0
cc_217 N_A0_c_261_n N_A1_M1005_g 7.88859e-19 $X=1.97 $Y=1.02 $X2=0 $Y2=0
cc_218 N_A0_c_262_n N_A1_M1005_g 0.0196805f $X=1.97 $Y=1.02 $X2=0 $Y2=0
cc_219 N_A0_M1013_g A1 6.52706e-19 $X=1.88 $Y=0.45 $X2=0 $Y2=0
cc_220 N_A0_c_261_n A1 0.0270768f $X=1.97 $Y=1.02 $X2=0 $Y2=0
cc_221 N_A0_c_262_n A1 0.0013991f $X=1.97 $Y=1.02 $X2=0 $Y2=0
cc_222 N_A0_c_266_n A1 2.1419e-19 $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_223 N_A0_c_263_n A1 0.0248491f $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_224 N_A0_c_260_n N_A1_c_316_n 0.00486777f $X=2.05 $Y=1.55 $X2=0 $Y2=0
cc_225 N_A0_c_266_n N_A1_c_316_n 0.00615004f $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_226 N_A0_c_263_n N_A1_c_316_n 0.0012601f $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_227 N_A0_M1004_g N_S_M1002_g 0.0362959f $X=2.465 $Y=2.565 $X2=0 $Y2=0
cc_228 N_A0_c_263_n S 0.015853f $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_229 N_A0_c_266_n N_S_c_374_n 0.0210467f $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_230 N_A0_c_263_n N_S_c_374_n 0.0066328f $X=2.485 $Y=1.92 $X2=0 $Y2=0
cc_231 N_A0_M1004_g N_VPWR_c_426_n 0.00181332f $X=2.465 $Y=2.565 $X2=0 $Y2=0
cc_232 N_A0_M1004_g N_VPWR_c_428_n 0.00502121f $X=2.465 $Y=2.565 $X2=0 $Y2=0
cc_233 N_A0_M1004_g N_VPWR_c_422_n 0.0052212f $X=2.465 $Y=2.565 $X2=0 $Y2=0
cc_234 N_A0_M1013_g N_VGND_c_506_n 0.00406358f $X=1.88 $Y=0.45 $X2=0 $Y2=0
cc_235 N_A0_M1013_g N_VGND_c_508_n 0.00589678f $X=1.88 $Y=0.45 $X2=0 $Y2=0
cc_236 N_A1_M1005_g N_S_c_367_n 0.051636f $X=2.42 $Y=0.45 $X2=-0.19 $Y2=-0.245
cc_237 A1 N_S_c_367_n 0.00791311f $X=2.555 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_238 N_A1_M1005_g N_S_c_368_n 0.00502219f $X=2.42 $Y=0.45 $X2=0 $Y2=0
cc_239 A1 N_S_c_368_n 0.00334389f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_240 N_A1_c_316_n N_S_c_368_n 0.0218337f $X=2.525 $Y=1.295 $X2=0 $Y2=0
cc_241 A1 N_S_M1009_g 7.94872e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_242 A1 N_S_c_371_n 0.00478559f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_243 N_A1_M1005_g S 2.62572e-19 $X=2.42 $Y=0.45 $X2=0 $Y2=0
cc_244 A1 S 0.0385141f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_245 N_A1_c_316_n S 0.00131793f $X=2.525 $Y=1.295 $X2=0 $Y2=0
cc_246 N_A1_c_316_n N_S_c_374_n 0.00316822f $X=2.525 $Y=1.295 $X2=0 $Y2=0
cc_247 N_A1_M1010_g N_VPWR_c_428_n 0.00401048f $X=2.035 $Y=2.565 $X2=0 $Y2=0
cc_248 N_A1_M1010_g N_VPWR_c_422_n 0.0052212f $X=2.035 $Y=2.565 $X2=0 $Y2=0
cc_249 N_A1_M1005_g N_VGND_c_506_n 0.00414516f $X=2.42 $Y=0.45 $X2=0 $Y2=0
cc_250 A1 N_VGND_c_506_n 0.00900946f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_251 N_A1_M1005_g N_VGND_c_508_n 0.00628744f $X=2.42 $Y=0.45 $X2=0 $Y2=0
cc_252 A1 N_VGND_c_508_n 0.0119235f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_253 A1 A_499_48# 0.00139886f $X=2.555 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_254 N_S_M1002_g N_VPWR_c_426_n 0.0121409f $X=2.935 $Y=2.565 $X2=0 $Y2=0
cc_255 N_S_M1012_g N_VPWR_c_426_n 0.0121445f $X=3.365 $Y=2.565 $X2=0 $Y2=0
cc_256 N_S_M1002_g N_VPWR_c_428_n 0.00435433f $X=2.935 $Y=2.565 $X2=0 $Y2=0
cc_257 N_S_M1012_g N_VPWR_c_429_n 0.00435433f $X=3.365 $Y=2.565 $X2=0 $Y2=0
cc_258 N_S_M1002_g N_VPWR_c_422_n 0.00438581f $X=2.935 $Y=2.565 $X2=0 $Y2=0
cc_259 N_S_M1012_g N_VPWR_c_422_n 0.0043858f $X=3.365 $Y=2.565 $X2=0 $Y2=0
cc_260 N_S_c_367_n N_VGND_c_504_n 0.00525435f $X=2.78 $Y=0.77 $X2=0 $Y2=0
cc_261 N_S_M1009_g N_VGND_c_504_n 0.00331318f $X=3.335 $Y=0.45 $X2=0 $Y2=0
cc_262 N_S_c_371_n N_VGND_c_504_n 0.00490739f $X=2.975 $Y=0.845 $X2=0 $Y2=0
cc_263 S N_VGND_c_504_n 0.0230334f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_264 N_S_c_374_n N_VGND_c_504_n 2.08436e-19 $X=3.12 $Y=1.345 $X2=0 $Y2=0
cc_265 N_S_c_367_n N_VGND_c_506_n 0.00544382f $X=2.78 $Y=0.77 $X2=0 $Y2=0
cc_266 N_S_c_371_n N_VGND_c_506_n 7.88586e-19 $X=2.975 $Y=0.845 $X2=0 $Y2=0
cc_267 N_S_M1009_g N_VGND_c_507_n 0.0058025f $X=3.335 $Y=0.45 $X2=0 $Y2=0
cc_268 N_S_c_367_n N_VGND_c_508_n 0.0099026f $X=2.78 $Y=0.77 $X2=0 $Y2=0
cc_269 N_S_M1009_g N_VGND_c_508_n 0.0115476f $X=3.335 $Y=0.45 $X2=0 $Y2=0
cc_270 N_S_c_371_n N_VGND_c_508_n 0.00109002f $X=2.975 $Y=0.845 $X2=0 $Y2=0
cc_271 N_S_c_372_n N_VGND_c_508_n 7.77756e-19 $X=3.35 $Y=0.94 $X2=0 $Y2=0
cc_272 S N_VGND_c_508_n 0.00257153f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_273 N_VPWR_c_422_n N_X_M1006_d 0.0041489f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_274 N_VPWR_c_427_n X 0.0136943f $X=0.985 $Y=3.33 $X2=0 $Y2=0
cc_275 N_VPWR_c_422_n X 0.00866444f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_276 N_VPWR_c_424_n N_X_c_476_n 0.045553f $X=0.29 $Y=1.98 $X2=0 $Y2=0
cc_277 N_X_c_494_p N_VGND_c_502_n 0.0295012f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_278 N_X_c_494_p N_VGND_c_505_n 0.0147587f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_279 N_X_M1007_d N_VGND_c_508_n 0.00310528f $X=0.58 $Y=0.235 $X2=0 $Y2=0
cc_280 N_X_c_494_p N_VGND_c_508_n 0.00983606f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_281 N_VGND_c_508_n A_319_48# 0.0023229f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_282 N_VGND_c_508_n A_499_48# 0.00198436f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
