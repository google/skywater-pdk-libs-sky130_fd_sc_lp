* File: sky130_fd_sc_lp__or4_m.pex.spice
* Created: Fri Aug 28 11:25:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4_M%D 1 5 9 14 16 18 19 20 21 22 29
r31 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r32 21 22 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r33 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r34 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r35 19 30 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.12
r36 18 30 10.8136 $w=1.98e-07 $l=1.95e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.12
r37 16 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.27 $Y2=1.12
r38 16 17 46.7501 $w=3.3e-07 $l=2.97405e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.285 $Y2=1.75
r39 12 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.105
+ $X2=0.27 $Y2=1.12
r40 12 14 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=0.27 $Y=1.03
+ $X2=0.625 $Y2=1.03
r41 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.92 $Y=1.825 $X2=0.92
+ $Y2=2.195
r42 3 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.625 $Y=0.955
+ $X2=0.625 $Y2=1.03
r43 3 5 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.625 $Y=0.955
+ $X2=0.625 $Y2=0.445
r44 2 17 12.8954 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.435 $Y=1.75
+ $X2=0.285 $Y2=1.75
r45 1 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.845 $Y=1.75
+ $X2=0.92 $Y2=1.825
r46 1 2 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.845 $Y=1.75
+ $X2=0.435 $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_M%C 3 5 8 10 11 12 13 18 20
r39 18 20 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.167 $Y=0.93
+ $X2=1.167 $Y2=0.765
r40 12 13 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=0.925
+ $X2=1.195 $Y2=1.295
r41 12 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.19
+ $Y=0.93 $X2=1.19 $Y2=0.93
r42 11 12 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=0.555
+ $X2=1.195 $Y2=0.925
r43 8 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.28 $Y=2.195
+ $X2=1.28 $Y2=1.435
r44 5 10 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=1.167 $Y=1.248
+ $X2=1.167 $Y2=1.435
r45 4 18 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=1.167 $Y=0.952
+ $X2=1.167 $Y2=0.93
r46 4 5 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=1.167 $Y=0.952
+ $X2=1.167 $Y2=1.248
r47 3 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.055 $Y=0.445
+ $X2=1.055 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_M%B 2 5 9 10 11 12 16 18
r39 16 18 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.742 $Y=0.93
+ $X2=1.742 $Y2=0.765
r40 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.73 $Y=0.925
+ $X2=1.73 $Y2=1.295
r41 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=0.93 $X2=1.73 $Y2=0.93
r42 9 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.845 $Y=0.445
+ $X2=1.845 $Y2=0.765
r43 5 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.64 $Y=2.195
+ $X2=1.64 $Y2=1.435
r44 2 10 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=1.742 $Y=1.258
+ $X2=1.742 $Y2=1.435
r45 1 16 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=1.742 $Y=0.942
+ $X2=1.742 $Y2=0.93
r46 1 2 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=1.742 $Y=0.942
+ $X2=1.742 $Y2=1.258
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_M%A 1 3 7 11 14 17 18
c45 7 0 5.77162e-20 $X=2.275 $Y=0.445
r46 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.295
+ $Y=1.085 $X2=2.295 $Y2=1.085
r47 14 18 3.16609 $w=5.08e-07 $l=1.35e-07 $layer=LI1_cond $X=2.16 $Y=1.255
+ $X2=2.295 $Y2=1.255
r48 13 17 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=0.92
+ $X2=2.295 $Y2=1.085
r49 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.295 $Y=1.425
+ $X2=2.295 $Y2=1.085
r50 7 13 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=2.275 $Y=0.445
+ $X2=2.275 $Y2=0.92
r51 1 11 63.1956 $w=2.25e-07 $l=5.27257e-07 $layer=POLY_cond $X=2 $Y=1.825
+ $X2=2.295 $Y2=1.425
r52 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2 $Y=1.825 $X2=2
+ $Y2=2.195
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_M%A_116_397# 1 2 3 10 15 18 22 26 28 32 37 39 41
+ 42 44 45 48 49
r100 45 47 11.5094 $w=2.65e-07 $l=2.5e-07 $layer=LI1_cond $X=0.762 $Y=1.88
+ $X2=0.762 $Y2=2.13
r101 43 44 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=2.725 $Y=0.82
+ $X2=2.725 $Y2=1.795
r102 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.64 $Y=0.735
+ $X2=2.725 $Y2=0.82
r103 41 42 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.64 $Y=0.735
+ $X2=2.245 $Y2=0.735
r104 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=1.88
+ $X2=1.94 $Y2=1.88
r105 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.64 $Y=1.88
+ $X2=2.725 $Y2=1.795
r106 39 40 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.64 $Y=1.88
+ $X2=2.105 $Y2=1.88
r107 35 42 17.761 $w=9e-08 $l=1.72337e-07 $layer=LI1_cond $X=2.11 $Y=0.65
+ $X2=2.245 $Y2=0.735
r108 35 37 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.11 $Y=0.65
+ $X2=2.11 $Y2=0.495
r109 33 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.94 $Y=2.94 $X2=1.94
+ $Y2=2.85
r110 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=2.94 $X2=1.94 $Y2=2.94
r111 30 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=1.965
+ $X2=1.94 $Y2=1.88
r112 30 32 34.0495 $w=3.28e-07 $l=9.75e-07 $layer=LI1_cond $X=1.94 $Y=1.965
+ $X2=1.94 $Y2=2.94
r113 29 45 3.33486 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=0.925 $Y=1.88
+ $X2=0.762 $Y2=1.88
r114 28 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.775 $Y=1.88
+ $X2=1.94 $Y2=1.88
r115 28 29 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.775 $Y=1.88
+ $X2=0.925 $Y2=1.88
r116 24 45 4.90929 $w=2.65e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.83 $Y=1.795
+ $X2=0.762 $Y2=1.88
r117 24 26 75.0096 $w=1.88e-07 $l=1.285e-06 $layer=LI1_cond $X=0.83 $Y=1.795
+ $X2=0.83 $Y2=0.51
r118 20 22 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.745 $Y=1.8
+ $X2=2.885 $Y2=1.8
r119 16 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=1.725
+ $X2=2.885 $Y2=1.8
r120 16 18 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=2.885 $Y=1.725
+ $X2=2.885 $Y2=0.445
r121 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.745 $Y=2.775
+ $X2=2.745 $Y2=2.195
r122 12 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.745 $Y=1.875
+ $X2=2.745 $Y2=1.8
r123 12 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.745 $Y=1.875
+ $X2=2.745 $Y2=2.195
r124 11 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.105 $Y=2.85
+ $X2=1.94 $Y2=2.85
r125 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.67 $Y=2.85
+ $X2=2.745 $Y2=2.775
r126 10 11 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.67 $Y=2.85
+ $X2=2.105 $Y2=2.85
r127 3 47 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.985 $X2=0.705 $Y2=2.13
r128 2 37 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.235 $X2=2.06 $Y2=0.495
r129 1 26 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.7
+ $Y=0.235 $X2=0.84 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_M%VPWR 1 6 9 10 11 21 22
r26 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r27 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r28 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 14 18 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 11 15 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 9 18 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.45 $Y2=3.33
r35 8 21 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=2.45 $Y2=3.33
r37 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=3.245 $X2=2.45
+ $Y2=3.33
r38 4 6 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=2.45 $Y=3.245
+ $X2=2.45 $Y2=2.26
r39 1 6 600 $w=1.7e-07 $l=4.9371e-07 $layer=licon1_PDIFF $count=1 $X=2.075
+ $Y=1.985 $X2=2.45 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_M%X 1 2 7 8 9 10 11 12 13 35 43
c20 43 0 5.77162e-20 $X=3.1 $Y=0.385
r21 35 36 5.79586 $w=4.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.03 $Y=2.26
+ $X2=3.03 $Y2=2.155
r22 12 13 9.41594 $w=4.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.03 $Y=2.405
+ $X2=3.03 $Y2=2.775
r23 12 35 3.69003 $w=4.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.03 $Y=2.405
+ $X2=3.03 $Y2=2.26
r24 11 36 6.01275 $w=2.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.15 $Y=2.035
+ $X2=3.15 $Y2=2.155
r25 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.15 $Y=1.665
+ $X2=3.15 $Y2=2.035
r26 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.15 $Y=1.295
+ $X2=3.15 $Y2=1.665
r27 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.15 $Y=0.925 $X2=3.15
+ $Y2=1.295
r28 7 43 2.83598 $w=3.98e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.47 $X2=3.1
+ $Y2=0.385
r29 7 8 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.15 $Y=0.555 $X2=3.15
+ $Y2=0.925
r30 2 35 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.82
+ $Y=1.985 $X2=2.96 $Y2=2.26
r31 1 43 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_M%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r53 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 37 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r56 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=2.59
+ $Y2=0
r58 34 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=3.12
+ $Y2=0
r59 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r60 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r61 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=1.63
+ $Y2=0
r62 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=2.16
+ $Y2=0
r63 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.59
+ $Y2=0
r64 29 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.16
+ $Y2=0
r65 28 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r66 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r67 25 40 4.53571 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.277
+ $Y2=0
r68 25 27 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=1.2
+ $Y2=0
r69 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.63
+ $Y2=0
r70 24 27 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.2
+ $Y2=0
r71 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r72 22 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r73 22 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0
r75 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0.36
r76 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0
r77 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0.38
r78 10 40 3.23047 $w=3.3e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.39 $Y=0.085
+ $X2=0.277 $Y2=0
r79 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.39 $Y=0.085
+ $X2=0.39 $Y2=0.38
r80 3 20 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.235 $X2=2.59 $Y2=0.36
r81 2 16 182 $w=1.7e-07 $l=5.67891e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.63 $Y2=0.38
r82 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.265
+ $Y=0.235 $X2=0.39 $Y2=0.38
.ends

