# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand2_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__nand2_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.440000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.189000 ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.930000 0.905000 1.220000 1.180000 ;
        RECT 0.930000 1.180000 1.315000 1.575000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.189000 ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.955000 0.400000 2.890000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.237300 ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 0.555000 1.300000 0.725000 ;
        RECT 0.580000 0.725000 0.750000 1.815000 ;
        RECT 0.580000 1.815000 1.315000 2.275000 ;
        RECT 0.970000 0.265000 1.300000 0.555000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.440000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.440000 0.085000 ;
      RECT 0.000000  3.245000 1.440000 3.415000 ;
      RECT 0.150000  0.085000 0.400000 0.725000 ;
      RECT 0.580000  2.505000 0.910000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
  END
END sky130_fd_sc_lp__nand2_lp
END LIBRARY
