* File: sky130_fd_sc_lp__nor2b_4.pex.spice
* Created: Wed Sep  2 10:08:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2B_4%B_N 3 7 9 10 11 15
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.46 $X2=0.27 $Y2=1.46
r29 11 15 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=1.46
r30 9 14 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=0.565 $Y=1.46
+ $X2=0.27 $Y2=1.46
r31 9 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.565 $Y=1.46
+ $X2=0.64 $Y2=1.46
r32 5 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=1.625
+ $X2=0.64 $Y2=1.46
r33 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.64 $Y=1.625 $X2=0.64
+ $Y2=2.465
r34 1 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.46
r35 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.64 $Y=1.295 $X2=0.64
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_4%A 3 7 11 15 19 23 27 31 37 38 41 42 46 47 48
+ 49 62 67 68 75
c158 62 0 1.143e-19 $X=2.87 $Y=1.51
c159 27 0 1.96167e-19 $X=4.16 $Y=0.655
r160 61 68 6.41701 $w=4.38e-07 $l=2.45e-07 $layer=LI1_cond $X=2.53 $Y=1.645
+ $X2=2.285 $Y2=1.645
r161 60 62 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.53 $Y=1.51
+ $X2=2.87 $Y2=1.51
r162 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.51 $X2=2.53 $Y2=1.51
r163 57 60 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.44 $Y=1.51 $X2=2.53
+ $Y2=1.51
r164 49 67 3.5359 $w=4.38e-07 $l=1.35e-07 $layer=LI1_cond $X=3.12 $Y=1.645
+ $X2=2.985 $Y2=1.645
r165 48 67 9.0362 $w=4.38e-07 $l=3.45e-07 $layer=LI1_cond $X=2.64 $Y=1.645
+ $X2=2.985 $Y2=1.645
r166 48 61 2.88111 $w=4.38e-07 $l=1.1e-07 $layer=LI1_cond $X=2.64 $Y=1.645
+ $X2=2.53 $Y2=1.645
r167 47 68 3.27399 $w=4.38e-07 $l=1.25e-07 $layer=LI1_cond $X=2.16 $Y=1.645
+ $X2=2.285 $Y2=1.645
r168 47 75 7.00188 $w=4.38e-07 $l=9.5e-08 $layer=LI1_cond $X=2.16 $Y=1.645
+ $X2=2.065 $Y2=1.645
r169 46 49 43.7401 $w=2.23e-07 $l=8.4e-07 $layer=LI1_cond $X=4.045 $Y=1.78
+ $X2=3.205 $Y2=1.78
r170 42 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.51
+ $X2=1.13 $Y2=1.675
r171 42 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.51
+ $X2=1.13 $Y2=1.345
r172 41 44 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.13 $Y=1.51
+ $X2=1.13 $Y2=1.78
r173 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.51 $X2=1.13 $Y2=1.51
r174 38 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.51
+ $X2=4.21 $Y2=1.675
r175 38 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.51
+ $X2=4.21 $Y2=1.345
r176 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.51 $X2=4.21 $Y2=1.51
r177 35 46 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.175 $Y=1.695
+ $X2=4.045 $Y2=1.78
r178 35 37 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=4.175 $Y=1.695
+ $X2=4.175 $Y2=1.51
r179 34 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=1.78
+ $X2=1.13 $Y2=1.78
r180 34 75 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.295 $Y=1.78
+ $X2=2.065 $Y2=1.78
r181 31 66 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.16 $Y=2.465
+ $X2=4.16 $Y2=1.675
r182 27 65 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.16 $Y=0.655
+ $X2=4.16 $Y2=1.345
r183 21 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.87 $Y=1.675
+ $X2=2.87 $Y2=1.51
r184 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.87 $Y=1.675
+ $X2=2.87 $Y2=2.465
r185 17 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.87 $Y=1.345
+ $X2=2.87 $Y2=1.51
r186 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.87 $Y=1.345
+ $X2=2.87 $Y2=0.655
r187 13 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.44 $Y=1.675
+ $X2=2.44 $Y2=1.51
r188 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.44 $Y=1.675
+ $X2=2.44 $Y2=2.465
r189 9 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.44 $Y=1.345
+ $X2=2.44 $Y2=1.51
r190 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.44 $Y=1.345
+ $X2=2.44 $Y2=0.655
r191 7 56 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.15 $Y=2.465
+ $X2=1.15 $Y2=1.675
r192 3 55 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.15 $Y=0.655
+ $X2=1.15 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_4%A_60_47# 1 2 7 9 12 14 16 19 21 23 26 28 30
+ 33 37 41 44 45 46 47 54 56 62 71 76
c160 62 0 6.01393e-20 $X=3.505 $Y=1.17
c161 56 0 5.41602e-20 $X=1.73 $Y=1.17
r162 66 76 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=3.47 $Y=1.35
+ $X2=3.73 $Y2=1.35
r163 66 73 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=3.47 $Y=1.35
+ $X2=3.3 $Y2=1.35
r164 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.47
+ $Y=1.35 $X2=3.47 $Y2=1.35
r165 62 65 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=3.505 $Y=1.17
+ $X2=3.505 $Y2=1.35
r166 60 71 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=1.73 $Y=1.35
+ $X2=2.01 $Y2=1.35
r167 60 68 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.73 $Y=1.35
+ $X2=1.58 $Y2=1.35
r168 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.35 $X2=1.73 $Y2=1.35
r169 56 59 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.73 $Y=1.17
+ $X2=1.73 $Y2=1.35
r170 48 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=1.17
+ $X2=1.73 $Y2=1.17
r171 47 62 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.375 $Y=1.17
+ $X2=3.505 $Y2=1.17
r172 47 48 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=3.375 $Y=1.17
+ $X2=1.895 $Y2=1.17
r173 46 50 5.55076 $w=1.95e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.785 $Y=1.17
+ $X2=0.7 $Y2=1.13
r174 45 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=1.17
+ $X2=1.73 $Y2=1.17
r175 45 46 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.565 $Y=1.17
+ $X2=0.785 $Y2=1.17
r176 44 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.93 $X2=0.7
+ $Y2=2.015
r177 43 50 1.54022 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.7 $Y=1.255
+ $X2=0.7 $Y2=1.13
r178 43 44 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.7 $Y=1.255
+ $X2=0.7 $Y2=1.93
r179 39 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.395 $Y=2.015
+ $X2=0.7 $Y2=2.015
r180 39 41 34.5733 $w=2.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.395 $Y=2.1
+ $X2=0.395 $Y2=2.91
r181 35 50 19.3949 $w=1.95e-07 $l=3.1e-07 $layer=LI1_cond $X=0.39 $Y=1.13
+ $X2=0.7 $Y2=1.13
r182 35 37 25.93 $w=2.58e-07 $l=5.85e-07 $layer=LI1_cond $X=0.39 $Y=1.005
+ $X2=0.39 $Y2=0.42
r183 31 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.515
+ $X2=3.73 $Y2=1.35
r184 31 33 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.73 $Y=1.515
+ $X2=3.73 $Y2=2.465
r185 28 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.185
+ $X2=3.73 $Y2=1.35
r186 28 30 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.73 $Y=1.185
+ $X2=3.73 $Y2=0.655
r187 24 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.515
+ $X2=3.3 $Y2=1.35
r188 24 26 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.3 $Y=1.515
+ $X2=3.3 $Y2=2.465
r189 21 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.185
+ $X2=3.3 $Y2=1.35
r190 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.3 $Y=1.185
+ $X2=3.3 $Y2=0.655
r191 17 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.515
+ $X2=2.01 $Y2=1.35
r192 17 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.01 $Y=1.515
+ $X2=2.01 $Y2=2.465
r193 14 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.01 $Y=1.185
+ $X2=2.01 $Y2=1.35
r194 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.01 $Y=1.185
+ $X2=2.01 $Y2=0.655
r195 10 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=1.35
r196 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=2.465
r197 7 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.185
+ $X2=1.58 $Y2=1.35
r198 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.58 $Y=1.185
+ $X2=1.58 $Y2=0.655
r199 2 39 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.835 $X2=0.425 $Y2=2.095
r200 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.835 $X2=0.425 $Y2=2.91
r201 1 37 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.3
+ $Y=0.235 $X2=0.425 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_4%VPWR 1 2 3 13 16 18 20 23 28 29 30 36 45
r73 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r74 42 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 41 42 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 38 41 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.08 $Y2=3.33
r77 38 39 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r78 36 44 4.4922 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.21 $Y=3.33
+ $X2=4.505 $Y2=3.33
r79 36 41 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.21 $Y=3.33
+ $X2=4.08 $Y2=3.33
r80 34 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r81 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r82 30 42 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=4.08 $Y2=3.33
r83 30 39 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r84 28 33 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.75 $Y=3.33 $X2=0.72
+ $Y2=3.33
r85 28 29 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.75 $Y=3.33 $X2=0.89
+ $Y2=3.33
r86 27 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.03 $Y=3.33 $X2=1.2
+ $Y2=3.33
r87 27 29 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.03 $Y=3.33 $X2=0.89
+ $Y2=3.33
r88 25 26 4.31382 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.915 $Y=2.54
+ $X2=0.915 $Y2=2.655
r89 23 25 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.915 $Y=2.38
+ $X2=0.915 $Y2=2.54
r90 18 44 3.27398 $w=3.3e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.375 $Y=3.245
+ $X2=4.505 $Y2=3.33
r91 18 20 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=4.375 $Y=3.245
+ $X2=4.375 $Y2=2.475
r92 14 25 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=2.54
+ $X2=0.915 $Y2=2.54
r93 14 16 78.9173 $w=2.28e-07 $l=1.575e-06 $layer=LI1_cond $X=1.08 $Y=2.54
+ $X2=2.655 $Y2=2.54
r94 13 26 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.89 $Y=2.95
+ $X2=0.89 $Y2=2.655
r95 11 29 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=3.33
r96 11 13 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=2.95
r97 3 20 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=4.235
+ $Y=1.835 $X2=4.375 $Y2=2.475
r98 2 16 600 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.835 $X2=2.655 $Y2=2.55
r99 1 23 600 $w=1.7e-07 $l=6.37201e-07 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=1.835 $X2=0.915 $Y2=2.38
r100 1 13 600 $w=1.7e-07 $l=1.21088e-06 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=1.835 $X2=0.915 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_4%A_245_367# 1 2 3 4 13 21 23 27 29
r36 25 27 19.1318 $w=1.98e-07 $l=3.45e-07 $layer=LI1_cond $X=3.94 $Y=2.885
+ $X2=3.94 $Y2=2.54
r37 24 29 4.95952 $w=2.1e-07 $l=1.14018e-07 $layer=LI1_cond $X=3.19 $Y=2.975
+ $X2=3.09 $Y2=2.945
r38 23 25 6.84108 $w=1.8e-07 $l=1.3784e-07 $layer=LI1_cond $X=3.84 $Y=2.975
+ $X2=3.94 $Y2=2.885
r39 23 24 40.0505 $w=1.78e-07 $l=6.5e-07 $layer=LI1_cond $X=3.84 $Y=2.975
+ $X2=3.19 $Y2=2.975
r40 19 29 1.51883 $w=2e-07 $l=1.2e-07 $layer=LI1_cond $X=3.09 $Y=2.825 $X2=3.09
+ $Y2=2.945
r41 19 21 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=3.09 $Y=2.825
+ $X2=3.09 $Y2=2.54
r42 15 18 41.2959 $w=2.38e-07 $l=8.6e-07 $layer=LI1_cond $X=1.365 $Y=2.945
+ $X2=2.225 $Y2=2.945
r43 13 29 4.95952 $w=2.1e-07 $l=1e-07 $layer=LI1_cond $X=2.99 $Y=2.945 $X2=3.09
+ $Y2=2.945
r44 13 18 36.7341 $w=2.38e-07 $l=7.65e-07 $layer=LI1_cond $X=2.99 $Y=2.945
+ $X2=2.225 $Y2=2.945
r45 4 27 300 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_PDIFF $count=2 $X=3.805
+ $Y=1.835 $X2=3.945 $Y2=2.54
r46 3 21 300 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_PDIFF $count=2 $X=2.945
+ $Y=1.835 $X2=3.085 $Y2=2.54
r47 2 18 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.085
+ $Y=1.835 $X2=2.225 $Y2=2.95
r48 1 15 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=1.835 $X2=1.365 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_4%Y 1 2 3 4 5 6 21 23 24 25 29 31 35 37 41 45
+ 47 52 53 54 56 57 64 65 66
c117 57 0 1.96167e-19 $X=3.935 $Y=0.83
r118 65 66 16.7488 $w=2.23e-07 $l=3.27e-07 $layer=LI1_cond $X=4.587 $Y=1.665
+ $X2=4.587 $Y2=1.992
r119 64 65 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=4.587 $Y=1.295
+ $X2=4.587 $Y2=1.665
r120 63 64 6.14636 $w=2.23e-07 $l=1.2e-07 $layer=LI1_cond $X=4.587 $Y=1.175
+ $X2=4.587 $Y2=1.295
r121 60 61 9.33971 $w=1.88e-07 $l=1.6e-07 $layer=LI1_cond $X=3.935 $Y=0.93
+ $X2=3.935 $Y2=1.09
r122 57 60 5.83732 $w=1.88e-07 $l=1e-07 $layer=LI1_cond $X=3.935 $Y=0.83
+ $X2=3.935 $Y2=0.93
r123 57 58 5.00416 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=0.83
+ $X2=3.935 $Y2=0.745
r124 55 66 39.9242 $w=2.53e-07 $l=8.55e-07 $layer=LI1_cond $X=3.62 $Y=2.12
+ $X2=4.475 $Y2=2.12
r125 55 56 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.62 $Y=2.12
+ $X2=3.515 $Y2=2.12
r126 50 52 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=2.145
+ $X2=1.96 $Y2=2.145
r127 48 61 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.03 $Y=1.09 $X2=3.935
+ $Y2=1.09
r128 47 63 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.475 $Y=1.09
+ $X2=4.587 $Y2=1.175
r129 47 48 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=4.475 $Y=1.09
+ $X2=4.03 $Y2=1.09
r130 45 58 20.0253 $w=1.78e-07 $l=3.25e-07 $layer=LI1_cond $X=3.94 $Y=0.42
+ $X2=3.94 $Y2=0.745
r131 39 56 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=2.205
+ $X2=3.515 $Y2=2.12
r132 39 41 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=3.515 $Y=2.205
+ $X2=3.515 $Y2=2.21
r133 38 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=0.83
+ $X2=3.085 $Y2=0.83
r134 37 57 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.84 $Y=0.83 $X2=3.935
+ $Y2=0.83
r135 37 38 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.84 $Y=0.83
+ $X2=3.25 $Y2=0.83
r136 33 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.745
+ $X2=3.085 $Y2=0.83
r137 33 35 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.085 $Y=0.745
+ $X2=3.085 $Y2=0.42
r138 32 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=0.83
+ $X2=2.225 $Y2=0.83
r139 31 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=0.83
+ $X2=3.085 $Y2=0.83
r140 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.92 $Y=0.83
+ $X2=2.39 $Y2=0.83
r141 27 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0.745
+ $X2=2.225 $Y2=0.83
r142 27 29 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.225 $Y=0.745
+ $X2=2.225 $Y2=0.42
r143 25 56 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.41 $Y=2.12
+ $X2=3.515 $Y2=2.12
r144 25 52 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=3.41 $Y=2.12
+ $X2=1.96 $Y2=2.12
r145 23 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=0.83
+ $X2=2.225 $Y2=0.83
r146 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.06 $Y=0.83
+ $X2=1.53 $Y2=0.83
r147 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.365 $Y=0.745
+ $X2=1.53 $Y2=0.83
r148 19 21 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.365 $Y=0.745
+ $X2=1.365 $Y2=0.42
r149 6 41 300 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=2 $X=3.375
+ $Y=1.835 $X2=3.515 $Y2=2.21
r150 5 50 600 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=1.835 $X2=1.795 $Y2=2.15
r151 4 60 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.805
+ $Y=0.235 $X2=3.945 $Y2=0.93
r152 4 45 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.805
+ $Y=0.235 $X2=3.945 $Y2=0.42
r153 3 35 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.235 $X2=3.085 $Y2=0.42
r154 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.085
+ $Y=0.235 $X2=2.225 $Y2=0.42
r155 1 21 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.225
+ $Y=0.235 $X2=1.365 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2B_4%VGND 1 2 3 4 5 20 24 26 30 34 36 38 40 41 43
+ 44 45 55 60 63 67
r80 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r81 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r82 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r83 58 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r84 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r85 55 66 4.4922 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.505
+ $Y2=0
r86 55 57 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.08
+ $Y2=0
r87 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r88 54 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r89 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r90 51 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.655
+ $Y2=0
r91 51 53 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=3.12
+ $Y2=0
r92 50 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r93 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r94 47 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=0.855
+ $Y2=0
r95 47 49 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.02 $Y=0 $X2=1.68
+ $Y2=0
r96 45 64 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r97 45 50 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r98 43 53 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.12
+ $Y2=0
r99 43 44 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.55
+ $Y2=0
r100 42 57 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.68 $Y=0 $X2=4.08
+ $Y2=0
r101 42 44 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.68 $Y=0 $X2=3.55
+ $Y2=0
r102 40 49 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.68
+ $Y2=0
r103 40 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.795
+ $Y2=0
r104 36 66 3.27398 $w=3.3e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.375 $Y=0.085
+ $X2=4.505 $Y2=0
r105 36 38 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.375 $Y=0.085
+ $X2=4.375 $Y2=0.38
r106 32 44 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r107 32 34 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.41
r108 28 63 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.655 $Y=0.085
+ $X2=2.655 $Y2=0
r109 28 30 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=2.655 $Y=0.085
+ $X2=2.655 $Y2=0.41
r110 27 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.795
+ $Y2=0
r111 26 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.655
+ $Y2=0
r112 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.56 $Y=0 $X2=1.89
+ $Y2=0
r113 22 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=0.085
+ $X2=1.795 $Y2=0
r114 22 24 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=1.795 $Y=0.085
+ $X2=1.795 $Y2=0.41
r115 18 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=0.085
+ $X2=0.855 $Y2=0
r116 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=0.085
+ $X2=0.855 $Y2=0.38
r117 5 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.235
+ $Y=0.235 $X2=4.375 $Y2=0.38
r118 4 34 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.235 $X2=3.515 $Y2=0.41
r119 3 30 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.235 $X2=2.655 $Y2=0.41
r120 2 24 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.235 $X2=1.795 $Y2=0.41
r121 1 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.715
+ $Y=0.235 $X2=0.855 $Y2=0.38
.ends

