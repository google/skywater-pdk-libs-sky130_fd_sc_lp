* File: sky130_fd_sc_lp__isobufsrc_1.pex.spice
* Created: Fri Aug 28 10:41:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_1%A 3 5 7 9 10
c25 10 0 6.58189e-20 $X=0.72 $Y=1.665
c26 3 0 2.76518e-19 $X=0.735 $Y=0.445
r27 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.51 $X2=0.64 $Y2=1.51
r28 10 15 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=0.72 $Y=1.587 $X2=0.64
+ $Y2=1.587
r29 9 15 14.1839 $w=3.23e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=1.587 $X2=0.64
+ $Y2=1.587
r30 5 14 38.9663 $w=3.64e-07 $l=2.18746e-07 $layer=POLY_cond $X=0.8 $Y=1.675
+ $X2=0.675 $Y2=1.51
r31 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.8 $Y=1.675 $X2=0.8
+ $Y2=2.045
r32 1 14 38.9663 $w=3.64e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.735 $Y=1.345
+ $X2=0.675 $Y2=1.51
r33 1 3 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=0.735 $Y=1.345 $X2=0.735
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_1%SLEEP 3 7 9 12 13
c34 7 0 6.58189e-20 $X=1.34 $Y=2.465
r35 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.51
+ $X2=1.25 $Y2=1.675
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.51
+ $X2=1.25 $Y2=1.345
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.51 $X2=1.25 $Y2=1.51
r38 9 13 4.70075 $w=3.78e-07 $l=1.55e-07 $layer=LI1_cond $X=1.225 $Y=1.665
+ $X2=1.225 $Y2=1.51
r39 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.34 $Y=2.465
+ $X2=1.34 $Y2=1.675
r40 3 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.34 $Y=0.655
+ $X2=1.34 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_1%A_79_47# 1 2 9 13 16 18 22 23 25 26 30
+ 33
c61 30 0 1.21421e-19 $X=1.79 $Y=1.35
r62 30 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.35
+ $X2=1.79 $Y2=1.515
r63 30 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.35
+ $X2=1.79 $Y2=1.185
r64 29 31 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=1.35
+ $X2=1.735 $Y2=1.515
r65 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.35 $X2=1.79 $Y2=1.35
r66 26 29 6.91466 $w=2.98e-07 $l=1.8e-07 $layer=LI1_cond $X=1.735 $Y=1.17
+ $X2=1.735 $Y2=1.35
r67 25 31 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.67 $Y=1.92
+ $X2=1.67 $Y2=1.515
r68 22 26 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.585 $Y=1.17 $X2=1.735
+ $Y2=1.17
r69 22 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.585 $Y=1.17
+ $X2=0.625 $Y2=1.17
r70 18 25 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.585 $Y=2.03
+ $X2=1.67 $Y2=1.92
r71 18 20 52.3838 $w=2.18e-07 $l=1e-06 $layer=LI1_cond $X=1.585 $Y=2.03
+ $X2=0.585 $Y2=2.03
r72 14 23 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.49 $Y=1.085
+ $X2=0.625 $Y2=1.17
r73 14 16 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.49 $Y=1.085
+ $X2=0.49 $Y2=0.45
r74 13 33 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.77 $Y=0.655
+ $X2=1.77 $Y2=1.185
r75 9 34 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.7 $Y=2.465 $X2=1.7
+ $Y2=1.515
r76 2 20 600 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=0.46
+ $Y=1.835 $X2=0.585 $Y2=2.03
r77 1 16 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.395
+ $Y=0.235 $X2=0.52 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_1%VPWR 1 6 8 10 17 18 21
r20 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r21 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.125 $Y2=3.33
r22 15 17 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=2.16 $Y2=3.33
r23 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r24 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=1.125 $Y2=3.33
r25 10 12 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r27 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.72
+ $Y2=3.33
r28 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r29 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=3.245
+ $X2=1.125 $Y2=3.33
r30 4 6 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=1.125 $Y=3.245
+ $X2=1.125 $Y2=2.42
r31 1 6 300 $w=1.7e-07 $l=6.9891e-07 $layer=licon1_PDIFF $count=2 $X=0.875
+ $Y=1.835 $X2=1.125 $Y2=2.42
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_1%X 1 2 7 9 11 15 16 17 18 19 20 29 32 40
c37 9 0 1.68039e-19 $X=1.555 $Y=0.42
c38 7 0 2.299e-19 $X=1.52 $Y=0.745
r39 38 40 0.738746 $w=3.88e-07 $l=2.5e-08 $layer=LI1_cond $X=2.12 $Y=2.01
+ $X2=2.12 $Y2=2.035
r40 29 32 0.443247 $w=2.58e-07 $l=1e-08 $layer=LI1_cond $X=2.185 $Y=0.915
+ $X2=2.185 $Y2=0.925
r41 20 47 3.98923 $w=3.88e-07 $l=1.35e-07 $layer=LI1_cond $X=2.12 $Y=2.775
+ $X2=2.12 $Y2=2.91
r42 19 20 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.12 $Y=2.405
+ $X2=2.12 $Y2=2.775
r43 18 38 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=2.12 $Y=1.98 $X2=2.12
+ $Y2=2.01
r44 18 52 6.15921 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=1.98
+ $X2=2.12 $Y2=1.815
r45 18 19 10.0469 $w=3.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.12 $Y=2.065
+ $X2=2.12 $Y2=2.405
r46 18 40 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=2.12 $Y=2.065
+ $X2=2.12 $Y2=2.035
r47 17 52 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=2.185 $Y=1.665
+ $X2=2.185 $Y2=1.815
r48 16 17 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.185 $Y=1.295
+ $X2=2.185 $Y2=1.665
r49 15 29 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=0.83
+ $X2=2.185 $Y2=0.915
r50 15 16 14.7601 $w=2.58e-07 $l=3.33e-07 $layer=LI1_cond $X=2.185 $Y=0.962
+ $X2=2.185 $Y2=1.295
r51 15 32 1.64002 $w=2.58e-07 $l=3.7e-08 $layer=LI1_cond $X=2.185 $Y=0.962
+ $X2=2.185 $Y2=0.925
r52 12 14 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.65 $Y=0.83 $X2=1.52
+ $Y2=0.83
r53 11 15 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.055 $Y=0.83
+ $X2=2.185 $Y2=0.83
r54 11 12 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.055 $Y=0.83
+ $X2=1.65 $Y2=0.83
r55 7 14 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=0.745 $X2=1.52
+ $Y2=0.83
r56 7 9 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=1.52 $Y=0.745
+ $X2=1.52 $Y2=0.42
r57 2 18 400 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=1.775
+ $Y=1.835 $X2=2.01 $Y2=1.98
r58 2 47 400 $w=1.7e-07 $l=1.1867e-06 $layer=licon1_PDIFF $count=1 $X=1.775
+ $Y=1.835 $X2=2.01 $Y2=2.91
r59 1 14 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.235 $X2=1.555 $Y2=0.83
r60 1 9 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.415
+ $Y=0.235 $X2=1.555 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__ISOBUFSRC_1%VGND 1 2 9 11 13 16 17 18 24 30
r34 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 27 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r36 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r37 24 29 4.50438 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=2.11
+ $Y2=0
r38 24 26 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=1.68
+ $Y2=0
r39 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r41 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r42 16 21 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.72
+ $Y2=0
r43 16 17 10.2049 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.007
+ $Y2=0
r44 15 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.68
+ $Y2=0
r45 15 17 10.2049 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.007
+ $Y2=0
r46 11 29 3.26179 $w=3.3e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.985 $Y=0.085
+ $X2=2.11 $Y2=0
r47 11 13 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.985 $Y=0.085
+ $X2=1.985 $Y2=0.45
r48 7 17 1.63918 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.007 $Y=0.085
+ $X2=1.007 $Y2=0
r49 7 9 7.99931 $w=4.23e-07 $l=2.95e-07 $layer=LI1_cond $X=1.007 $Y=0.085
+ $X2=1.007 $Y2=0.38
r50 2 13 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.235 $X2=1.985 $Y2=0.45
r51 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.81
+ $Y=0.235 $X2=0.95 $Y2=0.38
.ends

