* File: sky130_fd_sc_lp__xnor2_lp.pxi.spice
* Created: Wed Sep  2 10:40:24 2020
* 
x_PM_SKY130_FD_SC_LP__XNOR2_LP%A_82_66# N_A_82_66#_M1008_d N_A_82_66#_M1007_d
+ N_A_82_66#_M1009_g N_A_82_66#_M1000_g N_A_82_66#_c_63_n N_A_82_66#_c_69_n
+ N_A_82_66#_c_70_n N_A_82_66#_c_88_p N_A_82_66#_c_77_p N_A_82_66#_c_71_n
+ N_A_82_66#_c_64_n N_A_82_66#_c_73_n N_A_82_66#_c_65_n N_A_82_66#_c_66_n
+ PM_SKY130_FD_SC_LP__XNOR2_LP%A_82_66#
x_PM_SKY130_FD_SC_LP__XNOR2_LP%A N_A_M1002_g N_A_c_141_n N_A_M1004_g N_A_M1007_g
+ N_A_c_142_n N_A_M1005_g A N_A_c_143_n N_A_c_144_n
+ PM_SKY130_FD_SC_LP__XNOR2_LP%A
x_PM_SKY130_FD_SC_LP__XNOR2_LP%B N_B_M1006_g N_B_M1001_g N_B_c_194_n N_B_c_195_n
+ N_B_M1003_g N_B_M1008_g N_B_c_197_n B N_B_c_198_n N_B_c_199_n
+ PM_SKY130_FD_SC_LP__XNOR2_LP%B
x_PM_SKY130_FD_SC_LP__XNOR2_LP%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_M1003_d
+ N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_268_n
+ N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n VPWR N_VPWR_c_272_n
+ N_VPWR_c_263_n PM_SKY130_FD_SC_LP__XNOR2_LP%VPWR
x_PM_SKY130_FD_SC_LP__XNOR2_LP%Y N_Y_M1009_s N_Y_M1000_d N_Y_c_312_n N_Y_c_313_n
+ N_Y_c_320_n Y Y Y Y Y PM_SKY130_FD_SC_LP__XNOR2_LP%Y
x_PM_SKY130_FD_SC_LP__XNOR2_LP%A_112_92# N_A_112_92#_M1009_d N_A_112_92#_M1001_d
+ N_A_112_92#_c_345_n N_A_112_92#_c_346_n N_A_112_92#_c_347_n
+ N_A_112_92#_c_348_n PM_SKY130_FD_SC_LP__XNOR2_LP%A_112_92#
x_PM_SKY130_FD_SC_LP__XNOR2_LP%VGND N_VGND_M1001_s N_VGND_M1004_d N_VGND_c_374_n
+ N_VGND_c_375_n N_VGND_c_376_n VGND N_VGND_c_377_n N_VGND_c_378_n
+ N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n PM_SKY130_FD_SC_LP__XNOR2_LP%VGND
cc_1 VNB N_A_82_66#_M1009_g 0.0521091f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.67
cc_2 VNB N_A_82_66#_c_63_n 0.00513937f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.63
cc_3 VNB N_A_82_66#_c_64_n 0.0288692f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=2.02
cc_4 VNB N_A_82_66#_c_65_n 0.0280857f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.835
cc_5 VNB N_A_82_66#_c_66_n 0.0258312f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.63
cc_6 VNB N_A_c_141_n 0.0135832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_c_142_n 0.0130302f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.595
cc_8 VNB N_A_c_143_n 6.97565e-19 $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=2.02
cc_9 VNB N_A_c_144_n 0.0880156f $X=-0.19 $Y=-0.245 $X2=2.395 $Y2=2.105
cc_10 VNB N_B_M1006_g 0.0250869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_M1001_g 0.0314904f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.67
cc_12 VNB N_B_c_194_n 0.107095f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.67
cc_13 VNB N_B_c_195_n 0.011606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_M1008_g 0.0592368f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.63
cc_15 VNB N_B_c_197_n 0.0211529f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=2.02
cc_16 VNB N_B_c_198_n 0.0193663f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.24
cc_17 VNB N_B_c_199_n 0.00413684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_263_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB Y 0.0229391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB Y 0.0386738f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.24
cc_21 VNB N_A_112_92#_c_345_n 0.0131992f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.67
cc_22 VNB N_A_112_92#_c_346_n 0.0218816f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.795
cc_23 VNB N_A_112_92#_c_347_n 0.00429736f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.595
cc_24 VNB N_A_112_92#_c_348_n 0.00396962f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.63
cc_25 VNB N_VGND_c_374_n 0.0139622f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.67
cc_26 VNB N_VGND_c_375_n 0.0186281f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.795
cc_27 VNB N_VGND_c_376_n 0.0104951f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.63
cc_28 VNB N_VGND_c_377_n 0.0325812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_378_n 0.0317278f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.24
cc_30 VNB N_VGND_c_379_n 0.209859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_380_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=1.065
cc_32 VNB N_VGND_c_381_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=3.092 $Y2=0.835
cc_33 VPB N_A_82_66#_M1000_g 0.0380902f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=2.595
cc_34 VPB N_A_82_66#_c_63_n 0.00391534f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=1.63
cc_35 VPB N_A_82_66#_c_69_n 0.00207192f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=2.02
cc_36 VPB N_A_82_66#_c_70_n 0.00888168f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=2.105
cc_37 VPB N_A_82_66#_c_71_n 0.01323f $X=-0.19 $Y=1.655 $X2=3.1 $Y2=2.105
cc_38 VPB N_A_82_66#_c_64_n 0.01738f $X=-0.19 $Y=1.655 $X2=3.185 $Y2=2.02
cc_39 VPB N_A_82_66#_c_73_n 0.00572113f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.105
cc_40 VPB N_A_82_66#_c_66_n 0.0174328f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.63
cc_41 VPB N_A_M1002_g 0.038513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_M1007_g 0.038684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_c_143_n 0.00272477f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=2.02
cc_44 VPB N_A_c_144_n 0.00529095f $X=-0.19 $Y=1.655 $X2=2.395 $Y2=2.105
cc_45 VPB N_B_M1006_g 0.0390333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_B_M1003_g 0.0347017f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=2.595
cc_47 VPB N_B_c_198_n 0.0146948f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.24
cc_48 VPB N_B_c_199_n 0.00235259f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_264_n 0.0320215f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=2.595
cc_50 VPB N_VPWR_c_265_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.705 $Y2=1.63
cc_51 VPB N_VPWR_c_266_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=1.63
cc_52 VPB N_VPWR_c_267_n 0.0306765f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=1.795
cc_53 VPB N_VPWR_c_268_n 0.0121672f $X=-0.19 $Y=1.655 $X2=1.525 $Y2=2.105
cc_54 VPB N_VPWR_c_269_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.19
cc_55 VPB N_VPWR_c_270_n 0.0336396f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.24
cc_56 VPB N_VPWR_c_271_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_272_n 0.0180468f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.63
cc_58 VPB N_VPWR_c_263_n 0.0530199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_Y_c_312_n 0.00665348f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.465
cc_60 VPB N_Y_c_313_n 0.017193f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.67
cc_61 VPB Y 0.0171868f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.24
cc_62 N_A_82_66#_c_69_n N_A_M1002_g 0.00492462f $X=1.44 $Y=2.02 $X2=0 $Y2=0
cc_63 N_A_82_66#_c_70_n N_A_M1002_g 0.0287875f $X=2.395 $Y=2.105 $X2=0 $Y2=0
cc_64 N_A_82_66#_c_77_p N_A_M1002_g 8.96718e-19 $X=2.56 $Y=2.24 $X2=0 $Y2=0
cc_65 N_A_82_66#_c_70_n N_A_M1007_g 0.019614f $X=2.395 $Y=2.105 $X2=0 $Y2=0
cc_66 N_A_82_66#_c_77_p N_A_M1007_g 0.0186751f $X=2.56 $Y=2.24 $X2=0 $Y2=0
cc_67 N_A_82_66#_c_73_n N_A_M1007_g 0.00247044f $X=2.56 $Y=2.105 $X2=0 $Y2=0
cc_68 N_A_82_66#_c_65_n N_A_c_142_n 0.00135161f $X=3.08 $Y=0.835 $X2=0 $Y2=0
cc_69 N_A_82_66#_c_63_n N_A_c_143_n 0.0128152f $X=1.355 $Y=1.63 $X2=0 $Y2=0
cc_70 N_A_82_66#_c_70_n N_A_c_143_n 0.0198621f $X=2.395 $Y=2.105 $X2=0 $Y2=0
cc_71 N_A_82_66#_c_63_n N_A_c_144_n 0.00428614f $X=1.355 $Y=1.63 $X2=0 $Y2=0
cc_72 N_A_82_66#_c_70_n N_A_c_144_n 0.00139135f $X=2.395 $Y=2.105 $X2=0 $Y2=0
cc_73 N_A_82_66#_c_63_n N_B_M1006_g 0.0262684f $X=1.355 $Y=1.63 $X2=0 $Y2=0
cc_74 N_A_82_66#_c_69_n N_B_M1006_g 0.00573536f $X=1.44 $Y=2.02 $X2=0 $Y2=0
cc_75 N_A_82_66#_c_88_p N_B_M1006_g 0.00720587f $X=1.525 $Y=2.105 $X2=0 $Y2=0
cc_76 N_A_82_66#_c_66_n N_B_M1006_g 0.048292f $X=0.745 $Y=1.63 $X2=0 $Y2=0
cc_77 N_A_82_66#_c_77_p N_B_M1003_g 0.0235494f $X=2.56 $Y=2.24 $X2=0 $Y2=0
cc_78 N_A_82_66#_c_71_n N_B_M1003_g 0.0201967f $X=3.1 $Y=2.105 $X2=0 $Y2=0
cc_79 N_A_82_66#_c_64_n N_B_M1003_g 0.00664445f $X=3.185 $Y=2.02 $X2=0 $Y2=0
cc_80 N_A_82_66#_c_73_n N_B_M1003_g 0.00163487f $X=2.56 $Y=2.105 $X2=0 $Y2=0
cc_81 N_A_82_66#_c_64_n N_B_M1008_g 0.0153664f $X=3.185 $Y=2.02 $X2=0 $Y2=0
cc_82 N_A_82_66#_c_65_n N_B_M1008_g 0.0113826f $X=3.08 $Y=0.835 $X2=0 $Y2=0
cc_83 N_A_82_66#_M1009_g N_B_c_197_n 0.00684931f $X=0.485 $Y=0.67 $X2=0 $Y2=0
cc_84 N_A_82_66#_c_63_n N_B_c_197_n 9.33926e-19 $X=1.355 $Y=1.63 $X2=0 $Y2=0
cc_85 N_A_82_66#_c_71_n N_B_c_198_n 3.71629e-19 $X=3.1 $Y=2.105 $X2=0 $Y2=0
cc_86 N_A_82_66#_c_64_n N_B_c_198_n 0.00773251f $X=3.185 $Y=2.02 $X2=0 $Y2=0
cc_87 N_A_82_66#_c_73_n N_B_c_198_n 0.00162266f $X=2.56 $Y=2.105 $X2=0 $Y2=0
cc_88 N_A_82_66#_c_65_n N_B_c_198_n 6.59447e-19 $X=3.08 $Y=0.835 $X2=0 $Y2=0
cc_89 N_A_82_66#_c_71_n N_B_c_199_n 0.0132692f $X=3.1 $Y=2.105 $X2=0 $Y2=0
cc_90 N_A_82_66#_c_64_n N_B_c_199_n 0.0240488f $X=3.185 $Y=2.02 $X2=0 $Y2=0
cc_91 N_A_82_66#_c_73_n N_B_c_199_n 0.0164798f $X=2.56 $Y=2.105 $X2=0 $Y2=0
cc_92 N_A_82_66#_c_70_n N_VPWR_M1002_d 0.00180746f $X=2.395 $Y=2.105 $X2=0 $Y2=0
cc_93 N_A_82_66#_c_71_n N_VPWR_M1003_d 0.00291845f $X=3.1 $Y=2.105 $X2=0 $Y2=0
cc_94 N_A_82_66#_M1000_g N_VPWR_c_264_n 0.0208226f $X=0.745 $Y=2.595 $X2=0 $Y2=0
cc_95 N_A_82_66#_c_70_n N_VPWR_c_265_n 0.0163515f $X=2.395 $Y=2.105 $X2=0 $Y2=0
cc_96 N_A_82_66#_c_77_p N_VPWR_c_265_n 0.045794f $X=2.56 $Y=2.24 $X2=0 $Y2=0
cc_97 N_A_82_66#_c_77_p N_VPWR_c_267_n 0.045794f $X=2.56 $Y=2.24 $X2=0 $Y2=0
cc_98 N_A_82_66#_c_71_n N_VPWR_c_267_n 0.0223246f $X=3.1 $Y=2.105 $X2=0 $Y2=0
cc_99 N_A_82_66#_M1000_g N_VPWR_c_270_n 0.00840199f $X=0.745 $Y=2.595 $X2=0
+ $Y2=0
cc_100 N_A_82_66#_c_77_p N_VPWR_c_272_n 0.0177952f $X=2.56 $Y=2.24 $X2=0 $Y2=0
cc_101 N_A_82_66#_M1007_d N_VPWR_c_263_n 0.00223819f $X=2.42 $Y=2.095 $X2=0
+ $Y2=0
cc_102 N_A_82_66#_M1000_g N_VPWR_c_263_n 0.0136033f $X=0.745 $Y=2.595 $X2=0
+ $Y2=0
cc_103 N_A_82_66#_c_77_p N_VPWR_c_263_n 0.0123247f $X=2.56 $Y=2.24 $X2=0 $Y2=0
cc_104 N_A_82_66#_M1000_g N_Y_c_312_n 0.0218581f $X=0.745 $Y=2.595 $X2=0 $Y2=0
cc_105 N_A_82_66#_c_63_n N_Y_c_312_n 0.0486713f $X=1.355 $Y=1.63 $X2=0 $Y2=0
cc_106 N_A_82_66#_c_69_n N_Y_c_312_n 0.0032409f $X=1.44 $Y=2.02 $X2=0 $Y2=0
cc_107 N_A_82_66#_c_88_p N_Y_c_312_n 0.0101017f $X=1.525 $Y=2.105 $X2=0 $Y2=0
cc_108 N_A_82_66#_c_66_n N_Y_c_312_n 0.00719794f $X=0.745 $Y=1.63 $X2=0 $Y2=0
cc_109 N_A_82_66#_M1000_g N_Y_c_320_n 0.0243371f $X=0.745 $Y=2.595 $X2=0 $Y2=0
cc_110 N_A_82_66#_c_88_p N_Y_c_320_n 0.00339424f $X=1.525 $Y=2.105 $X2=0 $Y2=0
cc_111 N_A_82_66#_M1009_g Y 0.0079188f $X=0.485 $Y=0.67 $X2=0 $Y2=0
cc_112 N_A_82_66#_M1009_g Y 0.0256528f $X=0.485 $Y=0.67 $X2=0 $Y2=0
cc_113 N_A_82_66#_M1000_g Y 0.0061332f $X=0.745 $Y=2.595 $X2=0 $Y2=0
cc_114 N_A_82_66#_c_63_n Y 0.0252802f $X=1.355 $Y=1.63 $X2=0 $Y2=0
cc_115 N_A_82_66#_c_70_n A_280_419# 0.00217487f $X=2.395 $Y=2.105 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A_82_66#_c_88_p A_280_419# 0.00306752f $X=1.525 $Y=2.105 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_82_66#_M1009_g N_A_112_92#_c_345_n 0.0065332f $X=0.485 $Y=0.67 $X2=0
+ $Y2=0
cc_118 N_A_82_66#_c_63_n N_A_112_92#_c_346_n 0.0490043f $X=1.355 $Y=1.63 $X2=0
+ $Y2=0
cc_119 N_A_82_66#_M1009_g N_A_112_92#_c_347_n 0.00234871f $X=0.485 $Y=0.67 $X2=0
+ $Y2=0
cc_120 N_A_82_66#_c_63_n N_A_112_92#_c_347_n 0.0201951f $X=1.355 $Y=1.63 $X2=0
+ $Y2=0
cc_121 N_A_82_66#_c_66_n N_A_112_92#_c_347_n 0.00675115f $X=0.745 $Y=1.63 $X2=0
+ $Y2=0
cc_122 N_A_82_66#_M1009_g N_VGND_c_374_n 0.00366022f $X=0.485 $Y=0.67 $X2=0
+ $Y2=0
cc_123 N_A_82_66#_c_65_n N_VGND_c_376_n 0.00708585f $X=3.08 $Y=0.835 $X2=0 $Y2=0
cc_124 N_A_82_66#_M1009_g N_VGND_c_377_n 0.00491683f $X=0.485 $Y=0.67 $X2=0
+ $Y2=0
cc_125 N_A_82_66#_c_65_n N_VGND_c_378_n 0.00744886f $X=3.08 $Y=0.835 $X2=0 $Y2=0
cc_126 N_A_82_66#_M1009_g N_VGND_c_379_n 0.00517496f $X=0.485 $Y=0.67 $X2=0
+ $Y2=0
cc_127 N_A_82_66#_c_65_n N_VGND_c_379_n 0.0107293f $X=3.08 $Y=0.835 $X2=0 $Y2=0
cc_128 N_A_c_143_n N_B_M1006_g 7.98427e-19 $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_144_n N_B_M1006_g 0.102585f $X=2.295 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_141_n N_B_M1001_g 0.0118161f $X=2.045 $Y=1.12 $X2=0 $Y2=0
cc_131 N_A_c_141_n N_B_c_194_n 0.00894529f $X=2.045 $Y=1.12 $X2=0 $Y2=0
cc_132 N_A_c_142_n N_B_c_194_n 0.00907339f $X=2.475 $Y=1.12 $X2=0 $Y2=0
cc_133 N_A_M1007_g N_B_M1003_g 0.031542f $X=2.295 $Y=2.595 $X2=0 $Y2=0
cc_134 N_A_c_142_n N_B_M1008_g 0.0408321f $X=2.475 $Y=1.12 $X2=0 $Y2=0
cc_135 N_A_c_143_n N_B_M1008_g 0.00143915f $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_c_144_n N_B_M1008_g 0.00753084f $X=2.295 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_c_144_n N_B_c_197_n 0.00977923f $X=2.295 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_143_n N_B_c_198_n 2.53686e-19 $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_144_n N_B_c_198_n 0.0189629f $X=2.295 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_143_n N_B_c_199_n 0.0207474f $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_144_n N_B_c_199_n 0.00435693f $X=2.295 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_M1002_g N_VPWR_c_265_n 0.0198958f $X=1.765 $Y=2.595 $X2=0 $Y2=0
cc_143 N_A_M1007_g N_VPWR_c_265_n 0.0178867f $X=2.295 $Y=2.595 $X2=0 $Y2=0
cc_144 N_A_M1007_g N_VPWR_c_267_n 0.00120686f $X=2.295 $Y=2.595 $X2=0 $Y2=0
cc_145 N_A_M1002_g N_VPWR_c_270_n 0.008763f $X=1.765 $Y=2.595 $X2=0 $Y2=0
cc_146 N_A_M1007_g N_VPWR_c_272_n 0.00840199f $X=2.295 $Y=2.595 $X2=0 $Y2=0
cc_147 N_A_M1002_g N_VPWR_c_263_n 0.0144563f $X=1.765 $Y=2.595 $X2=0 $Y2=0
cc_148 N_A_M1007_g N_VPWR_c_263_n 0.0136033f $X=2.295 $Y=2.595 $X2=0 $Y2=0
cc_149 N_A_M1002_g N_Y_c_320_n 0.00381029f $X=1.765 $Y=2.595 $X2=0 $Y2=0
cc_150 N_A_c_143_n N_A_112_92#_c_346_n 0.0030491f $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_144_n N_A_112_92#_c_346_n 0.0213858f $X=2.295 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_141_n N_A_112_92#_c_348_n 0.00539947f $X=2.045 $Y=1.12 $X2=0 $Y2=0
cc_153 N_A_c_141_n N_VGND_c_374_n 5.6275e-19 $X=2.045 $Y=1.12 $X2=0 $Y2=0
cc_154 N_A_c_141_n N_VGND_c_376_n 0.0102118f $X=2.045 $Y=1.12 $X2=0 $Y2=0
cc_155 N_A_c_142_n N_VGND_c_376_n 0.00344526f $X=2.475 $Y=1.12 $X2=0 $Y2=0
cc_156 N_A_c_143_n N_VGND_c_376_n 0.0207027f $X=2.18 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_144_n N_VGND_c_376_n 0.00314735f $X=2.295 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_141_n N_VGND_c_379_n 7.97988e-19 $X=2.045 $Y=1.12 $X2=0 $Y2=0
cc_159 N_A_c_142_n N_VGND_c_379_n 9.49986e-19 $X=2.475 $Y=1.12 $X2=0 $Y2=0
cc_160 N_B_M1006_g N_VPWR_c_264_n 0.00121833f $X=1.275 $Y=2.595 $X2=0 $Y2=0
cc_161 N_B_M1006_g N_VPWR_c_265_n 0.00403993f $X=1.275 $Y=2.595 $X2=0 $Y2=0
cc_162 N_B_M1003_g N_VPWR_c_265_n 0.00120686f $X=2.825 $Y=2.595 $X2=0 $Y2=0
cc_163 N_B_M1003_g N_VPWR_c_267_n 0.0191563f $X=2.825 $Y=2.595 $X2=0 $Y2=0
cc_164 N_B_M1006_g N_VPWR_c_270_n 0.00939541f $X=1.275 $Y=2.595 $X2=0 $Y2=0
cc_165 N_B_M1003_g N_VPWR_c_272_n 0.00840199f $X=2.825 $Y=2.595 $X2=0 $Y2=0
cc_166 N_B_M1006_g N_VPWR_c_263_n 0.0161521f $X=1.275 $Y=2.595 $X2=0 $Y2=0
cc_167 N_B_M1003_g N_VPWR_c_263_n 0.0136033f $X=2.825 $Y=2.595 $X2=0 $Y2=0
cc_168 N_B_M1006_g N_Y_c_312_n 0.00455016f $X=1.275 $Y=2.595 $X2=0 $Y2=0
cc_169 N_B_M1006_g N_Y_c_320_n 0.0212894f $X=1.275 $Y=2.595 $X2=0 $Y2=0
cc_170 N_B_M1001_g N_A_112_92#_c_345_n 0.00531518f $X=1.455 $Y=0.835 $X2=0 $Y2=0
cc_171 N_B_M1006_g N_A_112_92#_c_346_n 0.00424692f $X=1.275 $Y=2.595 $X2=0 $Y2=0
cc_172 N_B_M1001_g N_A_112_92#_c_346_n 0.00595264f $X=1.455 $Y=0.835 $X2=0 $Y2=0
cc_173 N_B_c_197_n N_A_112_92#_c_346_n 0.0145114f $X=1.455 $Y=1.195 $X2=0 $Y2=0
cc_174 N_B_M1001_g N_A_112_92#_c_348_n 0.00467559f $X=1.455 $Y=0.835 $X2=0 $Y2=0
cc_175 N_B_c_194_n N_A_112_92#_c_348_n 0.00423145f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_176 N_B_M1001_g N_VGND_c_374_n 0.0239291f $X=1.455 $Y=0.835 $X2=0 $Y2=0
cc_177 N_B_c_195_n N_VGND_c_374_n 0.00763335f $X=1.53 $Y=0.18 $X2=0 $Y2=0
cc_178 N_B_c_197_n N_VGND_c_374_n 0.0015874f $X=1.455 $Y=1.195 $X2=0 $Y2=0
cc_179 N_B_c_195_n N_VGND_c_375_n 0.0223737f $X=1.53 $Y=0.18 $X2=0 $Y2=0
cc_180 N_B_M1001_g N_VGND_c_376_n 0.00631882f $X=1.455 $Y=0.835 $X2=0 $Y2=0
cc_181 N_B_c_194_n N_VGND_c_376_n 0.0211809f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_182 N_B_M1008_g N_VGND_c_376_n 0.00742201f $X=2.865 $Y=0.835 $X2=0 $Y2=0
cc_183 N_B_c_194_n N_VGND_c_378_n 0.0215943f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_184 N_B_c_194_n N_VGND_c_379_n 0.0529798f $X=2.79 $Y=0.18 $X2=0 $Y2=0
cc_185 N_B_c_195_n N_VGND_c_379_n 0.00749832f $X=1.53 $Y=0.18 $X2=0 $Y2=0
cc_186 N_VPWR_c_263_n N_Y_M1000_d 0.00223819f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_187 N_VPWR_M1000_s N_Y_c_312_n 0.0024817f $X=0.335 $Y=2.095 $X2=0 $Y2=0
cc_188 N_VPWR_c_264_n N_Y_c_312_n 0.017885f $X=0.48 $Y=2.49 $X2=0 $Y2=0
cc_189 N_VPWR_M1000_s N_Y_c_313_n 2.821e-19 $X=0.335 $Y=2.095 $X2=0 $Y2=0
cc_190 N_VPWR_c_264_n N_Y_c_313_n 0.00343641f $X=0.48 $Y=2.49 $X2=0 $Y2=0
cc_191 N_VPWR_c_264_n N_Y_c_320_n 0.0487591f $X=0.48 $Y=2.49 $X2=0 $Y2=0
cc_192 N_VPWR_c_270_n N_Y_c_320_n 0.0177952f $X=1.865 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_263_n N_Y_c_320_n 0.0123247f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_c_263_n A_280_419# 0.010279f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_195 Y N_A_112_92#_c_345_n 0.0179429f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_196 Y N_A_112_92#_c_345_n 0.0126887f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_197 Y N_A_112_92#_c_347_n 0.0109342f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_198 Y N_VGND_c_377_n 0.0105942f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_199 Y N_VGND_c_379_n 0.0113723f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_200 N_A_112_92#_c_345_n N_VGND_c_374_n 0.0348134f $X=0.7 $Y=0.67 $X2=0 $Y2=0
cc_201 N_A_112_92#_c_346_n N_VGND_c_374_n 0.0234162f $X=1.585 $Y=1.2 $X2=0 $Y2=0
cc_202 N_A_112_92#_c_348_n N_VGND_c_374_n 0.0125556f $X=1.75 $Y=0.835 $X2=0
+ $Y2=0
cc_203 N_A_112_92#_c_348_n N_VGND_c_375_n 0.00534397f $X=1.75 $Y=0.835 $X2=0
+ $Y2=0
cc_204 N_A_112_92#_c_348_n N_VGND_c_376_n 0.0247809f $X=1.75 $Y=0.835 $X2=0
+ $Y2=0
cc_205 N_A_112_92#_c_345_n N_VGND_c_377_n 0.00810947f $X=0.7 $Y=0.67 $X2=0 $Y2=0
cc_206 N_A_112_92#_c_345_n N_VGND_c_379_n 0.00864691f $X=0.7 $Y=0.67 $X2=0 $Y2=0
cc_207 N_A_112_92#_c_348_n N_VGND_c_379_n 0.00671416f $X=1.75 $Y=0.835 $X2=0
+ $Y2=0
