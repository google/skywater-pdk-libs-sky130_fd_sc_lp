* File: sky130_fd_sc_lp__dlrtp_lp.pxi.spice
* Created: Fri Aug 28 10:27:37 2020
* 
x_PM_SKY130_FD_SC_LP__DLRTP_LP%GATE N_GATE_M1010_g N_GATE_M1022_g N_GATE_M1001_g
+ N_GATE_M1018_g GATE GATE GATE N_GATE_c_169_n PM_SKY130_FD_SC_LP__DLRTP_LP%GATE
x_PM_SKY130_FD_SC_LP__DLRTP_LP%A_186_57# N_A_186_57#_M1001_d N_A_186_57#_M1018_d
+ N_A_186_57#_M1004_g N_A_186_57#_c_197_n N_A_186_57#_M1006_g
+ N_A_186_57#_c_198_n N_A_186_57#_M1002_g N_A_186_57#_M1005_g
+ N_A_186_57#_c_199_n N_A_186_57#_M1017_g N_A_186_57#_c_201_n
+ N_A_186_57#_c_202_n N_A_186_57#_M1028_g N_A_186_57#_c_203_n
+ N_A_186_57#_c_217_n N_A_186_57#_c_204_n N_A_186_57#_c_237_p
+ N_A_186_57#_c_205_n N_A_186_57#_c_206_n N_A_186_57#_c_219_n
+ N_A_186_57#_c_220_n N_A_186_57#_c_207_n N_A_186_57#_c_208_n
+ N_A_186_57#_c_209_n N_A_186_57#_c_210_n N_A_186_57#_c_211_n
+ N_A_186_57#_c_212_n N_A_186_57#_c_213_n PM_SKY130_FD_SC_LP__DLRTP_LP%A_186_57#
x_PM_SKY130_FD_SC_LP__DLRTP_LP%D N_D_M1019_g N_D_c_332_n N_D_M1008_g N_D_M1020_g
+ N_D_c_333_n N_D_M1011_g D N_D_c_330_n N_D_c_331_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP%D
x_PM_SKY130_FD_SC_LP__DLRTP_LP%A_294_547# N_A_294_547#_M1006_s
+ N_A_294_547#_M1004_s N_A_294_547#_c_374_n N_A_294_547#_M1027_g
+ N_A_294_547#_c_370_n N_A_294_547#_c_371_n N_A_294_547#_M1026_g
+ N_A_294_547#_c_373_n N_A_294_547#_c_379_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP%A_294_547#
x_PM_SKY130_FD_SC_LP__DLRTP_LP%A_638_73# N_A_638_73#_M1020_d N_A_638_73#_M1011_d
+ N_A_638_73#_M1014_g N_A_638_73#_M1000_g N_A_638_73#_c_437_n
+ N_A_638_73#_c_444_n N_A_638_73#_c_438_n N_A_638_73#_c_445_n
+ N_A_638_73#_c_439_n N_A_638_73#_c_440_n N_A_638_73#_c_448_n
+ N_A_638_73#_c_449_n N_A_638_73#_c_441_n N_A_638_73#_c_442_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP%A_638_73#
x_PM_SKY130_FD_SC_LP__DLRTP_LP%A_1208_75# N_A_1208_75#_M1015_s
+ N_A_1208_75#_M1013_d N_A_1208_75#_c_523_n N_A_1208_75#_M1029_g
+ N_A_1208_75#_c_524_n N_A_1208_75#_c_525_n N_A_1208_75#_M1009_g
+ N_A_1208_75#_c_527_n N_A_1208_75#_c_528_n N_A_1208_75#_M1016_g
+ N_A_1208_75#_c_529_n N_A_1208_75#_M1007_g N_A_1208_75#_c_541_n
+ N_A_1208_75#_M1023_g N_A_1208_75#_c_530_n N_A_1208_75#_c_531_n
+ N_A_1208_75#_M1024_g N_A_1208_75#_c_533_n N_A_1208_75#_c_534_n
+ N_A_1208_75#_c_560_p N_A_1208_75#_c_535_n N_A_1208_75#_c_544_n
+ N_A_1208_75#_c_536_n N_A_1208_75#_c_537_n N_A_1208_75#_c_546_n
+ N_A_1208_75#_c_538_n N_A_1208_75#_c_539_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP%A_1208_75#
x_PM_SKY130_FD_SC_LP__DLRTP_LP%A_887_343# N_A_887_343#_M1028_d
+ N_A_887_343#_M1017_d N_A_887_343#_M1025_g N_A_887_343#_M1015_g
+ N_A_887_343#_M1003_g N_A_887_343#_c_648_n N_A_887_343#_c_649_n
+ N_A_887_343#_c_650_n N_A_887_343#_c_651_n N_A_887_343#_c_652_n
+ N_A_887_343#_c_653_n N_A_887_343#_c_654_n N_A_887_343#_c_655_n
+ N_A_887_343#_c_656_n N_A_887_343#_c_657_n N_A_887_343#_c_658_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP%A_887_343#
x_PM_SKY130_FD_SC_LP__DLRTP_LP%RESET_B N_RESET_B_M1021_g N_RESET_B_M1012_g
+ N_RESET_B_M1013_g RESET_B N_RESET_B_c_766_n N_RESET_B_c_767_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP%RESET_B
x_PM_SKY130_FD_SC_LP__DLRTP_LP%VPWR N_VPWR_M1022_s N_VPWR_M1005_d N_VPWR_M1000_d
+ N_VPWR_M1025_d N_VPWR_M1023_s N_VPWR_c_811_n N_VPWR_c_812_n N_VPWR_c_813_n
+ N_VPWR_c_814_n N_VPWR_c_815_n N_VPWR_c_816_n N_VPWR_c_817_n N_VPWR_c_818_n
+ VPWR N_VPWR_c_819_n N_VPWR_c_820_n N_VPWR_c_821_n N_VPWR_c_822_n
+ N_VPWR_c_810_n N_VPWR_c_824_n N_VPWR_c_825_n N_VPWR_c_826_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DLRTP_LP%A_800_343# N_A_800_343#_M1017_s
+ N_A_800_343#_M1000_s N_A_800_343#_c_904_n N_A_800_343#_c_905_n
+ N_A_800_343#_c_906_n N_A_800_343#_c_907_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP%A_800_343#
x_PM_SKY130_FD_SC_LP__DLRTP_LP%A_996_343# N_A_996_343#_M1027_d
+ N_A_996_343#_M1009_d N_A_996_343#_c_928_n N_A_996_343#_c_929_n
+ N_A_996_343#_c_930_n PM_SKY130_FD_SC_LP__DLRTP_LP%A_996_343#
x_PM_SKY130_FD_SC_LP__DLRTP_LP%A_1420_367# N_A_1420_367#_M1025_s
+ N_A_1420_367#_M1003_d N_A_1420_367#_c_953_n N_A_1420_367#_c_954_n
+ N_A_1420_367#_c_960_n N_A_1420_367#_c_955_n N_A_1420_367#_c_956_n
+ N_A_1420_367#_c_957_n PM_SKY130_FD_SC_LP__DLRTP_LP%A_1420_367#
x_PM_SKY130_FD_SC_LP__DLRTP_LP%Q N_Q_M1007_d N_Q_M1024_d Q Q Q Q Q Q Q
+ N_Q_c_998_n PM_SKY130_FD_SC_LP__DLRTP_LP%Q
x_PM_SKY130_FD_SC_LP__DLRTP_LP%VGND N_VGND_M1010_s N_VGND_M1002_d N_VGND_M1014_d
+ N_VGND_M1021_d N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n
+ N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n VGND N_VGND_c_1023_n
+ N_VGND_c_1024_n N_VGND_c_1025_n N_VGND_c_1026_n N_VGND_c_1027_n
+ N_VGND_c_1028_n PM_SKY130_FD_SC_LP__DLRTP_LP%VGND
x_PM_SKY130_FD_SC_LP__DLRTP_LP%A_862_101# N_A_862_101#_M1028_s
+ N_A_862_101#_M1029_d N_A_862_101#_c_1110_n N_A_862_101#_c_1111_n
+ N_A_862_101#_c_1112_n N_A_862_101#_c_1113_n N_A_862_101#_c_1114_n
+ N_A_862_101#_c_1115_n N_A_862_101#_c_1116_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP%A_862_101#
cc_1 VNB N_GATE_M1010_g 0.0484835f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_2 VNB N_GATE_M1001_g 0.0383858f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_3 VNB GATE 0.0268452f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_GATE_c_169_n 0.0519144f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.345
cc_5 VNB N_A_186_57#_c_197_n 0.0178318f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_6 VNB N_A_186_57#_c_198_n 0.0159255f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.67
cc_7 VNB N_A_186_57#_c_199_n 0.0399066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_186_57#_M1017_g 0.023327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_186_57#_c_201_n 0.0262709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_186_57#_c_202_n 0.01796f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.345
cc_11 VNB N_A_186_57#_c_203_n 0.00634987f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.295
cc_12 VNB N_A_186_57#_c_204_n 0.0171128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_186_57#_c_205_n 4.07275e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_186_57#_c_206_n 0.0806715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_186_57#_c_207_n 0.00345107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_186_57#_c_208_n 0.00124242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_186_57#_c_209_n 0.00384978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_186_57#_c_210_n 0.0121953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_186_57#_c_211_n 0.0199836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_186_57#_c_212_n 0.00100562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_186_57#_c_213_n 0.0375205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_D_M1019_g 0.0248756f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_23 VNB N_D_M1020_g 0.0308305f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.495
cc_24 VNB N_D_c_330_n 0.00463365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_D_c_331_n 0.0598574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_294_547#_c_370_n 0.00814792f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.85
cc_27 VNB N_A_294_547#_c_371_n 0.00657817f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.67
cc_28 VNB N_A_294_547#_M1026_g 0.0377396f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_29 VNB N_A_294_547#_c_373_n 0.0122148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_638_73#_M1014_g 0.0374641f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.18
cc_31 VNB N_A_638_73#_M1000_g 0.00318212f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.67
cc_32 VNB N_A_638_73#_c_437_n 0.0273164f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_33 VNB N_A_638_73#_c_438_n 0.0161059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_638_73#_c_439_n 0.00462897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_638_73#_c_440_n 0.00374693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_638_73#_c_441_n 0.0162908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_638_73#_c_442_n 0.0109834f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.345
cc_38 VNB N_A_1208_75#_c_523_n 0.0182329f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.67
cc_39 VNB N_A_1208_75#_c_524_n 0.00933855f $X=-0.19 $Y=-0.245 $X2=0.855
+ $Y2=0.495
cc_40 VNB N_A_1208_75#_c_525_n 0.00887484f $X=-0.19 $Y=-0.245 $X2=0.855
+ $Y2=0.495
cc_41 VNB N_A_1208_75#_M1009_g 0.0348179f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.67
cc_42 VNB N_A_1208_75#_c_527_n 0.00961044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1208_75#_c_528_n 0.0192913f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_44 VNB N_A_1208_75#_c_529_n 0.0190533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1208_75#_c_530_n 0.0310303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1208_75#_c_531_n 0.0509022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1208_75#_M1024_g 0.0202105f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.345
cc_48 VNB N_A_1208_75#_c_533_n 0.00717486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1208_75#_c_534_n 0.0346068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1208_75#_c_535_n 0.0183284f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.665
cc_51 VNB N_A_1208_75#_c_536_n 0.00241369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1208_75#_c_537_n 0.0468189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1208_75#_c_538_n 0.0081523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1208_75#_c_539_n 0.00101923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_887_343#_M1025_g 0.0112658f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.18
cc_56 VNB N_A_887_343#_M1003_g 0.00173276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_887_343#_c_648_n 9.85018e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_887_343#_c_649_n 0.00594192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_887_343#_c_650_n 0.0387702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_887_343#_c_651_n 0.00993991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_887_343#_c_652_n 0.0039598f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.345
cc_62 VNB N_A_887_343#_c_653_n 0.0177693f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.345
cc_63 VNB N_A_887_343#_c_654_n 0.00124125f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.345
cc_64 VNB N_A_887_343#_c_655_n 0.00455982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_887_343#_c_656_n 0.0409408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_887_343#_c_657_n 0.0359155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_887_343#_c_658_n 0.0185667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_RESET_B_M1021_g 0.0286496f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_69 VNB N_RESET_B_c_766_n 0.037544f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_70 VNB N_RESET_B_c_767_n 0.00170088f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_71 VNB N_VPWR_c_810_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB Q 0.0245967f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.18
cc_73 VNB N_Q_c_998_n 0.0564616f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.665
cc_74 VNB N_VGND_c_1016_n 0.0113827f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.85
cc_75 VNB N_VGND_c_1017_n 0.0267104f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.67
cc_76 VNB N_VGND_c_1018_n 0.00383595f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_77 VNB N_VGND_c_1019_n 0.0124398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1020_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1021_n 0.0772001f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.345
cc_80 VNB N_VGND_c_1022_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.345
cc_81 VNB N_VGND_c_1023_n 0.0489774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1024_n 0.0492919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1025_n 0.0641299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1026_n 0.574559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1027_n 0.0059813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1028_n 0.00510127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_862_101#_c_1110_n 0.0128131f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.18
cc_88 VNB N_A_862_101#_c_1111_n 0.0127039f $X=-0.19 $Y=-0.245 $X2=0.855
+ $Y2=0.495
cc_89 VNB N_A_862_101#_c_1112_n 0.0108629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_862_101#_c_1113_n 0.00107216f $X=-0.19 $Y=-0.245 $X2=0.855
+ $Y2=2.67
cc_91 VNB N_A_862_101#_c_1114_n 0.0118439f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.67
cc_92 VNB N_A_862_101#_c_1115_n 0.00138846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_862_101#_c_1116_n 0.00700084f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_94 VPB N_GATE_M1022_g 0.0438416f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.67
cc_95 VPB N_GATE_M1018_g 0.0381401f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.67
cc_96 VPB GATE 0.0337091f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_97 VPB N_GATE_c_169_n 0.021817f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.345
cc_98 VPB N_A_186_57#_M1004_g 0.0212362f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.18
cc_99 VPB N_A_186_57#_M1005_g 0.0183994f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_100 VPB N_A_186_57#_M1017_g 0.0218428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_186_57#_c_217_n 0.0143224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_186_57#_c_206_n 0.00766614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_186_57#_c_219_n 0.00687046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_186_57#_c_220_n 8.1344e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_186_57#_c_211_n 0.0137765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_D_c_332_n 0.0150555f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.85
cc_107 VPB N_D_c_333_n 0.0146071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_D_c_331_n 0.00805965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_294_547#_c_374_n 0.233804f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.67
cc_110 VPB N_A_294_547#_M1027_g 0.0568481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_294_547#_c_370_n 0.0117486f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.85
cc_112 VPB N_A_294_547#_c_371_n 0.00274988f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.67
cc_113 VPB N_A_294_547#_c_373_n 0.0211979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_294_547#_c_379_n 0.0427294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_638_73#_M1000_g 0.0286382f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.67
cc_116 VPB N_A_638_73#_c_444_n 0.0601627f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_117 VPB N_A_638_73#_c_445_n 0.02984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_638_73#_c_439_n 0.0101846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_638_73#_c_440_n 4.57665e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_638_73#_c_448_n 0.0091832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_638_73#_c_449_n 0.0178057f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.345
cc_122 VPB N_A_1208_75#_M1009_g 0.0338575f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.67
cc_123 VPB N_A_1208_75#_c_541_n 0.0184194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_1208_75#_c_531_n 0.00785968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_1208_75#_M1024_g 0.0239117f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.345
cc_126 VPB N_A_1208_75#_c_544_n 0.0181128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_1208_75#_c_536_n 0.00417418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_1208_75#_c_546_n 0.004276f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_887_343#_M1025_g 0.0256005f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.18
cc_130 VPB N_A_887_343#_M1003_g 0.0239963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_887_343#_c_648_n 0.00522131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_RESET_B_M1012_g 0.0168623f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.67
cc_133 VPB N_RESET_B_M1013_g 0.0180175f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.495
cc_134 VPB N_RESET_B_c_766_n 0.00345318f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_135 VPB N_RESET_B_c_767_n 0.00494962f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_136 VPB N_VPWR_c_811_n 0.0117739f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_812_n 0.0367041f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_138 VPB N_VPWR_c_813_n 0.031787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_814_n 0.0316461f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_815_n 0.00238736f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.345
cc_141 VPB N_VPWR_c_816_n 0.0114857f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_817_n 0.0387563f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.665
cc_143 VPB N_VPWR_c_818_n 0.00356964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_819_n 0.0561353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_820_n 0.0812251f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_821_n 0.0427435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_822_n 0.0279832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_810_n 0.15632f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_824_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_825_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_826_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_800_343#_c_904_n 0.00582359f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.18
cc_153 VPB N_A_800_343#_c_905_n 0.0239402f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.495
cc_154 VPB N_A_800_343#_c_906_n 0.00425911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_800_343#_c_907_n 0.00447773f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.67
cc_156 VPB N_A_996_343#_c_928_n 0.0288637f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.67
cc_157 VPB N_A_996_343#_c_929_n 0.0174788f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.495
cc_158 VPB N_A_996_343#_c_930_n 0.00936114f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.85
cc_159 VPB N_A_1420_367#_c_953_n 0.00777283f $X=-0.19 $Y=1.655 $X2=0.855
+ $Y2=1.18
cc_160 VPB N_A_1420_367#_c_954_n 0.0217465f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.85
cc_161 VPB N_A_1420_367#_c_955_n 0.00312972f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.21
cc_162 VPB N_A_1420_367#_c_956_n 0.00515167f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_163 VPB N_A_1420_367#_c_957_n 0.00274001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB Q 0.0543794f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.18
cc_165 N_GATE_M1022_g N_A_186_57#_c_217_n 0.00185f $X=0.495 $Y=2.67 $X2=0 $Y2=0
cc_166 N_GATE_M1018_g N_A_186_57#_c_217_n 0.0129496f $X=0.855 $Y=2.67 $X2=0
+ $Y2=0
cc_167 N_GATE_M1010_g N_A_186_57#_c_210_n 0.00125204f $X=0.495 $Y=0.495 $X2=0
+ $Y2=0
cc_168 N_GATE_M1001_g N_A_186_57#_c_210_n 0.0101019f $X=0.855 $Y=0.495 $X2=0
+ $Y2=0
cc_169 N_GATE_M1001_g N_A_186_57#_c_211_n 0.0428073f $X=0.855 $Y=0.495 $X2=0
+ $Y2=0
cc_170 GATE N_A_186_57#_c_211_n 0.0616405f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_171 N_GATE_M1001_g N_A_294_547#_c_373_n 0.00421772f $X=0.855 $Y=0.495 $X2=0
+ $Y2=0
cc_172 N_GATE_M1018_g N_A_294_547#_c_373_n 0.00217183f $X=0.855 $Y=2.67 $X2=0
+ $Y2=0
cc_173 N_GATE_M1018_g N_A_294_547#_c_379_n 0.00342565f $X=0.855 $Y=2.67 $X2=0
+ $Y2=0
cc_174 N_GATE_M1022_g N_VPWR_c_812_n 0.0167131f $X=0.495 $Y=2.67 $X2=0 $Y2=0
cc_175 N_GATE_M1018_g N_VPWR_c_812_n 0.00252244f $X=0.855 $Y=2.67 $X2=0 $Y2=0
cc_176 GATE N_VPWR_c_812_n 0.0283856f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_177 N_GATE_M1022_g N_VPWR_c_819_n 0.0040395f $X=0.495 $Y=2.67 $X2=0 $Y2=0
cc_178 N_GATE_M1018_g N_VPWR_c_819_n 0.00457319f $X=0.855 $Y=2.67 $X2=0 $Y2=0
cc_179 N_GATE_M1022_g N_VPWR_c_810_n 0.00772493f $X=0.495 $Y=2.67 $X2=0 $Y2=0
cc_180 N_GATE_M1018_g N_VPWR_c_810_n 0.00904779f $X=0.855 $Y=2.67 $X2=0 $Y2=0
cc_181 N_GATE_M1010_g N_VGND_c_1017_n 0.0143087f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_182 N_GATE_M1001_g N_VGND_c_1017_n 0.002112f $X=0.855 $Y=0.495 $X2=0 $Y2=0
cc_183 GATE N_VGND_c_1017_n 0.0147872f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_184 N_GATE_M1010_g N_VGND_c_1023_n 0.00445056f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_185 N_GATE_M1001_g N_VGND_c_1023_n 0.00502664f $X=0.855 $Y=0.495 $X2=0 $Y2=0
cc_186 N_GATE_M1010_g N_VGND_c_1026_n 0.00796275f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_187 N_GATE_M1001_g N_VGND_c_1026_n 0.010303f $X=0.855 $Y=0.495 $X2=0 $Y2=0
cc_188 N_A_186_57#_c_198_n N_D_M1019_g 0.0137745f $X=2.325 $Y=0.895 $X2=0 $Y2=0
cc_189 N_A_186_57#_c_205_n N_D_M1019_g 9.1728e-19 $X=2.145 $Y=1.06 $X2=0 $Y2=0
cc_190 N_A_186_57#_c_206_n N_D_M1019_g 0.0106443f $X=2.145 $Y=1.06 $X2=0 $Y2=0
cc_191 N_A_186_57#_c_208_n N_D_M1019_g 9.44732e-19 $X=3.32 $Y=1.06 $X2=0 $Y2=0
cc_192 N_A_186_57#_M1005_g N_D_c_332_n 0.00982214f $X=2.355 $Y=2.045 $X2=0 $Y2=0
cc_193 N_A_186_57#_c_219_n N_D_c_332_n 0.0124848f $X=3.15 $Y=1.675 $X2=0 $Y2=0
cc_194 N_A_186_57#_c_208_n N_D_M1020_g 0.00664092f $X=3.32 $Y=1.06 $X2=0 $Y2=0
cc_195 N_A_186_57#_c_213_n N_D_M1020_g 0.0181479f $X=3.76 $Y=1.06 $X2=0 $Y2=0
cc_196 N_A_186_57#_c_219_n N_D_c_333_n 0.00420196f $X=3.15 $Y=1.675 $X2=0 $Y2=0
cc_197 N_A_186_57#_c_237_p N_D_c_330_n 0.022394f $X=2.145 $Y=1.59 $X2=0 $Y2=0
cc_198 N_A_186_57#_c_206_n N_D_c_330_n 0.00267252f $X=2.145 $Y=1.06 $X2=0 $Y2=0
cc_199 N_A_186_57#_c_219_n N_D_c_330_n 0.0323819f $X=3.15 $Y=1.675 $X2=0 $Y2=0
cc_200 N_A_186_57#_c_207_n N_D_c_330_n 0.0128896f $X=3.235 $Y=1.59 $X2=0 $Y2=0
cc_201 N_A_186_57#_c_208_n N_D_c_330_n 0.0111789f $X=3.32 $Y=1.06 $X2=0 $Y2=0
cc_202 N_A_186_57#_c_237_p N_D_c_331_n 0.00118505f $X=2.145 $Y=1.59 $X2=0 $Y2=0
cc_203 N_A_186_57#_c_206_n N_D_c_331_n 0.0314198f $X=2.145 $Y=1.06 $X2=0 $Y2=0
cc_204 N_A_186_57#_c_219_n N_D_c_331_n 0.0179689f $X=3.15 $Y=1.675 $X2=0 $Y2=0
cc_205 N_A_186_57#_c_207_n N_D_c_331_n 0.0205187f $X=3.235 $Y=1.59 $X2=0 $Y2=0
cc_206 N_A_186_57#_c_208_n N_D_c_331_n 0.00417158f $X=3.32 $Y=1.06 $X2=0 $Y2=0
cc_207 N_A_186_57#_c_209_n N_D_c_331_n 0.00462155f $X=3.595 $Y=1.06 $X2=0 $Y2=0
cc_208 N_A_186_57#_c_213_n N_D_c_331_n 9.3041e-19 $X=3.76 $Y=1.06 $X2=0 $Y2=0
cc_209 N_A_186_57#_c_204_n N_A_294_547#_M1006_s 0.00472846f $X=1.98 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_210 N_A_186_57#_M1005_g N_A_294_547#_c_374_n 0.00949186f $X=2.355 $Y=2.045
+ $X2=0 $Y2=0
cc_211 N_A_186_57#_M1017_g N_A_294_547#_c_374_n 0.00713917f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_212 N_A_186_57#_M1017_g N_A_294_547#_c_371_n 0.020676f $X=4.36 $Y=2.035 $X2=0
+ $Y2=0
cc_213 N_A_186_57#_c_201_n N_A_294_547#_c_371_n 0.00143727f $X=4.71 $Y=1.11
+ $X2=0 $Y2=0
cc_214 N_A_186_57#_M1017_g N_A_294_547#_M1026_g 0.00240397f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_215 N_A_186_57#_c_202_n N_A_294_547#_M1026_g 0.0193572f $X=4.785 $Y=1.035
+ $X2=0 $Y2=0
cc_216 N_A_186_57#_M1004_g N_A_294_547#_c_373_n 0.0225411f $X=1.845 $Y=2.045
+ $X2=0 $Y2=0
cc_217 N_A_186_57#_c_197_n N_A_294_547#_c_373_n 0.00895952f $X=1.965 $Y=0.895
+ $X2=0 $Y2=0
cc_218 N_A_186_57#_M1005_g N_A_294_547#_c_373_n 0.00271871f $X=2.355 $Y=2.045
+ $X2=0 $Y2=0
cc_219 N_A_186_57#_c_204_n N_A_294_547#_c_373_n 0.0242549f $X=1.98 $Y=0.35 $X2=0
+ $Y2=0
cc_220 N_A_186_57#_c_206_n N_A_294_547#_c_373_n 0.0217711f $X=2.145 $Y=1.06
+ $X2=0 $Y2=0
cc_221 N_A_186_57#_c_220_n N_A_294_547#_c_373_n 0.0136826f $X=2.31 $Y=1.675
+ $X2=0 $Y2=0
cc_222 N_A_186_57#_c_210_n N_A_294_547#_c_373_n 0.157073f $X=1.07 $Y=0.35 $X2=0
+ $Y2=0
cc_223 N_A_186_57#_c_212_n N_A_294_547#_c_373_n 0.0702876f $X=2.145 $Y=0.895
+ $X2=0 $Y2=0
cc_224 N_A_186_57#_M1004_g N_A_294_547#_c_379_n 0.00942354f $X=1.845 $Y=2.045
+ $X2=0 $Y2=0
cc_225 N_A_186_57#_c_217_n N_A_294_547#_c_379_n 0.00117448f $X=1.07 $Y=2.495
+ $X2=0 $Y2=0
cc_226 N_A_186_57#_c_199_n N_A_638_73#_c_438_n 0.00522237f $X=4.285 $Y=1.11
+ $X2=0 $Y2=0
cc_227 N_A_186_57#_c_209_n N_A_638_73#_c_438_n 0.0190769f $X=3.595 $Y=1.06 $X2=0
+ $Y2=0
cc_228 N_A_186_57#_c_213_n N_A_638_73#_c_438_n 0.00590329f $X=3.76 $Y=1.06 $X2=0
+ $Y2=0
cc_229 N_A_186_57#_M1017_g N_A_638_73#_c_445_n 0.00633523f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_230 N_A_186_57#_c_219_n N_A_638_73#_c_445_n 0.0119525f $X=3.15 $Y=1.675 $X2=0
+ $Y2=0
cc_231 N_A_186_57#_c_207_n N_A_638_73#_c_445_n 9.89606e-19 $X=3.235 $Y=1.59
+ $X2=0 $Y2=0
cc_232 N_A_186_57#_c_199_n N_A_638_73#_c_439_n 0.00580739f $X=4.285 $Y=1.11
+ $X2=0 $Y2=0
cc_233 N_A_186_57#_M1017_g N_A_638_73#_c_439_n 0.00389227f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_234 N_A_186_57#_c_209_n N_A_638_73#_c_439_n 6.83737e-19 $X=3.595 $Y=1.06
+ $X2=0 $Y2=0
cc_235 N_A_186_57#_c_213_n N_A_638_73#_c_439_n 2.20499e-19 $X=3.76 $Y=1.06 $X2=0
+ $Y2=0
cc_236 N_A_186_57#_c_207_n N_A_638_73#_c_440_n 0.0132435f $X=3.235 $Y=1.59 $X2=0
+ $Y2=0
cc_237 N_A_186_57#_c_209_n N_A_638_73#_c_440_n 0.0201951f $X=3.595 $Y=1.06 $X2=0
+ $Y2=0
cc_238 N_A_186_57#_c_213_n N_A_638_73#_c_440_n 0.00579521f $X=3.76 $Y=1.06 $X2=0
+ $Y2=0
cc_239 N_A_186_57#_c_199_n N_A_638_73#_c_441_n 0.0184747f $X=4.285 $Y=1.11 $X2=0
+ $Y2=0
cc_240 N_A_186_57#_M1017_g N_A_638_73#_c_441_n 0.00628049f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_241 N_A_186_57#_c_202_n N_A_638_73#_c_441_n 0.00220472f $X=4.785 $Y=1.035
+ $X2=0 $Y2=0
cc_242 N_A_186_57#_c_207_n N_A_638_73#_c_441_n 0.00547627f $X=3.235 $Y=1.59
+ $X2=0 $Y2=0
cc_243 N_A_186_57#_c_209_n N_A_638_73#_c_441_n 0.0243148f $X=3.595 $Y=1.06 $X2=0
+ $Y2=0
cc_244 N_A_186_57#_c_213_n N_A_638_73#_c_441_n 0.00111733f $X=3.76 $Y=1.06 $X2=0
+ $Y2=0
cc_245 N_A_186_57#_c_208_n N_A_638_73#_c_442_n 0.0105441f $X=3.32 $Y=1.06 $X2=0
+ $Y2=0
cc_246 N_A_186_57#_c_209_n N_A_638_73#_c_442_n 0.0135468f $X=3.595 $Y=1.06 $X2=0
+ $Y2=0
cc_247 N_A_186_57#_c_213_n N_A_638_73#_c_442_n 0.00145517f $X=3.76 $Y=1.06 $X2=0
+ $Y2=0
cc_248 N_A_186_57#_M1017_g N_A_887_343#_c_648_n 0.00505242f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_249 N_A_186_57#_M1017_g N_A_887_343#_c_649_n 0.00314361f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_250 N_A_186_57#_c_201_n N_A_887_343#_c_649_n 0.00881261f $X=4.71 $Y=1.11
+ $X2=0 $Y2=0
cc_251 N_A_186_57#_c_202_n N_A_887_343#_c_649_n 0.00896882f $X=4.785 $Y=1.035
+ $X2=0 $Y2=0
cc_252 N_A_186_57#_M1017_g N_A_887_343#_c_651_n 0.00262566f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_253 N_A_186_57#_c_201_n N_A_887_343#_c_651_n 0.0111441f $X=4.71 $Y=1.11 $X2=0
+ $Y2=0
cc_254 N_A_186_57#_c_219_n N_VPWR_M1005_d 0.00845669f $X=3.15 $Y=1.675 $X2=0
+ $Y2=0
cc_255 N_A_186_57#_c_217_n N_VPWR_c_812_n 0.0227343f $X=1.07 $Y=2.495 $X2=0
+ $Y2=0
cc_256 N_A_186_57#_M1004_g N_VPWR_c_813_n 0.00170859f $X=1.845 $Y=2.045 $X2=0
+ $Y2=0
cc_257 N_A_186_57#_M1005_g N_VPWR_c_813_n 0.013624f $X=2.355 $Y=2.045 $X2=0
+ $Y2=0
cc_258 N_A_186_57#_c_219_n N_VPWR_c_813_n 0.0210003f $X=3.15 $Y=1.675 $X2=0
+ $Y2=0
cc_259 N_A_186_57#_c_217_n N_VPWR_c_819_n 0.0165564f $X=1.07 $Y=2.495 $X2=0
+ $Y2=0
cc_260 N_A_186_57#_c_217_n N_VPWR_c_810_n 0.0122141f $X=1.07 $Y=2.495 $X2=0
+ $Y2=0
cc_261 N_A_186_57#_c_220_n A_384_345# 0.0113647f $X=2.31 $Y=1.675 $X2=-0.19
+ $Y2=-0.245
cc_262 N_A_186_57#_c_219_n A_617_345# 0.00423681f $X=3.15 $Y=1.675 $X2=-0.19
+ $Y2=-0.245
cc_263 N_A_186_57#_c_199_n N_A_800_343#_c_904_n 0.00429774f $X=4.285 $Y=1.11
+ $X2=0 $Y2=0
cc_264 N_A_186_57#_M1017_g N_A_800_343#_c_904_n 0.0144034f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_265 N_A_186_57#_M1017_g N_A_800_343#_c_905_n 0.00869532f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_266 N_A_186_57#_M1017_g N_A_800_343#_c_906_n 0.00236801f $X=4.36 $Y=2.035
+ $X2=0 $Y2=0
cc_267 N_A_186_57#_c_210_n N_VGND_c_1017_n 0.0153904f $X=1.07 $Y=0.35 $X2=0
+ $Y2=0
cc_268 N_A_186_57#_c_197_n N_VGND_c_1018_n 5.77822e-19 $X=1.965 $Y=0.895 $X2=0
+ $Y2=0
cc_269 N_A_186_57#_c_198_n N_VGND_c_1018_n 0.00878355f $X=2.325 $Y=0.895 $X2=0
+ $Y2=0
cc_270 N_A_186_57#_c_204_n N_VGND_c_1018_n 0.0114938f $X=1.98 $Y=0.35 $X2=0
+ $Y2=0
cc_271 N_A_186_57#_c_212_n N_VGND_c_1018_n 0.016633f $X=2.145 $Y=0.895 $X2=0
+ $Y2=0
cc_272 N_A_186_57#_c_202_n N_VGND_c_1021_n 7.10185e-19 $X=4.785 $Y=1.035 $X2=0
+ $Y2=0
cc_273 N_A_186_57#_c_197_n N_VGND_c_1023_n 0.00282277f $X=1.965 $Y=0.895 $X2=0
+ $Y2=0
cc_274 N_A_186_57#_c_198_n N_VGND_c_1023_n 0.00386543f $X=2.325 $Y=0.895 $X2=0
+ $Y2=0
cc_275 N_A_186_57#_c_204_n N_VGND_c_1023_n 0.0561449f $X=1.98 $Y=0.35 $X2=0
+ $Y2=0
cc_276 N_A_186_57#_c_210_n N_VGND_c_1023_n 0.0217285f $X=1.07 $Y=0.35 $X2=0
+ $Y2=0
cc_277 N_A_186_57#_c_197_n N_VGND_c_1026_n 0.00371134f $X=1.965 $Y=0.895 $X2=0
+ $Y2=0
cc_278 N_A_186_57#_c_198_n N_VGND_c_1026_n 0.00759904f $X=2.325 $Y=0.895 $X2=0
+ $Y2=0
cc_279 N_A_186_57#_c_204_n N_VGND_c_1026_n 0.0337288f $X=1.98 $Y=0.35 $X2=0
+ $Y2=0
cc_280 N_A_186_57#_c_210_n N_VGND_c_1026_n 0.0125175f $X=1.07 $Y=0.35 $X2=0
+ $Y2=0
cc_281 N_A_186_57#_c_204_n A_408_73# 6.67573e-19 $X=1.98 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_282 N_A_186_57#_c_212_n A_408_73# 0.00333377f $X=2.145 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_283 N_A_186_57#_c_202_n N_A_862_101#_c_1110_n 0.012303f $X=4.785 $Y=1.035
+ $X2=0 $Y2=0
cc_284 N_A_186_57#_c_203_n N_A_862_101#_c_1110_n 0.0133361f $X=4.36 $Y=1.11
+ $X2=0 $Y2=0
cc_285 N_A_186_57#_c_201_n N_A_862_101#_c_1111_n 0.00194999f $X=4.71 $Y=1.11
+ $X2=0 $Y2=0
cc_286 N_A_186_57#_c_202_n N_A_862_101#_c_1111_n 0.0111814f $X=4.785 $Y=1.035
+ $X2=0 $Y2=0
cc_287 N_A_186_57#_c_202_n N_A_862_101#_c_1113_n 6.38398e-19 $X=4.785 $Y=1.035
+ $X2=0 $Y2=0
cc_288 N_D_c_332_n N_A_294_547#_c_374_n 0.00972832f $X=3.01 $Y=1.615 $X2=0 $Y2=0
cc_289 N_D_c_333_n N_A_294_547#_c_374_n 0.00972832f $X=3.37 $Y=1.615 $X2=0 $Y2=0
cc_290 N_D_c_331_n N_A_638_73#_c_445_n 0.00883365f $X=3.115 $Y=1.347 $X2=0 $Y2=0
cc_291 N_D_c_331_n N_A_638_73#_c_440_n 0.00356167f $X=3.115 $Y=1.347 $X2=0 $Y2=0
cc_292 N_D_M1019_g N_A_638_73#_c_442_n 0.00100708f $X=2.755 $Y=0.575 $X2=0 $Y2=0
cc_293 N_D_M1020_g N_A_638_73#_c_442_n 0.00684272f $X=3.115 $Y=0.575 $X2=0 $Y2=0
cc_294 N_D_c_332_n N_VPWR_c_813_n 0.0137602f $X=3.01 $Y=1.615 $X2=0 $Y2=0
cc_295 N_D_M1019_g N_VGND_c_1018_n 0.0103492f $X=2.755 $Y=0.575 $X2=0 $Y2=0
cc_296 N_D_M1020_g N_VGND_c_1018_n 0.00159305f $X=3.115 $Y=0.575 $X2=0 $Y2=0
cc_297 N_D_c_330_n N_VGND_c_1018_n 0.00715721f $X=2.805 $Y=1.245 $X2=0 $Y2=0
cc_298 N_D_M1019_g N_VGND_c_1021_n 0.00386543f $X=2.755 $Y=0.575 $X2=0 $Y2=0
cc_299 N_D_M1020_g N_VGND_c_1021_n 0.00438034f $X=3.115 $Y=0.575 $X2=0 $Y2=0
cc_300 N_D_M1019_g N_VGND_c_1026_n 0.00759904f $X=2.755 $Y=0.575 $X2=0 $Y2=0
cc_301 N_D_M1020_g N_VGND_c_1026_n 0.00838734f $X=3.115 $Y=0.575 $X2=0 $Y2=0
cc_302 N_A_294_547#_M1026_g N_A_638_73#_M1014_g 0.0314599f $X=5.215 $Y=0.715
+ $X2=0 $Y2=0
cc_303 N_A_294_547#_c_370_n N_A_638_73#_c_437_n 0.0314599f $X=5.14 $Y=1.53 $X2=0
+ $Y2=0
cc_304 N_A_294_547#_c_374_n N_A_638_73#_c_444_n 0.00345459f $X=4.83 $Y=2.81
+ $X2=0 $Y2=0
cc_305 N_A_294_547#_c_374_n N_A_638_73#_c_448_n 0.0218378f $X=4.83 $Y=2.81 $X2=0
+ $Y2=0
cc_306 N_A_294_547#_c_374_n N_A_638_73#_c_449_n 0.057217f $X=4.83 $Y=2.81 $X2=0
+ $Y2=0
cc_307 N_A_294_547#_c_371_n N_A_887_343#_c_648_n 0.0101339f $X=4.98 $Y=1.53
+ $X2=0 $Y2=0
cc_308 N_A_294_547#_c_371_n N_A_887_343#_c_649_n 0.00142156f $X=4.98 $Y=1.53
+ $X2=0 $Y2=0
cc_309 N_A_294_547#_M1026_g N_A_887_343#_c_649_n 0.0071469f $X=5.215 $Y=0.715
+ $X2=0 $Y2=0
cc_310 N_A_294_547#_c_370_n N_A_887_343#_c_650_n 0.00418392f $X=5.14 $Y=1.53
+ $X2=0 $Y2=0
cc_311 N_A_294_547#_M1026_g N_A_887_343#_c_650_n 0.01071f $X=5.215 $Y=0.715
+ $X2=0 $Y2=0
cc_312 N_A_294_547#_c_370_n N_A_887_343#_c_651_n 0.00308211f $X=5.14 $Y=1.53
+ $X2=0 $Y2=0
cc_313 N_A_294_547#_c_371_n N_A_887_343#_c_651_n 0.0096929f $X=4.98 $Y=1.53
+ $X2=0 $Y2=0
cc_314 N_A_294_547#_c_374_n N_VPWR_c_813_n 0.0310734f $X=4.83 $Y=2.81 $X2=0
+ $Y2=0
cc_315 N_A_294_547#_c_373_n N_VPWR_c_813_n 0.0322564f $X=1.635 $Y=0.78 $X2=0
+ $Y2=0
cc_316 N_A_294_547#_c_379_n N_VPWR_c_813_n 0.00297747f $X=1.635 $Y=2.81 $X2=0
+ $Y2=0
cc_317 N_A_294_547#_c_374_n N_VPWR_c_819_n 0.0142367f $X=4.83 $Y=2.81 $X2=0
+ $Y2=0
cc_318 N_A_294_547#_c_373_n N_VPWR_c_819_n 0.021313f $X=1.635 $Y=0.78 $X2=0
+ $Y2=0
cc_319 N_A_294_547#_c_379_n N_VPWR_c_819_n 0.00212849f $X=1.635 $Y=2.81 $X2=0
+ $Y2=0
cc_320 N_A_294_547#_c_374_n N_VPWR_c_820_n 0.024142f $X=4.83 $Y=2.81 $X2=0 $Y2=0
cc_321 N_A_294_547#_c_374_n N_VPWR_c_810_n 0.0352282f $X=4.83 $Y=2.81 $X2=0
+ $Y2=0
cc_322 N_A_294_547#_c_373_n N_VPWR_c_810_n 0.0126816f $X=1.635 $Y=0.78 $X2=0
+ $Y2=0
cc_323 N_A_294_547#_M1027_g N_A_800_343#_c_904_n 9.30074e-19 $X=4.905 $Y=1.925
+ $X2=0 $Y2=0
cc_324 N_A_294_547#_c_374_n N_A_800_343#_c_905_n 0.00813227f $X=4.83 $Y=2.81
+ $X2=0 $Y2=0
cc_325 N_A_294_547#_M1027_g N_A_800_343#_c_905_n 0.0176462f $X=4.905 $Y=1.925
+ $X2=0 $Y2=0
cc_326 N_A_294_547#_c_374_n N_A_800_343#_c_906_n 0.00621727f $X=4.83 $Y=2.81
+ $X2=0 $Y2=0
cc_327 N_A_294_547#_M1027_g N_A_800_343#_c_907_n 0.00587337f $X=4.905 $Y=1.925
+ $X2=0 $Y2=0
cc_328 N_A_294_547#_M1027_g N_A_996_343#_c_930_n 0.00737697f $X=4.905 $Y=1.925
+ $X2=0 $Y2=0
cc_329 N_A_294_547#_c_370_n N_A_996_343#_c_930_n 0.00775368f $X=5.14 $Y=1.53
+ $X2=0 $Y2=0
cc_330 N_A_294_547#_M1026_g N_VGND_c_1019_n 3.71719e-19 $X=5.215 $Y=0.715 $X2=0
+ $Y2=0
cc_331 N_A_294_547#_M1026_g N_VGND_c_1021_n 7.27864e-19 $X=5.215 $Y=0.715 $X2=0
+ $Y2=0
cc_332 N_A_294_547#_M1026_g N_A_862_101#_c_1111_n 0.00983421f $X=5.215 $Y=0.715
+ $X2=0 $Y2=0
cc_333 N_A_294_547#_M1026_g N_A_862_101#_c_1113_n 0.0109202f $X=5.215 $Y=0.715
+ $X2=0 $Y2=0
cc_334 N_A_294_547#_M1026_g N_A_862_101#_c_1115_n 0.00386949f $X=5.215 $Y=0.715
+ $X2=0 $Y2=0
cc_335 N_A_638_73#_M1014_g N_A_1208_75#_c_523_n 0.0189652f $X=5.605 $Y=0.715
+ $X2=0 $Y2=0
cc_336 N_A_638_73#_M1014_g N_A_1208_75#_M1009_g 0.00435296f $X=5.605 $Y=0.715
+ $X2=0 $Y2=0
cc_337 N_A_638_73#_c_437_n N_A_1208_75#_M1009_g 0.0262304f $X=5.895 $Y=1.5 $X2=0
+ $Y2=0
cc_338 N_A_638_73#_c_439_n N_A_887_343#_c_648_n 0.00294002f $X=3.94 $Y=1.49
+ $X2=0 $Y2=0
cc_339 N_A_638_73#_M1014_g N_A_887_343#_c_650_n 0.00560766f $X=5.605 $Y=0.715
+ $X2=0 $Y2=0
cc_340 N_A_638_73#_c_437_n N_A_887_343#_c_650_n 0.0146777f $X=5.895 $Y=1.5 $X2=0
+ $Y2=0
cc_341 N_A_638_73#_c_439_n N_A_887_343#_c_651_n 0.00575908f $X=3.94 $Y=1.49
+ $X2=0 $Y2=0
cc_342 N_A_638_73#_c_441_n N_A_887_343#_c_651_n 0.00281784f $X=4.025 $Y=1.405
+ $X2=0 $Y2=0
cc_343 N_A_638_73#_M1000_g N_VPWR_c_814_n 0.0197414f $X=5.895 $Y=2.255 $X2=0
+ $Y2=0
cc_344 N_A_638_73#_c_444_n N_VPWR_c_814_n 0.0126542f $X=5.82 $Y=2.9 $X2=0 $Y2=0
cc_345 N_A_638_73#_c_449_n N_VPWR_c_814_n 0.0250026f $X=5.6 $Y=2.9 $X2=0 $Y2=0
cc_346 N_A_638_73#_c_444_n N_VPWR_c_820_n 0.0136565f $X=5.82 $Y=2.9 $X2=0 $Y2=0
cc_347 N_A_638_73#_c_448_n N_VPWR_c_820_n 0.0168561f $X=3.75 $Y=2.9 $X2=0 $Y2=0
cc_348 N_A_638_73#_c_449_n N_VPWR_c_820_n 0.126939f $X=5.6 $Y=2.9 $X2=0 $Y2=0
cc_349 N_A_638_73#_c_444_n N_VPWR_c_810_n 0.0167424f $X=5.82 $Y=2.9 $X2=0 $Y2=0
cc_350 N_A_638_73#_c_448_n N_VPWR_c_810_n 0.00967329f $X=3.75 $Y=2.9 $X2=0 $Y2=0
cc_351 N_A_638_73#_c_449_n N_VPWR_c_810_n 0.0762676f $X=5.6 $Y=2.9 $X2=0 $Y2=0
cc_352 N_A_638_73#_c_445_n N_A_800_343#_c_904_n 0.0415657f $X=3.585 $Y=1.87
+ $X2=0 $Y2=0
cc_353 N_A_638_73#_c_439_n N_A_800_343#_c_904_n 0.0114066f $X=3.94 $Y=1.49 $X2=0
+ $Y2=0
cc_354 N_A_638_73#_c_444_n N_A_800_343#_c_905_n 0.00750991f $X=5.82 $Y=2.9 $X2=0
+ $Y2=0
cc_355 N_A_638_73#_c_449_n N_A_800_343#_c_905_n 0.103305f $X=5.6 $Y=2.9 $X2=0
+ $Y2=0
cc_356 N_A_638_73#_c_445_n N_A_800_343#_c_906_n 0.0119252f $X=3.585 $Y=1.87
+ $X2=0 $Y2=0
cc_357 N_A_638_73#_c_449_n N_A_800_343#_c_906_n 0.0255786f $X=5.6 $Y=2.9 $X2=0
+ $Y2=0
cc_358 N_A_638_73#_M1000_g N_A_996_343#_c_928_n 0.0167789f $X=5.895 $Y=2.255
+ $X2=0 $Y2=0
cc_359 N_A_638_73#_c_437_n N_A_996_343#_c_928_n 0.00706626f $X=5.895 $Y=1.5
+ $X2=0 $Y2=0
cc_360 N_A_638_73#_M1000_g N_A_996_343#_c_929_n 9.5372e-19 $X=5.895 $Y=2.255
+ $X2=0 $Y2=0
cc_361 N_A_638_73#_M1000_g N_A_996_343#_c_930_n 0.00514523f $X=5.895 $Y=2.255
+ $X2=0 $Y2=0
cc_362 N_A_638_73#_c_442_n N_VGND_c_1018_n 0.0123792f $X=3.33 $Y=0.53 $X2=0
+ $Y2=0
cc_363 N_A_638_73#_M1014_g N_VGND_c_1019_n 0.00737328f $X=5.605 $Y=0.715 $X2=0
+ $Y2=0
cc_364 N_A_638_73#_M1014_g N_VGND_c_1021_n 0.00402651f $X=5.605 $Y=0.715 $X2=0
+ $Y2=0
cc_365 N_A_638_73#_c_438_n N_VGND_c_1021_n 0.01414f $X=3.94 $Y=0.63 $X2=0 $Y2=0
cc_366 N_A_638_73#_c_442_n N_VGND_c_1021_n 0.0142325f $X=3.33 $Y=0.53 $X2=0
+ $Y2=0
cc_367 N_A_638_73#_M1014_g N_VGND_c_1026_n 0.00423264f $X=5.605 $Y=0.715 $X2=0
+ $Y2=0
cc_368 N_A_638_73#_c_438_n N_VGND_c_1026_n 0.0191329f $X=3.94 $Y=0.63 $X2=0
+ $Y2=0
cc_369 N_A_638_73#_c_442_n N_VGND_c_1026_n 0.0117991f $X=3.33 $Y=0.53 $X2=0
+ $Y2=0
cc_370 N_A_638_73#_c_438_n N_A_862_101#_c_1110_n 0.0143282f $X=3.94 $Y=0.63
+ $X2=0 $Y2=0
cc_371 N_A_638_73#_c_441_n N_A_862_101#_c_1110_n 0.0174794f $X=4.025 $Y=1.405
+ $X2=0 $Y2=0
cc_372 N_A_638_73#_M1014_g N_A_862_101#_c_1111_n 4.7271e-19 $X=5.605 $Y=0.715
+ $X2=0 $Y2=0
cc_373 N_A_638_73#_M1014_g N_A_862_101#_c_1113_n 0.00648371f $X=5.605 $Y=0.715
+ $X2=0 $Y2=0
cc_374 N_A_638_73#_M1014_g N_A_862_101#_c_1114_n 0.0142893f $X=5.605 $Y=0.715
+ $X2=0 $Y2=0
cc_375 N_A_638_73#_c_437_n N_A_862_101#_c_1114_n 0.00164703f $X=5.895 $Y=1.5
+ $X2=0 $Y2=0
cc_376 N_A_638_73#_M1014_g N_A_862_101#_c_1116_n 8.62699e-19 $X=5.605 $Y=0.715
+ $X2=0 $Y2=0
cc_377 N_A_1208_75#_c_544_n N_A_887_343#_M1003_g 0.0105485f $X=9.075 $Y=1.9
+ $X2=0 $Y2=0
cc_378 N_A_1208_75#_c_536_n N_A_887_343#_M1003_g 0.00551413f $X=9.16 $Y=1.815
+ $X2=0 $Y2=0
cc_379 N_A_1208_75#_c_546_n N_A_887_343#_M1003_g 0.00878622f $X=8.465 $Y=1.9
+ $X2=0 $Y2=0
cc_380 N_A_1208_75#_c_525_n N_A_887_343#_c_650_n 0.0080377f $X=6.19 $Y=1.11
+ $X2=0 $Y2=0
cc_381 N_A_1208_75#_M1009_g N_A_887_343#_c_650_n 0.0135653f $X=6.44 $Y=2.145
+ $X2=0 $Y2=0
cc_382 N_A_1208_75#_c_527_n N_A_887_343#_c_650_n 0.0105539f $X=6.675 $Y=1.11
+ $X2=0 $Y2=0
cc_383 N_A_1208_75#_c_534_n N_A_887_343#_c_650_n 0.00103331f $X=6.84 $Y=0.77
+ $X2=0 $Y2=0
cc_384 N_A_1208_75#_c_535_n N_A_887_343#_c_650_n 0.0214407f $X=7.425 $Y=0.73
+ $X2=0 $Y2=0
cc_385 N_A_1208_75#_c_534_n N_A_887_343#_c_652_n 4.20366e-19 $X=6.84 $Y=0.77
+ $X2=0 $Y2=0
cc_386 N_A_1208_75#_c_528_n N_A_887_343#_c_653_n 0.00116143f $X=9.21 $Y=1.185
+ $X2=0 $Y2=0
cc_387 N_A_1208_75#_c_560_p N_A_887_343#_c_653_n 0.0835529f $X=9.075 $Y=0.73
+ $X2=0 $Y2=0
cc_388 N_A_1208_75#_c_546_n N_A_887_343#_c_653_n 0.00811187f $X=8.465 $Y=1.9
+ $X2=0 $Y2=0
cc_389 N_A_1208_75#_c_539_n N_A_887_343#_c_653_n 0.0135345f $X=9.27 $Y=1.185
+ $X2=0 $Y2=0
cc_390 N_A_1208_75#_M1015_s N_A_887_343#_c_654_n 0.0027075f $X=7.115 $Y=0.235
+ $X2=0 $Y2=0
cc_391 N_A_1208_75#_c_534_n N_A_887_343#_c_654_n 0.00417388f $X=6.84 $Y=0.77
+ $X2=0 $Y2=0
cc_392 N_A_1208_75#_c_560_p N_A_887_343#_c_654_n 0.00885917f $X=9.075 $Y=0.73
+ $X2=0 $Y2=0
cc_393 N_A_1208_75#_c_535_n N_A_887_343#_c_654_n 0.012199f $X=7.425 $Y=0.73
+ $X2=0 $Y2=0
cc_394 N_A_1208_75#_c_528_n N_A_887_343#_c_655_n 8.04527e-19 $X=9.21 $Y=1.185
+ $X2=0 $Y2=0
cc_395 N_A_1208_75#_c_531_n N_A_887_343#_c_655_n 2.4739e-19 $X=9.645 $Y=1.26
+ $X2=0 $Y2=0
cc_396 N_A_1208_75#_c_544_n N_A_887_343#_c_655_n 0.0187967f $X=9.075 $Y=1.9
+ $X2=0 $Y2=0
cc_397 N_A_1208_75#_c_546_n N_A_887_343#_c_655_n 0.00475343f $X=8.465 $Y=1.9
+ $X2=0 $Y2=0
cc_398 N_A_1208_75#_c_539_n N_A_887_343#_c_655_n 0.0351425f $X=9.27 $Y=1.185
+ $X2=0 $Y2=0
cc_399 N_A_1208_75#_c_531_n N_A_887_343#_c_656_n 0.0130017f $X=9.645 $Y=1.26
+ $X2=0 $Y2=0
cc_400 N_A_1208_75#_c_560_p N_A_887_343#_c_656_n 0.00119253f $X=9.075 $Y=0.73
+ $X2=0 $Y2=0
cc_401 N_A_1208_75#_c_544_n N_A_887_343#_c_656_n 9.56629e-19 $X=9.075 $Y=1.9
+ $X2=0 $Y2=0
cc_402 N_A_1208_75#_c_546_n N_A_887_343#_c_656_n 2.8376e-19 $X=8.465 $Y=1.9
+ $X2=0 $Y2=0
cc_403 N_A_1208_75#_c_538_n N_A_887_343#_c_656_n 0.00242304f $X=9.3 $Y=1.35
+ $X2=0 $Y2=0
cc_404 N_A_1208_75#_M1009_g N_A_887_343#_c_657_n 0.00528299f $X=6.44 $Y=2.145
+ $X2=0 $Y2=0
cc_405 N_A_1208_75#_c_535_n N_A_887_343#_c_657_n 7.72406e-19 $X=7.425 $Y=0.73
+ $X2=0 $Y2=0
cc_406 N_A_1208_75#_c_534_n N_A_887_343#_c_658_n 0.00459166f $X=6.84 $Y=0.77
+ $X2=0 $Y2=0
cc_407 N_A_1208_75#_c_560_p N_A_887_343#_c_658_n 0.00828538f $X=9.075 $Y=0.73
+ $X2=0 $Y2=0
cc_408 N_A_1208_75#_c_535_n N_A_887_343#_c_658_n 0.0108873f $X=7.425 $Y=0.73
+ $X2=0 $Y2=0
cc_409 N_A_1208_75#_c_537_n N_A_887_343#_c_658_n 0.0132571f $X=6.84 $Y=0.43
+ $X2=0 $Y2=0
cc_410 N_A_1208_75#_c_560_p N_RESET_B_M1021_g 0.0134579f $X=9.075 $Y=0.73 $X2=0
+ $Y2=0
cc_411 N_A_1208_75#_c_535_n N_RESET_B_M1021_g 0.00144747f $X=7.425 $Y=0.73 $X2=0
+ $Y2=0
cc_412 N_A_1208_75#_c_546_n N_RESET_B_M1012_g 0.00165516f $X=8.465 $Y=1.9 $X2=0
+ $Y2=0
cc_413 N_A_1208_75#_c_546_n N_RESET_B_M1013_g 0.00680138f $X=8.465 $Y=1.9 $X2=0
+ $Y2=0
cc_414 N_A_1208_75#_M1009_g N_VPWR_c_814_n 0.0059732f $X=6.44 $Y=2.145 $X2=0
+ $Y2=0
cc_415 N_A_1208_75#_c_541_n N_VPWR_c_816_n 0.0271902f $X=9.67 $Y=1.725 $X2=0
+ $Y2=0
cc_416 N_A_1208_75#_c_531_n N_VPWR_c_816_n 0.00456917f $X=9.645 $Y=1.26 $X2=0
+ $Y2=0
cc_417 N_A_1208_75#_M1024_g N_VPWR_c_816_n 0.00378397f $X=10.06 $Y=2.465 $X2=0
+ $Y2=0
cc_418 N_A_1208_75#_c_538_n N_VPWR_c_816_n 0.0049951f $X=9.3 $Y=1.35 $X2=0 $Y2=0
cc_419 N_A_1208_75#_c_541_n N_VPWR_c_822_n 0.00486043f $X=9.67 $Y=1.725 $X2=0
+ $Y2=0
cc_420 N_A_1208_75#_M1024_g N_VPWR_c_822_n 0.00549284f $X=10.06 $Y=2.465 $X2=0
+ $Y2=0
cc_421 N_A_1208_75#_M1013_d N_VPWR_c_810_n 0.00408795f $X=8.325 $Y=1.835 $X2=0
+ $Y2=0
cc_422 N_A_1208_75#_M1009_g N_VPWR_c_810_n 0.0038268f $X=6.44 $Y=2.145 $X2=0
+ $Y2=0
cc_423 N_A_1208_75#_c_541_n N_VPWR_c_810_n 0.00823808f $X=9.67 $Y=1.725 $X2=0
+ $Y2=0
cc_424 N_A_1208_75#_M1024_g N_VPWR_c_810_n 0.0108594f $X=10.06 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_1208_75#_M1009_g N_A_996_343#_c_928_n 0.0156731f $X=6.44 $Y=2.145
+ $X2=0 $Y2=0
cc_426 N_A_1208_75#_M1009_g N_A_996_343#_c_929_n 0.0108073f $X=6.44 $Y=2.145
+ $X2=0 $Y2=0
cc_427 N_A_1208_75#_c_544_n N_A_1420_367#_M1003_d 0.00334849f $X=9.075 $Y=1.9
+ $X2=0 $Y2=0
cc_428 N_A_1208_75#_M1009_g N_A_1420_367#_c_953_n 0.00123097f $X=6.44 $Y=2.145
+ $X2=0 $Y2=0
cc_429 N_A_1208_75#_M1013_d N_A_1420_367#_c_960_n 0.00513066f $X=8.325 $Y=1.835
+ $X2=0 $Y2=0
cc_430 N_A_1208_75#_c_544_n N_A_1420_367#_c_960_n 0.00484169f $X=9.075 $Y=1.9
+ $X2=0 $Y2=0
cc_431 N_A_1208_75#_c_546_n N_A_1420_367#_c_960_n 0.0154328f $X=8.465 $Y=1.9
+ $X2=0 $Y2=0
cc_432 N_A_1208_75#_c_544_n N_A_1420_367#_c_955_n 0.0193955f $X=9.075 $Y=1.9
+ $X2=0 $Y2=0
cc_433 N_A_1208_75#_c_541_n N_A_1420_367#_c_956_n 0.00143001f $X=9.67 $Y=1.725
+ $X2=0 $Y2=0
cc_434 N_A_1208_75#_M1009_g N_A_1420_367#_c_957_n 0.00317961f $X=6.44 $Y=2.145
+ $X2=0 $Y2=0
cc_435 N_A_1208_75#_c_529_n Q 0.00242057f $X=9.57 $Y=1.185 $X2=0 $Y2=0
cc_436 N_A_1208_75#_c_530_n Q 0.00835352f $X=9.985 $Y=1.26 $X2=0 $Y2=0
cc_437 N_A_1208_75#_c_531_n Q 0.00648652f $X=9.645 $Y=1.26 $X2=0 $Y2=0
cc_438 N_A_1208_75#_M1024_g Q 0.0431621f $X=10.06 $Y=2.465 $X2=0 $Y2=0
cc_439 N_A_1208_75#_c_538_n Q 0.00824897f $X=9.3 $Y=1.35 $X2=0 $Y2=0
cc_440 N_A_1208_75#_c_529_n N_Q_c_998_n 0.0028004f $X=9.57 $Y=1.185 $X2=0 $Y2=0
cc_441 N_A_1208_75#_c_530_n N_Q_c_998_n 0.0231955f $X=9.985 $Y=1.26 $X2=0 $Y2=0
cc_442 N_A_1208_75#_c_560_p N_Q_c_998_n 0.00563251f $X=9.075 $Y=0.73 $X2=0 $Y2=0
cc_443 N_A_1208_75#_c_539_n N_Q_c_998_n 0.0118778f $X=9.27 $Y=1.185 $X2=0 $Y2=0
cc_444 N_A_1208_75#_c_560_p N_VGND_M1021_d 0.0409926f $X=9.075 $Y=0.73 $X2=0
+ $Y2=0
cc_445 N_A_1208_75#_c_539_n N_VGND_M1021_d 0.00770091f $X=9.27 $Y=1.185 $X2=0
+ $Y2=0
cc_446 N_A_1208_75#_c_523_n N_VGND_c_1019_n 0.00488538f $X=6.115 $Y=1.035 $X2=0
+ $Y2=0
cc_447 N_A_1208_75#_c_537_n N_VGND_c_1019_n 0.00152724f $X=6.84 $Y=0.43 $X2=0
+ $Y2=0
cc_448 N_A_1208_75#_c_560_p N_VGND_c_1020_n 0.019543f $X=9.075 $Y=0.73 $X2=0
+ $Y2=0
cc_449 N_A_1208_75#_c_535_n N_VGND_c_1020_n 0.0067198f $X=7.425 $Y=0.73 $X2=0
+ $Y2=0
cc_450 N_A_1208_75#_c_523_n N_VGND_c_1024_n 0.00464519f $X=6.115 $Y=1.035 $X2=0
+ $Y2=0
cc_451 N_A_1208_75#_c_560_p N_VGND_c_1024_n 0.00721273f $X=9.075 $Y=0.73 $X2=0
+ $Y2=0
cc_452 N_A_1208_75#_c_535_n N_VGND_c_1024_n 0.0467013f $X=7.425 $Y=0.73 $X2=0
+ $Y2=0
cc_453 N_A_1208_75#_c_537_n N_VGND_c_1024_n 0.00210642f $X=6.84 $Y=0.43 $X2=0
+ $Y2=0
cc_454 N_A_1208_75#_c_528_n N_VGND_c_1025_n 0.00468809f $X=9.21 $Y=1.185 $X2=0
+ $Y2=0
cc_455 N_A_1208_75#_c_529_n N_VGND_c_1025_n 0.00585385f $X=9.57 $Y=1.185 $X2=0
+ $Y2=0
cc_456 N_A_1208_75#_c_560_p N_VGND_c_1025_n 0.0166923f $X=9.075 $Y=0.73 $X2=0
+ $Y2=0
cc_457 N_A_1208_75#_M1015_s N_VGND_c_1026_n 0.00232985f $X=7.115 $Y=0.235 $X2=0
+ $Y2=0
cc_458 N_A_1208_75#_c_523_n N_VGND_c_1026_n 0.00503886f $X=6.115 $Y=1.035 $X2=0
+ $Y2=0
cc_459 N_A_1208_75#_c_528_n N_VGND_c_1026_n 0.00855112f $X=9.21 $Y=1.185 $X2=0
+ $Y2=0
cc_460 N_A_1208_75#_c_529_n N_VGND_c_1026_n 0.0119619f $X=9.57 $Y=1.185 $X2=0
+ $Y2=0
cc_461 N_A_1208_75#_c_560_p N_VGND_c_1026_n 0.0422607f $X=9.075 $Y=0.73 $X2=0
+ $Y2=0
cc_462 N_A_1208_75#_c_535_n N_VGND_c_1026_n 0.0286033f $X=7.425 $Y=0.73 $X2=0
+ $Y2=0
cc_463 N_A_1208_75#_c_523_n N_A_862_101#_c_1114_n 0.00691791f $X=6.115 $Y=1.035
+ $X2=0 $Y2=0
cc_464 N_A_1208_75#_c_524_n N_A_862_101#_c_1114_n 0.00501898f $X=6.365 $Y=1.11
+ $X2=0 $Y2=0
cc_465 N_A_1208_75#_c_525_n N_A_862_101#_c_1114_n 0.00453389f $X=6.19 $Y=1.11
+ $X2=0 $Y2=0
cc_466 N_A_1208_75#_c_533_n N_A_862_101#_c_1114_n 0.0125605f $X=6.44 $Y=1.11
+ $X2=0 $Y2=0
cc_467 N_A_1208_75#_c_534_n N_A_862_101#_c_1114_n 0.00116806f $X=6.84 $Y=0.77
+ $X2=0 $Y2=0
cc_468 N_A_1208_75#_c_523_n N_A_862_101#_c_1116_n 0.00897202f $X=6.115 $Y=1.035
+ $X2=0 $Y2=0
cc_469 N_A_1208_75#_c_534_n N_A_862_101#_c_1116_n 0.00149445f $X=6.84 $Y=0.77
+ $X2=0 $Y2=0
cc_470 N_A_1208_75#_c_535_n N_A_862_101#_c_1116_n 0.0356169f $X=7.425 $Y=0.73
+ $X2=0 $Y2=0
cc_471 N_A_1208_75#_c_537_n N_A_862_101#_c_1116_n 0.00184718f $X=6.84 $Y=0.43
+ $X2=0 $Y2=0
cc_472 N_A_1208_75#_c_560_p A_1510_47# 0.0035945f $X=9.075 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_473 N_A_887_343#_c_652_n N_RESET_B_M1021_g 0.00115197f $X=7.385 $Y=1.345
+ $X2=0 $Y2=0
cc_474 N_A_887_343#_c_653_n N_RESET_B_M1021_g 0.0123392f $X=8.565 $Y=1.08 $X2=0
+ $Y2=0
cc_475 N_A_887_343#_c_655_n N_RESET_B_M1021_g 0.0032399f $X=8.73 $Y=1.46 $X2=0
+ $Y2=0
cc_476 N_A_887_343#_c_656_n N_RESET_B_M1021_g 0.0010385f $X=8.73 $Y=1.46 $X2=0
+ $Y2=0
cc_477 N_A_887_343#_c_658_n N_RESET_B_M1021_g 0.0384018f $X=7.385 $Y=1.185 $X2=0
+ $Y2=0
cc_478 N_A_887_343#_M1025_g N_RESET_B_M1012_g 0.0526651f $X=7.46 $Y=2.465 $X2=0
+ $Y2=0
cc_479 N_A_887_343#_M1025_g N_RESET_B_c_766_n 0.00872802f $X=7.46 $Y=2.465 $X2=0
+ $Y2=0
cc_480 N_A_887_343#_M1003_g N_RESET_B_c_766_n 0.0591893f $X=8.68 $Y=2.465 $X2=0
+ $Y2=0
cc_481 N_A_887_343#_c_652_n N_RESET_B_c_766_n 6.24677e-19 $X=7.385 $Y=1.345
+ $X2=0 $Y2=0
cc_482 N_A_887_343#_c_653_n N_RESET_B_c_766_n 0.00796505f $X=8.565 $Y=1.08 $X2=0
+ $Y2=0
cc_483 N_A_887_343#_c_655_n N_RESET_B_c_766_n 0.0012162f $X=8.73 $Y=1.46 $X2=0
+ $Y2=0
cc_484 N_A_887_343#_c_656_n N_RESET_B_c_766_n 0.00999409f $X=8.73 $Y=1.46 $X2=0
+ $Y2=0
cc_485 N_A_887_343#_c_657_n N_RESET_B_c_766_n 0.0384018f $X=7.385 $Y=1.35 $X2=0
+ $Y2=0
cc_486 N_A_887_343#_M1025_g N_RESET_B_c_767_n 0.00325478f $X=7.46 $Y=2.465 $X2=0
+ $Y2=0
cc_487 N_A_887_343#_M1003_g N_RESET_B_c_767_n 2.09187e-19 $X=8.68 $Y=2.465 $X2=0
+ $Y2=0
cc_488 N_A_887_343#_c_652_n N_RESET_B_c_767_n 0.0102874f $X=7.385 $Y=1.345 $X2=0
+ $Y2=0
cc_489 N_A_887_343#_c_653_n N_RESET_B_c_767_n 0.0236677f $X=8.565 $Y=1.08 $X2=0
+ $Y2=0
cc_490 N_A_887_343#_c_655_n N_RESET_B_c_767_n 0.00963847f $X=8.73 $Y=1.46 $X2=0
+ $Y2=0
cc_491 N_A_887_343#_c_656_n N_RESET_B_c_767_n 0.0010366f $X=8.73 $Y=1.46 $X2=0
+ $Y2=0
cc_492 N_A_887_343#_c_657_n N_RESET_B_c_767_n 2.17416e-19 $X=7.385 $Y=1.35 $X2=0
+ $Y2=0
cc_493 N_A_887_343#_M1025_g N_VPWR_c_815_n 0.0029516f $X=7.46 $Y=2.465 $X2=0
+ $Y2=0
cc_494 N_A_887_343#_M1003_g N_VPWR_c_816_n 0.00327672f $X=8.68 $Y=2.465 $X2=0
+ $Y2=0
cc_495 N_A_887_343#_M1025_g N_VPWR_c_817_n 0.00549284f $X=7.46 $Y=2.465 $X2=0
+ $Y2=0
cc_496 N_A_887_343#_M1003_g N_VPWR_c_821_n 0.00585385f $X=8.68 $Y=2.465 $X2=0
+ $Y2=0
cc_497 N_A_887_343#_M1025_g N_VPWR_c_810_n 0.00741697f $X=7.46 $Y=2.465 $X2=0
+ $Y2=0
cc_498 N_A_887_343#_M1003_g N_VPWR_c_810_n 0.00776999f $X=8.68 $Y=2.465 $X2=0
+ $Y2=0
cc_499 N_A_887_343#_c_648_n N_A_800_343#_c_905_n 0.0196829f $X=4.575 $Y=1.95
+ $X2=0 $Y2=0
cc_500 N_A_887_343#_M1025_g N_A_996_343#_c_928_n 0.00342072f $X=7.46 $Y=2.465
+ $X2=0 $Y2=0
cc_501 N_A_887_343#_c_650_n N_A_996_343#_c_928_n 0.110467f $X=7.22 $Y=1.43 $X2=0
+ $Y2=0
cc_502 N_A_887_343#_M1025_g N_A_996_343#_c_929_n 0.00108655f $X=7.46 $Y=2.465
+ $X2=0 $Y2=0
cc_503 N_A_887_343#_c_648_n N_A_996_343#_c_930_n 0.0292395f $X=4.575 $Y=1.95
+ $X2=0 $Y2=0
cc_504 N_A_887_343#_c_651_n N_A_996_343#_c_930_n 0.0243101f $X=5.085 $Y=1.43
+ $X2=0 $Y2=0
cc_505 N_A_887_343#_M1025_g N_A_1420_367#_c_953_n 0.0115777f $X=7.46 $Y=2.465
+ $X2=0 $Y2=0
cc_506 N_A_887_343#_c_650_n N_A_1420_367#_c_953_n 0.00787821f $X=7.22 $Y=1.43
+ $X2=0 $Y2=0
cc_507 N_A_887_343#_c_652_n N_A_1420_367#_c_953_n 0.0106885f $X=7.385 $Y=1.345
+ $X2=0 $Y2=0
cc_508 N_A_887_343#_c_657_n N_A_1420_367#_c_953_n 0.00121786f $X=7.385 $Y=1.35
+ $X2=0 $Y2=0
cc_509 N_A_887_343#_M1025_g N_A_1420_367#_c_954_n 0.00892791f $X=7.46 $Y=2.465
+ $X2=0 $Y2=0
cc_510 N_A_887_343#_M1025_g N_A_1420_367#_c_960_n 0.0123771f $X=7.46 $Y=2.465
+ $X2=0 $Y2=0
cc_511 N_A_887_343#_M1003_g N_A_1420_367#_c_960_n 0.0107014f $X=8.68 $Y=2.465
+ $X2=0 $Y2=0
cc_512 N_A_887_343#_M1025_g N_A_1420_367#_c_957_n 3.84191e-19 $X=7.46 $Y=2.465
+ $X2=0 $Y2=0
cc_513 N_A_887_343#_c_653_n N_VGND_M1021_d 0.0140407f $X=8.565 $Y=1.08 $X2=0
+ $Y2=0
cc_514 N_A_887_343#_c_658_n N_VGND_c_1020_n 0.00180232f $X=7.385 $Y=1.185 $X2=0
+ $Y2=0
cc_515 N_A_887_343#_c_658_n N_VGND_c_1024_n 0.0041543f $X=7.385 $Y=1.185 $X2=0
+ $Y2=0
cc_516 N_A_887_343#_c_658_n N_VGND_c_1026_n 0.00726304f $X=7.385 $Y=1.185 $X2=0
+ $Y2=0
cc_517 N_A_887_343#_c_649_n N_A_862_101#_c_1110_n 0.0209892f $X=5 $Y=0.78 $X2=0
+ $Y2=0
cc_518 N_A_887_343#_c_651_n N_A_862_101#_c_1110_n 0.00598905f $X=5.085 $Y=1.43
+ $X2=0 $Y2=0
cc_519 N_A_887_343#_c_649_n N_A_862_101#_c_1111_n 0.0159778f $X=5 $Y=0.78 $X2=0
+ $Y2=0
cc_520 N_A_887_343#_c_649_n N_A_862_101#_c_1113_n 0.0149126f $X=5 $Y=0.78 $X2=0
+ $Y2=0
cc_521 N_A_887_343#_c_650_n N_A_862_101#_c_1114_n 0.0757928f $X=7.22 $Y=1.43
+ $X2=0 $Y2=0
cc_522 N_A_887_343#_c_649_n N_A_862_101#_c_1115_n 0.0133775f $X=5 $Y=0.78 $X2=0
+ $Y2=0
cc_523 N_A_887_343#_c_650_n N_A_862_101#_c_1115_n 0.0135788f $X=7.22 $Y=1.43
+ $X2=0 $Y2=0
cc_524 N_A_887_343#_c_653_n A_1510_47# 0.00137516f $X=8.565 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_525 N_RESET_B_M1012_g N_VPWR_c_815_n 0.0121516f $X=7.89 $Y=2.465 $X2=0 $Y2=0
cc_526 N_RESET_B_M1013_g N_VPWR_c_815_n 0.00322247f $X=8.25 $Y=2.465 $X2=0 $Y2=0
cc_527 N_RESET_B_M1012_g N_VPWR_c_821_n 0.00486043f $X=7.89 $Y=2.465 $X2=0 $Y2=0
cc_528 N_RESET_B_M1013_g N_VPWR_c_821_n 0.00585385f $X=8.25 $Y=2.465 $X2=0 $Y2=0
cc_529 N_RESET_B_M1012_g N_VPWR_c_810_n 0.00439806f $X=7.89 $Y=2.465 $X2=0 $Y2=0
cc_530 N_RESET_B_M1013_g N_VPWR_c_810_n 0.00633756f $X=8.25 $Y=2.465 $X2=0 $Y2=0
cc_531 N_RESET_B_M1012_g N_A_1420_367#_c_953_n 0.00248418f $X=7.89 $Y=2.465
+ $X2=0 $Y2=0
cc_532 N_RESET_B_M1012_g N_A_1420_367#_c_954_n 0.00100275f $X=7.89 $Y=2.465
+ $X2=0 $Y2=0
cc_533 N_RESET_B_M1012_g N_A_1420_367#_c_960_n 0.0131077f $X=7.89 $Y=2.465 $X2=0
+ $Y2=0
cc_534 N_RESET_B_M1013_g N_A_1420_367#_c_960_n 0.0153692f $X=8.25 $Y=2.465 $X2=0
+ $Y2=0
cc_535 N_RESET_B_c_767_n N_A_1420_367#_c_960_n 0.00914201f $X=7.955 $Y=1.51
+ $X2=0 $Y2=0
cc_536 N_RESET_B_M1021_g N_VGND_c_1020_n 0.0100629f $X=7.865 $Y=0.655 $X2=0
+ $Y2=0
cc_537 N_RESET_B_M1021_g N_VGND_c_1024_n 0.00354752f $X=7.865 $Y=0.655 $X2=0
+ $Y2=0
cc_538 N_RESET_B_M1021_g N_VGND_c_1026_n 0.00413095f $X=7.865 $Y=0.655 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_814_n N_A_996_343#_c_928_n 0.0234047f $X=6.11 $Y=2.32 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_814_n N_A_996_343#_c_929_n 0.0214166f $X=6.11 $Y=2.32 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_810_n N_A_1420_367#_M1025_s 0.0023218f $X=10.32 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_542 N_VPWR_c_810_n N_A_1420_367#_M1003_d 0.00266738f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_817_n N_A_1420_367#_c_954_n 0.019758f $X=7.59 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_810_n N_A_1420_367#_c_954_n 0.012508f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_M1025_d N_A_1420_367#_c_960_n 0.00811522f $X=7.535 $Y=1.835 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_815_n N_A_1420_367#_c_960_n 0.0142991f $X=7.675 $Y=2.895 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_810_n N_A_1420_367#_c_960_n 0.0366801f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_816_n N_A_1420_367#_c_955_n 0.0227647f $X=9.455 $Y=2.33 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_816_n N_A_1420_367#_c_956_n 0.0376052f $X=9.455 $Y=2.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_821_n N_A_1420_367#_c_956_n 0.0163773f $X=9.29 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_810_n N_A_1420_367#_c_956_n 0.00959046f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_810_n A_1593_367# 0.00306596f $X=10.32 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_553 N_VPWR_c_810_n A_1949_367# 0.010279f $X=10.32 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_554 N_VPWR_c_810_n N_Q_M1024_d 0.0023218f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_555 N_VPWR_c_816_n Q 0.0285126f $X=9.455 $Y=2.33 $X2=0 $Y2=0
cc_556 N_VPWR_c_822_n Q 0.019758f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_557 N_VPWR_c_810_n Q 0.012508f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_558 N_A_800_343#_c_905_n N_A_996_343#_c_928_n 0.00796895f $X=5.515 $Y=2.47
+ $X2=0 $Y2=0
cc_559 N_A_800_343#_c_907_n N_A_996_343#_c_928_n 0.0192142f $X=5.68 $Y=2.3 $X2=0
+ $Y2=0
cc_560 N_A_800_343#_c_905_n N_A_996_343#_c_930_n 0.0214984f $X=5.515 $Y=2.47
+ $X2=0 $Y2=0
cc_561 N_A_800_343#_c_907_n N_A_996_343#_c_930_n 0.00726339f $X=5.68 $Y=2.3
+ $X2=0 $Y2=0
cc_562 N_A_996_343#_c_928_n N_A_1420_367#_c_953_n 0.00328588f $X=6.49 $Y=1.78
+ $X2=0 $Y2=0
cc_563 N_A_996_343#_c_929_n N_A_1420_367#_c_953_n 0.0284373f $X=6.655 $Y=2.145
+ $X2=0 $Y2=0
cc_564 N_A_996_343#_c_929_n N_A_1420_367#_c_957_n 0.00328588f $X=6.655 $Y=2.145
+ $X2=0 $Y2=0
cc_565 N_A_1420_367#_c_960_n A_1593_367# 0.00366956f $X=8.81 $Y=2.41 $X2=-0.19
+ $Y2=1.655
cc_566 N_Q_c_998_n N_VGND_c_1025_n 0.0512239f $X=9.81 $Y=0.43 $X2=0 $Y2=0
cc_567 N_Q_M1007_d N_VGND_c_1026_n 0.00253148f $X=9.645 $Y=0.235 $X2=0 $Y2=0
cc_568 N_Q_c_998_n N_VGND_c_1026_n 0.0306837f $X=9.81 $Y=0.43 $X2=0 $Y2=0
cc_569 N_VGND_c_1019_n N_A_862_101#_c_1111_n 0.0122875f $X=5.82 $Y=0.65 $X2=0
+ $Y2=0
cc_570 N_VGND_c_1021_n N_A_862_101#_c_1111_n 0.0505168f $X=5.655 $Y=0 $X2=0
+ $Y2=0
cc_571 N_VGND_c_1026_n N_A_862_101#_c_1111_n 0.0306752f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_572 N_VGND_c_1021_n N_A_862_101#_c_1112_n 0.0222501f $X=5.655 $Y=0 $X2=0
+ $Y2=0
cc_573 N_VGND_c_1026_n N_A_862_101#_c_1112_n 0.0127687f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_574 N_VGND_c_1019_n N_A_862_101#_c_1113_n 0.0230722f $X=5.82 $Y=0.65 $X2=0
+ $Y2=0
cc_575 N_VGND_c_1019_n N_A_862_101#_c_1114_n 0.0233214f $X=5.82 $Y=0.65 $X2=0
+ $Y2=0
cc_576 N_VGND_c_1019_n N_A_862_101#_c_1116_n 0.0125869f $X=5.82 $Y=0.65 $X2=0
+ $Y2=0
cc_577 N_VGND_c_1024_n N_A_862_101#_c_1116_n 0.00937762f $X=7.915 $Y=0 $X2=0
+ $Y2=0
cc_578 N_VGND_c_1026_n N_A_862_101#_c_1116_n 0.0110641f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_579 N_VGND_c_1026_n A_1510_47# 0.00282558f $X=10.32 $Y=0 $X2=-0.19 $Y2=-0.245
cc_580 N_VGND_c_1026_n A_1857_47# 0.00899413f $X=10.32 $Y=0 $X2=-0.19 $Y2=-0.245
cc_581 N_A_862_101#_c_1113_n A_1058_101# 0.0040322f $X=5.35 $Y=0.995 $X2=-0.19
+ $Y2=-0.245
