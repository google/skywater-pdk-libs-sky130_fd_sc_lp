* NGSPICE file created from sky130_fd_sc_lp__a2bb2oi_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2bb2oi_lp A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 VGND A1_N a_652_47# VNB nshort w=420000u l=150000u
+  ad=3.612e+11p pd=4.24e+06u as=8.82e+10p ps=1.26e+06u
M1001 Y B2 a_170_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.008e+11p ps=1.32e+06u
M1002 Y a_296_146# a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.8e+11p pd=2.56e+06u as=5.65e+11p ps=5.13e+06u
M1003 VPWR B1 a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1004 VGND a_296_146# a_334_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1005 a_652_47# A1_N a_296_146# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1006 a_334_47# a_296_146# Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_409# B2 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_296_146# A2_N a_456_339# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=5.7e+11p ps=5.14e+06u
M1009 VPWR A1_N a_456_339# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_170_47# B1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_494_47# A2_N VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1012 a_296_146# A2_N a_494_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

