# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o21bai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o21bai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 1.375000 2.795000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.580000 1.375000 2.255000 1.750000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.185000 0.515000 1.890000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.764400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.080000 0.255000 1.410000 1.015000 ;
        RECT 1.240000 1.015000 1.410000 1.930000 ;
        RECT 1.240000 1.930000 1.925000 2.100000 ;
        RECT 1.595000 2.100000 1.925000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.095000  0.385000 0.355000 0.845000 ;
      RECT 0.095000  0.845000 0.910000 1.015000 ;
      RECT 0.525000  0.085000 0.855000 0.675000 ;
      RECT 0.570000  2.060000 0.900000 2.390000 ;
      RECT 0.685000  1.015000 0.910000 1.185000 ;
      RECT 0.685000  1.185000 1.070000 1.515000 ;
      RECT 0.685000  1.515000 0.900000 2.060000 ;
      RECT 1.070000  2.270000 1.425000 3.245000 ;
      RECT 1.580000  0.255000 1.810000 1.035000 ;
      RECT 1.580000  1.035000 2.785000 1.205000 ;
      RECT 1.980000  0.085000 2.310000 0.865000 ;
      RECT 2.455000  1.920000 2.785000 3.245000 ;
      RECT 2.480000  0.255000 2.785000 1.035000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_lp__o21bai_1
END LIBRARY
