* File: sky130_fd_sc_lp__a2bb2o_lp.spice
* Created: Fri Aug 28 09:56:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2o_lp.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2o_lp  VNB VPB B2 B1 A1_N A2_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2_N	A2_N
* A1_N	A1_N
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1009 A_150_57# N_B2_M1009_g N_A_63_57#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_B1_M1007_g A_150_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1012 A_314_57# N_A_284_31#_M1012_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_63_57#_M1014_d N_A_284_31#_M1014_g A_314_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 A_584_74# N_A_63_57#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_63_57#_M1011_g A_584_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 A_742_74# N_A1_N_M1000_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1013 N_A_284_31#_M1013_d N_A1_N_M1013_g A_742_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 A_900_74# N_A2_N_M1001_g N_A_284_31#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A2_N_M1004_g A_900_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_B2_M1008_g N_A_43_408#_M1008_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1002 N_A_43_408#_M1002_d N_B1_M1002_g N_VPWR_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.1525 AS=0.14 PD=1.305 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1005 N_A_63_57#_M1005_d N_A_284_31#_M1005_g N_A_43_408#_M1002_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.59 AS=0.1525 PD=3.18 PS=1.305 NRD=60.0653 NRS=4.9053 M=1 R=4
+ SA=125001 SB=125000 A=0.25 P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_A_63_57#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.22 AS=0.285 PD=1.44 PS=2.57 NRD=15.7403 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1006 A_794_409# N_A1_N_M1006_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.22 PD=1.24 PS=1.44 NRD=12.7853 NRS=15.7403 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1015 N_A_284_31#_M1015_d N_A2_N_M1015_g A_794_409# VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.12 PD=2.57 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5559 P=15.05
c_98 VPB 0 1.45652e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a2bb2o_lp.pxi.spice"
*
.ends
*
*
