* File: sky130_fd_sc_lp__a2bb2oi_4.pex.spice
* Created: Fri Aug 28 09:56:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%B1 3 7 11 15 19 23 27 29 31 33 41 47 48 52
+ 61
c121 47 0 9.18783e-20 $X=3.6 $Y=1.295
c122 27 0 8.05408e-21 $X=3.72 $Y=0.655
r123 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=1.375 $X2=3.74 $Y2=1.375
r124 60 61 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.565 $Y=1.46
+ $X2=1.57 $Y2=1.46
r125 57 58 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.135 $Y=1.46
+ $X2=1.14 $Y2=1.46
r126 56 57 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=0.71 $Y=1.46
+ $X2=1.135 $Y2=1.46
r127 55 56 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.705 $Y=1.46
+ $X2=0.71 $Y2=1.46
r128 52 55 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.63 $Y=1.46
+ $X2=0.705 $Y2=1.46
r129 48 65 8.89542 $w=3.18e-07 $l=2.47e-07 $layer=LI1_cond $X=3.665 $Y=1.622
+ $X2=3.665 $Y2=1.375
r130 47 65 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=3.665 $Y=1.295
+ $X2=3.665 $Y2=1.375
r131 42 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=1.75
+ $X2=1.72 $Y2=1.75
r132 41 48 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.505 $Y=1.75
+ $X2=3.665 $Y2=1.75
r133 41 42 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=3.505 $Y=1.75
+ $X2=1.805 $Y2=1.75
r134 40 60 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.48 $Y=1.46
+ $X2=1.565 $Y2=1.46
r135 40 58 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.48 $Y=1.46
+ $X2=1.14 $Y2=1.46
r136 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.48
+ $Y=1.46 $X2=1.48 $Y2=1.46
r137 36 52 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.46 $Y=1.46
+ $X2=0.63 $Y2=1.46
r138 35 39 55.184 $w=2.03e-07 $l=1.02e-06 $layer=LI1_cond $X=0.46 $Y=1.452
+ $X2=1.48 $Y2=1.452
r139 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.46
+ $Y=1.46 $X2=0.46 $Y2=1.46
r140 33 45 19.4417 $w=1.68e-07 $l=2.98e-07 $layer=LI1_cond $X=1.72 $Y=1.452
+ $X2=1.72 $Y2=1.75
r141 33 39 8.38581 $w=2.03e-07 $l=1.55e-07 $layer=LI1_cond $X=1.635 $Y=1.452
+ $X2=1.48 $Y2=1.452
r142 29 64 38.7839 $w=3.5e-07 $l=2.14173e-07 $layer=POLY_cond $X=3.875 $Y=1.54
+ $X2=3.762 $Y2=1.375
r143 29 31 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.875 $Y=1.54
+ $X2=3.875 $Y2=2.465
r144 25 64 38.7839 $w=3.5e-07 $l=1.84811e-07 $layer=POLY_cond $X=3.72 $Y=1.21
+ $X2=3.762 $Y2=1.375
r145 25 27 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.72 $Y=1.21
+ $X2=3.72 $Y2=0.655
r146 21 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.295
+ $X2=1.57 $Y2=1.46
r147 21 23 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.57 $Y=1.295
+ $X2=1.57 $Y2=0.655
r148 17 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.565 $Y=1.625
+ $X2=1.565 $Y2=1.46
r149 17 19 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.565 $Y=1.625
+ $X2=1.565 $Y2=2.465
r150 13 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.295
+ $X2=1.14 $Y2=1.46
r151 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.14 $Y=1.295
+ $X2=1.14 $Y2=0.655
r152 9 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.625
+ $X2=1.135 $Y2=1.46
r153 9 11 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.135 $Y=1.625
+ $X2=1.135 $Y2=2.465
r154 5 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.71 $Y=1.295
+ $X2=0.71 $Y2=1.46
r155 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.71 $Y=1.295 $X2=0.71
+ $Y2=0.655
r156 1 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.705 $Y=1.625
+ $X2=0.705 $Y2=1.46
r157 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.705 $Y=1.625
+ $X2=0.705 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%B2 3 7 11 15 19 23 27 31 33 34 35 54 55 57
+ 69
c81 54 0 8.05408e-21 $X=3.17 $Y=1.4
c82 27 0 3.60491e-20 $X=3.285 $Y=2.465
r83 57 69 1.13539 $w=2.85e-07 $l=2.2e-08 $layer=LI1_cond $X=2.182 $Y=1.342
+ $X2=2.16 $Y2=1.342
r84 55 56 0.732523 $w=3.29e-07 $l=5e-09 $layer=POLY_cond $X=3.285 $Y=1.4
+ $X2=3.29 $Y2=1.4
r85 53 55 16.848 $w=3.29e-07 $l=1.15e-07 $layer=POLY_cond $X=3.17 $Y=1.4
+ $X2=3.285 $Y2=1.4
r86 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.4 $X2=3.17 $Y2=1.4
r87 51 53 45.4164 $w=3.29e-07 $l=3.1e-07 $layer=POLY_cond $X=2.86 $Y=1.4
+ $X2=3.17 $Y2=1.4
r88 50 51 0.732523 $w=3.29e-07 $l=5e-09 $layer=POLY_cond $X=2.855 $Y=1.4
+ $X2=2.86 $Y2=1.4
r89 48 50 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=2.83 $Y=1.4
+ $X2=2.855 $Y2=1.4
r90 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.83 $Y=1.4
+ $X2=2.83 $Y2=1.4
r91 46 48 58.6018 $w=3.29e-07 $l=4e-07 $layer=POLY_cond $X=2.43 $Y=1.4 $X2=2.83
+ $Y2=1.4
r92 45 46 0.732523 $w=3.29e-07 $l=5e-09 $layer=POLY_cond $X=2.425 $Y=1.4
+ $X2=2.43 $Y2=1.4
r93 44 69 0.484127 $w=2.52e-07 $l=1e-08 $layer=LI1_cond $X=2.15 $Y=1.342
+ $X2=2.16 $Y2=1.342
r94 43 45 40.2888 $w=3.29e-07 $l=2.75e-07 $layer=POLY_cond $X=2.15 $Y=1.4
+ $X2=2.425 $Y2=1.4
r95 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.4 $X2=2.15 $Y2=1.4
r96 41 43 21.9757 $w=3.29e-07 $l=1.5e-07 $layer=POLY_cond $X=2 $Y=1.4 $X2=2.15
+ $Y2=1.4
r97 40 41 0.732523 $w=3.29e-07 $l=5e-09 $layer=POLY_cond $X=1.995 $Y=1.4 $X2=2
+ $Y2=1.4
r98 35 54 2.02183 $w=2.83e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=1.342 $X2=3.17
+ $Y2=1.342
r99 35 49 11.7266 $w=2.83e-07 $l=2.9e-07 $layer=LI1_cond $X=3.12 $Y=1.342
+ $X2=2.83 $Y2=1.342
r100 34 49 7.68295 $w=2.83e-07 $l=1.9e-07 $layer=LI1_cond $X=2.64 $Y=1.342
+ $X2=2.83 $Y2=1.342
r101 33 44 1.06508 $w=2.52e-07 $l=2.2e-08 $layer=LI1_cond $X=2.128 $Y=1.342
+ $X2=2.15 $Y2=1.342
r102 33 34 17.2664 $w=2.83e-07 $l=4.27e-07 $layer=LI1_cond $X=2.213 $Y=1.342
+ $X2=2.64 $Y2=1.342
r103 33 57 1.25353 $w=2.83e-07 $l=3.1e-08 $layer=LI1_cond $X=2.213 $Y=1.342
+ $X2=2.182 $Y2=1.342
r104 29 56 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.29 $Y=1.235
+ $X2=3.29 $Y2=1.4
r105 29 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.29 $Y=1.235
+ $X2=3.29 $Y2=0.655
r106 25 55 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.565
+ $X2=3.285 $Y2=1.4
r107 25 27 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=3.285 $Y=1.565
+ $X2=3.285 $Y2=2.465
r108 21 51 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.86 $Y=1.235
+ $X2=2.86 $Y2=1.4
r109 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.86 $Y=1.235
+ $X2=2.86 $Y2=0.655
r110 17 50 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.565
+ $X2=2.855 $Y2=1.4
r111 17 19 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.855 $Y=1.565
+ $X2=2.855 $Y2=2.465
r112 13 46 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=1.235
+ $X2=2.43 $Y2=1.4
r113 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.43 $Y=1.235
+ $X2=2.43 $Y2=0.655
r114 9 45 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.425 $Y=1.565
+ $X2=2.425 $Y2=1.4
r115 9 11 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.425 $Y=1.565
+ $X2=2.425 $Y2=2.465
r116 5 41 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2 $Y=1.235 $X2=2
+ $Y2=1.4
r117 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2 $Y=1.235 $X2=2
+ $Y2=0.655
r118 1 40 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.995 $Y=1.565
+ $X2=1.995 $Y2=1.4
r119 1 3 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.995 $Y=1.565
+ $X2=1.995 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%A_832_21# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 56 59 62 64 65 68 70 72 76 80 82 84 85 88 92 94 96 99 103 104 108 109 113
+ 114 118 129
c193 129 0 2.77078e-19 $X=5.595 $Y=1.49
r194 128 129 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.525 $Y=1.49
+ $X2=5.595 $Y2=1.49
r195 127 128 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=5.165 $Y=1.49
+ $X2=5.525 $Y2=1.49
r196 126 127 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.095 $Y=1.49
+ $X2=5.165 $Y2=1.49
r197 123 124 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.665 $Y=1.49
+ $X2=4.735 $Y2=1.49
r198 119 121 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.235 $Y=1.49
+ $X2=4.305 $Y2=1.49
r199 114 116 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=9.265 $Y=0.955
+ $X2=9.265 $Y2=1.09
r200 114 115 4.75232 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=0.955
+ $X2=9.265 $Y2=0.87
r201 105 107 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.965 $Y=1.15
+ $X2=6.17 $Y2=1.15
r202 102 126 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.02 $Y=1.49
+ $X2=5.095 $Y2=1.49
r203 102 124 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=5.02 $Y=1.49
+ $X2=4.735 $Y2=1.49
r204 101 104 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=5.02 $Y=1.552
+ $X2=5.185 $Y2=1.552
r205 101 103 2.7521 $w=3.33e-07 $l=8e-08 $layer=LI1_cond $X=5.02 $Y=1.552
+ $X2=4.94 $Y2=1.552
r206 101 102 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.02
+ $Y=1.49 $X2=5.02 $Y2=1.49
r207 98 99 28.133 $w=2.03e-07 $l=5.2e-07 $layer=LI1_cond $X=9.832 $Y=1.175
+ $X2=9.832 $Y2=1.695
r208 97 118 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=9.475 $Y=1.785
+ $X2=9.345 $Y2=1.785
r209 96 99 6.85394 $w=1.8e-07 $l=1.39943e-07 $layer=LI1_cond $X=9.73 $Y=1.785
+ $X2=9.832 $Y2=1.695
r210 96 97 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=9.73 $Y=1.785
+ $X2=9.475 $Y2=1.785
r211 95 116 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=9.365 $Y=1.09
+ $X2=9.265 $Y2=1.09
r212 94 98 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=9.73 $Y=1.09
+ $X2=9.832 $Y2=1.175
r213 94 95 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.73 $Y=1.09
+ $X2=9.365 $Y2=1.09
r214 90 118 0.0585112 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=9.345 $Y=1.875
+ $X2=9.345 $Y2=1.785
r215 90 92 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=9.345 $Y=1.875
+ $X2=9.345 $Y2=1.98
r216 88 115 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=9.27 $Y=0.42
+ $X2=9.27 $Y2=0.87
r217 84 118 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=9.215 $Y=1.785
+ $X2=9.345 $Y2=1.785
r218 84 85 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=9.215 $Y=1.785
+ $X2=8.615 $Y2=1.785
r219 83 113 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=8.505 $Y=0.955
+ $X2=8.405 $Y2=0.955
r220 82 114 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=9.165 $Y=0.955
+ $X2=9.265 $Y2=0.955
r221 82 83 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=9.165 $Y=0.955
+ $X2=8.505 $Y2=0.955
r222 78 85 7.21025 $w=1.8e-07 $l=1.77381e-07 $layer=LI1_cond $X=8.477 $Y=1.875
+ $X2=8.615 $Y2=1.785
r223 78 80 4.40024 $w=2.73e-07 $l=1.05e-07 $layer=LI1_cond $X=8.477 $Y=1.875
+ $X2=8.477 $Y2=1.98
r224 74 113 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=0.87
+ $X2=8.405 $Y2=0.955
r225 74 76 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=8.405 $Y=0.87
+ $X2=8.405 $Y2=0.42
r226 73 109 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=0.955
+ $X2=7.955 $Y2=0.955
r227 72 113 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=8.305 $Y=0.955
+ $X2=8.405 $Y2=0.955
r228 72 73 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.305 $Y=0.955
+ $X2=8.04 $Y2=0.955
r229 71 108 5.34142 $w=1.82e-07 $l=9.5e-08 $layer=LI1_cond $X=7.125 $Y=1.137
+ $X2=7.03 $Y2=1.137
r230 70 109 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=7.955 $Y=1.137
+ $X2=7.955 $Y2=0.955
r231 70 71 42.373 $w=1.93e-07 $l=7.45e-07 $layer=LI1_cond $X=7.87 $Y=1.137
+ $X2=7.125 $Y2=1.137
r232 66 108 1.19794 $w=1.9e-07 $l=9.7e-08 $layer=LI1_cond $X=7.03 $Y=1.04
+ $X2=7.03 $Y2=1.137
r233 66 68 36.1914 $w=1.88e-07 $l=6.2e-07 $layer=LI1_cond $X=7.03 $Y=1.04
+ $X2=7.03 $Y2=0.42
r234 65 107 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.265 $Y=1.15
+ $X2=6.17 $Y2=1.15
r235 64 108 5.34142 $w=1.82e-07 $l=1.01292e-07 $layer=LI1_cond $X=6.935 $Y=1.15
+ $X2=7.03 $Y2=1.137
r236 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.935 $Y=1.15
+ $X2=6.265 $Y2=1.15
r237 60 107 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.17 $Y=1.065
+ $X2=6.17 $Y2=1.15
r238 60 62 27.7273 $w=1.88e-07 $l=4.75e-07 $layer=LI1_cond $X=6.17 $Y=1.065
+ $X2=6.17 $Y2=0.59
r239 58 105 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=1.235
+ $X2=5.965 $Y2=1.15
r240 58 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.965 $Y=1.235
+ $X2=5.965 $Y2=1.55
r241 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.88 $Y=1.635
+ $X2=5.965 $Y2=1.55
r242 56 104 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.88 $Y=1.635
+ $X2=5.185 $Y2=1.635
r243 54 123 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.5 $Y=1.49
+ $X2=4.665 $Y2=1.49
r244 54 121 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.5 $Y=1.49
+ $X2=4.305 $Y2=1.49
r245 53 103 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.5 $Y=1.55
+ $X2=4.94 $Y2=1.55
r246 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.5
+ $Y=1.49 $X2=4.5 $Y2=1.49
r247 47 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.595 $Y=1.655
+ $X2=5.595 $Y2=1.49
r248 47 49 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.595 $Y=1.655
+ $X2=5.595 $Y2=2.465
r249 43 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.525 $Y=1.325
+ $X2=5.525 $Y2=1.49
r250 43 45 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.525 $Y=1.325
+ $X2=5.525 $Y2=0.655
r251 39 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.165 $Y=1.655
+ $X2=5.165 $Y2=1.49
r252 39 41 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.165 $Y=1.655
+ $X2=5.165 $Y2=2.465
r253 35 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.095 $Y=1.325
+ $X2=5.095 $Y2=1.49
r254 35 37 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.095 $Y=1.325
+ $X2=5.095 $Y2=0.655
r255 31 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=1.655
+ $X2=4.735 $Y2=1.49
r256 31 33 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.735 $Y=1.655
+ $X2=4.735 $Y2=2.465
r257 27 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.665 $Y=1.325
+ $X2=4.665 $Y2=1.49
r258 27 29 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=4.665 $Y=1.325
+ $X2=4.665 $Y2=0.655
r259 23 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.655
+ $X2=4.305 $Y2=1.49
r260 23 25 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.305 $Y=1.655
+ $X2=4.305 $Y2=2.465
r261 19 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.325
+ $X2=4.235 $Y2=1.49
r262 19 21 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=4.235 $Y=1.325
+ $X2=4.235 $Y2=0.655
r263 6 92 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.2
+ $Y=1.835 $X2=9.34 $Y2=1.98
r264 5 80 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.34
+ $Y=1.835 $X2=8.48 $Y2=1.98
r265 4 88 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.13
+ $Y=0.235 $X2=9.27 $Y2=0.42
r266 3 76 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.27
+ $Y=0.235 $X2=8.41 $Y2=0.42
r267 2 68 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.89
+ $Y=0.235 $X2=7.03 $Y2=0.42
r268 1 62 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=6.03
+ $Y=0.235 $X2=6.17 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%A1_N 3 7 11 15 19 23 27 31 33 34 35 36 59
c93 36 0 8.22749e-20 $X=7.92 $Y=1.665
r94 57 59 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.745 $Y=1.51
+ $X2=7.835 $Y2=1.51
r95 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.745
+ $Y=1.51 $X2=7.745 $Y2=1.51
r96 54 57 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.405 $Y=1.51
+ $X2=7.745 $Y2=1.51
r97 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.405
+ $Y=1.51 $X2=7.405 $Y2=1.51
r98 52 54 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=7.245 $Y=1.51
+ $X2=7.405 $Y2=1.51
r99 51 52 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=6.975 $Y=1.51
+ $X2=7.245 $Y2=1.51
r100 50 51 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.815 $Y=1.51
+ $X2=6.975 $Y2=1.51
r101 48 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.725 $Y=1.51
+ $X2=6.815 $Y2=1.51
r102 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.725
+ $Y=1.51 $X2=6.725 $Y2=1.51
r103 46 48 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=6.545 $Y=1.51
+ $X2=6.725 $Y2=1.51
r104 44 46 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.385 $Y=1.51
+ $X2=6.545 $Y2=1.51
r105 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.385
+ $Y=1.51 $X2=6.385 $Y2=1.51
r106 41 44 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.955 $Y=1.51
+ $X2=6.385 $Y2=1.51
r107 36 58 5.76222 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=7.92 $Y=1.58
+ $X2=7.745 $Y2=1.58
r108 35 58 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=7.44 $Y=1.58
+ $X2=7.745 $Y2=1.58
r109 35 55 1.15244 $w=3.48e-07 $l=3.5e-08 $layer=LI1_cond $X=7.44 $Y=1.58
+ $X2=7.405 $Y2=1.58
r110 34 55 14.6525 $w=3.48e-07 $l=4.45e-07 $layer=LI1_cond $X=6.96 $Y=1.58
+ $X2=7.405 $Y2=1.58
r111 34 49 7.73783 $w=3.48e-07 $l=2.35e-07 $layer=LI1_cond $X=6.96 $Y=1.58
+ $X2=6.725 $Y2=1.58
r112 33 49 8.0671 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=6.48 $Y=1.58
+ $X2=6.725 $Y2=1.58
r113 33 45 3.12806 $w=3.48e-07 $l=9.5e-08 $layer=LI1_cond $X=6.48 $Y=1.58
+ $X2=6.385 $Y2=1.58
r114 29 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.835 $Y=1.675
+ $X2=7.835 $Y2=1.51
r115 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.835 $Y=1.675
+ $X2=7.835 $Y2=2.465
r116 25 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.405 $Y=1.675
+ $X2=7.405 $Y2=1.51
r117 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.405 $Y=1.675
+ $X2=7.405 $Y2=2.465
r118 21 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.245 $Y=1.345
+ $X2=7.245 $Y2=1.51
r119 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.245 $Y=1.345
+ $X2=7.245 $Y2=0.655
r120 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.975 $Y=1.675
+ $X2=6.975 $Y2=1.51
r121 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.975 $Y=1.675
+ $X2=6.975 $Y2=2.465
r122 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.815 $Y=1.345
+ $X2=6.815 $Y2=1.51
r123 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.815 $Y=1.345
+ $X2=6.815 $Y2=0.655
r124 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.545 $Y=1.675
+ $X2=6.545 $Y2=1.51
r125 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.545 $Y=1.675
+ $X2=6.545 $Y2=2.465
r126 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.385 $Y=1.345
+ $X2=6.385 $Y2=1.51
r127 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.385 $Y=1.345
+ $X2=6.385 $Y2=0.655
r128 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.345
+ $X2=5.955 $Y2=1.51
r129 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.955 $Y=1.345
+ $X2=5.955 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%A2_N 3 7 11 15 19 23 27 31 33 34 54 56 58
+ 70
r83 58 70 2.63416 $w=3.13e-07 $l=7.2e-08 $layer=LI1_cond $X=8.808 $Y=1.367
+ $X2=8.88 $Y2=1.367
r84 55 56 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=9.485 $Y=1.44
+ $X2=9.555 $Y2=1.44
r85 53 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.395 $Y=1.44
+ $X2=9.485 $Y2=1.44
r86 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.395
+ $Y=1.44 $X2=9.395 $Y2=1.44
r87 51 53 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=9.125 $Y=1.44
+ $X2=9.395 $Y2=1.44
r88 50 51 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=9.055 $Y=1.44
+ $X2=9.125 $Y2=1.44
r89 48 50 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.715 $Y=1.44
+ $X2=9.055 $Y2=1.44
r90 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.715
+ $Y=1.44 $X2=8.715 $Y2=1.44
r91 46 48 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=8.695 $Y=1.44
+ $X2=8.715 $Y2=1.44
r92 45 46 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.625 $Y=1.44
+ $X2=8.695 $Y2=1.44
r93 43 45 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=8.375 $Y=1.44
+ $X2=8.625 $Y2=1.44
r94 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.375
+ $Y=1.44 $X2=8.375 $Y2=1.44
r95 41 43 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.265 $Y=1.44
+ $X2=8.375 $Y2=1.44
r96 39 41 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.195 $Y=1.44
+ $X2=8.265 $Y2=1.44
r97 34 70 0.219513 $w=3.13e-07 $l=6e-09 $layer=LI1_cond $X=8.886 $Y=1.367
+ $X2=8.88 $Y2=1.367
r98 34 54 23.3881 $w=2.13e-07 $l=4.3e-07 $layer=LI1_cond $X=8.965 $Y=1.435
+ $X2=9.395 $Y2=1.435
r99 34 58 0.256098 $w=3.13e-07 $l=7e-09 $layer=LI1_cond $X=8.801 $Y=1.367
+ $X2=8.808 $Y2=1.367
r100 34 49 3.14635 $w=3.13e-07 $l=8.6e-08 $layer=LI1_cond $X=8.801 $Y=1.367
+ $X2=8.715 $Y2=1.367
r101 33 49 11.5244 $w=3.13e-07 $l=3.15e-07 $layer=LI1_cond $X=8.4 $Y=1.367
+ $X2=8.715 $Y2=1.367
r102 33 44 0.914637 $w=3.13e-07 $l=2.5e-08 $layer=LI1_cond $X=8.4 $Y=1.367
+ $X2=8.375 $Y2=1.367
r103 29 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.555 $Y=1.605
+ $X2=9.555 $Y2=1.44
r104 29 31 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=9.555 $Y=1.605
+ $X2=9.555 $Y2=2.465
r105 25 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.485 $Y=1.275
+ $X2=9.485 $Y2=1.44
r106 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=9.485 $Y=1.275
+ $X2=9.485 $Y2=0.655
r107 21 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.125 $Y=1.605
+ $X2=9.125 $Y2=1.44
r108 21 23 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=9.125 $Y=1.605
+ $X2=9.125 $Y2=2.465
r109 17 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.055 $Y=1.275
+ $X2=9.055 $Y2=1.44
r110 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=9.055 $Y=1.275
+ $X2=9.055 $Y2=0.655
r111 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.695 $Y=1.605
+ $X2=8.695 $Y2=1.44
r112 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.695 $Y=1.605
+ $X2=8.695 $Y2=2.465
r113 9 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.625 $Y=1.275
+ $X2=8.625 $Y2=1.44
r114 9 11 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.625 $Y=1.275
+ $X2=8.625 $Y2=0.655
r115 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.265 $Y=1.605
+ $X2=8.265 $Y2=1.44
r116 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.265 $Y=1.605
+ $X2=8.265 $Y2=2.465
r117 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.195 $Y=1.275
+ $X2=8.195 $Y2=1.44
r118 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.195 $Y=1.275
+ $X2=8.195 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%A_73_367# 1 2 3 4 5 6 7 24 28 29 32 34 38
+ 40 44 46 48 49 50 51 54 56 58 60 62 69 71 74
c90 48 0 3.60491e-20 $X=4.05 $Y=2.425
r91 66 67 4.61288 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=2.1 $X2=1.36
+ $Y2=2.185
r92 65 66 6.33766 $w=2.08e-07 $l=1.2e-07 $layer=LI1_cond $X=1.36 $Y=1.98
+ $X2=1.36 $Y2=2.1
r93 62 65 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=1.36 $Y=1.81
+ $X2=1.36 $Y2=1.98
r94 58 76 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=2.905
+ $X2=5.845 $Y2=2.99
r95 58 60 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=5.845 $Y=2.905
+ $X2=5.845 $Y2=2.055
r96 57 74 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.045 $Y=2.99
+ $X2=4.95 $Y2=2.99
r97 56 76 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.715 $Y=2.99
+ $X2=5.845 $Y2=2.99
r98 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.715 $Y=2.99
+ $X2=5.045 $Y2=2.99
r99 52 74 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=2.905
+ $X2=4.95 $Y2=2.99
r100 52 54 28.311 $w=1.88e-07 $l=4.85e-07 $layer=LI1_cond $X=4.95 $Y=2.905
+ $X2=4.95 $Y2=2.42
r101 50 74 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.855 $Y=2.99
+ $X2=4.95 $Y2=2.99
r102 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.855 $Y=2.99
+ $X2=4.185 $Y2=2.99
r103 49 51 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.05 $Y=2.905
+ $X2=4.185 $Y2=2.99
r104 48 49 20.4879 $w=2.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.05 $Y=2.425
+ $X2=4.05 $Y2=2.905
r105 47 71 3.81196 $w=2.85e-07 $l=1e-07 $layer=LI1_cond $X=3.175 $Y=2.215
+ $X2=3.075 $Y2=2.215
r106 46 48 18.2784 $w=4e-07 $l=6.31328e-07 $layer=LI1_cond $X=3.515 $Y=2.215
+ $X2=4.05 $Y2=2.425
r107 46 47 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=3.515 $Y=2.215
+ $X2=3.175 $Y2=2.215
r108 42 71 2.64391 $w=2e-07 $l=2e-07 $layer=LI1_cond $X=3.075 $Y=2.415 $X2=3.075
+ $Y2=2.215
r109 42 44 7.20909 $w=1.98e-07 $l=1.3e-07 $layer=LI1_cond $X=3.075 $Y=2.415
+ $X2=3.075 $Y2=2.545
r110 41 69 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.305 $Y=2.1
+ $X2=2.21 $Y2=2.1
r111 40 71 3.81196 $w=2.85e-07 $l=1.57242e-07 $layer=LI1_cond $X=2.975 $Y=2.1
+ $X2=3.075 $Y2=2.215
r112 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.975 $Y=2.1
+ $X2=2.305 $Y2=2.1
r113 36 69 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=2.185
+ $X2=2.21 $Y2=2.1
r114 36 38 42.3206 $w=1.88e-07 $l=7.25e-07 $layer=LI1_cond $X=2.21 $Y=2.185
+ $X2=2.21 $Y2=2.91
r115 35 66 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.465 $Y=2.1
+ $X2=1.36 $Y2=2.1
r116 34 69 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.115 $Y=2.1
+ $X2=2.21 $Y2=2.1
r117 34 35 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.115 $Y=2.1
+ $X2=1.465 $Y2=2.1
r118 32 67 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=1.35 $Y=2.44
+ $X2=1.35 $Y2=2.185
r119 28 62 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.255 $Y=1.81
+ $X2=1.36 $Y2=1.81
r120 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.255 $Y=1.81
+ $X2=0.585 $Y2=1.81
r121 24 26 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.455 $Y=1.98
+ $X2=0.455 $Y2=2.91
r122 22 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.455 $Y=1.895
+ $X2=0.585 $Y2=1.81
r123 22 24 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.455 $Y=1.895
+ $X2=0.455 $Y2=1.98
r124 7 76 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.67
+ $Y=1.835 $X2=5.81 $Y2=2.91
r125 7 60 400 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=5.67
+ $Y=1.835 $X2=5.81 $Y2=2.055
r126 6 54 300 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_PDIFF $count=2 $X=4.81
+ $Y=1.835 $X2=4.95 $Y2=2.42
r127 5 48 300 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_PDIFF $count=2 $X=3.95
+ $Y=1.835 $X2=4.09 $Y2=2.42
r128 4 71 600 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.835 $X2=3.07 $Y2=2.18
r129 4 44 300 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=2 $X=2.93
+ $Y=1.835 $X2=3.07 $Y2=2.545
r130 3 69 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=2.07
+ $Y=1.835 $X2=2.21 $Y2=2.18
r131 3 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.07
+ $Y=1.835 $X2=2.21 $Y2=2.91
r132 2 65 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.21
+ $Y=1.835 $X2=1.35 $Y2=1.98
r133 2 32 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=1.21
+ $Y=1.835 $X2=1.35 $Y2=2.44
r134 1 26 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.365
+ $Y=1.835 $X2=0.49 $Y2=2.91
r135 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.365
+ $Y=1.835 $X2=0.49 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 45 47
+ 48 50 51 53 54 55 61 66 85 86 89 92 95
r145 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r146 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r147 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r148 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r149 83 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=9.84 $Y2=3.33
r150 82 85 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=9.84 $Y2=3.33
r151 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r152 80 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r153 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r155 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r156 74 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r157 73 76 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=6.48 $Y2=3.33
r158 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r159 71 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.58 $Y2=3.33
r160 71 73 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=4.08 $Y2=3.33
r161 70 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r162 70 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r163 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r164 67 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.64 $Y2=3.33
r165 67 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=3.12 $Y2=3.33
r166 66 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.58 $Y2=3.33
r167 66 69 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.12 $Y2=3.33
r168 65 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r169 65 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r170 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r171 62 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=1.78 $Y2=3.33
r172 62 64 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=2.16 $Y2=3.33
r173 61 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.64 $Y2=3.33
r174 61 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=3.33
+ $X2=2.16 $Y2=3.33
r175 59 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r176 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r177 55 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r178 55 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r179 53 79 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.455 $Y=3.33
+ $X2=7.44 $Y2=3.33
r180 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=3.33
+ $X2=7.62 $Y2=3.33
r181 52 82 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.785 $Y=3.33
+ $X2=7.92 $Y2=3.33
r182 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.785 $Y=3.33
+ $X2=7.62 $Y2=3.33
r183 50 76 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.48 $Y2=3.33
r184 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.76 $Y2=3.33
r185 49 79 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.925 $Y=3.33
+ $X2=7.44 $Y2=3.33
r186 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.925 $Y=3.33
+ $X2=6.76 $Y2=3.33
r187 47 58 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.72 $Y2=3.33
r188 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.92 $Y2=3.33
r189 43 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.62 $Y=3.245
+ $X2=7.62 $Y2=3.33
r190 43 45 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.62 $Y=3.245
+ $X2=7.62 $Y2=2.375
r191 39 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=3.245
+ $X2=6.76 $Y2=3.33
r192 39 41 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.76 $Y=3.245
+ $X2=6.76 $Y2=2.375
r193 35 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.58 $Y2=3.33
r194 35 37 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.58 $Y2=2.67
r195 31 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=3.245
+ $X2=2.64 $Y2=3.33
r196 31 33 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=2.64 $Y=3.245
+ $X2=2.64 $Y2=2.44
r197 27 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=3.245
+ $X2=1.78 $Y2=3.33
r198 27 29 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=1.78 $Y=3.245
+ $X2=1.78 $Y2=2.44
r199 26 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.92 $Y2=3.33
r200 25 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=1.78 $Y2=3.33
r201 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=1.085 $Y2=3.33
r202 21 24 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=0.92 $Y=2.15 $X2=0.92
+ $Y2=2.95
r203 19 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=3.33
r204 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=2.95
r205 6 45 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=7.48
+ $Y=1.835 $X2=7.62 $Y2=2.375
r206 5 41 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=6.62
+ $Y=1.835 $X2=6.76 $Y2=2.375
r207 4 37 300 $w=1.7e-07 $l=9.38576e-07 $layer=licon1_PDIFF $count=2 $X=3.36
+ $Y=1.835 $X2=3.58 $Y2=2.67
r208 3 33 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=2.5
+ $Y=1.835 $X2=2.64 $Y2=2.44
r209 2 29 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=1.64
+ $Y=1.835 $X2=1.78 $Y2=2.44
r210 1 24 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.78
+ $Y=1.835 $X2=0.92 $Y2=2.95
r211 1 21 400 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_PDIFF $count=1 $X=0.78
+ $Y=1.835 $X2=0.92 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%Y 1 2 3 4 5 6 19 26 29 33 35 36 37 41 51
+ 53 54
r96 54 56 8.92683 $w=2.87e-07 $l=2.1e-07 $layer=LI1_cond $X=5.52 $Y=1.212
+ $X2=5.31 $Y2=1.212
r97 50 51 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=4.52 $Y=1.985
+ $X2=4.77 $Y2=1.985
r98 47 50 24.4 $w=1.98e-07 $l=4.4e-07 $layer=LI1_cond $X=4.08 $Y=1.985 $X2=4.52
+ $Y2=1.985
r99 39 56 3.15132 $w=1.9e-07 $l=1.67e-07 $layer=LI1_cond $X=5.31 $Y=1.045
+ $X2=5.31 $Y2=1.212
r100 39 41 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=5.31 $Y=1.045
+ $X2=5.31 $Y2=0.42
r101 37 53 4.65494 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=5.215 $Y=1.987
+ $X2=5.38 $Y2=1.987
r102 37 51 25.31 $w=1.93e-07 $l=4.45e-07 $layer=LI1_cond $X=5.215 $Y=1.987
+ $X2=4.77 $Y2=1.987
r103 36 46 7.2949 $w=3.42e-07 $l=1.95282e-07 $layer=LI1_cond $X=4.545 $Y=1.13
+ $X2=4.427 $Y2=0.985
r104 35 56 6.04938 $w=2.87e-07 $l=1.29673e-07 $layer=LI1_cond $X=5.215 $Y=1.13
+ $X2=5.31 $Y2=1.212
r105 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.215 $Y=1.13
+ $X2=4.545 $Y2=1.13
r106 33 50 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=4.52 $Y=2.65
+ $X2=4.52 $Y2=2.085
r107 27 46 2.95219 $w=2.35e-07 $l=2.3e-07 $layer=LI1_cond $X=4.427 $Y=0.755
+ $X2=4.427 $Y2=0.985
r108 27 29 16.4284 $w=2.33e-07 $l=3.35e-07 $layer=LI1_cond $X=4.427 $Y=0.755
+ $X2=4.427 $Y2=0.42
r109 26 47 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.08 $Y=1.885 $X2=4.08
+ $Y2=1.985
r110 25 46 12.3784 $w=3.42e-07 $l=3.47e-07 $layer=LI1_cond $X=4.08 $Y=0.985
+ $X2=4.427 $Y2=0.985
r111 25 26 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.08 $Y=1.03
+ $X2=4.08 $Y2=1.885
r112 21 24 36.04 $w=2.73e-07 $l=8.6e-07 $layer=LI1_cond $X=2.215 $Y=0.892
+ $X2=3.075 $Y2=0.892
r113 19 25 3.53581 $w=3.42e-07 $l=1.28662e-07 $layer=LI1_cond $X=3.995 $Y=0.892
+ $X2=4.08 $Y2=0.985
r114 19 24 38.5545 $w=2.73e-07 $l=9.2e-07 $layer=LI1_cond $X=3.995 $Y=0.892
+ $X2=3.075 $Y2=0.892
r115 6 53 300 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=2 $X=5.24
+ $Y=1.835 $X2=5.38 $Y2=2.055
r116 5 50 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.835 $X2=4.52 $Y2=1.97
r117 5 33 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.835 $X2=4.52 $Y2=2.65
r118 4 41 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.17
+ $Y=0.235 $X2=5.31 $Y2=0.42
r119 3 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.31
+ $Y=0.235 $X2=4.45 $Y2=0.42
r120 2 24 182 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_NDIFF $count=1 $X=2.935
+ $Y=0.235 $X2=3.075 $Y2=0.89
r121 1 21 182 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.235 $X2=2.215 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%A_1241_367# 1 2 3 4 5 16 18 20 24 26 28 29
+ 30 34 36 38 40 45 51
r56 38 53 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.79 $Y=2.905
+ $X2=9.79 $Y2=2.99
r57 38 40 27.6189 $w=2.88e-07 $l=6.95e-07 $layer=LI1_cond $X=9.79 $Y=2.905
+ $X2=9.79 $Y2=2.21
r58 37 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.045 $Y=2.99
+ $X2=8.915 $Y2=2.99
r59 36 53 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.645 $Y=2.99
+ $X2=9.79 $Y2=2.99
r60 36 37 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=9.645 $Y=2.99
+ $X2=9.045 $Y2=2.99
r61 32 51 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.915 $Y=2.905
+ $X2=8.915 $Y2=2.99
r62 32 34 30.8057 $w=2.58e-07 $l=6.95e-07 $layer=LI1_cond $X=8.915 $Y=2.905
+ $X2=8.915 $Y2=2.21
r63 31 49 3.88258 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=8.17 $Y=2.99
+ $X2=8.062 $Y2=2.99
r64 30 51 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.785 $Y=2.99
+ $X2=8.915 $Y2=2.99
r65 30 31 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=8.785 $Y=2.99
+ $X2=8.17 $Y2=2.99
r66 29 49 3.05574 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=8.062 $Y=2.905
+ $X2=8.062 $Y2=2.99
r67 28 47 3.07165 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=8.062 $Y=2.1
+ $X2=8.062 $Y2=2.015
r68 28 29 43.1496 $w=2.13e-07 $l=8.05e-07 $layer=LI1_cond $X=8.062 $Y=2.1
+ $X2=8.062 $Y2=2.905
r69 27 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.285 $Y=2.015
+ $X2=7.19 $Y2=2.015
r70 26 47 3.86667 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=7.955 $Y=2.015
+ $X2=8.062 $Y2=2.015
r71 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.955 $Y=2.015
+ $X2=7.285 $Y2=2.015
r72 22 45 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.19 $Y=2.1 $X2=7.19
+ $Y2=2.015
r73 22 24 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=7.19 $Y=2.1 $X2=7.19
+ $Y2=2.91
r74 21 43 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.425 $Y=2.015
+ $X2=6.295 $Y2=2.015
r75 20 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.095 $Y=2.015
+ $X2=7.19 $Y2=2.015
r76 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.095 $Y=2.015
+ $X2=6.425 $Y2=2.015
r77 16 43 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=2.1
+ $X2=6.295 $Y2=2.015
r78 16 18 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=6.295 $Y=2.1
+ $X2=6.295 $Y2=2.91
r79 5 53 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.63
+ $Y=1.835 $X2=9.77 $Y2=2.91
r80 5 40 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=9.63
+ $Y=1.835 $X2=9.77 $Y2=2.21
r81 4 51 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.835 $X2=8.91 $Y2=2.91
r82 4 34 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=8.77
+ $Y=1.835 $X2=8.91 $Y2=2.21
r83 3 49 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.91
+ $Y=1.835 $X2=8.05 $Y2=2.91
r84 3 47 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=7.91
+ $Y=1.835 $X2=8.05 $Y2=2.095
r85 2 45 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=7.05
+ $Y=1.835 $X2=7.19 $Y2=2.095
r86 2 24 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.05
+ $Y=1.835 $X2=7.19 $Y2=2.91
r87 1 43 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.835 $X2=6.33 $Y2=2.095
r88 1 18 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.835 $X2=6.33 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%VGND 1 2 3 4 5 6 7 8 9 30 32 36 40 44 48
+ 50 54 58 60 62 64 65 67 68 70 71 72 73 74 93 98 103 109 112 120 124 128
c159 48 0 1.94803e-19 $X=5.74 $Y=0.36
r160 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r161 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r162 120 122 6.92256 $w=7.49e-07 $l=5.37587e-07 $layer=LI1_cond $X=7.715 $Y=0.36
+ $X2=7.46 $Y2=0.785
r163 116 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r164 115 120 5.86382 $w=7.49e-07 $l=3.6e-07 $layer=LI1_cond $X=7.715 $Y=0
+ $X2=7.715 $Y2=0.36
r165 115 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r166 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r167 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r168 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r169 107 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r170 107 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r171 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r172 104 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.005 $Y=0
+ $X2=8.84 $Y2=0
r173 104 106 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.005 $Y=0
+ $X2=9.36 $Y2=0
r174 103 127 4.55259 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.807 $Y2=0
r175 103 106 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.36 $Y2=0
r176 102 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r177 102 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=7.92 $Y2=0
r178 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r179 99 115 9.76921 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=8.135 $Y=0
+ $X2=7.715 $Y2=0
r180 99 101 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.135 $Y=0
+ $X2=8.4 $Y2=0
r181 98 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.675 $Y=0
+ $X2=8.84 $Y2=0
r182 98 101 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=0
+ $X2=8.4 $Y2=0
r183 97 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r184 97 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r185 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r186 94 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=0 $X2=6.6
+ $Y2=0
r187 94 96 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.765 $Y=0
+ $X2=6.96 $Y2=0
r188 93 115 9.76921 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=7.295 $Y=0
+ $X2=7.715 $Y2=0
r189 93 96 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.295 $Y=0
+ $X2=6.96 $Y2=0
r190 92 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.48 $Y2=0
r191 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r192 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r193 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r194 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r195 83 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r196 83 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r197 82 85 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r198 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r199 80 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=0
+ $X2=1.355 $Y2=0
r200 80 82 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.68
+ $Y2=0
r201 78 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r202 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r203 74 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r204 74 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r205 72 91 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.575 $Y=0 $X2=5.52
+ $Y2=0
r206 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.575 $Y=0 $X2=5.74
+ $Y2=0
r207 70 88 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=4.56 $Y2=0
r208 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.88
+ $Y2=0
r209 69 91 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=5.52 $Y2=0
r210 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=0 $X2=4.88
+ $Y2=0
r211 67 85 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.6
+ $Y2=0
r212 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.975
+ $Y2=0
r213 66 88 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.56
+ $Y2=0
r214 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=3.975
+ $Y2=0
r215 64 77 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.33 $Y=0 $X2=0.24
+ $Y2=0
r216 64 65 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.33 $Y=0 $X2=0.475
+ $Y2=0
r217 60 127 3.21359 $w=3.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=9.7 $Y=0.085
+ $X2=9.807 $Y2=0
r218 60 62 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.7 $Y=0.085
+ $X2=9.7 $Y2=0.38
r219 56 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.84 $Y2=0
r220 56 58 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.84 $Y2=0.535
r221 52 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.6 $Y=0.085
+ $X2=6.6 $Y2=0
r222 52 54 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.6 $Y=0.085
+ $X2=6.6 $Y2=0.38
r223 51 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.905 $Y=0 $X2=5.74
+ $Y2=0
r224 50 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=0 $X2=6.6
+ $Y2=0
r225 50 51 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.435 $Y=0
+ $X2=5.905 $Y2=0
r226 46 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.74 $Y=0.085
+ $X2=5.74 $Y2=0
r227 46 48 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.74 $Y=0.085
+ $X2=5.74 $Y2=0.36
r228 42 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0
r229 42 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0.36
r230 38 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=0.085
+ $X2=3.975 $Y2=0
r231 38 40 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=3.975 $Y=0.085
+ $X2=3.975 $Y2=0.465
r232 34 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=0.085
+ $X2=1.355 $Y2=0
r233 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.355 $Y=0.085
+ $X2=1.355 $Y2=0.36
r234 33 65 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.475
+ $Y2=0
r235 32 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=0
+ $X2=1.355 $Y2=0
r236 32 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.19 $Y=0 $X2=0.62
+ $Y2=0
r237 28 65 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.475 $Y=0.085
+ $X2=0.475 $Y2=0
r238 28 30 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.475 $Y=0.085
+ $X2=0.475 $Y2=0.38
r239 9 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.56
+ $Y=0.235 $X2=9.7 $Y2=0.38
r240 8 58 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=8.7
+ $Y=0.235 $X2=8.84 $Y2=0.535
r241 7 122 121.333 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_NDIFF $count=1
+ $X=7.32 $Y=0.235 $X2=7.46 $Y2=0.785
r242 7 120 121.333 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1
+ $X=7.32 $Y=0.235 $X2=7.46 $Y2=0.36
r243 6 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.46
+ $Y=0.235 $X2=6.6 $Y2=0.38
r244 5 48 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.6
+ $Y=0.235 $X2=5.74 $Y2=0.36
r245 4 44 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.74
+ $Y=0.235 $X2=4.88 $Y2=0.36
r246 3 40 182 $w=1.7e-07 $l=3.07083e-07 $layer=licon1_NDIFF $count=1 $X=3.795
+ $Y=0.235 $X2=3.975 $Y2=0.465
r247 2 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.215
+ $Y=0.235 $X2=1.355 $Y2=0.36
r248 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.37
+ $Y=0.235 $X2=0.495 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_4%A_157_47# 1 2 3 4 15 17 18 19 27
r34 25 27 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.645 $Y=0.42
+ $X2=3.505 $Y2=0.42
r35 23 30 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.87 $Y=0.42 $X2=1.78
+ $Y2=0.42
r36 23 25 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=1.87 $Y=0.42
+ $X2=2.645 $Y2=0.42
r37 20 22 3.69697 $w=1.78e-07 $l=6e-08 $layer=LI1_cond $X=1.78 $Y=1.01 $X2=1.78
+ $Y2=0.95
r38 19 30 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0.585
+ $X2=1.78 $Y2=0.42
r39 19 22 22.4899 $w=1.78e-07 $l=3.65e-07 $layer=LI1_cond $X=1.78 $Y=0.585
+ $X2=1.78 $Y2=0.95
r40 17 20 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.69 $Y=1.095
+ $X2=1.78 $Y2=1.01
r41 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.69 $Y=1.095
+ $X2=1.02 $Y2=1.095
r42 13 18 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.905 $Y=1.01
+ $X2=1.02 $Y2=1.095
r43 13 15 29.5627 $w=2.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.905 $Y=1.01
+ $X2=0.905 $Y2=0.42
r44 4 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.505 $Y2=0.42
r45 3 25 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.505
+ $Y=0.235 $X2=2.645 $Y2=0.42
r46 2 30 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.235 $X2=1.785 $Y2=0.42
r47 2 22 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.235 $X2=1.785 $Y2=0.95
r48 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.785
+ $Y=0.235 $X2=0.925 $Y2=0.42
.ends

