# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfxtp_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfxtp_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.215000 2.295000 1.885000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.605000 1.920000 13.275000 2.960000 ;
        RECT 12.685000 0.325000 13.075000 0.785000 ;
        RECT 12.905000 0.785000 13.075000 1.920000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.245000 3.715000 1.915000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.689000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 1.515000 0.875000 1.845000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.950000 1.180000 4.280000 1.510000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.245000 13.920000 3.415000 ;
      RECT  0.115000  0.605000  0.670000 1.165000 ;
      RECT  0.115000  1.165000  1.755000 1.335000 ;
      RECT  0.115000  1.335000  0.365000 3.065000 ;
      RECT  0.645000  2.025000  0.975000 3.245000 ;
      RECT  1.160000  0.085000  1.490000 0.985000 ;
      RECT  1.200000  2.065000  1.530000 2.505000 ;
      RECT  1.200000  2.505000  3.590000 2.675000 ;
      RECT  1.200000  2.675000  1.530000 3.065000 ;
      RECT  1.425000  1.335000  1.755000 1.835000 ;
      RECT  1.730000  2.065000  2.645000 2.155000 ;
      RECT  1.730000  2.155000  6.885000 2.325000 ;
      RECT  2.200000  0.605000  2.645000 1.035000 ;
      RECT  2.475000  1.035000  2.645000 2.065000 ;
      RECT  2.730000  2.855000  3.060000 3.245000 ;
      RECT  3.090000  0.085000  3.420000 1.065000 ;
      RECT  3.260000  2.675000  3.590000 3.065000 ;
      RECT  3.645000  0.310000  3.975000 0.830000 ;
      RECT  3.645000  0.830000  5.045000 1.000000 ;
      RECT  3.905000  1.715000  4.630000 1.975000 ;
      RECT  4.435000  0.085000  4.765000 0.650000 ;
      RECT  4.435000  2.505000  4.765000 3.245000 ;
      RECT  4.460000  1.000000  5.045000 1.530000 ;
      RECT  4.460000  1.530000  4.630000 1.715000 ;
      RECT  4.965000  1.715000  5.820000 1.975000 ;
      RECT  5.225000  0.310000  5.555000 1.305000 ;
      RECT  5.225000  1.305000  5.820000 1.715000 ;
      RECT  5.780000  0.265000  7.825000 0.435000 ;
      RECT  5.780000  0.435000  6.030000 1.125000 ;
      RECT  6.210000  0.615000  7.320000 0.785000 ;
      RECT  6.210000  0.785000  6.380000 1.715000 ;
      RECT  6.210000  1.715000  6.885000 2.155000 ;
      RECT  6.555000  2.325000  6.885000 2.755000 ;
      RECT  6.560000  0.965000  6.890000 1.365000 ;
      RECT  6.560000  1.365000  7.415000 1.535000 ;
      RECT  7.070000  0.785000  7.320000 1.185000 ;
      RECT  7.085000  1.535000  7.415000 1.665000 ;
      RECT  7.085000  1.665000  8.790000 1.835000 ;
      RECT  7.085000  1.835000  7.415000 2.755000 ;
      RECT  7.575000  0.435000  7.825000 0.975000 ;
      RECT  7.880000  1.155000  8.210000 1.485000 ;
      RECT  8.040000  0.895000  9.275000 1.065000 ;
      RECT  8.040000  1.065000  8.210000 1.155000 ;
      RECT  8.080000  0.085000  8.410000 0.715000 ;
      RECT  8.105000  2.015000  8.435000 3.245000 ;
      RECT  8.460000  1.245000  8.790000 1.665000 ;
      RECT  8.945000  0.265000 10.685000 0.435000 ;
      RECT  8.945000  0.435000  9.275000 0.895000 ;
      RECT  9.105000  1.065000  9.275000 1.715000 ;
      RECT  9.105000  1.715000  9.435000 2.755000 ;
      RECT  9.530000  0.615000 11.160000 0.785000 ;
      RECT  9.530000  0.785000  9.770000 1.215000 ;
      RECT  9.840000  1.475000 11.675000 1.645000 ;
      RECT  9.840000  1.645000 10.170000 2.825000 ;
      RECT  9.940000  0.965000 10.270000 1.475000 ;
      RECT 10.775000  0.965000 12.725000 1.135000 ;
      RECT 10.775000  1.135000 11.105000 1.295000 ;
      RECT 10.910000  0.325000 11.160000 0.615000 ;
      RECT 10.965000  1.825000 11.295000 3.245000 ;
      RECT 11.340000  0.085000 11.670000 0.785000 ;
      RECT 11.345000  1.315000 11.675000 1.475000 ;
      RECT 11.570000  1.825000 12.025000 2.825000 ;
      RECT 11.855000  1.135000 12.025000 1.825000 ;
      RECT 12.130000  0.325000 12.460000 0.785000 ;
      RECT 12.130000  0.785000 12.300000 0.965000 ;
      RECT 12.395000  1.135000 12.725000 1.635000 ;
      RECT 13.475000  0.085000 13.805000 0.785000 ;
      RECT 13.475000  1.920000 13.805000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfxtp_lp
END LIBRARY
