* File: sky130_fd_sc_lp__sdfrbp_1.pex.spice
* Created: Wed Sep  2 10:34:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%SCE 3 5 6 8 9 11 12 14 16 21 23 25 26 29 30
+ 34 35 41 45 47 53 55
c104 29 0 5.71674e-20 $X=2.235 $Y=1.56
r105 47 53 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=1.14 $Y=1.7 $X2=1.2
+ $Y2=1.7
r106 39 41 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=0.97 $Y=1.7 $X2=1.07
+ $Y2=1.7
r107 35 55 5.94776 $w=3.28e-07 $l=9.3e-08 $layer=LI1_cond $X=1.212 $Y=1.7
+ $X2=1.305 $Y2=1.7
r108 35 53 0.41907 $w=3.28e-07 $l=1.2e-08 $layer=LI1_cond $X=1.212 $Y=1.7
+ $X2=1.2 $Y2=1.7
r109 35 47 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=1.07 $Y=1.7 $X2=1.14
+ $Y2=1.7
r110 35 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.07
+ $Y=1.7 $X2=1.07 $Y2=1.7
r111 34 35 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.72 $Y=1.7
+ $X2=1.07 $Y2=1.7
r112 30 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.56
+ $X2=2.235 $Y2=1.395
r113 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.56 $X2=2.235 $Y2=1.56
r114 26 29 8.04881 $w=3.13e-07 $l=2.2e-07 $layer=LI1_cond $X=2.227 $Y=1.78
+ $X2=2.227 $Y2=1.56
r115 26 55 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.07 $Y=1.78
+ $X2=1.305 $Y2=1.78
r116 25 45 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=2.325 $Y=1.21
+ $X2=2.325 $Y2=1.395
r117 24 25 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=2.345 $Y=1.06
+ $X2=2.345 $Y2=1.21
r118 21 24 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.365 $Y=0.615
+ $X2=2.365 $Y2=1.06
r119 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.4 $Y=2.345
+ $X2=1.4 $Y2=2.775
r120 13 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.045 $Y=2.27
+ $X2=0.97 $Y2=2.27
r121 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.325 $Y=2.27
+ $X2=1.4 $Y2=2.345
r122 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.325 $Y=2.27
+ $X2=1.045 $Y2=2.27
r123 9 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.97 $Y=2.345
+ $X2=0.97 $Y2=2.27
r124 9 11 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.97 $Y=2.345
+ $X2=0.97 $Y2=2.775
r125 8 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.97 $Y=2.195
+ $X2=0.97 $Y2=2.27
r126 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.865
+ $X2=0.97 $Y2=1.7
r127 7 8 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.97 $Y=1.865
+ $X2=0.97 $Y2=2.195
r128 5 39 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.895 $Y=1.7
+ $X2=0.97 $Y2=1.7
r129 5 6 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=0.895 $Y=1.7
+ $X2=0.55 $Y2=1.7
r130 1 6 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.475 $Y=1.535
+ $X2=0.55 $Y2=1.7
r131 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.475 $Y=1.535
+ $X2=0.475 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%A_27_75# 1 2 7 9 12 16 19 20 21 24 25 29 33
+ 34 36 37
c82 24 0 1.95141e-19 $X=1.07 $Y=1.07
r83 34 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=2.13
+ $X2=2.21 $Y2=2.295
r84 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=2.13 $X2=2.21 $Y2=2.13
r85 31 37 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=2.125
+ $X2=0.755 $Y2=2.125
r86 31 33 79.4848 $w=1.78e-07 $l=1.29e-06 $layer=LI1_cond $X=0.92 $Y=2.125
+ $X2=2.21 $Y2=2.125
r87 27 37 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.755 $Y=2.215
+ $X2=0.755 $Y2=2.125
r88 27 29 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.755 $Y=2.215
+ $X2=0.755 $Y2=2.6
r89 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.07 $X2=1.07 $Y2=1.07
r90 22 36 0.546715 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=0.365 $Y=1.07
+ $X2=0.26 $Y2=1.07
r91 22 24 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.365 $Y=1.07
+ $X2=1.07 $Y2=1.07
r92 20 37 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.59 $Y=2.125
+ $X2=0.755 $Y2=2.125
r93 20 21 16.3283 $w=1.78e-07 $l=2.65e-07 $layer=LI1_cond $X=0.59 $Y=2.125
+ $X2=0.325 $Y2=2.125
r94 19 21 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.325 $Y2=2.125
r95 18 36 7.95398 $w=1.9e-07 $l=1.74714e-07 $layer=LI1_cond $X=0.24 $Y=1.235
+ $X2=0.26 $Y2=1.07
r96 18 19 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.24 $Y=1.235 $X2=0.24
+ $Y2=2.035
r97 14 36 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=0.905
+ $X2=0.26 $Y2=1.07
r98 14 16 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=0.26 $Y=0.905
+ $X2=0.26 $Y2=0.65
r99 12 42 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.19 $Y=2.775
+ $X2=2.19 $Y2=2.295
r100 7 25 68.7189 $w=2.49e-07 $l=4.29651e-07 $layer=POLY_cond $X=1.425 $Y=0.905
+ $X2=1.07 $Y2=1.07
r101 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.425 $Y=0.905
+ $X2=1.425 $Y2=0.585
r102 2 29 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.63
+ $Y=2.455 $X2=0.755 $Y2=2.6
r103 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.375 $X2=0.26 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%D 1 3 7 9 10
c43 7 0 9.68398e-20 $X=1.935 $Y=0.615
c44 1 0 1.95141e-19 $X=1.76 $Y=1.595
r45 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.64
+ $Y=1.43 $X2=1.64 $Y2=1.43
r46 10 15 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.64 $Y=1.295
+ $X2=1.64 $Y2=1.43
r47 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.64 $Y=0.925
+ $X2=1.64 $Y2=1.295
r48 5 14 77.8315 $w=3.19e-07 $l=5.12494e-07 $layer=POLY_cond $X=1.935 $Y=1.005
+ $X2=1.742 $Y2=1.43
r49 5 7 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.935 $Y=1.005
+ $X2=1.935 $Y2=0.615
r50 1 14 38.5462 $w=3.19e-07 $l=1.73767e-07 $layer=POLY_cond $X=1.76 $Y=1.595
+ $X2=1.742 $Y2=1.43
r51 1 3 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.76 $Y=1.595
+ $X2=1.76 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%SCD 3 7 11 12 13 14 15 20
c46 7 0 2.40407e-19 $X=2.725 $Y=0.615
r47 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.775
+ $Y=1.615 $X2=2.775 $Y2=1.615
r48 14 15 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.707 $Y=1.665
+ $X2=2.707 $Y2=2.035
r49 14 21 1.88925 $w=3.03e-07 $l=5e-08 $layer=LI1_cond $X=2.707 $Y=1.665
+ $X2=2.707 $Y2=1.615
r50 13 21 12.0912 $w=3.03e-07 $l=3.2e-07 $layer=LI1_cond $X=2.707 $Y=1.295
+ $X2=2.707 $Y2=1.615
r51 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.775 $Y=1.955
+ $X2=2.775 $Y2=1.615
r52 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.955
+ $X2=2.775 $Y2=2.12
r53 10 20 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.45
+ $X2=2.775 $Y2=1.615
r54 7 10 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=2.725 $Y=0.615
+ $X2=2.725 $Y2=1.45
r55 3 12 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.685 $Y=2.775
+ $X2=2.685 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%CLK 3 7 11 13 15 17 31
c46 17 0 9.87826e-20 $X=4.56 $Y=1.665
c47 7 0 2.77195e-20 $X=4.555 $Y=0.805
r48 30 31 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=4.555 $Y=1.375
+ $X2=4.615 $Y2=1.375
r49 28 30 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=4.38 $Y=1.375
+ $X2=4.555 $Y2=1.375
r50 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.38
+ $Y=1.375 $X2=4.38 $Y2=1.375
r51 25 28 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=4.125 $Y=1.375
+ $X2=4.38 $Y2=1.375
r52 17 29 3.71197 $w=5.78e-07 $l=1.8e-07 $layer=LI1_cond $X=4.56 $Y=1.49
+ $X2=4.38 $Y2=1.49
r53 15 29 6.18661 $w=5.78e-07 $l=3e-07 $layer=LI1_cond $X=4.08 $Y=1.49 $X2=4.38
+ $Y2=1.49
r54 13 15 9.89858 $w=5.78e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.49 $X2=4.08
+ $Y2=1.49
r55 9 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.615 $Y=1.54
+ $X2=4.615 $Y2=1.375
r56 9 11 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=4.615 $Y=1.54
+ $X2=4.615 $Y2=2.465
r57 5 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.555 $Y=1.21
+ $X2=4.555 $Y2=1.375
r58 5 7 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.555 $Y=1.21
+ $X2=4.555 $Y2=0.805
r59 1 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.125 $Y=1.21
+ $X2=4.125 $Y2=1.375
r60 1 3 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.125 $Y=1.21
+ $X2=4.125 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%A_1024_367# 1 2 9 11 15 19 22 24 26 30 31
+ 33 34 35 38 41 42 44 48 49 52 53 58
c165 53 0 8.80756e-20 $X=6.025 $Y=1.525
c166 52 0 1.9886e-19 $X=9.635 $Y=2.155
c167 41 0 1.1867e-19 $X=9.265 $Y=1.255
c168 11 0 1.24503e-19 $X=7 $Y=1.525
r169 52 62 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=9.63 $Y=2.155
+ $X2=9.63 $Y2=2.32
r170 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.635
+ $Y=2.155 $X2=9.635 $Y2=2.155
r171 49 51 15.5951 $w=3.27e-07 $l=4.18e-07 $layer=LI1_cond $X=9.217 $Y=2.135
+ $X2=9.635 $Y2=2.135
r172 45 56 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=6.025 $Y=1.805
+ $X2=6.025 $Y2=1.97
r173 45 53 37.9812 $w=4.1e-07 $l=2.8e-07 $layer=POLY_cond $X=6.025 $Y=1.805
+ $X2=6.025 $Y2=1.525
r174 44 47 4.25178 $w=7.03e-07 $l=5.18218e-07 $layer=LI1_cond $X=5.67 $Y=1.805
+ $X2=5.26 $Y2=2.05
r175 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.985
+ $Y=1.805 $X2=5.985 $Y2=1.805
r176 42 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.265 $Y=1.255
+ $X2=9.265 $Y2=1.09
r177 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.265
+ $Y=1.255 $X2=9.265 $Y2=1.255
r178 39 49 1.98942 $w=2.65e-07 $l=1.85e-07 $layer=LI1_cond $X=9.217 $Y=1.95
+ $X2=9.217 $Y2=2.135
r179 39 41 30.2244 $w=2.63e-07 $l=6.95e-07 $layer=LI1_cond $X=9.217 $Y=1.95
+ $X2=9.217 $Y2=1.255
r180 38 48 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=9.217 $Y=1.222
+ $X2=9.217 $Y2=1.09
r181 38 41 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=9.217 $Y=1.222
+ $X2=9.217 $Y2=1.255
r182 36 48 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.17 $Y=0.89 $X2=9.17
+ $Y2=1.09
r183 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.085 $Y=0.805
+ $X2=9.17 $Y2=0.89
r184 34 35 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=9.085 $Y=0.805
+ $X2=7.78 $Y2=0.805
r185 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.695 $Y=0.72
+ $X2=7.78 $Y2=0.805
r186 32 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.695 $Y=0.425
+ $X2=7.695 $Y2=0.72
r187 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.61 $Y=0.34
+ $X2=7.695 $Y2=0.425
r188 30 31 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=7.61 $Y=0.34
+ $X2=6.175 $Y2=0.34
r189 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.09 $Y=0.425
+ $X2=6.175 $Y2=0.34
r190 24 44 19.8915 $w=7.03e-07 $l=8.59724e-07 $layer=LI1_cond $X=6.09 $Y=1.13
+ $X2=5.67 $Y2=1.805
r191 24 28 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.09 $Y=1.13
+ $X2=6.09 $Y2=0.425
r192 24 26 9.21954 $w=2.98e-07 $l=2.4e-07 $layer=LI1_cond $X=5.335 $Y=1.085
+ $X2=5.335 $Y2=0.845
r193 22 62 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.69 $Y=2.69
+ $X2=9.69 $Y2=2.32
r194 19 58 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.175 $Y=0.66
+ $X2=9.175 $Y2=1.09
r195 13 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=7.075 $Y=1.45
+ $X2=7.075 $Y2=0.805
r196 12 53 26.4667 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=6.23 $Y=1.525
+ $X2=6.025 $Y2=1.525
r197 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7 $Y=1.525
+ $X2=7.075 $Y2=1.45
r198 11 12 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7 $Y=1.525 $X2=6.23
+ $Y2=1.525
r199 9 56 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.155 $Y=2.525
+ $X2=6.155 $Y2=1.97
r200 2 47 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=5.12
+ $Y=1.835 $X2=5.26 $Y2=2.05
r201 1 26 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=5.18
+ $Y=0.595 $X2=5.32 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%A_1374_362# 1 2 9 13 17 18 20 21 22 24 26
+ 28
c85 22 0 1.9886e-19 $X=8.787 $Y=2.002
c86 18 0 8.87177e-20 $X=7.15 $Y=1.99
c87 17 0 6.31644e-20 $X=7.15 $Y=1.99
r88 26 30 4.0965 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=8.83 $Y=1.295
+ $X2=8.83 $Y2=1.177
r89 26 28 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=8.83 $Y=1.295
+ $X2=8.83 $Y2=1.875
r90 22 28 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=8.787 $Y=2.002
+ $X2=8.787 $Y2=1.875
r91 22 24 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=8.787 $Y=2.002
+ $X2=8.787 $Y2=2.04
r92 20 30 2.95087 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=1.177
+ $X2=8.83 $Y2=1.177
r93 20 21 73.5602 $w=2.33e-07 $l=1.5e-06 $layer=LI1_cond $X=8.745 $Y=1.177
+ $X2=7.245 $Y2=1.177
r94 18 31 31.0723 $w=3.18e-07 $l=2.05e-07 $layer=POLY_cond $X=7.15 $Y=1.925
+ $X2=6.945 $Y2=1.925
r95 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.15
+ $Y=1.99 $X2=7.15 $Y2=1.99
r96 15 21 5.60639 $w=2.58e-07 $l=1.56665e-07 $layer=LI1_cond $X=7.155 $Y=1.295
+ $X2=7.245 $Y2=1.177
r97 15 17 42.8232 $w=1.78e-07 $l=6.95e-07 $layer=LI1_cond $X=7.155 $Y=1.295
+ $X2=7.155 $Y2=1.99
r98 11 18 43.1981 $w=3.18e-07 $l=3.83112e-07 $layer=POLY_cond $X=7.435 $Y=1.695
+ $X2=7.15 $Y2=1.925
r99 11 13 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=7.435 $Y=1.695
+ $X2=7.435 $Y2=0.805
r100 7 31 20.3436 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.945 $Y=2.155
+ $X2=6.945 $Y2=1.925
r101 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.945 $Y=2.155
+ $X2=6.945 $Y2=2.525
r102 2 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.63
+ $Y=1.895 $X2=8.77 $Y2=2.04
r103 1 30 182 $w=1.7e-07 $l=9.08364e-07 $layer=licon1_NDIFF $count=1 $X=8.53
+ $Y=0.34 $X2=8.75 $Y2=1.145
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%RESET_B 4 7 9 10 11 13 17 20 22 28 31 32 33
+ 34 35 36 44 49 50 53 56 58 59 60
c210 58 0 1.13095e-19 $X=10.7 $Y=2.035
c211 56 0 8.87177e-20 $X=7.89 $Y=1.99
c212 53 0 2.28509e-19 $X=7.795 $Y=2.03
c213 35 0 3.13244e-19 $X=10.175 $Y=2.035
c214 31 0 5.68043e-20 $X=10.62 $Y=1.02
c215 28 0 1.03579e-19 $X=10.72 $Y=2.755
c216 22 0 2.45352e-20 $X=10.62 $Y=1.6
r217 59 69 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=10.7 $Y=2.035
+ $X2=10.32 $Y2=2.035
r218 58 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.7 $Y=2.035
+ $X2=10.7 $Y2=2.2
r219 58 60 44.2063 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.7 $Y=2.035
+ $X2=10.7 $Y2=1.87
r220 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.7
+ $Y=2.035 $X2=10.7 $Y2=2.035
r221 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.89
+ $Y=1.99 $X2=7.89 $Y2=1.99
r222 53 55 14.4448 $w=3.17e-07 $l=9.5e-08 $layer=POLY_cond $X=7.795 $Y=2.03
+ $X2=7.89 $Y2=2.03
r223 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.475
+ $Y=2.115 $X2=3.475 $Y2=2.115
r224 46 49 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.225 $Y=2.115
+ $X2=3.475 $Y2=2.115
r225 44 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=2.035
+ $X2=10.32 $Y2=2.035
r226 42 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r227 38 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=2.035
+ $X2=3.6 $Y2=2.035
r228 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r229 35 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.175 $Y=2.035
+ $X2=10.32 $Y2=2.035
r230 35 36 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=10.175 $Y=2.035
+ $X2=8.065 $Y2=2.035
r231 34 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=2.035
+ $X2=3.6 $Y2=2.035
r232 33 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r233 33 34 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=3.745 $Y2=2.035
r234 31 32 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=10.625 $Y=1.02
+ $X2=10.625 $Y2=1.52
r235 30 31 25.4904 $w=1.6e-07 $l=5.5e-08 $layer=POLY_cond $X=10.62 $Y=0.965
+ $X2=10.62 $Y2=1.02
r236 28 61 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=10.72 $Y=2.755
+ $X2=10.72 $Y2=2.2
r237 22 32 37.4638 $w=1.6e-07 $l=8e-08 $layer=POLY_cond $X=10.62 $Y=1.6
+ $X2=10.62 $Y2=1.52
r238 22 60 125.135 $w=1.6e-07 $l=2.7e-07 $layer=POLY_cond $X=10.62 $Y=1.6
+ $X2=10.62 $Y2=1.87
r239 20 30 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=10.615 $Y=0.55
+ $X2=10.615 $Y2=0.965
r240 15 53 20.269 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.795 $Y=1.82
+ $X2=7.795 $Y2=2.03
r241 15 17 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=7.795 $Y=1.82
+ $X2=7.795 $Y2=0.805
r242 14 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.795 $Y=0.255
+ $X2=7.795 $Y2=0.805
r243 11 53 28.8896 $w=3.17e-07 $l=2.89828e-07 $layer=POLY_cond $X=7.605 $Y=2.24
+ $X2=7.795 $Y2=2.03
r244 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.605 $Y=2.24
+ $X2=7.605 $Y2=2.525
r245 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.72 $Y=0.18
+ $X2=7.795 $Y2=0.255
r246 9 10 2266.43 $w=1.5e-07 $l=4.42e-06 $layer=POLY_cond $X=7.72 $Y=0.18
+ $X2=3.3 $Y2=0.18
r247 5 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=2.28
+ $X2=3.225 $Y2=2.115
r248 5 7 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.225 $Y=2.28
+ $X2=3.225 $Y2=2.775
r249 2 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=1.95
+ $X2=3.225 $Y2=2.115
r250 2 4 684.543 $w=1.5e-07 $l=1.335e-06 $layer=POLY_cond $X=3.225 $Y=1.95
+ $X2=3.225 $Y2=0.615
r251 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.225 $Y=0.255
+ $X2=3.3 $Y2=0.18
r252 1 4 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.225 $Y=0.255
+ $X2=3.225 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%A_1246_463# 1 2 3 12 16 18 23 24 27 28 30
+ 31 35 38 41 42
c116 31 0 1.55177e-19 $X=8.41 $Y=1.555
c117 30 0 1.65324e-20 $X=8.41 $Y=1.555
c118 28 0 1.24503e-19 $X=7.605 $Y=1.557
c119 23 0 3.43879e-19 $X=6.81 $Y=2.335
c120 18 0 1.2249e-19 $X=6.725 $Y=2.635
c121 12 0 1.1867e-19 $X=8.455 $Y=0.66
r122 38 40 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=0.815
+ $X2=6.835 $Y2=0.98
r123 33 42 3.64284 $w=2.7e-07 $l=2.52785e-07 $layer=LI1_cond $X=7.605 $Y=2.51
+ $X2=7.425 $Y2=2.335
r124 33 35 7.07929 $w=3.48e-07 $l=2.15e-07 $layer=LI1_cond $X=7.605 $Y=2.51
+ $X2=7.82 $Y2=2.51
r125 31 45 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=8.437 $Y=1.555
+ $X2=8.437 $Y2=1.72
r126 31 44 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=8.437 $Y=1.555
+ $X2=8.437 $Y2=1.39
r127 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.41
+ $Y=1.555 $X2=8.41 $Y2=1.555
r128 28 30 48.2604 $w=1.83e-07 $l=8.05e-07 $layer=LI1_cond $X=7.605 $Y=1.557
+ $X2=8.41 $Y2=1.557
r129 27 42 2.83584 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=7.515 $Y=2.335
+ $X2=7.425 $Y2=2.335
r130 26 28 6.81816 $w=1.85e-07 $l=1.30457e-07 $layer=LI1_cond $X=7.515 $Y=1.65
+ $X2=7.605 $Y2=1.557
r131 26 27 42.2071 $w=1.78e-07 $l=6.85e-07 $layer=LI1_cond $X=7.515 $Y=1.65
+ $X2=7.515 $Y2=2.335
r132 25 41 3.91525 $w=2.35e-07 $l=1.63936e-07 $layer=LI1_cond $X=6.905 $Y=2.43
+ $X2=6.815 $Y2=2.555
r133 24 42 3.64284 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.425 $Y=2.43
+ $X2=7.425 $Y2=2.335
r134 24 25 30.3541 $w=1.88e-07 $l=5.2e-07 $layer=LI1_cond $X=7.425 $Y=2.43
+ $X2=6.905 $Y2=2.43
r135 23 41 2.53056 $w=1.7e-07 $l=2.22486e-07 $layer=LI1_cond $X=6.81 $Y=2.335
+ $X2=6.815 $Y2=2.555
r136 23 40 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=6.81 $Y=2.335
+ $X2=6.81 $Y2=0.98
r137 18 41 3.91525 $w=2.35e-07 $l=1.23693e-07 $layer=LI1_cond $X=6.725 $Y=2.635
+ $X2=6.815 $Y2=2.555
r138 18 20 14.6113 $w=2.78e-07 $l=3.55e-07 $layer=LI1_cond $X=6.725 $Y=2.635
+ $X2=6.37 $Y2=2.635
r139 16 45 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=8.555 $Y=2.315
+ $X2=8.555 $Y2=1.72
r140 12 44 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=8.455 $Y=0.66
+ $X2=8.455 $Y2=1.39
r141 3 35 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=7.68
+ $Y=2.315 $X2=7.82 $Y2=2.52
r142 2 20 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=6.23
+ $Y=2.315 $X2=6.37 $Y2=2.595
r143 1 38 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=6.72
+ $Y=0.595 $X2=6.86 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%A_840_119# 1 2 9 13 15 17 19 20 21 22 23 26
+ 28 30 31 36 37 38 41 43 44 48 51 52 53 55
c175 55 0 2.77195e-20 $X=4.34 $Y=0.865
c176 52 0 8.80756e-20 $X=4.91 $Y=1.715
c177 38 0 1.65324e-20 $X=9.06 $Y=1.705
c178 9 0 9.87826e-20 $X=5.045 $Y=2.465
r179 60 61 2.14222 $w=4.5e-07 $l=2e-08 $layer=POLY_cond $X=5.065 $Y=1.382
+ $X2=5.045 $Y2=1.382
r180 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.065
+ $Y=1.51 $X2=5.065 $Y2=1.51
r181 52 59 10.3645 $w=3.61e-07 $l=2.56924e-07 $layer=LI1_cond $X=4.91 $Y=1.715
+ $X2=5.027 $Y2=1.51
r182 52 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.91 $Y=1.715
+ $X2=4.91 $Y2=1.95
r183 51 59 9.01265 $w=3.61e-07 $l=2.15708e-07 $layer=LI1_cond $X=4.91 $Y=1.345
+ $X2=5.027 $Y2=1.51
r184 50 51 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.91 $Y=1.03
+ $X2=4.91 $Y2=1.345
r185 49 55 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.425 $Y=0.945
+ $X2=4.34 $Y2=0.865
r186 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.825 $Y=0.945
+ $X2=4.91 $Y2=1.03
r187 48 49 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=4.825 $Y=0.945
+ $X2=4.425 $Y2=0.945
r188 44 53 7.24806 $w=2.65e-07 $l=1.69245e-07 $layer=LI1_cond $X=4.825 $Y=2.082
+ $X2=4.91 $Y2=1.95
r189 44 46 18.4826 $w=2.63e-07 $l=4.25e-07 $layer=LI1_cond $X=4.825 $Y=2.082
+ $X2=4.4 $Y2=2.082
r190 39 41 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=9.725 $Y=1.63
+ $X2=9.725 $Y2=0.55
r191 37 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.65 $Y=1.705
+ $X2=9.725 $Y2=1.63
r192 37 38 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=9.65 $Y=1.705
+ $X2=9.06 $Y2=1.705
r193 34 36 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.985 $Y=3.075
+ $X2=8.985 $Y2=2.315
r194 33 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.985 $Y=1.78
+ $X2=9.06 $Y2=1.705
r195 33 36 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=8.985 $Y=1.78
+ $X2=8.985 $Y2=2.315
r196 32 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.66 $Y=3.15
+ $X2=6.585 $Y2=3.15
r197 31 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.91 $Y=3.15
+ $X2=8.985 $Y2=3.075
r198 31 32 1153.72 $w=1.5e-07 $l=2.25e-06 $layer=POLY_cond $X=8.91 $Y=3.15
+ $X2=6.66 $Y2=3.15
r199 28 30 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.645 $Y=1.09
+ $X2=6.645 $Y2=0.805
r200 24 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.585 $Y=3.075
+ $X2=6.585 $Y2=3.15
r201 24 26 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.585 $Y=3.075
+ $X2=6.585 $Y2=2.525
r202 22 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.51 $Y=3.15
+ $X2=6.585 $Y2=3.15
r203 22 23 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=6.51 $Y=3.15 $X2=5.61
+ $Y2=3.15
r204 21 64 31.0404 $w=4.5e-07 $l=2.51722e-07 $layer=POLY_cond $X=5.61 $Y=1.165
+ $X2=5.535 $Y2=1.382
r205 20 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.57 $Y=1.165
+ $X2=6.645 $Y2=1.09
r206 20 21 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=6.57 $Y=1.165
+ $X2=5.61 $Y2=1.165
r207 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.535 $Y=3.075
+ $X2=5.61 $Y2=3.15
r208 18 64 28.7666 $w=1.5e-07 $l=2.93e-07 $layer=POLY_cond $X=5.535 $Y=1.675
+ $X2=5.535 $Y2=1.382
r209 18 19 717.872 $w=1.5e-07 $l=1.4e-06 $layer=POLY_cond $X=5.535 $Y=1.675
+ $X2=5.535 $Y2=3.075
r210 15 64 28.7666 $w=1.5e-07 $l=2.92e-07 $layer=POLY_cond $X=5.535 $Y=1.09
+ $X2=5.535 $Y2=1.382
r211 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.535 $Y=1.09
+ $X2=5.535 $Y2=0.805
r212 11 64 46.0578 $w=4.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.105 $Y=1.382
+ $X2=5.535 $Y2=1.382
r213 11 60 4.28444 $w=4.5e-07 $l=4e-08 $layer=POLY_cond $X=5.105 $Y=1.382
+ $X2=5.065 $Y2=1.382
r214 11 13 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.105 $Y=1.26
+ $X2=5.105 $Y2=0.805
r215 7 61 28.7666 $w=1.5e-07 $l=2.93e-07 $layer=POLY_cond $X=5.045 $Y=1.675
+ $X2=5.045 $Y2=1.382
r216 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.045 $Y=1.675
+ $X2=5.045 $Y2=2.465
r217 2 46 600 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.835 $X2=4.4 $Y2=2.08
r218 1 55 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.595 $X2=4.34 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%A_2002_42# 1 2 9 13 15 17 19 23 24 26 27 31
+ 34 36
c114 27 0 1.85637e-19 $X=10.17 $Y=1.08
c115 15 0 2.45352e-20 $X=10.635 $Y=1.08
r116 31 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.175 $Y=1.25
+ $X2=10.175 $Y2=1.415
r117 31 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.175 $Y=1.25
+ $X2=10.175 $Y2=1.085
r118 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.175
+ $Y=1.25 $X2=10.175 $Y2=1.25
r119 27 30 5.76222 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=10.17 $Y=1.08
+ $X2=10.17 $Y2=1.25
r120 25 34 9.71229 $w=3.58e-07 $l=2.85e-07 $layer=LI1_cond $X=11.475 $Y=0.837
+ $X2=11.19 $Y2=0.837
r121 25 26 35.5754 $w=2.28e-07 $l=7.1e-07 $layer=LI1_cond $X=11.475 $Y=0.975
+ $X2=11.475 $Y2=1.685
r122 23 26 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=11.36 $Y=1.77
+ $X2=11.475 $Y2=1.685
r123 23 24 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.36 $Y=1.77
+ $X2=11.135 $Y2=1.77
r124 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.05 $Y=1.855
+ $X2=11.135 $Y2=1.77
r125 21 36 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=11.05 $Y=1.855
+ $X2=11.05 $Y2=2.37
r126 17 36 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=10.962 $Y=2.542
+ $X2=10.962 $Y2=2.37
r127 17 19 7.11508 $w=3.43e-07 $l=2.13e-07 $layer=LI1_cond $X=10.962 $Y=2.542
+ $X2=10.962 $Y2=2.755
r128 16 27 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=10.34 $Y=1.08
+ $X2=10.17 $Y2=1.08
r129 15 34 22.2952 $w=3.58e-07 $l=6.655e-07 $layer=LI1_cond $X=10.635 $Y=1.08
+ $X2=11.19 $Y2=0.837
r130 15 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.635 $Y=1.08
+ $X2=10.34 $Y2=1.08
r131 13 39 653.777 $w=1.5e-07 $l=1.275e-06 $layer=POLY_cond $X=10.245 $Y=2.69
+ $X2=10.245 $Y2=1.415
r132 9 38 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=10.085 $Y=0.55
+ $X2=10.085 $Y2=1.085
r133 2 19 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=10.795
+ $Y=2.545 $X2=10.935 $Y2=2.755
r134 1 34 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=11.05
+ $Y=0.34 $X2=11.19 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%A_1812_379# 1 2 9 11 15 16 17 18 21 24 26
+ 28 31 35 37 38 41 43 45 50 52 53 55 59 62 64 70 71 76 82 83 87 88 96
c214 71 0 1.42329e-19 $X=10.595 $Y=1.43
r215 95 96 36.5941 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=11.15 $Y=1.31
+ $X2=11.26 $Y2=1.31
r216 88 99 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.33 $Y=1.51
+ $X2=13.33 $Y2=1.675
r217 88 98 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.33 $Y=1.51
+ $X2=13.33 $Y2=1.345
r218 87 88 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.33
+ $Y=1.51 $X2=13.33 $Y2=1.51
r219 84 87 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=13.135 $Y=1.51
+ $X2=13.33 $Y2=1.51
r220 82 83 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.135
+ $Y=2.6 $X2=12.135 $Y2=2.6
r221 77 95 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=11.095 $Y=1.31
+ $X2=11.15 $Y2=1.31
r222 77 92 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=11.095 $Y=1.31
+ $X2=10.985 $Y2=1.31
r223 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.095
+ $Y=1.31 $X2=11.095 $Y2=1.31
r224 71 73 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.595 $Y=1.43
+ $X2=10.595 $Y2=1.6
r225 69 70 4.92405 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=9.975 $Y=1.62
+ $X2=10.06 $Y2=1.62
r226 64 66 12.4904 $w=4.03e-07 $l=4e-07 $layer=LI1_cond $X=9.627 $Y=0.535
+ $X2=9.627 $Y2=0.935
r227 61 84 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=13.135 $Y=1.675
+ $X2=13.135 $Y2=1.51
r228 61 62 45.5311 $w=1.88e-07 $l=7.8e-07 $layer=LI1_cond $X=13.135 $Y=1.675
+ $X2=13.135 $Y2=2.455
r229 60 82 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.3 $Y=2.54
+ $X2=12.135 $Y2=2.54
r230 59 62 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=13.04 $Y=2.54
+ $X2=13.135 $Y2=2.455
r231 59 60 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=13.04 $Y=2.54
+ $X2=12.3 $Y2=2.54
r232 56 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.68 $Y=1.43
+ $X2=10.595 $Y2=1.43
r233 55 76 6.43224 $w=2.13e-07 $l=1.2e-07 $layer=LI1_cond $X=11.082 $Y=1.43
+ $X2=11.082 $Y2=1.31
r234 55 56 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.975 $Y=1.43
+ $X2=10.68 $Y2=1.43
r235 53 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.51 $Y=1.6
+ $X2=10.595 $Y2=1.6
r236 53 70 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=10.51 $Y=1.6
+ $X2=10.06 $Y2=1.6
r237 51 69 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=9.975 $Y=1.725
+ $X2=9.975 $Y2=1.62
r238 51 52 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=9.975 $Y=1.725
+ $X2=9.975 $Y2=2.495
r239 50 69 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=9.69 $Y=1.62
+ $X2=9.975 $Y2=1.62
r240 50 66 23.872 $w=2.78e-07 $l=5.8e-07 $layer=LI1_cond $X=9.69 $Y=1.515
+ $X2=9.69 $Y2=0.935
r241 45 52 8.58847 $w=4.25e-07 $l=2.50926e-07 $layer=LI1_cond $X=9.89 $Y=2.707
+ $X2=9.975 $Y2=2.495
r242 45 47 14.5072 $w=4.23e-07 $l=5.35e-07 $layer=LI1_cond $X=9.89 $Y=2.707
+ $X2=9.355 $Y2=2.707
r243 44 83 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=12.135 $Y=3.075
+ $X2=12.135 $Y2=2.6
r244 37 38 30.125 $w=1.6e-07 $l=6.5e-08 $layer=POLY_cond $X=10.98 $Y=0.835
+ $X2=10.98 $Y2=0.9
r245 35 98 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=13.31 $Y=0.795
+ $X2=13.31 $Y2=1.345
r246 31 99 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=13.28 $Y=2.465
+ $X2=13.28 $Y2=1.675
r247 26 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.925 $Y=0.765
+ $X2=11.925 $Y2=0.84
r248 26 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.925 $Y=0.765
+ $X2=11.925 $Y2=0.445
r249 22 43 18.1413 $w=1.72e-07 $l=8.57321e-08 $layer=POLY_cond $X=11.685
+ $Y=1.295 $X2=11.662 $Y2=1.22
r250 22 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.685 $Y=1.295
+ $X2=11.685 $Y2=1.955
r251 21 43 18.1413 $w=1.72e-07 $l=7.5e-08 $layer=POLY_cond $X=11.662 $Y=1.145
+ $X2=11.662 $Y2=1.22
r252 20 41 134.857 $w=1.5e-07 $l=2.63e-07 $layer=POLY_cond $X=11.662 $Y=0.84
+ $X2=11.925 $Y2=0.84
r253 20 21 78.2182 $w=1.95e-07 $l=2.3e-07 $layer=POLY_cond $X=11.662 $Y=0.915
+ $X2=11.662 $Y2=1.145
r254 18 43 7.3104 $w=1.5e-07 $l=9.7e-08 $layer=POLY_cond $X=11.565 $Y=1.22
+ $X2=11.662 $Y2=1.22
r255 18 96 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=11.565 $Y=1.22
+ $X2=11.26 $Y2=1.22
r256 16 44 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=11.97 $Y=3.15
+ $X2=12.135 $Y2=3.075
r257 16 17 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=11.97 $Y=3.15
+ $X2=11.225 $Y2=3.15
r258 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.15 $Y=3.075
+ $X2=11.225 $Y2=3.15
r259 13 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.15 $Y=3.075
+ $X2=11.15 $Y2=2.755
r260 12 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.15 $Y=1.475
+ $X2=11.15 $Y2=1.31
r261 12 15 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=11.15 $Y=1.475
+ $X2=11.15 $Y2=2.755
r262 11 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.985 $Y=1.145
+ $X2=10.985 $Y2=1.31
r263 11 38 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=10.985 $Y=1.145
+ $X2=10.985 $Y2=0.9
r264 9 37 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.975 $Y=0.55
+ $X2=10.975 $Y2=0.835
r265 2 47 600 $w=1.7e-07 $l=9.005e-07 $layer=licon1_PDIFF $count=1 $X=9.06
+ $Y=1.895 $X2=9.355 $Y2=2.66
r266 1 64 182 $w=1.7e-07 $l=3.43948e-07 $layer=licon1_NDIFF $count=1 $X=9.25
+ $Y=0.34 $X2=9.51 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%A_2352_327# 1 2 7 11 13 15 16 19 23 25
r51 25 26 6.69143 $w=4.98e-07 $l=1.65e-07 $layer=LI1_cond $X=12.055 $Y=1.78
+ $X2=12.055 $Y2=1.615
r52 23 30 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.16 $Y=1.31
+ $X2=12.16 $Y2=1.4
r53 22 26 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=12.175 $Y=1.31
+ $X2=12.175 $Y2=1.615
r54 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.16
+ $Y=1.31 $X2=12.16 $Y2=1.31
r55 19 22 38.3409 $w=2.58e-07 $l=8.65e-07 $layer=LI1_cond $X=12.175 $Y=0.445
+ $X2=12.175 $Y2=1.31
r56 13 16 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=12.88 $Y=1.325
+ $X2=12.865 $Y2=1.4
r57 13 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=12.88 $Y=1.325
+ $X2=12.88 $Y2=0.795
r58 9 16 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=12.85 $Y=1.475
+ $X2=12.865 $Y2=1.4
r59 9 11 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=12.85 $Y=1.475
+ $X2=12.85 $Y2=2.465
r60 8 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.325 $Y=1.4
+ $X2=12.16 $Y2=1.4
r61 7 16 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=12.775 $Y=1.4
+ $X2=12.865 $Y2=1.4
r62 7 8 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=12.775 $Y=1.4
+ $X2=12.325 $Y2=1.4
r63 2 25 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=11.76
+ $Y=1.635 $X2=11.9 $Y2=1.78
r64 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12
+ $Y=0.235 $X2=12.14 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 60 63 64 66 67 69 70 72 73 75 76 78 79 80 82 106 124 125 128 131
c180 54 0 1.03579e-19 $X=11.47 $Y=2.13
r181 131 132 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r182 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r183 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r184 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r185 121 122 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r186 119 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r187 118 121 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r188 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r189 116 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r190 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r191 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r192 113 132 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=8.4 $Y2=3.33
r193 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r194 110 131 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.48 $Y=3.33
+ $X2=8.365 $Y2=3.33
r195 110 112 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=8.48 $Y=3.33
+ $X2=10.32 $Y2=3.33
r196 109 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r197 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r198 106 131 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.25 $Y=3.33
+ $X2=8.365 $Y2=3.33
r199 106 108 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.25 $Y=3.33
+ $X2=7.92 $Y2=3.33
r200 101 104 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r201 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r202 99 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r203 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r204 96 99 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r205 95 98 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r206 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r207 93 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r208 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r209 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r210 90 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r212 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r213 87 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.22 $Y2=3.33
r214 87 89 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.68 $Y2=3.33
r215 85 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r216 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r217 82 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=1.22 $Y2=3.33
r218 82 84 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.72 $Y2=3.33
r219 80 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r220 80 102 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=5.04 $Y2=3.33
r221 80 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r222 78 121 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=12.9 $Y=3.33
+ $X2=12.72 $Y2=3.33
r223 78 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.9 $Y=3.33
+ $X2=13.065 $Y2=3.33
r224 77 124 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=13.23 $Y=3.33
+ $X2=13.68 $Y2=3.33
r225 77 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.23 $Y=3.33
+ $X2=13.065 $Y2=3.33
r226 75 115 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=11.305 $Y=3.33
+ $X2=11.28 $Y2=3.33
r227 75 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.305 $Y=3.33
+ $X2=11.47 $Y2=3.33
r228 74 118 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=11.635 $Y=3.33
+ $X2=11.76 $Y2=3.33
r229 74 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.635 $Y=3.33
+ $X2=11.47 $Y2=3.33
r230 72 112 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=10.35 $Y=3.33
+ $X2=10.32 $Y2=3.33
r231 72 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.35 $Y=3.33
+ $X2=10.48 $Y2=3.33
r232 71 115 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.61 $Y=3.33
+ $X2=11.28 $Y2=3.33
r233 71 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.61 $Y=3.33
+ $X2=10.48 $Y2=3.33
r234 69 104 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.075 $Y=3.33
+ $X2=6.96 $Y2=3.33
r235 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.075 $Y=3.33
+ $X2=7.24 $Y2=3.33
r236 68 108 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=7.405 $Y=3.33
+ $X2=7.92 $Y2=3.33
r237 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=3.33
+ $X2=7.24 $Y2=3.33
r238 66 98 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=4.56 $Y2=3.33
r239 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=4.83 $Y2=3.33
r240 65 101 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.995 $Y=3.33
+ $X2=5.04 $Y2=3.33
r241 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=3.33
+ $X2=4.83 $Y2=3.33
r242 63 92 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.64 $Y2=3.33
r243 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.94 $Y2=3.33
r244 62 95 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=3.12 $Y2=3.33
r245 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=2.94 $Y2=3.33
r246 58 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.065 $Y=3.245
+ $X2=13.065 $Y2=3.33
r247 58 60 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=13.065 $Y=3.245
+ $X2=13.065 $Y2=2.92
r248 54 57 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=11.47 $Y=2.13
+ $X2=11.47 $Y2=2.8
r249 52 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.47 $Y=3.245
+ $X2=11.47 $Y2=3.33
r250 52 57 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=11.47 $Y=3.245
+ $X2=11.47 $Y2=2.8
r251 48 73 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.48 $Y=3.245
+ $X2=10.48 $Y2=3.33
r252 48 50 23.7137 $w=2.58e-07 $l=5.35e-07 $layer=LI1_cond $X=10.48 $Y=3.245
+ $X2=10.48 $Y2=2.71
r253 44 131 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.365 $Y=3.245
+ $X2=8.365 $Y2=3.33
r254 44 46 60.378 $w=2.28e-07 $l=1.205e-06 $layer=LI1_cond $X=8.365 $Y=3.245
+ $X2=8.365 $Y2=2.04
r255 40 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=3.245
+ $X2=7.24 $Y2=3.33
r256 40 42 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=7.24 $Y=3.245
+ $X2=7.24 $Y2=2.79
r257 36 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.83 $Y=3.245
+ $X2=4.83 $Y2=3.33
r258 36 38 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.83 $Y=3.245
+ $X2=4.83 $Y2=2.895
r259 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=3.245
+ $X2=2.94 $Y2=3.33
r260 32 34 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=2.94 $Y=3.245
+ $X2=2.94 $Y2=2.895
r261 28 128 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r262 28 30 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.6
r263 9 60 600 $w=1.7e-07 $l=1.15288e-06 $layer=licon1_PDIFF $count=1 $X=12.925
+ $Y=1.835 $X2=13.065 $Y2=2.92
r264 8 54 600 $w=1.7e-07 $l=5.73738e-07 $layer=licon1_PDIFF $count=1 $X=11.3
+ $Y=1.635 $X2=11.47 $Y2=2.13
r265 7 57 600 $w=1.7e-07 $l=3.31134e-07 $layer=licon1_PDIFF $count=1 $X=11.225
+ $Y=2.545 $X2=11.4 $Y2=2.8
r266 6 50 600 $w=1.7e-07 $l=2.995e-07 $layer=licon1_PDIFF $count=1 $X=10.32
+ $Y=2.48 $X2=10.48 $Y2=2.71
r267 5 46 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=8.215
+ $Y=1.895 $X2=8.34 $Y2=2.04
r268 4 42 600 $w=1.7e-07 $l=5.74565e-07 $layer=licon1_PDIFF $count=1 $X=7.02
+ $Y=2.315 $X2=7.24 $Y2=2.79
r269 3 38 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=4.69
+ $Y=1.835 $X2=4.83 $Y2=2.895
r270 2 34 600 $w=1.7e-07 $l=5.22303e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=2.455 $X2=2.94 $Y2=2.895
r271 1 30 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=2.455 $X2=1.185 $Y2=2.6
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%A_367_491# 1 2 3 4 5 18 20 23 26 27 28 32
+ 35 37 43 44
c127 20 0 9.68398e-20 $X=3.04 $Y=0.9
r128 47 48 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=5.905 $Y=2.52
+ $X2=5.905 $Y2=2.535
r129 44 47 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=5.905 $Y=2.24
+ $X2=5.905 $Y2=2.52
r130 41 43 19.9119 $w=1.93e-07 $l=3.15e-07 $layer=LI1_cond $X=3.125 $Y=2.502
+ $X2=3.44 $Y2=2.502
r131 37 39 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.15 $Y=0.7 $X2=2.15
+ $Y2=0.9
r132 30 32 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=6.43 $Y=2.155
+ $X2=6.43 $Y2=0.865
r133 29 44 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.035 $Y=2.24
+ $X2=5.905 $Y2=2.24
r134 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.345 $Y=2.24
+ $X2=6.43 $Y2=2.155
r135 28 29 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.345 $Y=2.24
+ $X2=6.035 $Y2=2.24
r136 27 43 10.634 $w=1.93e-07 $l=1.80748e-07 $layer=LI1_cond $X=3.605 $Y=2.535
+ $X2=3.44 $Y2=2.502
r137 26 48 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.775 $Y=2.535
+ $X2=5.905 $Y2=2.535
r138 26 27 141.572 $w=1.68e-07 $l=2.17e-06 $layer=LI1_cond $X=5.775 $Y=2.535
+ $X2=3.605 $Y2=2.535
r139 23 41 1.47909 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=3.125 $Y=2.385
+ $X2=3.125 $Y2=2.502
r140 22 23 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.125 $Y=0.985
+ $X2=3.125 $Y2=2.385
r141 21 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0.9
+ $X2=2.15 $Y2=0.9
r142 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.04 $Y=0.9
+ $X2=3.125 $Y2=0.985
r143 20 21 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.04 $Y=0.9
+ $X2=2.315 $Y2=0.9
r144 19 35 4.12218 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=2.502
+ $X2=1.975 $Y2=2.502
r145 18 41 4.83854 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=2.502
+ $X2=3.125 $Y2=2.502
r146 18 19 44.1361 $w=2.33e-07 $l=9e-07 $layer=LI1_cond $X=3.04 $Y=2.502
+ $X2=2.14 $Y2=2.502
r147 5 47 600 $w=1.7e-07 $l=2.89914e-07 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=2.315 $X2=5.94 $Y2=2.52
r148 4 43 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.3
+ $Y=2.455 $X2=3.44 $Y2=2.6
r149 3 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.835
+ $Y=2.455 $X2=1.975 $Y2=2.6
r150 2 32 182 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_NDIFF $count=1 $X=6.305
+ $Y=0.595 $X2=6.43 $Y2=0.865
r151 1 37 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.01
+ $Y=0.405 $X2=2.15 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%Q 1 2 7 8 9 10 11
r19 10 11 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=12.647 $Y=1.665
+ $X2=12.647 $Y2=2.035
r20 9 10 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=12.647 $Y=1.295
+ $X2=12.647 $Y2=1.665
r21 8 9 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=12.647 $Y=0.925
+ $X2=12.647 $Y2=1.295
r22 7 8 13.5287 $w=3.43e-07 $l=4.05e-07 $layer=LI1_cond $X=12.647 $Y=0.52
+ $X2=12.647 $Y2=0.925
r23 2 11 600 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=12.51
+ $Y=1.835 $X2=12.635 $Y2=2.12
r24 1 7 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=12.54
+ $Y=0.375 $X2=12.665 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%Q_N 1 2 7 8 9 10 11 12 13 25 31 54
r20 52 54 0.473607 $w=3.63e-07 $l=1.5e-08 $layer=LI1_cond $X=13.582 $Y=2.02
+ $X2=13.582 $Y2=2.035
r21 38 54 0.0631476 $w=3.63e-07 $l=2e-09 $layer=LI1_cond $X=13.582 $Y=2.037
+ $X2=13.582 $Y2=2.035
r22 23 31 2.02456 $w=3.68e-07 $l=6.5e-08 $layer=LI1_cond $X=13.58 $Y=0.99
+ $X2=13.58 $Y2=0.925
r23 13 45 4.26246 $w=3.63e-07 $l=1.35e-07 $layer=LI1_cond $X=13.582 $Y=2.775
+ $X2=13.582 $Y2=2.91
r24 12 13 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=13.582 $Y=2.405
+ $X2=13.582 $Y2=2.775
r25 11 52 0.852492 $w=3.63e-07 $l=2.7e-08 $layer=LI1_cond $X=13.582 $Y=1.993
+ $X2=13.582 $Y2=2.02
r26 11 50 7.32 $w=3.63e-07 $l=1.38e-07 $layer=LI1_cond $X=13.582 $Y=1.993
+ $X2=13.582 $Y2=1.855
r27 11 12 10.3246 $w=3.63e-07 $l=3.27e-07 $layer=LI1_cond $X=13.582 $Y=2.078
+ $X2=13.582 $Y2=2.405
r28 11 38 1.29453 $w=3.63e-07 $l=4.1e-08 $layer=LI1_cond $X=13.582 $Y=2.078
+ $X2=13.582 $Y2=2.037
r29 10 50 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=13.675 $Y=1.665
+ $X2=13.675 $Y2=1.855
r30 9 10 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=13.675 $Y=1.295
+ $X2=13.675 $Y2=1.665
r31 9 48 7.39394 $w=1.78e-07 $l=1.2e-07 $layer=LI1_cond $X=13.675 $Y=1.295
+ $X2=13.675 $Y2=1.175
r32 8 48 8.49656 $w=3.68e-07 $l=1.75e-07 $layer=LI1_cond $X=13.58 $Y=1 $X2=13.58
+ $Y2=1.175
r33 8 23 0.311471 $w=3.68e-07 $l=1e-08 $layer=LI1_cond $X=13.58 $Y=1 $X2=13.58
+ $Y2=0.99
r34 8 31 0.311471 $w=3.68e-07 $l=1e-08 $layer=LI1_cond $X=13.58 $Y=0.915
+ $X2=13.58 $Y2=0.925
r35 7 8 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=13.58 $Y=0.555
+ $X2=13.58 $Y2=0.915
r36 7 25 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=13.58 $Y=0.555
+ $X2=13.58 $Y2=0.52
r37 2 52 400 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=13.355
+ $Y=1.835 $X2=13.495 $Y2=2.02
r38 2 45 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=13.355
+ $Y=1.835 $X2=13.495 $Y2=2.91
r39 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.385
+ $Y=0.375 $X2=13.525 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 55 58 59 61 62 64 65 67 68 69 71 76 94 101 111 112 115 118 121 124
c140 112 0 3.56444e-20 $X=13.68 $Y=0
c141 31 0 1.47595e-19 $X=3.44 $Y=0.56
r142 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r143 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r144 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r145 115 116 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r146 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r147 109 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.68 $Y2=0
r148 109 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=11.76 $Y2=0
r149 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r150 106 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.875 $Y=0
+ $X2=11.71 $Y2=0
r151 106 108 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=11.875 $Y=0
+ $X2=12.72 $Y2=0
r152 105 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r153 105 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r154 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r155 102 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.465 $Y=0
+ $X2=10.3 $Y2=0
r156 102 104 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=10.465 $Y=0
+ $X2=11.28 $Y2=0
r157 101 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.545 $Y=0
+ $X2=11.71 $Y2=0
r158 101 104 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.545 $Y=0
+ $X2=11.28 $Y2=0
r159 100 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r160 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r161 97 100 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=9.84 $Y2=0
r162 96 99 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=9.84
+ $Y2=0
r163 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r164 94 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.135 $Y=0
+ $X2=10.3 $Y2=0
r165 94 99 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.135 $Y=0
+ $X2=9.84 $Y2=0
r166 93 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r167 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r168 89 92 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=0 $X2=7.92
+ $Y2=0
r169 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r170 87 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r171 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r172 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r173 84 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r174 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r175 81 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=0
+ $X2=3.44 $Y2=0
r176 81 83 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.605 $Y=0
+ $X2=4.56 $Y2=0
r177 80 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r178 80 116 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=0.72 $Y2=0
r179 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r180 77 115 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=0.69 $Y2=0
r181 77 79 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=3.12 $Y2=0
r182 76 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=0
+ $X2=3.44 $Y2=0
r183 76 79 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=0
+ $X2=3.12 $Y2=0
r184 74 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r185 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r186 71 115 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=0
+ $X2=0.69 $Y2=0
r187 71 73 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r188 69 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r189 69 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6
+ $Y2=0
r190 67 108 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12.99 $Y=0
+ $X2=12.72 $Y2=0
r191 67 68 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=12.99 $Y=0
+ $X2=13.107 $Y2=0
r192 66 111 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=13.225 $Y=0
+ $X2=13.68 $Y2=0
r193 66 68 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=13.225 $Y=0
+ $X2=13.107 $Y2=0
r194 64 92 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=7.95 $Y=0 $X2=7.92
+ $Y2=0
r195 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.95 $Y=0 $X2=8.115
+ $Y2=0
r196 63 96 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.28 $Y=0 $X2=8.4
+ $Y2=0
r197 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=0 $X2=8.115
+ $Y2=0
r198 61 86 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.655 $Y=0
+ $X2=5.52 $Y2=0
r199 61 62 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.655 $Y=0 $X2=5.745
+ $Y2=0
r200 60 89 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=0 $X2=6
+ $Y2=0
r201 60 62 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.745
+ $Y2=0
r202 58 83 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.665 $Y=0
+ $X2=4.56 $Y2=0
r203 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=0 $X2=4.83
+ $Y2=0
r204 57 86 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.995 $Y=0
+ $X2=5.52 $Y2=0
r205 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=0 $X2=4.83
+ $Y2=0
r206 53 68 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=13.107 $Y=0.085
+ $X2=13.107 $Y2=0
r207 53 55 20.3517 $w=2.33e-07 $l=4.15e-07 $layer=LI1_cond $X=13.107 $Y=0.085
+ $X2=13.107 $Y2=0.5
r208 49 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.71 $Y=0.085
+ $X2=11.71 $Y2=0
r209 49 51 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=11.71 $Y=0.085
+ $X2=11.71 $Y2=0.44
r210 45 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.3 $Y=0.085
+ $X2=10.3 $Y2=0
r211 45 47 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=10.3 $Y=0.085
+ $X2=10.3 $Y2=0.505
r212 41 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0
r213 41 43 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=8.115 $Y=0.085
+ $X2=8.115 $Y2=0.465
r214 37 62 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=0.085
+ $X2=5.745 $Y2=0
r215 37 39 43.7475 $w=1.78e-07 $l=7.1e-07 $layer=LI1_cond $X=5.745 $Y=0.085
+ $X2=5.745 $Y2=0.795
r216 33 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.83 $Y=0.085
+ $X2=4.83 $Y2=0
r217 33 35 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=4.83 $Y=0.085
+ $X2=4.83 $Y2=0.605
r218 29 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=0.085
+ $X2=3.44 $Y2=0
r219 29 31 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=3.44 $Y=0.085
+ $X2=3.44 $Y2=0.56
r220 25 115 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r221 25 27 22.974 $w=2.08e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.52
r222 8 55 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=12.955
+ $Y=0.375 $X2=13.095 $Y2=0.5
r223 7 51 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=11.585
+ $Y=0.235 $X2=11.71 $Y2=0.44
r224 6 47 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=10.16
+ $Y=0.34 $X2=10.3 $Y2=0.505
r225 5 43 182 $w=1.7e-07 $l=3.03109e-07 $layer=licon1_NDIFF $count=1 $X=7.87
+ $Y=0.595 $X2=8.115 $Y2=0.465
r226 4 39 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.595 $X2=5.75 $Y2=0.795
r227 3 35 182 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_NDIFF $count=1 $X=4.63
+ $Y=0.595 $X2=4.83 $Y2=0.605
r228 2 31 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.3
+ $Y=0.405 $X2=3.44 $Y2=0.56
r229 1 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.375 $X2=0.69 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_1%noxref_25 1 2 9 11 12 13
r33 13 16 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.94 $Y=0.34 $X2=2.94
+ $Y2=0.54
r34 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0.34
+ $X2=2.94 $Y2=0.34
r35 11 12 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=2.775 $Y=0.34
+ $X2=1.305 $Y2=0.34
r36 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.175 $Y=0.425
+ $X2=1.305 $Y2=0.34
r37 7 9 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.175 $Y=0.425
+ $X2=1.175 $Y2=0.57
r38 2 16 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.405 $X2=2.94 $Y2=0.54
r39 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.375 $X2=1.21 $Y2=0.57
.ends

