* File: sky130_fd_sc_lp__mux2_0.pex.spice
* Created: Wed Sep  2 09:59:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2_0%A_89_200# 1 2 9 13 15 16 17 20 21 23 24 27 30
+ 33 36
c78 23 0 1.05174e-19 $X=1.845 $Y=0.955
r79 38 39 5.20126 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.955
+ $X2=1.98 $Y2=1.04
r80 36 38 5.12197 $w=2.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.98 $Y=0.835
+ $X2=1.98 $Y2=0.955
r81 30 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=1.815
+ $X2=2.03 $Y2=1.9
r82 30 39 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.03 $Y=1.815
+ $X2=2.03 $Y2=1.04
r83 25 33 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.73 $Y=1.9 $X2=2.03
+ $Y2=1.9
r84 25 27 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=2.625
r85 23 38 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.845 $Y=0.955
+ $X2=1.98 $Y2=0.955
r86 23 24 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=1.845 $Y=0.955
+ $X2=0.78 $Y2=0.955
r87 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.165 $X2=0.61 $Y2=1.165
r88 18 24 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.652 $Y=1.04
+ $X2=0.78 $Y2=0.955
r89 18 20 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.652 $Y=1.04
+ $X2=0.652 $Y2=1.165
r90 16 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.61 $Y=1.505
+ $X2=0.61 $Y2=1.165
r91 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.505
+ $X2=0.61 $Y2=1.67
r92 15 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1 $X2=0.61
+ $Y2=1.165
r93 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.7 $Y=0.68 $X2=0.7
+ $Y2=1
r94 9 17 566.606 $w=1.5e-07 $l=1.105e-06 $layer=POLY_cond $X=0.52 $Y=2.775
+ $X2=0.52 $Y2=1.67
r95 2 27 600 $w=1.7e-07 $l=3.08504e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.455 $X2=1.73 $Y2=2.625
r96 1 36 182 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_NDIFF $count=1 $X=1.795
+ $Y=0.625 $X2=2.01 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_0%S 5 7 9 12 16 20 24 26 27 30 33 34 35 37 38
+ 39 40 41 42 48 51
c118 48 0 9.82229e-20 $X=3.3 $Y=1.745
c119 39 0 1.58325e-19 $X=2.805 $Y=2.405
c120 26 0 1.57021e-19 $X=3.3 $Y=2.25
r121 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.3
+ $Y=1.745 $X2=3.3 $Y2=1.745
r122 41 42 7.05836 $w=5.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.185 $Y=2.035
+ $X2=3.185 $Y2=2.32
r123 41 49 8.35521 $w=3.98e-07 $l=2.9e-07 $layer=LI1_cond $X=3.185 $Y=2.035
+ $X2=3.185 $Y2=1.745
r124 40 49 2.30489 $w=3.98e-07 $l=8e-08 $layer=LI1_cond $X=3.185 $Y=1.665
+ $X2=3.185 $Y2=1.745
r125 38 42 5.87433 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.985 $Y=2.405
+ $X2=3.185 $Y2=2.405
r126 38 39 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.985 $Y=2.405
+ $X2=2.805 $Y2=2.405
r127 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=2.49
+ $X2=2.805 $Y2=2.405
r128 36 37 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.72 $Y=2.49
+ $X2=2.72 $Y2=2.905
r129 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.635 $Y=2.99
+ $X2=2.72 $Y2=2.905
r130 34 35 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=2.635 $Y=2.99
+ $X2=1.33 $Y2=2.99
r131 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.245 $Y=2.905
+ $X2=1.33 $Y2=2.99
r132 32 33 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.245 $Y=2.265
+ $X2=1.245 $Y2=2.905
r133 30 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=2.13
+ $X2=0.97 $Y2=2.295
r134 30 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=2.13
+ $X2=0.97 $Y2=1.965
r135 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=2.13 $X2=0.97 $Y2=2.13
r136 27 32 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.16 $Y=2.155
+ $X2=1.245 $Y2=2.265
r137 27 29 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=1.16 $Y=2.155
+ $X2=0.97 $Y2=2.155
r138 25 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.3 $Y=2.085
+ $X2=3.3 $Y2=1.745
r139 25 26 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=2.085
+ $X2=3.3 $Y2=2.25
r140 24 48 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.3 $Y=1.73 $X2=3.3
+ $Y2=1.745
r141 23 24 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.285 $Y=1.58
+ $X2=3.285 $Y2=1.73
r142 18 20 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.06 $Y=1.075
+ $X2=1.21 $Y2=1.075
r143 16 26 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=3.295 $Y=2.785
+ $X2=3.295 $Y2=2.25
r144 12 23 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.18 $Y=0.835
+ $X2=3.18 $Y2=1.58
r145 7 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.21 $Y=1 $X2=1.21
+ $Y2=1.075
r146 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.21 $Y=1 $X2=1.21
+ $Y2=0.68
r147 5 52 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.06 $Y=2.665
+ $X2=1.06 $Y2=2.295
r148 1 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.06 $Y=1.15
+ $X2=1.06 $Y2=1.075
r149 1 51 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=1.06 $Y=1.15
+ $X2=1.06 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_0%A1 3 6 8 11 15 19 23 24 27
c59 23 0 1.00552e-19 $X=2.24 $Y=2.25
c60 8 0 4.32955e-20 $X=2.295 $Y=0.382
c61 6 0 5.77732e-20 $X=2.04 $Y=2.785
r62 24 27 6.63084 $w=3.98e-07 $l=9.5e-08 $layer=LI1_cond $X=2.265 $Y=2.25
+ $X2=2.265 $Y2=2.155
r63 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=2.25 $X2=2.24 $Y2=2.25
r64 20 23 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=2.04 $Y=2.25 $X2=2.24
+ $Y2=2.25
r65 15 24 4.46572 $w=3.98e-07 $l=1.55e-07 $layer=LI1_cond $X=2.265 $Y=2.405
+ $X2=2.265 $Y2=2.25
r66 13 27 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=2.38 $Y=0.5
+ $X2=2.38 $Y2=2.155
r67 11 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=0.35
+ $X2=1.81 $Y2=0.515
r68 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=0.35 $X2=1.81 $Y2=0.35
r69 8 13 7.04737 $w=2.35e-07 $l=1.54771e-07 $layer=LI1_cond $X=2.295 $Y=0.382
+ $X2=2.38 $Y2=0.5
r70 8 10 23.7845 $w=2.33e-07 $l=4.85e-07 $layer=LI1_cond $X=2.295 $Y=0.382
+ $X2=1.81 $Y2=0.382
r71 4 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=2.415
+ $X2=2.04 $Y2=2.25
r72 4 6 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.04 $Y=2.415 $X2=2.04
+ $Y2=2.785
r73 3 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.72 $Y=0.835
+ $X2=1.72 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_0%A0 3 6 7 11 15 17 18 26
c50 11 0 3.29812e-19 $X=2.26 $Y=0.835
c51 7 0 1.05174e-19 $X=2.185 $Y=1.49
r52 24 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.6 $Y=1.55
+ $X2=1.765 $Y2=1.55
r53 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.55 $X2=1.6 $Y2=1.55
r54 21 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.51 $Y=1.55 $X2=1.6
+ $Y2=1.55
r55 18 25 2.11944 $w=4.33e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=1.427 $X2=1.6
+ $Y2=1.427
r56 17 25 10.5972 $w=4.33e-07 $l=4e-07 $layer=LI1_cond $X=1.2 $Y=1.427 $X2=1.6
+ $Y2=1.427
r57 13 15 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.42 $Y=1.985 $X2=1.51
+ $Y2=1.985
r58 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.26 $Y=1.415
+ $X2=2.26 $Y2=0.835
r59 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.185 $Y=1.49
+ $X2=2.26 $Y2=1.415
r60 7 26 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.185 $Y=1.49
+ $X2=1.765 $Y2=1.49
r61 6 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.51 $Y=1.91 $X2=1.51
+ $Y2=1.985
r62 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.51 $Y=1.715
+ $X2=1.51 $Y2=1.55
r63 5 6 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.51 $Y=1.715
+ $X2=1.51 $Y2=1.91
r64 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.42 $Y=2.06 $X2=1.42
+ $Y2=1.985
r65 1 3 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=1.42 $Y=2.06 $X2=1.42
+ $Y2=2.665
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_0%A_509_99# 1 2 9 12 15 17 20 22 23 25 26 33
c62 25 0 4.28035e-19 $X=2.73 $Y=1.34
c63 9 0 4.32955e-20 $X=2.62 $Y=0.835
r64 31 33 5.76222 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=3.51 $Y=2.8 $X2=3.65
+ $Y2=2.8
r65 28 29 10.3341 $w=4.25e-07 $l=3.6e-07 $layer=LI1_cond $X=3.485 $Y=0.9
+ $X2=3.485 $Y2=1.26
r66 26 36 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.72 $Y=1.34
+ $X2=2.72 $Y2=1.175
r67 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.73
+ $Y=1.34 $X2=2.73 $Y2=1.34
r68 23 33 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.65 $Y=2.66 $X2=3.65
+ $Y2=2.8
r69 22 29 6.97754 $w=4.25e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.65 $Y=1.345
+ $X2=3.485 $Y2=1.26
r70 22 23 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=3.65 $Y=1.345
+ $X2=3.65 $Y2=2.66
r71 21 25 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.815 $Y=1.26 $X2=2.725
+ $Y2=1.26
r72 20 29 6.14847 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=3.235 $Y=1.26
+ $X2=3.485 $Y2=1.26
r73 20 21 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.235 $Y=1.26
+ $X2=2.815 $Y2=1.26
r74 15 17 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.69 $Y=2.785 $X2=2.69
+ $Y2=1.845
r75 12 17 40.1627 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.72 $Y=1.67
+ $X2=2.72 $Y2=1.845
r76 11 26 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=2.72 $Y=1.35 $X2=2.72
+ $Y2=1.34
r77 11 12 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.72 $Y=1.35
+ $X2=2.72 $Y2=1.67
r78 9 36 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.62 $Y=0.835 $X2=2.62
+ $Y2=1.175
r79 2 31 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=3.37
+ $Y=2.575 $X2=3.51 $Y2=2.775
r80 1 28 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.625 $X2=3.4 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_0%X 1 2 9 11 12 13 14 15 16 17 26 38
r25 39 48 0.808207 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=0.277 $Y=2.627
+ $X2=0.277 $Y2=2.6
r26 38 46 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=2.405 $X2=0.22
+ $Y2=2.435
r27 17 39 4.43017 $w=3.83e-07 $l=1.48e-07 $layer=LI1_cond $X=0.277 $Y=2.775
+ $X2=0.277 $Y2=2.627
r28 16 48 4.13083 $w=3.83e-07 $l=1.38e-07 $layer=LI1_cond $X=0.277 $Y=2.462
+ $X2=0.277 $Y2=2.6
r29 16 46 1.84985 $w=3.83e-07 $l=2.7e-08 $layer=LI1_cond $X=0.277 $Y=2.462
+ $X2=0.277 $Y2=2.435
r30 16 38 1.19513 $w=2.68e-07 $l=2.8e-08 $layer=LI1_cond $X=0.22 $Y=2.377
+ $X2=0.22 $Y2=2.405
r31 15 16 14.5976 $w=2.68e-07 $l=3.42e-07 $layer=LI1_cond $X=0.22 $Y=2.035
+ $X2=0.22 $Y2=2.377
r32 14 15 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=2.035
r33 13 14 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.665
r34 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.925
+ $X2=0.22 $Y2=1.295
r35 12 26 9.60369 $w=2.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.22 $Y=0.925
+ $X2=0.22 $Y2=0.7
r36 11 26 3.16176 $w=2.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.22 $Y=0.585
+ $X2=0.22 $Y2=0.7
r37 7 11 3.71163 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=0.355 $Y=0.585
+ $X2=0.22 $Y2=0.585
r38 7 9 6.51381 $w=2.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.355 $Y=0.585
+ $X2=0.485 $Y2=0.585
r39 2 48 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.18
+ $Y=2.455 $X2=0.305 $Y2=2.6
r40 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.34
+ $Y=0.47 $X2=0.485 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_0%VPWR 1 2 11 15 18 19 20 30 31 34
c43 15 0 1.57021e-19 $X=3.08 $Y=2.825
r44 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r46 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 22 34 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.815 $Y2=3.33
r52 22 24 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 18 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 18 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.975 $Y=3.33 $X2=3.075
+ $Y2=3.33
r57 17 30 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 17 19 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.175 $Y=3.33 $X2=3.075
+ $Y2=3.33
r59 13 19 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=3.245
+ $X2=3.075 $Y2=3.33
r60 13 15 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=3.075 $Y=3.245
+ $X2=3.075 $Y2=2.825
r61 9 34 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r62 9 11 20.9086 $w=3.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.61
r63 2 15 600 $w=1.7e-07 $l=4.21871e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=2.575 $X2=3.08 $Y2=2.825
r64 1 11 300 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.455 $X2=0.845 $Y2=2.61
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_0%VGND 1 2 9 13 16 17 19 20 21 34 35
r40 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r41 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r42 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r44 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r46 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 21 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r48 21 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r49 19 31 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.64
+ $Y2=0
r50 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.9
+ $Y2=0
r51 18 34 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=3.6
+ $Y2=0
r52 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=2.9
+ $Y2=0
r53 16 24 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.72
+ $Y2=0
r54 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.995
+ $Y2=0
r55 15 28 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.2
+ $Y2=0
r56 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=0.995
+ $Y2=0
r57 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=0.085 $X2=2.9
+ $Y2=0
r58 11 13 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=2.9 $Y=0.085 $X2=2.9
+ $Y2=0.82
r59 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.995 $Y=0.085
+ $X2=0.995 $Y2=0
r60 7 9 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.995 $Y=0.085
+ $X2=0.995 $Y2=0.595
r61 2 13 182 $w=1.7e-07 $l=2.86356e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.625 $X2=2.9 $Y2=0.82
r62 1 9 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.47 $X2=0.995 $Y2=0.595
.ends

