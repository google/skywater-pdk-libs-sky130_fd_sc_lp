* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a221o_lp A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_322_419# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VGND C1 a_764_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_545_400# B1 a_322_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_162_66# a_96_183# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND A2 a_336_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_545_400# C1 a_96_183# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_336_66# A1 a_96_183# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR A2 a_322_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_322_419# B2 a_545_400# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_582_66# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 X a_96_183# a_162_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_96_183# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_764_66# C1 a_96_183# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_96_183# B1 a_582_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
