* File: sky130_fd_sc_lp__sdfrtp_lp2.pex.spice
* Created: Fri Aug 28 11:28:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_81_194# 1 2 9 12 14 18 19 21 25 28 31
+ 33 34 35 39 42
c113 39 0 1.06473e-19 $X=4.14 $Y=2.2
c114 25 0 2.94669e-20 $X=3.985 $Y=0.76
c115 12 0 2.78071e-21 $X=2.59 $Y=2.595
r116 37 39 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=4 $Y=2.2 $X2=4.14
+ $Y2=2.2
r117 31 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.135
+ $X2=0.57 $Y2=0.97
r118 30 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=1.135
+ $X2=0.735 $Y2=1.135
r119 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.57
+ $Y=1.135 $X2=0.57 $Y2=1.135
r120 28 39 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.14 $Y=2.075
+ $X2=4.14 $Y2=2.2
r121 27 35 3.27229 $w=2.87e-07 $l=1.54771e-07 $layer=LI1_cond $X=4.14 $Y=1.27
+ $X2=4.022 $Y2=1.185
r122 27 28 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=4.14 $Y=1.27
+ $X2=4.14 $Y2=2.075
r123 23 35 3.27229 $w=2.87e-07 $l=8.5e-08 $layer=LI1_cond $X=4.022 $Y=1.1
+ $X2=4.022 $Y2=1.185
r124 23 25 9.67483 $w=4.03e-07 $l=3.4e-07 $layer=LI1_cond $X=4.022 $Y=1.1
+ $X2=4.022 $Y2=0.76
r125 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.765 $Y=1.185
+ $X2=2.6 $Y2=1.185
r126 21 35 3.2872 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=3.82 $Y=1.185
+ $X2=4.022 $Y2=1.185
r127 21 22 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=3.82 $Y=1.185
+ $X2=2.765 $Y2=1.185
r128 19 46 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.615
+ $X2=2.6 $Y2=1.78
r129 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.6
+ $Y=1.615 $X2=2.6 $Y2=1.615
r130 16 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=1.27 $X2=2.6
+ $Y2=1.185
r131 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.6 $Y=1.27
+ $X2=2.6 $Y2=1.615
r132 14 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.435 $Y=1.185
+ $X2=2.6 $Y2=1.185
r133 14 33 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=2.435 $Y=1.185
+ $X2=0.735 $Y2=1.185
r134 12 46 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.59 $Y=2.595
+ $X2=2.59 $Y2=1.78
r135 9 42 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.63 $Y=0.65
+ $X2=0.63 $Y2=0.97
r136 2 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=2.095 $X2=4 $Y2=2.24
r137 1 25 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.845
+ $Y=0.595 $X2=3.985 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%D 1 3 6 8
c33 8 0 3.60011e-19 $X=0.72 $Y=1.665
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.74
+ $Y=1.675 $X2=0.74 $Y2=1.675
r35 4 11 39.2698 $w=3.83e-07 $l=2.43926e-07 $layer=POLY_cond $X=1.02 $Y=1.51
+ $X2=0.845 $Y2=1.675
r36 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.02 $Y=1.51 $X2=1.02
+ $Y2=0.65
r37 1 11 49.8545 $w=3.83e-07 $l=4.16233e-07 $layer=POLY_cond $X=0.99 $Y=2.025
+ $X2=0.845 $Y2=1.675
r38 1 3 109.896 $w=2.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.99 $Y=2.025 $X2=0.99
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%SCE 3 6 8 10 15 17 19 23 25 28 29 31 34
+ 37 39 45
c107 34 0 1.66642e-19 $X=1.52 $Y=1.77
c108 29 0 2.41669e-19 $X=3.71 $Y=1.72
c109 6 0 1.93369e-19 $X=1.61 $Y=0.65
r110 35 45 10.0259 $w=5.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=1.84
+ $X2=1.685 $Y2=1.84
r111 34 37 47.2437 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.52 $Y=1.77
+ $X2=1.52 $Y2=2.02
r112 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.77
+ $X2=1.52 $Y2=1.605
r113 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.77 $X2=1.52 $Y2=1.77
r114 31 35 6.59905 $w=5.78e-07 $l=3.2e-07 $layer=LI1_cond $X=1.2 $Y=1.84
+ $X2=1.52 $Y2=1.84
r115 29 40 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.72
+ $X2=3.71 $Y2=1.885
r116 29 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.72
+ $X2=3.71 $Y2=1.555
r117 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.71
+ $Y=1.72 $X2=3.71 $Y2=1.72
r118 25 28 13.3953 $w=2.96e-07 $l=4.11096e-07 $layer=LI1_cond $X=3.485 $Y=2.045
+ $X2=3.68 $Y2=1.72
r119 25 45 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=3.485 $Y=2.045
+ $X2=1.685 $Y2=2.045
r120 22 23 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.62 $Y=1.165
+ $X2=3.77 $Y2=1.165
r121 20 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.41 $Y=1.165
+ $X2=3.62 $Y2=1.165
r122 17 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=1.09
+ $X2=3.77 $Y2=1.165
r123 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.77 $Y=1.09
+ $X2=3.77 $Y2=0.805
r124 15 40 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.735 $Y=2.595
+ $X2=3.735 $Y2=1.885
r125 11 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.62 $Y=1.24
+ $X2=3.62 $Y2=1.165
r126 11 39 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=3.62 $Y=1.24
+ $X2=3.62 $Y2=1.555
r127 8 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.09
+ $X2=3.41 $Y2=1.165
r128 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.41 $Y=1.09 $X2=3.41
+ $Y2=0.805
r129 6 36 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=1.61 $Y=0.65
+ $X2=1.61 $Y2=1.605
r130 3 37 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.48 $Y=2.595
+ $X2=1.48 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%SCD 3 7 9 12
c35 3 0 1.2046e-19 $X=2 $Y=0.65
r36 12 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.615
+ $X2=2.06 $Y2=1.78
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.06 $Y=1.615
+ $X2=2.06 $Y2=1.45
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=1.615 $X2=2.06 $Y2=1.615
r39 9 13 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.16 $Y=1.615 $X2=2.06
+ $Y2=1.615
r40 7 15 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.07 $Y=2.595
+ $X2=2.07 $Y2=1.78
r41 3 14 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2 $Y=0.65 $X2=2
+ $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%CLK 3 7 11 13 18
c38 13 0 4.72961e-20 $X=5.04 $Y=1.295
r39 18 20 14.412 $w=3.01e-07 $l=9e-08 $layer=POLY_cond $X=4.99 $Y=1.335 $X2=5.08
+ $Y2=1.335
r40 16 18 22.4186 $w=3.01e-07 $l=1.4e-07 $layer=POLY_cond $X=4.85 $Y=1.335
+ $X2=4.99 $Y2=1.335
r41 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.335 $X2=4.99 $Y2=1.335
r42 9 20 19.0468 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.08 $Y=1.17
+ $X2=5.08 $Y2=1.335
r43 9 11 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=5.08 $Y=1.17 $X2=5.08
+ $Y2=0.805
r44 5 16 7.2153 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.5 $X2=4.85
+ $Y2=1.335
r45 5 7 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=4.85 $Y=1.5 $X2=4.85
+ $Y2=2.54
r46 1 16 20.8173 $w=3.01e-07 $l=2.20624e-07 $layer=POLY_cond $X=4.72 $Y=1.17
+ $X2=4.85 $Y2=1.335
r47 1 3 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=4.72 $Y=1.17 $X2=4.72
+ $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_1147_408# 1 2 7 9 11 12 14 17 18 21 22
+ 23 24 26 29 31 34 38 39 41 42 45 57 60 67 68
c174 60 0 1.47992e-19 $X=6.6 $Y=1.555
c175 45 0 1.02141e-19 $X=10.295 $Y=0.93
c176 39 0 1.46627e-19 $X=7.64 $Y=1.29
c177 38 0 2.22113e-19 $X=7.64 $Y=1.29
c178 12 0 1.31384e-19 $X=7.73 $Y=1.125
r179 67 68 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.295 $Y=0.805
+ $X2=10.295 $Y2=0.73
r180 58 60 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.6 $Y=1.615 $X2=6.6
+ $Y2=1.555
r181 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.6
+ $Y=1.615 $X2=6.6 $Y2=1.615
r182 46 67 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=10.295 $Y=0.93
+ $X2=10.295 $Y2=0.805
r183 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.295
+ $Y=0.93 $X2=10.295 $Y2=0.93
r184 43 45 7.23627 $w=2.13e-07 $l=1.35e-07 $layer=LI1_cond $X=10.317 $Y=0.795
+ $X2=10.317 $Y2=0.93
r185 41 43 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=10.21 $Y=0.71
+ $X2=10.317 $Y2=0.795
r186 41 42 162.123 $w=1.68e-07 $l=2.485e-06 $layer=LI1_cond $X=10.21 $Y=0.71
+ $X2=7.725 $Y2=0.71
r187 39 66 10.3286 $w=4.2e-07 $l=9e-08 $layer=POLY_cond $X=7.64 $Y=1.392
+ $X2=7.73 $Y2=1.392
r188 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.64
+ $Y=1.29 $X2=7.64 $Y2=1.29
r189 36 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.64 $Y=0.795
+ $X2=7.725 $Y2=0.71
r190 36 38 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.64 $Y=0.795
+ $X2=7.64 $Y2=1.29
r191 32 57 11.8038 $w=3.28e-07 $l=3.38e-07 $layer=LI1_cond $X=6.262 $Y=1.615
+ $X2=6.6 $Y2=1.615
r192 32 53 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.262 $Y=1.615
+ $X2=6.132 $Y2=1.615
r193 32 34 19.7562 $w=3.83e-07 $l=6.6e-07 $layer=LI1_cond $X=6.262 $Y=1.45
+ $X2=6.262 $Y2=0.79
r194 31 49 11.8471 $w=2.48e-07 $l=2.57e-07 $layer=LI1_cond $X=6.132 $Y=2.155
+ $X2=5.875 $Y2=2.155
r195 30 53 1.01705 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=6.132 $Y=1.78
+ $X2=6.132 $Y2=1.615
r196 30 31 9.14637 $w=3.13e-07 $l=2.5e-07 $layer=LI1_cond $X=6.132 $Y=1.78
+ $X2=6.132 $Y2=2.03
r197 27 29 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.86 $Y=1.63
+ $X2=11.86 $Y2=1.87
r198 24 29 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=11.81 $Y=1.995
+ $X2=11.81 $Y2=1.87
r199 24 26 115.68 $w=2.5e-07 $l=6e-07 $layer=POLY_cond $X=11.81 $Y=1.995
+ $X2=11.81 $Y2=2.595
r200 22 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.785 $Y=1.555
+ $X2=11.86 $Y2=1.63
r201 22 23 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=11.785 $Y=1.555
+ $X2=11.605 $Y2=1.555
r202 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.53 $Y=1.48
+ $X2=11.605 $Y2=1.555
r203 20 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=11.53 $Y=0.88
+ $X2=11.53 $Y2=1.48
r204 19 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.46 $Y=0.805
+ $X2=10.295 $Y2=0.805
r205 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.455 $Y=0.805
+ $X2=11.53 $Y2=0.88
r206 18 19 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=11.455 $Y=0.805
+ $X2=10.46 $Y2=0.805
r207 17 68 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.385 $Y=0.445
+ $X2=10.385 $Y2=0.73
r208 12 66 27.059 $w=1.5e-07 $l=2.67e-07 $layer=POLY_cond $X=7.73 $Y=1.125
+ $X2=7.73 $Y2=1.392
r209 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.73 $Y=1.125
+ $X2=7.73 $Y2=0.805
r210 9 39 32.1333 $w=4.2e-07 $l=3.91714e-07 $layer=POLY_cond $X=7.36 $Y=1.66
+ $X2=7.64 $Y2=1.392
r211 9 11 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.36 $Y=1.66
+ $X2=7.36 $Y2=2.235
r212 8 60 13.3611 $w=2.1e-07 $l=1.65e-07 $layer=POLY_cond $X=6.765 $Y=1.555
+ $X2=6.6 $Y2=1.555
r213 7 9 26.3872 $w=4.2e-07 $l=1.69558e-07 $layer=POLY_cond $X=7.235 $Y=1.555
+ $X2=7.36 $Y2=1.66
r214 7 8 148.42 $w=2.1e-07 $l=4.7e-07 $layer=POLY_cond $X=7.235 $Y=1.555
+ $X2=6.765 $Y2=1.555
r215 2 49 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=2.04 $X2=5.875 $Y2=2.195
r216 1 34 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=6.105
+ $Y=0.595 $X2=6.245 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_1605_93# 1 2 7 9 12 14 15 18 19 21 22
+ 23 27 30 35 37 41 43 44
c124 44 0 9.28545e-20 $X=10.812 $Y=1.685
c125 22 0 5.71004e-20 $X=8.555 $Y=1.06
c126 21 0 1.52796e-19 $X=9.87 $Y=1.06
c127 19 0 6.11131e-20 $X=8.44 $Y=1.29
r128 43 44 8.71334 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=10.812 $Y=1.85
+ $X2=10.812 $Y2=1.685
r129 37 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=9.955 $Y=1.06
+ $X2=9.955 $Y2=1.36
r130 33 43 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=10.812 $Y=1.892
+ $X2=10.812 $Y2=1.85
r131 33 35 18.5502 $w=4.13e-07 $l=6.68e-07 $layer=LI1_cond $X=10.812 $Y=1.892
+ $X2=10.812 $Y2=2.56
r132 31 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.69 $Y=1.445
+ $X2=10.69 $Y2=1.36
r133 31 44 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.69 $Y=1.445
+ $X2=10.69 $Y2=1.685
r134 30 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.69 $Y=1.275
+ $X2=10.69 $Y2=1.36
r135 29 30 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=10.69 $Y=0.445
+ $X2=10.69 $Y2=1.275
r136 28 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.04 $Y=1.36
+ $X2=9.955 $Y2=1.36
r137 27 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.605 $Y=1.36
+ $X2=10.69 $Y2=1.36
r138 27 28 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=10.605 $Y=1.36
+ $X2=10.04 $Y2=1.36
r139 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.605 $Y=0.36
+ $X2=10.69 $Y2=0.445
r140 23 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=10.605 $Y=0.36
+ $X2=10.17 $Y2=0.36
r141 21 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.87 $Y=1.06
+ $X2=9.955 $Y2=1.06
r142 21 22 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=9.87 $Y=1.06
+ $X2=8.555 $Y2=1.06
r143 19 47 8.00664 $w=3.01e-07 $l=5e-08 $layer=POLY_cond $X=8.44 $Y=1.29
+ $X2=8.49 $Y2=1.29
r144 19 45 54.4452 $w=3.01e-07 $l=3.4e-07 $layer=POLY_cond $X=8.44 $Y=1.29
+ $X2=8.1 $Y2=1.29
r145 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.44
+ $Y=1.29 $X2=8.44 $Y2=1.29
r146 16 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.39 $Y=1.145
+ $X2=8.555 $Y2=1.06
r147 16 18 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.39 $Y=1.145
+ $X2=8.39 $Y2=1.29
r148 12 15 31.5625 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=8.5 $Y=1.73
+ $X2=8.5 $Y2=1.605
r149 12 14 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.5 $Y=1.73 $X2=8.5
+ $Y2=2.235
r150 10 47 9.14644 $w=2.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.49 $Y=1.455
+ $X2=8.49 $Y2=1.29
r151 10 15 41.851 $w=2.3e-07 $l=1.5e-07 $layer=POLY_cond $X=8.49 $Y=1.455
+ $X2=8.49 $Y2=1.605
r152 7 45 19.0468 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.1 $Y=1.125
+ $X2=8.1 $Y2=1.29
r153 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.1 $Y=1.125 $X2=8.1
+ $Y2=0.805
r154 2 43 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=10.635
+ $Y=1.705 $X2=10.855 $Y2=1.85
r155 2 35 400 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=10.635
+ $Y=1.705 $X2=10.855 $Y2=2.56
r156 1 25 182 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_NDIFF $count=1 $X=9.89
+ $Y=0.235 $X2=10.17 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%RESET_B 4 5 6 7 8 13 18 20 21 23 27 31 33
+ 35 39 42 43 45 46 47 48 56 59 60 61 65 78
c267 43 0 8.70527e-20 $X=13.32 $Y=1.77
c268 21 0 7.98625e-20 $X=9.03 $Y=1.575
c269 7 0 2.94669e-20 $X=2.975 $Y=1.165
r270 75 78 6.54083 $w=2.33e-07 $l=1.15e-07 $layer=LI1_cond $X=12.72 $Y=1.667
+ $X2=12.835 $Y2=1.667
r271 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.995
+ $Y=1.41 $X2=8.995 $Y2=1.41
r272 59 62 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.14 $Y=1.615
+ $X2=3.14 $Y2=1.78
r273 59 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.14 $Y=1.615
+ $X2=3.14 $Y2=1.45
r274 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.14
+ $Y=1.615 $X2=3.14 $Y2=1.615
r275 56 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=1.665
+ $X2=12.72 $Y2=1.665
r276 55 65 7.23488 $w=4.3e-07 $l=2.55e-07 $layer=LI1_cond $X=8.982 $Y=1.665
+ $X2=8.982 $Y2=1.41
r277 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.665
r278 50 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r279 48 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.025 $Y=1.665
+ $X2=8.88 $Y2=1.665
r280 47 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.575 $Y=1.665
+ $X2=12.72 $Y2=1.665
r281 47 48 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=12.575 $Y=1.665
+ $X2=9.025 $Y2=1.665
r282 46 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r283 45 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=8.88 $Y2=1.665
r284 45 46 6.76979 $w=1.4e-07 $l=5.47e-06 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=3.265 $Y2=1.665
r285 43 68 31.8564 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=13.337 $Y=1.77
+ $X2=13.337 $Y2=1.935
r286 43 67 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=13.337 $Y=1.77
+ $X2=13.337 $Y2=1.605
r287 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.32
+ $Y=1.77 $X2=13.32 $Y2=1.77
r288 39 42 2.01678 $w=3.98e-07 $l=7e-08 $layer=LI1_cond $X=13.285 $Y=1.7
+ $X2=13.285 $Y2=1.77
r289 35 39 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=13.085 $Y=1.7
+ $X2=13.285 $Y2=1.7
r290 35 78 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.085 $Y=1.7
+ $X2=12.835 $Y2=1.7
r291 31 68 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.395 $Y=2.595
+ $X2=13.395 $Y2=1.935
r292 27 67 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=13.23 $Y=0.445
+ $X2=13.23 $Y2=1.605
r293 21 64 27.0909 $w=3.28e-07 $l=1.81659e-07 $layer=POLY_cond $X=9.03 $Y=1.575
+ $X2=8.995 $Y2=1.41
r294 21 23 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.03 $Y=1.575
+ $X2=9.03 $Y2=2.235
r295 20 64 30.3239 $w=3.28e-07 $l=2.0994e-07 $layer=POLY_cond $X=8.985 $Y=1.205
+ $X2=8.995 $Y2=1.41
r296 19 33 88.7014 $w=1.44e-07 $l=2.65e-07 $layer=POLY_cond $X=8.985 $Y=0.9
+ $X2=8.72 $Y2=0.9
r297 19 20 42.8128 $w=3.1e-07 $l=2.3e-07 $layer=POLY_cond $X=8.985 $Y=0.975
+ $X2=8.985 $Y2=1.205
r298 16 33 1.84115 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.72 $Y=0.825
+ $X2=8.72 $Y2=0.9
r299 16 18 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.72 $Y=0.825
+ $X2=8.72 $Y2=0.54
r300 15 18 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.72 $Y=0.255
+ $X2=8.72 $Y2=0.54
r301 13 62 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=3.12 $Y=2.595
+ $X2=3.12 $Y2=1.78
r302 9 61 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.05 $Y=1.24
+ $X2=3.05 $Y2=1.45
r303 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.975 $Y=1.165
+ $X2=3.05 $Y2=1.24
r304 7 8 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.975 $Y=1.165 $X2=2.505
+ $Y2=1.165
r305 5 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.645 $Y=0.18
+ $X2=8.72 $Y2=0.255
r306 5 6 3148.38 $w=1.5e-07 $l=6.14e-06 $layer=POLY_cond $X=8.645 $Y=0.18
+ $X2=2.505 $Y2=0.18
r307 2 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.43 $Y=1.09
+ $X2=2.505 $Y2=1.165
r308 2 4 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.43 $Y=1.09 $X2=2.43
+ $Y2=0.65
r309 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.43 $Y=0.255
+ $X2=2.505 $Y2=0.18
r310 1 4 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.43 $Y=0.255
+ $X2=2.43 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_1432_119# 1 2 3 10 12 15 16 17 20 24 28
+ 32 34 36 38 42 43 46
c113 43 0 1.02141e-19 $X=9.535 $Y=1.41
c114 34 0 7.98625e-20 $X=9.275 $Y=2.045
c115 24 0 1.95202e-19 $X=9.62 $Y=0.925
c116 16 0 3.6571e-20 $X=10.385 $Y=1.5
r117 50 51 5.33952 $w=3.77e-07 $l=1.65e-07 $layer=LI1_cond $X=9.487 $Y=1.88
+ $X2=9.487 $Y2=2.045
r118 46 48 3.43222 $w=5.73e-07 $l=1.65e-07 $layer=LI1_cond $X=7.502 $Y=1.88
+ $X2=7.502 $Y2=2.045
r119 46 47 8.43332 $w=5.73e-07 $l=9e-08 $layer=LI1_cond $X=7.502 $Y=1.88
+ $X2=7.502 $Y2=1.79
r120 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.535
+ $Y=1.41 $X2=9.535 $Y2=1.41
r121 40 50 5.56084 $w=3.77e-07 $l=1.8747e-07 $layer=LI1_cond $X=9.535 $Y=1.715
+ $X2=9.487 $Y2=1.88
r122 40 42 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=9.535 $Y=1.715
+ $X2=9.535 $Y2=1.41
r123 36 51 2.62512 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=9.487 $Y=2.13
+ $X2=9.487 $Y2=2.045
r124 36 38 2.84721 $w=4.23e-07 $l=1.05e-07 $layer=LI1_cond $X=9.487 $Y=2.13
+ $X2=9.487 $Y2=2.235
r125 35 48 8.04321 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=7.79 $Y=2.045
+ $X2=7.502 $Y2=2.045
r126 34 51 5.41993 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=9.275 $Y=2.045
+ $X2=9.487 $Y2=2.045
r127 34 35 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=9.275 $Y=2.045
+ $X2=7.79 $Y2=2.045
r128 30 48 1.76812 $w=5.73e-07 $l=8.5e-08 $layer=LI1_cond $X=7.502 $Y=2.13
+ $X2=7.502 $Y2=2.045
r129 30 32 2.18414 $w=5.73e-07 $l=1.05e-07 $layer=LI1_cond $X=7.502 $Y=2.13
+ $X2=7.502 $Y2=2.235
r130 28 47 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=7.3 $Y=0.79 $X2=7.3
+ $Y2=1.79
r131 25 43 1.54335 $w=5.2e-07 $l=1.5e-08 $layer=POLY_cond $X=9.63 $Y=1.425
+ $X2=9.63 $Y2=1.41
r132 24 43 49.9018 $w=5.2e-07 $l=4.85e-07 $layer=POLY_cond $X=9.63 $Y=0.925
+ $X2=9.63 $Y2=1.41
r133 18 20 156.526 $w=2.5e-07 $l=6.3e-07 $layer=POLY_cond $X=10.51 $Y=1.575
+ $X2=10.51 $Y2=2.205
r134 17 25 39.3537 $w=1.5e-07 $l=2.95127e-07 $layer=POLY_cond $X=9.89 $Y=1.5
+ $X2=9.63 $Y2=1.425
r135 16 18 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=10.385 $Y=1.5
+ $X2=10.51 $Y2=1.575
r136 16 17 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.385 $Y=1.5
+ $X2=9.89 $Y2=1.5
r137 10 24 29.5599 $w=5.2e-07 $l=1.95e-07 $layer=POLY_cond $X=9.62 $Y=0.73
+ $X2=9.62 $Y2=0.925
r138 10 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.815 $Y=0.73
+ $X2=9.815 $Y2=0.445
r139 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.425 $Y=0.73
+ $X2=9.425 $Y2=0.445
r140 3 50 600 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_PDIFF $count=1 $X=9.155
+ $Y=1.735 $X2=9.44 $Y2=1.88
r141 3 38 300 $w=1.7e-07 $l=6.26498e-07 $layer=licon1_PDIFF $count=2 $X=9.155
+ $Y=1.735 $X2=9.44 $Y2=2.235
r142 2 46 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.485
+ $Y=1.735 $X2=7.625 $Y2=1.88
r143 2 32 300 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=2 $X=7.485
+ $Y=1.735 $X2=7.625 $Y2=2.235
r144 1 28 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=0.595 $X2=7.3 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_876_119# 1 2 9 11 13 17 19 20 22 23 24
+ 26 29 31 36 39 41 44 48 50 54 55 57 60 62 64 65
c184 65 0 1.64983e-19 $X=11.98 $Y=1.075
c185 60 0 9.28545e-20 $X=11.08 $Y=1.285
c186 57 0 3.6571e-20 $X=11.815 $Y=1.285
c187 54 0 9.9346e-20 $X=5.64 $Y=1.345
c188 50 0 4.86458e-20 $X=5.475 $Y=1.765
c189 13 0 4.72961e-20 $X=5.67 $Y=0.805
c190 9 0 5.74786e-20 $X=5.61 $Y=2.54
r191 65 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.98 $Y=1.075
+ $X2=11.98 $Y2=0.91
r192 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.98
+ $Y=1.075 $X2=11.98 $Y2=1.075
r193 60 73 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.08 $Y=1.285
+ $X2=11.08 $Y2=1.45
r194 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.08
+ $Y=1.285 $X2=11.08 $Y2=1.285
r195 57 64 8.34528 $w=2.88e-07 $l=2.1e-07 $layer=LI1_cond $X=11.96 $Y=1.285
+ $X2=11.96 $Y2=1.075
r196 57 59 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=11.815 $Y=1.285
+ $X2=11.08 $Y2=1.285
r197 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.64
+ $Y=1.345 $X2=5.64 $Y2=1.345
r198 52 54 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.64 $Y=1.68
+ $X2=5.64 $Y2=1.345
r199 51 62 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.67 $Y=1.765
+ $X2=4.545 $Y2=1.765
r200 50 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.475 $Y=1.765
+ $X2=5.64 $Y2=1.68
r201 50 51 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=5.475 $Y=1.765
+ $X2=4.67 $Y2=1.765
r202 46 62 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=1.85
+ $X2=4.545 $Y2=1.765
r203 46 48 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.545 $Y=1.85
+ $X2=4.545 $Y2=2.185
r204 42 62 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.505 $Y=1.68
+ $X2=4.545 $Y2=1.765
r205 42 44 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=4.505 $Y=1.68
+ $X2=4.505 $Y2=0.805
r206 39 75 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.92 $Y=0.445
+ $X2=11.92 $Y2=0.91
r207 36 73 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=11.12 $Y=2.205
+ $X2=11.12 $Y2=1.45
r208 34 36 216.155 $w=2.5e-07 $l=8.7e-07 $layer=POLY_cond $X=11.12 $Y=3.075
+ $X2=11.12 $Y2=2.205
r209 32 41 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=8.165 $Y=3.15
+ $X2=8.04 $Y2=3.15
r210 31 34 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=10.995 $Y=3.15
+ $X2=11.12 $Y2=3.075
r211 31 32 1451.13 $w=1.5e-07 $l=2.83e-06 $layer=POLY_cond $X=10.995 $Y=3.15
+ $X2=8.165 $Y2=3.15
r212 27 41 1.63566 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.04 $Y=3.075
+ $X2=8.04 $Y2=3.15
r213 27 29 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.04 $Y=3.075
+ $X2=8.04 $Y2=2.235
r214 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.085 $Y=1.09
+ $X2=7.085 $Y2=0.805
r215 22 41 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=7.915 $Y=3.15
+ $X2=8.04 $Y2=3.15
r216 22 23 866.574 $w=1.5e-07 $l=1.69e-06 $layer=POLY_cond $X=7.915 $Y=3.15
+ $X2=6.225 $Y2=3.15
r217 21 55 12.5195 $w=6.93e-07 $l=4.56207e-07 $layer=POLY_cond $X=6.225 $Y=1.165
+ $X2=5.85 $Y2=1.345
r218 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.01 $Y=1.165
+ $X2=7.085 $Y2=1.09
r219 20 21 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=7.01 $Y=1.165
+ $X2=6.225 $Y2=1.165
r220 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.15 $Y=3.075
+ $X2=6.225 $Y2=3.15
r221 18 55 74.1003 $w=3.46e-07 $l=6.37593e-07 $layer=POLY_cond $X=6.15 $Y=1.85
+ $X2=5.85 $Y2=1.345
r222 18 19 628.138 $w=1.5e-07 $l=1.225e-06 $layer=POLY_cond $X=6.15 $Y=1.85
+ $X2=6.15 $Y2=3.075
r223 11 21 40.8047 $w=6.93e-07 $l=2.29456e-07 $layer=POLY_cond $X=6.03 $Y=1.09
+ $X2=6.225 $Y2=1.165
r224 11 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.03 $Y=1.09
+ $X2=6.03 $Y2=0.805
r225 11 13 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=5.67 $Y=1.18
+ $X2=5.67 $Y2=0.805
r226 7 55 71.076 $w=3.46e-07 $l=6.13372e-07 $layer=POLY_cond $X=5.61 $Y=1.85
+ $X2=5.85 $Y2=1.345
r227 7 9 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.61 $Y=1.85 $X2=5.61
+ $Y2=2.54
r228 2 48 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=4.44
+ $Y=2.04 $X2=4.585 $Y2=2.185
r229 1 44 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.595 $X2=4.505 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_2435_296# 1 2 9 13 20 26 30 33 34 35 37
+ 38 39 41
c97 13 0 3.96307e-21 $X=12.46 $Y=0.445
r98 37 38 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=13.665 $Y=2.28
+ $X2=13.665 $Y2=2.115
r99 34 35 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=13.015 $Y=1.237
+ $X2=13.185 $Y2=1.237
r100 32 33 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=14.11 $Y=0.51
+ $X2=14.11 $Y2=1.265
r101 31 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.835 $Y=1.35
+ $X2=13.75 $Y2=1.35
r102 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.025 $Y=1.35
+ $X2=14.11 $Y2=1.265
r103 30 31 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=14.025 $Y=1.35
+ $X2=13.835 $Y2=1.35
r104 26 32 6.93832 $w=2.15e-07 $l=1.44375e-07 $layer=LI1_cond $X=14.025 $Y=0.402
+ $X2=14.11 $Y2=0.51
r105 26 28 10.1844 $w=2.13e-07 $l=1.9e-07 $layer=LI1_cond $X=14.025 $Y=0.402
+ $X2=13.835 $Y2=0.402
r106 24 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.75 $Y=1.435
+ $X2=13.75 $Y2=1.35
r107 24 38 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=13.75 $Y=1.435
+ $X2=13.75 $Y2=2.115
r108 20 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.665 $Y=1.35
+ $X2=13.75 $Y2=1.35
r109 20 35 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=13.665 $Y=1.35
+ $X2=13.185 $Y2=1.35
r110 18 41 46.5982 $w=3.31e-07 $l=3.2e-07 $layer=POLY_cond $X=12.78 $Y=1.335
+ $X2=12.46 $Y2=1.335
r111 17 34 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=12.78 $Y=1.205
+ $X2=13.015 $Y2=1.205
r112 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.78
+ $Y=1.205 $X2=12.78 $Y2=1.205
r113 11 41 21.295 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=12.46 $Y=1.04
+ $X2=12.46 $Y2=1.335
r114 11 13 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=12.46 $Y=1.04
+ $X2=12.46 $Y2=0.445
r115 7 41 23.2991 $w=3.31e-07 $l=3.66367e-07 $layer=POLY_cond $X=12.3 $Y=1.63
+ $X2=12.46 $Y2=1.335
r116 7 9 239.758 $w=2.5e-07 $l=9.65e-07 $layer=POLY_cond $X=12.3 $Y=1.63
+ $X2=12.3 $Y2=2.595
r117 2 37 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=13.52
+ $Y=2.095 $X2=13.66 $Y2=2.28
r118 1 28 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=13.695
+ $Y=0.235 $X2=13.835 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_2092_47# 1 2 7 9 12 14 15 16 18 19 21
+ 23 25 29 31 35 37 40 41 46 50 53
c156 46 0 1.68946e-19 $X=11.675 $Y=0.47
c157 40 0 1.03775e-19 $X=12.37 $Y=1.685
c158 15 0 2.03987e-19 $X=14.05 $Y=1.02
r159 57 61 39.8953 $w=2.96e-07 $l=2.45e-07 $layer=POLY_cond $X=13.68 $Y=0.93
+ $X2=13.925 $Y2=0.93
r160 57 59 9.77027 $w=2.96e-07 $l=6e-08 $layer=POLY_cond $X=13.68 $Y=0.93
+ $X2=13.62 $Y2=0.93
r161 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.68
+ $Y=0.93 $X2=13.68 $Y2=0.93
r162 53 56 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=13.68 $Y=0.775
+ $X2=13.68 $Y2=0.93
r163 50 52 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=12.37 $Y=0.59
+ $X2=12.37 $Y2=0.775
r164 46 48 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=11.675 $Y=0.47
+ $X2=11.675 $Y2=0.59
r165 42 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.455 $Y=0.775
+ $X2=12.37 $Y2=0.775
r166 41 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.515 $Y=0.775
+ $X2=13.68 $Y2=0.775
r167 41 42 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=13.515 $Y=0.775
+ $X2=12.455 $Y2=0.775
r168 39 52 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=12.37 $Y=0.86
+ $X2=12.37 $Y2=0.775
r169 39 40 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=12.37 $Y=0.86
+ $X2=12.37 $Y2=1.685
r170 38 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.84 $Y=0.59
+ $X2=11.675 $Y2=0.59
r171 37 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.285 $Y=0.59
+ $X2=12.37 $Y2=0.59
r172 37 38 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=12.285 $Y=0.59
+ $X2=11.84 $Y2=0.59
r173 36 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.63 $Y=1.77
+ $X2=11.465 $Y2=1.77
r174 35 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.285 $Y=1.77
+ $X2=12.37 $Y2=1.685
r175 35 36 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=12.285 $Y=1.77
+ $X2=11.63 $Y2=1.77
r176 31 33 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=11.465 $Y=2.2
+ $X2=11.465 $Y2=2.9
r177 29 44 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.465 $Y=1.855
+ $X2=11.465 $Y2=1.77
r178 29 31 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=11.465 $Y=1.855
+ $X2=11.465 $Y2=2.2
r179 23 28 1.49928 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.035 $Y=0.945
+ $X2=15.035 $Y2=1.02
r180 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=15.035 $Y=0.945
+ $X2=15.035 $Y2=0.66
r181 19 28 6.78873 $w=1.42e-07 $l=2e-08 $layer=POLY_cond $X=15.015 $Y=1.02
+ $X2=15.035 $Y2=1.02
r182 19 26 115.408 $w=1.42e-07 $l=3.4e-07 $layer=POLY_cond $X=15.015 $Y=1.02
+ $X2=14.675 $Y2=1.02
r183 19 21 334.17 $w=2.5e-07 $l=1.345e-06 $layer=POLY_cond $X=15.015 $Y=1.095
+ $X2=15.015 $Y2=2.44
r184 16 26 1.49928 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.675 $Y=0.945
+ $X2=14.675 $Y2=1.02
r185 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=14.675 $Y=0.945
+ $X2=14.675 $Y2=0.66
r186 15 61 32.0583 $w=2.96e-07 $l=1.63936e-07 $layer=POLY_cond $X=14.05 $Y=1.02
+ $X2=13.925 $Y2=0.93
r187 14 26 24.2889 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.6 $Y=1.02
+ $X2=14.675 $Y2=1.02
r188 14 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=14.6 $Y=1.02
+ $X2=14.05 $Y2=1.02
r189 10 61 6.82538 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.925 $Y=1.095
+ $X2=13.925 $Y2=0.93
r190 10 12 372.68 $w=2.5e-07 $l=1.5e-06 $layer=POLY_cond $X=13.925 $Y=1.095
+ $X2=13.925 $Y2=2.595
r191 7 59 18.6531 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.62 $Y=0.765
+ $X2=13.62 $Y2=0.93
r192 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.62 $Y=0.765
+ $X2=13.62 $Y2=0.445
r193 2 44 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=11.245
+ $Y=1.705 $X2=11.465 $Y2=1.85
r194 2 33 600 $w=1.7e-07 $l=1.30036e-06 $layer=licon1_PDIFF $count=1 $X=11.245
+ $Y=1.705 $X2=11.465 $Y2=2.9
r195 2 31 300 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_PDIFF $count=2 $X=11.245
+ $Y=1.705 $X2=11.465 $Y2=2.2
r196 1 46 182 $w=1.7e-07 $l=1.32731e-06 $layer=licon1_NDIFF $count=1 $X=10.46
+ $Y=0.235 $X2=11.675 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_2863_90# 1 2 9 13 17 23 26 28 31 35 39
+ 40 45 47
c70 26 0 7.76453e-20 $X=15.515 $Y=1.74
r71 43 45 4.16027 $w=4.58e-07 $l=1.6e-07 $layer=LI1_cond $X=14.46 $Y=0.66
+ $X2=14.62 $Y2=0.66
r72 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=15.515
+ $Y=1.235 $X2=15.515 $Y2=1.235
r73 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=15.515 $Y=1.57
+ $X2=15.515 $Y2=1.235
r74 36 47 3.11956 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=14.915 $Y=1.655
+ $X2=14.725 $Y2=1.655
r75 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=15.35 $Y=1.655
+ $X2=15.515 $Y2=1.57
r76 35 36 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=15.35 $Y=1.655
+ $X2=14.915 $Y2=1.655
r77 31 33 21.5325 $w=3.78e-07 $l=7.1e-07 $layer=LI1_cond $X=14.725 $Y=2.085
+ $X2=14.725 $Y2=2.795
r78 29 47 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=14.725 $Y=1.74
+ $X2=14.725 $Y2=1.655
r79 29 31 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=14.725 $Y=1.74
+ $X2=14.725 $Y2=2.085
r80 28 47 3.40559 $w=2.75e-07 $l=1.41244e-07 $layer=LI1_cond $X=14.62 $Y=1.57
+ $X2=14.725 $Y2=1.655
r81 27 45 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=14.62 $Y=0.89
+ $X2=14.62 $Y2=0.66
r82 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=14.62 $Y=0.89
+ $X2=14.62 $Y2=1.57
r83 25 40 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=15.515 $Y=1.575
+ $X2=15.515 $Y2=1.235
r84 25 26 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.515 $Y=1.575
+ $X2=15.515 $Y2=1.74
r85 22 40 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=15.515 $Y=1.22
+ $X2=15.515 $Y2=1.235
r86 22 23 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=15.515 $Y=1.145
+ $X2=15.825 $Y2=1.145
r87 19 22 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=15.465 $Y=1.145
+ $X2=15.515 $Y2=1.145
r88 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.825 $Y=1.07
+ $X2=15.825 $Y2=1.145
r89 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=15.825 $Y=1.07
+ $X2=15.825 $Y2=0.66
r90 13 26 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=15.545 $Y=2.44
+ $X2=15.545 $Y2=1.74
r91 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.465 $Y=1.07
+ $X2=15.465 $Y2=1.145
r92 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=15.465 $Y=1.07
+ $X2=15.465 $Y2=0.66
r93 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=14.605
+ $Y=1.94 $X2=14.75 $Y2=2.795
r94 2 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=14.605
+ $Y=1.94 $X2=14.75 $Y2=2.085
r95 1 43 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=14.315
+ $Y=0.45 $X2=14.46 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%A_116_419# 1 2 3 4 5 19 20 24 27 28 29 31
+ 32 33 36 39 41 43 44 48 49 51 55 56
c137 56 0 8.95267e-20 $X=6.87 $Y=1.145
c138 36 0 1.31384e-19 $X=6.87 $Y=0.79
c139 28 0 5.74786e-20 $X=4.84 $Y=2.98
c140 24 0 1.37977e-19 $X=3.73 $Y=2.59
r141 54 55 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.855 $Y=2.475
+ $X2=2.855 $Y2=2.59
r142 51 54 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.855 $Y=2.395
+ $X2=2.855 $Y2=2.475
r143 48 49 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=0.74
+ $X2=1.15 $Y2=0.74
r144 43 45 2.3174 $w=7.98e-07 $l=1.55e-07 $layer=LI1_cond $X=0.49 $Y=2.24
+ $X2=0.49 $Y2=2.395
r145 43 44 11.434 $w=7.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.49 $Y=2.24
+ $X2=0.49 $Y2=2.075
r146 41 56 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=6.95 $Y=2.085
+ $X2=6.95 $Y2=1.145
r147 39 58 3.40825 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=6.95 $Y=2.46
+ $X2=6.95 $Y2=2.607
r148 39 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.95 $Y=2.46
+ $X2=6.95 $Y2=2.085
r149 34 56 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=0.98
+ $X2=6.87 $Y2=1.145
r150 34 36 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.87 $Y=0.98
+ $X2=6.87 $Y2=0.79
r151 32 58 3.40825 $w=1.7e-07 $l=1.11781e-07 $layer=LI1_cond $X=6.865 $Y=2.545
+ $X2=6.95 $Y2=2.607
r152 32 33 121.021 $w=1.68e-07 $l=1.855e-06 $layer=LI1_cond $X=6.865 $Y=2.545
+ $X2=5.01 $Y2=2.545
r153 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.925 $Y=2.63
+ $X2=5.01 $Y2=2.545
r154 30 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.925 $Y=2.63
+ $X2=4.925 $Y2=2.895
r155 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.84 $Y=2.98
+ $X2=4.925 $Y2=2.895
r156 28 29 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.84 $Y=2.98
+ $X2=3.9 $Y2=2.98
r157 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.815 $Y=2.895
+ $X2=3.9 $Y2=2.98
r158 26 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.815 $Y=2.675
+ $X2=3.815 $Y2=2.895
r159 25 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=2.59
+ $X2=2.855 $Y2=2.59
r160 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.73 $Y=2.59
+ $X2=3.815 $Y2=2.675
r161 24 25 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.73 $Y=2.59
+ $X2=3.02 $Y2=2.59
r162 21 45 10.2089 $w=1.7e-07 $l=4e-07 $layer=LI1_cond $X=0.89 $Y=2.395 $X2=0.49
+ $Y2=2.395
r163 20 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=2.395
+ $X2=2.855 $Y2=2.395
r164 20 21 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=2.69 $Y=2.395
+ $X2=0.89 $Y2=2.395
r165 19 49 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=0.26 $Y=0.705
+ $X2=1.15 $Y2=0.705
r166 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.175 $Y=0.79
+ $X2=0.26 $Y2=0.705
r167 16 44 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=0.175 $Y=0.79
+ $X2=0.175 $Y2=2.075
r168 5 58 600 $w=1.7e-07 $l=7.09753e-07 $layer=licon1_PDIFF $count=1 $X=6.825
+ $Y=1.94 $X2=6.95 $Y2=2.59
r169 5 41 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.825
+ $Y=1.94 $X2=6.95 $Y2=2.085
r170 4 54 300 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.715
+ $Y=2.095 $X2=2.855 $Y2=2.475
r171 3 43 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.095 $X2=0.725 $Y2=2.24
r172 2 36 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=6.725
+ $Y=0.595 $X2=6.87 $Y2=0.79
r173 1 48 182 $w=1.7e-07 $l=4.36348e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.44 $X2=1.315 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 49 55
+ 59 63 68 69 71 72 74 75 76 78 99 106 118 127 128 131 134 137 140 143
r173 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r174 141 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=15.12 $Y2=3.33
r175 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r176 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r177 134 135 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r178 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r179 128 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=15.12 $Y2=3.33
r180 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r181 125 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.445 $Y=3.33
+ $X2=15.28 $Y2=3.33
r182 125 127 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=15.445 $Y=3.33
+ $X2=16.08 $Y2=3.33
r183 124 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r184 123 124 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r185 121 124 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r186 120 123 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r187 120 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r188 118 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.025 $Y=3.33
+ $X2=14.19 $Y2=3.33
r189 118 123 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=14.025 $Y=3.33
+ $X2=13.68 $Y2=3.33
r190 117 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r191 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r192 114 117 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=12.24 $Y2=3.33
r193 114 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r194 113 116 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=10.8 $Y=3.33
+ $X2=12.24 $Y2=3.33
r195 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r196 111 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.41 $Y=3.33
+ $X2=10.245 $Y2=3.33
r197 111 113 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.41 $Y=3.33
+ $X2=10.8 $Y2=3.33
r198 110 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r199 110 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r200 109 110 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r201 107 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.915 $Y=3.33
+ $X2=8.75 $Y2=3.33
r202 107 109 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=8.915 $Y=3.33
+ $X2=9.84 $Y2=3.33
r203 106 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.08 $Y=3.33
+ $X2=10.245 $Y2=3.33
r204 106 109 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.08 $Y=3.33
+ $X2=9.84 $Y2=3.33
r205 105 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r206 104 105 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r207 101 104 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r208 101 102 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r209 99 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.585 $Y=3.33
+ $X2=8.75 $Y2=3.33
r210 99 104 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.585 $Y=3.33
+ $X2=8.4 $Y2=3.33
r211 98 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r212 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r213 95 98 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r214 94 97 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r215 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r216 92 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r217 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r218 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r219 89 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r220 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r221 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r222 86 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=3.33
+ $X2=1.745 $Y2=3.33
r223 86 88 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.91 $Y=3.33
+ $X2=2.16 $Y2=3.33
r224 85 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r226 81 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r227 80 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r228 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r229 78 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=3.33
+ $X2=1.745 $Y2=3.33
r230 78 84 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.58 $Y=3.33
+ $X2=1.2 $Y2=3.33
r231 76 105 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=8.4 $Y2=3.33
r232 76 102 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=5.52 $Y2=3.33
r233 74 116 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=12.4 $Y=3.33
+ $X2=12.24 $Y2=3.33
r234 74 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.4 $Y=3.33
+ $X2=12.525 $Y2=3.33
r235 73 120 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=12.65 $Y=3.33
+ $X2=12.72 $Y2=3.33
r236 73 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.65 $Y=3.33
+ $X2=12.525 $Y2=3.33
r237 71 97 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.04 $Y2=3.33
r238 71 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.345 $Y2=3.33
r239 70 101 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.51 $Y=3.33
+ $X2=5.52 $Y2=3.33
r240 70 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=3.33
+ $X2=5.345 $Y2=3.33
r241 68 91 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.22 $Y=3.33 $X2=3.12
+ $Y2=3.33
r242 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=3.33
+ $X2=3.385 $Y2=3.33
r243 67 94 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.55 $Y=3.33 $X2=3.6
+ $Y2=3.33
r244 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=3.33
+ $X2=3.385 $Y2=3.33
r245 63 66 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=15.28 $Y=2.085
+ $X2=15.28 $Y2=2.795
r246 61 143 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.28 $Y=3.245
+ $X2=15.28 $Y2=3.33
r247 61 66 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=15.28 $Y=3.245
+ $X2=15.28 $Y2=2.795
r248 60 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.355 $Y=3.33
+ $X2=14.19 $Y2=3.33
r249 59 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.115 $Y=3.33
+ $X2=15.28 $Y2=3.33
r250 59 60 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=15.115 $Y=3.33
+ $X2=14.355 $Y2=3.33
r251 55 58 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=14.19 $Y=2.24
+ $X2=14.19 $Y2=2.95
r252 53 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.19 $Y=3.245
+ $X2=14.19 $Y2=3.33
r253 53 58 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=14.19 $Y=3.245
+ $X2=14.19 $Y2=2.95
r254 49 52 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=12.525 $Y=2.24
+ $X2=12.525 $Y2=2.95
r255 47 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.525 $Y=3.245
+ $X2=12.525 $Y2=3.33
r256 47 52 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=12.525 $Y=3.245
+ $X2=12.525 $Y2=2.95
r257 43 46 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=10.245 $Y=1.85
+ $X2=10.245 $Y2=2.56
r258 41 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.245 $Y=3.245
+ $X2=10.245 $Y2=3.33
r259 41 46 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=10.245 $Y=3.245
+ $X2=10.245 $Y2=2.56
r260 37 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.75 $Y=3.245
+ $X2=8.75 $Y2=3.33
r261 37 39 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=8.75 $Y=3.245
+ $X2=8.75 $Y2=2.53
r262 33 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=3.245
+ $X2=5.345 $Y2=3.33
r263 33 35 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=5.345 $Y=3.245
+ $X2=5.345 $Y2=2.895
r264 29 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=3.245
+ $X2=3.385 $Y2=3.33
r265 29 31 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.385 $Y=3.245
+ $X2=3.385 $Y2=2.945
r266 25 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=3.245
+ $X2=1.745 $Y2=3.33
r267 25 27 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.745 $Y=3.245
+ $X2=1.745 $Y2=2.885
r268 8 66 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=15.14
+ $Y=1.94 $X2=15.28 $Y2=2.795
r269 8 63 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.14
+ $Y=1.94 $X2=15.28 $Y2=2.085
r270 7 58 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=14.05
+ $Y=2.095 $X2=14.19 $Y2=2.95
r271 7 55 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.05
+ $Y=2.095 $X2=14.19 $Y2=2.24
r272 6 52 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=12.425
+ $Y=2.095 $X2=12.565 $Y2=2.95
r273 6 49 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.425
+ $Y=2.095 $X2=12.565 $Y2=2.24
r274 5 46 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=1.705 $X2=10.245 $Y2=2.56
r275 5 43 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=1.705 $X2=10.245 $Y2=1.85
r276 4 39 600 $w=1.7e-07 $l=8.62163e-07 $layer=licon1_PDIFF $count=1 $X=8.625
+ $Y=1.735 $X2=8.765 $Y2=2.53
r277 3 35 600 $w=1.7e-07 $l=1.02341e-06 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=2.04 $X2=5.345 $Y2=2.895
r278 2 31 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=2.095 $X2=3.385 $Y2=2.945
r279 1 27 600 $w=1.7e-07 $l=8.57146e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=2.095 $X2=1.745 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%Q 1 2 7 8 9 10 11 12 13
c22 11 0 7.76453e-20 $X=16.08 $Y=2.035
r23 33 45 2.45623 $w=5.58e-07 $l=1.15e-07 $layer=LI1_cond $X=15.925 $Y=2.2
+ $X2=15.925 $Y2=2.085
r24 13 39 0.427171 $w=5.58e-07 $l=2e-08 $layer=LI1_cond $X=15.925 $Y=2.775
+ $X2=15.925 $Y2=2.795
r25 12 13 7.90266 $w=5.58e-07 $l=3.7e-07 $layer=LI1_cond $X=15.925 $Y=2.405
+ $X2=15.925 $Y2=2.775
r26 12 33 4.3785 $w=5.58e-07 $l=2.05e-07 $layer=LI1_cond $X=15.925 $Y=2.405
+ $X2=15.925 $Y2=2.2
r27 11 45 1.06793 $w=5.58e-07 $l=5e-08 $layer=LI1_cond $X=15.925 $Y=2.035
+ $X2=15.925 $Y2=2.085
r28 11 42 4.45725 $w=5.58e-07 $l=1.15e-07 $layer=LI1_cond $X=15.925 $Y=2.035
+ $X2=15.925 $Y2=1.92
r29 10 42 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=16.04 $Y=1.665
+ $X2=16.04 $Y2=1.92
r30 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=16.04 $Y=1.295
+ $X2=16.04 $Y2=1.665
r31 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=16.04 $Y=0.925
+ $X2=16.04 $Y2=1.295
r32 8 26 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=16.04 $Y=0.925
+ $X2=16.04 $Y2=0.66
r33 7 26 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=16.04 $Y=0.555
+ $X2=16.04 $Y2=0.66
r34 2 45 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.67
+ $Y=1.94 $X2=15.81 $Y2=2.085
r35 2 39 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=15.67
+ $Y=1.94 $X2=15.81 $Y2=2.795
r36 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=15.9
+ $Y=0.45 $X2=16.04 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%noxref_23 1 2 7 11 16
r28 14 16 10.4571 $w=1.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.335 $Y=0.352
+ $X2=0.5 $Y2=0.352
r29 9 11 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.215 $Y=0.435
+ $X2=2.215 $Y2=0.65
r30 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.05 $Y=0.35
+ $X2=2.215 $Y2=0.435
r31 7 16 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=2.05 $Y=0.35 $X2=0.5
+ $Y2=0.35
r32 2 11 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.44 $X2=2.215 $Y2=0.65
r33 1 14 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.205 $X2=0.335 $Y2=0.35
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_LP2%VGND 1 2 3 4 5 18 22 24 28 32 36 38 40 45
+ 53 61 68 69 72 75 78 81 84
c134 69 0 2.36927e-20 $X=16.08 $Y=0
c135 61 0 9.32417e-20 $X=15.085 $Y=0
c136 53 0 1.95202e-19 $X=12.635 $Y=0
c137 18 0 1.2046e-19 $X=2.725 $Y=0.65
r138 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r139 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r140 78 79 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r141 75 76 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r142 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r143 69 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=15.12 $Y2=0
r144 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r145 66 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.415 $Y=0
+ $X2=15.25 $Y2=0
r146 66 68 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=15.415 $Y=0
+ $X2=16.08 $Y2=0
r147 65 85 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=15.12 $Y2=0
r148 65 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r149 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r150 62 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.965 $Y=0
+ $X2=12.8 $Y2=0
r151 62 64 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=12.965 $Y=0
+ $X2=13.2 $Y2=0
r152 61 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.085 $Y=0
+ $X2=15.25 $Y2=0
r153 61 64 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=15.085 $Y=0
+ $X2=13.2 $Y2=0
r154 60 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r155 59 60 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r156 57 60 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=12.24 $Y2=0
r157 57 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r158 56 59 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=12.24 $Y2=0
r159 56 57 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r160 54 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.18 $Y=0 $X2=9.015
+ $Y2=0
r161 54 56 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=9.18 $Y=0 $X2=9.36
+ $Y2=0
r162 53 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.635 $Y=0
+ $X2=12.8 $Y2=0
r163 53 59 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.635 $Y=0
+ $X2=12.24 $Y2=0
r164 52 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r165 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r166 49 52 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=5.04 $Y2=0
r167 49 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r168 48 51 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r169 48 49 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r170 46 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.725
+ $Y2=0
r171 46 48 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.12
+ $Y2=0
r172 45 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.375
+ $Y2=0
r173 45 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.04
+ $Y2=0
r174 43 73 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r175 42 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r176 40 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=0 $X2=2.725
+ $Y2=0
r177 40 42 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=2.56 $Y=0 $X2=0.24
+ $Y2=0
r178 38 79 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=8.16 $Y=0 $X2=8.88
+ $Y2=0
r179 38 76 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=8.16 $Y=0 $X2=5.52
+ $Y2=0
r180 34 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.25 $Y=0.085
+ $X2=15.25 $Y2=0
r181 34 36 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=15.25 $Y=0.085
+ $X2=15.25 $Y2=0.66
r182 30 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.8 $Y=0.085
+ $X2=12.8 $Y2=0
r183 30 32 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=12.8 $Y=0.085
+ $X2=12.8 $Y2=0.4
r184 26 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.015 $Y=0.085
+ $X2=9.015 $Y2=0
r185 26 28 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=9.015 $Y=0.085
+ $X2=9.015 $Y2=0.28
r186 25 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=0 $X2=5.375
+ $Y2=0
r187 24 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.85 $Y=0 $X2=9.015
+ $Y2=0
r188 24 25 215.947 $w=1.68e-07 $l=3.31e-06 $layer=LI1_cond $X=8.85 $Y=0 $X2=5.54
+ $Y2=0
r189 20 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=0.085
+ $X2=5.375 $Y2=0
r190 20 22 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=5.375 $Y=0.085
+ $X2=5.375 $Y2=0.62
r191 16 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0
r192 16 18 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0.65
r193 5 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=15.11
+ $Y=0.45 $X2=15.25 $Y2=0.66
r194 4 32 182 $w=1.7e-07 $l=3.37565e-07 $layer=licon1_NDIFF $count=1 $X=12.535
+ $Y=0.235 $X2=12.8 $Y2=0.4
r195 3 28 182 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_NDIFF $count=1 $X=8.795
+ $Y=0.33 $X2=9.015 $Y2=0.28
r196 2 22 182 $w=1.7e-07 $l=2.32164e-07 $layer=licon1_NDIFF $count=1 $X=5.155
+ $Y=0.595 $X2=5.375 $Y2=0.62
r197 1 18 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=2.505
+ $Y=0.44 $X2=2.725 $Y2=0.65
.ends

