* NGSPICE file created from sky130_fd_sc_lp__or2_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or2_1 A B VGND VNB VPB VPWR X
M1000 X a_76_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=4.263e+11p ps=4.02e+06u
M1001 a_76_367# B VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1002 VGND A a_76_367# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_159_367# B a_76_367# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.113e+11p ps=1.37e+06u
M1004 X a_76_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=5.019e+11p ps=3.85e+06u
M1005 VPWR A a_159_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

