* File: sky130_fd_sc_lp__o32ai_2.spice
* Created: Fri Aug 28 11:18:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32ai_2.pex.spice"
.subckt sky130_fd_sc_lp__o32ai_2  VNB VPB B2 B1 A3 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1004 N_A_39_65#_M1004_d N_B2_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.9 A=0.126 P=1.98 MULT=1
MM1019 N_A_39_65#_M1019_d N_B2_M1019_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.4 A=0.126 P=1.98 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_A_39_65#_M1019_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1512 PD=1.2 PS=1.2 NRD=11.424 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75003.9 A=0.126 P=1.98 MULT=1
MM1012 N_Y_M1006_d N_B1_M1012_g N_A_39_65#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1512 PD=1.2 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75001.6
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1007 N_A_39_65#_M1012_s N_A3_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.3402 PD=1.2 PS=1.65 NRD=0 NRS=9.996 M=1 R=5.6 SA=75002.1
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1018 N_A_39_65#_M1018_d N_A3_M1018_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1218 AS=0.3402 PD=1.13 PS=1.65 NRD=0 NRS=0 M=1 R=5.6 SA=75003.1
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_39_65#_M1018_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1302 AS=0.1218 PD=1.15 PS=1.13 NRD=0 NRS=1.428 M=1 R=5.6 SA=75003.5
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1002_d N_A2_M1013_g N_A_39_65#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1302 AS=0.1176 PD=1.15 PS=1.12 NRD=4.284 NRS=0 M=1 R=5.6 SA=75004
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A1_M1001_g N_A_39_65#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.4
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1001_d N_A1_M1010_g N_A_39_65#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75004.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_39_367#_M1005_d N_B2_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1015 N_A_39_367#_M1015_d N_B2_M1015_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_A_39_367#_M1015_d N_B1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_A_39_367#_M1016_d N_B1_M1016_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1011 N_A_519_365#_M1011_d N_A3_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1017 N_A_519_365#_M1017_d N_A3_M1017_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 N_A_778_365#_M1003_d N_A2_M1003_g N_A_519_365#_M1017_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_A_778_365#_M1003_d N_A2_M1014_g N_A_519_365#_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_778_365#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g N_A_778_365#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3698 P=16.99
*
.include "sky130_fd_sc_lp__o32ai_2.pxi.spice"
*
.ends
*
*
