* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 VPWR a_221_70# a_372_397# VPB phighvt w=640000u l=150000u
+  ad=1.8268e+12p pd=1.445e+07u as=3.254e+11p ps=2.76e+06u
M1001 Q a_776_99# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=8.967e+11p ps=8.84e+06u
M1002 a_776_99# a_626_125# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1003 VGND D a_31_464# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1004 a_221_70# GATE_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 a_221_70# GATE_N VPWR VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1006 VGND a_776_99# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_582_473# a_31_464# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1008 Q a_776_99# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1009 a_626_125# a_372_397# a_582_473# VPB phighvt w=640000u l=150000u
+  ad=2.286e+11p pd=2.07e+06u as=0p ps=0u
M1010 VPWR RESET_B a_776_99# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND RESET_B a_996_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1012 a_763_473# a_221_70# a_626_125# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1013 VPWR D a_31_464# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1014 VPWR a_776_99# a_763_473# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_626_125# a_221_70# a_554_125# VNB nshort w=420000u l=150000u
+  ad=1.47e+11p pd=1.54e+06u as=8.82e+10p ps=1.26e+06u
M1016 a_726_125# a_372_397# a_626_125# VNB nshort w=420000u l=150000u
+  ad=1.05e+11p pd=1.34e+06u as=0p ps=0u
M1017 a_996_47# a_626_125# a_776_99# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1018 VGND a_221_70# a_372_397# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1019 a_554_125# a_31_464# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_776_99# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_776_99# a_726_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
