* File: sky130_fd_sc_lp__or2_lp.spice
* Created: Fri Aug 28 11:21:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2_lp.pex.spice"
.subckt sky130_fd_sc_lp__or2_lp  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 A_118_114# N_A_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_196_114#_M1001_d N_A_M1001_g A_118_114# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1002 A_282_114# N_B_M1002_g N_A_196_114#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_B_M1008_g A_282_114# VNB NSHORT L=0.15 W=0.42 AD=0.105
+ AS=0.0441 PD=0.92 PS=0.63 NRD=62.856 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1005 A_484_114# N_A_196_114#_M1005_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.105 PD=0.66 PS=0.92 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_196_114#_M1003_g A_484_114# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_154_468# N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_196_114#_M1000_d N_B_M1000_g A_154_468# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_435_490# N_A_196_114#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_X_M1007_d N_A_196_114#_M1007_g A_435_490# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__or2_lp.pxi.spice"
*
.ends
*
*
