* NGSPICE file created from sky130_fd_sc_lp__nand4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
M1000 a_324_45# a_217_69# a_842_67# VNB nshort w=840000u l=150000u
+  ad=1.6287e+12p pd=1.271e+07u as=9.408e+11p ps=8.96e+06u
M1001 a_842_67# C a_1251_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.1508e+12p ps=1.114e+07u
M1002 VPWR A_N a_44_69# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.6242e+12p pd=3.254e+07u as=3.339e+11p ps=3.05e+06u
M1003 Y D VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.8224e+12p pd=2.464e+07u as=0p ps=0u
M1004 a_217_69# B_N VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=7.056e+11p ps=6.72e+06u
M1005 Y a_217_69# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_44_69# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1251_47# D VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y C VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1251_47# D VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_217_69# B_N VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1012 a_842_67# a_217_69# a_324_45# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1251_47# C a_842_67# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_44_69# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y a_44_69# a_324_45# VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1016 a_324_45# a_44_69# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_842_67# C a_1251_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_217_69# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1251_47# C a_842_67# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y C VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR D Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_324_45# a_217_69# a_842_67# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_217_69# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND D a_1251_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y a_44_69# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR D Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y D VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y a_44_69# a_324_45# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_324_45# a_44_69# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_842_67# a_217_69# a_324_45# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 Y a_217_69# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND A_N a_44_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1033 VPWR C Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND D a_1251_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Y a_44_69# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

