* File: sky130_fd_sc_lp__o21ba_lp.pex.spice
* Created: Fri Aug 28 11:06:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BA_LP%A1 3 7 9 11 18
r28 18 21 65.0426 $w=5.55e-07 $l=5.05e-07 $layer=POLY_cond $X=0.497 $Y=1.28
+ $X2=0.497 $Y2=1.785
r29 18 20 48.1474 $w=5.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.497 $Y=1.28
+ $X2=0.497 $Y2=1.115
r30 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.28 $X2=0.385 $Y2=1.28
r31 11 19 5.98039 $w=6.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=1.45
+ $X2=0.385 $Y2=1.45
r32 9 19 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.45
+ $X2=0.385 $Y2=1.45
r33 7 21 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.65 $Y=2.445
+ $X2=0.65 $Y2=1.785
r34 3 20 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.53 $Y=0.485
+ $X2=0.53 $Y2=1.115
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_LP%A2 3 7 11 12 13 14 18
r40 13 14 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.18 $Y=1.28
+ $X2=1.18 $Y2=1.665
r41 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.18
+ $Y=1.28 $X2=1.18 $Y2=1.28
r42 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=1.28
r43 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.62
+ $X2=1.18 $Y2=1.785
r44 10 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.115
+ $X2=1.18 $Y2=1.28
r45 7 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.12 $Y=0.485
+ $X2=1.12 $Y2=1.115
r46 3 12 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.14 $Y=2.445
+ $X2=1.14 $Y2=1.785
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_LP%A_317_29# 1 2 9 13 15 16 17 18 23 26 28 29
+ 35
r68 32 35 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.54 $Y=2.09
+ $X2=2.665 $Y2=2.09
r69 28 31 16.9582 $w=5.93e-07 $l=5.05e-07 $layer=LI1_cond $X=2.327 $Y=1.07
+ $X2=2.327 $Y2=1.575
r70 28 30 5.67112 $w=5.93e-07 $l=1.65e-07 $layer=LI1_cond $X=2.327 $Y=1.07
+ $X2=2.327 $Y2=0.905
r71 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.195
+ $Y=1.07 $X2=2.195 $Y2=1.07
r72 26 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=1.925
+ $X2=2.54 $Y2=2.09
r73 26 31 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.54 $Y=1.925
+ $X2=2.54 $Y2=1.575
r74 23 30 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.46 $Y=0.585
+ $X2=2.46 $Y2=0.905
r75 20 29 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.195 $Y=1.425
+ $X2=2.195 $Y2=1.07
r76 19 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.195 $Y=1.055
+ $X2=2.195 $Y2=1.07
r77 17 20 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.03 $Y=1.5
+ $X2=2.195 $Y2=1.425
r78 17 18 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.03 $Y=1.5
+ $X2=1.835 $Y2=1.5
r79 15 19 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.03 $Y=0.98
+ $X2=2.195 $Y2=1.055
r80 15 16 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.03 $Y=0.98
+ $X2=1.735 $Y2=0.98
r81 11 18 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=1.71 $Y=1.575
+ $X2=1.835 $Y2=1.5
r82 11 13 216.155 $w=2.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.71 $Y=1.575
+ $X2=1.71 $Y2=2.445
r83 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.66 $Y=0.905
+ $X2=1.735 $Y2=0.98
r84 7 9 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.66 $Y=0.905 $X2=1.66
+ $Y2=0.485
r85 2 35 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.945 $X2=2.665 $Y2=2.09
r86 1 23 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.375 $X2=2.46 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_LP%B1_N 1 3 4 5 8 12 15 20 23 24 27
r61 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.985
+ $Y=1.24 $X2=2.985 $Y2=1.24
r62 24 28 2.41001 $w=6.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.12 $Y=1.41
+ $X2=2.985 $Y2=1.41
r63 22 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.985 $Y=1.58
+ $X2=2.985 $Y2=1.24
r64 22 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.985 $Y=1.58
+ $X2=2.985 $Y2=1.745
r65 19 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.985 $Y=1.225
+ $X2=2.985 $Y2=1.24
r66 19 20 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=2.985 $Y=1.15
+ $X2=3.035 $Y2=1.15
r67 16 19 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=2.675 $Y=1.15
+ $X2=2.985 $Y2=1.15
r68 15 23 653.777 $w=1.5e-07 $l=1.275e-06 $layer=POLY_cond $X=3.075 $Y=3.02
+ $X2=3.075 $Y2=1.745
r69 10 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.035 $Y=1.075
+ $X2=3.035 $Y2=1.15
r70 10 12 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.035 $Y=1.075
+ $X2=3.035 $Y2=0.585
r71 6 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.675 $Y=1.075
+ $X2=2.675 $Y2=1.15
r72 6 8 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.675 $Y=1.075
+ $X2=2.675 $Y2=0.585
r73 4 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3 $Y=3.095
+ $X2=3.075 $Y2=3.02
r74 4 5 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=3 $Y=3.095 $X2=2.525
+ $Y2=3.095
r75 1 5 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=2.4 $Y=3.02
+ $X2=2.525 $Y2=3.095
r76 1 3 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.4 $Y=3.02 $X2=2.4
+ $Y2=2.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_LP%A_253_389# 1 2 9 13 17 20 21 25 26 29 31 34
+ 37
r89 34 36 10.4318 $w=3.58e-07 $l=2.25e-07 $layer=LI1_cond $X=1.86 $Y=0.49
+ $X2=1.86 $Y2=0.715
r90 31 32 9.36614 $w=5.08e-07 $l=3.9e-07 $layer=LI1_cond $X=1.565 $Y=2.13
+ $X2=1.565 $Y2=2.52
r91 29 37 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.5 $Y=2.435 $X2=3.5
+ $Y2=1.665
r92 26 39 66.9034 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=3.645 $Y=1.16
+ $X2=3.645 $Y2=1.665
r93 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.58
+ $Y=1.16 $X2=3.58 $Y2=1.16
r94 23 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=1.5
+ $X2=3.58 $Y2=1.665
r95 23 25 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.58 $Y=1.5 $X2=3.58
+ $Y2=1.16
r96 22 32 7.25644 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=1.85 $Y=2.52
+ $X2=1.565 $Y2=2.52
r97 21 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.415 $Y=2.52
+ $X2=3.5 $Y2=2.435
r98 21 22 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=3.415 $Y=2.52
+ $X2=1.85 $Y2=2.52
r99 20 31 9.75777 $w=5.08e-07 $l=2.70185e-07 $layer=LI1_cond $X=1.765 $Y=1.965
+ $X2=1.565 $Y2=2.13
r100 20 36 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.765 $Y=1.965
+ $X2=1.765 $Y2=0.715
r101 15 26 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=3.825 $Y=0.995
+ $X2=3.645 $Y2=1.16
r102 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.825 $Y=0.995
+ $X2=3.825 $Y2=0.585
r103 13 39 231.062 $w=2.5e-07 $l=9.3e-07 $layer=POLY_cond $X=3.775 $Y=2.595
+ $X2=3.775 $Y2=1.665
r104 7 26 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=3.465 $Y=0.995
+ $X2=3.645 $Y2=1.16
r105 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.465 $Y=0.995
+ $X2=3.465 $Y2=0.585
r106 2 31 300 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_PDIFF $count=2 $X=1.265
+ $Y=1.945 $X2=1.445 $Y2=2.13
r107 1 34 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.735
+ $Y=0.275 $X2=1.875 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_LP%VPWR 1 2 3 10 12 16 20 23 24 25 27 40 41 47
r44 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r47 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 35 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=3.33
+ $X2=2.055 $Y2=3.33
r49 35 37 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.22 $Y=3.33 $X2=3.12
+ $Y2=3.33
r50 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 30 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r54 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 28 44 4.54404 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.275 $Y2=3.33
r56 28 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=2.055 $Y2=3.33
r58 27 33 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 25 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r60 25 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 25 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 23 37 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.51 $Y2=3.33
r64 22 40 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=3.51 $Y2=3.33
r66 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.51 $Y=3.245
+ $X2=3.51 $Y2=3.33
r67 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.51 $Y=3.245
+ $X2=3.51 $Y2=2.95
r68 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=3.33
r69 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=2.95
r70 10 44 3.22214 $w=3.3e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.385 $Y=3.245
+ $X2=0.275 $Y2=3.33
r71 10 12 38.9386 $w=3.28e-07 $l=1.115e-06 $layer=LI1_cond $X=0.385 $Y=3.245
+ $X2=0.385 $Y2=2.13
r72 3 20 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.365
+ $Y=2.095 $X2=3.51 $Y2=2.95
r73 2 16 600 $w=1.7e-07 $l=1.10956e-06 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=1.945 $X2=2.055 $Y2=2.95
r74 1 12 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.24
+ $Y=1.945 $X2=0.385 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_LP%X 1 2 9 12 13 14 15 16 30
r21 30 40 1.92074 $w=2.38e-07 $l=4e-08 $layer=LI1_cond $X=4.085 $Y=2.035
+ $X2=4.085 $Y2=2.075
r22 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.04 $Y=2.405
+ $X2=4.04 $Y2=2.775
r23 15 33 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.04 $Y=2.405
+ $X2=4.04 $Y2=2.24
r24 14 33 4.99392 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=4.04 $Y=2.097
+ $X2=4.04 $Y2=2.24
r25 14 40 1.64602 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=4.04 $Y=2.097
+ $X2=4.04 $Y2=2.075
r26 14 30 1.10442 $w=2.38e-07 $l=2.3e-08 $layer=LI1_cond $X=4.085 $Y=2.012
+ $X2=4.085 $Y2=2.035
r27 13 14 16.6624 $w=2.38e-07 $l=3.47e-07 $layer=LI1_cond $X=4.085 $Y=1.665
+ $X2=4.085 $Y2=2.012
r28 12 13 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.085 $Y=1.295
+ $X2=4.085 $Y2=1.665
r29 11 12 23.0489 $w=2.38e-07 $l=4.8e-07 $layer=LI1_cond $X=4.085 $Y=0.815
+ $X2=4.085 $Y2=1.295
r30 9 11 8.90991 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.04 $Y=0.585
+ $X2=4.04 $Y2=0.815
r31 2 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.9
+ $Y=2.095 $X2=4.04 $Y2=2.24
r32 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.375 $X2=4.04 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_LP%A_34_55# 1 2 9 11 12 15
r29 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.335 $Y=0.765
+ $X2=1.335 $Y2=0.49
r30 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=0.85
+ $X2=1.335 $Y2=0.765
r31 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.17 $Y=0.85 $X2=0.48
+ $Y2=0.85
r32 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.315 $Y=0.765
+ $X2=0.48 $Y2=0.85
r33 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.315 $Y=0.765
+ $X2=0.315 $Y2=0.49
r34 2 15 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.275 $X2=1.335 $Y2=0.49
r35 1 9 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.275 $X2=0.315 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_LP%VGND 1 2 11 15 17 19 26 27 30 33
r45 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 27 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r48 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r49 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.25
+ $Y2=0
r50 24 26 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=4.08
+ $Y2=0
r51 23 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 20 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.825
+ $Y2=0
r54 20 22 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r55 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.25
+ $Y2=0
r56 19 22 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=3.085 $Y=0 $X2=1.2
+ $Y2=0
r57 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r58 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r59 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0
r60 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=3.25 $Y=0.085 $X2=3.25
+ $Y2=0.585
r61 9 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r62 9 11 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.42
r63 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.11
+ $Y=0.375 $X2=3.25 $Y2=0.585
r64 1 11 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.275 $X2=0.825 $Y2=0.42
.ends

