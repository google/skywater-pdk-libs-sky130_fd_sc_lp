* NGSPICE file created from sky130_fd_sc_lp__sleep_pargate_plv_21.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sleep_pargate_plv_21 VIRTPWR VPWR SLEEP VPB
M1000 VIRTPWR SLEEP VPWR VPB phighvt w=7e+06u l=150000u
+  ad=3.815e+12p pd=2.909e+07u as=3.815e+12p ps=2.909e+07u
M1001 VIRTPWR SLEEP VPWR VPB phighvt w=7e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VPWR SLEEP VIRTPWR VPB phighvt w=7e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

