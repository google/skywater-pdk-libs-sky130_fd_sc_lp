* NGSPICE file created from sky130_fd_sc_lp__a31oi_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a31oi_0 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 Y A1 a_201_47# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=1.008e+11p ps=1.32e+06u
M1001 VPWR A2 a_110_473# VPB phighvt w=640000u l=150000u
+  ad=3.488e+11p pd=3.65e+06u as=3.584e+11p ps=3.68e+06u
M1002 a_123_47# A3 VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.226e+11p ps=2.74e+06u
M1003 VGND B1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B1 a_110_473# VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1005 a_110_473# A3 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_110_473# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_201_47# A2 a_123_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

