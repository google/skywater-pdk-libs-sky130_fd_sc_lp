* File: sky130_fd_sc_lp__o2111a_0.pex.spice
* Created: Fri Aug 28 10:59:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111A_0%A_80_21# 1 2 3 12 15 18 20 24 25 26 27 28
+ 29 32 36 38 42 44
c91 38 0 8.91973e-20 $X=2.51 $Y=2.125
c92 26 0 8.95018e-20 $X=1.12 $Y=0.825
r93 40 42 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.655 $Y=2.215
+ $X2=2.655 $Y2=2.55
r94 39 44 7.03415 $w=1.8e-07 $l=1.33e-07 $layer=LI1_cond $X=1.57 $Y=2.125
+ $X2=1.437 $Y2=2.125
r95 38 40 7.31368 $w=1.8e-07 $l=1.84594e-07 $layer=LI1_cond $X=2.51 $Y=2.125
+ $X2=2.655 $Y2=2.215
r96 38 39 57.9192 $w=1.78e-07 $l=9.4e-07 $layer=LI1_cond $X=2.51 $Y=2.125
+ $X2=1.57 $Y2=2.125
r97 34 44 0.00540396 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=1.437 $Y=2.215
+ $X2=1.437 $Y2=2.125
r98 34 36 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=1.437 $Y=2.215
+ $X2=1.437 $Y2=2.55
r99 30 32 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.247 $Y=0.74
+ $X2=1.247 $Y2=0.445
r100 28 44 7.03415 $w=1.8e-07 $l=1.32e-07 $layer=LI1_cond $X=1.305 $Y=2.125
+ $X2=1.437 $Y2=2.125
r101 28 29 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.305 $Y=2.125
+ $X2=0.795 $Y2=2.125
r102 26 30 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.12 $Y=0.825
+ $X2=1.247 $Y2=0.74
r103 26 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.12 $Y=0.825
+ $X2=0.795 $Y2=0.825
r104 25 46 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.71
+ $X2=0.597 $Y2=1.545
r105 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.71 $X2=0.63 $Y2=1.71
r106 22 29 7.17723 $w=1.8e-07 $l=1.74284e-07 $layer=LI1_cond $X=0.66 $Y=2.035
+ $X2=0.795 $Y2=2.125
r107 22 24 13.872 $w=2.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.66 $Y=2.035
+ $X2=0.66 $Y2=1.71
r108 21 27 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.66 $Y=0.91
+ $X2=0.795 $Y2=0.825
r109 21 24 34.1465 $w=2.68e-07 $l=8e-07 $layer=LI1_cond $X=0.66 $Y=0.91 $X2=0.66
+ $Y2=1.71
r110 18 20 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.72 $Y=2.725
+ $X2=0.72 $Y2=2.215
r111 15 20 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.597 $Y=2.018
+ $X2=0.597 $Y2=2.215
r112 14 25 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.597 $Y=1.742
+ $X2=0.597 $Y2=1.71
r113 14 15 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.597 $Y=1.742
+ $X2=0.597 $Y2=2.018
r114 12 46 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=1.545
r115 3 42 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=2.405 $X2=2.635 $Y2=2.55
r116 2 36 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.295
+ $Y=2.405 $X2=1.435 $Y2=2.55
r117 1 32 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.235 $X2=1.285 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_0%D1 3 7 9 11 12 13 16 18 19 23
c55 18 0 6.75915e-20 $X=1.2 $Y=1.295
r56 18 19 14.8931 $w=3.23e-07 $l=4.2e-07 $layer=LI1_cond $X=1.197 $Y=1.245
+ $X2=1.197 $Y2=1.665
r57 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2
+ $Y=1.245 $X2=1.2 $Y2=1.245
r58 14 16 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.29 $Y=0.84 $X2=1.5
+ $Y2=0.84
r59 12 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.2 $Y=1.585 $X2=1.2
+ $Y2=1.245
r60 12 13 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.585
+ $X2=1.2 $Y2=1.75
r61 11 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.08 $X2=1.2
+ $Y2=1.245
r62 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.5 $Y=0.765 $X2=1.5
+ $Y2=0.84
r63 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.5 $Y=0.765 $X2=1.5
+ $Y2=0.445
r64 5 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=0.915
+ $X2=1.29 $Y2=0.84
r65 5 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=0.915
+ $X2=1.29 $Y2=1.08
r66 3 13 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=1.22 $Y=2.725
+ $X2=1.22 $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_0%C1 2 5 9 11 12 13 14 15 21
c49 12 0 1.15369e-19 $X=1.68 $Y=0.555
c50 9 0 1.57093e-19 $X=1.86 $Y=0.445
c51 5 0 1.21157e-19 $X=1.65 $Y=2.725
r52 21 23 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.32
+ $X2=1.755 $Y2=1.155
r53 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.77
+ $Y=1.32 $X2=1.77 $Y2=1.32
r54 15 22 12.8256 $w=3.08e-07 $l=3.45e-07 $layer=LI1_cond $X=1.7 $Y=1.665
+ $X2=1.7 $Y2=1.32
r55 14 22 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=1.7 $Y=1.295 $X2=1.7
+ $Y2=1.32
r56 13 14 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.7 $Y=0.925 $X2=1.7
+ $Y2=1.295
r57 12 13 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.7 $Y=0.555 $X2=1.7
+ $Y2=0.925
r58 9 23 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.86 $Y=0.445
+ $X2=1.86 $Y2=1.155
r59 5 11 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.65 $Y=2.725 $X2=1.65
+ $Y2=1.825
r60 2 11 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.755 $Y=1.645
+ $X2=1.755 $Y2=1.825
r61 1 21 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.755 $Y=1.335
+ $X2=1.755 $Y2=1.32
r62 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.755 $Y=1.335
+ $X2=1.755 $Y2=1.645
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_0%B1 3 6 9 11 12 13 17
c41 12 0 1.21157e-19 $X=2.16 $Y=1.295
c42 11 0 1.15369e-19 $X=2.325 $Y=1.865
c43 3 0 5.11591e-20 $X=2.22 $Y=0.445
r44 17 19 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.36
+ $X2=2.325 $Y2=1.195
r45 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.34
+ $Y=1.36 $X2=2.34 $Y2=1.36
r46 13 18 7.52173 $w=4.83e-07 $l=3.05e-07 $layer=LI1_cond $X=2.267 $Y=1.665
+ $X2=2.267 $Y2=1.36
r47 12 18 1.60299 $w=4.83e-07 $l=6.5e-08 $layer=LI1_cond $X=2.267 $Y=1.295
+ $X2=2.267 $Y2=1.36
r48 9 11 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.42 $Y=2.725
+ $X2=2.42 $Y2=1.865
r49 6 11 47.2362 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=2.325 $Y=1.685
+ $X2=2.325 $Y2=1.865
r50 5 17 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=2.325 $Y=1.375
+ $X2=2.325 $Y2=1.36
r51 5 6 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=2.325 $Y=1.375
+ $X2=2.325 $Y2=1.685
r52 3 19 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.22 $Y=0.445
+ $X2=2.22 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_0%A2 1 3 8 12 15 16 17 18 19 23
c50 18 0 5.11591e-20 $X=3.12 $Y=1.295
c51 16 0 1.4009e-19 $X=2.88 $Y=1.66
c52 12 0 3.0424e-20 $X=2.79 $Y=0.84
r53 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.88
+ $Y=1.32 $X2=2.88 $Y2=1.32
r54 19 24 8.25294 $w=4.98e-07 $l=3.45e-07 $layer=LI1_cond $X=2.965 $Y=1.665
+ $X2=2.965 $Y2=1.32
r55 18 24 0.598039 $w=4.98e-07 $l=2.5e-08 $layer=LI1_cond $X=2.965 $Y=1.295
+ $X2=2.965 $Y2=1.32
r56 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.88 $Y=1.66
+ $X2=2.88 $Y2=1.32
r57 16 17 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.66
+ $X2=2.88 $Y2=1.825
r58 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.155
+ $X2=2.88 $Y2=1.32
r59 10 12 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.65 $Y=0.84
+ $X2=2.79 $Y2=0.84
r60 8 17 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.85 $Y=2.725 $X2=2.85
+ $Y2=1.825
r61 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.79 $Y=0.915
+ $X2=2.79 $Y2=0.84
r62 4 15 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.79 $Y=0.915
+ $X2=2.79 $Y2=1.155
r63 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.65 $Y=0.765
+ $X2=2.65 $Y2=0.84
r64 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.65 $Y=0.765 $X2=2.65
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_0%A1 1 3 6 8 9 11 14 16 17 18 19 26
c40 11 0 8.91973e-20 $X=3.39 $Y=2.065
c41 8 0 2.12886e-20 $X=3.515 $Y=1.155
r42 18 19 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=2.035
r43 17 18 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.295
+ $X2=3.57 $Y2=1.665
r44 17 26 5.45074 $w=3.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.57 $Y=1.295
+ $X2=3.57 $Y2=1.12
r45 12 14 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.21 $Y=2.14
+ $X2=3.39 $Y2=2.14
r46 11 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.39 $Y=2.065
+ $X2=3.39 $Y2=2.14
r47 11 16 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.39 $Y=2.065
+ $X2=3.39 $Y2=1.625
r48 9 16 50.5417 $w=4e-07 $l=2e-07 $layer=POLY_cond $X=3.515 $Y=1.425 $X2=3.515
+ $Y2=1.625
r49 8 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.55 $Y=1.12
+ $X2=3.55 $Y2=1.12
r50 8 9 37.5404 $w=4e-07 $l=2.7e-07 $layer=POLY_cond $X=3.515 $Y=1.155 $X2=3.515
+ $Y2=1.425
r51 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.21 $Y=2.215
+ $X2=3.21 $Y2=2.14
r52 4 6 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.21 $Y=2.215 $X2=3.21
+ $Y2=2.725
r53 1 8 78.1911 $w=2.25e-07 $l=4.52106e-07 $layer=POLY_cond $X=3.15 $Y=0.765
+ $X2=3.515 $Y2=0.96
r54 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.15 $Y=0.765 $X2=3.15
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_0%X 1 2 7 8 9 10 11 12 13 24 38
r17 38 39 3.90788 $w=5.83e-07 $l=2e-08 $layer=LI1_cond $X=0.377 $Y=2.405
+ $X2=0.377 $Y2=2.385
r18 13 42 4.6003 $w=5.83e-07 $l=2.25e-07 $layer=LI1_cond $X=0.377 $Y=2.775
+ $X2=0.377 $Y2=2.55
r19 12 42 2.31037 $w=5.83e-07 $l=1.13e-07 $layer=LI1_cond $X=0.377 $Y=2.437
+ $X2=0.377 $Y2=2.55
r20 12 38 0.654265 $w=5.83e-07 $l=3.2e-08 $layer=LI1_cond $X=0.377 $Y=2.437
+ $X2=0.377 $Y2=2.405
r21 12 39 1.40854 $w=2.68e-07 $l=3.3e-08 $layer=LI1_cond $X=0.22 $Y=2.352
+ $X2=0.22 $Y2=2.385
r22 11 12 13.5305 $w=2.68e-07 $l=3.17e-07 $layer=LI1_cond $X=0.22 $Y=2.035
+ $X2=0.22 $Y2=2.352
r23 10 11 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=2.035
r24 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.665
r25 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.925 $X2=0.22
+ $Y2=1.295
r26 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.555 $X2=0.22
+ $Y2=0.925
r27 7 24 4.69514 $w=2.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.22 $Y=0.555
+ $X2=0.22 $Y2=0.445
r28 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.38
+ $Y=2.405 $X2=0.505 $Y2=2.55
r29 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_0%VPWR 1 2 3 12 16 18 20 23 24 25 31 35 41 45
r44 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 36 41 12.559 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=2.34 $Y=3.33 $X2=2.04
+ $Y2=3.33
r50 36 38 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 35 44 4.50438 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=3.26 $Y=3.33 $X2=3.55
+ $Y2=3.33
r52 35 38 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.26 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 31 41 12.559 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=1.74 $Y=3.33 $X2=2.04
+ $Y2=3.33
r55 31 33 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.74 $Y=3.33 $X2=1.68
+ $Y2=3.33
r56 29 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 25 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 25 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 23 28 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.84 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 23 24 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.84 $Y=3.33
+ $X2=0.987 $Y2=3.33
r62 22 33 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 22 24 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=0.987 $Y2=3.33
r64 18 44 3.26179 $w=3.3e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.55 $Y2=3.33
r65 18 20 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.425 $Y=3.245
+ $X2=3.425 $Y2=2.55
r66 14 41 2.52064 $w=6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=3.245 $X2=2.04
+ $Y2=3.33
r67 14 16 13.8546 $w=5.98e-07 $l=6.95e-07 $layer=LI1_cond $X=2.04 $Y=3.245
+ $X2=2.04 $Y2=2.55
r68 10 24 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.987 $Y=3.245
+ $X2=0.987 $Y2=3.33
r69 10 12 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=0.987 $Y=3.245
+ $X2=0.987 $Y2=2.55
r70 3 20 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.285
+ $Y=2.405 $X2=3.425 $Y2=2.55
r71 2 16 150 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=4 $X=1.725
+ $Y=2.405 $X2=2.205 $Y2=2.55
r72 1 12 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.795
+ $Y=2.405 $X2=0.97 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_0%VGND 1 2 9 13 16 17 18 20 33 34 37
c54 34 0 2.12886e-20 $X=3.6 $Y=0
c55 16 0 3.0424e-20 $X=2.735 $Y=0
r56 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r58 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r59 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r60 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r61 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r62 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r63 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r64 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r65 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r66 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r67 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r68 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r69 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r70 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r71 16 30 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.64
+ $Y2=0
r72 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.9
+ $Y2=0
r73 15 33 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=3.6
+ $Y2=0
r74 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.065 $Y=0 $X2=2.9
+ $Y2=0
r75 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=0.085 $X2=2.9
+ $Y2=0
r76 11 13 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.9 $Y=0.085
+ $X2=2.9 $Y2=0.41
r77 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r78 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0.445
r79 2 13 182 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_NDIFF $count=1 $X=2.725
+ $Y=0.235 $X2=2.9 $Y2=0.41
r80 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_0%A_459_47# 1 2 9 11 12 15
r31 13 15 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=3.39 $Y=0.695
+ $X2=3.39 $Y2=0.445
r32 11 13 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.25 $Y=0.78
+ $X2=3.39 $Y2=0.695
r33 11 12 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.25 $Y=0.78
+ $X2=2.565 $Y2=0.78
r34 7 12 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=2.417 $Y=0.695
+ $X2=2.565 $Y2=0.78
r35 7 9 9.76647 $w=2.93e-07 $l=2.5e-07 $layer=LI1_cond $X=2.417 $Y=0.695
+ $X2=2.417 $Y2=0.445
r36 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.235 $X2=3.365 $Y2=0.445
r37 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.235 $X2=2.435 $Y2=0.445
.ends

