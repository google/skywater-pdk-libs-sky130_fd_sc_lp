* File: sky130_fd_sc_lp__nand2b_m.pxi.spice
* Created: Wed Sep  2 10:03:54 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2B_M%A_N N_A_N_M1004_g N_A_N_c_54_n N_A_N_M1005_g
+ N_A_N_c_55_n A_N A_N A_N A_N A_N N_A_N_c_57_n PM_SKY130_FD_SC_LP__NAND2B_M%A_N
x_PM_SKY130_FD_SC_LP__NAND2B_M%B N_B_M1003_g N_B_M1001_g N_B_c_92_n N_B_c_93_n
+ N_B_c_94_n B B N_B_c_96_n PM_SKY130_FD_SC_LP__NAND2B_M%B
x_PM_SKY130_FD_SC_LP__NAND2B_M%A_46_54# N_A_46_54#_M1004_s N_A_46_54#_M1005_s
+ N_A_46_54#_M1000_g N_A_46_54#_M1002_g N_A_46_54#_c_137_n N_A_46_54#_c_143_n
+ N_A_46_54#_c_144_n N_A_46_54#_c_138_n N_A_46_54#_c_139_n N_A_46_54#_c_140_n
+ N_A_46_54#_c_146_n N_A_46_54#_c_147_n N_A_46_54#_c_148_n N_A_46_54#_c_149_n
+ N_A_46_54#_c_170_n N_A_46_54#_c_150_n N_A_46_54#_c_151_n
+ PM_SKY130_FD_SC_LP__NAND2B_M%A_46_54#
x_PM_SKY130_FD_SC_LP__NAND2B_M%VPWR N_VPWR_M1005_d N_VPWR_M1000_d N_VPWR_c_206_n
+ N_VPWR_c_207_n N_VPWR_c_208_n N_VPWR_c_209_n N_VPWR_c_210_n N_VPWR_c_211_n
+ VPWR N_VPWR_c_212_n N_VPWR_c_205_n PM_SKY130_FD_SC_LP__NAND2B_M%VPWR
x_PM_SKY130_FD_SC_LP__NAND2B_M%Y N_Y_M1002_d N_Y_M1003_d N_Y_c_248_n N_Y_c_242_n
+ Y Y Y Y Y Y N_Y_c_241_n N_Y_c_245_n Y PM_SKY130_FD_SC_LP__NAND2B_M%Y
x_PM_SKY130_FD_SC_LP__NAND2B_M%VGND N_VGND_M1004_d N_VGND_c_277_n N_VGND_c_278_n
+ N_VGND_c_279_n VGND N_VGND_c_280_n N_VGND_c_281_n
+ PM_SKY130_FD_SC_LP__NAND2B_M%VGND
cc_1 VNB N_A_N_M1004_g 0.0349731f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.48
cc_2 VNB N_A_N_c_54_n 0.0236294f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.523
cc_3 VNB N_A_N_c_55_n 0.010935f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.71
cc_4 VNB A_N 0.00323738f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB N_A_N_c_57_n 0.0231163f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.205
cc_6 VNB N_B_M1003_g 0.0104329f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.48
cc_7 VNB N_B_c_92_n 0.0185864f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.87
cc_8 VNB N_B_c_93_n 0.0241346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B_c_94_n 0.0175794f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.71
cc_10 VNB B 0.0031332f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_11 VNB N_B_c_96_n 0.0177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_46_54#_c_137_n 0.041136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_46_54#_c_138_n 0.0196257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_46_54#_c_139_n 0.0114071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_46_54#_c_140_n 0.046005f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.205
cc_16 VNB N_VPWR_c_205_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.712 $Y2=1.295
cc_17 VNB Y 0.00205552f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_18 VNB Y 0.0512422f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_19 VNB N_Y_c_241_n 0.0111748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_277_n 0.00601167f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.523
cc_21 VNB N_VGND_c_278_n 0.030974f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.87
cc_22 VNB N_VGND_c_279_n 0.00401293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_280_n 0.0372199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_281_n 0.182433f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.205
cc_25 VPB N_A_N_M1005_g 0.0705234f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.87
cc_26 VPB N_A_N_c_55_n 0.0118182f $X=-0.19 $Y=1.655 $X2=0.682 $Y2=1.71
cc_27 VPB A_N 0.00479347f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_28 VPB N_B_M1003_g 0.0612492f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.48
cc_29 VPB N_A_46_54#_M1000_g 0.0291107f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.87
cc_30 VPB N_A_46_54#_c_137_n 0.00332352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_A_46_54#_c_143_n 0.0260429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_46_54#_c_144_n 0.0171098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_A_46_54#_c_140_n 0.0320291f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=1.205
cc_34 VPB N_A_46_54#_c_146_n 0.00957747f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_46_54#_c_147_n 0.00661101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A_46_54#_c_148_n 0.0178592f $X=-0.19 $Y=1.655 $X2=0.712 $Y2=1.205
cc_37 VPB N_A_46_54#_c_149_n 0.0107864f $X=-0.19 $Y=1.655 $X2=0.712 $Y2=1.295
cc_38 VPB N_A_46_54#_c_150_n 0.0227256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_46_54#_c_151_n 0.00828103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_206_n 0.00467824f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.87
cc_41 VPB N_VPWR_c_207_n 0.0133303f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_42 VPB N_VPWR_c_208_n 0.0293489f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_43 VPB N_VPWR_c_209_n 0.00401228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_210_n 0.0155832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_211_n 0.00521708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_212_n 0.0128905f $X=-0.19 $Y=1.655 $X2=0.712 $Y2=1.205
cc_47 VPB N_VPWR_c_205_n 0.0647161f $X=-0.19 $Y=1.655 $X2=0.712 $Y2=1.295
cc_48 VPB N_Y_c_242_n 0.00384295f $X=-0.19 $Y=1.655 $X2=0.682 $Y2=1.71
cc_49 VPB Y 0.0399758f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_50 VPB Y 0.0130766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_Y_c_245_n 0.0103428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 N_A_N_c_54_n N_B_M1003_g 0.0618167f $X=0.682 $Y=1.523 $X2=0 $Y2=0
cc_53 A_N N_B_M1003_g 0.00357886f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_54 N_A_N_M1004_g N_B_c_92_n 0.00679495f $X=0.57 $Y=0.48 $X2=0 $Y2=0
cc_55 A_N N_B_c_92_n 0.00377894f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_56 A_N N_B_c_93_n 0.00139163f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_57 N_A_N_c_57_n N_B_c_93_n 0.013438f $X=0.705 $Y=1.205 $X2=0 $Y2=0
cc_58 N_A_N_c_54_n N_B_c_94_n 0.013438f $X=0.682 $Y=1.523 $X2=0 $Y2=0
cc_59 N_A_N_M1004_g B 2.36585e-19 $X=0.57 $Y=0.48 $X2=0 $Y2=0
cc_60 A_N B 0.0296515f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_61 N_A_N_c_57_n B 0.00152034f $X=0.705 $Y=1.205 $X2=0 $Y2=0
cc_62 N_A_N_M1004_g N_B_c_96_n 0.00559302f $X=0.57 $Y=0.48 $X2=0 $Y2=0
cc_63 A_N N_B_c_96_n 0.00190905f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_64 N_A_N_M1004_g N_A_46_54#_c_140_n 0.025516f $X=0.57 $Y=0.48 $X2=0 $Y2=0
cc_65 N_A_N_M1005_g N_A_46_54#_c_140_n 0.00599763f $X=0.795 $Y=2.87 $X2=0 $Y2=0
cc_66 A_N N_A_46_54#_c_140_n 0.108114f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_67 N_A_N_M1005_g N_A_46_54#_c_146_n 0.00561436f $X=0.795 $Y=2.87 $X2=0 $Y2=0
cc_68 N_A_N_M1005_g N_A_46_54#_c_147_n 0.0149736f $X=0.795 $Y=2.87 $X2=0 $Y2=0
cc_69 N_A_N_c_55_n N_A_46_54#_c_148_n 0.00367615f $X=0.682 $Y=1.71 $X2=0 $Y2=0
cc_70 A_N N_A_46_54#_c_148_n 0.0141035f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_71 N_A_N_M1005_g N_A_46_54#_c_151_n 0.00201618f $X=0.795 $Y=2.87 $X2=0 $Y2=0
cc_72 N_A_N_M1005_g N_VPWR_c_206_n 0.00280554f $X=0.795 $Y=2.87 $X2=0 $Y2=0
cc_73 N_A_N_M1005_g N_VPWR_c_208_n 0.00570116f $X=0.795 $Y=2.87 $X2=0 $Y2=0
cc_74 N_A_N_M1005_g N_VPWR_c_205_n 0.00751744f $X=0.795 $Y=2.87 $X2=0 $Y2=0
cc_75 A_N N_VGND_M1004_d 0.00418334f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_76 N_A_N_M1004_g N_VGND_c_277_n 0.00530658f $X=0.57 $Y=0.48 $X2=0 $Y2=0
cc_77 A_N N_VGND_c_277_n 0.00782932f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_78 N_A_N_M1004_g N_VGND_c_278_n 0.00521889f $X=0.57 $Y=0.48 $X2=0 $Y2=0
cc_79 A_N N_VGND_c_278_n 0.00449085f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_80 N_A_N_M1004_g N_VGND_c_281_n 0.0110722f $X=0.57 $Y=0.48 $X2=0 $Y2=0
cc_81 A_N N_VGND_c_281_n 0.00613101f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_82 N_B_M1003_g N_A_46_54#_M1000_g 0.0215288f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_83 N_B_M1003_g N_A_46_54#_c_137_n 0.00992388f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_84 B N_A_46_54#_c_137_n 0.00283196f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_85 N_B_c_96_n N_A_46_54#_c_137_n 0.0279607f $X=1.245 $Y=0.965 $X2=0 $Y2=0
cc_86 N_B_c_92_n N_A_46_54#_c_138_n 0.0254113f $X=1.245 $Y=0.8 $X2=0 $Y2=0
cc_87 B N_A_46_54#_c_139_n 8.46157e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_88 N_B_c_96_n N_A_46_54#_c_139_n 0.0254113f $X=1.245 $Y=0.965 $X2=0 $Y2=0
cc_89 N_B_M1003_g N_A_46_54#_c_149_n 0.0150659f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_90 N_B_c_94_n N_A_46_54#_c_149_n 0.00216786f $X=1.245 $Y=1.47 $X2=0 $Y2=0
cc_91 B N_A_46_54#_c_149_n 0.00435963f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_92 N_B_M1003_g N_A_46_54#_c_170_n 0.00219519f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_93 N_B_M1003_g N_A_46_54#_c_150_n 0.0377617f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_94 N_B_M1003_g N_A_46_54#_c_151_n 0.00581625f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_95 N_B_c_94_n N_A_46_54#_c_151_n 0.00114197f $X=1.245 $Y=1.47 $X2=0 $Y2=0
cc_96 B N_A_46_54#_c_151_n 0.00111561f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_97 N_B_M1003_g N_VPWR_c_206_n 0.00145709f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_98 N_B_M1003_g N_VPWR_c_207_n 7.52553e-19 $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_99 N_B_M1003_g N_VPWR_c_210_n 0.00570116f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_100 N_B_M1003_g N_VPWR_c_205_n 0.0105051f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_101 N_B_M1003_g N_Y_c_242_n 0.00287294f $X=1.225 $Y=2.87 $X2=0 $Y2=0
cc_102 N_B_c_92_n Y 7.40936e-19 $X=1.245 $Y=0.8 $X2=0 $Y2=0
cc_103 N_B_c_92_n N_VGND_c_277_n 0.00776291f $X=1.245 $Y=0.8 $X2=0 $Y2=0
cc_104 B N_VGND_c_277_n 0.00527585f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_105 N_B_c_96_n N_VGND_c_277_n 0.00220941f $X=1.245 $Y=0.965 $X2=0 $Y2=0
cc_106 N_B_c_92_n N_VGND_c_280_n 0.00550375f $X=1.245 $Y=0.8 $X2=0 $Y2=0
cc_107 N_B_c_92_n N_VGND_c_281_n 0.00879549f $X=1.245 $Y=0.8 $X2=0 $Y2=0
cc_108 B N_VGND_c_281_n 0.0050172f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_109 N_A_46_54#_c_147_n N_VPWR_c_206_n 0.00336215f $X=0.985 $Y=2.385 $X2=0
+ $Y2=0
cc_110 N_A_46_54#_c_151_n N_VPWR_c_206_n 0.00614722f $X=1.07 $Y=2.215 $X2=0
+ $Y2=0
cc_111 N_A_46_54#_M1000_g N_VPWR_c_207_n 0.00870102f $X=1.655 $Y=2.87 $X2=0
+ $Y2=0
cc_112 N_A_46_54#_c_146_n N_VPWR_c_208_n 0.00810105f $X=0.58 $Y=2.805 $X2=0
+ $Y2=0
cc_113 N_A_46_54#_M1000_g N_VPWR_c_210_n 0.00348402f $X=1.655 $Y=2.87 $X2=0
+ $Y2=0
cc_114 N_A_46_54#_M1000_g N_VPWR_c_205_n 0.00423222f $X=1.655 $Y=2.87 $X2=0
+ $Y2=0
cc_115 N_A_46_54#_c_146_n N_VPWR_c_205_n 0.00755621f $X=0.58 $Y=2.805 $X2=0
+ $Y2=0
cc_116 N_A_46_54#_c_147_n N_VPWR_c_205_n 3.21265e-19 $X=0.985 $Y=2.385 $X2=0
+ $Y2=0
cc_117 N_A_46_54#_c_148_n N_VPWR_c_205_n 0.0141156f $X=0.685 $Y=2.385 $X2=0
+ $Y2=0
cc_118 N_A_46_54#_c_151_n N_VPWR_c_205_n 0.00198333f $X=1.07 $Y=2.215 $X2=0
+ $Y2=0
cc_119 N_A_46_54#_M1000_g N_Y_c_248_n 2.03427e-19 $X=1.655 $Y=2.87 $X2=0 $Y2=0
cc_120 N_A_46_54#_c_146_n N_Y_c_248_n 2.5226e-19 $X=0.58 $Y=2.805 $X2=0 $Y2=0
cc_121 N_A_46_54#_c_146_n N_Y_c_242_n 0.00558332f $X=0.58 $Y=2.805 $X2=0 $Y2=0
cc_122 N_A_46_54#_c_149_n N_Y_c_242_n 0.0150051f $X=1.54 $Y=2.215 $X2=0 $Y2=0
cc_123 N_A_46_54#_c_138_n Y 0.00514268f $X=1.71 $Y=0.8 $X2=0 $Y2=0
cc_124 N_A_46_54#_M1000_g Y 0.00281355f $X=1.655 $Y=2.87 $X2=0 $Y2=0
cc_125 N_A_46_54#_c_143_n Y 0.00114707f $X=1.705 $Y=2.215 $X2=0 $Y2=0
cc_126 N_A_46_54#_c_144_n Y 0.00289409f $X=1.705 $Y=2.38 $X2=0 $Y2=0
cc_127 N_A_46_54#_c_138_n Y 0.00383122f $X=1.71 $Y=0.8 $X2=0 $Y2=0
cc_128 N_A_46_54#_c_139_n Y 0.0279082f $X=1.71 $Y=0.95 $X2=0 $Y2=0
cc_129 N_A_46_54#_c_149_n Y 0.0117991f $X=1.54 $Y=2.215 $X2=0 $Y2=0
cc_130 N_A_46_54#_c_170_n Y 0.0221382f $X=1.705 $Y=1.875 $X2=0 $Y2=0
cc_131 N_A_46_54#_c_150_n Y 0.0103241f $X=1.705 $Y=1.875 $X2=0 $Y2=0
cc_132 N_A_46_54#_M1000_g Y 0.0132129f $X=1.655 $Y=2.87 $X2=0 $Y2=0
cc_133 N_A_46_54#_c_144_n Y 0.00512433f $X=1.705 $Y=2.38 $X2=0 $Y2=0
cc_134 N_A_46_54#_c_149_n Y 0.02513f $X=1.54 $Y=2.215 $X2=0 $Y2=0
cc_135 N_A_46_54#_c_140_n N_VGND_c_278_n 0.00725068f $X=0.355 $Y=0.545 $X2=0
+ $Y2=0
cc_136 N_A_46_54#_c_138_n N_VGND_c_280_n 0.0051993f $X=1.71 $Y=0.8 $X2=0 $Y2=0
cc_137 N_A_46_54#_c_138_n N_VGND_c_281_n 0.010453f $X=1.71 $Y=0.8 $X2=0 $Y2=0
cc_138 N_A_46_54#_c_140_n N_VGND_c_281_n 0.00680975f $X=0.355 $Y=0.545 $X2=0
+ $Y2=0
cc_139 N_VPWR_c_210_n N_Y_c_248_n 0.00725617f $X=1.705 $Y=3.33 $X2=0 $Y2=0
cc_140 N_VPWR_c_205_n N_Y_c_248_n 0.0068189f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_141 N_VPWR_c_207_n Y 0.0219898f $X=1.87 $Y=2.935 $X2=0 $Y2=0
cc_142 N_VPWR_c_210_n Y 0.00273981f $X=1.705 $Y=3.33 $X2=0 $Y2=0
cc_143 N_VPWR_c_212_n Y 6.4789e-19 $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_144 N_VPWR_c_205_n Y 0.00688563f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_145 N_VPWR_c_212_n N_Y_c_245_n 0.00312529f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_146 N_VPWR_c_205_n N_Y_c_245_n 0.00497556f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_147 Y N_VGND_c_277_n 0.00428711f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_148 Y N_VGND_c_280_n 0.00890169f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_149 N_Y_c_241_n N_VGND_c_280_n 0.00555891f $X=2.16 $Y=0.65 $X2=0 $Y2=0
cc_150 Y N_VGND_c_281_n 0.0108779f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_151 N_Y_c_241_n N_VGND_c_281_n 0.00592732f $X=2.16 $Y=0.65 $X2=0 $Y2=0
