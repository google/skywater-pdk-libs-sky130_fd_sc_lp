* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fa_m A B CIN VGND VNB VPB VPWR COUT SUM
X0 VGND A a_843_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_385_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_1101_119# SUM VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 COUT a_80_241# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1101_119# CIN a_1195_391# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1195_391# B a_1267_391# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_1267_391# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_227_125# B a_80_241# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_1267_119# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 COUT a_80_241# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_843_391# CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_385_125# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR B a_385_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 VGND A a_227_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND B a_843_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1195_119# B a_1267_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND B a_385_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR A a_227_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_227_367# B a_80_241# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_80_241# CIN a_385_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_843_391# a_80_241# a_1101_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VPWR A a_843_391# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_1101_119# CIN a_1195_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_843_119# CIN VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_80_241# CIN a_385_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_843_119# a_80_241# a_1101_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR B a_843_391# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 VPWR a_1101_119# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
