* File: sky130_fd_sc_lp__o21a_2.spice
* Created: Fri Aug 28 11:03:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21a_2.pex.spice"
.subckt sky130_fd_sc_lp__o21a_2  VNB VPB B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_X_M1004_d N_A_86_21#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_X_M1004_d N_A_86_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_392_51#_M1000_d N_B1_M1000_g N_A_86_21#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_392_51#_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1002 N_A_392_51#_M1002_d N_A1_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1344 PD=2.21 PS=1.16 NRD=0 NRS=2.856 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_X_M1003_d N_A_86_21#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1008 N_X_M1003_d N_A_86_21#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.504 PD=1.54 PS=2.06 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6 SB=75002
+ A=0.189 P=2.82 MULT=1
MM1001 N_A_86_21#_M1001_d N_B1_M1001_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.504 PD=1.54 PS=2.06 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6 SB=75001.1
+ A=0.189 P=2.82 MULT=1
MM1009 A_478_367# N_A2_M1009_g N_A_86_21#_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=16.4101 NRS=0 M=1 R=8.4 SA=75002
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g A_478_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2016 PD=3.05 PS=1.58 NRD=0 NRS=16.4101 M=1 R=8.4 SA=75002.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o21a_2.pxi.spice"
*
.ends
*
*
