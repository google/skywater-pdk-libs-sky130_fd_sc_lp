* File: sky130_fd_sc_lp__clkbuflp_2.pxi.spice
* Created: Fri Aug 28 10:15:45 2020
* 
x_PM_SKY130_FD_SC_LP__CLKBUFLP_2%A N_A_c_41_n N_A_M1003_g N_A_M1001_g N_A_c_43_n
+ N_A_M1000_g A A N_A_c_45_n PM_SKY130_FD_SC_LP__CLKBUFLP_2%A
x_PM_SKY130_FD_SC_LP__CLKBUFLP_2%A_27_47# N_A_27_47#_M1003_s N_A_27_47#_M1001_s
+ N_A_27_47#_M1002_g N_A_27_47#_M1005_g N_A_27_47#_M1004_g N_A_27_47#_M1008_g
+ N_A_27_47#_M1006_g N_A_27_47#_M1007_g N_A_27_47#_c_86_n N_A_27_47#_c_92_n
+ N_A_27_47#_c_87_n N_A_27_47#_c_88_n N_A_27_47#_c_89_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_2%A_27_47#
x_PM_SKY130_FD_SC_LP__CLKBUFLP_2%VPWR N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_c_156_n N_VPWR_c_157_n N_VPWR_c_158_n N_VPWR_c_159_n VPWR
+ N_VPWR_c_160_n N_VPWR_c_161_n N_VPWR_c_155_n N_VPWR_c_163_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_2%VPWR
x_PM_SKY130_FD_SC_LP__CLKBUFLP_2%X N_X_M1004_s N_X_M1002_s N_X_c_191_n X X X X
+ N_X_c_188_n X PM_SKY130_FD_SC_LP__CLKBUFLP_2%X
x_PM_SKY130_FD_SC_LP__CLKBUFLP_2%VGND N_VGND_M1000_d N_VGND_M1007_d
+ N_VGND_c_221_n N_VGND_c_222_n VGND N_VGND_c_223_n N_VGND_c_224_n
+ N_VGND_c_225_n N_VGND_c_226_n N_VGND_c_227_n N_VGND_c_228_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_2%VGND
cc_1 VNB N_A_c_41_n 0.019034f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.775
cc_2 VNB N_A_M1001_g 0.0378259f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.585
cc_3 VNB N_A_c_43_n 0.0159515f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.775
cc_4 VNB A 0.00518384f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.84
cc_5 VNB N_A_c_45_n 0.0379586f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.94
cc_6 VNB N_A_27_47#_M1002_g 0.00688641f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.445
cc_7 VNB N_A_27_47#_M1005_g 0.035638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_M1004_g 0.0341497f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.94
cc_9 VNB N_A_27_47#_M1008_g 0.00745847f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.94
cc_10 VNB N_A_27_47#_M1006_g 0.0317695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1007_g 0.0544535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_86_n 0.0489388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_87_n 0.0049056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_88_n 0.0224862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_89_n 0.111813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_155_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_X_c_188_n 0.0117552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_221_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.445
cc_19 VNB N_VGND_c_222_n 0.0185162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_223_n 0.0266942f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.94
cc_21 VNB N_VGND_c_224_n 0.0310424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_225_n 0.0201227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_226_n 0.207405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_227_n 0.00436918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_228_n 0.00510891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VPB N_A_M1001_g 0.0505034f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.585
cc_27 VPB N_A_27_47#_M1002_g 0.0412807f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.445
cc_28 VPB N_A_27_47#_M1008_g 0.0516166f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.94
cc_29 VPB N_A_27_47#_c_92_n 0.0496575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_A_27_47#_c_88_n 0.0163566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_156_n 0.00451604f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.445
cc_32 VPB N_VPWR_c_157_n 0.0437034f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.94
cc_33 VPB N_VPWR_c_158_n 0.0240299f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.94
cc_34 VPB N_VPWR_c_159_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.94
cc_35 VPB N_VPWR_c_160_n 0.0175811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_161_n 0.0387386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_155_n 0.0961094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_163_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB X 0.017829f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.94
cc_40 VPB N_X_c_188_n 0.00257184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 N_A_M1001_g N_A_27_47#_M1002_g 0.0315964f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_42 N_A_c_43_n N_A_27_47#_M1005_g 0.0254156f $X=0.835 $Y=0.775 $X2=0 $Y2=0
cc_43 A N_A_27_47#_M1005_g 0.0149455f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_44 N_A_c_45_n N_A_27_47#_M1005_g 0.0062355f $X=0.72 $Y=0.94 $X2=0 $Y2=0
cc_45 A N_A_27_47#_M1004_g 9.69255e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_46 N_A_c_41_n N_A_27_47#_c_86_n 0.0152463f $X=0.475 $Y=0.775 $X2=0 $Y2=0
cc_47 N_A_M1001_g N_A_27_47#_c_86_n 0.00615549f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_48 A N_A_27_47#_c_86_n 0.0260286f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_49 N_A_M1001_g N_A_27_47#_c_92_n 0.0273906f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_50 N_A_M1001_g N_A_27_47#_c_87_n 0.0217094f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_51 A N_A_27_47#_c_87_n 0.0542086f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_52 N_A_c_45_n N_A_27_47#_c_87_n 4.02914e-19 $X=0.72 $Y=0.94 $X2=0 $Y2=0
cc_53 N_A_M1001_g N_A_27_47#_c_88_n 0.0200833f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_54 A N_A_27_47#_c_88_n 0.00528913f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_55 N_A_c_45_n N_A_27_47#_c_88_n 0.00858934f $X=0.72 $Y=0.94 $X2=0 $Y2=0
cc_56 N_A_M1001_g N_A_27_47#_c_89_n 0.0229188f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_57 A N_A_27_47#_c_89_n 0.00363089f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_58 N_A_M1001_g N_VPWR_c_156_n 0.0242966f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VPWR_c_158_n 0.00839865f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_60 N_A_M1001_g N_VPWR_c_155_n 0.0147894f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_X_c_191_n 2.45109e-19 $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_62 N_A_M1001_g X 0.0016204f $X=0.72 $Y=2.585 $X2=0 $Y2=0
cc_63 A N_X_c_188_n 0.0217535f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_64 N_A_c_41_n N_VGND_c_221_n 0.00223338f $X=0.475 $Y=0.775 $X2=0 $Y2=0
cc_65 N_A_c_43_n N_VGND_c_221_n 0.0114645f $X=0.835 $Y=0.775 $X2=0 $Y2=0
cc_66 A N_VGND_c_221_n 0.022081f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A_c_41_n N_VGND_c_223_n 0.00585385f $X=0.475 $Y=0.775 $X2=0 $Y2=0
cc_68 N_A_c_43_n N_VGND_c_223_n 0.00486043f $X=0.835 $Y=0.775 $X2=0 $Y2=0
cc_69 N_A_c_45_n N_VGND_c_223_n 5.88488e-19 $X=0.72 $Y=0.94 $X2=0 $Y2=0
cc_70 N_A_c_41_n N_VGND_c_226_n 0.0117282f $X=0.475 $Y=0.775 $X2=0 $Y2=0
cc_71 N_A_c_43_n N_VGND_c_226_n 0.00427207f $X=0.835 $Y=0.775 $X2=0 $Y2=0
cc_72 A N_VGND_c_226_n 0.0158594f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_73 N_A_c_45_n N_VGND_c_226_n 7.97054e-19 $X=0.72 $Y=0.94 $X2=0 $Y2=0
cc_74 N_A_27_47#_M1002_g N_VPWR_c_156_n 0.0221364f $X=1.25 $Y=2.585 $X2=0 $Y2=0
cc_75 N_A_27_47#_M1008_g N_VPWR_c_156_n 0.00115344f $X=1.78 $Y=2.585 $X2=0 $Y2=0
cc_76 N_A_27_47#_c_92_n N_VPWR_c_156_n 0.0665496f $X=0.455 $Y=2.23 $X2=0 $Y2=0
cc_77 N_A_27_47#_c_87_n N_VPWR_c_156_n 0.0122463f $X=1.22 $Y=1.38 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_89_n N_VPWR_c_156_n 0.00130351f $X=2.415 $Y=1.375 $X2=0 $Y2=0
cc_79 N_A_27_47#_M1002_g N_VPWR_c_157_n 9.25377e-19 $X=1.25 $Y=2.585 $X2=0 $Y2=0
cc_80 N_A_27_47#_M1008_g N_VPWR_c_157_n 0.0236177f $X=1.78 $Y=2.585 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_89_n N_VPWR_c_157_n 0.00109948f $X=2.415 $Y=1.375 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_92_n N_VPWR_c_158_n 0.0210467f $X=0.455 $Y=2.23 $X2=0 $Y2=0
cc_83 N_A_27_47#_M1002_g N_VPWR_c_160_n 0.00794322f $X=1.25 $Y=2.585 $X2=0 $Y2=0
cc_84 N_A_27_47#_M1008_g N_VPWR_c_160_n 0.00839865f $X=1.78 $Y=2.585 $X2=0 $Y2=0
cc_85 N_A_27_47#_M1001_s N_VPWR_c_155_n 0.00212301f $X=0.33 $Y=2.085 $X2=0 $Y2=0
cc_86 N_A_27_47#_M1002_g N_VPWR_c_155_n 0.012523f $X=1.25 $Y=2.585 $X2=0 $Y2=0
cc_87 N_A_27_47#_M1008_g N_VPWR_c_155_n 0.0136348f $X=1.78 $Y=2.585 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_92_n N_VPWR_c_155_n 0.0125689f $X=0.455 $Y=2.23 $X2=0 $Y2=0
cc_89 N_A_27_47#_M1002_g N_X_c_191_n 0.0258353f $X=1.25 $Y=2.585 $X2=0 $Y2=0
cc_90 N_A_27_47#_M1008_g N_X_c_191_n 0.0294899f $X=1.78 $Y=2.585 $X2=0 $Y2=0
cc_91 N_A_27_47#_M1002_g X 0.00691419f $X=1.25 $Y=2.585 $X2=0 $Y2=0
cc_92 N_A_27_47#_M1008_g X 0.0204325f $X=1.78 $Y=2.585 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_87_n X 0.00506752f $X=1.22 $Y=1.38 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_89_n X 0.00440205f $X=2.415 $Y=1.375 $X2=0 $Y2=0
cc_95 N_A_27_47#_M1002_g N_X_c_188_n 0.0043779f $X=1.25 $Y=2.585 $X2=0 $Y2=0
cc_96 N_A_27_47#_M1005_g N_X_c_188_n 0.00387231f $X=1.265 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_27_47#_M1004_g N_X_c_188_n 0.0291408f $X=1.625 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_27_47#_M1008_g N_X_c_188_n 0.00800349f $X=1.78 $Y=2.585 $X2=0 $Y2=0
cc_99 N_A_27_47#_M1006_g N_X_c_188_n 0.0264249f $X=2.055 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_27_47#_M1007_g N_X_c_188_n 0.0205347f $X=2.415 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_87_n N_X_c_188_n 0.0218147f $X=1.22 $Y=1.38 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_89_n N_X_c_188_n 0.057353f $X=2.415 $Y=1.375 $X2=0 $Y2=0
cc_103 N_A_27_47#_M1005_g N_VGND_c_221_n 0.0104103f $X=1.265 $Y=0.445 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_M1004_g N_VGND_c_221_n 0.00214138f $X=1.625 $Y=0.445 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_M1006_g N_VGND_c_222_n 0.00155937f $X=2.055 $Y=0.445 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_M1007_g N_VGND_c_222_n 0.0114035f $X=2.415 $Y=0.445 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_86_n N_VGND_c_223_n 0.0174096f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_108 N_A_27_47#_M1005_g N_VGND_c_224_n 0.00486043f $X=1.265 $Y=0.445 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_M1004_g N_VGND_c_224_n 0.00368782f $X=1.625 $Y=0.445 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_M1006_g N_VGND_c_224_n 0.00359757f $X=2.055 $Y=0.445 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_M1007_g N_VGND_c_224_n 0.00486043f $X=2.415 $Y=0.445 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_M1003_s N_VGND_c_226_n 0.00302351f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_M1005_g N_VGND_c_226_n 0.00473304f $X=1.265 $Y=0.445 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_M1004_g N_VGND_c_226_n 0.00542579f $X=1.625 $Y=0.445 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_M1006_g N_VGND_c_226_n 0.0052035f $X=2.055 $Y=0.445 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_M1007_g N_VGND_c_226_n 0.00814425f $X=2.415 $Y=0.445 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_c_86_n N_VGND_c_226_n 0.0107567f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_118 N_VPWR_c_155_n N_X_M1002_s 0.00223559f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_119 N_VPWR_c_156_n N_X_c_191_n 0.0763033f $X=0.985 $Y=2.23 $X2=0 $Y2=0
cc_120 N_VPWR_c_157_n N_X_c_191_n 0.0656691f $X=2.045 $Y=2.23 $X2=0 $Y2=0
cc_121 N_VPWR_c_160_n N_X_c_191_n 0.0209688f $X=1.88 $Y=3.33 $X2=0 $Y2=0
cc_122 N_VPWR_c_155_n N_X_c_191_n 0.013415f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_123 N_VPWR_c_157_n X 0.023516f $X=2.045 $Y=2.23 $X2=0 $Y2=0
cc_124 N_X_c_188_n N_VGND_c_221_n 0.0155556f $X=1.84 $Y=0.44 $X2=0 $Y2=0
cc_125 N_X_c_188_n N_VGND_c_222_n 0.0252484f $X=1.84 $Y=0.44 $X2=0 $Y2=0
cc_126 N_X_c_188_n N_VGND_c_224_n 0.0408566f $X=1.84 $Y=0.44 $X2=0 $Y2=0
cc_127 N_X_M1004_s N_VGND_c_226_n 0.00223819f $X=1.7 $Y=0.235 $X2=0 $Y2=0
cc_128 N_X_c_188_n N_VGND_c_226_n 0.0260885f $X=1.84 $Y=0.44 $X2=0 $Y2=0
cc_129 N_X_c_188_n A_426_47# 0.00452967f $X=1.84 $Y=0.44 $X2=-0.19 $Y2=-0.245
cc_130 A_110_47# N_VGND_c_226_n 0.00302274f $X=0.55 $Y=0.235 $X2=3.12 $Y2=0
cc_131 N_VGND_c_226_n A_268_47# 0.00899413f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_132 N_VGND_c_226_n A_426_47# 0.00415997f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
