* File: sky130_fd_sc_lp__and3b_lp.pxi.spice
* Created: Wed Sep  2 09:32:25 2020
* 
x_PM_SKY130_FD_SC_LP__AND3B_LP%A_N N_A_N_c_81_n N_A_N_M1005_g N_A_N_M1009_g
+ N_A_N_c_83_n N_A_N_c_84_n N_A_N_M1011_g N_A_N_c_85_n N_A_N_c_86_n A_N A_N
+ N_A_N_c_87_n N_A_N_c_88_n PM_SKY130_FD_SC_LP__AND3B_LP%A_N
x_PM_SKY130_FD_SC_LP__AND3B_LP%A_137_408# N_A_137_408#_M1011_d
+ N_A_137_408#_M1009_d N_A_137_408#_M1008_g N_A_137_408#_c_123_n
+ N_A_137_408#_M1001_g N_A_137_408#_c_124_n N_A_137_408#_c_130_n
+ N_A_137_408#_c_131_n N_A_137_408#_c_125_n N_A_137_408#_c_132_n
+ N_A_137_408#_c_126_n N_A_137_408#_c_127_n N_A_137_408#_c_128_n
+ PM_SKY130_FD_SC_LP__AND3B_LP%A_137_408#
x_PM_SKY130_FD_SC_LP__AND3B_LP%B N_B_c_188_n N_B_M1003_g N_B_M1006_g N_B_c_185_n
+ B B N_B_c_186_n N_B_c_187_n PM_SKY130_FD_SC_LP__AND3B_LP%B
x_PM_SKY130_FD_SC_LP__AND3B_LP%C N_C_M1007_g N_C_M1010_g N_C_c_229_n N_C_c_234_n
+ C C N_C_c_231_n PM_SKY130_FD_SC_LP__AND3B_LP%C
x_PM_SKY130_FD_SC_LP__AND3B_LP%A_248_409# N_A_248_409#_M1001_s
+ N_A_248_409#_M1008_s N_A_248_409#_M1003_d N_A_248_409#_c_274_n
+ N_A_248_409#_M1000_g N_A_248_409#_M1004_g N_A_248_409#_c_276_n
+ N_A_248_409#_M1002_g N_A_248_409#_c_286_n N_A_248_409#_c_277_n
+ N_A_248_409#_c_287_n N_A_248_409#_c_288_n N_A_248_409#_c_278_n
+ N_A_248_409#_c_279_n N_A_248_409#_c_289_n N_A_248_409#_c_290_n
+ N_A_248_409#_c_280_n N_A_248_409#_c_281_n N_A_248_409#_c_282_n
+ N_A_248_409#_c_292_n N_A_248_409#_c_283_n N_A_248_409#_c_284_n
+ PM_SKY130_FD_SC_LP__AND3B_LP%A_248_409#
x_PM_SKY130_FD_SC_LP__AND3B_LP%VPWR N_VPWR_M1009_s N_VPWR_M1008_d N_VPWR_M1010_d
+ N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n
+ N_VPWR_c_393_n VPWR N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_387_n
+ N_VPWR_c_397_n PM_SKY130_FD_SC_LP__AND3B_LP%VPWR
x_PM_SKY130_FD_SC_LP__AND3B_LP%X N_X_M1002_d N_X_M1004_d N_X_c_434_n X X X X X X
+ PM_SKY130_FD_SC_LP__AND3B_LP%X
x_PM_SKY130_FD_SC_LP__AND3B_LP%VGND N_VGND_M1005_s N_VGND_M1007_d N_VGND_c_461_n
+ N_VGND_c_462_n N_VGND_c_463_n N_VGND_c_464_n N_VGND_c_465_n VGND
+ N_VGND_c_466_n N_VGND_c_467_n PM_SKY130_FD_SC_LP__AND3B_LP%VGND
cc_1 VNB N_A_N_c_81_n 0.0177984f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.78
cc_2 VNB N_A_N_M1009_g 0.00611216f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.54
cc_3 VNB N_A_N_c_83_n 0.0249772f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.855
cc_4 VNB N_A_N_c_84_n 0.0177835f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.78
cc_5 VNB N_A_N_c_85_n 0.022979f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=0.855
cc_6 VNB N_A_N_c_86_n 0.0317491f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.575
cc_7 VNB N_A_N_c_87_n 0.0628848f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_8 VNB N_A_N_c_88_n 0.00298149f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.07
cc_9 VNB N_A_137_408#_c_123_n 0.0180638f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=0.93
cc_10 VNB N_A_137_408#_c_124_n 0.0209739f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A_137_408#_c_125_n 0.0141405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_137_408#_c_126_n 0.00973294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_137_408#_c_127_n 0.0704719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_137_408#_c_128_n 0.015417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_M1006_g 0.0340016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_185_n 0.0185722f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.495
cc_17 VNB N_B_c_186_n 0.0143138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_187_n 0.00486564f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.07
cc_19 VNB N_C_M1007_g 0.035953f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_20 VNB N_C_c_229_n 0.0209572f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.495
cc_21 VNB C 0.00528809f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=0.93
cc_22 VNB N_C_c_231_n 0.0157274f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB N_A_248_409#_c_274_n 0.0176761f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.78
cc_24 VNB N_A_248_409#_M1004_g 0.0106126f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.425
cc_25 VNB N_A_248_409#_c_276_n 0.0198928f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.575
cc_26 VNB N_A_248_409#_c_277_n 0.00712279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_248_409#_c_278_n 0.0289982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_248_409#_c_279_n 0.00319676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_248_409#_c_280_n 0.00230529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_248_409#_c_281_n 0.00300595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_248_409#_c_282_n 0.00100691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_248_409#_c_283_n 0.0777877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_248_409#_c_284_n 0.00143055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_387_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_434_n 0.0388766f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.855
cc_36 VNB X 0.0217459f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.495
cc_37 VNB X 0.0121436f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.495
cc_38 VNB N_VGND_c_461_n 0.0113827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_462_n 0.0242568f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.855
cc_40 VNB N_VGND_c_463_n 0.00424508f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=0.93
cc_41 VNB N_VGND_c_464_n 0.063465f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.425
cc_42 VNB N_VGND_c_465_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.575
cc_43 VNB N_VGND_c_466_n 0.0398494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_467_n 0.274829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A_N_M1009_g 0.0550817f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.54
cc_46 VPB N_A_N_c_88_n 0.00821726f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_47 VPB N_A_137_408#_M1008_g 0.0334232f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.855
cc_48 VPB N_A_137_408#_c_130_n 0.0070336f $X=-0.19 $Y=1.655 $X2=0.355 $Y2=1.07
cc_49 VPB N_A_137_408#_c_131_n 0.0100497f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_50 VPB N_A_137_408#_c_132_n 0.00409336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_137_408#_c_126_n 0.0129427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_137_408#_c_127_n 0.0324078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_B_c_188_n 0.0116807f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.78
cc_54 VPB N_B_M1003_g 0.0283856f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.495
cc_55 VPB N_B_c_185_n 0.00110618f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.495
cc_56 VPB N_B_c_187_n 0.00348556f $X=-0.19 $Y=1.655 $X2=0.355 $Y2=1.07
cc_57 VPB N_C_M1010_g 0.0294875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_C_c_229_n 0.00127079f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.495
cc_59 VPB N_C_c_234_n 0.0132791f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.495
cc_60 VPB C 0.00246418f $X=-0.19 $Y=1.655 $X2=0.355 $Y2=0.93
cc_61 VPB N_A_248_409#_M1004_g 0.0448556f $X=-0.19 $Y=1.655 $X2=0.355 $Y2=1.425
cc_62 VPB N_A_248_409#_c_286_n 0.0100935f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_63 VPB N_A_248_409#_c_287_n 0.00249329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_248_409#_c_288_n 0.00426456f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_248_409#_c_289_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_248_409#_c_290_n 0.00669005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_248_409#_c_282_n 0.00297842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_248_409#_c_292_n 0.00818658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_388_n 0.0117708f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.78
cc_70 VPB N_VPWR_c_389_n 0.0468447f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.495
cc_71 VPB N_VPWR_c_390_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_72 VPB N_VPWR_c_391_n 0.00418937f $X=-0.19 $Y=1.655 $X2=0.355 $Y2=1.07
cc_73 VPB N_VPWR_c_392_n 0.0335618f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.07
cc_74 VPB N_VPWR_c_393_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_394_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_395_n 0.0327924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_387_n 0.0718979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_397_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB X 0.0247296f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.495
cc_80 VPB X 0.067762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 N_A_N_c_83_n N_A_137_408#_c_124_n 0.00164789f $X=0.81 $Y=0.855 $X2=0 $Y2=0
cc_82 N_A_N_M1009_g N_A_137_408#_c_130_n 0.00446174f $X=0.56 $Y=2.54 $X2=0 $Y2=0
cc_83 N_A_N_M1009_g N_A_137_408#_c_131_n 0.0158747f $X=0.56 $Y=2.54 $X2=0 $Y2=0
cc_84 N_A_N_c_81_n N_A_137_408#_c_125_n 0.00190711f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_85 N_A_N_c_83_n N_A_137_408#_c_125_n 0.0146711f $X=0.81 $Y=0.855 $X2=0 $Y2=0
cc_86 N_A_N_c_84_n N_A_137_408#_c_125_n 0.0151837f $X=0.885 $Y=0.78 $X2=0 $Y2=0
cc_87 N_A_N_c_87_n N_A_137_408#_c_125_n 0.00881756f $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_88 N_A_N_c_88_n N_A_137_408#_c_125_n 0.0405655f $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_89 N_A_N_M1009_g N_A_137_408#_c_132_n 0.00631733f $X=0.56 $Y=2.54 $X2=0 $Y2=0
cc_90 N_A_N_c_86_n N_A_137_408#_c_126_n 0.00631733f $X=0.405 $Y=1.575 $X2=0
+ $Y2=0
cc_91 N_A_N_c_86_n N_A_137_408#_c_127_n 0.0120876f $X=0.405 $Y=1.575 $X2=0 $Y2=0
cc_92 N_A_N_c_87_n N_A_137_408#_c_127_n 0.00536727f $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_93 N_A_N_c_88_n N_A_137_408#_c_127_n 4.50434e-19 $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_94 N_A_N_M1009_g N_A_248_409#_c_286_n 0.00168543f $X=0.56 $Y=2.54 $X2=0 $Y2=0
cc_95 N_A_N_c_84_n N_A_248_409#_c_277_n 0.0012685f $X=0.885 $Y=0.78 $X2=0 $Y2=0
cc_96 N_A_N_M1009_g N_A_248_409#_c_288_n 3.95513e-19 $X=0.56 $Y=2.54 $X2=0 $Y2=0
cc_97 N_A_N_c_83_n N_A_248_409#_c_279_n 3.03943e-19 $X=0.81 $Y=0.855 $X2=0 $Y2=0
cc_98 N_A_N_M1009_g N_VPWR_c_389_n 0.0253197f $X=0.56 $Y=2.54 $X2=0 $Y2=0
cc_99 N_A_N_c_86_n N_VPWR_c_389_n 0.00151284f $X=0.405 $Y=1.575 $X2=0 $Y2=0
cc_100 N_A_N_c_88_n N_VPWR_c_389_n 0.023553f $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_101 N_A_N_M1009_g N_VPWR_c_392_n 0.00762416f $X=0.56 $Y=2.54 $X2=0 $Y2=0
cc_102 N_A_N_M1009_g N_VPWR_c_387_n 0.0142699f $X=0.56 $Y=2.54 $X2=0 $Y2=0
cc_103 N_A_N_c_81_n N_VGND_c_462_n 0.0134067f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_104 N_A_N_c_84_n N_VGND_c_462_n 0.00205514f $X=0.885 $Y=0.78 $X2=0 $Y2=0
cc_105 N_A_N_c_85_n N_VGND_c_462_n 0.00930805f $X=0.355 $Y=0.855 $X2=0 $Y2=0
cc_106 N_A_N_c_88_n N_VGND_c_462_n 0.0270319f $X=0.29 $Y=1.07 $X2=0 $Y2=0
cc_107 N_A_N_c_81_n N_VGND_c_464_n 0.00445056f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_108 N_A_N_c_83_n N_VGND_c_464_n 9.15697e-19 $X=0.81 $Y=0.855 $X2=0 $Y2=0
cc_109 N_A_N_c_84_n N_VGND_c_464_n 0.00342832f $X=0.885 $Y=0.78 $X2=0 $Y2=0
cc_110 N_A_N_c_81_n N_VGND_c_467_n 0.00802306f $X=0.495 $Y=0.78 $X2=0 $Y2=0
cc_111 N_A_N_c_83_n N_VGND_c_467_n 0.00126624f $X=0.81 $Y=0.855 $X2=0 $Y2=0
cc_112 N_A_N_c_84_n N_VGND_c_467_n 0.0061026f $X=0.885 $Y=0.78 $X2=0 $Y2=0
cc_113 N_A_137_408#_M1008_g N_B_M1003_g 0.030269f $X=1.65 $Y=2.545 $X2=0 $Y2=0
cc_114 N_A_137_408#_c_123_n N_B_M1006_g 0.0423428f $X=1.88 $Y=0.78 $X2=0 $Y2=0
cc_115 N_A_137_408#_c_128_n N_B_M1006_g 0.00782887f $X=1.415 $Y=1.17 $X2=0 $Y2=0
cc_116 N_A_137_408#_c_126_n N_B_c_186_n 2.62814e-19 $X=1.22 $Y=1.335 $X2=0 $Y2=0
cc_117 N_A_137_408#_c_127_n N_B_c_186_n 0.0369754f $X=1.22 $Y=1.335 $X2=0 $Y2=0
cc_118 N_A_137_408#_c_124_n N_B_c_187_n 0.0012154f $X=1.88 $Y=0.855 $X2=0 $Y2=0
cc_119 N_A_137_408#_c_126_n N_B_c_187_n 0.0529807f $X=1.22 $Y=1.335 $X2=0 $Y2=0
cc_120 N_A_137_408#_c_127_n N_B_c_187_n 0.0358333f $X=1.22 $Y=1.335 $X2=0 $Y2=0
cc_121 N_A_137_408#_M1008_g N_A_248_409#_c_286_n 0.0158404f $X=1.65 $Y=2.545
+ $X2=0 $Y2=0
cc_122 N_A_137_408#_c_131_n N_A_248_409#_c_286_n 0.0586203f $X=0.825 $Y=2.895
+ $X2=0 $Y2=0
cc_123 N_A_137_408#_c_123_n N_A_248_409#_c_277_n 0.0118015f $X=1.88 $Y=0.78
+ $X2=0 $Y2=0
cc_124 N_A_137_408#_c_124_n N_A_248_409#_c_277_n 0.00593998f $X=1.88 $Y=0.855
+ $X2=0 $Y2=0
cc_125 N_A_137_408#_c_125_n N_A_248_409#_c_277_n 0.0376839f $X=1.1 $Y=0.495
+ $X2=0 $Y2=0
cc_126 N_A_137_408#_M1008_g N_A_248_409#_c_287_n 0.0182823f $X=1.65 $Y=2.545
+ $X2=0 $Y2=0
cc_127 N_A_137_408#_M1008_g N_A_248_409#_c_288_n 0.00216931f $X=1.65 $Y=2.545
+ $X2=0 $Y2=0
cc_128 N_A_137_408#_c_130_n N_A_248_409#_c_288_n 0.0121278f $X=0.825 $Y=2.185
+ $X2=0 $Y2=0
cc_129 N_A_137_408#_c_126_n N_A_248_409#_c_288_n 0.0139887f $X=1.22 $Y=1.335
+ $X2=0 $Y2=0
cc_130 N_A_137_408#_c_127_n N_A_248_409#_c_288_n 0.00796888f $X=1.22 $Y=1.335
+ $X2=0 $Y2=0
cc_131 N_A_137_408#_c_124_n N_A_248_409#_c_278_n 0.00713002f $X=1.88 $Y=0.855
+ $X2=0 $Y2=0
cc_132 N_A_137_408#_c_124_n N_A_248_409#_c_279_n 0.00439916f $X=1.88 $Y=0.855
+ $X2=0 $Y2=0
cc_133 N_A_137_408#_c_125_n N_A_248_409#_c_279_n 0.0122422f $X=1.1 $Y=0.495
+ $X2=0 $Y2=0
cc_134 N_A_137_408#_c_127_n N_A_248_409#_c_279_n 0.00472649f $X=1.22 $Y=1.335
+ $X2=0 $Y2=0
cc_135 N_A_137_408#_c_128_n N_A_248_409#_c_279_n 0.00499769f $X=1.415 $Y=1.17
+ $X2=0 $Y2=0
cc_136 N_A_137_408#_M1008_g N_A_248_409#_c_289_n 8.94979e-19 $X=1.65 $Y=2.545
+ $X2=0 $Y2=0
cc_137 N_A_137_408#_c_130_n N_VPWR_c_389_n 0.0684934f $X=0.825 $Y=2.185 $X2=0
+ $Y2=0
cc_138 N_A_137_408#_M1008_g N_VPWR_c_390_n 0.0174514f $X=1.65 $Y=2.545 $X2=0
+ $Y2=0
cc_139 N_A_137_408#_M1008_g N_VPWR_c_392_n 0.00769046f $X=1.65 $Y=2.545 $X2=0
+ $Y2=0
cc_140 N_A_137_408#_c_131_n N_VPWR_c_392_n 0.021393f $X=0.825 $Y=2.895 $X2=0
+ $Y2=0
cc_141 N_A_137_408#_M1008_g N_VPWR_c_387_n 0.0143431f $X=1.65 $Y=2.545 $X2=0
+ $Y2=0
cc_142 N_A_137_408#_c_131_n N_VPWR_c_387_n 0.0125495f $X=0.825 $Y=2.895 $X2=0
+ $Y2=0
cc_143 N_A_137_408#_c_125_n N_VGND_c_462_n 0.0187024f $X=1.1 $Y=0.495 $X2=0
+ $Y2=0
cc_144 N_A_137_408#_c_123_n N_VGND_c_464_n 0.00502664f $X=1.88 $Y=0.78 $X2=0
+ $Y2=0
cc_145 N_A_137_408#_c_124_n N_VGND_c_464_n 3.83046e-19 $X=1.88 $Y=0.855 $X2=0
+ $Y2=0
cc_146 N_A_137_408#_c_125_n N_VGND_c_464_n 0.0293877f $X=1.1 $Y=0.495 $X2=0
+ $Y2=0
cc_147 N_A_137_408#_c_123_n N_VGND_c_467_n 0.00659248f $X=1.88 $Y=0.78 $X2=0
+ $Y2=0
cc_148 N_A_137_408#_c_125_n N_VGND_c_467_n 0.0165008f $X=1.1 $Y=0.495 $X2=0
+ $Y2=0
cc_149 N_B_M1006_g N_C_M1007_g 0.0233696f $X=2.27 $Y=0.495 $X2=0 $Y2=0
cc_150 N_B_M1003_g N_C_M1010_g 0.0173741f $X=2.18 $Y=2.545 $X2=0 $Y2=0
cc_151 N_B_c_185_n N_C_c_229_n 0.0233696f $X=2.18 $Y=1.675 $X2=0 $Y2=0
cc_152 N_B_c_188_n N_C_c_234_n 0.0233696f $X=2.18 $Y=1.84 $X2=0 $Y2=0
cc_153 N_B_c_186_n C 0.00235811f $X=2.18 $Y=1.335 $X2=0 $Y2=0
cc_154 N_B_c_187_n C 0.0542827f $X=2.18 $Y=1.335 $X2=0 $Y2=0
cc_155 N_B_c_186_n N_C_c_231_n 0.0233696f $X=2.18 $Y=1.335 $X2=0 $Y2=0
cc_156 N_B_c_187_n N_C_c_231_n 7.48751e-19 $X=2.18 $Y=1.335 $X2=0 $Y2=0
cc_157 N_B_M1003_g N_A_248_409#_c_286_n 8.94979e-19 $X=2.18 $Y=2.545 $X2=0 $Y2=0
cc_158 N_B_M1006_g N_A_248_409#_c_277_n 0.00274521f $X=2.27 $Y=0.495 $X2=0 $Y2=0
cc_159 N_B_c_188_n N_A_248_409#_c_287_n 0.00103139f $X=2.18 $Y=1.84 $X2=0 $Y2=0
cc_160 N_B_M1003_g N_A_248_409#_c_287_n 0.0178604f $X=2.18 $Y=2.545 $X2=0 $Y2=0
cc_161 N_B_c_187_n N_A_248_409#_c_287_n 0.0538265f $X=2.18 $Y=1.335 $X2=0 $Y2=0
cc_162 N_B_M1006_g N_A_248_409#_c_278_n 0.0116782f $X=2.27 $Y=0.495 $X2=0 $Y2=0
cc_163 N_B_c_186_n N_A_248_409#_c_278_n 0.00469578f $X=2.18 $Y=1.335 $X2=0 $Y2=0
cc_164 N_B_c_187_n N_A_248_409#_c_278_n 0.0394278f $X=2.18 $Y=1.335 $X2=0 $Y2=0
cc_165 N_B_c_187_n N_A_248_409#_c_279_n 0.0220658f $X=2.18 $Y=1.335 $X2=0 $Y2=0
cc_166 N_B_M1003_g N_A_248_409#_c_289_n 0.0156803f $X=2.18 $Y=2.545 $X2=0 $Y2=0
cc_167 N_B_c_188_n N_A_248_409#_c_292_n 0.00108331f $X=2.18 $Y=1.84 $X2=0 $Y2=0
cc_168 N_B_M1003_g N_A_248_409#_c_292_n 0.00104211f $X=2.18 $Y=2.545 $X2=0 $Y2=0
cc_169 N_B_c_187_n N_A_248_409#_c_292_n 0.00540441f $X=2.18 $Y=1.335 $X2=0 $Y2=0
cc_170 N_B_M1003_g N_VPWR_c_390_n 0.0164386f $X=2.18 $Y=2.545 $X2=0 $Y2=0
cc_171 N_B_M1003_g N_VPWR_c_391_n 8.50498e-19 $X=2.18 $Y=2.545 $X2=0 $Y2=0
cc_172 N_B_M1003_g N_VPWR_c_394_n 0.00769046f $X=2.18 $Y=2.545 $X2=0 $Y2=0
cc_173 N_B_M1003_g N_VPWR_c_387_n 0.0134474f $X=2.18 $Y=2.545 $X2=0 $Y2=0
cc_174 N_B_M1006_g N_VGND_c_463_n 0.00268914f $X=2.27 $Y=0.495 $X2=0 $Y2=0
cc_175 N_B_M1006_g N_VGND_c_464_n 0.0053602f $X=2.27 $Y=0.495 $X2=0 $Y2=0
cc_176 N_B_M1006_g N_VGND_c_467_n 0.00582628f $X=2.27 $Y=0.495 $X2=0 $Y2=0
cc_177 N_C_M1007_g N_A_248_409#_c_274_n 0.012269f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_178 N_C_M1010_g N_A_248_409#_M1004_g 0.0271467f $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_179 N_C_c_229_n N_A_248_409#_M1004_g 0.0133955f $X=2.75 $Y=1.675 $X2=0 $Y2=0
cc_180 C N_A_248_409#_M1004_g 3.63567e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_181 N_C_M1007_g N_A_248_409#_c_278_n 0.0120711f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_182 C N_A_248_409#_c_278_n 0.0293571f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_183 N_C_c_231_n N_A_248_409#_c_278_n 0.00123061f $X=2.75 $Y=1.335 $X2=0 $Y2=0
cc_184 N_C_M1010_g N_A_248_409#_c_289_n 0.0161384f $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_185 N_C_M1010_g N_A_248_409#_c_290_n 0.0183402f $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_186 N_C_c_234_n N_A_248_409#_c_290_n 5.43485e-19 $X=2.75 $Y=1.84 $X2=0 $Y2=0
cc_187 C N_A_248_409#_c_290_n 0.0223517f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_188 N_C_M1007_g N_A_248_409#_c_281_n 0.00367096f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_189 C N_A_248_409#_c_281_n 0.0502547f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_190 N_C_c_231_n N_A_248_409#_c_281_n 0.00141048f $X=2.75 $Y=1.335 $X2=0 $Y2=0
cc_191 N_C_M1010_g N_A_248_409#_c_282_n 0.00356794f $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_192 N_C_c_234_n N_A_248_409#_c_282_n 0.00141048f $X=2.75 $Y=1.84 $X2=0 $Y2=0
cc_193 N_C_M1010_g N_A_248_409#_c_292_n 0.00104103f $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_194 C N_A_248_409#_c_292_n 0.00731937f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_195 N_C_M1007_g N_A_248_409#_c_283_n 0.00874737f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_196 C N_A_248_409#_c_283_n 3.61519e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_197 N_C_c_231_n N_A_248_409#_c_283_n 0.0169083f $X=2.75 $Y=1.335 $X2=0 $Y2=0
cc_198 N_C_c_229_n N_A_248_409#_c_284_n 0.00141048f $X=2.75 $Y=1.675 $X2=0 $Y2=0
cc_199 N_C_M1010_g N_VPWR_c_390_n 8.50498e-19 $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_200 N_C_M1010_g N_VPWR_c_391_n 0.0165581f $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_201 N_C_M1010_g N_VPWR_c_394_n 0.00769046f $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_202 N_C_M1010_g N_VPWR_c_387_n 0.0134474f $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_203 N_C_M1010_g X 9.7864e-19 $X=2.71 $Y=2.545 $X2=0 $Y2=0
cc_204 N_C_M1007_g N_VGND_c_463_n 0.01151f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_205 N_C_M1007_g N_VGND_c_464_n 0.00445056f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_206 N_C_M1007_g N_VGND_c_467_n 0.00426841f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_207 N_A_248_409#_c_287_n N_VPWR_M1008_d 0.00180746f $X=2.28 $Y=2.105 $X2=0
+ $Y2=0
cc_208 N_A_248_409#_c_290_n N_VPWR_M1010_d 0.0039802f $X=3.095 $Y=2.105 $X2=0
+ $Y2=0
cc_209 N_A_248_409#_c_286_n N_VPWR_c_390_n 0.045794f $X=1.385 $Y=2.9 $X2=0 $Y2=0
cc_210 N_A_248_409#_c_287_n N_VPWR_c_390_n 0.0163515f $X=2.28 $Y=2.105 $X2=0
+ $Y2=0
cc_211 N_A_248_409#_c_289_n N_VPWR_c_390_n 0.045794f $X=2.445 $Y=2.9 $X2=0 $Y2=0
cc_212 N_A_248_409#_M1004_g N_VPWR_c_391_n 0.0102656f $X=3.345 $Y=2.545 $X2=0
+ $Y2=0
cc_213 N_A_248_409#_c_289_n N_VPWR_c_391_n 0.045794f $X=2.445 $Y=2.9 $X2=0 $Y2=0
cc_214 N_A_248_409#_c_290_n N_VPWR_c_391_n 0.0212953f $X=3.095 $Y=2.105 $X2=0
+ $Y2=0
cc_215 N_A_248_409#_c_286_n N_VPWR_c_392_n 0.0220321f $X=1.385 $Y=2.9 $X2=0
+ $Y2=0
cc_216 N_A_248_409#_c_289_n N_VPWR_c_394_n 0.021949f $X=2.445 $Y=2.9 $X2=0 $Y2=0
cc_217 N_A_248_409#_M1004_g N_VPWR_c_395_n 0.0086001f $X=3.345 $Y=2.545 $X2=0
+ $Y2=0
cc_218 N_A_248_409#_M1004_g N_VPWR_c_387_n 0.0168033f $X=3.345 $Y=2.545 $X2=0
+ $Y2=0
cc_219 N_A_248_409#_c_286_n N_VPWR_c_387_n 0.0125808f $X=1.385 $Y=2.9 $X2=0
+ $Y2=0
cc_220 N_A_248_409#_c_289_n N_VPWR_c_387_n 0.0124703f $X=2.445 $Y=2.9 $X2=0
+ $Y2=0
cc_221 N_A_248_409#_c_274_n N_X_c_434_n 0.00200943f $X=3.255 $Y=0.82 $X2=0 $Y2=0
cc_222 N_A_248_409#_c_276_n N_X_c_434_n 0.0135409f $X=3.615 $Y=0.82 $X2=0 $Y2=0
cc_223 N_A_248_409#_c_280_n N_X_c_434_n 0.0129587f $X=3.29 $Y=0.99 $X2=0 $Y2=0
cc_224 N_A_248_409#_c_281_n N_X_c_434_n 0.0184961f $X=3.29 $Y=1.295 $X2=0 $Y2=0
cc_225 N_A_248_409#_c_283_n N_X_c_434_n 0.0132611f $X=3.32 $Y=0.985 $X2=0 $Y2=0
cc_226 N_A_248_409#_c_283_n X 0.0105016f $X=3.32 $Y=0.985 $X2=0 $Y2=0
cc_227 N_A_248_409#_c_284_n X 0.0184961f $X=3.29 $Y=1.49 $X2=0 $Y2=0
cc_228 N_A_248_409#_M1004_g X 0.0129763f $X=3.345 $Y=2.545 $X2=0 $Y2=0
cc_229 N_A_248_409#_c_290_n X 2.04298e-19 $X=3.095 $Y=2.105 $X2=0 $Y2=0
cc_230 N_A_248_409#_c_282_n X 0.0220582f $X=3.18 $Y=2.02 $X2=0 $Y2=0
cc_231 N_A_248_409#_c_283_n X 0.00234697f $X=3.32 $Y=0.985 $X2=0 $Y2=0
cc_232 N_A_248_409#_M1004_g X 0.0197318f $X=3.345 $Y=2.545 $X2=0 $Y2=0
cc_233 N_A_248_409#_c_290_n X 0.0132745f $X=3.095 $Y=2.105 $X2=0 $Y2=0
cc_234 N_A_248_409#_c_283_n X 0.00607155f $X=3.32 $Y=0.985 $X2=0 $Y2=0
cc_235 N_A_248_409#_c_284_n X 0.00131253f $X=3.29 $Y=1.49 $X2=0 $Y2=0
cc_236 N_A_248_409#_c_274_n N_VGND_c_463_n 0.00741322f $X=3.255 $Y=0.82 $X2=0
+ $Y2=0
cc_237 N_A_248_409#_c_278_n N_VGND_c_463_n 0.0226313f $X=3.095 $Y=0.905 $X2=0
+ $Y2=0
cc_238 N_A_248_409#_c_277_n N_VGND_c_464_n 0.0220321f $X=1.665 $Y=0.495 $X2=0
+ $Y2=0
cc_239 N_A_248_409#_c_274_n N_VGND_c_466_n 0.0053602f $X=3.255 $Y=0.82 $X2=0
+ $Y2=0
cc_240 N_A_248_409#_c_276_n N_VGND_c_466_n 0.00502664f $X=3.615 $Y=0.82 $X2=0
+ $Y2=0
cc_241 N_A_248_409#_c_274_n N_VGND_c_467_n 0.00604995f $X=3.255 $Y=0.82 $X2=0
+ $Y2=0
cc_242 N_A_248_409#_c_276_n N_VGND_c_467_n 0.0101575f $X=3.615 $Y=0.82 $X2=0
+ $Y2=0
cc_243 N_A_248_409#_c_277_n N_VGND_c_467_n 0.0125808f $X=1.665 $Y=0.495 $X2=0
+ $Y2=0
cc_244 N_A_248_409#_c_278_n N_VGND_c_467_n 0.0311385f $X=3.095 $Y=0.905 $X2=0
+ $Y2=0
cc_245 N_A_248_409#_c_280_n N_VGND_c_467_n 0.0137708f $X=3.29 $Y=0.99 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_391_n X 0.036413f $X=2.975 $Y=2.535 $X2=0 $Y2=0
cc_247 N_VPWR_c_395_n X 0.0503504f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_248 N_VPWR_c_387_n X 0.0288319f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_249 N_X_c_434_n N_VGND_c_463_n 0.0104189f $X=3.83 $Y=0.495 $X2=0 $Y2=0
cc_250 N_X_c_434_n N_VGND_c_466_n 0.0220321f $X=3.83 $Y=0.495 $X2=0 $Y2=0
cc_251 N_X_c_434_n N_VGND_c_467_n 0.0125808f $X=3.83 $Y=0.495 $X2=0 $Y2=0
