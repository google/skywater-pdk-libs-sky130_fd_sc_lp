# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o221a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o221a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.370000 1.075000 5.030000 1.245000 ;
        RECT 3.370000 1.245000 3.690000 1.515000 ;
        RECT 4.465000 1.245000 5.030000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.860000 1.425000 4.295000 1.760000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.210000 3.155000 1.245000 ;
        RECT 1.035000 1.245000 1.820000 1.605000 ;
        RECT 1.595000 1.075000 3.155000 1.210000 ;
        RECT 2.905000 1.245000 3.155000 1.605000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.425000 2.735000 1.760000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.350000 1.350000 ;
        RECT 0.085000 1.350000 0.435000 1.785000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.465000 0.255000 5.695000 1.045000 ;
        RECT 5.465000 1.045000 7.115000 1.215000 ;
        RECT 5.540000 1.755000 7.115000 1.925000 ;
        RECT 5.540000 1.925000 5.730000 3.075000 ;
        RECT 6.365000 0.255000 6.555000 1.045000 ;
        RECT 6.400000 1.925000 6.590000 3.075000 ;
        RECT 6.865000 1.215000 7.115000 1.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
        RECT 3.245000  0.085000 3.575000 0.540000 ;
        RECT 4.105000  0.085000 4.435000 0.540000 ;
        RECT 5.035000  0.085000 5.295000 0.905000 ;
        RECT 5.865000  0.085000 6.195000 0.865000 ;
        RECT 6.725000  0.085000 7.055000 0.875000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.200000 3.415000 ;
        RECT 0.105000 1.955000 0.435000 3.245000 ;
        RECT 0.985000 2.270000 1.315000 3.245000 ;
        RECT 2.725000 2.270000 3.505000 3.245000 ;
        RECT 4.970000 2.270000 5.300000 3.245000 ;
        RECT 5.900000 2.105000 6.230000 3.245000 ;
        RECT 6.760000 2.105000 7.090000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105000 0.255000 3.055000 0.425000 ;
      RECT 0.105000 0.425000 0.365000 1.040000 ;
      RECT 0.535000 0.595000 0.865000 1.145000 ;
      RECT 0.605000 1.145000 0.865000 1.930000 ;
      RECT 0.605000 1.930000 5.370000 2.100000 ;
      RECT 0.605000 2.100000 0.815000 3.075000 ;
      RECT 1.035000 0.425000 3.055000 0.540000 ;
      RECT 1.035000 0.540000 1.265000 0.975000 ;
      RECT 1.435000 0.710000 2.645000 0.725000 ;
      RECT 1.435000 0.725000 4.865000 0.905000 ;
      RECT 1.485000 2.270000 1.695000 2.905000 ;
      RECT 1.485000 2.905000 2.555000 3.075000 ;
      RECT 1.865000 2.100000 2.195000 2.735000 ;
      RECT 2.365000 2.270000 2.555000 2.905000 ;
      RECT 2.725000 0.540000 3.055000 0.555000 ;
      RECT 3.135000 0.710000 4.865000 0.725000 ;
      RECT 3.675000 2.270000 3.865000 2.905000 ;
      RECT 3.675000 2.905000 4.795000 3.075000 ;
      RECT 4.035000 2.100000 4.365000 2.735000 ;
      RECT 4.535000 2.280000 4.795000 2.905000 ;
      RECT 5.200000 1.385000 6.695000 1.585000 ;
      RECT 5.200000 1.585000 5.370000 1.930000 ;
  END
END sky130_fd_sc_lp__o221a_4
