* File: sky130_fd_sc_lp__a21bo_4.spice
* Created: Wed Sep  2 09:18:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21bo_4.pex.spice"
.subckt sky130_fd_sc_lp__a21bo_4  VNB VPB B1_N A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_B1_N_M1013_g N_A_42_47#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.2226 PD=1.46 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75005.4 A=0.126 P=1.98 MULT=1
MM1001 N_X_M1001_d N_A_188_315#_M1001_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2604 PD=1.12 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75001 SB=75004.6
+ A=0.126 P=1.98 MULT=1
MM1011 N_X_M1001_d N_A_188_315#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75004.2 A=0.126 P=1.98 MULT=1
MM1018 N_X_M1018_d N_A_188_315#_M1018_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1218 AS=0.1176 PD=1.13 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.8
+ SB=75003.8 A=0.126 P=1.98 MULT=1
MM1019 N_X_M1018_d N_A_188_315#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1218 AS=0.3171 PD=1.13 PS=1.595 NRD=1.428 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1005 N_A_188_315#_M1005_d N_A_42_47#_M1005_g N_VGND_M1019_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.3171 PD=1.12 PS=1.595 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1020 N_A_188_315#_M1005_d N_A_42_47#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1002 N_A_908_47#_M1002_d N_A2_M1002_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6 SA=75004.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1012 N_A_188_315#_M1012_d N_A1_M1012_g N_A_908_47#_M1002_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1014 N_A_188_315#_M1012_d N_A1_M1014_g N_A_908_47#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1007 N_A_908_47#_M1014_s N_A2_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75005.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_VPWR_M1021_d N_B1_N_M1021_g N_A_42_47#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1021_d N_A_188_315#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A_188_315#_M1003_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1003_d N_A_188_315#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_A_188_315#_M1016_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1004 N_A_188_315#_M1004_d N_A_42_47#_M1004_g N_A_645_367#_M1004_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1017 N_A_188_315#_M1004_d N_A_42_47#_M1017_g N_A_645_367#_M1017_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75002 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_645_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_A_645_367#_M1006_d N_A1_M1006_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=6.2449 M=1 R=8.4
+ SA=75001.5 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1015 N_A_645_367#_M1006_d N_A1_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1015_s N_A2_M1010_g N_A_645_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX22_noxref VNB VPB NWDIODE A=12.3463 P=16.97
*
.include "sky130_fd_sc_lp__a21bo_4.pxi.spice"
*
.ends
*
*
