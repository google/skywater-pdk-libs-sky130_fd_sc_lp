* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 a_454_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND A1 a_819_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_27_47# C1 a_454_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_454_47# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_819_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_1210_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR A1 a_1210_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_819_47# B1 a_454_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Y A2 a_1210_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_1210_367# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_454_47# B1 a_819_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_819_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 VGND A1 a_819_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_819_47# B1 a_454_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VGND A2 a_819_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_819_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_1210_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 a_1210_367# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 Y A2 a_1210_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_819_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 VGND A2 a_819_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 Y D1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 a_454_47# B1 a_819_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 VPWR A1 a_1210_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 a_27_47# D1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 a_27_47# C1 a_454_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
