* File: sky130_fd_sc_lp__a221o_1.pex.spice
* Created: Wed Sep  2 09:21:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221O_1%A_80_21# 1 2 3 12 16 20 21 23 24 26 27 29 33
+ 37 39 42 46
c107 20 0 1.10918e-19 $X=0.6 $Y=1.47
r108 44 45 8.64507 $w=6.43e-07 $l=9e-08 $layer=LI1_cond $X=2.257 $Y=0.925
+ $X2=2.257 $Y2=1.015
r109 42 44 9.36465 $w=6.43e-07 $l=5.05e-07 $layer=LI1_cond $X=2.257 $Y=0.42
+ $X2=2.257 $Y2=0.925
r110 37 48 2.87089 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=3.835 $Y=0.835
+ $X2=3.835 $Y2=0.925
r111 37 39 17.7135 $w=2.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.835 $Y=0.835
+ $X2=3.835 $Y2=0.42
r112 33 35 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=3.805 $Y=1.98
+ $X2=3.805 $Y2=2.91
r113 31 33 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.805 $Y=1.855
+ $X2=3.805 $Y2=1.98
r114 30 44 8.41465 $w=1.8e-07 $l=3.23e-07 $layer=LI1_cond $X=2.58 $Y=0.925
+ $X2=2.257 $Y2=0.925
r115 29 48 4.30634 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=3.7 $Y=0.925
+ $X2=3.835 $Y2=0.925
r116 29 30 69.0101 $w=1.78e-07 $l=1.12e-06 $layer=LI1_cond $X=3.7 $Y=0.925
+ $X2=2.58 $Y2=0.925
r117 28 46 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.205 $Y=1.77
+ $X2=2.115 $Y2=1.77
r118 27 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.64 $Y=1.77
+ $X2=3.805 $Y2=1.855
r119 27 28 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=3.64 $Y=1.77
+ $X2=2.205 $Y2=1.77
r120 26 46 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=1.685
+ $X2=2.115 $Y2=1.77
r121 26 45 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=1.685
+ $X2=2.115 $Y2=1.015
r122 23 46 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.025 $Y=1.77
+ $X2=2.115 $Y2=1.77
r123 23 24 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=2.025 $Y=1.77
+ $X2=0.765 $Y2=1.77
r124 21 51 52.9909 $w=3.65e-07 $l=2.05e-07 $layer=POLY_cond $X=0.582 $Y=1.47
+ $X2=0.582 $Y2=1.675
r125 21 50 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.582 $Y=1.47
+ $X2=0.582 $Y2=1.305
r126 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.47 $X2=0.6 $Y2=1.47
r127 18 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.64 $Y=1.685
+ $X2=0.765 $Y2=1.77
r128 18 20 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=0.64 $Y=1.685
+ $X2=0.64 $Y2=1.47
r129 16 51 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.675
r130 12 50 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=0.475 $Y=0.655
+ $X2=0.475 $Y2=1.305
r131 3 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.665
+ $Y=1.835 $X2=3.805 $Y2=2.91
r132 3 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.665
+ $Y=1.835 $X2=3.805 $Y2=1.98
r133 2 48 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.235 $X2=3.805 $Y2=0.93
r134 2 39 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.235 $X2=3.805 $Y2=0.42
r135 1 42 45.5 $w=1.7e-07 $l=7.46793e-07 $layer=licon1_NDIFF $count=4 $X=1.755
+ $Y=0.235 $X2=2.415 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%A2 3 6 8 9 10 15 17
r38 15 18 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.147 $Y=1.35
+ $X2=1.147 $Y2=1.515
r39 15 17 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.147 $Y=1.35
+ $X2=1.147 $Y2=1.185
r40 10 26 4.55463 $w=3.08e-07 $l=1.1e-07 $layer=LI1_cond $X=1.21 $Y=1.295
+ $X2=1.21 $Y2=1.185
r41 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.35 $X2=1.14 $Y2=1.35
r42 9 26 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=1.24 $Y=0.925
+ $X2=1.24 $Y2=1.185
r43 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.24 $Y=0.555 $X2=1.24
+ $Y2=0.925
r44 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.245 $Y=2.465
+ $X2=1.245 $Y2=1.515
r45 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.245 $Y=0.655
+ $X2=1.245 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%A1 3 6 8 9 10 15 17
r37 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.35
+ $X2=1.77 $Y2=1.515
r38 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.35
+ $X2=1.77 $Y2=1.185
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.35 $X2=1.77 $Y2=1.35
r40 10 16 1.98076 $w=3.18e-07 $l=5.5e-08 $layer=LI1_cond $X=1.695 $Y=1.295
+ $X2=1.695 $Y2=1.35
r41 10 26 4.89143 $w=3.18e-07 $l=1.1e-07 $layer=LI1_cond $X=1.695 $Y=1.295
+ $X2=1.695 $Y2=1.185
r42 9 26 13.0276 $w=2.28e-07 $l=2.6e-07 $layer=LI1_cond $X=1.65 $Y=0.925
+ $X2=1.65 $Y2=1.185
r43 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=0.555 $X2=1.65
+ $Y2=0.925
r44 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.68 $Y=2.465
+ $X2=1.68 $Y2=1.515
r45 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.68 $Y=0.655
+ $X2=1.68 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%B1 3 6 7 10 12 13
r34 10 13 74.8734 $w=4e-07 $l=3.75e-07 $layer=POLY_cond $X=2.505 $Y=1.35
+ $X2=2.505 $Y2=1.725
r35 10 12 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=1.35
+ $X2=2.505 $Y2=1.185
r36 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.35 $X2=2.47 $Y2=1.35
r37 7 11 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.64 $Y=1.35 $X2=2.47
+ $Y2=1.35
r38 6 13 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.63 $Y=2.465
+ $X2=2.63 $Y2=1.725
r39 3 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.63 $Y=0.655
+ $X2=2.63 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%B2 1 3 4 6 8
r34 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.35 $X2=3.11 $Y2=1.35
r35 4 11 38.7084 $w=3.43e-07 $l=1.86145e-07 $layer=POLY_cond $X=3.14 $Y=1.515
+ $X2=3.095 $Y2=1.35
r36 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.14 $Y=1.515 $X2=3.14
+ $Y2=2.465
r37 1 11 38.7084 $w=3.43e-07 $l=2.11069e-07 $layer=POLY_cond $X=2.99 $Y=1.185
+ $X2=3.095 $Y2=1.35
r38 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.99 $Y=1.185 $X2=2.99
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%C1 3 6 8 9 13 15
r24 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.35
+ $X2=3.68 $Y2=1.515
r25 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.35
+ $X2=3.68 $Y2=1.185
r26 8 9 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.31 $X2=4.08
+ $Y2=1.31
r27 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.68
+ $Y=1.35 $X2=3.68 $Y2=1.35
r28 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.59 $Y=2.465
+ $X2=3.59 $Y2=1.515
r29 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.59 $Y=0.655
+ $X2=3.59 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%X 1 2 7 8 9 10 11 12 13 24 45
r16 22 45 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=0.255 $Y=0.905
+ $X2=0.255 $Y2=0.925
r17 13 42 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.215 $Y=2.775
+ $X2=0.215 $Y2=2.91
r18 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=2.405
+ $X2=0.215 $Y2=2.775
r19 11 12 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=0.215 $Y=1.98
+ $X2=0.215 $Y2=2.405
r20 10 11 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.215 $Y=1.665
+ $X2=0.215 $Y2=1.98
r21 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=1.295
+ $X2=0.215 $Y2=1.665
r22 9 47 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.215 $Y=1.295
+ $X2=0.215 $Y2=1.075
r23 8 47 4.66638 $w=3.38e-07 $l=1.18e-07 $layer=LI1_cond $X=0.255 $Y=0.957
+ $X2=0.255 $Y2=1.075
r24 8 45 1.08465 $w=3.38e-07 $l=3.2e-08 $layer=LI1_cond $X=0.255 $Y=0.957
+ $X2=0.255 $Y2=0.925
r25 8 22 1.11855 $w=3.38e-07 $l=3.3e-08 $layer=LI1_cond $X=0.255 $Y=0.872
+ $X2=0.255 $Y2=0.905
r26 7 8 10.7448 $w=3.38e-07 $l=3.17e-07 $layer=LI1_cond $X=0.255 $Y=0.555
+ $X2=0.255 $Y2=0.872
r27 7 24 5.76222 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=0.555
+ $X2=0.255 $Y2=0.385
r28 2 42 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r29 2 11 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
r30 1 24 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r55 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 30 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 27 39 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=0.86 $Y2=3.33
r61 27 29 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 22 39 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.86 $Y2=3.33
r65 22 24 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 20 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 20 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 20 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 18 29 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.73 $Y=3.33 $X2=1.68
+ $Y2=3.33
r70 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=1.895 $Y2=3.33
r71 17 32 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.06 $Y=3.33 $X2=2.16
+ $Y2=3.33
r72 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=3.33
+ $X2=1.895 $Y2=3.33
r73 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=3.245
+ $X2=1.895 $Y2=3.33
r74 13 15 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.895 $Y=3.245
+ $X2=1.895 $Y2=2.48
r75 9 12 14.9956 $w=6.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.86 $Y=2.11 $X2=0.86
+ $Y2=2.95
r76 7 39 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=3.245 $X2=0.86
+ $Y2=3.33
r77 7 12 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.86 $Y=3.245
+ $X2=0.86 $Y2=2.95
r78 2 15 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=1.755
+ $Y=1.835 $X2=1.895 $Y2=2.48
r79 1 12 200 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.95
r80 1 9 200 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=3 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%A_264_367# 1 2 7 9 11 13 15
r23 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=2.195
+ $X2=2.915 $Y2=2.11
r24 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.915 $Y=2.195
+ $X2=2.915 $Y2=2.625
r25 12 18 3.67268 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.56 $Y=2.11
+ $X2=1.462 $Y2=2.11
r26 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=2.11
+ $X2=2.915 $Y2=2.11
r27 11 12 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.75 $Y=2.11
+ $X2=1.56 $Y2=2.11
r28 7 18 3.18549 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.462 $Y=2.195
+ $X2=1.462 $Y2=2.11
r29 7 9 40.6667 $w=1.93e-07 $l=7.15e-07 $layer=LI1_cond $X=1.462 $Y=2.195
+ $X2=1.462 $Y2=2.91
r30 2 20 600 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.835 $X2=2.915 $Y2=2.11
r31 2 15 600 $w=1.7e-07 $l=8.88819e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=1.835 $X2=2.915 $Y2=2.625
r32 1 18 400 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=1.32
+ $Y=1.835 $X2=1.465 $Y2=2.19
r33 1 9 400 $w=1.7e-07 $l=1.14521e-06 $layer=licon1_PDIFF $count=1 $X=1.32
+ $Y=1.835 $X2=1.465 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%A_458_367# 1 2 9 11 12 13 15
r25 13 18 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=2.905
+ $X2=3.36 $Y2=2.99
r26 13 15 37.4544 $w=2.18e-07 $l=7.15e-07 $layer=LI1_cond $X=3.36 $Y=2.905
+ $X2=3.36 $Y2=2.19
r27 11 18 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.25 $Y=2.99 $X2=3.36
+ $Y2=2.99
r28 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.25 $Y=2.99
+ $X2=2.58 $Y2=2.99
r29 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=2.905
+ $X2=2.58 $Y2=2.99
r30 7 9 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.415 $Y=2.905
+ $X2=2.415 $Y2=2.48
r31 2 18 400 $w=1.7e-07 $l=1.14521e-06 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.835 $X2=3.36 $Y2=2.91
r32 2 15 400 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.835 $X2=3.36 $Y2=2.19
r33 1 9 300 $w=1.7e-07 $l=7.04734e-07 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=1.835 $X2=2.415 $Y2=2.48
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r47 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r49 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r50 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r51 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 27 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r53 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r55 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r56 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r57 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r59 20 22 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r60 18 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r61 18 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r62 16 30 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.13 $Y=0 $X2=3.12
+ $Y2=0
r63 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=3.295
+ $Y2=0
r64 15 33 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.46 $Y=0 $X2=4.08
+ $Y2=0
r65 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=0 $X2=3.295
+ $Y2=0
r66 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=0.085
+ $X2=3.295 $Y2=0
r67 11 13 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.295 $Y=0.085
+ $X2=3.295 $Y2=0.525
r68 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r69 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.38
r70 2 13 182 $w=1.7e-07 $l=3.8833e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.295 $Y2=0.525
r71 1 9 91 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.78 $Y2=0.38
.ends

