# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__o32ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o32ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.815000 1.210000 6.155000 1.525000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.210000 4.645000 1.525000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.000000 1.415000 2.835000 1.750000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.425000 1.830000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.425000 1.295000 1.750000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.243200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 0.595000 0.915000 1.075000 ;
        RECT 0.585000 1.075000 3.335000 1.245000 ;
        RECT 0.585000 1.920000 3.335000 2.090000 ;
        RECT 0.585000 2.090000 0.915000 2.735000 ;
        RECT 1.605000 0.595000 1.935000 1.075000 ;
        RECT 3.005000 1.245000 3.335000 1.920000 ;
        RECT 3.005000 2.090000 3.335000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 6.240000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 6.430000 3.520000 ;
        RECT  2.415000 1.645000 4.765000 1.655000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.155000  0.255000 2.445000 0.425000 ;
      RECT 0.155000  0.425000 0.415000 1.185000 ;
      RECT 0.155000  1.920000 0.415000 2.905000 ;
      RECT 0.155000  2.905000 1.275000 3.075000 ;
      RECT 1.085000  2.260000 2.205000 2.450000 ;
      RECT 1.085000  2.450000 1.275000 2.905000 ;
      RECT 1.095000  0.425000 1.425000 0.905000 ;
      RECT 1.445000  2.620000 1.775000 3.245000 ;
      RECT 1.945000  2.450000 2.205000 3.075000 ;
      RECT 2.115000  0.425000 2.445000 0.735000 ;
      RECT 2.115000  0.735000 3.775000 0.870000 ;
      RECT 2.115000  0.870000 5.595000 0.905000 ;
      RECT 2.555000  2.260000 2.825000 2.905000 ;
      RECT 2.555000  2.905000 4.625000 3.075000 ;
      RECT 2.615000  0.085000 3.405000 0.565000 ;
      RECT 3.505000  0.905000 5.595000 1.040000 ;
      RECT 3.505000  1.815000 3.695000 2.905000 ;
      RECT 3.575000  0.315000 3.775000 0.735000 ;
      RECT 3.865000  1.705000 5.540000 1.875000 ;
      RECT 3.865000  1.875000 4.195000 2.735000 ;
      RECT 3.945000  0.085000 4.275000 0.700000 ;
      RECT 4.365000  2.045000 4.625000 2.905000 ;
      RECT 4.465000  0.315000 4.665000 0.870000 ;
      RECT 4.815000  2.045000 5.145000 3.245000 ;
      RECT 4.835000  0.085000 5.165000 0.700000 ;
      RECT 5.315000  1.875000 5.540000 3.075000 ;
      RECT 5.335000  0.315000 5.595000 0.870000 ;
      RECT 5.710000  1.815000 6.005000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__o32ai_2
END LIBRARY
