* File: sky130_fd_sc_lp__conb_1.spice
* Created: Fri Aug 28 10:19:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__conb_1.pex.spice"
.subckt sky130_fd_sc_lp__conb_1  VNB VPB HI LO VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* LO	LO
* HI	HI
* VPB	VPB
* VNB	VNB
MM1001 N_LO_M1001_d N_HI_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_LO_M1003_g N_LO_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_HI_M1002_d N_HI_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_LO_M1000_g N_HI_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__conb_1.pxi.spice"
*
.ends
*
*
