* NGSPICE file created from sky130_fd_sc_lp__a41o_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_550_47# A2 a_478_47# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=1.764e+11p ps=2.1e+06u
M1001 VGND a_113_237# X VNB nshort w=840000u l=150000u
+  ad=8.736e+11p pd=5.44e+06u as=2.226e+11p ps=2.21e+06u
M1002 a_478_47# A1 a_113_237# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=2.8e+06u
M1003 a_346_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0395e+12p pd=9.21e+06u as=1.5183e+12p ps=9.97e+06u
M1004 a_658_47# A3 a_550_47# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=0p ps=0u
M1005 VPWR A1 a_346_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_346_367# A4 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A4 a_658_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_113_237# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1009 VPWR A3 a_346_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_113_237# B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_346_367# B1 a_113_237# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

