* File: sky130_fd_sc_lp__invkapwr_8.pxi.spice
* Created: Fri Aug 28 10:39:23 2020
* 
x_PM_SKY130_FD_SC_LP__INVKAPWR_8%A N_A_M1000_g N_A_M1003_g N_A_M1001_g
+ N_A_M1005_g N_A_M1002_g N_A_M1007_g N_A_M1004_g N_A_M1008_g N_A_M1006_g
+ N_A_M1010_g N_A_M1009_g N_A_M1012_g N_A_M1011_g N_A_M1014_g N_A_M1013_g
+ N_A_M1015_g N_A_M1018_g N_A_M1016_g N_A_M1017_g N_A_M1019_g A A A A A A A A A
+ A N_A_c_109_n PM_SKY130_FD_SC_LP__INVKAPWR_8%A
x_PM_SKY130_FD_SC_LP__INVKAPWR_8%KAPWR N_KAPWR_M1000_s N_KAPWR_M1003_s
+ N_KAPWR_M1007_s N_KAPWR_M1010_s N_KAPWR_M1014_s N_KAPWR_M1016_s
+ N_KAPWR_M1019_s KAPWR N_KAPWR_c_268_n N_KAPWR_c_293_p N_KAPWR_c_298_p
+ N_KAPWR_c_303_p N_KAPWR_c_308_p N_KAPWR_c_313_p N_KAPWR_c_318_p
+ N_KAPWR_c_269_n PM_SKY130_FD_SC_LP__INVKAPWR_8%KAPWR
x_PM_SKY130_FD_SC_LP__INVKAPWR_8%Y N_Y_M1001_s N_Y_M1004_s N_Y_M1009_s
+ N_Y_M1013_s N_Y_M1000_d N_Y_M1005_d N_Y_M1008_d N_Y_M1012_d N_Y_M1015_d
+ N_Y_M1017_d N_Y_c_345_n N_Y_c_346_n N_Y_c_347_n N_Y_c_363_n N_Y_c_364_n
+ N_Y_c_385_n N_Y_c_365_n N_Y_c_348_n N_Y_c_393_n N_Y_c_349_n N_Y_c_366_n
+ N_Y_c_350_n N_Y_c_405_n N_Y_c_351_n N_Y_c_367_n N_Y_c_352_n N_Y_c_417_n
+ N_Y_c_353_n N_Y_c_368_n N_Y_c_354_n N_Y_c_429_n N_Y_c_369_n N_Y_c_435_n
+ N_Y_c_370_n N_Y_c_371_n N_Y_c_355_n N_Y_c_372_n N_Y_c_356_n N_Y_c_373_n
+ N_Y_c_357_n N_Y_c_374_n N_Y_c_358_n N_Y_c_375_n N_Y_c_376_n Y Y N_Y_c_361_n
+ PM_SKY130_FD_SC_LP__INVKAPWR_8%Y
x_PM_SKY130_FD_SC_LP__INVKAPWR_8%VGND N_VGND_M1001_d N_VGND_M1002_d
+ N_VGND_M1006_d N_VGND_M1011_d N_VGND_M1018_d N_VGND_c_542_n N_VGND_c_543_n
+ N_VGND_c_544_n N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n N_VGND_c_548_n
+ N_VGND_c_549_n N_VGND_c_550_n N_VGND_c_551_n N_VGND_c_552_n N_VGND_c_553_n
+ VGND N_VGND_c_554_n N_VGND_c_555_n N_VGND_c_556_n N_VGND_c_557_n
+ N_VGND_c_558_n PM_SKY130_FD_SC_LP__INVKAPWR_8%VGND
x_PM_SKY130_FD_SC_LP__INVKAPWR_8%VPWR VPWR N_VPWR_c_605_n VPWR
+ PM_SKY130_FD_SC_LP__INVKAPWR_8%VPWR
cc_1 VNB N_A_M1000_g 0.00628988f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_2 VNB N_A_M1003_g 0.00579465f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_3 VNB N_A_M1001_g 0.0432088f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=0.56
cc_4 VNB N_A_M1005_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_5 VNB N_A_M1002_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.56
cc_6 VNB N_A_M1007_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_7 VNB N_A_M1004_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=0.56
cc_8 VNB N_A_M1008_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=2.465
cc_9 VNB N_A_M1006_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=0.56
cc_10 VNB N_A_M1010_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=2.465
cc_11 VNB N_A_M1009_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=0.56
cc_12 VNB N_A_M1012_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=2.465
cc_13 VNB N_A_M1011_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=0.56
cc_14 VNB N_A_M1014_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=2.465
cc_15 VNB N_A_M1013_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=0.56
cc_16 VNB N_A_M1015_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=2.465
cc_17 VNB N_A_M1018_g 0.0432088f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=0.56
cc_18 VNB N_A_M1016_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=2.465
cc_19 VNB N_A_M1017_g 0.00579365f $X=-0.19 $Y=-0.245 $X2=4.845 $Y2=2.465
cc_20 VNB N_A_M1019_g 0.00625137f $X=-0.19 $Y=-0.245 $X2=5.275 $Y2=2.465
cc_21 VNB N_A_c_109_n 0.275358f $X=-0.19 $Y=-0.245 $X2=5.275 $Y2=1.375
cc_22 VNB N_Y_c_345_n 0.0333088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_346_n 0.0278014f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=1.21
cc_24 VNB N_Y_c_347_n 0.0128703f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=0.56
cc_25 VNB N_Y_c_348_n 0.00119645f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=2.465
cc_26 VNB N_Y_c_349_n 0.00538522f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=2.465
cc_27 VNB N_Y_c_350_n 0.00110053f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.54
cc_28 VNB N_Y_c_351_n 0.00538522f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=1.54
cc_29 VNB N_Y_c_352_n 0.00110053f $X=-0.19 $Y=-0.245 $X2=4.845 $Y2=2.465
cc_30 VNB N_Y_c_353_n 0.00538522f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_31 VNB N_Y_c_354_n 0.00119645f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.21
cc_32 VNB N_Y_c_355_n 0.00205825f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=1.375
cc_33 VNB N_Y_c_356_n 0.00205825f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=1.375
cc_34 VNB N_Y_c_357_n 0.00205825f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.375
cc_35 VNB N_Y_c_358_n 0.00205825f $X=-0.19 $Y=-0.245 $X2=4.845 $Y2=1.375
cc_36 VNB Y 0.0263263f $X=-0.19 $Y=-0.245 $X2=5.275 $Y2=1.375
cc_37 VNB Y 0.0337179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_361_n 0.0132875f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.375
cc_39 VNB N_VGND_c_542_n 0.0235135f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.56
cc_40 VNB N_VGND_c_543_n 0.00698312f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_41 VNB N_VGND_c_544_n 0.00698312f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=0.56
cc_42 VNB N_VGND_c_545_n 0.00698312f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=2.465
cc_43 VNB N_VGND_c_546_n 0.0171844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_547_n 0.0235135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_548_n 0.0171844f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=2.465
cc_46 VNB N_VGND_c_549_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_550_n 0.0171844f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=0.56
cc_48 VNB N_VGND_c_551_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=0.56
cc_49 VNB N_VGND_c_552_n 0.0171844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_553_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=1.54
cc_51 VNB N_VGND_c_554_n 0.0347608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_555_n 0.0328515f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=1.21
cc_53 VNB N_VGND_c_556_n 0.326397f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=0.56
cc_54 VNB N_VGND_c_557_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=1.54
cc_55 VNB N_VGND_c_558_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB VPWR 0.243291f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.54
cc_57 VPB N_A_M1000_g 0.0234928f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_58 VPB N_A_M1003_g 0.018718f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_59 VPB N_A_M1005_g 0.0187369f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.465
cc_60 VPB N_A_M1007_g 0.0187369f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_61 VPB N_A_M1008_g 0.0187369f $X=-0.19 $Y=1.655 $X2=2.265 $Y2=2.465
cc_62 VPB N_A_M1010_g 0.0187369f $X=-0.19 $Y=1.655 $X2=2.695 $Y2=2.465
cc_63 VPB N_A_M1012_g 0.0187369f $X=-0.19 $Y=1.655 $X2=3.125 $Y2=2.465
cc_64 VPB N_A_M1014_g 0.0187369f $X=-0.19 $Y=1.655 $X2=3.555 $Y2=2.465
cc_65 VPB N_A_M1015_g 0.0187369f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=2.465
cc_66 VPB N_A_M1016_g 0.0187369f $X=-0.19 $Y=1.655 $X2=4.415 $Y2=2.465
cc_67 VPB N_A_M1017_g 0.0187175f $X=-0.19 $Y=1.655 $X2=4.845 $Y2=2.465
cc_68 VPB N_A_M1019_g 0.0234742f $X=-0.19 $Y=1.655 $X2=5.275 $Y2=2.465
cc_69 VPB N_KAPWR_c_268_n 0.0311165f $X=-0.19 $Y=1.655 $X2=2.265 $Y2=1.21
cc_70 VPB N_KAPWR_c_269_n 0.0294445f $X=-0.19 $Y=1.655 $X2=5.275 $Y2=1.54
cc_71 VPB N_Y_c_345_n 0.0025871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_Y_c_363_n 0.00201395f $X=-0.19 $Y=1.655 $X2=2.695 $Y2=0.56
cc_73 VPB N_Y_c_364_n 0.00873266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_Y_c_365_n 0.00243013f $X=-0.19 $Y=1.655 $X2=3.125 $Y2=0.56
cc_75 VPB N_Y_c_366_n 0.00243013f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=1.21
cc_76 VPB N_Y_c_367_n 0.00243013f $X=-0.19 $Y=1.655 $X2=4.415 $Y2=2.465
cc_77 VPB N_Y_c_368_n 0.00243013f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.21
cc_78 VPB N_Y_c_369_n 0.00242094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_Y_c_370_n 0.0089125f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.375
cc_80 VPB N_Y_c_371_n 0.00206951f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=1.375
cc_81 VPB N_Y_c_372_n 0.00206951f $X=-0.19 $Y=1.655 $X2=2.265 $Y2=1.375
cc_82 VPB N_Y_c_373_n 0.00206951f $X=-0.19 $Y=1.655 $X2=3.125 $Y2=1.375
cc_83 VPB N_Y_c_374_n 0.00206951f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=1.375
cc_84 VPB N_Y_c_375_n 0.00206951f $X=-0.19 $Y=1.655 $X2=5.1 $Y2=1.375
cc_85 VPB N_Y_c_376_n 0.00211646f $X=-0.19 $Y=1.655 $X2=5.1 $Y2=1.375
cc_86 VPB Y 0.00255258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB VPWR 0.0441237f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.54
cc_88 VPB N_VPWR_c_605_n 0.15719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 N_A_M1000_g N_KAPWR_c_269_n 0.00731133f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A_M1003_g N_KAPWR_c_269_n 0.00731133f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_91 N_A_M1005_g N_KAPWR_c_269_n 0.00731133f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A_M1007_g N_KAPWR_c_269_n 0.00731133f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_93 N_A_M1008_g N_KAPWR_c_269_n 0.00731133f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_M1010_g N_KAPWR_c_269_n 0.00731133f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A_M1012_g N_KAPWR_c_269_n 0.00731133f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A_M1014_g N_KAPWR_c_269_n 0.00731133f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A_M1015_g N_KAPWR_c_269_n 0.00731133f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_M1016_g N_KAPWR_c_269_n 0.00731133f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_M1017_g N_KAPWR_c_269_n 0.00731133f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_M1019_g N_KAPWR_c_269_n 0.00731133f $X=5.275 $Y=2.465 $X2=0 $Y2=0
cc_101 A N_Y_c_345_n 0.0262109f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_102 N_A_c_109_n N_Y_c_345_n 0.0152693f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_103 N_A_M1001_g N_Y_c_346_n 0.0155371f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_104 A N_Y_c_346_n 0.073583f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A_c_109_n N_Y_c_346_n 0.0221841f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_106 N_A_M1000_g N_Y_c_363_n 0.0165938f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_107 A N_Y_c_363_n 0.00860651f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_108 N_A_M1000_g N_Y_c_385_n 8.21354e-19 $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_M1003_g N_Y_c_385_n 8.21794e-19 $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A_M1003_g N_Y_c_365_n 0.0146426f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_M1005_g N_Y_c_365_n 0.0146426f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_112 A N_Y_c_365_n 0.0443704f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_113 N_A_c_109_n N_Y_c_365_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_114 N_A_M1001_g N_Y_c_348_n 0.00194229f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_115 N_A_M1002_g N_Y_c_348_n 0.00105846f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A_M1005_g N_Y_c_393_n 8.21354e-19 $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_M1007_g N_Y_c_393_n 8.21794e-19 $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_M1002_g N_Y_c_349_n 0.0131322f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_119 N_A_M1004_g N_Y_c_349_n 0.0131322f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_120 A N_Y_c_349_n 0.0444367f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_121 N_A_c_109_n N_Y_c_349_n 0.00225043f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_122 N_A_M1007_g N_Y_c_366_n 0.0146426f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_M1008_g N_Y_c_366_n 0.0146426f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_124 A N_Y_c_366_n 0.0443704f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A_c_109_n N_Y_c_366_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_126 N_A_M1004_g N_Y_c_350_n 0.00105846f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_127 N_A_M1006_g N_Y_c_350_n 0.00105846f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_128 N_A_M1008_g N_Y_c_405_n 8.21354e-19 $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A_M1010_g N_Y_c_405_n 8.21794e-19 $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A_M1006_g N_Y_c_351_n 0.0131322f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_131 N_A_M1009_g N_Y_c_351_n 0.0131322f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_132 A N_Y_c_351_n 0.0444367f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_133 N_A_c_109_n N_Y_c_351_n 0.00225043f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_134 N_A_M1010_g N_Y_c_367_n 0.0146426f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_M1012_g N_Y_c_367_n 0.0146426f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_136 A N_Y_c_367_n 0.0443704f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_137 N_A_c_109_n N_Y_c_367_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_138 N_A_M1009_g N_Y_c_352_n 0.00105846f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_139 N_A_M1011_g N_Y_c_352_n 0.00105846f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A_M1012_g N_Y_c_417_n 8.21354e-19 $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_M1014_g N_Y_c_417_n 8.21794e-19 $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_M1011_g N_Y_c_353_n 0.0131322f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_143 N_A_M1013_g N_Y_c_353_n 0.0131322f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_144 A N_Y_c_353_n 0.0444367f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_145 N_A_c_109_n N_Y_c_353_n 0.00225043f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_146 N_A_M1014_g N_Y_c_368_n 0.0146426f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_M1015_g N_Y_c_368_n 0.0146426f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_148 A N_Y_c_368_n 0.0443704f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A_c_109_n N_Y_c_368_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_150 N_A_M1013_g N_Y_c_354_n 0.00105846f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A_M1018_g N_Y_c_354_n 0.00194229f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A_M1015_g N_Y_c_429_n 8.21354e-19 $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_M1016_g N_Y_c_429_n 8.21794e-19 $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_M1016_g N_Y_c_369_n 0.0146426f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_M1017_g N_Y_c_369_n 0.0146085f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_156 A N_Y_c_369_n 0.0439938f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A_c_109_n N_Y_c_369_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_158 N_A_M1017_g N_Y_c_435_n 8.22659e-19 $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A_M1019_g N_Y_c_435_n 8.22659e-19 $X=5.275 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A_M1019_g N_Y_c_370_n 0.0170121f $X=5.275 $Y=2.465 $X2=0 $Y2=0
cc_161 A N_Y_c_370_n 0.00536724f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_162 A N_Y_c_371_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A_c_109_n N_Y_c_371_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_164 A N_Y_c_355_n 0.0218346f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A_c_109_n N_Y_c_355_n 0.00232201f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_166 A N_Y_c_372_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_167 N_A_c_109_n N_Y_c_372_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_168 A N_Y_c_356_n 0.0218346f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_169 N_A_c_109_n N_Y_c_356_n 0.00232201f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_170 A N_Y_c_373_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A_c_109_n N_Y_c_373_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_172 A N_Y_c_357_n 0.0218346f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A_c_109_n N_Y_c_357_n 0.00232201f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_174 A N_Y_c_374_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A_c_109_n N_Y_c_374_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_176 A N_Y_c_358_n 0.0218346f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A_c_109_n N_Y_c_358_n 0.00232201f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_178 A N_Y_c_375_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A_c_109_n N_Y_c_375_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_180 A N_Y_c_376_n 0.0219298f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_181 N_A_c_109_n N_Y_c_376_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_182 N_A_M1018_g Y 0.0155371f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_183 A Y 0.0705391f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A_c_109_n Y 0.0223886f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_185 A Y 0.0263702f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A_c_109_n Y 0.0160643f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_187 N_A_M1001_g N_VGND_c_542_n 0.0038152f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A_M1002_g N_VGND_c_543_n 0.00181038f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A_M1004_g N_VGND_c_543_n 0.00181038f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_190 N_A_M1006_g N_VGND_c_544_n 0.00181038f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A_M1009_g N_VGND_c_544_n 0.00181038f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A_M1011_g N_VGND_c_545_n 0.00181038f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_193 N_A_M1013_g N_VGND_c_545_n 0.00181038f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_194 N_A_M1013_g N_VGND_c_546_n 0.00478016f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_195 N_A_M1018_g N_VGND_c_546_n 0.00478016f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_196 N_A_M1018_g N_VGND_c_547_n 0.0038152f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A_M1001_g N_VGND_c_548_n 0.00478016f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A_M1002_g N_VGND_c_548_n 0.00478016f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_199 N_A_M1004_g N_VGND_c_550_n 0.00478016f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_200 N_A_M1006_g N_VGND_c_550_n 0.00478016f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_201 N_A_M1009_g N_VGND_c_552_n 0.00478016f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_202 N_A_M1011_g N_VGND_c_552_n 0.00478016f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A_M1001_g N_VGND_c_556_n 0.0051579f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_204 N_A_M1002_g N_VGND_c_556_n 0.00490796f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_205 N_A_M1004_g N_VGND_c_556_n 0.00490796f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_206 N_A_M1006_g N_VGND_c_556_n 0.00490796f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A_M1009_g N_VGND_c_556_n 0.00490796f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_208 N_A_M1011_g N_VGND_c_556_n 0.00490796f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_209 N_A_M1013_g N_VGND_c_556_n 0.00490796f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_210 N_A_M1018_g N_VGND_c_556_n 0.0051579f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_211 N_A_M1000_g VPWR 0.00631531f $X=0.545 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_212 N_A_M1003_g VPWR 0.0053229f $X=0.975 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_213 N_A_M1005_g VPWR 0.0053229f $X=1.405 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_214 N_A_M1007_g VPWR 0.0053229f $X=1.835 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_215 N_A_M1008_g VPWR 0.0053229f $X=2.265 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_216 N_A_M1010_g VPWR 0.0053229f $X=2.695 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_217 N_A_M1012_g VPWR 0.0053229f $X=3.125 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_218 N_A_M1014_g VPWR 0.0053229f $X=3.555 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_219 N_A_M1015_g VPWR 0.0053229f $X=3.985 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_220 N_A_M1016_g VPWR 0.0053229f $X=4.415 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_221 N_A_M1017_g VPWR 0.0053229f $X=4.845 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_222 N_A_M1019_g VPWR 0.00626484f $X=5.275 $Y=2.465 $X2=-0.19 $Y2=-0.245
cc_223 N_A_M1000_g N_VPWR_c_605_n 0.00585385f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_M1003_g N_VPWR_c_605_n 0.00585385f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A_M1005_g N_VPWR_c_605_n 0.00585385f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A_M1007_g N_VPWR_c_605_n 0.00585385f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_227 N_A_M1008_g N_VPWR_c_605_n 0.00585385f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A_M1010_g N_VPWR_c_605_n 0.00585385f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A_M1012_g N_VPWR_c_605_n 0.00585385f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A_M1014_g N_VPWR_c_605_n 0.00585385f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_M1015_g N_VPWR_c_605_n 0.00585385f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A_M1016_g N_VPWR_c_605_n 0.00585385f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A_M1017_g N_VPWR_c_605_n 0.00585385f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A_M1019_g N_VPWR_c_605_n 0.00585385f $X=5.275 $Y=2.465 $X2=0 $Y2=0
cc_235 N_KAPWR_c_269_n N_Y_M1000_d 9.4832e-19 $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_236 N_KAPWR_c_269_n N_Y_M1005_d 9.4832e-19 $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_237 N_KAPWR_c_269_n N_Y_M1008_d 9.4832e-19 $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_238 N_KAPWR_c_269_n N_Y_M1012_d 9.4832e-19 $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_239 N_KAPWR_c_269_n N_Y_M1015_d 9.4832e-19 $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_240 N_KAPWR_c_269_n N_Y_M1017_d 7.22529e-19 $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_241 N_KAPWR_M1000_s N_Y_c_363_n 7.1286e-19 $X=0.205 $Y=1.835 $X2=0 $Y2=0
cc_242 N_KAPWR_c_268_n N_Y_c_363_n 0.00550656f $X=0.33 $Y=2.22 $X2=0 $Y2=0
cc_243 N_KAPWR_M1000_s N_Y_c_364_n 0.00178451f $X=0.205 $Y=1.835 $X2=0 $Y2=0
cc_244 N_KAPWR_c_268_n N_Y_c_364_n 0.0129974f $X=0.33 $Y=2.22 $X2=0 $Y2=0
cc_245 N_KAPWR_c_268_n N_Y_c_385_n 0.00885226f $X=0.33 $Y=2.22 $X2=0 $Y2=0
cc_246 N_KAPWR_c_293_p N_Y_c_385_n 0.0091127f $X=1.19 $Y=2.22 $X2=0 $Y2=0
cc_247 N_KAPWR_c_269_n N_Y_c_385_n 0.0284615f $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_248 N_KAPWR_M1003_s N_Y_c_365_n 0.00176619f $X=1.05 $Y=1.835 $X2=0 $Y2=0
cc_249 N_KAPWR_c_293_p N_Y_c_365_n 0.0135319f $X=1.19 $Y=2.22 $X2=0 $Y2=0
cc_250 N_KAPWR_c_293_p N_Y_c_393_n 0.00885226f $X=1.19 $Y=2.22 $X2=0 $Y2=0
cc_251 N_KAPWR_c_298_p N_Y_c_393_n 0.0091127f $X=2.05 $Y=2.22 $X2=0 $Y2=0
cc_252 N_KAPWR_c_269_n N_Y_c_393_n 0.0284615f $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_253 N_KAPWR_M1007_s N_Y_c_366_n 0.00176619f $X=1.91 $Y=1.835 $X2=0 $Y2=0
cc_254 N_KAPWR_c_298_p N_Y_c_366_n 0.0135319f $X=2.05 $Y=2.22 $X2=0 $Y2=0
cc_255 N_KAPWR_c_298_p N_Y_c_405_n 0.00885226f $X=2.05 $Y=2.22 $X2=0 $Y2=0
cc_256 N_KAPWR_c_303_p N_Y_c_405_n 0.0091127f $X=2.91 $Y=2.22 $X2=0 $Y2=0
cc_257 N_KAPWR_c_269_n N_Y_c_405_n 0.0284615f $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_258 N_KAPWR_M1010_s N_Y_c_367_n 0.00176619f $X=2.77 $Y=1.835 $X2=0 $Y2=0
cc_259 N_KAPWR_c_303_p N_Y_c_367_n 0.0135319f $X=2.91 $Y=2.22 $X2=0 $Y2=0
cc_260 N_KAPWR_c_303_p N_Y_c_417_n 0.00885226f $X=2.91 $Y=2.22 $X2=0 $Y2=0
cc_261 N_KAPWR_c_308_p N_Y_c_417_n 0.0091127f $X=3.77 $Y=2.22 $X2=0 $Y2=0
cc_262 N_KAPWR_c_269_n N_Y_c_417_n 0.0284615f $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_263 N_KAPWR_M1014_s N_Y_c_368_n 0.00176619f $X=3.63 $Y=1.835 $X2=0 $Y2=0
cc_264 N_KAPWR_c_308_p N_Y_c_368_n 0.0135319f $X=3.77 $Y=2.22 $X2=0 $Y2=0
cc_265 N_KAPWR_c_308_p N_Y_c_429_n 0.00885226f $X=3.77 $Y=2.22 $X2=0 $Y2=0
cc_266 N_KAPWR_c_313_p N_Y_c_429_n 0.0091127f $X=4.63 $Y=2.22 $X2=0 $Y2=0
cc_267 N_KAPWR_c_269_n N_Y_c_429_n 0.0284615f $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_268 N_KAPWR_M1016_s N_Y_c_369_n 0.00176619f $X=4.49 $Y=1.835 $X2=0 $Y2=0
cc_269 N_KAPWR_c_313_p N_Y_c_369_n 0.0135319f $X=4.63 $Y=2.22 $X2=0 $Y2=0
cc_270 N_KAPWR_c_313_p N_Y_c_435_n 0.00911549f $X=4.63 $Y=2.22 $X2=0 $Y2=0
cc_271 N_KAPWR_c_318_p N_Y_c_435_n 0.0091127f $X=5.49 $Y=2.22 $X2=0 $Y2=0
cc_272 N_KAPWR_c_269_n N_Y_c_435_n 0.0288605f $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_273 N_KAPWR_M1019_s N_Y_c_370_n 0.00250337f $X=5.35 $Y=1.835 $X2=0 $Y2=0
cc_274 N_KAPWR_c_318_p N_Y_c_370_n 0.0183848f $X=5.49 $Y=2.22 $X2=0 $Y2=0
cc_275 N_KAPWR_M1000_s VPWR 0.00114602f $X=0.205 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_276 N_KAPWR_M1003_s VPWR 0.00121489f $X=1.05 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_277 N_KAPWR_M1007_s VPWR 0.00121489f $X=1.91 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_278 N_KAPWR_M1010_s VPWR 0.00121489f $X=2.77 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_279 N_KAPWR_M1014_s VPWR 0.00121489f $X=3.63 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_280 N_KAPWR_M1016_s VPWR 0.00121489f $X=4.49 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_281 N_KAPWR_M1019_s VPWR 0.00114194f $X=5.35 $Y=1.835 $X2=-0.19 $Y2=1.655
cc_282 N_KAPWR_c_268_n VPWR 0.00242444f $X=0.33 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_283 N_KAPWR_c_293_p VPWR 0.00242444f $X=1.19 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_284 N_KAPWR_c_298_p VPWR 0.00242444f $X=2.05 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_285 N_KAPWR_c_303_p VPWR 0.00242444f $X=2.91 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_286 N_KAPWR_c_308_p VPWR 0.00242444f $X=3.77 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_287 N_KAPWR_c_313_p VPWR 0.00242444f $X=4.63 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_288 N_KAPWR_c_318_p VPWR 0.00237745f $X=5.49 $Y=2.22 $X2=-0.19 $Y2=1.655
cc_289 N_KAPWR_c_269_n VPWR 0.581884f $X=5.495 $Y=2.81 $X2=-0.19 $Y2=1.655
cc_290 N_KAPWR_c_268_n N_VPWR_c_605_n 0.0165439f $X=0.33 $Y=2.22 $X2=0 $Y2=0
cc_291 N_KAPWR_c_293_p N_VPWR_c_605_n 0.0149362f $X=1.19 $Y=2.22 $X2=0 $Y2=0
cc_292 N_KAPWR_c_298_p N_VPWR_c_605_n 0.0149362f $X=2.05 $Y=2.22 $X2=0 $Y2=0
cc_293 N_KAPWR_c_303_p N_VPWR_c_605_n 0.0149362f $X=2.91 $Y=2.22 $X2=0 $Y2=0
cc_294 N_KAPWR_c_308_p N_VPWR_c_605_n 0.0149362f $X=3.77 $Y=2.22 $X2=0 $Y2=0
cc_295 N_KAPWR_c_313_p N_VPWR_c_605_n 0.0149362f $X=4.63 $Y=2.22 $X2=0 $Y2=0
cc_296 N_KAPWR_c_318_p N_VPWR_c_605_n 0.0161868f $X=5.49 $Y=2.22 $X2=0 $Y2=0
cc_297 N_KAPWR_c_269_n N_VPWR_c_605_n 0.0137776f $X=5.495 $Y=2.81 $X2=0 $Y2=0
cc_298 N_Y_c_346_n N_VGND_c_542_n 0.0219547f $X=1.49 $Y=0.94 $X2=0 $Y2=0
cc_299 N_Y_c_349_n N_VGND_c_543_n 0.0169602f $X=2.35 $Y=0.94 $X2=0 $Y2=0
cc_300 N_Y_c_351_n N_VGND_c_544_n 0.0169602f $X=3.21 $Y=0.94 $X2=0 $Y2=0
cc_301 N_Y_c_353_n N_VGND_c_545_n 0.0169602f $X=4.07 $Y=0.94 $X2=0 $Y2=0
cc_302 N_Y_c_354_n N_VGND_c_546_n 0.00786011f $X=4.2 $Y=0.56 $X2=0 $Y2=0
cc_303 Y N_VGND_c_547_n 0.0219547f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_304 N_Y_c_348_n N_VGND_c_548_n 0.00786011f $X=1.62 $Y=0.56 $X2=0 $Y2=0
cc_305 N_Y_c_350_n N_VGND_c_550_n 0.00786011f $X=2.48 $Y=0.56 $X2=0 $Y2=0
cc_306 N_Y_c_352_n N_VGND_c_552_n 0.00786011f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_307 N_Y_c_346_n N_VGND_c_556_n 0.0297069f $X=1.49 $Y=0.94 $X2=0 $Y2=0
cc_308 N_Y_c_347_n N_VGND_c_556_n 0.00670311f $X=0.345 $Y=0.94 $X2=0 $Y2=0
cc_309 N_Y_c_348_n N_VGND_c_556_n 0.00924776f $X=1.62 $Y=0.56 $X2=0 $Y2=0
cc_310 N_Y_c_349_n N_VGND_c_556_n 0.0106287f $X=2.35 $Y=0.94 $X2=0 $Y2=0
cc_311 N_Y_c_350_n N_VGND_c_556_n 0.00924776f $X=2.48 $Y=0.56 $X2=0 $Y2=0
cc_312 N_Y_c_351_n N_VGND_c_556_n 0.0106287f $X=3.21 $Y=0.94 $X2=0 $Y2=0
cc_313 N_Y_c_352_n N_VGND_c_556_n 0.00924776f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_314 N_Y_c_353_n N_VGND_c_556_n 0.0106287f $X=4.07 $Y=0.94 $X2=0 $Y2=0
cc_315 N_Y_c_354_n N_VGND_c_556_n 0.00924776f $X=4.2 $Y=0.56 $X2=0 $Y2=0
cc_316 Y N_VGND_c_556_n 0.0283045f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_317 N_Y_c_361_n N_VGND_c_556_n 0.00729456f $X=5.527 $Y=1.04 $X2=0 $Y2=0
cc_318 N_Y_M1000_d VPWR 0.00125588f $X=0.62 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_319 N_Y_M1005_d VPWR 0.00125588f $X=1.48 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_320 N_Y_M1008_d VPWR 0.00125588f $X=2.34 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_321 N_Y_M1012_d VPWR 0.00125588f $X=3.2 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_322 N_Y_M1015_d VPWR 0.00125588f $X=4.06 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_323 N_Y_M1017_d VPWR 0.0012358f $X=4.92 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_324 N_Y_c_385_n VPWR 0.0024325f $X=0.76 $Y=2 $X2=-0.19 $Y2=-0.245
cc_325 N_Y_c_393_n VPWR 0.0024325f $X=1.62 $Y=2 $X2=-0.19 $Y2=-0.245
cc_326 N_Y_c_405_n VPWR 0.0024325f $X=2.48 $Y=2 $X2=-0.19 $Y2=-0.245
cc_327 N_Y_c_417_n VPWR 0.0024325f $X=3.34 $Y=2 $X2=-0.19 $Y2=-0.245
cc_328 N_Y_c_429_n VPWR 0.0024325f $X=4.2 $Y=2 $X2=-0.19 $Y2=-0.245
cc_329 N_Y_c_435_n VPWR 0.00248057f $X=5.06 $Y=2 $X2=-0.19 $Y2=-0.245
cc_330 N_Y_c_385_n N_VPWR_c_605_n 0.0124051f $X=0.76 $Y=2 $X2=0 $Y2=0
cc_331 N_Y_c_393_n N_VPWR_c_605_n 0.0124051f $X=1.62 $Y=2 $X2=0 $Y2=0
cc_332 N_Y_c_405_n N_VPWR_c_605_n 0.0124051f $X=2.48 $Y=2 $X2=0 $Y2=0
cc_333 N_Y_c_417_n N_VPWR_c_605_n 0.0124051f $X=3.34 $Y=2 $X2=0 $Y2=0
cc_334 N_Y_c_429_n N_VPWR_c_605_n 0.0124051f $X=4.2 $Y=2 $X2=0 $Y2=0
cc_335 N_Y_c_435_n N_VPWR_c_605_n 0.012556f $X=5.06 $Y=2 $X2=0 $Y2=0
