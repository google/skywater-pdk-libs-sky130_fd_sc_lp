* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__maj3_4 A B C VGND VNB VPB VPWR X
X0 a_65_367# C a_154_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR A a_318_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_65_367# C a_154_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_318_47# B a_65_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_65_367# B a_482_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR a_65_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 X a_65_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_482_367# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND A a_318_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_154_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 X a_65_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND a_65_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_318_367# B a_65_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VGND a_65_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VPWR a_65_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_154_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_482_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_65_367# B a_482_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 X a_65_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 X a_65_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
