* File: sky130_fd_sc_lp__a311o_4.pxi.spice
* Created: Wed Sep  2 09:25:14 2020
* 
x_PM_SKY130_FD_SC_LP__A311O_4%C1 N_C1_M1002_g N_C1_M1013_g N_C1_M1010_g
+ N_C1_M1026_g C1 C1 N_C1_c_138_n PM_SKY130_FD_SC_LP__A311O_4%C1
x_PM_SKY130_FD_SC_LP__A311O_4%B1 N_B1_M1024_g N_B1_M1000_g N_B1_c_181_n
+ N_B1_M1020_g N_B1_M1027_g B1 B1 N_B1_c_183_n PM_SKY130_FD_SC_LP__A311O_4%B1
x_PM_SKY130_FD_SC_LP__A311O_4%A_111_47# N_A_111_47#_M1002_d N_A_111_47#_M1000_d
+ N_A_111_47#_M1004_s N_A_111_47#_M1013_s N_A_111_47#_M1011_g
+ N_A_111_47#_M1012_g N_A_111_47#_M1001_g N_A_111_47#_M1014_g
+ N_A_111_47#_M1003_g N_A_111_47#_M1021_g N_A_111_47#_c_251_n
+ N_A_111_47#_M1009_g N_A_111_47#_c_238_n N_A_111_47#_c_239_n
+ N_A_111_47#_M1015_g N_A_111_47#_c_422_p N_A_111_47#_c_240_n
+ N_A_111_47#_c_241_n N_A_111_47#_c_419_p N_A_111_47#_c_242_n
+ N_A_111_47#_c_322_p N_A_111_47#_c_256_n N_A_111_47#_c_243_n
+ N_A_111_47#_c_332_p N_A_111_47#_c_327_p N_A_111_47#_c_285_p
+ N_A_111_47#_c_244_n N_A_111_47#_c_296_p N_A_111_47#_c_245_n
+ N_A_111_47#_c_246_n N_A_111_47#_c_247_n N_A_111_47#_c_375_p
+ N_A_111_47#_c_286_p N_A_111_47#_c_248_n PM_SKY130_FD_SC_LP__A311O_4%A_111_47#
x_PM_SKY130_FD_SC_LP__A311O_4%A3 N_A3_c_434_n N_A3_M1005_g N_A3_c_435_n
+ N_A3_c_436_n N_A3_c_437_n N_A3_M1016_g N_A3_M1007_g N_A3_M1023_g A3 A3
+ N_A3_c_439_n PM_SKY130_FD_SC_LP__A311O_4%A3
x_PM_SKY130_FD_SC_LP__A311O_4%A2 N_A2_M1006_g N_A2_M1017_g N_A2_M1025_g
+ N_A2_M1018_g A2 N_A2_c_499_n N_A2_c_500_n PM_SKY130_FD_SC_LP__A311O_4%A2
x_PM_SKY130_FD_SC_LP__A311O_4%A1 N_A1_c_545_n N_A1_M1004_g N_A1_M1008_g
+ N_A1_c_547_n N_A1_M1022_g N_A1_M1019_g A1 A1 N_A1_c_550_n
+ PM_SKY130_FD_SC_LP__A311O_4%A1
x_PM_SKY130_FD_SC_LP__A311O_4%A_28_367# N_A_28_367#_M1013_d N_A_28_367#_M1026_d
+ N_A_28_367#_M1027_d N_A_28_367#_c_592_n N_A_28_367#_c_593_n
+ N_A_28_367#_c_599_n N_A_28_367#_c_601_n N_A_28_367#_c_608_n
+ N_A_28_367#_c_610_n N_A_28_367#_c_603_n PM_SKY130_FD_SC_LP__A311O_4%A_28_367#
x_PM_SKY130_FD_SC_LP__A311O_4%A_283_367# N_A_283_367#_M1024_s
+ N_A_283_367#_M1007_s N_A_283_367#_M1017_s N_A_283_367#_M1008_s
+ N_A_283_367#_c_635_n N_A_283_367#_c_636_n N_A_283_367#_c_637_n
+ N_A_283_367#_c_638_n N_A_283_367#_c_697_p N_A_283_367#_c_664_n
+ N_A_283_367#_c_704_p N_A_283_367#_c_665_n N_A_283_367#_c_705_p
+ N_A_283_367#_c_639_n N_A_283_367#_c_644_n N_A_283_367#_c_669_n
+ N_A_283_367#_c_672_n PM_SKY130_FD_SC_LP__A311O_4%A_283_367#
x_PM_SKY130_FD_SC_LP__A311O_4%VPWR N_VPWR_M1001_d N_VPWR_M1003_d N_VPWR_M1015_d
+ N_VPWR_M1023_d N_VPWR_M1025_d N_VPWR_M1019_d N_VPWR_c_719_n N_VPWR_c_720_n
+ N_VPWR_c_721_n N_VPWR_c_722_n N_VPWR_c_723_n N_VPWR_c_724_n N_VPWR_c_725_n
+ N_VPWR_c_726_n N_VPWR_c_727_n N_VPWR_c_728_n VPWR N_VPWR_c_729_n
+ N_VPWR_c_730_n N_VPWR_c_731_n N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n
+ N_VPWR_c_735_n N_VPWR_c_736_n N_VPWR_c_718_n PM_SKY130_FD_SC_LP__A311O_4%VPWR
x_PM_SKY130_FD_SC_LP__A311O_4%X N_X_M1011_d N_X_M1014_d N_X_M1001_s N_X_M1009_s
+ N_X_c_897_p N_X_c_837_n N_X_c_838_n N_X_c_843_n N_X_c_894_p N_X_c_839_n
+ N_X_c_840_n N_X_c_841_n X N_X_c_842_n PM_SKY130_FD_SC_LP__A311O_4%X
x_PM_SKY130_FD_SC_LP__A311O_4%VGND N_VGND_M1002_s N_VGND_M1010_s N_VGND_M1020_s
+ N_VGND_M1012_s N_VGND_M1021_s N_VGND_M1016_s N_VGND_c_906_n N_VGND_c_907_n
+ N_VGND_c_908_n N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n N_VGND_c_912_n
+ N_VGND_c_913_n N_VGND_c_914_n N_VGND_c_915_n N_VGND_c_916_n N_VGND_c_917_n
+ VGND N_VGND_c_918_n N_VGND_c_919_n N_VGND_c_920_n N_VGND_c_921_n
+ N_VGND_c_922_n N_VGND_c_923_n N_VGND_c_924_n PM_SKY130_FD_SC_LP__A311O_4%VGND
x_PM_SKY130_FD_SC_LP__A311O_4%A_877_47# N_A_877_47#_M1005_d N_A_877_47#_M1006_s
+ N_A_877_47#_c_1036_n N_A_877_47#_c_1013_n N_A_877_47#_c_1014_n
+ N_A_877_47#_c_1044_p N_A_877_47#_c_1015_n N_A_877_47#_c_1016_n
+ PM_SKY130_FD_SC_LP__A311O_4%A_877_47#
x_PM_SKY130_FD_SC_LP__A311O_4%A_1098_69# N_A_1098_69#_M1006_d
+ N_A_1098_69#_M1018_d N_A_1098_69#_M1022_d N_A_1098_69#_c_1045_n
+ N_A_1098_69#_c_1046_n N_A_1098_69#_c_1047_n N_A_1098_69#_c_1051_n
+ N_A_1098_69#_c_1048_n N_A_1098_69#_c_1049_n N_A_1098_69#_c_1050_n
+ PM_SKY130_FD_SC_LP__A311O_4%A_1098_69#
cc_1 VNB N_C1_M1002_g 0.0231841f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.655
cc_2 VNB N_C1_M1013_g 0.00703468f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_3 VNB N_C1_M1010_g 0.0166425f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.655
cc_4 VNB N_C1_M1026_g 0.00493246f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_5 VNB C1 0.0201069f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_C1_c_138_n 0.0629515f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.375
cc_7 VNB N_B1_M1000_g 0.0207369f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_8 VNB N_B1_c_181_n 0.044964f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.21
cc_9 VNB N_B1_M1020_g 0.0200516f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.655
cc_10 VNB N_B1_c_183_n 0.0019519f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.375
cc_11 VNB N_A_111_47#_M1011_g 0.0203838f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_12 VNB N_A_111_47#_M1012_g 0.0200476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_111_47#_M1014_g 0.0200544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_111_47#_M1021_g 0.0233758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_111_47#_c_238_n 0.0156564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_111_47#_c_239_n 0.0906629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_111_47#_c_240_n 0.00134204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_111_47#_c_241_n 0.00731317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_111_47#_c_242_n 0.00613969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_111_47#_c_243_n 9.74151e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_111_47#_c_244_n 4.69647e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_111_47#_c_245_n 0.0014391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_111_47#_c_246_n 0.00167068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_111_47#_c_247_n 0.00465761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_111_47#_c_248_n 0.00896824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A3_c_434_n 0.0167854f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.21
cc_27 VNB N_A3_c_435_n 0.0132036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A3_c_436_n 0.0102946f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.54
cc_29 VNB N_A3_c_437_n 0.0172446f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_30 VNB A3 0.00476478f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB N_A3_c_439_n 0.0720228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_M1006_g 0.0229828f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.655
cc_33 VNB N_A2_M1018_g 0.019905f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_34 VNB N_A2_c_499_n 0.00162563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_c_500_n 0.0404894f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.375
cc_36 VNB N_A1_c_545_n 0.0159789f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.21
cc_37 VNB N_A1_M1008_g 0.00122435f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_38 VNB N_A1_c_547_n 0.0191005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A1_M1019_g 0.00149052f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.54
cc_40 VNB A1 0.0201525f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=2.465
cc_41 VNB N_A1_c_550_n 0.0687329f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.375
cc_42 VNB N_VPWR_c_718_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_837_n 0.00304439f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_44 VNB N_X_c_838_n 0.00226637f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_45 VNB N_X_c_839_n 0.00613616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_X_c_840_n 0.00532738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_X_c_841_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0.257 $Y2=1.665
cc_48 VNB N_X_c_842_n 0.00639593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_906_n 0.0105251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_907_n 0.0340281f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.375
cc_51 VNB N_VGND_c_908_n 0.00215937f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.375
cc_52 VNB N_VGND_c_909_n 3.15299e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_910_n 3.10897e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_911_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_912_n 0.00174197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_913_n 0.00275589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_914_n 0.0145469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_915_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_916_n 0.013305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_917_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_918_n 0.013276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_919_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_920_n 0.0630861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_921_n 0.391148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_922_n 0.00522308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_923_n 0.010461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_924_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_877_47#_c_1013_n 5.21048e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_877_47#_c_1014_n 0.00377476f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.54
cc_70 VNB N_A_877_47#_c_1015_n 0.00202686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_877_47#_c_1016_n 0.00807867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1098_69#_c_1045_n 0.00489145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1098_69#_c_1046_n 0.00259172f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.465
cc_74 VNB N_A_1098_69#_c_1047_n 0.00434252f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=2.465
cc_75 VNB N_A_1098_69#_c_1048_n 0.011971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1098_69#_c_1049_n 0.023359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1098_69#_c_1050_n 0.00167433f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=1.375
cc_78 VPB N_C1_M1013_g 0.0259851f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_79 VPB N_C1_M1026_g 0.0195402f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_80 VPB C1 0.00714594f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_81 VPB N_B1_M1024_g 0.0192422f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.655
cc_82 VPB N_B1_c_181_n 0.0073844f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.21
cc_83 VPB N_B1_M1027_g 0.0270413f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_84 VPB N_B1_c_183_n 0.00682947f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.375
cc_85 VPB N_A_111_47#_M1001_g 0.0214627f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.375
cc_86 VPB N_A_111_47#_M1003_g 0.0201418f $X=-0.19 $Y=1.655 $X2=0.257 $Y2=1.665
cc_87 VPB N_A_111_47#_c_251_n 0.0167539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_111_47#_c_238_n 0.0152813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_111_47#_c_239_n 0.0349134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_111_47#_M1015_g 0.0195108f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_111_47#_c_240_n 0.00339243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_111_47#_c_256_n 0.00686688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_111_47#_c_244_n 0.00141617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A3_M1007_g 0.0185025f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.655
cc_95 VPB N_A3_M1023_g 0.0185253f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_96 VPB A3 0.0049778f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_97 VPB N_A3_c_439_n 0.00373829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A2_M1017_g 0.0184976f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_99 VPB N_A2_M1025_g 0.0190886f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.655
cc_100 VPB N_A2_c_499_n 0.00346618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A2_c_500_n 0.00807368f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.375
cc_102 VPB N_A1_M1008_g 0.0198797f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_103 VPB N_A1_M1019_g 0.0244545f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.54
cc_104 VPB A1 0.00754493f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_105 VPB N_A_28_367#_c_592_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.655
cc_106 VPB N_A_28_367#_c_593_n 0.0384572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_283_367#_c_635_n 0.0105539f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.465
cc_108 VPB N_A_283_367#_c_636_n 0.00994071f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_109 VPB N_A_283_367#_c_637_n 0.00210573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_283_367#_c_638_n 0.00450419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_283_367#_c_639_n 0.00179998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_719_n 0.0093642f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.375
cc_113 VPB N_VPWR_c_720_n 0.0068491f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.375
cc_114 VPB N_VPWR_c_721_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_722_n 0.0121672f $X=-0.19 $Y=1.655 $X2=0.257 $Y2=1.665
cc_116 VPB N_VPWR_c_723_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_724_n 0.00431378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_725_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_726_n 0.0482594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_727_n 0.0202541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_728_n 0.00436154f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_729_n 0.0601954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_730_n 0.0186999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_731_n 0.0149122f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_732_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_733_n 0.00631443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_734_n 0.00631443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_735_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_736_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_718_n 0.0586719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_X_c_843_n 0.00657499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_X_c_842_n 0.00401287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 N_C1_M1026_g N_B1_M1024_g 0.019907f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_134 N_C1_M1010_g N_B1_M1000_g 0.0182554f $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_135 N_C1_c_138_n N_B1_c_181_n 0.0260575f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_136 N_C1_M1026_g N_B1_c_183_n 0.00433734f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_137 N_C1_c_138_n N_B1_c_183_n 0.00337638f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_138 N_C1_M1013_g N_A_111_47#_c_240_n 0.00423221f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_139 N_C1_M1026_g N_A_111_47#_c_240_n 0.00427902f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_140 C1 N_A_111_47#_c_240_n 0.0372118f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_141 N_C1_c_138_n N_A_111_47#_c_240_n 0.0160369f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_142 N_C1_M1010_g N_A_111_47#_c_241_n 0.0112003f $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_143 N_C1_c_138_n N_A_111_47#_c_241_n 0.008348f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_144 N_C1_M1002_g N_A_111_47#_c_245_n 0.0042928f $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_145 C1 N_A_111_47#_c_245_n 0.00280287f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_146 N_C1_c_138_n N_A_111_47#_c_245_n 0.00442282f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_147 N_C1_M1013_g N_A_28_367#_c_592_n 5.81207e-19 $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_148 N_C1_M1013_g N_A_28_367#_c_593_n 0.0140518f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_149 N_C1_M1026_g N_A_28_367#_c_593_n 6.6542e-19 $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_150 C1 N_A_28_367#_c_593_n 0.026915f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_151 N_C1_c_138_n N_A_28_367#_c_593_n 0.00108305f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_152 N_C1_M1013_g N_A_28_367#_c_599_n 0.0105205f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_153 N_C1_M1026_g N_A_28_367#_c_599_n 0.0105205f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_154 N_C1_M1013_g N_A_28_367#_c_601_n 6.6542e-19 $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_155 N_C1_M1026_g N_A_28_367#_c_601_n 0.0131354f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_156 N_C1_M1026_g N_A_28_367#_c_603_n 5.89773e-19 $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_157 N_C1_M1013_g N_VPWR_c_729_n 0.00357842f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_158 N_C1_M1026_g N_VPWR_c_729_n 0.00357842f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_159 N_C1_M1013_g N_VPWR_c_718_n 0.00628849f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_160 N_C1_M1026_g N_VPWR_c_718_n 0.00537652f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_161 N_C1_M1002_g N_VGND_c_907_n 0.016591f $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_162 N_C1_M1010_g N_VGND_c_907_n 6.78137e-19 $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_163 C1 N_VGND_c_907_n 0.02584f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_164 N_C1_c_138_n N_VGND_c_907_n 0.00176637f $X=0.91 $Y=1.375 $X2=0 $Y2=0
cc_165 N_C1_M1002_g N_VGND_c_908_n 6.16093e-19 $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_166 N_C1_M1010_g N_VGND_c_908_n 0.0103732f $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_167 N_C1_M1002_g N_VGND_c_918_n 0.00486043f $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_168 N_C1_M1010_g N_VGND_c_918_n 0.00544582f $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_169 N_C1_M1002_g N_VGND_c_921_n 0.00824727f $X=0.48 $Y=0.655 $X2=0 $Y2=0
cc_170 N_C1_M1010_g N_VGND_c_921_n 0.009174f $X=0.91 $Y=0.655 $X2=0 $Y2=0
cc_171 N_B1_M1020_g N_A_111_47#_M1011_g 0.0167953f $X=1.81 $Y=0.655 $X2=0 $Y2=0
cc_172 N_B1_c_181_n N_A_111_47#_c_239_n 0.0167953f $X=1.81 $Y=1.29 $X2=0 $Y2=0
cc_173 N_B1_c_183_n N_A_111_47#_c_239_n 3.73173e-19 $X=1.7 $Y=1.5 $X2=0 $Y2=0
cc_174 N_B1_c_181_n N_A_111_47#_c_240_n 7.21418e-19 $X=1.81 $Y=1.29 $X2=0 $Y2=0
cc_175 N_B1_c_183_n N_A_111_47#_c_240_n 0.0251678f $X=1.7 $Y=1.5 $X2=0 $Y2=0
cc_176 N_B1_M1000_g N_A_111_47#_c_241_n 0.0152057f $X=1.38 $Y=0.655 $X2=0 $Y2=0
cc_177 N_B1_c_181_n N_A_111_47#_c_241_n 0.00309106f $X=1.81 $Y=1.29 $X2=0 $Y2=0
cc_178 N_B1_c_183_n N_A_111_47#_c_241_n 0.0382103f $X=1.7 $Y=1.5 $X2=0 $Y2=0
cc_179 N_B1_M1020_g N_A_111_47#_c_242_n 0.0138701f $X=1.81 $Y=0.655 $X2=0 $Y2=0
cc_180 N_B1_c_183_n N_A_111_47#_c_242_n 0.0126439f $X=1.7 $Y=1.5 $X2=0 $Y2=0
cc_181 N_B1_c_181_n N_A_111_47#_c_246_n 0.00278388f $X=1.81 $Y=1.29 $X2=0 $Y2=0
cc_182 N_B1_c_183_n N_A_111_47#_c_246_n 0.0181513f $X=1.7 $Y=1.5 $X2=0 $Y2=0
cc_183 N_B1_M1020_g N_A_111_47#_c_247_n 0.00527857f $X=1.81 $Y=0.655 $X2=0 $Y2=0
cc_184 N_B1_c_183_n N_A_111_47#_c_247_n 0.0135054f $X=1.7 $Y=1.5 $X2=0 $Y2=0
cc_185 N_B1_M1024_g N_A_28_367#_c_601_n 0.0131668f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B1_c_181_n N_A_28_367#_c_601_n 2.98561e-19 $X=1.81 $Y=1.29 $X2=0 $Y2=0
cc_187 N_B1_M1027_g N_A_28_367#_c_601_n 6.09902e-19 $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_188 N_B1_c_183_n N_A_28_367#_c_601_n 0.0222158f $X=1.7 $Y=1.5 $X2=0 $Y2=0
cc_189 N_B1_M1024_g N_A_28_367#_c_608_n 0.0106991f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_190 N_B1_M1027_g N_A_28_367#_c_608_n 0.0113012f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B1_M1024_g N_A_28_367#_c_610_n 5.67876e-19 $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_192 N_B1_M1027_g N_A_28_367#_c_610_n 0.0100161f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_193 N_B1_M1024_g N_A_28_367#_c_603_n 5.89773e-19 $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_194 N_B1_M1027_g N_A_283_367#_c_635_n 0.014386f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_195 N_B1_c_183_n N_A_283_367#_c_635_n 0.0111388f $X=1.7 $Y=1.5 $X2=0 $Y2=0
cc_196 N_B1_M1027_g N_A_283_367#_c_636_n 0.00257507f $X=1.81 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_B1_M1027_g N_A_283_367#_c_638_n 5.40627e-19 $X=1.81 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_B1_c_181_n N_A_283_367#_c_644_n 8.88905e-19 $X=1.81 $Y=1.29 $X2=0 $Y2=0
cc_199 N_B1_c_183_n N_A_283_367#_c_644_n 0.0188835f $X=1.7 $Y=1.5 $X2=0 $Y2=0
cc_200 N_B1_M1027_g N_VPWR_c_719_n 0.00198836f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_201 N_B1_M1024_g N_VPWR_c_729_n 0.00357842f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B1_M1027_g N_VPWR_c_729_n 0.00357842f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B1_M1024_g N_VPWR_c_718_n 0.00548485f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B1_M1027_g N_VPWR_c_718_n 0.0067592f $X=1.81 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B1_M1000_g N_VGND_c_908_n 0.00204792f $X=1.38 $Y=0.655 $X2=0 $Y2=0
cc_206 N_B1_M1000_g N_VGND_c_909_n 6.44001e-19 $X=1.38 $Y=0.655 $X2=0 $Y2=0
cc_207 N_B1_M1020_g N_VGND_c_909_n 0.0115568f $X=1.81 $Y=0.655 $X2=0 $Y2=0
cc_208 N_B1_M1000_g N_VGND_c_914_n 0.00583607f $X=1.38 $Y=0.655 $X2=0 $Y2=0
cc_209 N_B1_M1020_g N_VGND_c_914_n 0.00486043f $X=1.81 $Y=0.655 $X2=0 $Y2=0
cc_210 N_B1_M1000_g N_VGND_c_921_n 0.0106071f $X=1.38 $Y=0.655 $X2=0 $Y2=0
cc_211 N_B1_M1020_g N_VGND_c_921_n 0.00824727f $X=1.81 $Y=0.655 $X2=0 $Y2=0
cc_212 N_A_111_47#_M1021_g N_A3_c_434_n 0.00621809f $X=3.54 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_111_47#_c_238_n N_A3_c_436_n 0.0239735f $X=4.465 $Y=1.625 $X2=0 $Y2=0
cc_214 N_A_111_47#_c_239_n N_A3_c_436_n 0.00159971f $X=3.995 $Y=1.625 $X2=0
+ $Y2=0
cc_215 N_A_111_47#_M1015_g N_A3_M1007_g 0.0301524f $X=4.54 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A_111_47#_c_285_p N_A3_M1007_g 0.0109148f $X=6.545 $Y=2.005 $X2=0 $Y2=0
cc_217 N_A_111_47#_c_286_p N_A3_M1007_g 0.00441725f $X=4.65 $Y=2.005 $X2=0 $Y2=0
cc_218 N_A_111_47#_c_285_p N_A3_M1023_g 0.0103994f $X=6.545 $Y=2.005 $X2=0 $Y2=0
cc_219 N_A_111_47#_c_238_n A3 2.05054e-19 $X=4.465 $Y=1.625 $X2=0 $Y2=0
cc_220 N_A_111_47#_c_285_p A3 0.0472385f $X=6.545 $Y=2.005 $X2=0 $Y2=0
cc_221 N_A_111_47#_c_238_n N_A3_c_439_n 0.0301524f $X=4.465 $Y=1.625 $X2=0 $Y2=0
cc_222 N_A_111_47#_c_285_p N_A3_c_439_n 0.00387168f $X=6.545 $Y=2.005 $X2=0
+ $Y2=0
cc_223 N_A_111_47#_c_286_p N_A3_c_439_n 3.36791e-19 $X=4.65 $Y=2.005 $X2=0 $Y2=0
cc_224 N_A_111_47#_c_285_p N_A2_M1017_g 0.011041f $X=6.545 $Y=2.005 $X2=0 $Y2=0
cc_225 N_A_111_47#_c_285_p N_A2_M1025_g 0.0108435f $X=6.545 $Y=2.005 $X2=0 $Y2=0
cc_226 N_A_111_47#_c_244_n N_A2_M1025_g 0.00368345f $X=6.63 $Y=1.92 $X2=0 $Y2=0
cc_227 N_A_111_47#_c_296_p N_A2_M1018_g 9.66569e-19 $X=6.98 $Y=0.68 $X2=0 $Y2=0
cc_228 N_A_111_47#_c_285_p N_A2_c_499_n 0.0401834f $X=6.545 $Y=2.005 $X2=0 $Y2=0
cc_229 N_A_111_47#_c_244_n N_A2_c_499_n 0.00860235f $X=6.63 $Y=1.92 $X2=0 $Y2=0
cc_230 N_A_111_47#_c_248_n N_A2_c_499_n 0.0259449f $X=6.98 $Y=1.495 $X2=0 $Y2=0
cc_231 N_A_111_47#_c_285_p N_A2_c_500_n 0.00288103f $X=6.545 $Y=2.005 $X2=0
+ $Y2=0
cc_232 N_A_111_47#_c_244_n N_A2_c_500_n 2.20623e-19 $X=6.63 $Y=1.92 $X2=0 $Y2=0
cc_233 N_A_111_47#_c_248_n N_A2_c_500_n 0.002445f $X=6.98 $Y=1.495 $X2=0 $Y2=0
cc_234 N_A_111_47#_c_296_p N_A1_c_545_n 0.00966336f $X=6.98 $Y=0.68 $X2=-0.19
+ $Y2=-0.245
cc_235 N_A_111_47#_c_285_p N_A1_M1008_g 0.004475f $X=6.545 $Y=2.005 $X2=0 $Y2=0
cc_236 N_A_111_47#_c_244_n N_A1_M1008_g 0.00657276f $X=6.63 $Y=1.92 $X2=0 $Y2=0
cc_237 N_A_111_47#_c_248_n N_A1_M1008_g 0.0042375f $X=6.98 $Y=1.495 $X2=0 $Y2=0
cc_238 N_A_111_47#_c_296_p N_A1_c_547_n 0.0146316f $X=6.98 $Y=0.68 $X2=0 $Y2=0
cc_239 N_A_111_47#_c_244_n N_A1_M1019_g 6.69384e-19 $X=6.63 $Y=1.92 $X2=0 $Y2=0
cc_240 N_A_111_47#_c_248_n N_A1_M1019_g 0.00158502f $X=6.98 $Y=1.495 $X2=0 $Y2=0
cc_241 N_A_111_47#_c_244_n A1 0.002998f $X=6.63 $Y=1.92 $X2=0 $Y2=0
cc_242 N_A_111_47#_c_296_p A1 0.0103071f $X=6.98 $Y=0.68 $X2=0 $Y2=0
cc_243 N_A_111_47#_c_248_n A1 0.0233062f $X=6.98 $Y=1.495 $X2=0 $Y2=0
cc_244 N_A_111_47#_c_296_p N_A1_c_550_n 0.00646747f $X=6.98 $Y=0.68 $X2=0 $Y2=0
cc_245 N_A_111_47#_c_248_n N_A1_c_550_n 0.0261836f $X=6.98 $Y=1.495 $X2=0 $Y2=0
cc_246 N_A_111_47#_M1013_s N_A_28_367#_c_599_n 0.00332344f $X=0.555 $Y=1.835
+ $X2=0 $Y2=0
cc_247 N_A_111_47#_c_240_n N_A_28_367#_c_599_n 0.0126348f $X=0.695 $Y=2.095
+ $X2=0 $Y2=0
cc_248 N_A_111_47#_c_241_n N_A_28_367#_c_601_n 2.15591e-19 $X=1.475 $Y=1.16
+ $X2=0 $Y2=0
cc_249 N_A_111_47#_c_285_p N_A_283_367#_M1007_s 0.00333177f $X=6.545 $Y=2.005
+ $X2=0 $Y2=0
cc_250 N_A_111_47#_c_285_p N_A_283_367#_M1017_s 0.00332475f $X=6.545 $Y=2.005
+ $X2=0 $Y2=0
cc_251 N_A_111_47#_c_239_n N_A_283_367#_c_635_n 0.00692364f $X=3.995 $Y=1.625
+ $X2=0 $Y2=0
cc_252 N_A_111_47#_c_242_n N_A_283_367#_c_635_n 0.00377709f $X=2.035 $Y=1.16
+ $X2=0 $Y2=0
cc_253 N_A_111_47#_c_322_p N_A_283_367#_c_635_n 0.0121501f $X=2.64 $Y=1.475
+ $X2=0 $Y2=0
cc_254 N_A_111_47#_c_256_n N_A_283_367#_c_635_n 0.0135569f $X=2.725 $Y=2.185
+ $X2=0 $Y2=0
cc_255 N_A_111_47#_c_247_n N_A_283_367#_c_635_n 0.00834694f $X=2.12 $Y=1.16
+ $X2=0 $Y2=0
cc_256 N_A_111_47#_M1001_g N_A_283_367#_c_636_n 0.00540788f $X=2.94 $Y=2.405
+ $X2=0 $Y2=0
cc_257 N_A_111_47#_c_256_n N_A_283_367#_c_636_n 0.00667094f $X=2.725 $Y=2.185
+ $X2=0 $Y2=0
cc_258 N_A_111_47#_c_327_p N_A_283_367#_c_636_n 0.0134822f $X=2.81 $Y=2.27 $X2=0
+ $Y2=0
cc_259 N_A_111_47#_M1001_g N_A_283_367#_c_637_n 0.013664f $X=2.94 $Y=2.405 $X2=0
+ $Y2=0
cc_260 N_A_111_47#_M1003_g N_A_283_367#_c_637_n 0.012421f $X=3.37 $Y=2.405 $X2=0
+ $Y2=0
cc_261 N_A_111_47#_c_251_n N_A_283_367#_c_637_n 0.0133381f $X=3.92 $Y=1.7 $X2=0
+ $Y2=0
cc_262 N_A_111_47#_M1015_g N_A_283_367#_c_637_n 0.0124752f $X=4.54 $Y=2.465
+ $X2=0 $Y2=0
cc_263 N_A_111_47#_c_332_p N_A_283_367#_c_637_n 0.0959669f $X=4.565 $Y=2.27
+ $X2=0 $Y2=0
cc_264 N_A_111_47#_c_327_p N_A_283_367#_c_637_n 0.0136234f $X=2.81 $Y=2.27 $X2=0
+ $Y2=0
cc_265 N_A_111_47#_c_285_p N_A_283_367#_c_637_n 0.00770503f $X=6.545 $Y=2.005
+ $X2=0 $Y2=0
cc_266 N_A_111_47#_c_286_p N_A_283_367#_c_637_n 0.00846276f $X=4.65 $Y=2.005
+ $X2=0 $Y2=0
cc_267 N_A_111_47#_c_285_p N_A_283_367#_c_664_n 0.0323235f $X=6.545 $Y=2.005
+ $X2=0 $Y2=0
cc_268 N_A_111_47#_c_285_p N_A_283_367#_c_665_n 0.0299276f $X=6.545 $Y=2.005
+ $X2=0 $Y2=0
cc_269 N_A_111_47#_c_248_n N_A_283_367#_c_665_n 0.00315294f $X=6.98 $Y=1.495
+ $X2=0 $Y2=0
cc_270 N_A_111_47#_c_244_n N_A_283_367#_c_639_n 0.00425162f $X=6.63 $Y=1.92
+ $X2=0 $Y2=0
cc_271 N_A_111_47#_c_248_n N_A_283_367#_c_639_n 0.0165165f $X=6.98 $Y=1.495
+ $X2=0 $Y2=0
cc_272 N_A_111_47#_M1015_g N_A_283_367#_c_669_n 9.99886e-19 $X=4.54 $Y=2.465
+ $X2=0 $Y2=0
cc_273 N_A_111_47#_c_285_p N_A_283_367#_c_669_n 0.0152279f $X=6.545 $Y=2.005
+ $X2=0 $Y2=0
cc_274 N_A_111_47#_c_286_p N_A_283_367#_c_669_n 0.00463238f $X=4.65 $Y=2.005
+ $X2=0 $Y2=0
cc_275 N_A_111_47#_c_285_p N_A_283_367#_c_672_n 0.0135055f $X=6.545 $Y=2.005
+ $X2=0 $Y2=0
cc_276 N_A_111_47#_c_256_n N_VPWR_M1001_d 0.0107934f $X=2.725 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_277 N_A_111_47#_c_327_p N_VPWR_M1001_d 0.004208f $X=2.81 $Y=2.27 $X2=-0.19
+ $Y2=-0.245
cc_278 N_A_111_47#_c_332_p N_VPWR_M1003_d 0.00624971f $X=4.565 $Y=2.27 $X2=0
+ $Y2=0
cc_279 N_A_111_47#_c_285_p N_VPWR_M1015_d 0.00382665f $X=6.545 $Y=2.005 $X2=0
+ $Y2=0
cc_280 N_A_111_47#_c_286_p N_VPWR_M1015_d 0.00471232f $X=4.65 $Y=2.005 $X2=0
+ $Y2=0
cc_281 N_A_111_47#_c_285_p N_VPWR_M1023_d 0.00609528f $X=6.545 $Y=2.005 $X2=0
+ $Y2=0
cc_282 N_A_111_47#_c_285_p N_VPWR_M1025_d 0.0070001f $X=6.545 $Y=2.005 $X2=0
+ $Y2=0
cc_283 N_A_111_47#_c_244_n N_VPWR_M1025_d 0.00100244f $X=6.63 $Y=1.92 $X2=0
+ $Y2=0
cc_284 N_A_111_47#_M1001_g N_VPWR_c_719_n 0.0117977f $X=2.94 $Y=2.405 $X2=0
+ $Y2=0
cc_285 N_A_111_47#_M1003_g N_VPWR_c_720_n 0.00437514f $X=3.37 $Y=2.405 $X2=0
+ $Y2=0
cc_286 N_A_111_47#_c_251_n N_VPWR_c_720_n 0.00437514f $X=3.92 $Y=1.7 $X2=0 $Y2=0
cc_287 N_A_111_47#_M1015_g N_VPWR_c_720_n 0.00132311f $X=4.54 $Y=2.465 $X2=0
+ $Y2=0
cc_288 N_A_111_47#_c_251_n N_VPWR_c_721_n 0.00145215f $X=3.92 $Y=1.7 $X2=0 $Y2=0
cc_289 N_A_111_47#_M1015_g N_VPWR_c_721_n 0.00993247f $X=4.54 $Y=2.465 $X2=0
+ $Y2=0
cc_290 N_A_111_47#_c_251_n N_VPWR_c_727_n 0.00377654f $X=3.92 $Y=1.7 $X2=0 $Y2=0
cc_291 N_A_111_47#_M1015_g N_VPWR_c_727_n 0.00353537f $X=4.54 $Y=2.465 $X2=0
+ $Y2=0
cc_292 N_A_111_47#_M1001_g N_VPWR_c_730_n 0.00377654f $X=2.94 $Y=2.405 $X2=0
+ $Y2=0
cc_293 N_A_111_47#_M1003_g N_VPWR_c_730_n 0.00377654f $X=3.37 $Y=2.405 $X2=0
+ $Y2=0
cc_294 N_A_111_47#_M1013_s N_VPWR_c_718_n 0.00225186f $X=0.555 $Y=1.835 $X2=0
+ $Y2=0
cc_295 N_A_111_47#_M1001_g N_VPWR_c_718_n 0.00608061f $X=2.94 $Y=2.405 $X2=0
+ $Y2=0
cc_296 N_A_111_47#_M1003_g N_VPWR_c_718_n 0.00535745f $X=3.37 $Y=2.405 $X2=0
+ $Y2=0
cc_297 N_A_111_47#_c_251_n N_VPWR_c_718_n 0.00561339f $X=3.92 $Y=1.7 $X2=0 $Y2=0
cc_298 N_A_111_47#_M1015_g N_VPWR_c_718_n 0.00504766f $X=4.54 $Y=2.465 $X2=0
+ $Y2=0
cc_299 N_A_111_47#_c_332_p N_X_M1001_s 0.00343895f $X=4.565 $Y=2.27 $X2=0 $Y2=0
cc_300 N_A_111_47#_c_332_p N_X_M1009_s 0.00832484f $X=4.565 $Y=2.27 $X2=0 $Y2=0
cc_301 N_A_111_47#_M1012_g N_X_c_837_n 0.0133482f $X=2.68 $Y=0.655 $X2=0 $Y2=0
cc_302 N_A_111_47#_M1014_g N_X_c_837_n 0.0136472f $X=3.11 $Y=0.655 $X2=0 $Y2=0
cc_303 N_A_111_47#_c_239_n N_X_c_837_n 0.00280857f $X=3.995 $Y=1.625 $X2=0 $Y2=0
cc_304 N_A_111_47#_c_322_p N_X_c_837_n 0.00562838f $X=2.64 $Y=1.475 $X2=0 $Y2=0
cc_305 N_A_111_47#_c_243_n N_X_c_837_n 0.0294091f $X=3.7 $Y=1.45 $X2=0 $Y2=0
cc_306 N_A_111_47#_c_375_p N_X_c_837_n 0.0131564f $X=2.68 $Y=1.45 $X2=0 $Y2=0
cc_307 N_A_111_47#_M1011_g N_X_c_838_n 9.75596e-19 $X=2.25 $Y=0.655 $X2=0 $Y2=0
cc_308 N_A_111_47#_c_239_n N_X_c_838_n 0.00256759f $X=3.995 $Y=1.625 $X2=0 $Y2=0
cc_309 N_A_111_47#_c_322_p N_X_c_838_n 0.015182f $X=2.64 $Y=1.475 $X2=0 $Y2=0
cc_310 N_A_111_47#_c_247_n N_X_c_838_n 0.00963391f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A_111_47#_M1001_g N_X_c_843_n 0.00388757f $X=2.94 $Y=2.405 $X2=0 $Y2=0
cc_312 N_A_111_47#_M1003_g N_X_c_843_n 0.0125462f $X=3.37 $Y=2.405 $X2=0 $Y2=0
cc_313 N_A_111_47#_c_251_n N_X_c_843_n 0.0170616f $X=3.92 $Y=1.7 $X2=0 $Y2=0
cc_314 N_A_111_47#_c_239_n N_X_c_843_n 0.00849333f $X=3.995 $Y=1.625 $X2=0 $Y2=0
cc_315 N_A_111_47#_c_256_n N_X_c_843_n 0.0114138f $X=2.725 $Y=2.185 $X2=0 $Y2=0
cc_316 N_A_111_47#_c_243_n N_X_c_843_n 0.0536652f $X=3.7 $Y=1.45 $X2=0 $Y2=0
cc_317 N_A_111_47#_c_332_p N_X_c_843_n 0.0572542f $X=4.565 $Y=2.27 $X2=0 $Y2=0
cc_318 N_A_111_47#_M1021_g N_X_c_839_n 0.0149436f $X=3.54 $Y=0.655 $X2=0 $Y2=0
cc_319 N_A_111_47#_c_238_n N_X_c_839_n 0.00155307f $X=4.465 $Y=1.625 $X2=0 $Y2=0
cc_320 N_A_111_47#_c_239_n N_X_c_839_n 0.0101235f $X=3.995 $Y=1.625 $X2=0 $Y2=0
cc_321 N_A_111_47#_c_243_n N_X_c_839_n 0.0312279f $X=3.7 $Y=1.45 $X2=0 $Y2=0
cc_322 N_A_111_47#_M1021_g N_X_c_840_n 0.00151396f $X=3.54 $Y=0.655 $X2=0 $Y2=0
cc_323 N_A_111_47#_c_239_n N_X_c_840_n 0.00256769f $X=3.995 $Y=1.625 $X2=0 $Y2=0
cc_324 N_A_111_47#_c_243_n N_X_c_840_n 0.00277424f $X=3.7 $Y=1.45 $X2=0 $Y2=0
cc_325 N_A_111_47#_c_239_n N_X_c_841_n 0.00299787f $X=3.995 $Y=1.625 $X2=0 $Y2=0
cc_326 N_A_111_47#_c_243_n N_X_c_841_n 0.0153308f $X=3.7 $Y=1.45 $X2=0 $Y2=0
cc_327 N_A_111_47#_M1003_g N_X_c_842_n 3.33936e-19 $X=3.37 $Y=2.405 $X2=0 $Y2=0
cc_328 N_A_111_47#_c_251_n N_X_c_842_n 0.00164598f $X=3.92 $Y=1.7 $X2=0 $Y2=0
cc_329 N_A_111_47#_c_238_n N_X_c_842_n 0.0259365f $X=4.465 $Y=1.625 $X2=0 $Y2=0
cc_330 N_A_111_47#_c_239_n N_X_c_842_n 0.00347889f $X=3.995 $Y=1.625 $X2=0 $Y2=0
cc_331 N_A_111_47#_M1015_g N_X_c_842_n 0.0114364f $X=4.54 $Y=2.465 $X2=0 $Y2=0
cc_332 N_A_111_47#_c_243_n N_X_c_842_n 0.0103452f $X=3.7 $Y=1.45 $X2=0 $Y2=0
cc_333 N_A_111_47#_c_332_p N_X_c_842_n 0.0322705f $X=4.565 $Y=2.27 $X2=0 $Y2=0
cc_334 N_A_111_47#_c_286_p N_X_c_842_n 0.0181961f $X=4.65 $Y=2.005 $X2=0 $Y2=0
cc_335 N_A_111_47#_c_247_n N_VGND_M1020_s 0.00152477f $X=2.12 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_A_111_47#_c_241_n N_VGND_c_908_n 0.0219498f $X=1.475 $Y=1.16 $X2=0
+ $Y2=0
cc_337 N_A_111_47#_M1011_g N_VGND_c_909_n 0.0108669f $X=2.25 $Y=0.655 $X2=0
+ $Y2=0
cc_338 N_A_111_47#_M1012_g N_VGND_c_909_n 6.36634e-19 $X=2.68 $Y=0.655 $X2=0
+ $Y2=0
cc_339 N_A_111_47#_c_242_n N_VGND_c_909_n 0.0116313f $X=2.035 $Y=1.16 $X2=0
+ $Y2=0
cc_340 N_A_111_47#_c_247_n N_VGND_c_909_n 0.0108185f $X=2.12 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_111_47#_M1011_g N_VGND_c_910_n 6.23761e-19 $X=2.25 $Y=0.655 $X2=0
+ $Y2=0
cc_342 N_A_111_47#_M1012_g N_VGND_c_910_n 0.0104024f $X=2.68 $Y=0.655 $X2=0
+ $Y2=0
cc_343 N_A_111_47#_M1014_g N_VGND_c_910_n 0.0103791f $X=3.11 $Y=0.655 $X2=0
+ $Y2=0
cc_344 N_A_111_47#_M1021_g N_VGND_c_910_n 6.19666e-19 $X=3.54 $Y=0.655 $X2=0
+ $Y2=0
cc_345 N_A_111_47#_M1014_g N_VGND_c_911_n 0.00486043f $X=3.11 $Y=0.655 $X2=0
+ $Y2=0
cc_346 N_A_111_47#_M1021_g N_VGND_c_911_n 0.00486043f $X=3.54 $Y=0.655 $X2=0
+ $Y2=0
cc_347 N_A_111_47#_M1014_g N_VGND_c_912_n 6.33625e-19 $X=3.11 $Y=0.655 $X2=0
+ $Y2=0
cc_348 N_A_111_47#_M1021_g N_VGND_c_912_n 0.0113684f $X=3.54 $Y=0.655 $X2=0
+ $Y2=0
cc_349 N_A_111_47#_c_238_n N_VGND_c_912_n 4.50224e-19 $X=4.465 $Y=1.625 $X2=0
+ $Y2=0
cc_350 N_A_111_47#_c_419_p N_VGND_c_914_n 0.0133395f $X=1.595 $Y=0.42 $X2=0
+ $Y2=0
cc_351 N_A_111_47#_M1011_g N_VGND_c_916_n 0.00525069f $X=2.25 $Y=0.655 $X2=0
+ $Y2=0
cc_352 N_A_111_47#_M1012_g N_VGND_c_916_n 0.00486043f $X=2.68 $Y=0.655 $X2=0
+ $Y2=0
cc_353 N_A_111_47#_c_422_p N_VGND_c_918_n 0.0129847f $X=0.695 $Y=0.42 $X2=0
+ $Y2=0
cc_354 N_A_111_47#_M1002_d N_VGND_c_921_n 0.00484465f $X=0.555 $Y=0.235 $X2=0
+ $Y2=0
cc_355 N_A_111_47#_M1000_d N_VGND_c_921_n 0.00449678f $X=1.455 $Y=0.235 $X2=0
+ $Y2=0
cc_356 N_A_111_47#_M1011_g N_VGND_c_921_n 0.00886509f $X=2.25 $Y=0.655 $X2=0
+ $Y2=0
cc_357 N_A_111_47#_M1012_g N_VGND_c_921_n 0.00824727f $X=2.68 $Y=0.655 $X2=0
+ $Y2=0
cc_358 N_A_111_47#_M1014_g N_VGND_c_921_n 0.00824727f $X=3.11 $Y=0.655 $X2=0
+ $Y2=0
cc_359 N_A_111_47#_M1021_g N_VGND_c_921_n 0.00824727f $X=3.54 $Y=0.655 $X2=0
+ $Y2=0
cc_360 N_A_111_47#_c_422_p N_VGND_c_921_n 0.00789217f $X=0.695 $Y=0.42 $X2=0
+ $Y2=0
cc_361 N_A_111_47#_c_419_p N_VGND_c_921_n 0.00828095f $X=1.595 $Y=0.42 $X2=0
+ $Y2=0
cc_362 N_A_111_47#_c_248_n N_A_1098_69#_c_1051_n 0.00802942f $X=6.98 $Y=1.495
+ $X2=0 $Y2=0
cc_363 N_A_111_47#_M1004_s N_A_1098_69#_c_1048_n 0.00176461f $X=6.84 $Y=0.345
+ $X2=0 $Y2=0
cc_364 N_A_111_47#_c_296_p N_A_1098_69#_c_1048_n 0.0159805f $X=6.98 $Y=0.68
+ $X2=0 $Y2=0
cc_365 N_A3_c_439_n N_A2_M1006_g 0.0393034f $X=5.185 $Y=1.5 $X2=0 $Y2=0
cc_366 A3 N_A2_c_499_n 0.0293434f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_367 N_A3_c_439_n N_A2_c_499_n 8.1329e-19 $X=5.185 $Y=1.5 $X2=0 $Y2=0
cc_368 N_A3_M1023_g N_A2_c_500_n 0.034875f $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_369 A3 N_A2_c_500_n 0.00258367f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_370 N_A3_M1007_g N_A_283_367#_c_637_n 0.0101224f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_371 N_A3_M1023_g N_A_283_367#_c_664_n 0.0122129f $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_372 N_A3_M1007_g N_A_283_367#_c_669_n 0.00744216f $X=4.97 $Y=2.465 $X2=0
+ $Y2=0
cc_373 N_A3_M1007_g N_VPWR_c_721_n 0.00639943f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A3_M1023_g N_VPWR_c_721_n 5.09333e-19 $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_375 N_A3_M1007_g N_VPWR_c_722_n 0.00354582f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_376 N_A3_M1023_g N_VPWR_c_722_n 0.00486043f $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_377 N_A3_M1007_g N_VPWR_c_723_n 6.27441e-19 $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_378 N_A3_M1023_g N_VPWR_c_723_n 0.0111421f $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_379 N_A3_M1007_g N_VPWR_c_718_n 0.00410364f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A3_M1023_g N_VPWR_c_718_n 0.00824727f $X=5.4 $Y=2.465 $X2=0 $Y2=0
cc_381 N_A3_c_434_n N_X_c_839_n 0.00221777f $X=4.31 $Y=1.16 $X2=0 $Y2=0
cc_382 N_A3_c_436_n N_X_c_840_n 0.00392268f $X=4.385 $Y=1.25 $X2=0 $Y2=0
cc_383 N_A3_c_439_n N_X_c_840_n 0.00156373f $X=5.185 $Y=1.5 $X2=0 $Y2=0
cc_384 N_A3_c_436_n N_X_c_842_n 0.0100872f $X=4.385 $Y=1.25 $X2=0 $Y2=0
cc_385 A3 N_X_c_842_n 0.0296865f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_386 N_A3_c_439_n N_X_c_842_n 0.00234234f $X=5.185 $Y=1.5 $X2=0 $Y2=0
cc_387 N_A3_c_434_n N_VGND_c_912_n 0.0115447f $X=4.31 $Y=1.16 $X2=0 $Y2=0
cc_388 N_A3_c_437_n N_VGND_c_912_n 6.33625e-19 $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A3_c_434_n N_VGND_c_913_n 6.16837e-19 $X=4.31 $Y=1.16 $X2=0 $Y2=0
cc_390 N_A3_c_437_n N_VGND_c_913_n 0.0113905f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_391 N_A3_c_439_n N_VGND_c_913_n 0.0016113f $X=5.185 $Y=1.5 $X2=0 $Y2=0
cc_392 N_A3_c_434_n N_VGND_c_919_n 0.00486043f $X=4.31 $Y=1.16 $X2=0 $Y2=0
cc_393 N_A3_c_437_n N_VGND_c_919_n 0.00486043f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_394 N_A3_c_434_n N_VGND_c_921_n 0.00824727f $X=4.31 $Y=1.16 $X2=0 $Y2=0
cc_395 N_A3_c_437_n N_VGND_c_921_n 0.00824727f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_396 N_A3_c_434_n N_A_877_47#_c_1013_n 7.44201e-19 $X=4.31 $Y=1.16 $X2=0 $Y2=0
cc_397 N_A3_c_435_n N_A_877_47#_c_1013_n 0.00595186f $X=4.665 $Y=1.25 $X2=0
+ $Y2=0
cc_398 A3 N_A_877_47#_c_1014_n 0.0134395f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_399 N_A3_c_439_n N_A_877_47#_c_1014_n 0.0026089f $X=5.185 $Y=1.5 $X2=0 $Y2=0
cc_400 N_A3_c_435_n N_A_877_47#_c_1015_n 6.40952e-19 $X=4.665 $Y=1.25 $X2=0
+ $Y2=0
cc_401 N_A3_c_437_n N_A_877_47#_c_1015_n 0.0102265f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_402 A3 N_A_877_47#_c_1015_n 0.033765f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_403 N_A3_c_439_n N_A_877_47#_c_1015_n 0.021352f $X=5.185 $Y=1.5 $X2=0 $Y2=0
cc_404 N_A3_c_437_n N_A_877_47#_c_1016_n 0.00114292f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_405 N_A3_c_439_n N_A_877_47#_c_1016_n 0.00585389f $X=5.185 $Y=1.5 $X2=0 $Y2=0
cc_406 N_A2_M1018_g N_A1_c_545_n 0.0181985f $X=6.335 $Y=0.765 $X2=-0.19
+ $Y2=-0.245
cc_407 N_A2_M1025_g N_A1_M1008_g 0.0374041f $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_408 N_A2_c_499_n N_A1_M1008_g 2.47102e-19 $X=6.28 $Y=1.51 $X2=0 $Y2=0
cc_409 N_A2_c_499_n N_A1_c_550_n 2.55592e-19 $X=6.28 $Y=1.51 $X2=0 $Y2=0
cc_410 N_A2_c_500_n N_A1_c_550_n 0.0177423f $X=6.335 $Y=1.51 $X2=0 $Y2=0
cc_411 N_A2_M1017_g N_A_283_367#_c_664_n 0.012172f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_412 N_A2_M1025_g N_A_283_367#_c_665_n 0.0133505f $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_413 N_A2_M1017_g N_VPWR_c_723_n 0.0111872f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_414 N_A2_M1025_g N_VPWR_c_723_n 5.98522e-19 $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_415 N_A2_M1025_g N_VPWR_c_724_n 0.00272396f $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_416 N_A2_M1017_g N_VPWR_c_731_n 0.00486043f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_417 N_A2_M1025_g N_VPWR_c_731_n 0.00585385f $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_418 N_A2_M1017_g N_VPWR_c_718_n 0.00824727f $X=5.83 $Y=2.465 $X2=0 $Y2=0
cc_419 N_A2_M1025_g N_VPWR_c_718_n 0.0108404f $X=6.26 $Y=2.465 $X2=0 $Y2=0
cc_420 N_A2_M1006_g N_VGND_c_913_n 0.00225064f $X=5.83 $Y=0.765 $X2=0 $Y2=0
cc_421 N_A2_M1006_g N_VGND_c_920_n 0.0029147f $X=5.83 $Y=0.765 $X2=0 $Y2=0
cc_422 N_A2_M1018_g N_VGND_c_920_n 0.0029147f $X=6.335 $Y=0.765 $X2=0 $Y2=0
cc_423 N_A2_M1006_g N_VGND_c_921_n 0.00432836f $X=5.83 $Y=0.765 $X2=0 $Y2=0
cc_424 N_A2_M1018_g N_VGND_c_921_n 0.00403428f $X=6.335 $Y=0.765 $X2=0 $Y2=0
cc_425 N_A2_M1006_g N_A_877_47#_c_1014_n 0.0130041f $X=5.83 $Y=0.765 $X2=0 $Y2=0
cc_426 N_A2_c_499_n N_A_877_47#_c_1014_n 0.0332889f $X=6.28 $Y=1.51 $X2=0 $Y2=0
cc_427 N_A2_c_500_n N_A_877_47#_c_1014_n 0.00135247f $X=6.335 $Y=1.51 $X2=0
+ $Y2=0
cc_428 N_A2_M1006_g N_A_877_47#_c_1016_n 0.00151407f $X=5.83 $Y=0.765 $X2=0
+ $Y2=0
cc_429 N_A2_M1006_g N_A_1098_69#_c_1046_n 0.0130765f $X=5.83 $Y=0.765 $X2=0
+ $Y2=0
cc_430 N_A2_M1018_g N_A_1098_69#_c_1046_n 0.0132699f $X=6.335 $Y=0.765 $X2=0
+ $Y2=0
cc_431 N_A1_M1008_g N_A_283_367#_c_665_n 0.0150801f $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_432 N_A1_M1008_g N_A_283_367#_c_639_n 4.85022e-19 $X=6.765 $Y=2.465 $X2=0
+ $Y2=0
cc_433 N_A1_M1019_g N_A_283_367#_c_639_n 8.1712e-19 $X=7.195 $Y=2.465 $X2=0
+ $Y2=0
cc_434 N_A1_c_550_n N_A_283_367#_c_639_n 7.50045e-19 $X=7.41 $Y=1.46 $X2=0 $Y2=0
cc_435 N_A1_M1008_g N_VPWR_c_724_n 0.00269764f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_436 N_A1_M1008_g N_VPWR_c_726_n 6.48903e-19 $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_437 N_A1_M1019_g N_VPWR_c_726_n 0.0213301f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_438 A1 N_VPWR_c_726_n 0.0228788f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_439 N_A1_c_550_n N_VPWR_c_726_n 0.00147549f $X=7.41 $Y=1.46 $X2=0 $Y2=0
cc_440 N_A1_M1008_g N_VPWR_c_732_n 0.00585385f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_441 N_A1_M1019_g N_VPWR_c_732_n 0.00486043f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_442 N_A1_M1008_g N_VPWR_c_718_n 0.0108541f $X=6.765 $Y=2.465 $X2=0 $Y2=0
cc_443 N_A1_M1019_g N_VPWR_c_718_n 0.00824727f $X=7.195 $Y=2.465 $X2=0 $Y2=0
cc_444 N_A1_c_545_n N_VGND_c_920_n 0.0029147f $X=6.765 $Y=1.295 $X2=0 $Y2=0
cc_445 N_A1_c_547_n N_VGND_c_920_n 0.0029147f $X=7.195 $Y=1.295 $X2=0 $Y2=0
cc_446 N_A1_c_545_n N_VGND_c_921_n 0.00399217f $X=6.765 $Y=1.295 $X2=0 $Y2=0
cc_447 N_A1_c_547_n N_VGND_c_921_n 0.00420369f $X=7.195 $Y=1.295 $X2=0 $Y2=0
cc_448 N_A1_c_545_n N_A_1098_69#_c_1048_n 0.0121173f $X=6.765 $Y=1.295 $X2=0
+ $Y2=0
cc_449 N_A1_c_547_n N_A_1098_69#_c_1048_n 0.0128685f $X=7.195 $Y=1.295 $X2=0
+ $Y2=0
cc_450 A1 N_A_1098_69#_c_1049_n 0.0228786f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_451 N_A1_c_550_n N_A_1098_69#_c_1049_n 0.00161388f $X=7.41 $Y=1.46 $X2=0
+ $Y2=0
cc_452 N_A_28_367#_c_608_n N_A_283_367#_M1024_s 0.00412427f $X=1.86 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_453 N_A_28_367#_M1027_d N_A_283_367#_c_635_n 0.00749058f $X=1.885 $Y=1.835
+ $X2=0 $Y2=0
cc_454 N_A_28_367#_c_610_n N_A_283_367#_c_635_n 0.0161865f $X=2.025 $Y=2.425
+ $X2=0 $Y2=0
cc_455 N_A_28_367#_c_610_n N_A_283_367#_c_636_n 0.0201954f $X=2.025 $Y=2.425
+ $X2=0 $Y2=0
cc_456 N_A_28_367#_c_610_n N_A_283_367#_c_638_n 0.014539f $X=2.025 $Y=2.425
+ $X2=0 $Y2=0
cc_457 N_A_28_367#_c_608_n N_A_283_367#_c_644_n 0.0156793f $X=1.86 $Y=2.99 $X2=0
+ $Y2=0
cc_458 N_A_28_367#_c_608_n N_VPWR_c_719_n 0.00887173f $X=1.86 $Y=2.99 $X2=0
+ $Y2=0
cc_459 N_A_28_367#_c_610_n N_VPWR_c_719_n 0.00191791f $X=2.025 $Y=2.425 $X2=0
+ $Y2=0
cc_460 N_A_28_367#_c_592_n N_VPWR_c_729_n 0.0211538f $X=0.265 $Y=2.905 $X2=0
+ $Y2=0
cc_461 N_A_28_367#_c_599_n N_VPWR_c_729_n 0.0298674f $X=0.96 $Y=2.99 $X2=0 $Y2=0
cc_462 N_A_28_367#_c_608_n N_VPWR_c_729_n 0.0485798f $X=1.86 $Y=2.99 $X2=0 $Y2=0
cc_463 N_A_28_367#_c_603_n N_VPWR_c_729_n 0.01906f $X=1.125 $Y=2.91 $X2=0 $Y2=0
cc_464 N_A_28_367#_M1013_d N_VPWR_c_718_n 0.00215158f $X=0.14 $Y=1.835 $X2=0
+ $Y2=0
cc_465 N_A_28_367#_M1026_d N_VPWR_c_718_n 0.00223559f $X=0.985 $Y=1.835 $X2=0
+ $Y2=0
cc_466 N_A_28_367#_M1027_d N_VPWR_c_718_n 0.00319521f $X=1.885 $Y=1.835 $X2=0
+ $Y2=0
cc_467 N_A_28_367#_c_592_n N_VPWR_c_718_n 0.0126374f $X=0.265 $Y=2.905 $X2=0
+ $Y2=0
cc_468 N_A_28_367#_c_599_n N_VPWR_c_718_n 0.0187823f $X=0.96 $Y=2.99 $X2=0 $Y2=0
cc_469 N_A_28_367#_c_608_n N_VPWR_c_718_n 0.0302021f $X=1.86 $Y=2.99 $X2=0 $Y2=0
cc_470 N_A_28_367#_c_603_n N_VPWR_c_718_n 0.0124545f $X=1.125 $Y=2.91 $X2=0
+ $Y2=0
cc_471 N_A_283_367#_c_637_n N_VPWR_M1001_d 0.0117792f $X=5.02 $Y=2.61 $X2=-0.19
+ $Y2=1.655
cc_472 N_A_283_367#_c_637_n N_VPWR_M1003_d 0.00634171f $X=5.02 $Y=2.61 $X2=0
+ $Y2=0
cc_473 N_A_283_367#_c_637_n N_VPWR_M1015_d 0.00408251f $X=5.02 $Y=2.61 $X2=0
+ $Y2=0
cc_474 N_A_283_367#_c_664_n N_VPWR_M1023_d 0.00353353f $X=5.95 $Y=2.345 $X2=0
+ $Y2=0
cc_475 N_A_283_367#_c_665_n N_VPWR_M1025_d 0.00506674f $X=6.845 $Y=2.345 $X2=0
+ $Y2=0
cc_476 N_A_283_367#_c_637_n N_VPWR_c_719_n 0.0251179f $X=5.02 $Y=2.61 $X2=0
+ $Y2=0
cc_477 N_A_283_367#_c_637_n N_VPWR_c_720_n 0.0218033f $X=5.02 $Y=2.61 $X2=0
+ $Y2=0
cc_478 N_A_283_367#_c_637_n N_VPWR_c_721_n 0.0159984f $X=5.02 $Y=2.61 $X2=0
+ $Y2=0
cc_479 N_A_283_367#_c_637_n N_VPWR_c_722_n 0.00162329f $X=5.02 $Y=2.61 $X2=0
+ $Y2=0
cc_480 N_A_283_367#_c_697_p N_VPWR_c_722_n 0.0124525f $X=5.185 $Y=2.91 $X2=0
+ $Y2=0
cc_481 N_A_283_367#_c_669_n N_VPWR_c_722_n 8.58849e-19 $X=5.185 $Y=2.345 $X2=0
+ $Y2=0
cc_482 N_A_283_367#_c_664_n N_VPWR_c_723_n 0.0170777f $X=5.95 $Y=2.345 $X2=0
+ $Y2=0
cc_483 N_A_283_367#_c_665_n N_VPWR_c_724_n 0.0196074f $X=6.845 $Y=2.345 $X2=0
+ $Y2=0
cc_484 N_A_283_367#_c_637_n N_VPWR_c_727_n 0.0121469f $X=5.02 $Y=2.61 $X2=0
+ $Y2=0
cc_485 N_A_283_367#_c_638_n N_VPWR_c_729_n 0.00344284f $X=2.46 $Y=2.61 $X2=0
+ $Y2=0
cc_486 N_A_283_367#_c_637_n N_VPWR_c_730_n 0.0100216f $X=5.02 $Y=2.61 $X2=0
+ $Y2=0
cc_487 N_A_283_367#_c_704_p N_VPWR_c_731_n 0.0131621f $X=6.045 $Y=2.91 $X2=0
+ $Y2=0
cc_488 N_A_283_367#_c_705_p N_VPWR_c_732_n 0.0138717f $X=6.98 $Y=2.45 $X2=0
+ $Y2=0
cc_489 N_A_283_367#_M1024_s N_VPWR_c_718_n 0.00257355f $X=1.415 $Y=1.835 $X2=0
+ $Y2=0
cc_490 N_A_283_367#_M1007_s N_VPWR_c_718_n 0.00395019f $X=5.045 $Y=1.835 $X2=0
+ $Y2=0
cc_491 N_A_283_367#_M1017_s N_VPWR_c_718_n 0.00467071f $X=5.905 $Y=1.835 $X2=0
+ $Y2=0
cc_492 N_A_283_367#_M1008_s N_VPWR_c_718_n 0.00397496f $X=6.84 $Y=1.835 $X2=0
+ $Y2=0
cc_493 N_A_283_367#_c_637_n N_VPWR_c_718_n 0.0460987f $X=5.02 $Y=2.61 $X2=0
+ $Y2=0
cc_494 N_A_283_367#_c_638_n N_VPWR_c_718_n 0.00515889f $X=2.46 $Y=2.61 $X2=0
+ $Y2=0
cc_495 N_A_283_367#_c_697_p N_VPWR_c_718_n 0.00730901f $X=5.185 $Y=2.91 $X2=0
+ $Y2=0
cc_496 N_A_283_367#_c_704_p N_VPWR_c_718_n 0.00808656f $X=6.045 $Y=2.91 $X2=0
+ $Y2=0
cc_497 N_A_283_367#_c_705_p N_VPWR_c_718_n 0.00886411f $X=6.98 $Y=2.45 $X2=0
+ $Y2=0
cc_498 N_A_283_367#_c_669_n N_VPWR_c_718_n 0.00188717f $X=5.185 $Y=2.345 $X2=0
+ $Y2=0
cc_499 N_A_283_367#_c_637_n N_X_M1001_s 0.00465938f $X=5.02 $Y=2.61 $X2=0 $Y2=0
cc_500 N_A_283_367#_c_637_n N_X_M1009_s 0.0110153f $X=5.02 $Y=2.61 $X2=0 $Y2=0
cc_501 N_VPWR_c_718_n N_X_M1009_s 0.00422337f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_502 N_VPWR_M1003_d N_X_c_843_n 0.00361877f $X=3.445 $Y=1.775 $X2=0 $Y2=0
cc_503 N_X_c_837_n N_VGND_M1012_s 0.00176461f $X=3.23 $Y=1.11 $X2=0 $Y2=0
cc_504 N_X_c_839_n N_VGND_M1021_s 0.00639547f $X=4.06 $Y=1.11 $X2=0 $Y2=0
cc_505 N_X_c_837_n N_VGND_c_910_n 0.0170777f $X=3.23 $Y=1.11 $X2=0 $Y2=0
cc_506 N_X_c_894_p N_VGND_c_911_n 0.0124525f $X=3.325 $Y=0.42 $X2=0 $Y2=0
cc_507 N_X_c_839_n N_VGND_c_912_n 0.0439558f $X=4.06 $Y=1.11 $X2=0 $Y2=0
cc_508 N_X_c_842_n N_VGND_c_912_n 9.51516e-19 $X=4.392 $Y=1.882 $X2=0 $Y2=0
cc_509 N_X_c_897_p N_VGND_c_916_n 0.0122751f $X=2.465 $Y=0.42 $X2=0 $Y2=0
cc_510 N_X_M1011_d N_VGND_c_921_n 0.0055404f $X=2.325 $Y=0.235 $X2=0 $Y2=0
cc_511 N_X_M1014_d N_VGND_c_921_n 0.00536646f $X=3.185 $Y=0.235 $X2=0 $Y2=0
cc_512 N_X_c_897_p N_VGND_c_921_n 0.00711462f $X=2.465 $Y=0.42 $X2=0 $Y2=0
cc_513 N_X_c_894_p N_VGND_c_921_n 0.00730901f $X=3.325 $Y=0.42 $X2=0 $Y2=0
cc_514 N_X_c_839_n N_A_877_47#_c_1013_n 0.00976354f $X=4.06 $Y=1.11 $X2=0 $Y2=0
cc_515 N_X_c_840_n N_A_877_47#_c_1013_n 0.0027916f $X=4.145 $Y=1.405 $X2=0 $Y2=0
cc_516 N_X_c_842_n N_A_877_47#_c_1013_n 0.0160744f $X=4.392 $Y=1.882 $X2=0 $Y2=0
cc_517 N_X_c_842_n N_A_877_47#_c_1015_n 0.00792768f $X=4.392 $Y=1.882 $X2=0
+ $Y2=0
cc_518 N_VGND_c_921_n N_A_877_47#_M1005_d 0.00536646f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_519 N_VGND_c_919_n N_A_877_47#_c_1036_n 0.0124525f $X=4.79 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_921_n N_A_877_47#_c_1036_n 0.00730901f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_M1016_s N_A_877_47#_c_1015_n 0.00412166f $X=4.815 $Y=0.235 $X2=0
+ $Y2=0
cc_522 N_VGND_c_913_n N_A_877_47#_c_1015_n 0.018043f $X=4.955 $Y=0.38 $X2=0
+ $Y2=0
cc_523 N_VGND_c_913_n N_A_1098_69#_c_1045_n 0.0206777f $X=4.955 $Y=0.38 $X2=0
+ $Y2=0
cc_524 N_VGND_c_920_n N_A_1098_69#_c_1046_n 0.0422287f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_921_n N_A_1098_69#_c_1046_n 0.0238173f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_913_n N_A_1098_69#_c_1047_n 0.0091975f $X=4.955 $Y=0.38 $X2=0
+ $Y2=0
cc_527 N_VGND_c_920_n N_A_1098_69#_c_1047_n 0.0208969f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_c_921_n N_A_1098_69#_c_1047_n 0.0114218f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_529 N_VGND_c_920_n N_A_1098_69#_c_1048_n 0.0608672f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_530 N_VGND_c_921_n N_A_1098_69#_c_1048_n 0.0339255f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_531 N_VGND_c_920_n N_A_1098_69#_c_1050_n 0.016488f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_921_n N_A_1098_69#_c_1050_n 0.00894187f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_533 N_A_877_47#_c_1014_n N_A_1098_69#_M1006_d 0.00797757f $X=5.915 $Y=1.09
+ $X2=-0.19 $Y2=-0.245
cc_534 N_A_877_47#_c_1014_n N_A_1098_69#_c_1045_n 0.0199559f $X=5.915 $Y=1.09
+ $X2=0 $Y2=0
cc_535 N_A_877_47#_M1006_s N_A_1098_69#_c_1046_n 0.00256188f $X=5.905 $Y=0.345
+ $X2=0 $Y2=0
cc_536 N_A_877_47#_c_1014_n N_A_1098_69#_c_1046_n 0.0036834f $X=5.915 $Y=1.09
+ $X2=0 $Y2=0
cc_537 N_A_877_47#_c_1044_p N_A_1098_69#_c_1046_n 0.0181205f $X=6.08 $Y=0.68
+ $X2=0 $Y2=0
