* File: sky130_fd_sc_lp__a311o_1.spice
* Created: Wed Sep  2 09:25:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311o_1.pex.spice"
.subckt sky130_fd_sc_lp__a311o_1  VNB VPB A3 A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_80_21#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2793 AS=0.2226 PD=1.505 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75003
+ A=0.126 P=1.98 MULT=1
MM1009 A_273_47# N_A3_M1009_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84 AD=0.126
+ AS=0.2793 PD=1.14 PS=1.505 NRD=13.56 NRS=0 M=1 R=5.6 SA=75001 SB=75002.2
+ A=0.126 P=1.98 MULT=1
MM1001 A_363_47# N_A2_M1001_g A_273_47# VNB NSHORT L=0.15 W=0.84 AD=0.126
+ AS=0.126 PD=1.14 PS=1.14 NRD=13.56 NRS=13.56 M=1 R=5.6 SA=75001.5 SB=75001.8
+ A=0.126 P=1.98 MULT=1
MM1002 N_A_80_21#_M1002_d N_A1_M1002_g A_363_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.189 AS=0.126 PD=1.29 PS=1.14 NRD=12.132 NRS=13.56 M=1 R=5.6 SA=75001.9
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_B1_M1007_g N_A_80_21#_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.189 PD=1.23 PS=1.29 NRD=5.712 NRS=12.132 M=1 R=5.6 SA=75002.5
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_A_80_21#_M1008_d N_C1_M1008_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75003
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.3339 PD=1.61 PS=3.05 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1005 N_A_259_367#_M1005_d N_A3_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2205 PD=1.54 PS=1.61 NRD=0 NRS=4.6886 M=1 R=8.4
+ SA=75000.7 SB=75002.3 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_259_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3969 AS=0.1764 PD=1.89 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1006 N_A_259_367#_M1006_d N_A1_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.3969 PD=1.65 PS=1.89 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 A_609_367# N_B1_M1011_g N_A_259_367#_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.2457 PD=1.47 PS=1.65 NRD=7.8012 NRS=6.2449 M=1 R=8.4 SA=75002.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_A_80_21#_M1010_d N_C1_M1010_g A_609_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75002.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a311o_1.pxi.spice"
*
.ends
*
*
