# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand2b_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nand2b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.185000 0.840000 1.515000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 1.075000 2.695000 1.245000 ;
        RECT 1.010000 1.245000 1.300000 1.515000 ;
        RECT 2.365000 1.245000 2.695000 1.515000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.970200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.230000 2.035000 3.275000 2.120000 ;
        RECT 1.230000 2.120000 2.320000 2.205000 ;
        RECT 1.230000 2.205000 1.460000 3.075000 ;
        RECT 1.630000 0.655000 1.960000 0.725000 ;
        RECT 1.630000 0.725000 3.275000 0.905000 ;
        RECT 1.970000 1.830000 3.275000 2.035000 ;
        RECT 2.130000 2.205000 2.320000 3.075000 ;
        RECT 2.875000 0.905000 3.275000 1.830000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.090000  0.685000 0.355000 1.015000 ;
      RECT 0.090000  1.015000 0.260000 1.695000 ;
      RECT 0.090000  1.695000 1.800000 1.865000 ;
      RECT 0.090000  1.865000 0.505000 2.210000 ;
      RECT 0.525000  0.085000 0.950000 0.905000 ;
      RECT 0.525000  0.905000 0.855000 0.995000 ;
      RECT 0.675000  2.035000 1.060000 3.245000 ;
      RECT 1.120000  0.255000 2.390000 0.485000 ;
      RECT 1.120000  0.485000 1.450000 0.905000 ;
      RECT 1.470000  1.415000 1.800000 1.695000 ;
      RECT 1.630000  2.375000 1.960000 3.245000 ;
      RECT 2.490000  2.290000 2.820000 3.245000 ;
      RECT 2.560000  0.085000 2.820000 0.555000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__nand2b_2
END LIBRARY
