* NGSPICE file created from sky130_fd_sc_lp__or4bb_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or4bb_m A B C_N D_N VGND VNB VPB VPWR X
M1000 X a_336_439# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.961e+11p ps=3.09e+06u
M1001 a_196_530# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=5.292e+11p ps=5.88e+06u
M1002 a_336_439# a_196_530# VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=0p ps=0u
M1003 VGND A a_336_439# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_419_439# a_196_530# a_336_439# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1005 a_491_439# a_27_530# a_419_439# VPB phighvt w=420000u l=150000u
+  ad=1.834e+11p pd=2.02e+06u as=0p ps=0u
M1006 a_196_530# D_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 a_593_485# B a_491_439# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 VPWR A a_593_485# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_530# a_336_439# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C_N a_27_530# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 VPWR C_N a_27_530# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 X a_336_439# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 a_336_439# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

