* File: sky130_fd_sc_lp__a21bo_lp.spice
* Created: Fri Aug 28 09:49:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21bo_lp.pex.spice"
.subckt sky130_fd_sc_lp__a21bo_lp  VNB VPB A2 A1 B1_N X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1_N	B1_N
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1007 A_114_55# N_A_84_29#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_84_29#_M1001_g A_114_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1008 A_272_55# N_A2_M1008_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_84_29#_M1009_d N_A1_M1009_g A_272_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 A_436_55# N_A_308_364#_M1000_g N_A_84_29#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_308_364#_M1012_g A_436_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1002 A_594_55# N_B1_N_M1002_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_308_364#_M1003_d N_B1_N_M1003_g A_594_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_84_29#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.145 AS=0.285 PD=1.29 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1011 N_A_252_409#_M1011_d N_A2_M1011_g N_VPWR_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.145 PD=1.28 PS=1.29 NRD=0 NRS=1.9503 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1006 N_A_84_29#_M1006_d N_A_308_364#_M1006_g N_A_252_409#_M1011_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_252_409#_M1010_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1005 N_A_308_364#_M1005_d N_B1_N_M1005_g N_VPWR_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a21bo_lp.pxi.spice"
*
.ends
*
*
