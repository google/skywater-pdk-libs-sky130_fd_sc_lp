* File: sky130_fd_sc_lp__iso1p_lp.pxi.spice
* Created: Wed Sep  2 09:58:22 2020
* 
x_PM_SKY130_FD_SC_LP__ISO1P_LP%A N_A_c_42_n N_A_M1007_g N_A_c_43_n N_A_M1005_g
+ N_A_c_45_n N_A_M1008_g A A PM_SKY130_FD_SC_LP__ISO1P_LP%A
x_PM_SKY130_FD_SC_LP__ISO1P_LP%SLEEP N_SLEEP_M1000_g N_SLEEP_M1001_g
+ N_SLEEP_M1009_g SLEEP N_SLEEP_c_83_n N_SLEEP_c_81_n
+ PM_SKY130_FD_SC_LP__ISO1P_LP%SLEEP
x_PM_SKY130_FD_SC_LP__ISO1P_LP%A_161_489# N_A_161_489#_M1008_d
+ N_A_161_489#_M1005_s N_A_161_489#_c_119_n N_A_161_489#_M1002_g
+ N_A_161_489#_M1003_g N_A_161_489#_c_120_n N_A_161_489#_M1004_g
+ N_A_161_489#_M1006_g N_A_161_489#_c_127_n N_A_161_489#_c_128_n
+ N_A_161_489#_c_129_n N_A_161_489#_c_121_n N_A_161_489#_c_122_n
+ N_A_161_489#_c_123_n N_A_161_489#_c_168_p N_A_161_489#_c_152_n
+ N_A_161_489#_c_124_n PM_SKY130_FD_SC_LP__ISO1P_LP%A_161_489#
x_PM_SKY130_FD_SC_LP__ISO1P_LP%KAPWR N_KAPWR_M1000_d KAPWR N_KAPWR_c_188_n
+ N_KAPWR_c_189_n PM_SKY130_FD_SC_LP__ISO1P_LP%KAPWR
x_PM_SKY130_FD_SC_LP__ISO1P_LP%X N_X_M1004_d N_X_M1006_d X X X X X N_X_c_216_n X
+ X X X X PM_SKY130_FD_SC_LP__ISO1P_LP%X
x_PM_SKY130_FD_SC_LP__ISO1P_LP%VGND N_VGND_M1007_s N_VGND_M1009_d N_VGND_c_229_n
+ N_VGND_c_230_n VGND N_VGND_c_231_n N_VGND_c_232_n N_VGND_c_233_n
+ N_VGND_c_234_n N_VGND_c_235_n N_VGND_c_236_n PM_SKY130_FD_SC_LP__ISO1P_LP%VGND
x_PM_SKY130_FD_SC_LP__ISO1P_LP%VPWR VPWR N_VPWR_c_266_n VPWR
+ PM_SKY130_FD_SC_LP__ISO1P_LP%VPWR
cc_1 VNB N_A_c_42_n 0.0174937f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.96
cc_2 VNB N_A_c_43_n 0.100216f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.645
cc_3 VNB N_A_M1005_g 4.92816e-19 $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.655
cc_4 VNB N_A_c_45_n 0.0141934f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.96
cc_5 VNB A 0.0235969f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_6 VNB N_SLEEP_M1000_g 5.47148e-19 $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.675
cc_7 VNB N_SLEEP_M1001_g 0.0301649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SLEEP_M1009_g 0.0292713f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_9 VNB N_SLEEP_c_81_n 0.054154f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=1.665
cc_10 VNB N_A_161_489#_c_119_n 0.0156843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_161_489#_c_120_n 0.020326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_161_489#_c_121_n 0.00525468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_161_489#_c_122_n 0.0206002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_161_489#_c_123_n 0.00879765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_161_489#_c_124_n 0.0632971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_X_c_216_n 0.0692912f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_17 VNB N_VGND_c_229_n 0.0316526f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.675
cc_18 VNB N_VGND_c_230_n 0.0116388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_231_n 0.0167814f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.48
cc_20 VNB N_VGND_c_232_n 0.0383522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_233_n 0.0319968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_234_n 0.252491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_235_n 0.00577043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_236_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB VPWR 0.143779f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.96
cc_26 VPB N_A_M1005_g 0.0641941f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=2.655
cc_27 VPB A 0.0161359f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_28 VPB N_SLEEP_M1000_g 0.0658945f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.675
cc_29 VPB N_SLEEP_c_83_n 0.00582997f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=1.48
cc_30 VPB N_A_161_489#_M1003_g 0.0227029f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_31 VPB N_A_161_489#_M1006_g 0.0203893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_161_489#_c_127_n 0.0241388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_A_161_489#_c_128_n 0.0196027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_A_161_489#_c_129_n 0.00984468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_161_489#_c_124_n 0.00293676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_KAPWR_c_188_n 0.054445f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_37 VPB N_KAPWR_c_189_n 0.0142089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_X_c_216_n 0.0621984f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.295
cc_39 VPB VPWR 0.0582378f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.96
cc_40 VPB N_VPWR_c_266_n 0.0977898f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=0.96
cc_41 N_A_M1005_g N_SLEEP_M1000_g 0.0532446f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_42 N_A_c_43_n N_SLEEP_M1001_g 0.00938378f $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_43 N_A_c_45_n N_SLEEP_M1001_g 0.0171659f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_44 A N_SLEEP_M1001_g 4.46117e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_45 N_A_c_43_n N_SLEEP_c_83_n 4.97555e-19 $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_46 A N_SLEEP_c_83_n 0.0282905f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_47 N_A_c_43_n N_SLEEP_c_81_n 0.0532446f $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_48 A N_SLEEP_c_81_n 0.00161646f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_49 N_A_M1005_g N_A_161_489#_c_127_n 0.0176365f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_50 N_A_M1005_g N_A_161_489#_c_128_n 0.00816541f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_51 A N_A_161_489#_c_128_n 0.00780975f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_52 N_A_c_43_n N_A_161_489#_c_129_n 0.00183499f $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_53 N_A_M1005_g N_A_161_489#_c_129_n 0.00423371f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_54 A N_A_161_489#_c_129_n 0.0260029f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_55 N_A_c_45_n N_A_161_489#_c_121_n 0.00377352f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_56 N_A_c_43_n N_A_161_489#_c_123_n 0.00533946f $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_57 A N_A_161_489#_c_123_n 8.46245e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_58 N_A_M1005_g N_KAPWR_c_188_n 0.00440736f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_59 N_A_M1005_g N_KAPWR_c_189_n 0.00267943f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_60 N_A_c_42_n N_VGND_c_229_n 0.0124306f $X=0.81 $Y=0.96 $X2=0 $Y2=0
cc_61 N_A_c_43_n N_VGND_c_229_n 8.10401e-19 $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_62 N_A_c_45_n N_VGND_c_229_n 0.0016536f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_63 A N_VGND_c_229_n 0.00995469f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_64 N_A_c_42_n N_VGND_c_232_n 0.00424179f $X=0.81 $Y=0.96 $X2=0 $Y2=0
cc_65 N_A_c_45_n N_VGND_c_232_n 0.00510437f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_66 N_A_c_42_n N_VGND_c_234_n 0.0043341f $X=0.81 $Y=0.96 $X2=0 $Y2=0
cc_67 N_A_c_45_n N_VGND_c_234_n 0.00515964f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_68 N_A_M1005_g VPWR 0.00310524f $X=1.15 $Y=2.655 $X2=-0.19 $Y2=-0.245
cc_69 N_A_M1005_g N_VPWR_c_266_n 0.00489592f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_70 N_SLEEP_M1009_g N_A_161_489#_c_119_n 0.0280814f $X=1.96 $Y=0.675 $X2=0
+ $Y2=0
cc_71 N_SLEEP_M1000_g N_A_161_489#_c_127_n 0.00236308f $X=1.51 $Y=2.655 $X2=0
+ $Y2=0
cc_72 N_SLEEP_M1000_g N_A_161_489#_c_128_n 0.013341f $X=1.51 $Y=2.655 $X2=0
+ $Y2=0
cc_73 N_SLEEP_c_83_n N_A_161_489#_c_128_n 0.0460501f $X=1.94 $Y=1.48 $X2=0 $Y2=0
cc_74 N_SLEEP_c_81_n N_A_161_489#_c_128_n 0.0027233f $X=1.96 $Y=1.48 $X2=0 $Y2=0
cc_75 N_SLEEP_M1001_g N_A_161_489#_c_121_n 0.00370726f $X=1.6 $Y=0.675 $X2=0
+ $Y2=0
cc_76 N_SLEEP_M1001_g N_A_161_489#_c_122_n 0.0140103f $X=1.6 $Y=0.675 $X2=0
+ $Y2=0
cc_77 N_SLEEP_M1009_g N_A_161_489#_c_122_n 0.01362f $X=1.96 $Y=0.675 $X2=0 $Y2=0
cc_78 N_SLEEP_c_83_n N_A_161_489#_c_122_n 0.0459044f $X=1.94 $Y=1.48 $X2=0 $Y2=0
cc_79 N_SLEEP_c_81_n N_A_161_489#_c_122_n 0.00330876f $X=1.96 $Y=1.48 $X2=0
+ $Y2=0
cc_80 N_SLEEP_c_83_n N_A_161_489#_c_123_n 0.00463681f $X=1.94 $Y=1.48 $X2=0
+ $Y2=0
cc_81 N_SLEEP_c_81_n N_A_161_489#_c_123_n 0.00158276f $X=1.96 $Y=1.48 $X2=0
+ $Y2=0
cc_82 N_SLEEP_M1009_g N_A_161_489#_c_152_n 7.7944e-19 $X=1.96 $Y=0.675 $X2=0
+ $Y2=0
cc_83 N_SLEEP_c_83_n N_A_161_489#_c_152_n 0.0241847f $X=1.94 $Y=1.48 $X2=0 $Y2=0
cc_84 N_SLEEP_c_81_n N_A_161_489#_c_152_n 0.0013583f $X=1.96 $Y=1.48 $X2=0 $Y2=0
cc_85 N_SLEEP_c_83_n N_A_161_489#_c_124_n 0.00338649f $X=1.94 $Y=1.48 $X2=0
+ $Y2=0
cc_86 N_SLEEP_c_81_n N_A_161_489#_c_124_n 0.0223211f $X=1.96 $Y=1.48 $X2=0 $Y2=0
cc_87 N_SLEEP_M1000_g N_KAPWR_c_188_n 0.00365957f $X=1.51 $Y=2.655 $X2=0 $Y2=0
cc_88 N_SLEEP_M1000_g N_KAPWR_c_189_n 0.0194223f $X=1.51 $Y=2.655 $X2=0 $Y2=0
cc_89 N_SLEEP_M1001_g N_VGND_c_230_n 0.00165191f $X=1.6 $Y=0.675 $X2=0 $Y2=0
cc_90 N_SLEEP_M1009_g N_VGND_c_230_n 0.0111446f $X=1.96 $Y=0.675 $X2=0 $Y2=0
cc_91 N_SLEEP_M1001_g N_VGND_c_232_n 0.00510437f $X=1.6 $Y=0.675 $X2=0 $Y2=0
cc_92 N_SLEEP_M1009_g N_VGND_c_232_n 0.00424179f $X=1.96 $Y=0.675 $X2=0 $Y2=0
cc_93 N_SLEEP_M1001_g N_VGND_c_234_n 0.00515964f $X=1.6 $Y=0.675 $X2=0 $Y2=0
cc_94 N_SLEEP_M1009_g N_VGND_c_234_n 0.0043341f $X=1.96 $Y=0.675 $X2=0 $Y2=0
cc_95 N_SLEEP_M1000_g VPWR 0.0025877f $X=1.51 $Y=2.655 $X2=-0.19 $Y2=-0.245
cc_96 N_SLEEP_M1000_g N_VPWR_c_266_n 0.00438266f $X=1.51 $Y=2.655 $X2=0 $Y2=0
cc_97 N_A_161_489#_c_128_n N_KAPWR_M1000_d 0.00935341f $X=2.35 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_161_489#_M1003_g N_KAPWR_c_188_n 0.00320298f $X=2.39 $Y=2.465 $X2=0
+ $Y2=0
cc_99 N_A_161_489#_M1006_g N_KAPWR_c_188_n 0.009404f $X=2.75 $Y=2.465 $X2=0
+ $Y2=0
cc_100 N_A_161_489#_c_127_n N_KAPWR_c_188_n 0.0357314f $X=0.935 $Y=2.655 $X2=0
+ $Y2=0
cc_101 N_A_161_489#_c_128_n N_KAPWR_c_188_n 0.0282029f $X=2.35 $Y=2.04 $X2=0
+ $Y2=0
cc_102 N_A_161_489#_M1003_g N_KAPWR_c_189_n 0.018678f $X=2.39 $Y=2.465 $X2=0
+ $Y2=0
cc_103 N_A_161_489#_M1006_g N_KAPWR_c_189_n 0.00245424f $X=2.75 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_A_161_489#_c_127_n N_KAPWR_c_189_n 0.015825f $X=0.935 $Y=2.655 $X2=0
+ $Y2=0
cc_105 N_A_161_489#_c_128_n N_KAPWR_c_189_n 0.0599322f $X=2.35 $Y=2.04 $X2=0
+ $Y2=0
cc_106 N_A_161_489#_c_128_n A_493_367# 0.00216169f $X=2.35 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_107 N_A_161_489#_c_120_n N_X_c_216_n 0.0332622f $X=2.75 $Y=1.005 $X2=0 $Y2=0
cc_108 N_A_161_489#_c_168_p N_X_c_216_n 0.0145272f $X=2.517 $Y=1.18 $X2=0 $Y2=0
cc_109 N_A_161_489#_c_152_n N_X_c_216_n 0.0572537f $X=2.517 $Y=1.955 $X2=0 $Y2=0
cc_110 N_A_161_489#_c_121_n N_VGND_c_229_n 0.00635101f $X=1.385 $Y=0.72 $X2=0
+ $Y2=0
cc_111 N_A_161_489#_c_119_n N_VGND_c_230_n 0.0111236f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_112 N_A_161_489#_c_120_n N_VGND_c_230_n 0.00170417f $X=2.75 $Y=1.005 $X2=0
+ $Y2=0
cc_113 N_A_161_489#_c_121_n N_VGND_c_230_n 0.00643814f $X=1.385 $Y=0.72 $X2=0
+ $Y2=0
cc_114 N_A_161_489#_c_122_n N_VGND_c_230_n 0.0216087f $X=2.35 $Y=1.095 $X2=0
+ $Y2=0
cc_115 N_A_161_489#_c_121_n N_VGND_c_232_n 0.00680149f $X=1.385 $Y=0.72 $X2=0
+ $Y2=0
cc_116 N_A_161_489#_c_119_n N_VGND_c_233_n 0.00424179f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_117 N_A_161_489#_c_120_n N_VGND_c_233_n 0.00510437f $X=2.75 $Y=1.005 $X2=0
+ $Y2=0
cc_118 N_A_161_489#_c_119_n N_VGND_c_234_n 0.0043341f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_119 N_A_161_489#_c_120_n N_VGND_c_234_n 0.00515964f $X=2.75 $Y=1.005 $X2=0
+ $Y2=0
cc_120 N_A_161_489#_c_121_n N_VGND_c_234_n 0.00725225f $X=1.385 $Y=0.72 $X2=0
+ $Y2=0
cc_121 N_A_161_489#_M1003_g VPWR 0.00637747f $X=2.39 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_161_489#_M1006_g VPWR 0.00633226f $X=2.75 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_161_489#_c_127_n VPWR 0.00145921f $X=0.935 $Y=2.655 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_161_489#_M1003_g N_VPWR_c_266_n 0.00509549f $X=2.39 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_161_489#_M1006_g N_VPWR_c_266_n 0.00585385f $X=2.75 $Y=2.465 $X2=0
+ $Y2=0
cc_126 N_A_161_489#_c_127_n N_VPWR_c_266_n 0.00840241f $X=0.935 $Y=2.655 $X2=0
+ $Y2=0
cc_127 A_245_489# N_KAPWR_c_188_n 0.00269277f $X=1.225 $Y=2.445 $X2=2.155
+ $Y2=2.775
cc_128 N_KAPWR_c_188_n A_493_367# 0.00411194f $X=2.155 $Y=2.775 $X2=-0.19
+ $Y2=1.655
cc_129 N_KAPWR_c_188_n N_X_M1006_d 0.00127496f $X=2.155 $Y=2.775 $X2=0 $Y2=0
cc_130 N_KAPWR_c_188_n N_X_c_216_n 0.0481095f $X=2.155 $Y=2.775 $X2=0 $Y2=0
cc_131 N_KAPWR_c_189_n N_X_c_216_n 0.0129498f $X=2.175 $Y=2.38 $X2=0 $Y2=0
cc_132 N_KAPWR_M1000_d VPWR 0.00121531f $X=1.585 $Y=2.445 $X2=-0.19 $Y2=1.655
cc_133 N_KAPWR_c_188_n VPWR 0.294444f $X=2.155 $Y=2.775 $X2=-0.19 $Y2=1.655
cc_134 N_KAPWR_c_189_n VPWR 0.00867316f $X=2.175 $Y=2.38 $X2=-0.19 $Y2=1.655
cc_135 N_KAPWR_c_188_n N_VPWR_c_266_n 0.0106586f $X=2.155 $Y=2.775 $X2=0 $Y2=0
cc_136 N_KAPWR_c_189_n N_VPWR_c_266_n 0.0548023f $X=2.175 $Y=2.38 $X2=0 $Y2=0
cc_137 A_493_367# VPWR 0.00190157f $X=2.465 $Y=1.835 $X2=1.245 $Y2=0.465
cc_138 N_X_c_216_n N_VGND_c_233_n 0.0121076f $X=2.965 $Y=0.72 $X2=0 $Y2=0
cc_139 N_X_c_216_n N_VGND_c_234_n 0.0143287f $X=2.965 $Y=0.72 $X2=0 $Y2=0
cc_140 N_X_M1006_d VPWR 0.00135204f $X=2.825 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_141 N_X_c_216_n VPWR 0.00454457f $X=2.965 $Y=0.72 $X2=-0.19 $Y2=-0.245
cc_142 N_X_c_216_n N_VPWR_c_266_n 0.0287379f $X=2.965 $Y=0.72 $X2=0 $Y2=0
