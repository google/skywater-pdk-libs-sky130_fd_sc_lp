* File: sky130_fd_sc_lp__or3b_4.pex.spice
* Created: Fri Aug 28 11:24:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3B_4%C_N 3 6 8 9 10 11 12 19 21
r30 19 22 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.697 $Y=1.36
+ $X2=0.697 $Y2=1.525
r31 19 21 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.697 $Y=1.36
+ $X2=0.697 $Y2=1.195
r32 11 12 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.035
r33 10 11 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=1.295
+ $X2=0.73 $Y2=1.665
r34 10 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.36 $X2=0.72 $Y2=1.36
r35 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=0.925
+ $X2=0.73 $Y2=1.295
r36 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=0.555 $X2=0.73
+ $Y2=0.925
r37 6 22 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.585 $Y=2.045
+ $X2=0.585 $Y2=1.525
r38 3 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.585 $Y=0.875
+ $X2=0.585 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_4%A_253_23# 1 2 3 12 16 20 24 28 32 36 40 42 51
+ 52 53 56 58 62 68 70 71 73 75 76 85
c138 68 0 3.91013e-20 $X=3.362 $Y=1.09
r139 85 86 5.19077 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=2.63 $Y=1.51
+ $X2=2.665 $Y2=1.51
r140 82 83 5.19077 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=2.2 $Y=1.51
+ $X2=2.235 $Y2=1.51
r141 81 82 58.5815 $w=3.25e-07 $l=3.95e-07 $layer=POLY_cond $X=1.805 $Y=1.51
+ $X2=2.2 $Y2=1.51
r142 80 81 5.19077 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=1.77 $Y=1.51
+ $X2=1.805 $Y2=1.51
r143 77 78 5.19077 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=1.34 $Y=1.51
+ $X2=1.375 $Y2=1.51
r144 75 76 8.83418 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=1.98
+ $X2=4.485 $Y2=1.815
r145 70 71 3.69584 $w=5.53e-07 $l=1.5e-07 $layer=LI1_cond $X=4.432 $Y=2.91
+ $X2=4.432 $Y2=2.76
r146 66 73 2.68319 $w=3.57e-07 $l=2.16365e-07 $layer=LI1_cond $X=4.62 $Y=1.175
+ $X2=4.442 $Y2=1.09
r147 66 76 39.4343 $w=1.78e-07 $l=6.4e-07 $layer=LI1_cond $X=4.62 $Y=1.175
+ $X2=4.62 $Y2=1.815
r148 64 75 1.59477 $w=4.48e-07 $l=6e-08 $layer=LI1_cond $X=4.485 $Y=2.04
+ $X2=4.485 $Y2=1.98
r149 64 71 19.1373 $w=4.48e-07 $l=7.2e-07 $layer=LI1_cond $X=4.485 $Y=2.04
+ $X2=4.485 $Y2=2.76
r150 60 73 2.68319 $w=3.57e-07 $l=8.5e-08 $layer=LI1_cond $X=4.442 $Y=1.005
+ $X2=4.442 $Y2=1.09
r151 60 62 13.0786 $w=5.33e-07 $l=5.85e-07 $layer=LI1_cond $X=4.442 $Y=1.005
+ $X2=4.442 $Y2=0.42
r152 59 68 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.505 $Y=1.09
+ $X2=3.362 $Y2=1.09
r153 58 73 4.11427 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=4.175 $Y=1.09
+ $X2=4.442 $Y2=1.09
r154 58 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.175 $Y=1.09
+ $X2=3.505 $Y2=1.09
r155 54 68 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.362 $Y=1.005
+ $X2=3.362 $Y2=1.09
r156 54 56 23.6554 $w=2.83e-07 $l=5.85e-07 $layer=LI1_cond $X=3.362 $Y=1.005
+ $X2=3.362 $Y2=0.42
r157 52 68 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.22 $Y=1.09
+ $X2=3.362 $Y2=1.09
r158 52 53 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.22 $Y=1.09
+ $X2=2.85 $Y2=1.09
r159 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.765 $Y=1.175
+ $X2=2.85 $Y2=1.09
r160 50 51 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.765 $Y=1.175
+ $X2=2.765 $Y2=1.415
r161 49 85 13.3477 $w=3.25e-07 $l=9e-08 $layer=POLY_cond $X=2.54 $Y=1.51
+ $X2=2.63 $Y2=1.51
r162 49 83 45.2338 $w=3.25e-07 $l=3.05e-07 $layer=POLY_cond $X=2.54 $Y=1.51
+ $X2=2.235 $Y2=1.51
r163 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.54
+ $Y=1.51 $X2=2.54 $Y2=1.51
r164 45 80 37.0769 $w=3.25e-07 $l=2.5e-07 $layer=POLY_cond $X=1.52 $Y=1.51
+ $X2=1.77 $Y2=1.51
r165 45 78 21.5046 $w=3.25e-07 $l=1.45e-07 $layer=POLY_cond $X=1.52 $Y=1.51
+ $X2=1.375 $Y2=1.51
r166 44 48 51.1083 $w=2.28e-07 $l=1.02e-06 $layer=LI1_cond $X=1.52 $Y=1.53
+ $X2=2.54 $Y2=1.53
r167 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.52
+ $Y=1.51 $X2=1.52 $Y2=1.51
r168 42 51 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.68 $Y=1.53
+ $X2=2.765 $Y2=1.415
r169 42 48 7.01487 $w=2.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.68 $Y=1.53
+ $X2=2.54 $Y2=1.53
r170 38 86 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=1.675
+ $X2=2.665 $Y2=1.51
r171 38 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.665 $Y=1.675
+ $X2=2.665 $Y2=2.465
r172 34 85 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.63 $Y=1.345
+ $X2=2.63 $Y2=1.51
r173 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.63 $Y=1.345
+ $X2=2.63 $Y2=0.665
r174 30 83 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.675
+ $X2=2.235 $Y2=1.51
r175 30 32 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.235 $Y=1.675
+ $X2=2.235 $Y2=2.465
r176 26 82 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.345 $X2=2.2
+ $Y2=1.51
r177 26 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.2 $Y=1.345
+ $X2=2.2 $Y2=0.665
r178 22 81 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.675
+ $X2=1.805 $Y2=1.51
r179 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.805 $Y=1.675
+ $X2=1.805 $Y2=2.465
r180 18 80 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.345
+ $X2=1.77 $Y2=1.51
r181 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.77 $Y=1.345
+ $X2=1.77 $Y2=0.665
r182 14 78 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.675
+ $X2=1.375 $Y2=1.51
r183 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.375 $Y=1.675
+ $X2=1.375 $Y2=2.465
r184 10 77 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.345
+ $X2=1.34 $Y2=1.51
r185 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.34 $Y=1.345
+ $X2=1.34 $Y2=0.665
r186 3 75 300 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=2 $X=4.18
+ $Y=1.835 $X2=4.345 $Y2=1.98
r187 3 70 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.835 $X2=4.32 $Y2=2.91
r188 2 62 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=4.18
+ $Y=0.245 $X2=4.32 $Y2=0.42
r189 1 56 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.215
+ $Y=0.245 $X2=3.355 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_4%A 3 7 9 10 14 15
r39 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.51
+ $X2=3.115 $Y2=1.675
r40 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.51
+ $X2=3.115 $Y2=1.345
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.115
+ $Y=1.51 $X2=3.115 $Y2=1.51
r42 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.147 $Y=1.665
+ $X2=3.147 $Y2=2.035
r43 9 15 7.00505 $w=2.53e-07 $l=1.55e-07 $layer=LI1_cond $X=3.147 $Y=1.665
+ $X2=3.147 $Y2=1.51
r44 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.205 $Y=2.465
+ $X2=3.205 $Y2=1.675
r45 3 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.14 $Y=0.665
+ $X2=3.14 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_4%B 3 7 9 10 14 15
c38 14 0 2.2542e-19 $X=3.655 $Y=1.51
r39 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.51
+ $X2=3.655 $Y2=1.675
r40 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.51
+ $X2=3.655 $Y2=1.345
r41 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=1.51 $X2=3.655 $Y2=1.51
r42 9 10 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=3.592 $Y=1.665
+ $X2=3.592 $Y2=2.035
r43 9 15 6.05521 $w=2.93e-07 $l=1.55e-07 $layer=LI1_cond $X=3.592 $Y=1.665
+ $X2=3.592 $Y2=1.51
r44 7 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.57 $Y=0.665
+ $X2=3.57 $Y2=1.345
r45 3 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.565 $Y=2.465
+ $X2=3.565 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_4%A_49_133# 1 2 9 13 17 21 22 24 28 29
c75 24 0 1.86319e-19 $X=4.005 $Y=2.315
r76 29 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.195 $Y=1.51
+ $X2=4.195 $Y2=1.675
r77 29 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.195 $Y=1.51
+ $X2=4.195 $Y2=1.345
r78 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.195
+ $Y=1.51 $X2=4.195 $Y2=1.51
r79 25 28 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=4.005 $Y=1.495
+ $X2=4.195 $Y2=1.495
r80 23 25 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.005 $Y=1.645
+ $X2=4.005 $Y2=1.495
r81 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.005 $Y=1.645
+ $X2=4.005 $Y2=2.315
r82 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=2.4
+ $X2=4.005 $Y2=2.315
r83 21 22 226.059 $w=1.68e-07 $l=3.465e-06 $layer=LI1_cond $X=3.92 $Y=2.4
+ $X2=0.455 $Y2=2.4
r84 17 20 53.9343 $w=2.48e-07 $l=1.17e-06 $layer=LI1_cond $X=0.33 $Y=0.875
+ $X2=0.33 $Y2=2.045
r85 15 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.33 $Y=2.315
+ $X2=0.455 $Y2=2.4
r86 15 20 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=0.33 $Y=2.315
+ $X2=0.33 $Y2=2.045
r87 13 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.105 $Y=2.465
+ $X2=4.105 $Y2=1.675
r88 9 32 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.105 $Y=0.665
+ $X2=4.105 $Y2=1.345
r89 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.045
r90 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.665 $X2=0.37 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_4%VPWR 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r54 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 44 47 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 43 46 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 41 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r60 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 38 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.16 $Y2=3.33
r64 35 37 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 33 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.16 $Y2=3.33
r68 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 28 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r70 28 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 26 40 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.64 $Y2=3.33
r72 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.935 $Y2=3.33
r73 25 43 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.1 $Y=3.33 $X2=3.12
+ $Y2=3.33
r74 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.1 $Y=3.33
+ $X2=2.935 $Y2=3.33
r75 23 37 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=3.33
+ $X2=2.02 $Y2=3.33
r77 22 40 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=2.02 $Y2=3.33
r79 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=3.245
+ $X2=2.935 $Y2=3.33
r80 18 20 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.935 $Y=3.245
+ $X2=2.935 $Y2=2.78
r81 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=3.245
+ $X2=2.02 $Y2=3.33
r82 14 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.02 $Y=3.245
+ $X2=2.02 $Y2=2.78
r83 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=3.245
+ $X2=1.16 $Y2=3.33
r84 10 12 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.16 $Y=3.245
+ $X2=1.16 $Y2=2.78
r85 3 20 600 $w=1.7e-07 $l=1.03793e-06 $layer=licon1_PDIFF $count=1 $X=2.74
+ $Y=1.835 $X2=2.935 $Y2=2.78
r86 2 16 600 $w=1.7e-07 $l=1.01258e-06 $layer=licon1_PDIFF $count=1 $X=1.88
+ $Y=1.835 $X2=2.02 $Y2=2.78
r87 1 12 600 $w=1.7e-07 $l=1.16856e-06 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=1.16 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_4%X 1 2 3 4 14 15 16 19 21 25 27 28 29 30 31 39
r56 37 39 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.185 $Y=1.98
+ $X2=1.2 $Y2=1.98
r57 31 48 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.64 $Y=1.98
+ $X2=2.45 $Y2=1.98
r58 30 48 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.16 $Y=1.98
+ $X2=2.45 $Y2=1.98
r59 29 30 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.98
+ $X2=2.16 $Y2=1.98
r60 29 42 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.68 $Y=1.98 $X2=1.59
+ $Y2=1.98
r61 28 37 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.095 $Y=1.98 $X2=1.185
+ $Y2=1.98
r62 28 42 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.235 $Y=1.98
+ $X2=1.59 $Y2=1.98
r63 28 39 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.235 $Y=1.98
+ $X2=1.2 $Y2=1.98
r64 23 25 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=2.415 $Y=1.075
+ $X2=2.415 $Y2=0.42
r65 22 27 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.65 $Y=1.16 $X2=1.54
+ $Y2=1.16
r66 21 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.32 $Y=1.16
+ $X2=2.415 $Y2=1.075
r67 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.32 $Y=1.16
+ $X2=1.65 $Y2=1.16
r68 17 27 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=1.075
+ $X2=1.54 $Y2=1.16
r69 17 19 34.3114 $w=2.18e-07 $l=6.55e-07 $layer=LI1_cond $X=1.54 $Y=1.075
+ $X2=1.54 $Y2=0.42
r70 15 27 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.43 $Y=1.16 $X2=1.54
+ $Y2=1.16
r71 15 16 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.43 $Y=1.16
+ $X2=1.185 $Y2=1.16
r72 14 28 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=1.815
+ $X2=1.095 $Y2=1.98
r73 13 16 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.095 $Y=1.245
+ $X2=1.185 $Y2=1.16
r74 13 14 35.1212 $w=1.78e-07 $l=5.7e-07 $layer=LI1_cond $X=1.095 $Y=1.245
+ $X2=1.095 $Y2=1.815
r75 4 48 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.31
+ $Y=1.835 $X2=2.45 $Y2=1.98
r76 3 42 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.835 $X2=1.59 $Y2=1.98
r77 2 25 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.275
+ $Y=0.245 $X2=2.415 $Y2=0.42
r78 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.415
+ $Y=0.245 $X2=1.555 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37 39
+ 40 41 57 58
r70 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r71 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r72 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r73 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r74 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r75 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r76 45 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r77 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r78 41 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r79 41 49 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r80 39 54 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.6
+ $Y2=0
r81 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=0 $X2=3.84
+ $Y2=0
r82 38 57 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.56
+ $Y2=0
r83 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=3.84
+ $Y2=0
r84 36 51 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.64
+ $Y2=0
r85 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.885
+ $Y2=0
r86 35 54 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=3.6
+ $Y2=0
r87 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=0 $X2=2.885
+ $Y2=0
r88 33 48 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=1.68
+ $Y2=0
r89 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=1.985
+ $Y2=0
r90 32 51 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.64
+ $Y2=0
r91 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=1.985
+ $Y2=0
r92 30 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.72
+ $Y2=0
r93 30 31 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.132
+ $Y2=0
r94 29 48 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.68
+ $Y2=0
r95 29 31 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.132
+ $Y2=0
r96 25 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=0.085
+ $X2=3.84 $Y2=0
r97 25 27 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.84 $Y=0.085
+ $X2=3.84 $Y2=0.37
r98 21 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=0.085
+ $X2=2.885 $Y2=0
r99 21 23 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.885 $Y=0.085
+ $X2=2.885 $Y2=0.37
r100 17 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.085
+ $X2=1.985 $Y2=0
r101 17 19 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0.085
+ $X2=1.985 $Y2=0.39
r102 13 31 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.132 $Y=0.085
+ $X2=1.132 $Y2=0
r103 13 15 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=1.132 $Y=0.085
+ $X2=1.132 $Y2=0.39
r104 4 27 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=3.645
+ $Y=0.245 $X2=3.84 $Y2=0.37
r105 3 23 91 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=2 $X=2.705
+ $Y=0.245 $X2=2.885 $Y2=0.37
r106 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.845
+ $Y=0.245 $X2=1.985 $Y2=0.39
r107 1 15 91 $w=1.7e-07 $l=5.866e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.665 $X2=1.125 $Y2=0.39
.ends

