* File: sky130_fd_sc_lp__o211ai_lp.pxi.spice
* Created: Fri Aug 28 11:03:17 2020
* 
x_PM_SKY130_FD_SC_LP__O211AI_LP%A1 N_A1_M1007_g N_A1_M1004_g N_A1_c_61_n
+ N_A1_c_66_n A1 A1 N_A1_c_63_n PM_SKY130_FD_SC_LP__O211AI_LP%A1
x_PM_SKY130_FD_SC_LP__O211AI_LP%A2 N_A2_M1003_g N_A2_M1005_g N_A2_c_93_n
+ N_A2_c_98_n A2 A2 N_A2_c_95_n PM_SKY130_FD_SC_LP__O211AI_LP%A2
x_PM_SKY130_FD_SC_LP__O211AI_LP%B1 N_B1_M1001_g N_B1_M1006_g N_B1_c_134_n
+ N_B1_c_139_n B1 B1 N_B1_c_136_n PM_SKY130_FD_SC_LP__O211AI_LP%B1
x_PM_SKY130_FD_SC_LP__O211AI_LP%C1 N_C1_c_176_n N_C1_M1002_g N_C1_M1000_g
+ N_C1_c_177_n N_C1_c_178_n N_C1_c_179_n N_C1_c_180_n C1 C1 N_C1_c_182_n
+ PM_SKY130_FD_SC_LP__O211AI_LP%C1
x_PM_SKY130_FD_SC_LP__O211AI_LP%VPWR N_VPWR_M1007_s N_VPWR_M1006_d
+ N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n N_VPWR_c_225_n N_VPWR_c_226_n
+ VPWR N_VPWR_c_227_n N_VPWR_c_221_n PM_SKY130_FD_SC_LP__O211AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O211AI_LP%Y N_Y_M1002_d N_Y_M1003_d N_Y_M1000_d
+ N_Y_c_255_n N_Y_c_256_n N_Y_c_257_n N_Y_c_258_n N_Y_c_252_n N_Y_c_253_n
+ N_Y_c_260_n Y Y N_Y_c_254_n PM_SKY130_FD_SC_LP__O211AI_LP%Y
x_PM_SKY130_FD_SC_LP__O211AI_LP%A_38_57# N_A_38_57#_M1004_s N_A_38_57#_M1005_d
+ N_A_38_57#_c_302_n N_A_38_57#_c_303_n N_A_38_57#_c_304_n N_A_38_57#_c_305_n
+ PM_SKY130_FD_SC_LP__O211AI_LP%A_38_57#
x_PM_SKY130_FD_SC_LP__O211AI_LP%VGND N_VGND_M1004_d N_VGND_c_333_n VGND
+ N_VGND_c_334_n N_VGND_c_335_n N_VGND_c_336_n
+ PM_SKY130_FD_SC_LP__O211AI_LP%VGND
cc_1 VNB N_A1_M1004_g 0.048725f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.495
cc_2 VNB N_A1_c_61_n 0.0267375f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.69
cc_3 VNB A1 0.0237208f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_63_n 0.0189674f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.335
cc_5 VNB N_A2_M1005_g 0.0367589f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.495
cc_6 VNB N_A2_c_93_n 0.0213176f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.69
cc_7 VNB A2 0.00529762f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.84
cc_8 VNB N_A2_c_95_n 0.016135f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.335
cc_9 VNB N_B1_M1001_g 0.0351404f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.545
cc_10 VNB N_B1_c_134_n 0.0225403f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.69
cc_11 VNB B1 0.00727708f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.84
cc_12 VNB N_B1_c_136_n 0.0167676f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.335
cc_13 VNB N_C1_c_176_n 0.0180782f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.84
cc_14 VNB N_C1_c_177_n 0.0257324f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.69
cc_15 VNB N_C1_c_178_n 0.0116789f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_C1_c_179_n 0.0240236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C1_c_180_n 0.00284303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB C1 0.00655194f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.335
cc_19 VNB N_C1_c_182_n 0.0172288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_221_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_252_n 0.0228865f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.335
cc_22 VNB N_Y_c_253_n 0.0455834f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.665
cc_23 VNB N_Y_c_254_n 0.0191225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_38_57#_c_302_n 0.0238089f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.335
cc_25 VNB N_A_38_57#_c_303_n 0.0246724f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.69
cc_26 VNB N_A_38_57#_c_304_n 0.010032f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.69
cc_27 VNB N_A_38_57#_c_305_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_VGND_c_333_n 0.00712794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_334_n 0.0517616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_335_n 0.193123f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.335
cc_31 VNB N_VGND_c_336_n 0.0271037f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.295
cc_32 VPB N_A1_M1007_g 0.0360071f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_33 VPB N_A1_c_61_n 0.00284976f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.69
cc_34 VPB N_A1_c_66_n 0.0204975f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.84
cc_35 VPB A1 0.0103901f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_36 VPB N_A2_M1003_g 0.0292916f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_37 VPB N_A2_c_93_n 0.0012697f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.69
cc_38 VPB N_A2_c_98_n 0.012962f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.69
cc_39 VPB A2 0.00294695f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.84
cc_40 VPB N_B1_M1006_g 0.0294035f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.495
cc_41 VPB N_B1_c_134_n 0.00134252f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.69
cc_42 VPB N_B1_c_139_n 0.0139235f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.69
cc_43 VPB B1 7.56276e-19 $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.84
cc_44 VPB N_C1_M1000_g 0.03758f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_C1_c_180_n 0.0111394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB C1 0.00188859f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.335
cc_47 VPB N_VPWR_c_222_n 0.0117329f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.495
cc_48 VPB N_VPWR_c_223_n 0.0466159f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.335
cc_49 VPB N_VPWR_c_224_n 0.00416546f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_50 VPB N_VPWR_c_225_n 0.0355708f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.335
cc_51 VPB N_VPWR_c_226_n 0.00544869f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.335
cc_52 VPB N_VPWR_c_227_n 0.0242841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_221_n 0.0627537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_Y_c_255_n 0.00252852f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_55 VPB N_Y_c_256_n 0.00830824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_Y_c_257_n 0.00871349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_258_n 0.0422771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_Y_c_253_n 0.0180321f $X=-0.19 $Y=1.655 $X2=0.375 $Y2=1.665
cc_59 VPB N_Y_c_260_n 0.0163354f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 N_A1_M1007_g N_A2_M1003_g 0.041607f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_61 N_A1_M1004_g N_A2_M1005_g 0.0240233f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_62 N_A1_c_61_n N_A2_c_93_n 0.0101924f $X=0.49 $Y=1.69 $X2=0 $Y2=0
cc_63 N_A1_c_66_n N_A2_c_98_n 0.041607f $X=0.49 $Y=1.84 $X2=0 $Y2=0
cc_64 N_A1_c_66_n A2 5.90806e-19 $X=0.49 $Y=1.84 $X2=0 $Y2=0
cc_65 A1 A2 0.033285f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A1_c_63_n A2 0.00205502f $X=0.46 $Y=1.335 $X2=0 $Y2=0
cc_67 A1 N_A2_c_95_n 0.00255585f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A1_c_63_n N_A2_c_95_n 0.0101924f $X=0.46 $Y=1.335 $X2=0 $Y2=0
cc_69 N_A1_M1007_g N_VPWR_c_223_n 0.0267198f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_70 N_A1_c_66_n N_VPWR_c_223_n 0.00108458f $X=0.49 $Y=1.84 $X2=0 $Y2=0
cc_71 A1 N_VPWR_c_223_n 0.0280391f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A1_M1007_g N_VPWR_c_225_n 0.00802402f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_73 N_A1_M1007_g N_VPWR_c_221_n 0.0142664f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_74 N_A1_M1004_g N_A_38_57#_c_302_n 0.0111794f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_75 N_A1_M1004_g N_A_38_57#_c_303_n 0.00926821f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_76 A1 N_A_38_57#_c_303_n 0.00897633f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A1_M1004_g N_A_38_57#_c_304_n 0.004207f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_78 A1 N_A_38_57#_c_304_n 0.0285986f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A1_c_63_n N_A_38_57#_c_304_n 0.00139878f $X=0.46 $Y=1.335 $X2=0 $Y2=0
cc_80 N_A1_M1004_g N_A_38_57#_c_305_n 8.85777e-19 $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_81 N_A1_M1004_g N_VGND_c_333_n 0.00507706f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_82 N_A1_M1004_g N_VGND_c_335_n 0.00656529f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_83 N_A1_M1004_g N_VGND_c_336_n 0.00502664f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_84 N_A2_M1005_g N_B1_M1001_g 0.0296364f $X=1.14 $Y=0.495 $X2=0 $Y2=0
cc_85 N_A2_M1003_g N_B1_M1006_g 0.0151052f $X=1.05 $Y=2.545 $X2=0 $Y2=0
cc_86 N_A2_c_93_n N_B1_c_134_n 0.0117523f $X=1.09 $Y=1.675 $X2=0 $Y2=0
cc_87 N_A2_c_98_n N_B1_c_139_n 0.0117523f $X=1.09 $Y=1.84 $X2=0 $Y2=0
cc_88 A2 B1 0.0514086f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A2_c_95_n B1 7.56445e-19 $X=1.09 $Y=1.335 $X2=0 $Y2=0
cc_90 A2 N_B1_c_136_n 0.00411743f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A2_c_95_n N_B1_c_136_n 0.0117523f $X=1.09 $Y=1.335 $X2=0 $Y2=0
cc_92 N_A2_M1003_g N_VPWR_c_223_n 0.00519241f $X=1.05 $Y=2.545 $X2=0 $Y2=0
cc_93 N_A2_M1003_g N_VPWR_c_224_n 7.97642e-19 $X=1.05 $Y=2.545 $X2=0 $Y2=0
cc_94 N_A2_M1003_g N_VPWR_c_225_n 0.00893366f $X=1.05 $Y=2.545 $X2=0 $Y2=0
cc_95 N_A2_M1003_g N_VPWR_c_221_n 0.016682f $X=1.05 $Y=2.545 $X2=0 $Y2=0
cc_96 N_A2_M1003_g N_Y_c_255_n 5.70164e-19 $X=1.05 $Y=2.545 $X2=0 $Y2=0
cc_97 N_A2_M1003_g N_Y_c_257_n 8.32582e-19 $X=1.05 $Y=2.545 $X2=0 $Y2=0
cc_98 N_A2_c_98_n N_Y_c_257_n 5.05028e-19 $X=1.09 $Y=1.84 $X2=0 $Y2=0
cc_99 A2 N_Y_c_257_n 0.010844f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A2_M1005_g N_A_38_57#_c_302_n 8.85777e-19 $X=1.14 $Y=0.495 $X2=0 $Y2=0
cc_101 N_A2_M1005_g N_A_38_57#_c_303_n 0.0120381f $X=1.14 $Y=0.495 $X2=0 $Y2=0
cc_102 A2 N_A_38_57#_c_303_n 0.0304022f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_A2_c_95_n N_A_38_57#_c_303_n 0.00126602f $X=1.09 $Y=1.335 $X2=0 $Y2=0
cc_104 N_A2_M1005_g N_A_38_57#_c_305_n 0.00978191f $X=1.14 $Y=0.495 $X2=0 $Y2=0
cc_105 N_A2_M1005_g N_VGND_c_333_n 0.00507706f $X=1.14 $Y=0.495 $X2=0 $Y2=0
cc_106 N_A2_M1005_g N_VGND_c_334_n 0.00502664f $X=1.14 $Y=0.495 $X2=0 $Y2=0
cc_107 N_A2_M1005_g N_VGND_c_335_n 0.00589314f $X=1.14 $Y=0.495 $X2=0 $Y2=0
cc_108 N_B1_M1001_g N_C1_c_176_n 0.0402196f $X=1.57 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_109 N_B1_M1006_g N_C1_M1000_g 0.0261747f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_110 B1 N_C1_M1000_g 4.04747e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B1_M1001_g N_C1_c_178_n 0.00744953f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_112 N_B1_c_134_n N_C1_c_179_n 0.0119227f $X=1.66 $Y=1.675 $X2=0 $Y2=0
cc_113 N_B1_c_139_n N_C1_c_180_n 0.0119227f $X=1.66 $Y=1.84 $X2=0 $Y2=0
cc_114 N_B1_M1001_g C1 0.00114765f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_115 B1 C1 0.0399467f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_116 N_B1_c_136_n C1 0.00373413f $X=1.66 $Y=1.335 $X2=0 $Y2=0
cc_117 B1 N_C1_c_182_n 7.49315e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B1_c_136_n N_C1_c_182_n 0.0119227f $X=1.66 $Y=1.335 $X2=0 $Y2=0
cc_119 N_B1_M1006_g N_VPWR_c_224_n 0.0164699f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_120 N_B1_M1006_g N_VPWR_c_225_n 0.00769046f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_121 N_B1_M1006_g N_VPWR_c_221_n 0.0135127f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_122 N_B1_M1006_g N_Y_c_255_n 0.0158534f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_123 N_B1_M1006_g N_Y_c_256_n 0.0180783f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_124 N_B1_c_139_n N_Y_c_256_n 5.43485e-19 $X=1.66 $Y=1.84 $X2=0 $Y2=0
cc_125 B1 N_Y_c_256_n 0.0223517f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B1_M1006_g N_Y_c_257_n 0.0010172f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_127 B1 N_Y_c_257_n 0.00193735f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_128 N_B1_M1006_g N_Y_c_258_n 8.9454e-19 $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_129 N_B1_M1001_g N_Y_c_254_n 0.00129114f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_130 N_B1_M1001_g N_A_38_57#_c_303_n 0.00578619f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_131 B1 N_A_38_57#_c_303_n 0.00193735f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_M1001_g N_A_38_57#_c_305_n 0.011386f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_133 N_B1_M1001_g N_VGND_c_334_n 0.00502664f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_134 N_B1_M1001_g N_VGND_c_335_n 0.00950403f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_135 N_C1_M1000_g N_VPWR_c_224_n 0.00298779f $X=2.19 $Y=2.545 $X2=0 $Y2=0
cc_136 N_C1_M1000_g N_VPWR_c_227_n 0.0086001f $X=2.19 $Y=2.545 $X2=0 $Y2=0
cc_137 N_C1_M1000_g N_VPWR_c_221_n 0.0163435f $X=2.19 $Y=2.545 $X2=0 $Y2=0
cc_138 N_C1_M1000_g N_Y_c_255_n 8.62562e-19 $X=2.19 $Y=2.545 $X2=0 $Y2=0
cc_139 N_C1_M1000_g N_Y_c_256_n 0.0193288f $X=2.19 $Y=2.545 $X2=0 $Y2=0
cc_140 C1 N_Y_c_256_n 0.0142099f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_141 N_C1_M1000_g N_Y_c_258_n 0.0143167f $X=2.19 $Y=2.545 $X2=0 $Y2=0
cc_142 N_C1_c_176_n N_Y_c_253_n 0.00124366f $X=1.96 $Y=0.78 $X2=0 $Y2=0
cc_143 N_C1_M1000_g N_Y_c_253_n 0.00779971f $X=2.19 $Y=2.545 $X2=0 $Y2=0
cc_144 N_C1_c_177_n N_Y_c_253_n 0.00951333f $X=2.14 $Y=0.855 $X2=0 $Y2=0
cc_145 C1 N_Y_c_253_n 0.0464518f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_146 N_C1_c_182_n N_Y_c_253_n 0.0147882f $X=2.23 $Y=1.275 $X2=0 $Y2=0
cc_147 N_C1_M1000_g N_Y_c_260_n 0.00134807f $X=2.19 $Y=2.545 $X2=0 $Y2=0
cc_148 N_C1_c_180_n N_Y_c_260_n 5.9401e-19 $X=2.23 $Y=1.78 $X2=0 $Y2=0
cc_149 C1 N_Y_c_260_n 0.00702626f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_150 N_C1_c_176_n N_Y_c_254_n 0.0105535f $X=1.96 $Y=0.78 $X2=0 $Y2=0
cc_151 N_C1_c_177_n N_Y_c_254_n 0.00616548f $X=2.14 $Y=0.855 $X2=0 $Y2=0
cc_152 C1 N_Y_c_254_n 0.0162955f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_153 N_C1_c_182_n N_Y_c_254_n 0.00118553f $X=2.23 $Y=1.275 $X2=0 $Y2=0
cc_154 N_C1_c_177_n N_A_38_57#_c_303_n 5.8374e-19 $X=2.14 $Y=0.855 $X2=0 $Y2=0
cc_155 N_C1_c_178_n N_A_38_57#_c_303_n 2.69321e-19 $X=2.23 $Y=1.11 $X2=0 $Y2=0
cc_156 N_C1_c_176_n N_A_38_57#_c_305_n 0.00178748f $X=1.96 $Y=0.78 $X2=0 $Y2=0
cc_157 N_C1_c_176_n N_VGND_c_334_n 0.00501304f $X=1.96 $Y=0.78 $X2=0 $Y2=0
cc_158 N_C1_c_176_n N_VGND_c_335_n 0.0103493f $X=1.96 $Y=0.78 $X2=0 $Y2=0
cc_159 N_VPWR_c_224_n N_Y_c_255_n 0.045794f $X=1.885 $Y=2.535 $X2=0 $Y2=0
cc_160 N_VPWR_c_225_n N_Y_c_255_n 0.0220321f $X=1.72 $Y=3.33 $X2=0 $Y2=0
cc_161 N_VPWR_c_221_n N_Y_c_255_n 0.0125808f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_162 N_VPWR_M1006_d N_Y_c_256_n 0.00224299f $X=1.745 $Y=2.045 $X2=0 $Y2=0
cc_163 N_VPWR_c_224_n N_Y_c_256_n 0.017764f $X=1.885 $Y=2.535 $X2=0 $Y2=0
cc_164 N_VPWR_c_224_n N_Y_c_258_n 0.0214848f $X=1.885 $Y=2.535 $X2=0 $Y2=0
cc_165 N_VPWR_c_227_n N_Y_c_258_n 0.0311344f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_166 N_VPWR_c_221_n N_Y_c_258_n 0.0178044f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_167 N_Y_c_254_n N_A_38_57#_c_305_n 0.0153883f $X=2.585 $Y=0.495 $X2=0 $Y2=0
cc_168 N_Y_c_252_n N_VGND_c_334_n 0.0114622f $X=2.67 $Y=0.725 $X2=0 $Y2=0
cc_169 N_Y_c_254_n N_VGND_c_334_n 0.0373076f $X=2.585 $Y=0.495 $X2=0 $Y2=0
cc_170 N_Y_c_252_n N_VGND_c_335_n 0.00657784f $X=2.67 $Y=0.725 $X2=0 $Y2=0
cc_171 N_Y_c_254_n N_VGND_c_335_n 0.0218851f $X=2.585 $Y=0.495 $X2=0 $Y2=0
cc_172 N_A_38_57#_c_302_n N_VGND_c_333_n 0.0141997f $X=0.335 $Y=0.495 $X2=0
+ $Y2=0
cc_173 N_A_38_57#_c_303_n N_VGND_c_333_n 0.0251886f $X=1.19 $Y=0.905 $X2=0 $Y2=0
cc_174 N_A_38_57#_c_305_n N_VGND_c_333_n 0.0141997f $X=1.355 $Y=0.495 $X2=0
+ $Y2=0
cc_175 N_A_38_57#_c_305_n N_VGND_c_334_n 0.021949f $X=1.355 $Y=0.495 $X2=0 $Y2=0
cc_176 N_A_38_57#_c_302_n N_VGND_c_335_n 0.0125808f $X=0.335 $Y=0.495 $X2=0
+ $Y2=0
cc_177 N_A_38_57#_c_303_n N_VGND_c_335_n 0.0120154f $X=1.19 $Y=0.905 $X2=0 $Y2=0
cc_178 N_A_38_57#_c_305_n N_VGND_c_335_n 0.0124703f $X=1.355 $Y=0.495 $X2=0
+ $Y2=0
cc_179 N_A_38_57#_c_302_n N_VGND_c_336_n 0.0220321f $X=0.335 $Y=0.495 $X2=0
+ $Y2=0
