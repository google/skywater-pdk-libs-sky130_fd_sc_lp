* File: sky130_fd_sc_lp__and4bb_1.pxi.spice
* Created: Fri Aug 28 10:09:03 2020
* 
x_PM_SKY130_FD_SC_LP__AND4BB_1%A_N N_A_N_M1009_g N_A_N_M1003_g N_A_N_c_99_n A_N
+ A_N N_A_N_c_100_n N_A_N_c_101_n A_N PM_SKY130_FD_SC_LP__AND4BB_1%A_N
x_PM_SKY130_FD_SC_LP__AND4BB_1%B_N N_B_N_M1000_g N_B_N_M1005_g N_B_N_c_138_n
+ N_B_N_c_144_n B_N N_B_N_c_139_n N_B_N_c_140_n N_B_N_c_141_n
+ PM_SKY130_FD_SC_LP__AND4BB_1%B_N
x_PM_SKY130_FD_SC_LP__AND4BB_1%A_27_51# N_A_27_51#_M1009_s N_A_27_51#_M1003_s
+ N_A_27_51#_c_185_n N_A_27_51#_M1006_g N_A_27_51#_M1013_g N_A_27_51#_c_188_n
+ N_A_27_51#_c_189_n N_A_27_51#_c_190_n N_A_27_51#_c_191_n N_A_27_51#_c_192_n
+ N_A_27_51#_c_198_n N_A_27_51#_c_193_n N_A_27_51#_c_194_n N_A_27_51#_c_195_n
+ PM_SKY130_FD_SC_LP__AND4BB_1%A_27_51#
x_PM_SKY130_FD_SC_LP__AND4BB_1%A_196_51# N_A_196_51#_M1000_d N_A_196_51#_M1005_d
+ N_A_196_51#_M1007_g N_A_196_51#_M1004_g N_A_196_51#_c_272_n
+ N_A_196_51#_c_264_n N_A_196_51#_c_273_n N_A_196_51#_c_274_n
+ N_A_196_51#_c_265_n N_A_196_51#_c_266_n N_A_196_51#_c_267_n
+ N_A_196_51#_c_268_n N_A_196_51#_c_269_n N_A_196_51#_c_270_n
+ PM_SKY130_FD_SC_LP__AND4BB_1%A_196_51#
x_PM_SKY130_FD_SC_LP__AND4BB_1%C N_C_M1001_g N_C_M1002_g C C N_C_c_347_n
+ N_C_c_348_n PM_SKY130_FD_SC_LP__AND4BB_1%C
x_PM_SKY130_FD_SC_LP__AND4BB_1%D N_D_M1010_g N_D_M1008_g D N_D_c_383_n
+ PM_SKY130_FD_SC_LP__AND4BB_1%D
x_PM_SKY130_FD_SC_LP__AND4BB_1%A_344_131# N_A_344_131#_M1013_s
+ N_A_344_131#_M1006_d N_A_344_131#_M1001_d N_A_344_131#_M1012_g
+ N_A_344_131#_M1011_g N_A_344_131#_c_408_n N_A_344_131#_c_409_n
+ N_A_344_131#_c_414_n N_A_344_131#_c_415_n N_A_344_131#_c_416_n
+ N_A_344_131#_c_417_n N_A_344_131#_c_410_n N_A_344_131#_c_411_n
+ N_A_344_131#_c_420_n N_A_344_131#_c_421_n
+ PM_SKY130_FD_SC_LP__AND4BB_1%A_344_131#
x_PM_SKY130_FD_SC_LP__AND4BB_1%VPWR N_VPWR_M1003_d N_VPWR_M1006_s N_VPWR_M1004_d
+ N_VPWR_M1008_d N_VPWR_c_482_n N_VPWR_c_483_n N_VPWR_c_484_n N_VPWR_c_485_n
+ N_VPWR_c_486_n N_VPWR_c_532_n VPWR N_VPWR_c_487_n N_VPWR_c_488_n
+ N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_481_n N_VPWR_c_492_n N_VPWR_c_493_n
+ N_VPWR_c_494_n N_VPWR_c_495_n PM_SKY130_FD_SC_LP__AND4BB_1%VPWR
x_PM_SKY130_FD_SC_LP__AND4BB_1%X N_X_M1012_d N_X_M1011_d N_X_c_542_n N_X_c_543_n
+ N_X_c_539_n X X N_X_c_541_n X PM_SKY130_FD_SC_LP__AND4BB_1%X
x_PM_SKY130_FD_SC_LP__AND4BB_1%VGND N_VGND_M1009_d N_VGND_M1010_d N_VGND_c_559_n
+ N_VGND_c_560_n VGND N_VGND_c_561_n N_VGND_c_562_n N_VGND_c_563_n
+ N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n PM_SKY130_FD_SC_LP__AND4BB_1%VGND
cc_1 VNB N_A_N_M1009_g 0.0702375f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.465
cc_2 VNB N_B_N_c_138_n 0.0301742f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.67
cc_3 VNB N_B_N_c_139_n 0.0332817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_4 VNB N_B_N_c_140_n 0.00791639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_B_N_c_141_n 0.0200929f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.835
cc_6 VNB N_A_27_51#_c_185_n 0.0214859f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.865
cc_7 VNB N_A_27_51#_M1006_g 0.00740161f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.175
cc_8 VNB N_A_27_51#_M1013_g 0.0247896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_51#_c_188_n 0.0103974f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.835
cc_10 VNB N_A_27_51#_c_189_n 0.0505613f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.005
cc_11 VNB N_A_27_51#_c_190_n 0.00740553f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.062
cc_12 VNB N_A_27_51#_c_191_n 0.00716999f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.977
cc_13 VNB N_A_27_51#_c_192_n 0.0121549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_51#_c_193_n 0.0075431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_51#_c_194_n 0.00238558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_51#_c_195_n 0.0263563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_196_51#_M1007_g 0.035715f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.835
cc_18 VNB N_A_196_51#_c_264_n 0.0117156f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.835
cc_19 VNB N_A_196_51#_c_265_n 0.031174f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.062
cc_20 VNB N_A_196_51#_c_266_n 0.0489373f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.405
cc_21 VNB N_A_196_51#_c_267_n 0.0094115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_196_51#_c_268_n 0.00393145f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.835
cc_23 VNB N_A_196_51#_c_269_n 0.00461729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_196_51#_c_270_n 0.0110052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C_M1001_g 0.00773869f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.465
cc_26 VNB C 0.0064456f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.67
cc_27 VNB N_C_c_347_n 0.0279135f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.835
cc_28 VNB N_C_c_348_n 0.0165075f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.835
cc_29 VNB N_D_M1010_g 0.0393043f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.465
cc_30 VNB N_A_344_131#_M1012_g 0.0320822f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_31 VNB N_A_344_131#_c_408_n 0.00281335f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.835
cc_32 VNB N_A_344_131#_c_409_n 0.00500651f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.062
cc_33 VNB N_A_344_131#_c_410_n 0.00222647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_344_131#_c_411_n 0.028459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_481_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_539_n 0.0280384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB X 0.010088f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.835
cc_38 VNB N_X_c_541_n 0.0268936f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.062
cc_39 VNB N_VGND_c_559_n 0.00586594f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.835
cc_40 VNB N_VGND_c_560_n 0.0227161f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_41 VNB N_VGND_c_561_n 0.0173198f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.835
cc_42 VNB N_VGND_c_562_n 0.065042f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.405
cc_43 VNB N_VGND_c_563_n 0.0172252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_564_n 0.253296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_565_n 0.00497591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_566_n 0.00615512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VPB N_A_N_M1009_g 8.34254e-19 $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.465
cc_48 VPB N_A_N_M1003_g 0.0228055f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.865
cc_49 VPB N_A_N_c_99_n 0.0491544f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.175
cc_50 VPB N_A_N_c_100_n 0.016348f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.835
cc_51 VPB N_A_N_c_101_n 0.0061067f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.005
cc_52 VPB A_N 0.00847724f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.035
cc_53 VPB N_B_N_M1005_g 0.044906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B_N_c_138_n 0.0168913f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.67
cc_55 VPB N_B_N_c_144_n 0.0104883f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.175
cc_56 VPB N_A_27_51#_M1006_g 0.0334591f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.175
cc_57 VPB N_A_27_51#_c_190_n 0.0492883f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.062
cc_58 VPB N_A_27_51#_c_198_n 0.0156757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_27_51#_c_195_n 0.00983237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_196_51#_M1007_g 0.0279097f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.835
cc_61 VPB N_A_196_51#_c_272_n 0.0231662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_196_51#_c_273_n 0.0152964f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.835
cc_63 VPB N_A_196_51#_c_274_n 0.0046449f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.005
cc_64 VPB N_A_196_51#_c_269_n 0.00369093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_C_M1001_g 0.0287143f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.465
cc_66 VPB N_D_M1010_g 0.0388515f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.465
cc_67 VPB D 0.00750014f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.865
cc_68 VPB N_D_c_383_n 0.0496531f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_69 VPB N_A_344_131#_M1011_g 0.0245544f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_344_131#_c_409_n 7.67686e-19 $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.062
cc_71 VPB N_A_344_131#_c_414_n 0.00144289f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_344_131#_c_415_n 0.00987183f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.977
cc_73 VPB N_A_344_131#_c_416_n 0.00158757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_344_131#_c_417_n 0.00550809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_344_131#_c_410_n 3.00451e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_344_131#_c_411_n 0.00674388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_344_131#_c_420_n 0.00148998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_344_131#_c_421_n 0.00230243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_482_n 8.60259e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_483_n 0.0176419f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.835
cc_81 VPB N_VPWR_c_484_n 0.0270275f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=2.035
cc_82 VPB N_VPWR_c_485_n 0.0248916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_486_n 0.00507937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_487_n 0.0179742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_488_n 0.0172794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_489_n 0.0186178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_490_n 0.0172252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_481_n 0.0858255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_492_n 0.00461449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_493_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_494_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_495_n 0.00458712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_X_c_542_n 0.00601347f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.865
cc_94 VPB N_X_c_543_n 0.0346529f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.835
cc_95 VPB N_X_c_539_n 0.0160993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 N_A_N_M1003_g N_B_N_M1005_g 0.0141636f $X=0.575 $Y=2.865 $X2=0 $Y2=0
cc_97 N_A_N_c_99_n N_B_N_M1005_g 0.0203407f $X=0.525 $Y=2.175 $X2=0 $Y2=0
cc_98 A_N N_B_N_M1005_g 0.00391571f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A_N_M1009_g N_B_N_c_138_n 0.0192382f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_100 N_A_N_c_100_n N_B_N_c_138_n 0.0119082f $X=0.525 $Y=1.835 $X2=0 $Y2=0
cc_101 N_A_N_c_101_n N_B_N_c_138_n 0.00268771f $X=0.66 $Y=2.005 $X2=0 $Y2=0
cc_102 N_A_N_c_99_n N_B_N_c_144_n 0.0119082f $X=0.525 $Y=2.175 $X2=0 $Y2=0
cc_103 A_N N_B_N_c_144_n 6.1274e-19 $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_104 N_A_N_M1009_g N_B_N_c_140_n 0.00281502f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_105 N_A_N_M1009_g N_B_N_c_141_n 0.0260517f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_106 N_A_N_M1009_g N_A_27_51#_c_189_n 0.0225793f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_107 N_A_N_M1009_g N_A_27_51#_c_190_n 0.00479712f $X=0.475 $Y=0.465 $X2=0
+ $Y2=0
cc_108 N_A_N_M1003_g N_A_27_51#_c_190_n 0.00492848f $X=0.575 $Y=2.865 $X2=0
+ $Y2=0
cc_109 N_A_N_c_99_n N_A_27_51#_c_190_n 0.00113928f $X=0.525 $Y=2.175 $X2=0 $Y2=0
cc_110 N_A_N_c_100_n N_A_27_51#_c_190_n 0.0163603f $X=0.525 $Y=1.835 $X2=0 $Y2=0
cc_111 N_A_N_c_101_n N_A_27_51#_c_190_n 0.0243715f $X=0.66 $Y=2.005 $X2=0 $Y2=0
cc_112 A_N N_A_27_51#_c_190_n 0.0393837f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_113 N_A_N_c_100_n N_A_27_51#_c_192_n 0.00143974f $X=0.525 $Y=1.835 $X2=0
+ $Y2=0
cc_114 N_A_N_c_99_n N_A_27_51#_c_198_n 0.0029681f $X=0.525 $Y=2.175 $X2=0 $Y2=0
cc_115 A_N N_A_27_51#_c_198_n 6.96421e-19 $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_116 N_A_N_M1009_g N_A_27_51#_c_193_n 0.0180238f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_117 N_A_N_c_100_n N_A_27_51#_c_193_n 0.00136753f $X=0.525 $Y=1.835 $X2=0
+ $Y2=0
cc_118 N_A_N_c_101_n N_A_27_51#_c_193_n 0.0307588f $X=0.66 $Y=2.005 $X2=0 $Y2=0
cc_119 N_A_N_M1009_g N_A_27_51#_c_194_n 4.32637e-19 $X=0.475 $Y=0.465 $X2=0
+ $Y2=0
cc_120 N_A_N_c_101_n N_A_196_51#_c_272_n 0.00321533f $X=0.66 $Y=2.005 $X2=0
+ $Y2=0
cc_121 A_N N_A_196_51#_c_272_n 0.0339469f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_122 N_A_N_c_101_n N_A_196_51#_c_274_n 0.0119035f $X=0.66 $Y=2.005 $X2=0 $Y2=0
cc_123 N_A_N_M1003_g N_VPWR_c_482_n 0.0109733f $X=0.575 $Y=2.865 $X2=0 $Y2=0
cc_124 A_N N_VPWR_c_482_n 0.0196053f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_125 N_A_N_M1003_g N_VPWR_c_487_n 0.00469214f $X=0.575 $Y=2.865 $X2=0 $Y2=0
cc_126 N_A_N_M1003_g N_VPWR_c_481_n 0.00536787f $X=0.575 $Y=2.865 $X2=0 $Y2=0
cc_127 A_N N_VPWR_c_481_n 0.00700273f $X=0.72 $Y=2.035 $X2=0 $Y2=0
cc_128 N_A_N_M1009_g N_VGND_c_559_n 0.00303117f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_129 N_A_N_M1009_g N_VGND_c_561_n 0.00565115f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_130 N_A_N_M1009_g N_VGND_c_564_n 0.0114017f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_131 N_B_N_c_140_n N_A_27_51#_c_189_n 0.0281934f $X=0.995 $Y=0.95 $X2=0 $Y2=0
cc_132 N_B_N_c_139_n N_A_27_51#_c_191_n 0.00211276f $X=0.995 $Y=0.95 $X2=0 $Y2=0
cc_133 N_B_N_c_138_n N_A_27_51#_c_193_n 0.00410577f $X=0.99 $Y=1.925 $X2=0 $Y2=0
cc_134 N_B_N_c_139_n N_A_27_51#_c_193_n 0.00178607f $X=0.995 $Y=0.95 $X2=0 $Y2=0
cc_135 N_B_N_c_140_n N_A_27_51#_c_193_n 0.0336815f $X=0.995 $Y=0.95 $X2=0 $Y2=0
cc_136 N_B_N_c_138_n N_A_27_51#_c_194_n 0.015091f $X=0.99 $Y=1.925 $X2=0 $Y2=0
cc_137 N_B_N_c_144_n N_A_27_51#_c_194_n 0.00112893f $X=0.99 $Y=2.075 $X2=0 $Y2=0
cc_138 N_B_N_c_139_n N_A_27_51#_c_194_n 0.00123045f $X=0.995 $Y=0.95 $X2=0 $Y2=0
cc_139 N_B_N_c_138_n N_A_27_51#_c_195_n 0.0217969f $X=0.99 $Y=1.925 $X2=0 $Y2=0
cc_140 N_B_N_c_144_n N_A_196_51#_c_272_n 0.0191414f $X=0.99 $Y=2.075 $X2=0 $Y2=0
cc_141 N_B_N_c_139_n N_A_196_51#_c_264_n 0.00701101f $X=0.995 $Y=0.95 $X2=0
+ $Y2=0
cc_142 N_B_N_c_140_n N_A_196_51#_c_264_n 0.0174619f $X=0.995 $Y=0.95 $X2=0 $Y2=0
cc_143 N_B_N_c_141_n N_A_196_51#_c_264_n 0.00437359f $X=0.995 $Y=0.785 $X2=0
+ $Y2=0
cc_144 N_B_N_c_138_n N_A_196_51#_c_274_n 0.00332703f $X=0.99 $Y=1.925 $X2=0
+ $Y2=0
cc_145 N_B_N_c_144_n N_A_196_51#_c_274_n 7.70472e-19 $X=0.99 $Y=2.075 $X2=0
+ $Y2=0
cc_146 N_B_N_c_138_n N_A_196_51#_c_268_n 0.00498903f $X=0.99 $Y=1.925 $X2=0
+ $Y2=0
cc_147 N_B_N_c_139_n N_A_196_51#_c_268_n 7.51442e-19 $X=0.995 $Y=0.95 $X2=0
+ $Y2=0
cc_148 N_B_N_c_140_n N_A_196_51#_c_268_n 0.00188088f $X=0.995 $Y=0.95 $X2=0
+ $Y2=0
cc_149 N_B_N_c_139_n N_A_196_51#_c_270_n 0.00543552f $X=0.995 $Y=0.95 $X2=0
+ $Y2=0
cc_150 N_B_N_c_140_n N_A_196_51#_c_270_n 0.00491754f $X=0.995 $Y=0.95 $X2=0
+ $Y2=0
cc_151 N_B_N_M1005_g N_VPWR_c_482_n 0.00985813f $X=1.005 $Y=2.865 $X2=0 $Y2=0
cc_152 N_B_N_M1005_g N_VPWR_c_483_n 0.00469214f $X=1.005 $Y=2.865 $X2=0 $Y2=0
cc_153 N_B_N_M1005_g N_VPWR_c_484_n 0.00324015f $X=1.005 $Y=2.865 $X2=0 $Y2=0
cc_154 N_B_N_M1005_g N_VPWR_c_481_n 0.00945295f $X=1.005 $Y=2.865 $X2=0 $Y2=0
cc_155 N_B_N_c_140_n N_VGND_c_559_n 0.0176204f $X=0.995 $Y=0.95 $X2=0 $Y2=0
cc_156 N_B_N_c_141_n N_VGND_c_559_n 0.00303117f $X=0.995 $Y=0.785 $X2=0 $Y2=0
cc_157 N_B_N_c_141_n N_VGND_c_562_n 0.00565115f $X=0.995 $Y=0.785 $X2=0 $Y2=0
cc_158 N_B_N_c_139_n N_VGND_c_564_n 2.64147e-19 $X=0.995 $Y=0.95 $X2=0 $Y2=0
cc_159 N_B_N_c_140_n N_VGND_c_564_n 0.00650556f $X=0.995 $Y=0.95 $X2=0 $Y2=0
cc_160 N_B_N_c_141_n N_VGND_c_564_n 0.00715583f $X=0.995 $Y=0.785 $X2=0 $Y2=0
cc_161 N_A_27_51#_M1006_g N_A_196_51#_M1007_g 0.0232918f $X=1.99 $Y=2.175 $X2=0
+ $Y2=0
cc_162 N_A_27_51#_c_188_n N_A_196_51#_M1007_g 0.029116f $X=2.025 $Y=1.43 $X2=0
+ $Y2=0
cc_163 N_A_27_51#_M1006_g N_A_196_51#_c_272_n 0.00406608f $X=1.99 $Y=2.175 $X2=0
+ $Y2=0
cc_164 N_A_27_51#_M1013_g N_A_196_51#_c_264_n 0.00275566f $X=2.06 $Y=0.865 $X2=0
+ $Y2=0
cc_165 N_A_27_51#_c_185_n N_A_196_51#_c_273_n 0.00355672f $X=1.915 $Y=1.43 $X2=0
+ $Y2=0
cc_166 N_A_27_51#_M1006_g N_A_196_51#_c_273_n 0.00617381f $X=1.99 $Y=2.175 $X2=0
+ $Y2=0
cc_167 N_A_27_51#_c_191_n N_A_196_51#_c_273_n 0.0147434f $X=1.425 $Y=1.52 $X2=0
+ $Y2=0
cc_168 N_A_27_51#_c_195_n N_A_196_51#_c_273_n 0.00499008f $X=1.425 $Y=1.43 $X2=0
+ $Y2=0
cc_169 N_A_27_51#_c_191_n N_A_196_51#_c_274_n 0.0216471f $X=1.425 $Y=1.52 $X2=0
+ $Y2=0
cc_170 N_A_27_51#_c_195_n N_A_196_51#_c_274_n 0.00317024f $X=1.425 $Y=1.43 $X2=0
+ $Y2=0
cc_171 N_A_27_51#_M1013_g N_A_196_51#_c_265_n 0.00476174f $X=2.06 $Y=0.865 $X2=0
+ $Y2=0
cc_172 N_A_27_51#_M1013_g N_A_196_51#_c_266_n 0.029116f $X=2.06 $Y=0.865 $X2=0
+ $Y2=0
cc_173 N_A_27_51#_M1013_g N_A_196_51#_c_267_n 0.00394147f $X=2.06 $Y=0.865 $X2=0
+ $Y2=0
cc_174 N_A_27_51#_c_191_n N_A_196_51#_c_267_n 0.00645161f $X=1.425 $Y=1.52 $X2=0
+ $Y2=0
cc_175 N_A_27_51#_c_195_n N_A_196_51#_c_267_n 0.00666476f $X=1.425 $Y=1.43 $X2=0
+ $Y2=0
cc_176 N_A_27_51#_c_191_n N_A_196_51#_c_268_n 0.0137437f $X=1.425 $Y=1.52 $X2=0
+ $Y2=0
cc_177 N_A_27_51#_c_195_n N_A_196_51#_c_268_n 0.00429589f $X=1.425 $Y=1.43 $X2=0
+ $Y2=0
cc_178 N_A_27_51#_c_185_n N_A_196_51#_c_269_n 0.0109167f $X=1.915 $Y=1.43 $X2=0
+ $Y2=0
cc_179 N_A_27_51#_M1006_g N_A_196_51#_c_269_n 0.00601331f $X=1.99 $Y=2.175 $X2=0
+ $Y2=0
cc_180 N_A_27_51#_M1013_g N_A_196_51#_c_269_n 0.00219834f $X=2.06 $Y=0.865 $X2=0
+ $Y2=0
cc_181 N_A_27_51#_c_188_n N_A_196_51#_c_269_n 0.00273114f $X=2.025 $Y=1.43 $X2=0
+ $Y2=0
cc_182 N_A_27_51#_c_191_n N_A_196_51#_c_269_n 0.0140713f $X=1.425 $Y=1.52 $X2=0
+ $Y2=0
cc_183 N_A_27_51#_c_194_n N_A_196_51#_c_269_n 0.00274132f $X=1.095 $Y=1.472
+ $X2=0 $Y2=0
cc_184 N_A_27_51#_c_195_n N_A_196_51#_c_269_n 0.00189618f $X=1.425 $Y=1.43 $X2=0
+ $Y2=0
cc_185 N_A_27_51#_M1013_g N_A_196_51#_c_270_n 0.00251105f $X=2.06 $Y=0.865 $X2=0
+ $Y2=0
cc_186 N_A_27_51#_c_185_n N_A_344_131#_c_408_n 7.97138e-19 $X=1.915 $Y=1.43
+ $X2=0 $Y2=0
cc_187 N_A_27_51#_M1013_g N_A_344_131#_c_408_n 0.0117284f $X=2.06 $Y=0.865 $X2=0
+ $Y2=0
cc_188 N_A_27_51#_M1006_g N_A_344_131#_c_409_n 0.00144148f $X=1.99 $Y=2.175
+ $X2=0 $Y2=0
cc_189 N_A_27_51#_M1013_g N_A_344_131#_c_409_n 0.00920283f $X=2.06 $Y=0.865
+ $X2=0 $Y2=0
cc_190 N_A_27_51#_c_188_n N_A_344_131#_c_409_n 0.00394312f $X=2.025 $Y=1.43
+ $X2=0 $Y2=0
cc_191 N_A_27_51#_M1006_g N_A_344_131#_c_414_n 8.70795e-19 $X=1.99 $Y=2.175
+ $X2=0 $Y2=0
cc_192 N_A_27_51#_M1006_g N_A_344_131#_c_420_n 0.00140038f $X=1.99 $Y=2.175
+ $X2=0 $Y2=0
cc_193 N_A_27_51#_c_185_n N_VPWR_c_484_n 6.17285e-19 $X=1.915 $Y=1.43 $X2=0
+ $Y2=0
cc_194 N_A_27_51#_M1006_g N_VPWR_c_484_n 0.00882102f $X=1.99 $Y=2.175 $X2=0
+ $Y2=0
cc_195 N_A_27_51#_M1006_g N_VPWR_c_485_n 5.20255e-19 $X=1.99 $Y=2.175 $X2=0
+ $Y2=0
cc_196 N_A_27_51#_c_198_n N_VPWR_c_487_n 0.0186542f $X=0.36 $Y=2.865 $X2=0 $Y2=0
cc_197 N_A_27_51#_M1006_g N_VPWR_c_481_n 0.00327084f $X=1.99 $Y=2.175 $X2=0
+ $Y2=0
cc_198 N_A_27_51#_c_198_n N_VPWR_c_481_n 0.0135709f $X=0.36 $Y=2.865 $X2=0 $Y2=0
cc_199 N_A_27_51#_c_189_n N_VGND_c_561_n 0.0162918f $X=0.26 $Y=0.45 $X2=0 $Y2=0
cc_200 N_A_27_51#_c_189_n N_VGND_c_564_n 0.0114155f $X=0.26 $Y=0.45 $X2=0 $Y2=0
cc_201 N_A_196_51#_M1007_g N_C_M1001_g 0.0226319f $X=2.42 $Y=0.865 $X2=0 $Y2=0
cc_202 N_A_196_51#_M1007_g C 0.00751424f $X=2.42 $Y=0.865 $X2=0 $Y2=0
cc_203 N_A_196_51#_c_265_n C 0.00667789f $X=2.51 $Y=0.38 $X2=0 $Y2=0
cc_204 N_A_196_51#_c_266_n C 0.00281563f $X=2.51 $Y=0.38 $X2=0 $Y2=0
cc_205 N_A_196_51#_M1007_g N_C_c_347_n 0.0193021f $X=2.42 $Y=0.865 $X2=0 $Y2=0
cc_206 N_A_196_51#_M1007_g N_C_c_348_n 0.018227f $X=2.42 $Y=0.865 $X2=0 $Y2=0
cc_207 N_A_196_51#_c_266_n N_C_c_348_n 0.00140261f $X=2.51 $Y=0.38 $X2=0 $Y2=0
cc_208 N_A_196_51#_c_264_n N_A_344_131#_c_408_n 0.019181f $X=1.415 $Y=1.085
+ $X2=0 $Y2=0
cc_209 N_A_196_51#_c_265_n N_A_344_131#_c_408_n 0.0427339f $X=2.51 $Y=0.38 $X2=0
+ $Y2=0
cc_210 N_A_196_51#_c_267_n N_A_344_131#_c_408_n 0.0208497f $X=1.77 $Y=1.17 $X2=0
+ $Y2=0
cc_211 N_A_196_51#_M1007_g N_A_344_131#_c_409_n 0.00866863f $X=2.42 $Y=0.865
+ $X2=0 $Y2=0
cc_212 N_A_196_51#_c_264_n N_A_344_131#_c_409_n 0.00464822f $X=1.415 $Y=1.085
+ $X2=0 $Y2=0
cc_213 N_A_196_51#_c_267_n N_A_344_131#_c_409_n 0.0137322f $X=1.77 $Y=1.17 $X2=0
+ $Y2=0
cc_214 N_A_196_51#_c_269_n N_A_344_131#_c_409_n 0.0318791f $X=1.855 $Y=1.785
+ $X2=0 $Y2=0
cc_215 N_A_196_51#_M1007_g N_A_344_131#_c_414_n 0.00131565f $X=2.42 $Y=0.865
+ $X2=0 $Y2=0
cc_216 N_A_196_51#_c_273_n N_A_344_131#_c_414_n 0.00644078f $X=1.77 $Y=1.87
+ $X2=0 $Y2=0
cc_217 N_A_196_51#_M1007_g N_A_344_131#_c_415_n 0.0188948f $X=2.42 $Y=0.865
+ $X2=0 $Y2=0
cc_218 N_A_196_51#_c_273_n N_A_344_131#_c_420_n 0.00802274f $X=1.77 $Y=1.87
+ $X2=0 $Y2=0
cc_219 N_A_196_51#_c_269_n N_A_344_131#_c_420_n 0.00641961f $X=1.855 $Y=1.785
+ $X2=0 $Y2=0
cc_220 N_A_196_51#_c_272_n N_VPWR_c_483_n 0.0138111f $X=1.22 $Y=2.865 $X2=0
+ $Y2=0
cc_221 N_A_196_51#_M1007_g N_VPWR_c_484_n 5.14407e-19 $X=2.42 $Y=0.865 $X2=0
+ $Y2=0
cc_222 N_A_196_51#_c_272_n N_VPWR_c_484_n 0.0608512f $X=1.22 $Y=2.865 $X2=0
+ $Y2=0
cc_223 N_A_196_51#_c_273_n N_VPWR_c_484_n 0.0258815f $X=1.77 $Y=1.87 $X2=0 $Y2=0
cc_224 N_A_196_51#_M1007_g N_VPWR_c_485_n 0.00763203f $X=2.42 $Y=0.865 $X2=0
+ $Y2=0
cc_225 N_A_196_51#_M1007_g N_VPWR_c_481_n 0.00366023f $X=2.42 $Y=0.865 $X2=0
+ $Y2=0
cc_226 N_A_196_51#_c_272_n N_VPWR_c_481_n 0.00980511f $X=1.22 $Y=2.865 $X2=0
+ $Y2=0
cc_227 N_A_196_51#_c_266_n N_VGND_c_562_n 0.00612417f $X=2.51 $Y=0.38 $X2=0
+ $Y2=0
cc_228 N_A_196_51#_c_270_n N_VGND_c_562_n 0.109572f $X=1.5 $Y=0.435 $X2=0 $Y2=0
cc_229 N_A_196_51#_c_266_n N_VGND_c_564_n 0.00874097f $X=2.51 $Y=0.38 $X2=0
+ $Y2=0
cc_230 N_A_196_51#_c_270_n N_VGND_c_564_n 0.0625425f $X=1.5 $Y=0.435 $X2=0 $Y2=0
cc_231 N_C_M1001_g N_D_M1010_g 0.0264237f $X=2.89 $Y=2.175 $X2=0 $Y2=0
cc_232 C N_D_M1010_g 0.0185867f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_233 N_C_c_348_n N_D_M1010_g 0.0632312f $X=2.87 $Y=1.185 $X2=0 $Y2=0
cc_234 C N_A_344_131#_M1012_g 0.00121971f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_235 C N_A_344_131#_c_409_n 0.0345581f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_236 N_C_M1001_g N_A_344_131#_c_415_n 0.0151001f $X=2.89 $Y=2.175 $X2=0 $Y2=0
cc_237 C N_A_344_131#_c_415_n 0.0315447f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_238 N_C_c_347_n N_A_344_131#_c_415_n 0.00295182f $X=2.87 $Y=1.35 $X2=0 $Y2=0
cc_239 N_C_M1001_g N_A_344_131#_c_416_n 0.00138675f $X=2.89 $Y=2.175 $X2=0 $Y2=0
cc_240 C N_A_344_131#_c_417_n 0.00174113f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_241 C N_A_344_131#_c_410_n 0.00759618f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_242 C N_A_344_131#_c_411_n 4.83351e-19 $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_243 C N_A_344_131#_c_421_n 0.0216489f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_244 N_C_c_347_n N_A_344_131#_c_421_n 0.00134164f $X=2.87 $Y=1.35 $X2=0 $Y2=0
cc_245 N_C_M1001_g N_VPWR_c_485_n 0.00390786f $X=2.89 $Y=2.175 $X2=0 $Y2=0
cc_246 N_C_M1001_g N_VPWR_c_481_n 0.00389386f $X=2.89 $Y=2.175 $X2=0 $Y2=0
cc_247 C N_VGND_c_560_n 0.0153763f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_248 C N_VGND_c_562_n 0.00740976f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_249 N_C_c_348_n N_VGND_c_562_n 0.00315876f $X=2.87 $Y=1.185 $X2=0 $Y2=0
cc_250 C N_VGND_c_564_n 0.0165687f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_251 N_C_c_348_n N_VGND_c_564_n 0.0046122f $X=2.87 $Y=1.185 $X2=0 $Y2=0
cc_252 C A_499_131# 0.00964043f $X=3.035 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_253 C A_607_131# 0.00198184f $X=3.035 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_254 N_D_M1010_g N_A_344_131#_M1012_g 0.015856f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_255 N_D_M1010_g N_A_344_131#_M1011_g 0.0234046f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_256 N_D_M1010_g N_A_344_131#_c_416_n 0.00249778f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_257 D N_A_344_131#_c_416_n 0.0128016f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_258 N_D_c_383_n N_A_344_131#_c_416_n 0.00109632f $X=3.32 $Y=2.92 $X2=0 $Y2=0
cc_259 N_D_M1010_g N_A_344_131#_c_417_n 0.0194659f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_260 N_D_M1010_g N_A_344_131#_c_410_n 0.00229257f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_261 N_D_M1010_g N_A_344_131#_c_411_n 0.0203042f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_262 N_D_M1010_g N_VPWR_c_485_n 0.00394549f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_263 D N_VPWR_c_485_n 0.0377148f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_264 N_D_c_383_n N_VPWR_c_485_n 0.00257728f $X=3.32 $Y=2.92 $X2=0 $Y2=0
cc_265 N_D_M1010_g N_VPWR_c_486_n 0.0100111f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_266 D N_VPWR_c_486_n 0.0342813f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_267 D N_VPWR_c_489_n 0.0237895f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_268 N_D_c_383_n N_VPWR_c_489_n 0.00724997f $X=3.32 $Y=2.92 $X2=0 $Y2=0
cc_269 D N_VPWR_c_481_n 0.0122685f $X=3.035 $Y=2.69 $X2=0 $Y2=0
cc_270 N_D_c_383_n N_VPWR_c_481_n 0.0128422f $X=3.32 $Y=2.92 $X2=0 $Y2=0
cc_271 N_D_M1010_g N_VGND_c_560_n 0.00432875f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_272 N_D_M1010_g N_VGND_c_562_n 0.0038866f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_273 N_D_M1010_g N_VGND_c_564_n 0.0046122f $X=3.32 $Y=0.865 $X2=0 $Y2=0
cc_274 N_A_344_131#_c_417_n N_VPWR_M1008_d 0.00224329f $X=3.605 $Y=1.79 $X2=0
+ $Y2=0
cc_275 N_A_344_131#_c_415_n N_VPWR_c_485_n 0.0219498f $X=2.985 $Y=1.79 $X2=0
+ $Y2=0
cc_276 N_A_344_131#_M1011_g N_VPWR_c_486_n 0.00699041f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_277 N_A_344_131#_c_417_n N_VPWR_c_532_n 0.0233069f $X=3.605 $Y=1.79 $X2=0
+ $Y2=0
cc_278 N_A_344_131#_c_411_n N_VPWR_c_532_n 6.53598e-19 $X=3.77 $Y=1.51 $X2=0
+ $Y2=0
cc_279 N_A_344_131#_M1011_g N_VPWR_c_490_n 0.00585385f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_280 N_A_344_131#_M1011_g N_VPWR_c_481_n 0.0127684f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_281 N_A_344_131#_M1012_g N_X_c_539_n 0.00937997f $X=3.845 $Y=0.655 $X2=0
+ $Y2=0
cc_282 N_A_344_131#_M1011_g N_X_c_539_n 0.00959542f $X=3.845 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_A_344_131#_c_417_n N_X_c_539_n 0.0137394f $X=3.605 $Y=1.79 $X2=0 $Y2=0
cc_284 N_A_344_131#_c_410_n N_X_c_539_n 0.0268611f $X=3.77 $Y=1.51 $X2=0 $Y2=0
cc_285 N_A_344_131#_c_411_n N_X_c_539_n 0.00817612f $X=3.77 $Y=1.51 $X2=0 $Y2=0
cc_286 N_A_344_131#_M1012_g X 0.0029015f $X=3.845 $Y=0.655 $X2=0 $Y2=0
cc_287 N_A_344_131#_c_411_n X 3.6706e-19 $X=3.77 $Y=1.51 $X2=0 $Y2=0
cc_288 N_A_344_131#_M1012_g N_VGND_c_560_n 0.00802989f $X=3.845 $Y=0.655 $X2=0
+ $Y2=0
cc_289 N_A_344_131#_c_417_n N_VGND_c_560_n 0.00583569f $X=3.605 $Y=1.79 $X2=0
+ $Y2=0
cc_290 N_A_344_131#_c_410_n N_VGND_c_560_n 0.00969967f $X=3.77 $Y=1.51 $X2=0
+ $Y2=0
cc_291 N_A_344_131#_c_411_n N_VGND_c_560_n 0.00111769f $X=3.77 $Y=1.51 $X2=0
+ $Y2=0
cc_292 N_A_344_131#_M1012_g N_VGND_c_563_n 0.00585385f $X=3.845 $Y=0.655 $X2=0
+ $Y2=0
cc_293 N_A_344_131#_M1012_g N_VGND_c_564_n 0.0127684f $X=3.845 $Y=0.655 $X2=0
+ $Y2=0
cc_294 N_A_344_131#_c_408_n A_427_131# 0.00103069f $X=2.11 $Y=0.795 $X2=-0.19
+ $Y2=-0.245
cc_295 N_VPWR_c_481_n N_X_M1011_d 0.00232552f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_296 N_VPWR_c_490_n N_X_c_543_n 0.0199472f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_297 N_VPWR_c_481_n N_X_c_543_n 0.0119743f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_298 X N_VGND_c_560_n 0.00156984f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_299 N_X_c_541_n N_VGND_c_563_n 0.0199472f $X=4.06 $Y=0.42 $X2=0 $Y2=0
cc_300 N_X_M1012_d N_VGND_c_564_n 0.00232552f $X=3.92 $Y=0.235 $X2=0 $Y2=0
cc_301 N_X_c_541_n N_VGND_c_564_n 0.0119743f $X=4.06 $Y=0.42 $X2=0 $Y2=0
