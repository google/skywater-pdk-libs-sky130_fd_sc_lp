* File: sky130_fd_sc_lp__nand4_4.pex.spice
* Created: Fri Aug 28 10:51:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4_4%D 3 7 11 15 19 23 27 31 33 34 35 36 55
c74 36 0 5.72698e-20 $X=1.68 $Y=1.665
c75 27 0 5.09472e-20 $X=1.765 $Y=0.745
r76 55 56 7.4613 $w=3.23e-07 $l=5e-08 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.815 $Y2=1.51
r77 53 55 26.8607 $w=3.23e-07 $l=1.8e-07 $layer=POLY_cond $X=1.585 $Y=1.51
+ $X2=1.765 $Y2=1.51
r78 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=1.51 $X2=1.585 $Y2=1.51
r79 51 53 29.8452 $w=3.23e-07 $l=2e-07 $layer=POLY_cond $X=1.385 $Y=1.51
+ $X2=1.585 $Y2=1.51
r80 50 51 7.4613 $w=3.23e-07 $l=5e-08 $layer=POLY_cond $X=1.335 $Y=1.51
+ $X2=1.385 $Y2=1.51
r81 49 54 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.245 $Y=1.587
+ $X2=1.585 $Y2=1.587
r82 48 50 13.4303 $w=3.23e-07 $l=9e-08 $layer=POLY_cond $X=1.245 $Y=1.51
+ $X2=1.335 $Y2=1.51
r83 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.245
+ $Y=1.51 $X2=1.245 $Y2=1.51
r84 46 48 43.2755 $w=3.23e-07 $l=2.9e-07 $layer=POLY_cond $X=0.955 $Y=1.51
+ $X2=1.245 $Y2=1.51
r85 44 46 7.4613 $w=3.23e-07 $l=5e-08 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=0.955 $Y2=1.51
r86 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.905
+ $Y=1.51 $X2=0.905 $Y2=1.51
r87 42 44 56.7059 $w=3.23e-07 $l=3.8e-07 $layer=POLY_cond $X=0.525 $Y=1.51
+ $X2=0.905 $Y2=1.51
r88 41 42 7.4613 $w=3.23e-07 $l=5e-08 $layer=POLY_cond $X=0.475 $Y=1.51
+ $X2=0.525 $Y2=1.51
r89 36 54 3.36868 $w=3.23e-07 $l=9.5e-08 $layer=LI1_cond $X=1.68 $Y=1.587
+ $X2=1.585 $Y2=1.587
r90 35 49 1.59569 $w=3.23e-07 $l=4.5e-08 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.245 $Y2=1.587
r91 35 45 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=0.905 $Y2=1.587
r92 34 45 6.56006 $w=3.23e-07 $l=1.85e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=0.905 $Y2=1.587
r93 33 34 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.587
+ $X2=0.72 $Y2=1.587
r94 29 56 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.675
+ $X2=1.815 $Y2=1.51
r95 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.815 $Y=1.675
+ $X2=1.815 $Y2=2.465
r96 25 55 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=1.51
r97 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=0.745
r98 21 51 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.675
+ $X2=1.385 $Y2=1.51
r99 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.385 $Y=1.675
+ $X2=1.385 $Y2=2.465
r100 17 50 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.345
+ $X2=1.335 $Y2=1.51
r101 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.335 $Y=1.345
+ $X2=1.335 $Y2=0.745
r102 13 46 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.675
+ $X2=0.955 $Y2=1.51
r103 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.955 $Y=1.675
+ $X2=0.955 $Y2=2.465
r104 9 44 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=1.51
r105 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=0.745
r106 5 42 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.675
+ $X2=0.525 $Y2=1.51
r107 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.525 $Y=1.675
+ $X2=0.525 $Y2=2.465
r108 1 41 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=1.51
r109 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.475 $Y=1.345 $X2=0.475
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_4%C 3 7 11 15 19 23 27 31 33 34 35 50 51 53
c94 51 0 1.74102e-19 $X=3.485 $Y=1.51
c95 27 0 2.40437e-20 $X=3.485 $Y=0.745
c96 7 0 1.91748e-19 $X=2.405 $Y=2.465
r97 49 51 31.4007 $w=3.07e-07 $l=2e-07 $layer=POLY_cond $X=3.285 $Y=1.51
+ $X2=3.485 $Y2=1.51
r98 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.285
+ $Y=1.51 $X2=3.285 $Y2=1.51
r99 47 49 3.14007 $w=3.07e-07 $l=2e-08 $layer=POLY_cond $X=3.265 $Y=1.51
+ $X2=3.285 $Y2=1.51
r100 46 47 32.9707 $w=3.07e-07 $l=2.1e-07 $layer=POLY_cond $X=3.055 $Y=1.51
+ $X2=3.265 $Y2=1.51
r101 45 46 34.5407 $w=3.07e-07 $l=2.2e-07 $layer=POLY_cond $X=2.835 $Y=1.51
+ $X2=3.055 $Y2=1.51
r102 44 45 32.9707 $w=3.07e-07 $l=2.1e-07 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.835 $Y2=1.51
r103 43 44 34.5407 $w=3.07e-07 $l=2.2e-07 $layer=POLY_cond $X=2.405 $Y=1.51
+ $X2=2.625 $Y2=1.51
r104 42 53 4.0014 $w=3.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.265 $Y=1.565
+ $X2=2.385 $Y2=1.565
r105 41 43 21.9805 $w=3.07e-07 $l=1.4e-07 $layer=POLY_cond $X=2.265 $Y=1.51
+ $X2=2.405 $Y2=1.51
r106 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.265
+ $Y=1.51 $X2=2.265 $Y2=1.51
r107 39 41 10.9902 $w=3.07e-07 $l=7e-08 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.265 $Y2=1.51
r108 35 50 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.285 $Y2=1.565
r109 34 35 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r110 34 53 7.94251 $w=3.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.385 $Y2=1.565
r111 33 42 3.64957 $w=3.51e-07 $l=1.05e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.265 $Y2=1.565
r112 29 51 32.9707 $w=3.07e-07 $l=2.80624e-07 $layer=POLY_cond $X=3.695 $Y=1.675
+ $X2=3.485 $Y2=1.51
r113 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.695 $Y=1.675
+ $X2=3.695 $Y2=2.465
r114 25 51 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.345
+ $X2=3.485 $Y2=1.51
r115 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.485 $Y=1.345
+ $X2=3.485 $Y2=0.745
r116 21 47 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.265 $Y=1.675
+ $X2=3.265 $Y2=1.51
r117 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.265 $Y=1.675
+ $X2=3.265 $Y2=2.465
r118 17 46 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.345
+ $X2=3.055 $Y2=1.51
r119 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.055 $Y=1.345
+ $X2=3.055 $Y2=0.745
r120 13 45 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.675
+ $X2=2.835 $Y2=1.51
r121 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.835 $Y=1.675
+ $X2=2.835 $Y2=2.465
r122 9 44 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=1.51
r123 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=0.745
r124 5 43 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.675
+ $X2=2.405 $Y2=1.51
r125 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.405 $Y=1.675
+ $X2=2.405 $Y2=2.465
r126 1 39 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=1.51
r127 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.195 $Y=1.345 $X2=2.195
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_4%B 3 7 11 15 19 23 27 31 33 34 35 36 60 61
c77 60 0 1.74102e-19 $X=5.845 $Y=1.51
r78 59 61 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.845 $Y=1.51
+ $X2=5.865 $Y2=1.51
r79 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.845
+ $Y=1.51 $X2=5.845 $Y2=1.51
r80 57 59 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=5.435 $Y=1.51
+ $X2=5.845 $Y2=1.51
r81 56 57 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.415 $Y=1.51
+ $X2=5.435 $Y2=1.51
r82 54 56 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.165 $Y=1.51
+ $X2=5.415 $Y2=1.51
r83 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.165
+ $Y=1.51 $X2=5.165 $Y2=1.51
r84 52 54 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.005 $Y=1.51
+ $X2=5.165 $Y2=1.51
r85 51 52 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.985 $Y=1.51
+ $X2=5.005 $Y2=1.51
r86 49 51 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=4.825 $Y=1.51
+ $X2=4.985 $Y2=1.51
r87 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.825
+ $Y=1.51 $X2=4.825 $Y2=1.51
r88 47 49 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=4.575 $Y=1.51
+ $X2=4.825 $Y2=1.51
r89 46 47 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.555 $Y=1.51
+ $X2=4.575 $Y2=1.51
r90 44 46 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.485 $Y=1.51
+ $X2=4.555 $Y2=1.51
r91 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.485
+ $Y=1.51 $X2=4.485 $Y2=1.51
r92 41 44 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.125 $Y=1.51
+ $X2=4.485 $Y2=1.51
r93 36 60 11.5244 $w=3.23e-07 $l=3.25e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.845 $Y2=1.587
r94 36 55 12.5882 $w=3.23e-07 $l=3.55e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.165 $Y2=1.587
r95 35 55 4.43247 $w=3.23e-07 $l=1.25e-07 $layer=LI1_cond $X=5.04 $Y=1.587
+ $X2=5.165 $Y2=1.587
r96 35 50 7.62385 $w=3.23e-07 $l=2.15e-07 $layer=LI1_cond $X=5.04 $Y=1.587
+ $X2=4.825 $Y2=1.587
r97 34 50 9.39684 $w=3.23e-07 $l=2.65e-07 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.825 $Y2=1.587
r98 34 45 2.65948 $w=3.23e-07 $l=7.5e-08 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.485 $Y2=1.587
r99 33 45 14.3612 $w=3.23e-07 $l=4.05e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.485 $Y2=1.587
r100 29 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.865 $Y=1.345
+ $X2=5.865 $Y2=1.51
r101 29 31 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.865 $Y=1.345
+ $X2=5.865 $Y2=0.755
r102 25 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.435 $Y=1.345
+ $X2=5.435 $Y2=1.51
r103 25 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.435 $Y=1.345
+ $X2=5.435 $Y2=0.755
r104 21 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.415 $Y=1.675
+ $X2=5.415 $Y2=1.51
r105 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.415 $Y=1.675
+ $X2=5.415 $Y2=2.465
r106 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.005 $Y=1.345
+ $X2=5.005 $Y2=1.51
r107 17 19 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.005 $Y=1.345
+ $X2=5.005 $Y2=0.755
r108 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.675
+ $X2=4.985 $Y2=1.51
r109 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.985 $Y=1.675
+ $X2=4.985 $Y2=2.465
r110 9 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.575 $Y=1.345
+ $X2=4.575 $Y2=1.51
r111 9 11 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.575 $Y=1.345
+ $X2=4.575 $Y2=0.755
r112 5 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.555 $Y=1.675
+ $X2=4.555 $Y2=1.51
r113 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.555 $Y=1.675
+ $X2=4.555 $Y2=2.465
r114 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.125 $Y=1.675
+ $X2=4.125 $Y2=1.51
r115 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.125 $Y=1.675
+ $X2=4.125 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_4%A 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 43
r77 45 46 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=7.745
+ $Y=1.51 $X2=7.745 $Y2=1.51
r78 43 45 20.7312 $w=3.72e-07 $l=1.6e-07 $layer=POLY_cond $X=7.585 $Y=1.535
+ $X2=7.745 $Y2=1.535
r79 42 43 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=7.155 $Y=1.535
+ $X2=7.585 $Y2=1.535
r80 41 42 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=6.725 $Y=1.535
+ $X2=7.155 $Y2=1.535
r81 39 41 44.0538 $w=3.72e-07 $l=3.4e-07 $layer=POLY_cond $X=6.385 $Y=1.535
+ $X2=6.725 $Y2=1.535
r82 39 40 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.385
+ $Y=1.51 $X2=6.385 $Y2=1.51
r83 37 39 11.6613 $w=3.72e-07 $l=9e-08 $layer=POLY_cond $X=6.295 $Y=1.535
+ $X2=6.385 $Y2=1.535
r84 32 46 6.20546 $w=3.23e-07 $l=1.75e-07 $layer=LI1_cond $X=7.92 $Y=1.587
+ $X2=7.745 $Y2=1.587
r85 31 46 10.8152 $w=3.23e-07 $l=3.05e-07 $layer=LI1_cond $X=7.44 $Y=1.587
+ $X2=7.745 $Y2=1.587
r86 30 31 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.587
+ $X2=7.44 $Y2=1.587
r87 29 30 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.587
+ $X2=6.96 $Y2=1.587
r88 29 40 3.36868 $w=3.23e-07 $l=9.5e-08 $layer=LI1_cond $X=6.48 $Y=1.587
+ $X2=6.385 $Y2=1.587
r89 26 43 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.585 $Y=1.725
+ $X2=7.585 $Y2=1.535
r90 26 28 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.585 $Y=1.725
+ $X2=7.585 $Y2=2.465
r91 22 43 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.585 $Y=1.345
+ $X2=7.585 $Y2=1.535
r92 22 24 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=7.585 $Y=1.345
+ $X2=7.585 $Y2=0.755
r93 19 42 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.155 $Y=1.725
+ $X2=7.155 $Y2=1.535
r94 19 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.155 $Y=1.725
+ $X2=7.155 $Y2=2.465
r95 15 42 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.155 $Y=1.345
+ $X2=7.155 $Y2=1.535
r96 15 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=7.155 $Y=1.345
+ $X2=7.155 $Y2=0.755
r97 12 41 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.725 $Y=1.725
+ $X2=6.725 $Y2=1.535
r98 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.725 $Y=1.725
+ $X2=6.725 $Y2=2.465
r99 8 41 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.725 $Y=1.345
+ $X2=6.725 $Y2=1.535
r100 8 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.725 $Y=1.345
+ $X2=6.725 $Y2=0.755
r101 5 37 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.295 $Y=1.725
+ $X2=6.295 $Y2=1.535
r102 5 7 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.295 $Y=1.725
+ $X2=6.295 $Y2=2.465
r103 1 37 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.295 $Y=1.345
+ $X2=6.295 $Y2=1.535
r104 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.295 $Y=1.345
+ $X2=6.295 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 40 44 48 52
+ 54 58 62 64 66 71 72 73 74 75 77 82 87 99 104 113 116 119 122 127 131
r130 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r132 123 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r133 122 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r134 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r135 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r136 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 108 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r140 108 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r141 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r142 105 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.105 $Y=3.33
+ $X2=6.94 $Y2=3.33
r143 105 107 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.105 $Y=3.33
+ $X2=7.44 $Y2=3.33
r144 104 130 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=7.635 $Y=3.33
+ $X2=7.897 $Y2=3.33
r145 104 107 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.635 $Y=3.33
+ $X2=7.44 $Y2=3.33
r146 103 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r147 103 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r148 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r149 100 122 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=6.245 $Y=3.33
+ $X2=5.855 $Y2=3.33
r150 100 102 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.245 $Y=3.33
+ $X2=6.48 $Y2=3.33
r151 99 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=3.33
+ $X2=6.94 $Y2=3.33
r152 99 102 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.775 $Y=3.33
+ $X2=6.48 $Y2=3.33
r153 98 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r154 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r155 95 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r156 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r157 92 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=3.33
+ $X2=3.05 $Y2=3.33
r158 92 94 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=3.33
+ $X2=3.6 $Y2=3.33
r159 91 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r160 91 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r161 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r162 88 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.11 $Y2=3.33
r163 88 90 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.64 $Y2=3.33
r164 87 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=3.33
+ $X2=3.05 $Y2=3.33
r165 87 90 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.885 $Y=3.33
+ $X2=2.64 $Y2=3.33
r166 86 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r167 86 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r169 83 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r170 83 85 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r171 82 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=2.11 $Y2=3.33
r172 82 85 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=1.68 $Y2=3.33
r173 81 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r174 81 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r175 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r176 78 110 4.36354 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.22 $Y2=3.33
r177 78 80 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r178 77 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r179 77 80 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r180 75 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r181 75 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r182 73 97 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.56 $Y2=3.33
r183 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.77 $Y2=3.33
r184 71 94 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.6 $Y2=3.33
r185 71 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.91 $Y2=3.33
r186 70 97 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=4.56 $Y2=3.33
r187 70 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=3.91 $Y2=3.33
r188 66 69 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=7.8 $Y=2.01 $X2=7.8
+ $Y2=2.95
r189 64 130 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=7.8 $Y=3.245
+ $X2=7.897 $Y2=3.33
r190 64 69 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.8 $Y=3.245
+ $X2=7.8 $Y2=2.95
r191 60 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.94 $Y=3.245
+ $X2=6.94 $Y2=3.33
r192 60 62 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=6.94 $Y=3.245
+ $X2=6.94 $Y2=2.36
r193 56 122 3.08259 $w=7.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.855 $Y=3.245
+ $X2=5.855 $Y2=3.33
r194 56 58 13.5709 $w=7.78e-07 $l=8.85e-07 $layer=LI1_cond $X=5.855 $Y=3.245
+ $X2=5.855 $Y2=2.36
r195 55 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=4.77 $Y2=3.33
r196 54 122 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=5.465 $Y=3.33
+ $X2=5.855 $Y2=3.33
r197 54 55 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.465 $Y=3.33
+ $X2=4.935 $Y2=3.33
r198 50 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=3.33
r199 50 52 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=2.36
r200 46 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=3.245
+ $X2=3.91 $Y2=3.33
r201 46 48 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=3.91 $Y=3.245
+ $X2=3.91 $Y2=2.36
r202 42 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=3.245
+ $X2=3.05 $Y2=3.33
r203 42 44 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=3.05 $Y=3.245
+ $X2=3.05 $Y2=2.36
r204 38 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.11 $Y2=3.33
r205 38 40 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.11 $Y2=2.36
r206 34 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r207 34 36 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.39
r208 30 33 33.792 $w=2.93e-07 $l=8.65e-07 $layer=LI1_cond $X=0.292 $Y=2.085
+ $X2=0.292 $Y2=2.95
r209 28 110 3.11398 $w=2.95e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.292 $Y=3.245
+ $X2=0.22 $Y2=3.33
r210 28 33 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.292 $Y=3.245
+ $X2=0.292 $Y2=2.95
r211 9 69 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.66
+ $Y=1.835 $X2=7.8 $Y2=2.95
r212 9 66 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=7.66
+ $Y=1.835 $X2=7.8 $Y2=2.01
r213 8 62 300 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_PDIFF $count=2 $X=6.8
+ $Y=1.835 $X2=6.94 $Y2=2.36
r214 7 58 150 $w=1.7e-07 $l=8.1108e-07 $layer=licon1_PDIFF $count=4 $X=5.49
+ $Y=1.835 $X2=6.08 $Y2=2.36
r215 6 52 300 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_PDIFF $count=2 $X=4.63
+ $Y=1.835 $X2=4.77 $Y2=2.36
r216 5 48 300 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_PDIFF $count=2 $X=3.77
+ $Y=1.835 $X2=3.91 $Y2=2.36
r217 4 44 300 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=1.835 $X2=3.05 $Y2=2.36
r218 3 40 300 $w=1.7e-07 $l=6.254e-07 $layer=licon1_PDIFF $count=2 $X=1.89
+ $Y=1.835 $X2=2.11 $Y2=2.36
r219 2 36 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.39
r220 1 33 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=2.95
r221 1 30 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 39 42 43 44 45
+ 46 49 51 55 57 61 65 67 69 73 75 77 79 81 86 88 89 91 94 95 96 103 109 114
c151 96 0 1.34478e-19 $X=1.68 $Y=2.035
r152 96 103 6.78838 $w=1.85e-07 $l=1.3e-07 $layer=LI1_cond $X=1.635 $Y=2.02
+ $X2=1.505 $Y2=2.02
r153 96 114 22.9606 $w=4.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.635 $Y=2.12
+ $X2=1.635 $Y2=2.91
r154 95 103 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=2.02
+ $X2=1.505 $Y2=2.02
r155 95 104 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=1.2 $Y=2.02
+ $X2=0.835 $Y2=2.02
r156 94 104 3.63256 $w=2e-07 $l=1.13e-07 $layer=LI1_cond $X=0.722 $Y=2.02
+ $X2=0.835 $Y2=2.02
r157 94 109 25.1657 $w=3.93e-07 $l=7.9e-07 $layer=LI1_cond $X=0.722 $Y=2.12
+ $X2=0.722 $Y2=2.91
r158 83 84 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.48 $Y=2.005
+ $X2=3.715 $Y2=2.005
r159 79 96 26.5861 $w=3.08e-07 $l=6.8e-07 $layer=LI1_cond $X=2.445 $Y=2.005
+ $X2=1.765 $Y2=2.005
r160 79 81 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.445 $Y=2.005
+ $X2=2.58 $Y2=2.005
r161 75 93 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.37 $Y=2.09
+ $X2=7.37 $Y2=2.005
r162 75 77 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=7.37 $Y=2.09
+ $X2=7.37 $Y2=2.91
r163 71 73 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=7.37 $Y=1.085
+ $X2=7.37 $Y2=0.71
r164 70 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=1.17
+ $X2=6.51 $Y2=1.17
r165 69 71 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.205 $Y=1.17
+ $X2=7.37 $Y2=1.085
r166 69 70 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.205 $Y=1.17
+ $X2=6.675 $Y2=1.17
r167 68 91 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.605 $Y=2.005
+ $X2=6.51 $Y2=2.005
r168 67 93 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.275 $Y=2.005
+ $X2=7.37 $Y2=2.005
r169 67 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.275 $Y=2.005
+ $X2=6.605 $Y2=2.005
r170 63 91 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.51 $Y=2.09
+ $X2=6.51 $Y2=2.005
r171 63 65 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=6.51 $Y=2.09
+ $X2=6.51 $Y2=2.91
r172 59 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.51 $Y=1.085
+ $X2=6.51 $Y2=1.17
r173 59 61 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=6.51 $Y=1.085
+ $X2=6.51 $Y2=0.71
r174 58 88 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.295 $Y=2.005
+ $X2=5.2 $Y2=2.005
r175 57 91 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.415 $Y=2.005
+ $X2=6.51 $Y2=2.005
r176 57 58 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=6.415 $Y=2.005
+ $X2=5.295 $Y2=2.005
r177 53 88 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.2 $Y=2.09 $X2=5.2
+ $Y2=2.005
r178 53 55 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=5.2 $Y=2.09 $X2=5.2
+ $Y2=2.91
r179 52 86 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.435 $Y=2.005
+ $X2=4.34 $Y2=2.005
r180 51 88 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.105 $Y=2.005
+ $X2=5.2 $Y2=2.005
r181 51 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.105 $Y=2.005
+ $X2=4.435 $Y2=2.005
r182 47 86 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=2.09
+ $X2=4.34 $Y2=2.005
r183 47 49 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=4.34 $Y=2.09
+ $X2=4.34 $Y2=2.91
r184 46 84 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=2.005
+ $X2=3.715 $Y2=2.005
r185 45 86 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.245 $Y=2.005
+ $X2=4.34 $Y2=2.005
r186 45 46 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=4.245 $Y=2.005
+ $X2=3.8 $Y2=2.005
r187 43 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.345 $Y=1.17
+ $X2=6.51 $Y2=1.17
r188 43 44 166.037 $w=1.68e-07 $l=2.545e-06 $layer=LI1_cond $X=6.345 $Y=1.17
+ $X2=3.8 $Y2=1.17
r189 42 84 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=1.92
+ $X2=3.715 $Y2=2.005
r190 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.715 $Y=1.255
+ $X2=3.8 $Y2=1.17
r191 41 42 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.715 $Y=1.255
+ $X2=3.715 $Y2=1.92
r192 37 83 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=2.09
+ $X2=3.48 $Y2=2.005
r193 37 39 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=3.48 $Y=2.09
+ $X2=3.48 $Y2=2.91
r194 36 81 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.715 $Y=2.005
+ $X2=2.58 $Y2=2.005
r195 35 83 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.385 $Y=2.005
+ $X2=3.48 $Y2=2.005
r196 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.385 $Y=2.005
+ $X2=2.715 $Y2=2.005
r197 31 81 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=2.09
+ $X2=2.58 $Y2=2.005
r198 31 33 35.0001 $w=2.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.58 $Y=2.09
+ $X2=2.58 $Y2=2.91
r199 10 93 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.835 $X2=7.37 $Y2=2.085
r200 10 77 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.835 $X2=7.37 $Y2=2.91
r201 9 91 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=6.37
+ $Y=1.835 $X2=6.51 $Y2=2.085
r202 9 65 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.37
+ $Y=1.835 $X2=6.51 $Y2=2.91
r203 8 88 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=5.06
+ $Y=1.835 $X2=5.2 $Y2=2.085
r204 8 55 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.06
+ $Y=1.835 $X2=5.2 $Y2=2.91
r205 7 86 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=4.2
+ $Y=1.835 $X2=4.34 $Y2=2.085
r206 7 49 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.2
+ $Y=1.835 $X2=4.34 $Y2=2.91
r207 6 83 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=1.835 $X2=3.48 $Y2=2.085
r208 6 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.34
+ $Y=1.835 $X2=3.48 $Y2=2.91
r209 5 81 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2.085
r210 5 33 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2.91
r211 4 96 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.085
r212 4 114 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.91
r213 3 94 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.74 $Y2=2.085
r214 3 109 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.74 $Y2=2.91
r215 2 73 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=7.23
+ $Y=0.335 $X2=7.37 $Y2=0.71
r216 1 61 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=6.37
+ $Y=0.335 $X2=6.51 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_4%A_27_65# 1 2 3 4 5 18 20 21 24 26 32 33 36
+ 38 40 41 42
r71 42 45 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.78 $Y=0.35 $X2=3.78
+ $Y2=0.45
r72 39 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.935 $Y=0.35
+ $X2=2.84 $Y2=0.35
r73 38 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0.35
+ $X2=3.78 $Y2=0.35
r74 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.615 $Y=0.35
+ $X2=2.935 $Y2=0.35
r75 34 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.435
+ $X2=2.84 $Y2=0.35
r76 34 36 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=2.84 $Y=0.435
+ $X2=2.84 $Y2=0.7
r77 32 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.745 $Y=0.35
+ $X2=2.84 $Y2=0.35
r78 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.745 $Y=0.35
+ $X2=2.075 $Y2=0.35
r79 29 31 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=1.98 $Y=1.085
+ $X2=1.98 $Y2=0.45
r80 28 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.98 $Y=0.435
+ $X2=2.075 $Y2=0.35
r81 28 31 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=1.98 $Y=0.435
+ $X2=1.98 $Y2=0.45
r82 27 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.215 $Y=1.17
+ $X2=1.12 $Y2=1.17
r83 26 29 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.885 $Y=1.17
+ $X2=1.98 $Y2=1.085
r84 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.885 $Y=1.17
+ $X2=1.215 $Y2=1.17
r85 22 40 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=1.085
+ $X2=1.12 $Y2=1.17
r86 22 24 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=1.12 $Y=1.085
+ $X2=1.12 $Y2=0.47
r87 20 40 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.025 $Y=1.17
+ $X2=1.12 $Y2=1.17
r88 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=1.17
+ $X2=0.355 $Y2=1.17
r89 16 21 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.255 $Y=1.085
+ $X2=0.355 $Y2=1.17
r90 16 18 34.1045 $w=1.98e-07 $l=6.15e-07 $layer=LI1_cond $X=0.255 $Y=1.085
+ $X2=0.255 $Y2=0.47
r91 5 45 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.325 $X2=3.78 $Y2=0.45
r92 4 36 182 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.325 $X2=2.84 $Y2=0.7
r93 3 31 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.325 $X2=1.98 $Y2=0.45
r94 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.325 $X2=1.12 $Y2=0.47
r95 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.325 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_4%VGND 1 2 9 13 15 17 22 29 30 33 36
r81 36 37 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r82 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r83 29 30 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r84 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=0 $X2=1.55
+ $Y2=0
r85 27 29 404.818 $w=1.68e-07 $l=6.205e-06 $layer=LI1_cond $X=1.715 $Y=0
+ $X2=7.92 $Y2=0
r86 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r87 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r88 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r89 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r90 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r91 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.55
+ $Y2=0
r92 22 25 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.2
+ $Y2=0
r93 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r94 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r95 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r96 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r97 15 30 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=7.92
+ $Y2=0
r98 15 37 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=1.68
+ $Y2=0
r99 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0
r100 11 13 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0.45
r101 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r102 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.45
r103 2 13 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.325 $X2=1.55 $Y2=0.45
r104 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.325 $X2=0.69 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_4%A_454_65# 1 2 3 4 15 17 18 23 26
c52 18 0 5.09472e-20 $X=2.575 $Y=1.12
c53 17 0 2.40437e-20 $X=3.105 $Y=1.12
r54 28 29 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.27 $Y=0.83
+ $X2=3.27 $Y2=1.12
r55 26 28 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.27 $Y=0.69
+ $X2=3.27 $Y2=0.83
r56 21 23 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=4.79 $Y=0.83 $X2=5.65
+ $Y2=0.83
r57 19 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0.83
+ $X2=3.27 $Y2=0.83
r58 19 21 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=3.435 $Y=0.83
+ $X2=4.79 $Y2=0.83
r59 17 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=1.12
+ $X2=3.27 $Y2=1.12
r60 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.105 $Y=1.12
+ $X2=2.575 $Y2=1.12
r61 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.41 $Y=1.035
+ $X2=2.575 $Y2=1.12
r62 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.41 $Y=1.035
+ $X2=2.41 $Y2=0.69
r63 4 23 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=5.51
+ $Y=0.335 $X2=5.65 $Y2=0.83
r64 3 21 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=4.65
+ $Y=0.335 $X2=4.79 $Y2=0.83
r65 2 26 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.325 $X2=3.27 $Y2=0.69
r66 1 15 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.325 $X2=2.41 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_4%A_843_67# 1 2 3 4 5 16 24 26 30 32 36 38 39
r49 34 36 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=7.835 $Y=0.445
+ $X2=7.835 $Y2=0.48
r50 33 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.035 $Y=0.36
+ $X2=6.94 $Y2=0.36
r51 32 34 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.705 $Y=0.36
+ $X2=7.835 $Y2=0.445
r52 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.705 $Y=0.36
+ $X2=7.035 $Y2=0.36
r53 28 39 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.94 $Y=0.445
+ $X2=6.94 $Y2=0.36
r54 28 30 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=6.94 $Y=0.445
+ $X2=6.94 $Y2=0.75
r55 27 38 4.31353 $w=2.35e-07 $l=1.23288e-07 $layer=LI1_cond $X=6.175 $Y=0.36
+ $X2=6.08 $Y2=0.425
r56 26 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.845 $Y=0.36
+ $X2=6.94 $Y2=0.36
r57 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.845 $Y=0.36
+ $X2=6.175 $Y2=0.36
r58 22 38 2.11804 $w=1.9e-07 $l=1.5e-07 $layer=LI1_cond $X=6.08 $Y=0.575
+ $X2=6.08 $Y2=0.425
r59 22 24 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=6.08 $Y=0.575
+ $X2=6.08 $Y2=0.75
r60 18 21 33.0367 $w=2.98e-07 $l=8.6e-07 $layer=LI1_cond $X=4.36 $Y=0.425
+ $X2=5.22 $Y2=0.425
r61 16 38 4.31353 $w=2.35e-07 $l=9.5e-08 $layer=LI1_cond $X=5.985 $Y=0.425
+ $X2=6.08 $Y2=0.425
r62 16 21 29.3873 $w=2.98e-07 $l=7.65e-07 $layer=LI1_cond $X=5.985 $Y=0.425
+ $X2=5.22 $Y2=0.425
r63 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.66
+ $Y=0.335 $X2=7.8 $Y2=0.48
r64 4 30 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=6.8
+ $Y=0.335 $X2=6.94 $Y2=0.75
r65 3 24 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=5.94
+ $Y=0.335 $X2=6.08 $Y2=0.75
r66 2 21 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.08
+ $Y=0.335 $X2=5.22 $Y2=0.46
r67 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.215
+ $Y=0.335 $X2=4.36 $Y2=0.46
.ends

