* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__srsdfrtn_1 CLK_N D RESET_B SCD SCE SLEEP_B KAPWR VGND VNB
+ VPB VPWR Q
M1000 a_1041_419# a_742_63# a_305_97# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=4.078e+11p ps=3.91e+06u
M1001 VGND SCE a_27_55# VNB nshort w=420000u l=150000u
+  ad=1.322e+12p pd=1.296e+07u as=1.155e+11p ps=1.39e+06u
M1002 a_2951_99# a_666_89# a_2879_99# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_469_97# a_27_55# a_391_97# VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=1.008e+11p ps=1.32e+06u
M1004 a_411_491# a_27_55# a_305_97# VPB phighvt w=640000u l=150000u
+  ad=3.136e+11p pd=2.26e+06u as=0p ps=0u
M1005 a_2999_73# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.4703e+12p ps=1.248e+07u
M1006 a_2480_97# SLEEP_B VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 a_1453_77# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=2.331e+11p pd=2.79e+06u as=0p ps=0u
M1008 a_3115_99# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 a_2999_73# a_2717_427# a_3115_99# VNB nshort w=420000u l=150000u
+  ad=1.68e+11p pd=1.64e+06u as=0p ps=0u
M1010 KAPWR a_1343_51# a_1242_419# VPB phighvt w=1e+06u l=250000u
+  ad=1.68302e+12p pd=1.137e+07u as=5.15e+11p ps=3.03e+06u
M1011 a_1682_341# RESET_B a_1113_419# VPB phighvt w=1e+06u l=250000u
+  ad=2.1e+11p pd=2.42e+06u as=5.962e+11p ps=5.32e+06u
M1012 a_1373_77# a_1343_51# a_1009_107# VNB nshort w=420000u l=150000u
+  ad=1.05e+11p pd=1.34e+06u as=4.293e+11p ps=4.11e+06u
M1013 a_2879_99# a_666_89# a_2717_427# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.51e+11p ps=2.14e+06u
M1014 KAPWR a_1724_21# a_1682_341# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1343_51# a_666_89# a_2717_427# VPB phighvt w=840000u l=150000u
+  ad=8.3315e+11p pd=5.66e+06u as=2.688e+11p ps=2.43e+06u
M1016 VPWR SCE a_27_55# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1017 a_1724_21# SLEEP_B KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.65e+11p pd=2.53e+06u as=0p ps=0u
M1018 VGND a_742_63# a_666_89# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.513e+11p ps=3.02e+06u
M1019 KAPWR SLEEP_B a_742_63# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1020 a_1724_21# SLEEP_B a_2480_97# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1021 VPWR a_742_63# a_666_89# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1022 a_220_97# SCD a_469_97# VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=0p ps=0u
M1023 a_305_97# SCE a_220_97# VNB nshort w=420000u l=150000u
+  ad=2.331e+11p pd=2.79e+06u as=0p ps=0u
M1024 Q a_3368_57# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.465e+11p pd=3.07e+06u as=0p ps=0u
M1025 a_247_491# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1026 a_305_97# D a_247_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_1724_21# a_1453_77# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_469_97# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1343_51# a_1113_419# KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_2717_427# a_742_63# a_2645_427# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1031 VPWR a_2999_73# a_2562_427# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.31e+11p ps=2.78e+06u
M1032 a_1343_51# a_1113_419# a_1840_47# VNB nshort w=420000u l=150000u
+  ad=3.245e+11p pd=3.33e+06u as=8.82e+10p ps=1.26e+06u
M1033 Q a_3368_57# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1034 a_305_97# a_666_89# a_1201_215# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1035 a_1453_77# a_1343_51# a_1373_77# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND a_2717_427# a_3368_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1037 a_1113_419# a_742_63# a_1041_419# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_2198_97# CLK_N a_742_63# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.666e+11p ps=2.32e+06u
M1039 a_2276_97# SLEEP_B a_2198_97# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1040 a_391_97# D a_305_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1113_419# a_742_63# a_1009_107# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1042 a_742_63# CLK_N KAPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND SLEEP_B a_2276_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_2717_427# a_742_63# a_1343_51# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_1201_215# a_666_89# a_1113_419# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 VPWR a_2717_427# a_2999_73# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR a_2717_427# a_3368_57# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1048 a_1840_47# a_1113_419# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 a_305_97# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_2645_427# a_742_63# a_2562_427# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 VGND a_2999_73# a_2951_99# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1052 VPWR SCD a_411_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1053 a_1242_419# a_666_89# a_1113_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends
