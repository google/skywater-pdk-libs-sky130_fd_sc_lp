* File: sky130_fd_sc_lp__a21bo_lp.pxi.spice
* Created: Fri Aug 28 09:49:30 2020
* 
x_PM_SKY130_FD_SC_LP__A21BO_LP%A_84_29# N_A_84_29#_M1009_d N_A_84_29#_M1006_d
+ N_A_84_29#_M1007_g N_A_84_29#_c_82_n N_A_84_29#_M1004_g N_A_84_29#_M1001_g
+ N_A_84_29#_c_85_n N_A_84_29#_c_144_p N_A_84_29#_c_86_n N_A_84_29#_c_87_n
+ N_A_84_29#_c_88_n N_A_84_29#_c_94_n N_A_84_29#_c_140_p N_A_84_29#_c_89_n
+ N_A_84_29#_c_95_n N_A_84_29#_c_90_n N_A_84_29#_c_91_n
+ PM_SKY130_FD_SC_LP__A21BO_LP%A_84_29#
x_PM_SKY130_FD_SC_LP__A21BO_LP%A2 N_A2_M1011_g N_A2_M1008_g N_A2_c_176_n
+ N_A2_c_177_n A2 N_A2_c_178_n N_A2_c_179_n N_A2_c_180_n
+ PM_SKY130_FD_SC_LP__A21BO_LP%A2
x_PM_SKY130_FD_SC_LP__A21BO_LP%A1 N_A1_M1009_g N_A1_M1010_g N_A1_c_224_n
+ N_A1_c_225_n A1 N_A1_c_226_n N_A1_c_227_n N_A1_c_228_n
+ PM_SKY130_FD_SC_LP__A21BO_LP%A1
x_PM_SKY130_FD_SC_LP__A21BO_LP%A_308_364# N_A_308_364#_M1003_d
+ N_A_308_364#_M1005_d N_A_308_364#_c_293_n N_A_308_364#_M1006_g
+ N_A_308_364#_c_294_n N_A_308_364#_c_295_n N_A_308_364#_c_284_n
+ N_A_308_364#_M1000_g N_A_308_364#_c_285_n N_A_308_364#_c_286_n
+ N_A_308_364#_M1012_g N_A_308_364#_c_287_n N_A_308_364#_c_288_n
+ N_A_308_364#_c_297_n N_A_308_364#_c_289_n N_A_308_364#_c_290_n
+ N_A_308_364#_c_291_n N_A_308_364#_c_292_n
+ PM_SKY130_FD_SC_LP__A21BO_LP%A_308_364#
x_PM_SKY130_FD_SC_LP__A21BO_LP%B1_N N_B1_N_M1002_g N_B1_N_M1005_g N_B1_N_M1003_g
+ B1_N B1_N N_B1_N_c_379_n N_B1_N_c_380_n PM_SKY130_FD_SC_LP__A21BO_LP%B1_N
x_PM_SKY130_FD_SC_LP__A21BO_LP%X N_X_M1007_s N_X_M1004_s N_X_c_420_n N_X_c_421_n
+ N_X_c_418_n X PM_SKY130_FD_SC_LP__A21BO_LP%X
x_PM_SKY130_FD_SC_LP__A21BO_LP%VPWR N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_c_445_n
+ N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n VPWR N_VPWR_c_449_n
+ N_VPWR_c_444_n N_VPWR_c_451_n PM_SKY130_FD_SC_LP__A21BO_LP%VPWR
x_PM_SKY130_FD_SC_LP__A21BO_LP%A_252_409# N_A_252_409#_M1011_d
+ N_A_252_409#_M1010_s N_A_252_409#_c_492_n N_A_252_409#_c_488_n
+ N_A_252_409#_c_489_n N_A_252_409#_c_490_n
+ PM_SKY130_FD_SC_LP__A21BO_LP%A_252_409#
x_PM_SKY130_FD_SC_LP__A21BO_LP%VGND N_VGND_M1001_d N_VGND_M1012_d N_VGND_c_519_n
+ N_VGND_c_520_n VGND N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n
+ N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n PM_SKY130_FD_SC_LP__A21BO_LP%VGND
cc_1 VNB N_A_84_29#_M1007_g 0.0247405f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.485
cc_2 VNB N_A_84_29#_c_82_n 0.0156913f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.565
cc_3 VNB N_A_84_29#_M1004_g 0.00572722f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.545
cc_4 VNB N_A_84_29#_M1001_g 0.0196379f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_5 VNB N_A_84_29#_c_85_n 0.020089f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.04
cc_6 VNB N_A_84_29#_c_86_n 0.00319029f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.363
cc_7 VNB N_A_84_29#_c_87_n 5.42725e-19 $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.96
cc_8 VNB N_A_84_29#_c_88_n 0.0297631f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=0.98
cc_9 VNB N_A_84_29#_c_89_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=0.49
cc_10 VNB N_A_84_29#_c_90_n 0.0270086f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.06
cc_11 VNB N_A_84_29#_c_91_n 0.00166494f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.565
cc_12 VNB N_A2_M1011_g 0.0032861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_176_n 0.0142328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_177_n 0.00791574f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.565
cc_15 VNB N_A2_c_178_n 0.032392f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.89
cc_16 VNB N_A2_c_179_n 0.00229272f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_17 VNB N_A2_c_180_n 0.0184075f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_18 VNB N_A1_M1009_g 0.037972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_224_n 0.00236148f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.545
cc_20 VNB N_A1_c_225_n 0.0315117f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.545
cc_21 VNB N_A1_c_226_n 0.0103911f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.363
cc_22 VNB N_A1_c_227_n 0.0134855f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.96
cc_23 VNB N_A1_c_228_n 0.00504637f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.045
cc_24 VNB N_A_308_364#_c_284_n 0.0152458f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.545
cc_25 VNB N_A_308_364#_c_285_n 0.0361216f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_26 VNB N_A_308_364#_c_286_n 0.0144368f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_27 VNB N_A_308_364#_c_287_n 0.0112149f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.89
cc_28 VNB N_A_308_364#_c_288_n 0.0181973f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.363
cc_29 VNB N_A_308_364#_c_289_n 0.00456026f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=0.49
cc_30 VNB N_A_308_364#_c_290_n 0.0422418f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=2.19
cc_31 VNB N_A_308_364#_c_291_n 0.015895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_308_364#_c_292_n 0.0380201f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=0.98
cc_33 VNB N_B1_N_M1002_g 0.0249221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B1_N_M1005_g 0.00736955f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.89
cc_35 VNB N_B1_N_M1003_g 0.0326389f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.565
cc_36 VNB N_B1_N_c_379_n 0.00803285f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.89
cc_37 VNB N_B1_N_c_380_n 0.0622642f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.04
cc_38 VNB N_X_c_418_n 0.0443486f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.89
cc_39 VNB X 0.0263965f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_40 VNB N_VPWR_c_444_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=0.895
cc_41 VNB N_VGND_c_519_n 0.00381386f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.485
cc_42 VNB N_VGND_c_520_n 0.00151893f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.545
cc_43 VNB N_VGND_c_521_n 0.0269021f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.485
cc_44 VNB N_VGND_c_522_n 0.0350157f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.39
cc_45 VNB N_VGND_c_523_n 0.0278027f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.045
cc_46 VNB N_VGND_c_524_n 0.24098f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.045
cc_47 VNB N_VGND_c_525_n 0.0048828f $X=-0.19 $Y=-0.245 $X2=1.89 $Y2=0.49
cc_48 VNB N_VGND_c_526_n 0.00485212f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=2.19
cc_49 VPB N_A_84_29#_M1004_g 0.0445401f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.545
cc_50 VPB N_A_84_29#_c_87_n 0.00247453f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=1.96
cc_51 VPB N_A_84_29#_c_94_n 0.0150521f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.045
cc_52 VPB N_A_84_29#_c_95_n 0.00531502f $X=-0.19 $Y=1.655 $X2=1.93 $Y2=2.19
cc_53 VPB N_A2_M1011_g 0.0423032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A2_c_179_n 0.00380602f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.485
cc_55 VPB N_A1_M1010_g 0.0297685f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.89
cc_56 VPB N_A1_c_224_n 0.00278567f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.545
cc_57 VPB N_A1_c_226_n 0.00229381f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.363
cc_58 VPB N_A1_c_227_n 0.0230212f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=1.96
cc_59 VPB N_A1_c_228_n 0.00521269f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.045
cc_60 VPB N_A_308_364#_c_293_n 0.0234163f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.89
cc_61 VPB N_A_308_364#_c_294_n 0.0362208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_308_364#_c_295_n 0.013466f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.565
cc_63 VPB N_A_308_364#_c_285_n 0.0114124f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.485
cc_64 VPB N_A_308_364#_c_297_n 0.0432703f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.98
cc_65 VPB N_A_308_364#_c_292_n 0.0201097f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=0.98
cc_66 VPB N_B1_N_M1005_g 0.0489126f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.89
cc_67 VPB N_B1_N_c_379_n 0.00264904f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.89
cc_68 VPB N_X_c_420_n 0.0377814f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.565
cc_69 VPB N_X_c_421_n 0.015625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_X_c_418_n 0.0179656f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.89
cc_71 VPB N_VPWR_c_445_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.565
cc_72 VPB N_VPWR_c_446_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.89
cc_73 VPB N_VPWR_c_447_n 0.0433031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_448_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.04
cc_75 VPB N_VPWR_c_449_n 0.0189139f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.045
cc_76 VPB N_VPWR_c_444_n 0.0547389f $X=-0.19 $Y=1.655 $X2=1.89 $Y2=0.895
cc_77 VPB N_VPWR_c_451_n 0.024803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_252_409#_c_488_n 0.0138356f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.565
cc_79 VPB N_A_252_409#_c_489_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.545
cc_80 VPB N_A_252_409#_c_490_n 0.00825655f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.89
cc_81 N_A_84_29#_c_94_n N_A2_M1011_g 0.0217848f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_82 N_A_84_29#_c_95_n N_A2_M1011_g 8.26284e-19 $X=1.93 $Y=2.19 $X2=0 $Y2=0
cc_83 N_A_84_29#_c_91_n N_A2_M1011_g 0.0034979f $X=0.642 $Y=1.565 $X2=0 $Y2=0
cc_84 N_A_84_29#_M1001_g N_A2_c_176_n 0.0108719f $X=0.855 $Y=0.485 $X2=0 $Y2=0
cc_85 N_A_84_29#_c_89_n N_A2_c_176_n 0.00216292f $X=1.89 $Y=0.49 $X2=0 $Y2=0
cc_86 N_A_84_29#_M1001_g N_A2_c_177_n 0.0065895f $X=0.855 $Y=0.485 $X2=0 $Y2=0
cc_87 N_A_84_29#_c_88_n N_A2_c_177_n 0.00691064f $X=1.725 $Y=0.98 $X2=0 $Y2=0
cc_88 N_A_84_29#_M1004_g N_A2_c_178_n 0.0376583f $X=0.595 $Y=2.545 $X2=0 $Y2=0
cc_89 N_A_84_29#_c_86_n N_A2_c_178_n 0.0034979f $X=0.642 $Y=1.363 $X2=0 $Y2=0
cc_90 N_A_84_29#_c_88_n N_A2_c_178_n 0.0018185f $X=1.725 $Y=0.98 $X2=0 $Y2=0
cc_91 N_A_84_29#_c_94_n N_A2_c_178_n 4.33375e-19 $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_92 N_A_84_29#_c_90_n N_A2_c_178_n 0.015028f $X=0.605 $Y=1.06 $X2=0 $Y2=0
cc_93 N_A_84_29#_M1004_g N_A2_c_179_n 2.17164e-19 $X=0.595 $Y=2.545 $X2=0 $Y2=0
cc_94 N_A_84_29#_c_86_n N_A2_c_179_n 0.0373286f $X=0.642 $Y=1.363 $X2=0 $Y2=0
cc_95 N_A_84_29#_c_88_n N_A2_c_179_n 0.02085f $X=1.725 $Y=0.98 $X2=0 $Y2=0
cc_96 N_A_84_29#_c_94_n N_A2_c_179_n 0.0240247f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_97 N_A_84_29#_c_90_n N_A2_c_179_n 3.07878e-19 $X=0.605 $Y=1.06 $X2=0 $Y2=0
cc_98 N_A_84_29#_c_85_n N_A2_c_180_n 0.0065895f $X=0.675 $Y=1.04 $X2=0 $Y2=0
cc_99 N_A_84_29#_c_86_n N_A2_c_180_n 0.00444278f $X=0.642 $Y=1.363 $X2=0 $Y2=0
cc_100 N_A_84_29#_c_88_n N_A2_c_180_n 0.00756033f $X=1.725 $Y=0.98 $X2=0 $Y2=0
cc_101 N_A_84_29#_c_90_n N_A2_c_180_n 0.00550782f $X=0.605 $Y=1.06 $X2=0 $Y2=0
cc_102 N_A_84_29#_c_88_n N_A1_M1009_g 0.0138276f $X=1.725 $Y=0.98 $X2=0 $Y2=0
cc_103 N_A_84_29#_c_89_n N_A1_M1009_g 0.0136339f $X=1.89 $Y=0.49 $X2=0 $Y2=0
cc_104 N_A_84_29#_c_94_n N_A1_M1010_g 0.00406235f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_105 N_A_84_29#_c_95_n N_A1_M1010_g 0.00151067f $X=1.93 $Y=2.19 $X2=0 $Y2=0
cc_106 N_A_84_29#_c_88_n N_A1_c_224_n 0.024979f $X=1.725 $Y=0.98 $X2=0 $Y2=0
cc_107 N_A_84_29#_c_94_n N_A1_c_224_n 0.0207657f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_108 N_A_84_29#_c_88_n N_A1_c_225_n 0.00136218f $X=1.725 $Y=0.98 $X2=0 $Y2=0
cc_109 N_A_84_29#_c_94_n N_A1_c_225_n 2.69898e-19 $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_110 N_A_84_29#_c_88_n N_A1_c_228_n 0.00530346f $X=1.725 $Y=0.98 $X2=0 $Y2=0
cc_111 N_A_84_29#_c_94_n N_A1_c_228_n 0.0104686f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_112 N_A_84_29#_c_94_n N_A_308_364#_c_293_n 0.0162153f $X=1.765 $Y=2.045 $X2=0
+ $Y2=0
cc_113 N_A_84_29#_c_95_n N_A_308_364#_c_293_n 0.0107492f $X=1.93 $Y=2.19 $X2=0
+ $Y2=0
cc_114 N_A_84_29#_c_94_n N_A_308_364#_c_294_n 0.0109161f $X=1.765 $Y=2.045 $X2=0
+ $Y2=0
cc_115 N_A_84_29#_c_94_n N_A_308_364#_c_295_n 0.00435706f $X=1.765 $Y=2.045
+ $X2=0 $Y2=0
cc_116 N_A_84_29#_c_89_n N_A_308_364#_c_284_n 0.0101247f $X=1.89 $Y=0.49 $X2=0
+ $Y2=0
cc_117 N_A_84_29#_c_89_n N_A_308_364#_c_286_n 0.00165313f $X=1.89 $Y=0.49 $X2=0
+ $Y2=0
cc_118 N_A_84_29#_c_88_n N_A_308_364#_c_289_n 0.0126551f $X=1.725 $Y=0.98 $X2=0
+ $Y2=0
cc_119 N_A_84_29#_c_89_n N_A_308_364#_c_289_n 0.0145356f $X=1.89 $Y=0.49 $X2=0
+ $Y2=0
cc_120 N_A_84_29#_c_88_n N_A_308_364#_c_290_n 0.00340271f $X=1.725 $Y=0.98 $X2=0
+ $Y2=0
cc_121 N_A_84_29#_c_89_n N_A_308_364#_c_290_n 0.00260777f $X=1.89 $Y=0.49 $X2=0
+ $Y2=0
cc_122 N_A_84_29#_M1004_g N_X_c_420_n 0.0150657f $X=0.595 $Y=2.545 $X2=0 $Y2=0
cc_123 N_A_84_29#_c_82_n N_X_c_421_n 9.45561e-19 $X=0.595 $Y=1.565 $X2=0 $Y2=0
cc_124 N_A_84_29#_M1004_g N_X_c_421_n 0.00470913f $X=0.595 $Y=2.545 $X2=0 $Y2=0
cc_125 N_A_84_29#_c_140_p N_X_c_421_n 0.00812422f $X=0.845 $Y=2.045 $X2=0 $Y2=0
cc_126 N_A_84_29#_c_91_n N_X_c_421_n 0.00212147f $X=0.642 $Y=1.565 $X2=0 $Y2=0
cc_127 N_A_84_29#_M1007_g N_X_c_418_n 0.0202005f $X=0.495 $Y=0.485 $X2=0 $Y2=0
cc_128 N_A_84_29#_M1004_g N_X_c_418_n 0.00928062f $X=0.595 $Y=2.545 $X2=0 $Y2=0
cc_129 N_A_84_29#_c_144_p N_X_c_418_n 0.012967f $X=0.642 $Y=1.065 $X2=0 $Y2=0
cc_130 N_A_84_29#_c_86_n N_X_c_418_n 0.0364526f $X=0.642 $Y=1.363 $X2=0 $Y2=0
cc_131 N_A_84_29#_c_87_n N_X_c_418_n 0.0144799f $X=0.76 $Y=1.96 $X2=0 $Y2=0
cc_132 N_A_84_29#_c_140_p N_X_c_418_n 6.10912e-19 $X=0.845 $Y=2.045 $X2=0 $Y2=0
cc_133 N_A_84_29#_M1007_g X 0.00978536f $X=0.495 $Y=0.485 $X2=0 $Y2=0
cc_134 N_A_84_29#_M1001_g X 0.00122413f $X=0.855 $Y=0.485 $X2=0 $Y2=0
cc_135 N_A_84_29#_c_94_n N_VPWR_M1004_d 0.00116505f $X=1.765 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_84_29#_c_140_p N_VPWR_M1004_d 7.70949e-19 $X=0.845 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_84_29#_M1004_g N_VPWR_c_445_n 0.0189731f $X=0.595 $Y=2.545 $X2=0
+ $Y2=0
cc_138 N_A_84_29#_c_94_n N_VPWR_c_445_n 0.0093622f $X=1.765 $Y=2.045 $X2=0 $Y2=0
cc_139 N_A_84_29#_c_140_p N_VPWR_c_445_n 0.00777198f $X=0.845 $Y=2.045 $X2=0
+ $Y2=0
cc_140 N_A_84_29#_M1004_g N_VPWR_c_444_n 0.0141137f $X=0.595 $Y=2.545 $X2=0
+ $Y2=0
cc_141 N_A_84_29#_M1004_g N_VPWR_c_451_n 0.00769046f $X=0.595 $Y=2.545 $X2=0
+ $Y2=0
cc_142 N_A_84_29#_c_94_n N_A_252_409#_M1011_d 0.00180746f $X=1.765 $Y=2.045
+ $X2=-0.19 $Y2=-0.245
cc_143 N_A_84_29#_c_94_n N_A_252_409#_c_492_n 0.0163515f $X=1.765 $Y=2.045 $X2=0
+ $Y2=0
cc_144 N_A_84_29#_c_95_n N_A_252_409#_c_492_n 0.0266857f $X=1.93 $Y=2.19 $X2=0
+ $Y2=0
cc_145 N_A_84_29#_M1006_d N_A_252_409#_c_488_n 0.00334849f $X=1.79 $Y=2.045
+ $X2=0 $Y2=0
cc_146 N_A_84_29#_c_95_n N_A_252_409#_c_488_n 0.0195854f $X=1.93 $Y=2.19 $X2=0
+ $Y2=0
cc_147 N_A_84_29#_c_94_n N_A_252_409#_c_490_n 0.00107309f $X=1.765 $Y=2.045
+ $X2=0 $Y2=0
cc_148 N_A_84_29#_c_95_n N_A_252_409#_c_490_n 0.0394061f $X=1.93 $Y=2.19 $X2=0
+ $Y2=0
cc_149 N_A_84_29#_M1007_g N_VGND_c_519_n 0.00216919f $X=0.495 $Y=0.485 $X2=0
+ $Y2=0
cc_150 N_A_84_29#_M1001_g N_VGND_c_519_n 0.0125847f $X=0.855 $Y=0.485 $X2=0
+ $Y2=0
cc_151 N_A_84_29#_c_88_n N_VGND_c_519_n 0.0261819f $X=1.725 $Y=0.98 $X2=0 $Y2=0
cc_152 N_A_84_29#_c_89_n N_VGND_c_519_n 0.0142563f $X=1.89 $Y=0.49 $X2=0 $Y2=0
cc_153 N_A_84_29#_c_89_n N_VGND_c_520_n 0.00802976f $X=1.89 $Y=0.49 $X2=0 $Y2=0
cc_154 N_A_84_29#_M1007_g N_VGND_c_521_n 0.00511657f $X=0.495 $Y=0.485 $X2=0
+ $Y2=0
cc_155 N_A_84_29#_M1001_g N_VGND_c_521_n 0.00452967f $X=0.855 $Y=0.485 $X2=0
+ $Y2=0
cc_156 N_A_84_29#_c_89_n N_VGND_c_522_n 0.021949f $X=1.89 $Y=0.49 $X2=0 $Y2=0
cc_157 N_A_84_29#_M1007_g N_VGND_c_524_n 0.010231f $X=0.495 $Y=0.485 $X2=0 $Y2=0
cc_158 N_A_84_29#_M1001_g N_VGND_c_524_n 0.00799963f $X=0.855 $Y=0.485 $X2=0
+ $Y2=0
cc_159 N_A_84_29#_c_89_n N_VGND_c_524_n 0.0124703f $X=1.89 $Y=0.49 $X2=0 $Y2=0
cc_160 N_A2_c_176_n N_A1_M1009_g 0.0398149f $X=1.282 $Y=0.77 $X2=0 $Y2=0
cc_161 N_A2_c_180_n N_A1_M1009_g 0.0182666f $X=1.182 $Y=1.28 $X2=0 $Y2=0
cc_162 N_A2_M1011_g N_A1_c_224_n 6.25964e-19 $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_163 N_A2_c_178_n N_A1_c_224_n 6.60303e-19 $X=1.19 $Y=1.445 $X2=0 $Y2=0
cc_164 N_A2_c_179_n N_A1_c_224_n 0.0261275f $X=1.19 $Y=1.445 $X2=0 $Y2=0
cc_165 N_A2_c_180_n N_A1_c_224_n 0.00130558f $X=1.182 $Y=1.28 $X2=0 $Y2=0
cc_166 N_A2_c_179_n N_A1_c_225_n 0.00110444f $X=1.19 $Y=1.445 $X2=0 $Y2=0
cc_167 N_A2_c_180_n N_A1_c_225_n 0.0172357f $X=1.182 $Y=1.28 $X2=0 $Y2=0
cc_168 N_A2_M1011_g N_A_308_364#_c_295_n 0.031184f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_169 N_A2_M1011_g N_X_c_420_n 2.06137e-19 $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_170 N_A2_M1011_g N_X_c_421_n 7.68609e-19 $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_171 N_A2_M1011_g N_VPWR_c_445_n 0.0170675f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_172 N_A2_M1011_g N_VPWR_c_447_n 0.00803391f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_173 N_A2_M1011_g N_VPWR_c_444_n 0.0140321f $X=1.135 $Y=2.545 $X2=0 $Y2=0
cc_174 N_A2_M1011_g N_A_252_409#_c_492_n 0.0107683f $X=1.135 $Y=2.545 $X2=0
+ $Y2=0
cc_175 N_A2_M1011_g N_A_252_409#_c_489_n 0.0034262f $X=1.135 $Y=2.545 $X2=0
+ $Y2=0
cc_176 N_A2_c_176_n N_VGND_c_519_n 0.0128898f $X=1.282 $Y=0.77 $X2=0 $Y2=0
cc_177 N_A2_c_176_n N_VGND_c_522_n 0.00452967f $X=1.282 $Y=0.77 $X2=0 $Y2=0
cc_178 N_A2_c_176_n N_VGND_c_524_n 0.00809218f $X=1.282 $Y=0.77 $X2=0 $Y2=0
cc_179 N_A1_M1010_g N_A_308_364#_c_294_n 0.00165492f $X=2.755 $Y=2.595 $X2=0
+ $Y2=0
cc_180 N_A1_c_228_n N_A_308_364#_c_294_n 0.00514458f $X=2.495 $Y=1.742 $X2=0
+ $Y2=0
cc_181 N_A1_c_224_n N_A_308_364#_c_295_n 0.00280433f $X=1.76 $Y=1.415 $X2=0
+ $Y2=0
cc_182 N_A1_c_225_n N_A_308_364#_c_295_n 0.0174782f $X=1.76 $Y=1.415 $X2=0 $Y2=0
cc_183 N_A1_M1009_g N_A_308_364#_c_284_n 0.0195831f $X=1.675 $Y=0.485 $X2=0
+ $Y2=0
cc_184 N_A1_c_224_n N_A_308_364#_c_285_n 0.00263535f $X=1.76 $Y=1.415 $X2=0
+ $Y2=0
cc_185 N_A1_c_225_n N_A_308_364#_c_285_n 0.0211979f $X=1.76 $Y=1.415 $X2=0 $Y2=0
cc_186 N_A1_c_226_n N_A_308_364#_c_285_n 0.00154476f $X=2.66 $Y=1.77 $X2=0 $Y2=0
cc_187 N_A1_c_227_n N_A_308_364#_c_285_n 0.021056f $X=2.755 $Y=1.77 $X2=0 $Y2=0
cc_188 N_A1_c_228_n N_A_308_364#_c_285_n 0.0192893f $X=2.495 $Y=1.742 $X2=0
+ $Y2=0
cc_189 N_A1_M1010_g N_A_308_364#_c_297_n 4.70481e-19 $X=2.755 $Y=2.595 $X2=0
+ $Y2=0
cc_190 N_A1_M1009_g N_A_308_364#_c_289_n 5.03381e-19 $X=1.675 $Y=0.485 $X2=0
+ $Y2=0
cc_191 N_A1_c_228_n N_A_308_364#_c_289_n 0.0130443f $X=2.495 $Y=1.742 $X2=0
+ $Y2=0
cc_192 N_A1_M1009_g N_A_308_364#_c_290_n 0.00990693f $X=1.675 $Y=0.485 $X2=0
+ $Y2=0
cc_193 N_A1_c_227_n N_A_308_364#_c_290_n 0.00184401f $X=2.755 $Y=1.77 $X2=0
+ $Y2=0
cc_194 N_A1_c_228_n N_A_308_364#_c_290_n 0.00381916f $X=2.495 $Y=1.742 $X2=0
+ $Y2=0
cc_195 N_A1_c_226_n N_B1_N_M1005_g 0.00136429f $X=2.66 $Y=1.77 $X2=0 $Y2=0
cc_196 N_A1_c_227_n N_B1_N_M1005_g 0.0417501f $X=2.755 $Y=1.77 $X2=0 $Y2=0
cc_197 N_A1_c_226_n N_B1_N_c_379_n 0.0183965f $X=2.66 $Y=1.77 $X2=0 $Y2=0
cc_198 N_A1_c_227_n N_B1_N_c_379_n 0.00130551f $X=2.755 $Y=1.77 $X2=0 $Y2=0
cc_199 N_A1_c_227_n N_B1_N_c_380_n 0.00258884f $X=2.755 $Y=1.77 $X2=0 $Y2=0
cc_200 N_A1_M1010_g N_VPWR_c_446_n 0.0271319f $X=2.755 $Y=2.595 $X2=0 $Y2=0
cc_201 N_A1_M1010_g N_VPWR_c_447_n 0.00838695f $X=2.755 $Y=2.595 $X2=0 $Y2=0
cc_202 N_A1_M1010_g N_VPWR_c_444_n 0.01486f $X=2.755 $Y=2.595 $X2=0 $Y2=0
cc_203 N_A1_M1010_g N_A_252_409#_c_488_n 0.00315189f $X=2.755 $Y=2.595 $X2=0
+ $Y2=0
cc_204 N_A1_M1010_g N_A_252_409#_c_490_n 0.0180531f $X=2.755 $Y=2.595 $X2=0
+ $Y2=0
cc_205 N_A1_c_226_n N_A_252_409#_c_490_n 0.0101402f $X=2.66 $Y=1.77 $X2=0 $Y2=0
cc_206 N_A1_c_227_n N_A_252_409#_c_490_n 0.00294988f $X=2.755 $Y=1.77 $X2=0
+ $Y2=0
cc_207 N_A1_c_228_n N_A_252_409#_c_490_n 0.00764414f $X=2.495 $Y=1.742 $X2=0
+ $Y2=0
cc_208 N_A1_M1009_g N_VGND_c_519_n 0.00218527f $X=1.675 $Y=0.485 $X2=0 $Y2=0
cc_209 N_A1_M1009_g N_VGND_c_522_n 0.00511657f $X=1.675 $Y=0.485 $X2=0 $Y2=0
cc_210 N_A1_M1009_g N_VGND_c_524_n 0.00961146f $X=1.675 $Y=0.485 $X2=0 $Y2=0
cc_211 N_A_308_364#_c_286_n N_B1_N_M1002_g 0.014791f $X=2.465 $Y=0.805 $X2=0
+ $Y2=0
cc_212 N_A_308_364#_c_287_n N_B1_N_M1002_g 0.0149001f $X=3.305 $Y=0.77 $X2=0
+ $Y2=0
cc_213 N_A_308_364#_c_288_n N_B1_N_M1002_g 0.00155292f $X=3.47 $Y=0.49 $X2=0
+ $Y2=0
cc_214 N_A_308_364#_c_289_n N_B1_N_M1002_g 0.00173551f $X=2.415 $Y=0.77 $X2=0
+ $Y2=0
cc_215 N_A_308_364#_c_290_n N_B1_N_M1002_g 0.0188655f $X=2.415 $Y=0.97 $X2=0
+ $Y2=0
cc_216 N_A_308_364#_c_297_n N_B1_N_M1005_g 0.0239682f $X=3.55 $Y=2.24 $X2=0
+ $Y2=0
cc_217 N_A_308_364#_c_287_n N_B1_N_M1003_g 0.00818279f $X=3.305 $Y=0.77 $X2=0
+ $Y2=0
cc_218 N_A_308_364#_c_288_n N_B1_N_M1003_g 0.00771803f $X=3.47 $Y=0.49 $X2=0
+ $Y2=0
cc_219 N_A_308_364#_c_291_n N_B1_N_M1003_g 0.00437795f $X=3.51 $Y=0.77 $X2=0
+ $Y2=0
cc_220 N_A_308_364#_c_292_n N_B1_N_M1003_g 0.00422422f $X=3.55 $Y=2.075 $X2=0
+ $Y2=0
cc_221 N_A_308_364#_c_287_n N_B1_N_c_379_n 0.0223763f $X=3.305 $Y=0.77 $X2=0
+ $Y2=0
cc_222 N_A_308_364#_c_289_n N_B1_N_c_379_n 0.00357866f $X=2.415 $Y=0.77 $X2=0
+ $Y2=0
cc_223 N_A_308_364#_c_290_n N_B1_N_c_379_n 2.93574e-19 $X=2.415 $Y=0.97 $X2=0
+ $Y2=0
cc_224 N_A_308_364#_c_291_n N_B1_N_c_379_n 0.00233735f $X=3.51 $Y=0.77 $X2=0
+ $Y2=0
cc_225 N_A_308_364#_c_292_n N_B1_N_c_379_n 0.0477474f $X=3.55 $Y=2.075 $X2=0
+ $Y2=0
cc_226 N_A_308_364#_c_285_n N_B1_N_c_380_n 0.00557293f $X=2.21 $Y=1.82 $X2=0
+ $Y2=0
cc_227 N_A_308_364#_c_287_n N_B1_N_c_380_n 2.08868e-19 $X=3.305 $Y=0.77 $X2=0
+ $Y2=0
cc_228 N_A_308_364#_c_291_n N_B1_N_c_380_n 0.00233943f $X=3.51 $Y=0.77 $X2=0
+ $Y2=0
cc_229 N_A_308_364#_c_292_n N_B1_N_c_380_n 0.0259081f $X=3.55 $Y=2.075 $X2=0
+ $Y2=0
cc_230 N_A_308_364#_c_293_n N_VPWR_c_445_n 8.69147e-19 $X=1.665 $Y=1.97 $X2=0
+ $Y2=0
cc_231 N_A_308_364#_c_297_n N_VPWR_c_446_n 0.0625632f $X=3.55 $Y=2.24 $X2=0
+ $Y2=0
cc_232 N_A_308_364#_c_293_n N_VPWR_c_447_n 0.00546179f $X=1.665 $Y=1.97 $X2=0
+ $Y2=0
cc_233 N_A_308_364#_c_297_n N_VPWR_c_449_n 0.019758f $X=3.55 $Y=2.24 $X2=0 $Y2=0
cc_234 N_A_308_364#_M1005_d N_VPWR_c_444_n 0.0023218f $X=3.41 $Y=2.095 $X2=0
+ $Y2=0
cc_235 N_A_308_364#_c_293_n N_VPWR_c_444_n 0.00832053f $X=1.665 $Y=1.97 $X2=0
+ $Y2=0
cc_236 N_A_308_364#_c_297_n N_VPWR_c_444_n 0.012508f $X=3.55 $Y=2.24 $X2=0 $Y2=0
cc_237 N_A_308_364#_c_293_n N_A_252_409#_c_492_n 0.0158233f $X=1.665 $Y=1.97
+ $X2=0 $Y2=0
cc_238 N_A_308_364#_c_293_n N_A_252_409#_c_488_n 0.0185974f $X=1.665 $Y=1.97
+ $X2=0 $Y2=0
cc_239 N_A_308_364#_c_293_n N_A_252_409#_c_489_n 8.05528e-19 $X=1.665 $Y=1.97
+ $X2=0 $Y2=0
cc_240 N_A_308_364#_c_293_n N_A_252_409#_c_490_n 0.0044139f $X=1.665 $Y=1.97
+ $X2=0 $Y2=0
cc_241 N_A_308_364#_c_287_n N_VGND_M1012_d 0.00175078f $X=3.305 $Y=0.77 $X2=0
+ $Y2=0
cc_242 N_A_308_364#_c_284_n N_VGND_c_520_n 0.00159761f $X=2.105 $Y=0.805 $X2=0
+ $Y2=0
cc_243 N_A_308_364#_c_286_n N_VGND_c_520_n 0.00862393f $X=2.465 $Y=0.805 $X2=0
+ $Y2=0
cc_244 N_A_308_364#_c_287_n N_VGND_c_520_n 0.0138269f $X=3.305 $Y=0.77 $X2=0
+ $Y2=0
cc_245 N_A_308_364#_c_288_n N_VGND_c_520_n 0.00802976f $X=3.47 $Y=0.49 $X2=0
+ $Y2=0
cc_246 N_A_308_364#_c_289_n N_VGND_c_520_n 0.00173106f $X=2.415 $Y=0.77 $X2=0
+ $Y2=0
cc_247 N_A_308_364#_c_284_n N_VGND_c_522_n 0.00511657f $X=2.105 $Y=0.805 $X2=0
+ $Y2=0
cc_248 N_A_308_364#_c_286_n N_VGND_c_522_n 0.00332032f $X=2.465 $Y=0.805 $X2=0
+ $Y2=0
cc_249 N_A_308_364#_c_289_n N_VGND_c_522_n 0.00381057f $X=2.415 $Y=0.77 $X2=0
+ $Y2=0
cc_250 N_A_308_364#_c_287_n N_VGND_c_523_n 0.00611534f $X=3.305 $Y=0.77 $X2=0
+ $Y2=0
cc_251 N_A_308_364#_c_288_n N_VGND_c_523_n 0.0218625f $X=3.47 $Y=0.49 $X2=0
+ $Y2=0
cc_252 N_A_308_364#_c_291_n N_VGND_c_523_n 0.00146557f $X=3.51 $Y=0.77 $X2=0
+ $Y2=0
cc_253 N_A_308_364#_c_284_n N_VGND_c_524_n 0.00951891f $X=2.105 $Y=0.805 $X2=0
+ $Y2=0
cc_254 N_A_308_364#_c_286_n N_VGND_c_524_n 0.00393697f $X=2.465 $Y=0.805 $X2=0
+ $Y2=0
cc_255 N_A_308_364#_c_287_n N_VGND_c_524_n 0.0125194f $X=3.305 $Y=0.77 $X2=0
+ $Y2=0
cc_256 N_A_308_364#_c_288_n N_VGND_c_524_n 0.0125454f $X=3.47 $Y=0.49 $X2=0
+ $Y2=0
cc_257 N_A_308_364#_c_289_n N_VGND_c_524_n 0.00724832f $X=2.415 $Y=0.77 $X2=0
+ $Y2=0
cc_258 N_A_308_364#_c_291_n N_VGND_c_524_n 0.00233963f $X=3.51 $Y=0.77 $X2=0
+ $Y2=0
cc_259 N_A_308_364#_c_289_n A_436_55# 0.00164821f $X=2.415 $Y=0.77 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_308_364#_c_287_n A_594_55# 0.00176688f $X=3.305 $Y=0.77 $X2=-0.19
+ $Y2=-0.245
cc_261 N_B1_N_M1005_g N_VPWR_c_446_n 0.0264975f $X=3.285 $Y=2.595 $X2=0 $Y2=0
cc_262 N_B1_N_c_379_n N_VPWR_c_446_n 0.00828734f $X=3.17 $Y=1.2 $X2=0 $Y2=0
cc_263 N_B1_N_M1005_g N_VPWR_c_449_n 0.00840199f $X=3.285 $Y=2.595 $X2=0 $Y2=0
cc_264 N_B1_N_M1005_g N_VPWR_c_444_n 0.0145332f $X=3.285 $Y=2.595 $X2=0 $Y2=0
cc_265 N_B1_N_M1005_g N_A_252_409#_c_490_n 2.95915e-19 $X=3.285 $Y=2.595 $X2=0
+ $Y2=0
cc_266 N_B1_N_M1002_g N_VGND_c_520_n 0.00862492f $X=2.895 $Y=0.485 $X2=0 $Y2=0
cc_267 N_B1_N_M1003_g N_VGND_c_520_n 0.00159761f $X=3.255 $Y=0.485 $X2=0 $Y2=0
cc_268 N_B1_N_M1002_g N_VGND_c_523_n 0.00332138f $X=2.895 $Y=0.485 $X2=0 $Y2=0
cc_269 N_B1_N_M1003_g N_VGND_c_523_n 0.00389854f $X=3.255 $Y=0.485 $X2=0 $Y2=0
cc_270 N_B1_N_M1002_g N_VGND_c_524_n 0.00393904f $X=2.895 $Y=0.485 $X2=0 $Y2=0
cc_271 N_B1_N_M1003_g N_VGND_c_524_n 0.00621052f $X=3.255 $Y=0.485 $X2=0 $Y2=0
cc_272 N_X_c_420_n N_VPWR_c_445_n 0.0505393f $X=0.33 $Y=2.9 $X2=0 $Y2=0
cc_273 N_X_c_420_n N_VPWR_c_444_n 0.0154828f $X=0.33 $Y=2.9 $X2=0 $Y2=0
cc_274 N_X_c_420_n N_VPWR_c_451_n 0.0270889f $X=0.33 $Y=2.9 $X2=0 $Y2=0
cc_275 X N_VGND_c_519_n 0.0151404f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_276 X N_VGND_c_521_n 0.0233465f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_277 X N_VGND_c_524_n 0.0134709f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_278 N_VPWR_c_444_n N_A_252_409#_M1010_s 0.0023218f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_279 N_VPWR_c_445_n N_A_252_409#_c_492_n 0.0370422f $X=0.86 $Y=2.475 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_446_n N_A_252_409#_c_488_n 0.0119061f $X=3.02 $Y=2.28 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_447_n N_A_252_409#_c_488_n 0.0652481f $X=2.855 $Y=3.33 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_444_n N_A_252_409#_c_488_n 0.0399424f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_283 N_VPWR_c_445_n N_A_252_409#_c_489_n 0.0114492f $X=0.86 $Y=2.475 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_447_n N_A_252_409#_c_489_n 0.0220769f $X=2.855 $Y=3.33 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_444_n N_A_252_409#_c_489_n 0.0125384f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_286 N_VPWR_c_446_n N_A_252_409#_c_490_n 0.0513618f $X=3.02 $Y=2.28 $X2=0
+ $Y2=0
