# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__bufinv_16
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__bufinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.945000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.415000 1.570000 1.760000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  4.704000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.640000 1.920000 10.950000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.520000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.520000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.245000 11.520000 3.415000 ;
      RECT  0.275000  0.315000  0.570000 1.075000 ;
      RECT  0.275000  1.075000  1.920000 1.245000 ;
      RECT  0.275000  1.930000  1.920000 2.100000 ;
      RECT  0.275000  2.100000  0.570000 3.025000 ;
      RECT  0.740000  0.085000  1.000000 0.905000 ;
      RECT  0.740000  2.270000  1.000000 3.245000 ;
      RECT  1.170000  0.315000  1.430000 1.075000 ;
      RECT  1.170000  2.100000  1.430000 3.025000 ;
      RECT  1.600000  0.085000  1.870000 0.905000 ;
      RECT  1.600000  2.270000  1.905000 3.245000 ;
      RECT  1.750000  1.245000  1.920000 1.395000 ;
      RECT  1.750000  1.395000  4.170000 1.585000 ;
      RECT  1.750000  1.585000  1.920000 1.930000 ;
      RECT  2.090000  0.315000  2.335000 1.055000 ;
      RECT  2.090000  1.055000  4.520000 1.225000 ;
      RECT  2.090000  1.755000  4.520000 1.925000 ;
      RECT  2.090000  1.925000  2.335000 3.025000 ;
      RECT  2.505000  0.085000  2.765000 0.885000 ;
      RECT  2.505000  2.105000  2.765000 3.245000 ;
      RECT  2.935000  0.315000  3.195000 1.055000 ;
      RECT  2.935000  1.925000  3.195000 3.025000 ;
      RECT  3.365000  0.085000  3.625000 0.885000 ;
      RECT  3.365000  2.105000  3.625000 3.245000 ;
      RECT  3.795000  0.315000  4.055000 1.055000 ;
      RECT  3.795000  1.925000  4.055000 3.025000 ;
      RECT  4.225000  0.085000  4.485000 0.885000 ;
      RECT  4.225000  2.105000  4.485000 3.245000 ;
      RECT  4.340000  1.225000  4.520000 1.755000 ;
      RECT  4.690000  0.315000  4.915000 3.025000 ;
      RECT  5.085000  0.085000  5.345000 1.080000 ;
      RECT  5.085000  1.345000  5.345000 1.785000 ;
      RECT  5.085000  1.955000  5.345000 3.245000 ;
      RECT  5.515000  0.315000  5.775000 3.025000 ;
      RECT  5.945000  0.085000  6.205000 1.080000 ;
      RECT  5.945000  1.345000  6.205000 1.785000 ;
      RECT  5.945000  1.955000  6.205000 3.245000 ;
      RECT  6.375000  0.315000  6.635000 3.025000 ;
      RECT  6.805000  0.085000  7.065000 1.080000 ;
      RECT  6.805000  1.345000  7.065000 1.785000 ;
      RECT  6.805000  1.955000  7.065000 3.245000 ;
      RECT  7.235000  0.315000  7.495000 3.025000 ;
      RECT  7.665000  0.085000  7.925000 1.080000 ;
      RECT  7.665000  1.345000  7.925000 1.785000 ;
      RECT  7.665000  1.955000  7.925000 3.245000 ;
      RECT  8.095000  0.315000  8.355000 3.025000 ;
      RECT  8.525000  0.085000  8.785000 1.080000 ;
      RECT  8.525000  1.345000  8.785000 1.785000 ;
      RECT  8.525000  1.955000  8.785000 3.245000 ;
      RECT  8.955000  0.315000  9.215000 3.025000 ;
      RECT  9.385000  0.085000  9.645000 1.080000 ;
      RECT  9.385000  1.345000  9.645000 1.785000 ;
      RECT  9.385000  1.955000  9.645000 3.245000 ;
      RECT  9.815000  0.315000 10.075000 3.025000 ;
      RECT 10.245000  0.085000 10.505000 1.080000 ;
      RECT 10.245000  1.345000 10.505000 1.785000 ;
      RECT 10.245000  1.955000 10.505000 3.245000 ;
      RECT 10.675000  0.315000 10.935000 3.025000 ;
      RECT 11.105000  0.085000 11.400000 1.080000 ;
      RECT 11.105000  1.955000 11.400000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.350000  1.580000  4.520000 1.750000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.700000  1.950000  4.870000 2.120000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.130000  1.580000  5.300000 1.750000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.560000  1.950000  5.730000 2.120000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  5.990000  1.580000  6.160000 1.750000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.420000  1.950000  6.590000 2.120000 ;
      RECT  6.850000  1.580000  7.020000 1.750000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.280000  1.950000  7.450000 2.120000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.710000  1.580000  7.880000 1.750000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.140000  1.950000  8.310000 2.120000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.570000  1.580000  8.740000 1.750000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.000000  1.950000  9.170000 2.120000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.430000  1.580000  9.600000 1.750000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT  9.860000  1.950000 10.030000 2.120000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.290000  1.580000 10.460000 1.750000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 10.720000  1.950000 10.890000 2.120000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
    LAYER met1 ;
      RECT 4.290000 1.550000 10.520000 1.780000 ;
  END
END sky130_fd_sc_lp__bufinv_16
END LIBRARY
