* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311a_lp A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR B1 a_84_115# VPB phighvt w=1e+06u l=250000u
+  ad=6.45e+11p pd=5.29e+06u as=5.75e+11p ps=5.15e+06u
M1001 a_114_141# a_84_115# X VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1002 VGND A2 a_273_141# VNB nshort w=420000u l=150000u
+  ad=3.045e+11p pd=3.13e+06u as=2.352e+11p ps=2.8e+06u
M1003 a_356_419# A2 a_258_419# VPB phighvt w=1e+06u l=250000u
+  ad=2.9e+11p pd=2.58e+06u as=2.4e+11p ps=2.48e+06u
M1004 a_84_115# C1 a_563_141# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1005 a_84_115# C1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_273_141# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_273_141# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_563_141# B1 a_273_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_84_115# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1010 a_84_115# A3 a_356_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_84_115# a_114_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_258_419# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends
