* File: sky130_fd_sc_lp__einvn_lp.pex.spice
* Created: Fri Aug 28 10:33:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVN_LP%TE_B 3 5 7 10 12 14 15 21 22
c43 21 0 7.36295e-20 $X=0.77 $Y=1.745
r44 20 22 14.1765 $w=3.06e-07 $l=9e-08 $layer=POLY_cond $X=0.77 $Y=1.787
+ $X2=0.86 $Y2=1.787
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.745 $X2=0.77 $Y2=1.745
r46 18 20 25.9902 $w=3.06e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.787
+ $X2=0.77 $Y2=1.787
r47 17 18 16.5392 $w=3.06e-07 $l=1.05e-07 $layer=POLY_cond $X=0.5 $Y=1.787
+ $X2=0.605 $Y2=1.787
r48 15 21 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.77 $Y=2.035
+ $X2=0.77 $Y2=1.745
r49 12 22 43.317 $w=3.06e-07 $l=3.64452e-07 $layer=POLY_cond $X=1.135 $Y=1.995
+ $X2=0.86 $Y2=1.787
r50 12 14 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.135 $Y=1.995
+ $X2=1.135 $Y2=2.57
r51 8 22 19.4347 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.86 $Y=1.58
+ $X2=0.86 $Y2=1.787
r52 8 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.86 $Y=1.58 $X2=0.86
+ $Y2=0.95
r53 5 18 7.59805 $w=2.5e-07 $l=2.08e-07 $layer=POLY_cond $X=0.605 $Y=1.995
+ $X2=0.605 $Y2=1.787
r54 5 7 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=0.605 $Y=1.995
+ $X2=0.605 $Y2=2.57
r55 1 17 19.4347 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.5 $Y=1.58 $X2=0.5
+ $Y2=1.787
r56 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.5 $Y=1.58 $X2=0.5
+ $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_LP%A_28_148# 1 2 9 12 16 20 22 23 27 30
c45 27 0 7.36295e-20 $X=1.34 $Y=1.435
r46 27 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=1.435
+ $X2=1.34 $Y2=1.27
r47 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.34
+ $Y=1.435 $X2=1.34 $Y2=1.435
r48 23 26 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.34 $Y=1.315
+ $X2=1.34 $Y2=1.435
r49 21 22 3.66292 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=1.315
+ $X2=0.285 $Y2=1.315
r50 20 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=1.315
+ $X2=1.34 $Y2=1.315
r51 20 21 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.175 $Y=1.315
+ $X2=0.45 $Y2=1.315
r52 16 18 25.8827 $w=3.03e-07 $l=6.85e-07 $layer=LI1_cond $X=0.272 $Y=2.215
+ $X2=0.272 $Y2=2.9
r53 14 22 2.99104 $w=3.17e-07 $l=9.12688e-08 $layer=LI1_cond $X=0.272 $Y=1.4
+ $X2=0.285 $Y2=1.315
r54 14 16 30.7948 $w=3.03e-07 $l=8.15e-07 $layer=LI1_cond $X=0.272 $Y=1.4
+ $X2=0.272 $Y2=2.215
r55 10 22 2.99104 $w=3.17e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=1.23
+ $X2=0.285 $Y2=1.315
r56 10 12 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.285 $Y=1.23
+ $X2=0.285 $Y2=0.95
r57 9 30 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.345 $Y=0.95
+ $X2=1.345 $Y2=1.27
r58 2 18 400 $w=1.7e-07 $l=8.99583e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=2.07 $X2=0.34 $Y2=2.9
r59 2 16 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=2.07 $X2=0.34 $Y2=2.215
r60 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.74 $X2=0.285 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_LP%A 1 3 7 10 12 13 19
r29 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.945
+ $Y=0.465 $X2=1.945 $Y2=0.465
r30 16 19 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.82 $Y=0.465
+ $X2=1.945 $Y2=0.465
r31 13 20 8.89153 $w=2.95e-07 $l=2.15e-07 $layer=LI1_cond $X=2.16 $Y=0.485
+ $X2=1.945 $Y2=0.485
r32 12 20 10.9593 $w=2.95e-07 $l=2.65e-07 $layer=LI1_cond $X=1.68 $Y=0.485
+ $X2=1.945 $Y2=0.485
r33 5 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.82 $Y=1.84 $X2=1.82
+ $Y2=1.915
r34 5 7 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.82 $Y=1.84 $X2=1.82
+ $Y2=0.95
r35 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=0.63
+ $X2=1.82 $Y2=0.465
r36 4 7 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.82 $Y=0.63 $X2=1.82
+ $Y2=0.95
r37 1 10 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=1.625 $Y=1.915
+ $X2=1.82 $Y2=1.915
r38 1 3 111.824 $w=2.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.625 $Y=1.99
+ $X2=1.625 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_LP%VPWR 1 8 10 17 18 21
r21 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r22 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r23 14 17 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r24 12 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.87 $Y2=3.33
r25 12 14 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.2 $Y2=3.33
r26 10 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 10 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r29 6 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=3.245 $X2=0.87
+ $Y2=3.33
r30 6 8 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.87 $Y=3.245 $X2=0.87
+ $Y2=2.495
r31 1 8 300 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=2 $X=0.73
+ $Y=2.07 $X2=0.87 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_LP%Z 1 2 7 8 9 10 11 17
r17 11 29 2.71836 $w=5.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2 $Y=2.775 $X2=2
+ $Y2=2.9
r18 10 11 8.04635 $w=5.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2 $Y=2.405 $X2=2
+ $Y2=2.775
r19 10 23 4.13191 $w=5.48e-07 $l=1.9e-07 $layer=LI1_cond $X=2 $Y=2.405 $X2=2
+ $Y2=2.215
r20 9 23 3.91444 $w=5.48e-07 $l=1.8e-07 $layer=LI1_cond $X=2 $Y=2.035 $X2=2
+ $Y2=2.215
r21 8 9 8.04635 $w=5.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2 $Y=1.665 $X2=2
+ $Y2=2.035
r22 8 17 4.56684 $w=5.48e-07 $l=2.1e-07 $layer=LI1_cond $X=2 $Y=1.665 $X2=2
+ $Y2=1.455
r23 7 17 3.63656 $w=5.5e-07 $l=1.6e-07 $layer=LI1_cond $X=2 $Y=1.295 $X2=2
+ $Y2=1.455
r24 7 32 6.7112 $w=5.09e-07 $l=2.8e-07 $layer=LI1_cond $X=2 $Y=1.295 $X2=2
+ $Y2=1.015
r25 2 29 400 $w=1.7e-07 $l=8.97274e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=2.07 $X2=1.89 $Y2=2.9
r26 2 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=2.07 $X2=1.89 $Y2=2.215
r27 1 32 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.74 $X2=2.035 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_LP%VGND 1 6 8 10 17 18 21
r26 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.075
+ $Y2=0
r28 15 17 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=2.16
+ $Y2=0
r29 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.075
+ $Y2=0
r31 10 12 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.72
+ $Y2=0
r32 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r33 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r34 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.075 $Y=0.085
+ $X2=1.075 $Y2=0
r36 4 6 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=1.075 $Y=0.085 $X2=1.075
+ $Y2=0.885
r37 1 6 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.935
+ $Y=0.74 $X2=1.075 $Y2=0.885
.ends

