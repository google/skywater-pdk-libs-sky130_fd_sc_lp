* File: sky130_fd_sc_lp__lsbuf_lp.spice
* Created: Wed Sep  2 09:58:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__lsbuf_lp.pex.spice"
.subckt sky130_fd_sc_lp__lsbuf_lp  VGND VPB DESTVPB A VPWR DESTPWR X
* 
* X	X
* DESTPWR	DESTPWR
* VPWR	VPWR
* A	A
* DESTVPB	DESTVPB
* VPB	VPB
* VGND	VGND
MM1011 A_206_446# N_A_M1011_g N_VGND_M1011_s N_VGND_M1011_b NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 A_276_718# N_A_M1010_g N_A_193_718#_M1010_s N_VGND_M1011_b NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1008 N_A_278_47#_M1008_d N_A_M1008_g A_206_446# N_VGND_M1011_b NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g A_276_718# N_VGND_M1011_b NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.0882 PD=1.12 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1007 A_434_718# N_A_278_47#_M1007_g N_VGND_M1005_d N_VGND_M1011_b NSHORT
+ L=0.15 W=0.84 AD=0.0882 AS=0.1176 PD=1.05 PS=1.12 NRD=7.14 NRS=0 M=1 R=5.6
+ SA=75001 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1002 N_A_246_987#_M1002_d N_A_278_47#_M1002_g A_434_718# N_VGND_M1011_b NSHORT
+ L=0.15 W=0.84 AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6
+ SA=75001.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 A_712_718# N_A_193_718#_M1000_g N_VGND_M1000_s N_VGND_M1011_b NSHORT
+ L=0.15 W=0.84 AD=0.0882 AS=0.2394 PD=1.05 PS=2.25 NRD=7.14 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1013 N_X_M1013_d N_A_193_718#_M1013_g A_712_718# N_VGND_M1011_b NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 A_206_47# N_A_M1009_g N_VPWR_M1009_s N_VPB_M1009_b PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.5 A=0.15 P=2.3 MULT=1
MM1014 A_276_1085# N_A_246_987#_M1014_g N_A_193_718#_M1014_s N_DESTVPB_M1014_b
+ PHIGHVT L=0.15 W=1 AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=9.8303 NRS=0 M=1
+ R=6.66667 SA=75000.2 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1001 N_A_278_47#_M1001_d N_A_M1001_g A_206_47# N_VPB_M1009_b PHIGHVT L=0.15
+ W=1 AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667
+ SA=75000.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1015 N_DESTPWR_M1015_d N_A_246_987#_M1015_g A_276_1085# N_DESTVPB_M1014_b
+ PHIGHVT L=0.15 W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=9.8303 M=1
+ R=6.66667 SA=75000.5 SB=75001 A=0.15 P=2.3 MULT=1
MM1006 A_434_1085# N_A_193_718#_M1006_g N_DESTPWR_M1015_d N_DESTVPB_M1014_b
+ PHIGHVT L=0.15 W=1 AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=9.8303 NRS=0 M=1
+ R=6.66667 SA=75001 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1012 N_A_246_987#_M1012_d N_A_193_718#_M1012_g A_434_1085# N_DESTVPB_M1014_b
+ PHIGHVT L=0.15 W=1 AD=0.285 AS=0.105 PD=2.57 PS=1.21 NRD=0 NRS=9.8303 M=1
+ R=6.66667 SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1004 A_712_1085# N_A_193_718#_M1004_g N_DESTPWR_M1004_s N_DESTVPB_M1014_b
+ PHIGHVT L=0.15 W=1 AD=0.105 AS=0.285 PD=1.21 PS=2.57 NRD=9.8303 NRS=0 M=1
+ R=6.66667 SA=75000.2 SB=75000.5 A=0.15 P=2.3 MULT=1
MM1003 N_X_M1003_d N_A_193_718#_M1003_g A_712_1085# N_DESTVPB_M1014_b PHIGHVT
+ L=0.15 W=1 AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667
+ SA=75000.6 SB=75000.2 A=0.15 P=2.3 MULT=1
DX16_noxref N_VGND_M1011_b N_VPB_M1009_b NWDIODE A=9.04525 P=13.43
DX17_noxref N_VGND_M1011_b N_DESTVPB_M1014_b NWDIODE A=9.04525 P=13.43
*
.include "sky130_fd_sc_lp__lsbuf_lp.pxi.spice"
*
.ends
*
*
