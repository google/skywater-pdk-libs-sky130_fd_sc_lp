* File: sky130_fd_sc_lp__dfxbp_1.pxi.spice
* Created: Wed Sep  2 09:44:47 2020
* 
x_PM_SKY130_FD_SC_LP__DFXBP_1%CLK N_CLK_c_181_n N_CLK_M1004_g N_CLK_M1026_g
+ N_CLK_c_183_n CLK CLK CLK CLK N_CLK_c_185_n N_CLK_c_186_n
+ PM_SKY130_FD_SC_LP__DFXBP_1%CLK
x_PM_SKY130_FD_SC_LP__DFXBP_1%D N_D_M1023_g N_D_M1022_g N_D_c_210_n N_D_c_214_n
+ D D D N_D_c_212_n PM_SKY130_FD_SC_LP__DFXBP_1%D
x_PM_SKY130_FD_SC_LP__DFXBP_1%A_217_463# N_A_217_463#_M1008_s
+ N_A_217_463#_M1002_s N_A_217_463#_M1027_g N_A_217_463#_M1014_g
+ N_A_217_463#_M1018_g N_A_217_463#_c_253_n N_A_217_463#_M1019_g
+ N_A_217_463#_c_262_n N_A_217_463#_c_263_n N_A_217_463#_c_254_n
+ N_A_217_463#_c_265_n N_A_217_463#_c_266_n N_A_217_463#_c_267_n
+ N_A_217_463#_c_268_n N_A_217_463#_c_269_n N_A_217_463#_c_324_p
+ N_A_217_463#_c_270_n N_A_217_463#_c_255_n N_A_217_463#_c_272_n
+ N_A_217_463#_c_273_n N_A_217_463#_c_326_p N_A_217_463#_c_256_n
+ N_A_217_463#_c_257_n PM_SKY130_FD_SC_LP__DFXBP_1%A_217_463#
x_PM_SKY130_FD_SC_LP__DFXBP_1%A_697_93# N_A_697_93#_M1024_d N_A_697_93#_M1013_d
+ N_A_697_93#_c_418_n N_A_697_93#_M1005_g N_A_697_93#_M1001_g
+ N_A_697_93#_c_425_n N_A_697_93#_c_426_n N_A_697_93#_c_419_n
+ N_A_697_93#_c_420_n N_A_697_93#_c_421_n N_A_697_93#_c_422_n
+ N_A_697_93#_c_423_n PM_SKY130_FD_SC_LP__DFXBP_1%A_697_93#
x_PM_SKY130_FD_SC_LP__DFXBP_1%A_526_463# N_A_526_463#_M1010_d
+ N_A_526_463#_M1027_d N_A_526_463#_M1024_g N_A_526_463#_M1013_g
+ N_A_526_463#_c_495_n N_A_526_463#_c_489_n N_A_526_463#_c_490_n
+ N_A_526_463#_c_517_n N_A_526_463#_c_491_n N_A_526_463#_c_492_n
+ N_A_526_463#_c_493_n PM_SKY130_FD_SC_LP__DFXBP_1%A_526_463#
x_PM_SKY130_FD_SC_LP__DFXBP_1%A_110_82# N_A_110_82#_M1004_d N_A_110_82#_M1026_d
+ N_A_110_82#_c_570_n N_A_110_82#_c_571_n N_A_110_82#_M1002_g
+ N_A_110_82#_M1008_g N_A_110_82#_c_586_n N_A_110_82#_c_587_n
+ N_A_110_82#_c_574_n N_A_110_82#_c_575_n N_A_110_82#_M1010_g
+ N_A_110_82#_c_577_n N_A_110_82#_M1016_g N_A_110_82#_c_589_n
+ N_A_110_82#_M1025_g N_A_110_82#_M1000_g N_A_110_82#_c_579_n
+ N_A_110_82#_c_580_n N_A_110_82#_c_591_n N_A_110_82#_c_592_n
+ N_A_110_82#_c_593_n N_A_110_82#_c_581_n N_A_110_82#_c_582_n
+ N_A_110_82#_c_594_n N_A_110_82#_c_583_n N_A_110_82#_c_584_n
+ N_A_110_82#_c_596_n PM_SKY130_FD_SC_LP__DFXBP_1%A_110_82#
x_PM_SKY130_FD_SC_LP__DFXBP_1%A_1149_93# N_A_1149_93#_M1006_d
+ N_A_1149_93#_M1020_d N_A_1149_93#_c_708_n N_A_1149_93#_M1009_g
+ N_A_1149_93#_c_709_n N_A_1149_93#_M1003_g N_A_1149_93#_c_710_n
+ N_A_1149_93#_M1011_g N_A_1149_93#_M1021_g N_A_1149_93#_c_711_n
+ N_A_1149_93#_M1015_g N_A_1149_93#_M1017_g N_A_1149_93#_c_712_n
+ N_A_1149_93#_c_713_n N_A_1149_93#_c_714_n N_A_1149_93#_c_724_n
+ N_A_1149_93#_c_715_n N_A_1149_93#_c_716_n N_A_1149_93#_c_725_n
+ N_A_1149_93#_c_726_n N_A_1149_93#_c_727_n N_A_1149_93#_c_728_n
+ N_A_1149_93#_c_717_n N_A_1149_93#_c_718_n
+ PM_SKY130_FD_SC_LP__DFXBP_1%A_1149_93#
x_PM_SKY130_FD_SC_LP__DFXBP_1%A_997_119# N_A_997_119#_M1018_d
+ N_A_997_119#_M1025_d N_A_997_119#_M1006_g N_A_997_119#_M1020_g
+ N_A_997_119#_c_838_n N_A_997_119#_c_839_n N_A_997_119#_c_831_n
+ N_A_997_119#_c_832_n N_A_997_119#_c_833_n N_A_997_119#_c_834_n
+ N_A_997_119#_c_835_n N_A_997_119#_c_836_n
+ PM_SKY130_FD_SC_LP__DFXBP_1%A_997_119#
x_PM_SKY130_FD_SC_LP__DFXBP_1%A_1401_22# N_A_1401_22#_M1011_s
+ N_A_1401_22#_M1021_s N_A_1401_22#_c_902_n N_A_1401_22#_c_903_n
+ N_A_1401_22#_M1012_g N_A_1401_22#_M1007_g N_A_1401_22#_c_905_n
+ N_A_1401_22#_c_906_n N_A_1401_22#_c_907_n N_A_1401_22#_c_908_n
+ N_A_1401_22#_c_909_n N_A_1401_22#_c_912_n
+ PM_SKY130_FD_SC_LP__DFXBP_1%A_1401_22#
x_PM_SKY130_FD_SC_LP__DFXBP_1%VPWR N_VPWR_M1026_s N_VPWR_M1002_d N_VPWR_M1001_d
+ N_VPWR_M1003_d N_VPWR_M1021_d N_VPWR_M1017_s N_VPWR_c_967_n N_VPWR_c_968_n
+ N_VPWR_c_969_n N_VPWR_c_970_n N_VPWR_c_971_n N_VPWR_c_972_n N_VPWR_c_973_n
+ N_VPWR_c_974_n N_VPWR_c_975_n N_VPWR_c_976_n VPWR N_VPWR_c_977_n
+ N_VPWR_c_978_n N_VPWR_c_979_n N_VPWR_c_980_n N_VPWR_c_966_n N_VPWR_c_982_n
+ N_VPWR_c_983_n N_VPWR_c_984_n N_VPWR_c_985_n PM_SKY130_FD_SC_LP__DFXBP_1%VPWR
x_PM_SKY130_FD_SC_LP__DFXBP_1%A_440_463# N_A_440_463#_M1022_d
+ N_A_440_463#_M1023_d N_A_440_463#_c_1064_n N_A_440_463#_c_1070_n
+ PM_SKY130_FD_SC_LP__DFXBP_1%A_440_463#
x_PM_SKY130_FD_SC_LP__DFXBP_1%Q_N N_Q_N_M1012_d N_Q_N_M1007_d Q_N Q_N Q_N Q_N
+ N_Q_N_c_1084_n PM_SKY130_FD_SC_LP__DFXBP_1%Q_N
x_PM_SKY130_FD_SC_LP__DFXBP_1%Q N_Q_M1015_d N_Q_M1017_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DFXBP_1%Q
x_PM_SKY130_FD_SC_LP__DFXBP_1%VGND N_VGND_M1004_s N_VGND_M1008_d N_VGND_M1005_d
+ N_VGND_M1009_d N_VGND_M1011_d N_VGND_M1015_s N_VGND_c_1108_n N_VGND_c_1109_n
+ N_VGND_c_1110_n N_VGND_c_1111_n N_VGND_c_1112_n N_VGND_c_1113_n
+ N_VGND_c_1114_n N_VGND_c_1115_n N_VGND_c_1116_n N_VGND_c_1117_n
+ N_VGND_c_1118_n VGND N_VGND_c_1119_n N_VGND_c_1120_n N_VGND_c_1121_n
+ N_VGND_c_1122_n N_VGND_c_1123_n N_VGND_c_1124_n N_VGND_c_1125_n
+ N_VGND_c_1126_n PM_SKY130_FD_SC_LP__DFXBP_1%VGND
cc_1 VNB N_CLK_c_181_n 0.0258149f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.423
cc_2 VNB N_CLK_M1026_g 0.00272334f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_3 VNB N_CLK_c_183_n 0.0225363f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.61
cc_4 VNB CLK 0.0333978f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_CLK_c_185_n 0.0235693f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.105
cc_6 VNB N_CLK_c_186_n 0.0232437f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=0.94
cc_7 VNB N_D_M1022_g 0.0216572f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_8 VNB N_D_c_210_n 0.0382701f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB D 0.0110089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_D_c_212_n 0.0229021f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_11 VNB N_A_217_463#_M1014_g 0.0459739f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_A_217_463#_M1018_g 0.0233362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_217_463#_c_253_n 0.0363475f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.105
cc_14 VNB N_A_217_463#_c_254_n 0.00565121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_217_463#_c_255_n 0.00164299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_217_463#_c_256_n 0.00252178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_217_463#_c_257_n 0.0365912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_697_93#_c_418_n 0.0161649f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_19 VNB N_A_697_93#_c_419_n 0.00923025f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_20 VNB N_A_697_93#_c_420_n 0.0017708f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.295
cc_21 VNB N_A_697_93#_c_421_n 0.00229537f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_22 VNB N_A_697_93#_c_422_n 0.0106122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_697_93#_c_423_n 0.0382474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_526_463#_M1024_g 0.0207253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_526_463#_c_489_n 0.00742147f $X=-0.19 $Y=-0.245 $X2=0.362
+ $Y2=1.105
cc_26 VNB N_A_526_463#_c_490_n 0.00645847f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=0.94
cc_27 VNB N_A_526_463#_c_491_n 0.00402353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_526_463#_c_492_n 0.0221756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_526_463#_c_493_n 0.0118505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_110_82#_c_570_n 0.0138954f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_31 VNB N_A_110_82#_c_571_n 0.0185408f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_32 VNB N_A_110_82#_M1002_g 0.0136875f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_33 VNB N_A_110_82#_M1008_g 0.0404758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_110_82#_c_574_n 0.0793586f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.105
cc_35 VNB N_A_110_82#_c_575_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.105
cc_36 VNB N_A_110_82#_M1010_g 0.0383741f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_37 VNB N_A_110_82#_c_577_n 0.199944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_110_82#_M1000_g 0.034638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_110_82#_c_579_n 0.0159677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_110_82#_c_580_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_110_82#_c_581_n 0.0136128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_110_82#_c_582_n 0.00132319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_110_82#_c_583_n 0.00802094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_110_82#_c_584_n 0.0178338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1149_93#_c_708_n 0.0188136f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_46 VNB N_A_1149_93#_c_709_n 0.0546827f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.61
cc_47 VNB N_A_1149_93#_c_710_n 0.0188945f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_48 VNB N_A_1149_93#_c_711_n 0.0213689f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.105
cc_49 VNB N_A_1149_93#_c_712_n 0.0536772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1149_93#_c_713_n 0.0151489f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_51 VNB N_A_1149_93#_c_714_n 0.0025344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1149_93#_c_715_n 0.0116436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1149_93#_c_716_n 0.00741052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1149_93#_c_717_n 0.0212459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1149_93#_c_718_n 0.0406543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_997_119#_M1020_g 0.0109374f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_57 VNB N_A_997_119#_c_831_n 0.00252575f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.105
cc_58 VNB N_A_997_119#_c_832_n 0.0250537f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=0.94
cc_59 VNB N_A_997_119#_c_833_n 0.00300456f $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=1.295
cc_60 VNB N_A_997_119#_c_834_n 0.00185087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_997_119#_c_835_n 0.0341773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_997_119#_c_836_n 0.0202718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1401_22#_c_902_n 0.0655262f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_64 VNB N_A_1401_22#_c_903_n 0.0214302f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_65 VNB N_A_1401_22#_M1012_g 0.0348495f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_66 VNB N_A_1401_22#_c_905_n 0.00447349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1401_22#_c_906_n 0.00122914f $X=-0.19 $Y=-0.245 $X2=0.362
+ $Y2=1.105
cc_68 VNB N_A_1401_22#_c_907_n 0.0430358f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=0.94
cc_69 VNB N_A_1401_22#_c_908_n 0.00477366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1401_22#_c_909_n 0.00278683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VPWR_c_966_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_440_463#_c_1064_n 0.0117125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_Q_N_c_1084_n 0.0231091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB Q 0.0577545f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_75 VNB N_VGND_c_1108_n 0.0115788f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.105
cc_76 VNB N_VGND_c_1109_n 0.0235691f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.105
cc_77 VNB N_VGND_c_1110_n 0.0104291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1111_n 0.0194616f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_79 VNB N_VGND_c_1112_n 0.0135165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1113_n 0.0197892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1114_n 0.0195566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1115_n 0.0385116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1116_n 0.00426141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1117_n 0.0506667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1118_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1119_n 0.0433858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1120_n 0.0376879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1121_n 0.0176971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1122_n 0.0187657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1123_n 0.514705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1124_n 0.00965476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1125_n 0.00418557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1126_n 0.00519339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VPB N_CLK_M1026_g 0.0629221f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_95 VPB CLK 0.023901f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_96 VPB N_D_M1023_g 0.0350245f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.94
cc_97 VPB N_D_c_214_n 0.0207993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB D 0.00873157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_D_c_212_n 0.00289276f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_100 VPB N_A_217_463#_M1027_g 0.0204348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_217_463#_M1014_g 0.0107243f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_102 VPB N_A_217_463#_c_253_n 0.00656602f $X=-0.19 $Y=1.655 $X2=0.362
+ $Y2=1.105
cc_103 VPB N_A_217_463#_M1019_g 0.0258157f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_104 VPB N_A_217_463#_c_262_n 0.0193986f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_217_463#_c_263_n 0.0571006f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.105
cc_106 VPB N_A_217_463#_c_254_n 0.00574356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_217_463#_c_265_n 6.22156e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_217_463#_c_266_n 8.79799e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_217_463#_c_267_n 0.0208649f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_217_463#_c_268_n 0.00164809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_217_463#_c_269_n 0.00449348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_217_463#_c_270_n 0.00202686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_217_463#_c_255_n 0.00351589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_217_463#_c_272_n 0.013809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_217_463#_c_273_n 0.00195066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_697_93#_M1001_g 0.0216538f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_117 VPB N_A_697_93#_c_425_n 0.0313829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_697_93#_c_426_n 0.00705916f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.105
cc_119 VPB N_A_697_93#_c_422_n 0.00977617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_526_463#_M1013_g 0.0226717f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_121 VPB N_A_526_463#_c_495_n 0.00420899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_526_463#_c_490_n 0.00330586f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=0.94
cc_123 VPB N_A_526_463#_c_491_n 9.27686e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_526_463#_c_492_n 0.010629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_526_463#_c_493_n 0.0108555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_110_82#_M1002_g 0.0518063f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_127 VPB N_A_110_82#_c_586_n 0.110269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_110_82#_c_587_n 0.0126359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_110_82#_M1016_g 0.0206395f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.665
cc_130 VPB N_A_110_82#_c_589_n 0.139463f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=2.035
cc_131 VPB N_A_110_82#_M1025_g 0.0444854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_110_82#_c_591_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_110_82#_c_592_n 0.0018152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_110_82#_c_593_n 0.00223325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_110_82#_c_594_n 0.00930579f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_110_82#_c_584_n 0.0239365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_110_82#_c_596_n 0.0112791f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_1149_93#_c_709_n 0.0100678f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.61
cc_139 VPB N_A_1149_93#_M1003_g 0.0219158f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_140 VPB N_A_1149_93#_M1021_g 0.0259202f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.105
cc_141 VPB N_A_1149_93#_M1017_g 0.0251997f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.105
cc_142 VPB N_A_1149_93#_c_714_n 0.00271448f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_1149_93#_c_724_n 0.0098419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_1149_93#_c_725_n 0.0329717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_1149_93#_c_726_n 0.014557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_1149_93#_c_727_n 0.00832627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_1149_93#_c_728_n 0.00279688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_1149_93#_c_717_n 0.00186203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_1149_93#_c_718_n 0.0113933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_997_119#_M1020_g 0.0298434f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_151 VPB N_A_997_119#_c_838_n 0.00124651f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_152 VPB N_A_997_119#_c_839_n 0.0102183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_997_119#_c_833_n 0.00381825f $X=-0.19 $Y=1.655 $X2=0.255
+ $Y2=1.295
cc_154 VPB N_A_1401_22#_M1012_g 0.0258855f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_155 VPB N_A_1401_22#_c_906_n 0.00233933f $X=-0.19 $Y=1.655 $X2=0.362
+ $Y2=1.105
cc_156 VPB N_A_1401_22#_c_912_n 0.00408125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_967_n 0.0108797f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.105
cc_158 VPB N_VPWR_c_968_n 0.0399719f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.105
cc_159 VPB N_VPWR_c_969_n 0.00159471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_970_n 0.0142103f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.665
cc_161 VPB N_VPWR_c_971_n 0.0396373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_972_n 0.0176656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_973_n 0.0208467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_974_n 0.00495479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_975_n 0.0523199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_976_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_977_n 0.0300879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_978_n 0.0526134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_979_n 0.0422123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_980_n 0.0182379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_966_n 0.107027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_982_n 0.00317016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_983_n 0.00436716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_984_n 0.00510939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_985_n 0.00401177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_440_463#_c_1064_n 0.0127221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_Q_N_c_1084_n 0.00848805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB Q 0.05656f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_179 N_CLK_c_181_n N_A_110_82#_c_571_n 0.0170892f $X=0.362 $Y=1.423 $X2=0
+ $Y2=0
cc_180 CLK N_A_110_82#_c_571_n 5.02322e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_181 N_CLK_M1026_g N_A_110_82#_c_592_n 6.96261e-19 $X=0.475 $Y=2.66 $X2=0
+ $Y2=0
cc_182 CLK N_A_110_82#_c_581_n 0.103665f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_183 N_CLK_c_186_n N_A_110_82#_c_581_n 0.00566627f $X=0.362 $Y=0.94 $X2=0
+ $Y2=0
cc_184 N_CLK_c_181_n N_A_110_82#_c_582_n 0.00566627f $X=0.362 $Y=1.423 $X2=0
+ $Y2=0
cc_185 N_CLK_M1026_g N_A_110_82#_c_594_n 0.00566627f $X=0.475 $Y=2.66 $X2=0
+ $Y2=0
cc_186 N_CLK_c_185_n N_A_110_82#_c_583_n 0.00566627f $X=0.34 $Y=1.105 $X2=0
+ $Y2=0
cc_187 N_CLK_c_183_n N_A_110_82#_c_584_n 0.0170892f $X=0.362 $Y=1.61 $X2=0 $Y2=0
cc_188 N_CLK_c_183_n N_A_110_82#_c_596_n 0.00566627f $X=0.362 $Y=1.61 $X2=0
+ $Y2=0
cc_189 N_CLK_M1026_g N_VPWR_c_968_n 0.00577183f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_190 CLK N_VPWR_c_968_n 0.0274534f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_191 N_CLK_M1026_g N_VPWR_c_977_n 0.00478016f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_192 N_CLK_M1026_g N_VPWR_c_966_n 0.00978454f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_193 CLK N_VGND_c_1109_n 0.0266998f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_194 N_CLK_c_185_n N_VGND_c_1109_n 0.0012272f $X=0.34 $Y=1.105 $X2=0 $Y2=0
cc_195 N_CLK_c_186_n N_VGND_c_1109_n 0.0131656f $X=0.362 $Y=0.94 $X2=0 $Y2=0
cc_196 N_CLK_c_186_n N_VGND_c_1115_n 0.00455951f $X=0.362 $Y=0.94 $X2=0 $Y2=0
cc_197 CLK N_VGND_c_1123_n 0.0015796f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_198 N_CLK_c_186_n N_VGND_c_1123_n 0.00447788f $X=0.362 $Y=0.94 $X2=0 $Y2=0
cc_199 N_D_M1023_g N_A_217_463#_M1027_g 0.0129178f $X=2.125 $Y=2.525 $X2=0 $Y2=0
cc_200 N_D_M1022_g N_A_217_463#_M1014_g 0.00200785f $X=2.34 $Y=0.805 $X2=0 $Y2=0
cc_201 N_D_c_214_n N_A_217_463#_c_262_n 0.0129178f $X=2.012 $Y=1.88 $X2=0 $Y2=0
cc_202 N_D_M1023_g N_A_217_463#_c_254_n 8.54962e-19 $X=2.125 $Y=2.525 $X2=0
+ $Y2=0
cc_203 N_D_c_210_n N_A_217_463#_c_254_n 5.01242e-19 $X=2.34 $Y=1.285 $X2=0 $Y2=0
cc_204 D N_A_217_463#_c_254_n 0.0732464f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_205 N_D_M1023_g N_A_217_463#_c_265_n 0.00522547f $X=2.125 $Y=2.525 $X2=0
+ $Y2=0
cc_206 N_D_c_214_n N_A_217_463#_c_265_n 8.34593e-19 $X=2.012 $Y=1.88 $X2=0 $Y2=0
cc_207 D N_A_217_463#_c_265_n 0.0388579f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_208 N_D_M1023_g N_A_217_463#_c_266_n 0.00960633f $X=2.125 $Y=2.525 $X2=0
+ $Y2=0
cc_209 N_D_M1023_g N_A_217_463#_c_267_n 0.00337338f $X=2.125 $Y=2.525 $X2=0
+ $Y2=0
cc_210 N_D_M1023_g N_A_217_463#_c_268_n 2.20287e-19 $X=2.125 $Y=2.525 $X2=0
+ $Y2=0
cc_211 N_D_M1022_g N_A_526_463#_c_489_n 9.86949e-19 $X=2.34 $Y=0.805 $X2=0 $Y2=0
cc_212 N_D_M1023_g N_A_110_82#_M1002_g 0.0144855f $X=2.125 $Y=2.525 $X2=0 $Y2=0
cc_213 D N_A_110_82#_M1002_g 0.00668621f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_214 N_D_c_212_n N_A_110_82#_M1002_g 0.0169093f $X=1.99 $Y=1.375 $X2=0 $Y2=0
cc_215 N_D_M1022_g N_A_110_82#_M1008_g 0.00814899f $X=2.34 $Y=0.805 $X2=0 $Y2=0
cc_216 N_D_c_210_n N_A_110_82#_M1008_g 0.00503f $X=2.34 $Y=1.285 $X2=0 $Y2=0
cc_217 D N_A_110_82#_M1008_g 0.00124597f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_218 N_D_M1023_g N_A_110_82#_c_586_n 0.008966f $X=2.125 $Y=2.525 $X2=0 $Y2=0
cc_219 N_D_M1022_g N_A_110_82#_c_574_n 0.00978449f $X=2.34 $Y=0.805 $X2=0 $Y2=0
cc_220 N_D_M1022_g N_A_110_82#_M1010_g 0.0128449f $X=2.34 $Y=0.805 $X2=0 $Y2=0
cc_221 D N_A_110_82#_c_579_n 0.00446809f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_222 N_D_c_212_n N_A_110_82#_c_579_n 0.00503f $X=1.99 $Y=1.375 $X2=0 $Y2=0
cc_223 N_D_M1023_g N_VPWR_c_969_n 6.02314e-19 $X=2.125 $Y=2.525 $X2=0 $Y2=0
cc_224 N_D_M1022_g N_A_440_463#_c_1064_n 0.00791795f $X=2.34 $Y=0.805 $X2=0
+ $Y2=0
cc_225 N_D_c_210_n N_A_440_463#_c_1064_n 0.0105372f $X=2.34 $Y=1.285 $X2=0 $Y2=0
cc_226 D N_A_440_463#_c_1064_n 0.0723017f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_227 N_D_c_212_n N_A_440_463#_c_1064_n 0.0190257f $X=1.99 $Y=1.375 $X2=0 $Y2=0
cc_228 N_D_M1022_g N_A_440_463#_c_1070_n 0.0105946f $X=2.34 $Y=0.805 $X2=0 $Y2=0
cc_229 N_D_M1022_g N_VGND_c_1110_n 0.00591105f $X=2.34 $Y=0.805 $X2=0 $Y2=0
cc_230 N_D_c_210_n N_VGND_c_1110_n 0.00187654f $X=2.34 $Y=1.285 $X2=0 $Y2=0
cc_231 D N_VGND_c_1110_n 0.0219461f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_232 N_D_M1022_g N_VGND_c_1123_n 9.39239e-19 $X=2.34 $Y=0.805 $X2=0 $Y2=0
cc_233 N_A_217_463#_c_270_n N_A_697_93#_M1013_d 0.0172919f $X=4.865 $Y=2.5 $X2=0
+ $Y2=0
cc_234 N_A_217_463#_c_255_n N_A_697_93#_M1013_d 0.0056368f $X=4.95 $Y=2.415
+ $X2=0 $Y2=0
cc_235 N_A_217_463#_M1014_g N_A_697_93#_c_418_n 0.0590957f $X=3.2 $Y=0.805 $X2=0
+ $Y2=0
cc_236 N_A_217_463#_c_269_n N_A_697_93#_M1001_g 0.00516789f $X=3.215 $Y=2.415
+ $X2=0 $Y2=0
cc_237 N_A_217_463#_c_270_n N_A_697_93#_M1001_g 0.0129435f $X=4.865 $Y=2.5 $X2=0
+ $Y2=0
cc_238 N_A_217_463#_c_263_n N_A_697_93#_c_425_n 0.0213092f $X=3.125 $Y=1.99
+ $X2=0 $Y2=0
cc_239 N_A_217_463#_c_270_n N_A_697_93#_c_425_n 7.96576e-19 $X=4.865 $Y=2.5
+ $X2=0 $Y2=0
cc_240 N_A_217_463#_c_273_n N_A_697_93#_c_425_n 9.00155e-19 $X=3.215 $Y=2.025
+ $X2=0 $Y2=0
cc_241 N_A_217_463#_c_263_n N_A_697_93#_c_426_n 3.04749e-19 $X=3.125 $Y=1.99
+ $X2=0 $Y2=0
cc_242 N_A_217_463#_c_269_n N_A_697_93#_c_426_n 0.00605517f $X=3.215 $Y=2.415
+ $X2=0 $Y2=0
cc_243 N_A_217_463#_c_270_n N_A_697_93#_c_426_n 0.0747444f $X=4.865 $Y=2.5 $X2=0
+ $Y2=0
cc_244 N_A_217_463#_c_255_n N_A_697_93#_c_426_n 0.027499f $X=4.95 $Y=2.415 $X2=0
+ $Y2=0
cc_245 N_A_217_463#_c_273_n N_A_697_93#_c_426_n 0.0197092f $X=3.215 $Y=2.025
+ $X2=0 $Y2=0
cc_246 N_A_217_463#_M1018_g N_A_697_93#_c_419_n 0.00219379f $X=4.91 $Y=0.805
+ $X2=0 $Y2=0
cc_247 N_A_217_463#_c_256_n N_A_697_93#_c_419_n 0.0024515f $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_248 N_A_217_463#_M1018_g N_A_697_93#_c_420_n 0.00537708f $X=4.91 $Y=0.805
+ $X2=0 $Y2=0
cc_249 N_A_217_463#_M1014_g N_A_697_93#_c_421_n 9.00231e-19 $X=3.2 $Y=0.805
+ $X2=0 $Y2=0
cc_250 N_A_217_463#_M1014_g N_A_697_93#_c_422_n 0.0115062f $X=3.2 $Y=0.805 $X2=0
+ $Y2=0
cc_251 N_A_217_463#_c_267_n N_A_526_463#_M1027_d 0.00606583f $X=3.13 $Y=2.97
+ $X2=0 $Y2=0
cc_252 N_A_217_463#_M1018_g N_A_526_463#_M1024_g 0.0112984f $X=4.91 $Y=0.805
+ $X2=0 $Y2=0
cc_253 N_A_217_463#_c_256_n N_A_526_463#_M1024_g 9.8051e-19 $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_254 N_A_217_463#_c_270_n N_A_526_463#_M1013_g 0.0136635f $X=4.865 $Y=2.5
+ $X2=0 $Y2=0
cc_255 N_A_217_463#_c_255_n N_A_526_463#_M1013_g 0.00302014f $X=4.95 $Y=2.415
+ $X2=0 $Y2=0
cc_256 N_A_217_463#_M1027_g N_A_526_463#_c_495_n 0.00588126f $X=2.555 $Y=2.525
+ $X2=0 $Y2=0
cc_257 N_A_217_463#_M1014_g N_A_526_463#_c_495_n 0.00281318f $X=3.2 $Y=0.805
+ $X2=0 $Y2=0
cc_258 N_A_217_463#_c_262_n N_A_526_463#_c_495_n 0.00375549f $X=2.63 $Y=1.99
+ $X2=0 $Y2=0
cc_259 N_A_217_463#_c_263_n N_A_526_463#_c_495_n 0.0156177f $X=3.125 $Y=1.99
+ $X2=0 $Y2=0
cc_260 N_A_217_463#_c_269_n N_A_526_463#_c_495_n 0.00942883f $X=3.215 $Y=2.415
+ $X2=0 $Y2=0
cc_261 N_A_217_463#_c_273_n N_A_526_463#_c_495_n 0.0186297f $X=3.215 $Y=2.025
+ $X2=0 $Y2=0
cc_262 N_A_217_463#_M1014_g N_A_526_463#_c_489_n 0.0250473f $X=3.2 $Y=0.805
+ $X2=0 $Y2=0
cc_263 N_A_217_463#_M1014_g N_A_526_463#_c_490_n 0.00493873f $X=3.2 $Y=0.805
+ $X2=0 $Y2=0
cc_264 N_A_217_463#_c_262_n N_A_526_463#_c_490_n 7.97484e-19 $X=2.63 $Y=1.99
+ $X2=0 $Y2=0
cc_265 N_A_217_463#_c_263_n N_A_526_463#_c_490_n 0.00855999f $X=3.125 $Y=1.99
+ $X2=0 $Y2=0
cc_266 N_A_217_463#_c_273_n N_A_526_463#_c_490_n 0.0256699f $X=3.215 $Y=2.025
+ $X2=0 $Y2=0
cc_267 N_A_217_463#_M1027_g N_A_526_463#_c_517_n 0.0084155f $X=2.555 $Y=2.525
+ $X2=0 $Y2=0
cc_268 N_A_217_463#_c_263_n N_A_526_463#_c_517_n 0.00553428f $X=3.125 $Y=1.99
+ $X2=0 $Y2=0
cc_269 N_A_217_463#_c_267_n N_A_526_463#_c_517_n 0.0241152f $X=3.13 $Y=2.97
+ $X2=0 $Y2=0
cc_270 N_A_217_463#_c_269_n N_A_526_463#_c_517_n 0.00363146f $X=3.215 $Y=2.415
+ $X2=0 $Y2=0
cc_271 N_A_217_463#_c_324_p N_A_526_463#_c_517_n 0.00811983f $X=3.215 $Y=2.865
+ $X2=0 $Y2=0
cc_272 N_A_217_463#_c_273_n N_A_526_463#_c_517_n 9.72715e-19 $X=3.215 $Y=2.025
+ $X2=0 $Y2=0
cc_273 N_A_217_463#_c_326_p N_A_526_463#_c_517_n 0.0141544f $X=3.215 $Y=2.5
+ $X2=0 $Y2=0
cc_274 N_A_217_463#_c_256_n N_A_526_463#_c_491_n 0.0116923f $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_275 N_A_217_463#_c_257_n N_A_526_463#_c_491_n 6.3201e-19 $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_276 N_A_217_463#_c_255_n N_A_526_463#_c_492_n 0.00436395f $X=4.95 $Y=2.415
+ $X2=0 $Y2=0
cc_277 N_A_217_463#_c_257_n N_A_526_463#_c_492_n 0.0112984f $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_278 N_A_217_463#_M1014_g N_A_526_463#_c_493_n 0.0109425f $X=3.2 $Y=0.805
+ $X2=0 $Y2=0
cc_279 N_A_217_463#_c_254_n N_A_110_82#_c_570_n 0.00833681f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_280 N_A_217_463#_c_254_n N_A_110_82#_M1002_g 0.0241835f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_281 N_A_217_463#_c_265_n N_A_110_82#_M1002_g 0.00966381f $X=1.905 $Y=2.4
+ $X2=0 $Y2=0
cc_282 N_A_217_463#_c_266_n N_A_110_82#_M1002_g 0.00125737f $X=1.99 $Y=2.865
+ $X2=0 $Y2=0
cc_283 N_A_217_463#_c_268_n N_A_110_82#_M1002_g 7.40958e-19 $X=2.075 $Y=2.97
+ $X2=0 $Y2=0
cc_284 N_A_217_463#_c_272_n N_A_110_82#_M1002_g 0.00416435f $X=1.21 $Y=2.46
+ $X2=0 $Y2=0
cc_285 N_A_217_463#_c_254_n N_A_110_82#_M1008_g 0.00820761f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_286 N_A_217_463#_M1027_g N_A_110_82#_c_586_n 0.00881263f $X=2.555 $Y=2.525
+ $X2=0 $Y2=0
cc_287 N_A_217_463#_c_265_n N_A_110_82#_c_586_n 0.00420732f $X=1.905 $Y=2.4
+ $X2=0 $Y2=0
cc_288 N_A_217_463#_c_267_n N_A_110_82#_c_586_n 0.0175078f $X=3.13 $Y=2.97 $X2=0
+ $Y2=0
cc_289 N_A_217_463#_c_268_n N_A_110_82#_c_586_n 0.00378523f $X=2.075 $Y=2.97
+ $X2=0 $Y2=0
cc_290 N_A_217_463#_M1014_g N_A_110_82#_M1010_g 0.0131001f $X=3.2 $Y=0.805 $X2=0
+ $Y2=0
cc_291 N_A_217_463#_c_263_n N_A_110_82#_M1010_g 0.0017789f $X=3.125 $Y=1.99
+ $X2=0 $Y2=0
cc_292 N_A_217_463#_M1014_g N_A_110_82#_c_577_n 0.0102728f $X=3.2 $Y=0.805 $X2=0
+ $Y2=0
cc_293 N_A_217_463#_M1018_g N_A_110_82#_c_577_n 0.0104164f $X=4.91 $Y=0.805
+ $X2=0 $Y2=0
cc_294 N_A_217_463#_M1027_g N_A_110_82#_M1016_g 0.0106918f $X=2.555 $Y=2.525
+ $X2=0 $Y2=0
cc_295 N_A_217_463#_c_263_n N_A_110_82#_M1016_g 0.00998904f $X=3.125 $Y=1.99
+ $X2=0 $Y2=0
cc_296 N_A_217_463#_c_267_n N_A_110_82#_M1016_g 0.0125711f $X=3.13 $Y=2.97 $X2=0
+ $Y2=0
cc_297 N_A_217_463#_c_269_n N_A_110_82#_M1016_g 0.00221071f $X=3.215 $Y=2.415
+ $X2=0 $Y2=0
cc_298 N_A_217_463#_c_324_p N_A_110_82#_M1016_g 0.00811154f $X=3.215 $Y=2.865
+ $X2=0 $Y2=0
cc_299 N_A_217_463#_c_273_n N_A_110_82#_M1016_g 3.08802e-19 $X=3.215 $Y=2.025
+ $X2=0 $Y2=0
cc_300 N_A_217_463#_c_326_p N_A_110_82#_M1016_g 0.00525746f $X=3.215 $Y=2.5
+ $X2=0 $Y2=0
cc_301 N_A_217_463#_c_267_n N_A_110_82#_c_589_n 4.19731e-19 $X=3.13 $Y=2.97
+ $X2=0 $Y2=0
cc_302 N_A_217_463#_c_270_n N_A_110_82#_c_589_n 0.0159993f $X=4.865 $Y=2.5 $X2=0
+ $Y2=0
cc_303 N_A_217_463#_M1019_g N_A_110_82#_M1025_g 0.0109703f $X=5.61 $Y=2.105
+ $X2=0 $Y2=0
cc_304 N_A_217_463#_c_270_n N_A_110_82#_M1025_g 0.00558655f $X=4.865 $Y=2.5
+ $X2=0 $Y2=0
cc_305 N_A_217_463#_c_255_n N_A_110_82#_M1025_g 0.0149361f $X=4.95 $Y=2.415
+ $X2=0 $Y2=0
cc_306 N_A_217_463#_c_256_n N_A_110_82#_M1025_g 4.54815e-19 $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_307 N_A_217_463#_c_257_n N_A_110_82#_M1025_g 0.0107853f $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_308 N_A_217_463#_M1018_g N_A_110_82#_M1000_g 0.0147702f $X=4.91 $Y=0.805
+ $X2=0 $Y2=0
cc_309 N_A_217_463#_c_253_n N_A_110_82#_M1000_g 0.00727039f $X=5.385 $Y=1.48
+ $X2=0 $Y2=0
cc_310 N_A_217_463#_c_254_n N_A_110_82#_c_579_n 0.00450737f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_311 N_A_217_463#_c_267_n N_A_110_82#_c_591_n 0.00102791f $X=3.13 $Y=2.97
+ $X2=0 $Y2=0
cc_312 N_A_217_463#_c_272_n N_A_110_82#_c_593_n 0.0286402f $X=1.21 $Y=2.46 $X2=0
+ $Y2=0
cc_313 N_A_217_463#_c_254_n N_A_110_82#_c_581_n 0.0279798f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_314 N_A_217_463#_c_254_n N_A_110_82#_c_594_n 0.0171021f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_315 N_A_217_463#_c_272_n N_A_110_82#_c_594_n 0.0121643f $X=1.21 $Y=2.46 $X2=0
+ $Y2=0
cc_316 N_A_217_463#_c_254_n N_A_110_82#_c_583_n 0.0516544f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_317 N_A_217_463#_c_254_n N_A_110_82#_c_584_n 0.00345003f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_318 N_A_217_463#_c_272_n N_A_110_82#_c_584_n 0.00276968f $X=1.21 $Y=2.46
+ $X2=0 $Y2=0
cc_319 N_A_217_463#_c_253_n N_A_1149_93#_c_709_n 0.0321884f $X=5.385 $Y=1.48
+ $X2=0 $Y2=0
cc_320 N_A_217_463#_c_257_n N_A_1149_93#_c_709_n 6.85733e-19 $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_321 N_A_217_463#_M1019_g N_A_1149_93#_M1003_g 0.0278103f $X=5.61 $Y=2.105
+ $X2=0 $Y2=0
cc_322 N_A_217_463#_c_253_n N_A_1149_93#_c_728_n 0.00126605f $X=5.385 $Y=1.48
+ $X2=0 $Y2=0
cc_323 N_A_217_463#_c_253_n N_A_997_119#_c_838_n 0.00206676f $X=5.385 $Y=1.48
+ $X2=0 $Y2=0
cc_324 N_A_217_463#_c_255_n N_A_997_119#_c_838_n 0.0190293f $X=4.95 $Y=2.415
+ $X2=0 $Y2=0
cc_325 N_A_217_463#_M1018_g N_A_997_119#_c_831_n 0.00310273f $X=4.91 $Y=0.805
+ $X2=0 $Y2=0
cc_326 N_A_217_463#_c_253_n N_A_997_119#_c_831_n 0.00289635f $X=5.385 $Y=1.48
+ $X2=0 $Y2=0
cc_327 N_A_217_463#_c_256_n N_A_997_119#_c_831_n 0.0100408f $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_328 N_A_217_463#_c_257_n N_A_997_119#_c_831_n 0.00432339f $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_329 N_A_217_463#_c_253_n N_A_997_119#_c_832_n 0.0076208f $X=5.385 $Y=1.48
+ $X2=0 $Y2=0
cc_330 N_A_217_463#_c_253_n N_A_997_119#_c_833_n 0.0197912f $X=5.385 $Y=1.48
+ $X2=0 $Y2=0
cc_331 N_A_217_463#_M1019_g N_A_997_119#_c_833_n 0.0139969f $X=5.61 $Y=2.105
+ $X2=0 $Y2=0
cc_332 N_A_217_463#_c_255_n N_A_997_119#_c_833_n 0.0192616f $X=4.95 $Y=2.415
+ $X2=0 $Y2=0
cc_333 N_A_217_463#_c_256_n N_A_997_119#_c_833_n 0.0186468f $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_334 N_A_217_463#_c_257_n N_A_997_119#_c_833_n 0.00268696f $X=5 $Y=1.39 $X2=0
+ $Y2=0
cc_335 N_A_217_463#_c_265_n N_VPWR_M1002_d 0.0103486f $X=1.905 $Y=2.4 $X2=0
+ $Y2=0
cc_336 N_A_217_463#_c_266_n N_VPWR_M1002_d 0.00320389f $X=1.99 $Y=2.865 $X2=0
+ $Y2=0
cc_337 N_A_217_463#_c_270_n N_VPWR_M1001_d 0.0113511f $X=4.865 $Y=2.5 $X2=0
+ $Y2=0
cc_338 N_A_217_463#_c_265_n N_VPWR_c_969_n 0.014347f $X=1.905 $Y=2.4 $X2=0 $Y2=0
cc_339 N_A_217_463#_c_266_n N_VPWR_c_969_n 0.0157928f $X=1.99 $Y=2.865 $X2=0
+ $Y2=0
cc_340 N_A_217_463#_c_268_n N_VPWR_c_969_n 0.0180344f $X=2.075 $Y=2.97 $X2=0
+ $Y2=0
cc_341 N_A_217_463#_c_272_n N_VPWR_c_969_n 0.0114431f $X=1.21 $Y=2.46 $X2=0
+ $Y2=0
cc_342 N_A_217_463#_c_267_n N_VPWR_c_970_n 0.00637086f $X=3.13 $Y=2.97 $X2=0
+ $Y2=0
cc_343 N_A_217_463#_c_270_n N_VPWR_c_970_n 0.0240132f $X=4.865 $Y=2.5 $X2=0
+ $Y2=0
cc_344 N_A_217_463#_c_270_n N_VPWR_c_975_n 0.0095277f $X=4.865 $Y=2.5 $X2=0
+ $Y2=0
cc_345 N_A_217_463#_c_272_n N_VPWR_c_977_n 0.0116922f $X=1.21 $Y=2.46 $X2=0
+ $Y2=0
cc_346 N_A_217_463#_c_267_n N_VPWR_c_978_n 0.0803534f $X=3.13 $Y=2.97 $X2=0
+ $Y2=0
cc_347 N_A_217_463#_c_268_n N_VPWR_c_978_n 0.0115893f $X=2.075 $Y=2.97 $X2=0
+ $Y2=0
cc_348 N_A_217_463#_c_270_n N_VPWR_c_978_n 0.00799375f $X=4.865 $Y=2.5 $X2=0
+ $Y2=0
cc_349 N_A_217_463#_M1019_g N_VPWR_c_966_n 0.00373935f $X=5.61 $Y=2.105 $X2=0
+ $Y2=0
cc_350 N_A_217_463#_c_265_n N_VPWR_c_966_n 0.00803593f $X=1.905 $Y=2.4 $X2=0
+ $Y2=0
cc_351 N_A_217_463#_c_267_n N_VPWR_c_966_n 0.0413849f $X=3.13 $Y=2.97 $X2=0
+ $Y2=0
cc_352 N_A_217_463#_c_268_n N_VPWR_c_966_n 0.00583135f $X=2.075 $Y=2.97 $X2=0
+ $Y2=0
cc_353 N_A_217_463#_c_270_n N_VPWR_c_966_n 0.032634f $X=4.865 $Y=2.5 $X2=0 $Y2=0
cc_354 N_A_217_463#_c_272_n N_VPWR_c_966_n 0.0133089f $X=1.21 $Y=2.46 $X2=0
+ $Y2=0
cc_355 N_A_217_463#_M1014_g N_A_440_463#_c_1064_n 0.00189017f $X=3.2 $Y=0.805
+ $X2=0 $Y2=0
cc_356 N_A_217_463#_c_262_n N_A_440_463#_c_1064_n 0.00422119f $X=2.63 $Y=1.99
+ $X2=0 $Y2=0
cc_357 N_A_217_463#_c_267_n N_A_440_463#_c_1064_n 0.0140252f $X=3.13 $Y=2.97
+ $X2=0 $Y2=0
cc_358 N_A_217_463#_c_270_n A_650_499# 0.00971595f $X=4.865 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_359 N_A_217_463#_M1014_g N_VGND_c_1111_n 0.0015955f $X=3.2 $Y=0.805 $X2=0
+ $Y2=0
cc_360 N_A_217_463#_M1018_g N_VGND_c_1111_n 6.26645e-19 $X=4.91 $Y=0.805 $X2=0
+ $Y2=0
cc_361 N_A_217_463#_c_254_n N_VGND_c_1115_n 0.0038632f $X=1.325 $Y=0.805 $X2=0
+ $Y2=0
cc_362 N_A_217_463#_M1014_g N_VGND_c_1123_n 9.39239e-19 $X=3.2 $Y=0.805 $X2=0
+ $Y2=0
cc_363 N_A_217_463#_M1018_g N_VGND_c_1123_n 9.39239e-19 $X=4.91 $Y=0.805 $X2=0
+ $Y2=0
cc_364 N_A_217_463#_c_254_n N_VGND_c_1123_n 0.00628885f $X=1.325 $Y=0.805 $X2=0
+ $Y2=0
cc_365 N_A_697_93#_c_418_n N_A_526_463#_M1024_g 0.00414465f $X=3.56 $Y=1.125
+ $X2=0 $Y2=0
cc_366 N_A_697_93#_c_419_n N_A_526_463#_M1024_g 0.0130693f $X=4.505 $Y=1.17
+ $X2=0 $Y2=0
cc_367 N_A_697_93#_c_421_n N_A_526_463#_M1024_g 8.50044e-19 $X=3.71 $Y=1.17
+ $X2=0 $Y2=0
cc_368 N_A_697_93#_c_423_n N_A_526_463#_M1024_g 0.00790135f $X=3.75 $Y=1.29
+ $X2=0 $Y2=0
cc_369 N_A_697_93#_M1001_g N_A_526_463#_M1013_g 0.0151736f $X=3.685 $Y=2.525
+ $X2=0 $Y2=0
cc_370 N_A_697_93#_c_426_n N_A_526_463#_M1013_g 0.0149426f $X=4.6 $Y=2.07 $X2=0
+ $Y2=0
cc_371 N_A_697_93#_c_422_n N_A_526_463#_M1013_g 0.01034f $X=3.66 $Y=1.825 $X2=0
+ $Y2=0
cc_372 N_A_697_93#_c_418_n N_A_526_463#_c_489_n 0.00295618f $X=3.56 $Y=1.125
+ $X2=0 $Y2=0
cc_373 N_A_697_93#_c_421_n N_A_526_463#_c_489_n 0.0115428f $X=3.71 $Y=1.17 $X2=0
+ $Y2=0
cc_374 N_A_697_93#_c_422_n N_A_526_463#_c_489_n 4.67066e-19 $X=3.66 $Y=1.825
+ $X2=0 $Y2=0
cc_375 N_A_697_93#_c_419_n N_A_526_463#_c_491_n 0.0240603f $X=4.505 $Y=1.17
+ $X2=0 $Y2=0
cc_376 N_A_697_93#_c_422_n N_A_526_463#_c_491_n 6.13233e-19 $X=3.66 $Y=1.825
+ $X2=0 $Y2=0
cc_377 N_A_697_93#_c_423_n N_A_526_463#_c_491_n 2.04346e-19 $X=3.75 $Y=1.29
+ $X2=0 $Y2=0
cc_378 N_A_697_93#_c_426_n N_A_526_463#_c_492_n 0.00400328f $X=4.6 $Y=2.07 $X2=0
+ $Y2=0
cc_379 N_A_697_93#_c_419_n N_A_526_463#_c_492_n 0.00413151f $X=4.505 $Y=1.17
+ $X2=0 $Y2=0
cc_380 N_A_697_93#_c_422_n N_A_526_463#_c_492_n 0.0111255f $X=3.66 $Y=1.825
+ $X2=0 $Y2=0
cc_381 N_A_697_93#_c_423_n N_A_526_463#_c_492_n 0.00277893f $X=3.75 $Y=1.29
+ $X2=0 $Y2=0
cc_382 N_A_697_93#_c_425_n N_A_526_463#_c_493_n 0.0015833f $X=3.66 $Y=1.99 $X2=0
+ $Y2=0
cc_383 N_A_697_93#_c_426_n N_A_526_463#_c_493_n 0.0710483f $X=4.6 $Y=2.07 $X2=0
+ $Y2=0
cc_384 N_A_697_93#_c_419_n N_A_526_463#_c_493_n 0.0129261f $X=4.505 $Y=1.17
+ $X2=0 $Y2=0
cc_385 N_A_697_93#_c_421_n N_A_526_463#_c_493_n 0.0240324f $X=3.71 $Y=1.17 $X2=0
+ $Y2=0
cc_386 N_A_697_93#_c_422_n N_A_526_463#_c_493_n 0.0111472f $X=3.66 $Y=1.825
+ $X2=0 $Y2=0
cc_387 N_A_697_93#_c_423_n N_A_526_463#_c_493_n 0.00416253f $X=3.75 $Y=1.29
+ $X2=0 $Y2=0
cc_388 N_A_697_93#_c_418_n N_A_110_82#_c_577_n 0.0103107f $X=3.56 $Y=1.125 $X2=0
+ $Y2=0
cc_389 N_A_697_93#_c_420_n N_A_110_82#_c_577_n 0.00377174f $X=4.6 $Y=0.75 $X2=0
+ $Y2=0
cc_390 N_A_697_93#_M1001_g N_A_110_82#_M1016_g 0.015285f $X=3.685 $Y=2.525 $X2=0
+ $Y2=0
cc_391 N_A_697_93#_M1001_g N_A_110_82#_c_589_n 0.00993882f $X=3.685 $Y=2.525
+ $X2=0 $Y2=0
cc_392 N_A_697_93#_c_426_n N_A_110_82#_M1025_g 0.00113649f $X=4.6 $Y=2.07 $X2=0
+ $Y2=0
cc_393 N_A_697_93#_c_419_n N_A_997_119#_c_831_n 0.00517836f $X=4.505 $Y=1.17
+ $X2=0 $Y2=0
cc_394 N_A_697_93#_c_420_n N_A_997_119#_c_831_n 0.00275687f $X=4.6 $Y=0.75 $X2=0
+ $Y2=0
cc_395 N_A_697_93#_c_426_n N_VPWR_M1001_d 0.00789805f $X=4.6 $Y=2.07 $X2=0 $Y2=0
cc_396 N_A_697_93#_M1001_g N_VPWR_c_970_n 0.00136086f $X=3.685 $Y=2.525 $X2=0
+ $Y2=0
cc_397 N_A_697_93#_M1001_g N_VPWR_c_966_n 9.39239e-19 $X=3.685 $Y=2.525 $X2=0
+ $Y2=0
cc_398 N_A_697_93#_c_419_n N_VGND_M1005_d 0.00283787f $X=4.505 $Y=1.17 $X2=0
+ $Y2=0
cc_399 N_A_697_93#_c_418_n N_VGND_c_1111_n 0.0107665f $X=3.56 $Y=1.125 $X2=0
+ $Y2=0
cc_400 N_A_697_93#_c_419_n N_VGND_c_1111_n 0.0327659f $X=4.505 $Y=1.17 $X2=0
+ $Y2=0
cc_401 N_A_697_93#_c_420_n N_VGND_c_1111_n 0.0141797f $X=4.6 $Y=0.75 $X2=0 $Y2=0
cc_402 N_A_697_93#_c_421_n N_VGND_c_1111_n 0.0199755f $X=3.71 $Y=1.17 $X2=0
+ $Y2=0
cc_403 N_A_697_93#_c_423_n N_VGND_c_1111_n 0.00152496f $X=3.75 $Y=1.29 $X2=0
+ $Y2=0
cc_404 N_A_697_93#_c_420_n N_VGND_c_1117_n 0.00422723f $X=4.6 $Y=0.75 $X2=0
+ $Y2=0
cc_405 N_A_697_93#_c_418_n N_VGND_c_1123_n 7.88961e-19 $X=3.56 $Y=1.125 $X2=0
+ $Y2=0
cc_406 N_A_697_93#_c_420_n N_VGND_c_1123_n 0.0051697f $X=4.6 $Y=0.75 $X2=0 $Y2=0
cc_407 N_A_526_463#_c_489_n N_A_110_82#_M1010_g 0.00166186f $X=2.985 $Y=0.8
+ $X2=0 $Y2=0
cc_408 N_A_526_463#_c_490_n N_A_110_82#_M1010_g 0.00300657f $X=3.16 $Y=1.64
+ $X2=0 $Y2=0
cc_409 N_A_526_463#_M1024_g N_A_110_82#_c_577_n 0.0103107f $X=4.385 $Y=0.915
+ $X2=0 $Y2=0
cc_410 N_A_526_463#_c_489_n N_A_110_82#_c_577_n 0.00343726f $X=2.985 $Y=0.8
+ $X2=0 $Y2=0
cc_411 N_A_526_463#_c_517_n N_A_110_82#_M1016_g 0.0027175f $X=2.865 $Y=2.53
+ $X2=0 $Y2=0
cc_412 N_A_526_463#_M1013_g N_A_110_82#_c_589_n 0.00993882f $X=4.385 $Y=2.315
+ $X2=0 $Y2=0
cc_413 N_A_526_463#_M1013_g N_A_110_82#_M1025_g 0.0177833f $X=4.385 $Y=2.315
+ $X2=0 $Y2=0
cc_414 N_A_526_463#_M1013_g N_VPWR_c_970_n 0.00310929f $X=4.385 $Y=2.315 $X2=0
+ $Y2=0
cc_415 N_A_526_463#_M1013_g N_VPWR_c_966_n 9.39239e-19 $X=4.385 $Y=2.315 $X2=0
+ $Y2=0
cc_416 N_A_526_463#_c_495_n N_A_440_463#_c_1064_n 0.0445726f $X=2.69 $Y=2.365
+ $X2=0 $Y2=0
cc_417 N_A_526_463#_c_489_n N_A_440_463#_c_1064_n 0.0224603f $X=2.985 $Y=0.8
+ $X2=0 $Y2=0
cc_418 N_A_526_463#_c_490_n N_A_440_463#_c_1064_n 0.0142973f $X=3.16 $Y=1.64
+ $X2=0 $Y2=0
cc_419 N_A_526_463#_c_490_n N_A_440_463#_c_1070_n 0.00194998f $X=3.16 $Y=1.64
+ $X2=0 $Y2=0
cc_420 N_A_526_463#_M1024_g N_VGND_c_1111_n 0.00912344f $X=4.385 $Y=0.915 $X2=0
+ $Y2=0
cc_421 N_A_526_463#_c_489_n N_VGND_c_1111_n 0.0100248f $X=2.985 $Y=0.8 $X2=0
+ $Y2=0
cc_422 N_A_526_463#_c_489_n N_VGND_c_1119_n 0.00471174f $X=2.985 $Y=0.8 $X2=0
+ $Y2=0
cc_423 N_A_526_463#_M1024_g N_VGND_c_1123_n 7.88961e-19 $X=4.385 $Y=0.915 $X2=0
+ $Y2=0
cc_424 N_A_526_463#_c_489_n N_VGND_c_1123_n 0.00768442f $X=2.985 $Y=0.8 $X2=0
+ $Y2=0
cc_425 N_A_110_82#_M1000_g N_A_1149_93#_c_708_n 0.0389023f $X=5.45 $Y=0.805
+ $X2=0 $Y2=0
cc_426 N_A_110_82#_M1025_g N_A_997_119#_c_838_n 0.00162397f $X=5.085 $Y=2.315
+ $X2=0 $Y2=0
cc_427 N_A_110_82#_c_577_n N_A_997_119#_c_831_n 0.00492963f $X=5.375 $Y=0.18
+ $X2=0 $Y2=0
cc_428 N_A_110_82#_M1000_g N_A_997_119#_c_831_n 0.0201767f $X=5.45 $Y=0.805
+ $X2=0 $Y2=0
cc_429 N_A_110_82#_M1000_g N_A_997_119#_c_832_n 0.00330148f $X=5.45 $Y=0.805
+ $X2=0 $Y2=0
cc_430 N_A_110_82#_M1025_g N_A_997_119#_c_833_n 9.11673e-19 $X=5.085 $Y=2.315
+ $X2=0 $Y2=0
cc_431 N_A_110_82#_c_592_n N_VPWR_c_968_n 0.00225185f $X=0.677 $Y=2.437 $X2=0
+ $Y2=0
cc_432 N_A_110_82#_M1002_g N_VPWR_c_969_n 0.00951081f $X=1.425 $Y=2.635 $X2=0
+ $Y2=0
cc_433 N_A_110_82#_c_586_n N_VPWR_c_969_n 0.0144762f $X=3.1 $Y=3.15 $X2=0 $Y2=0
cc_434 N_A_110_82#_c_587_n N_VPWR_c_969_n 0.00320181f $X=1.5 $Y=3.15 $X2=0 $Y2=0
cc_435 N_A_110_82#_M1016_g N_VPWR_c_970_n 0.00109031f $X=3.175 $Y=2.705 $X2=0
+ $Y2=0
cc_436 N_A_110_82#_c_589_n N_VPWR_c_970_n 0.0249093f $X=5.01 $Y=3.15 $X2=0 $Y2=0
cc_437 N_A_110_82#_c_589_n N_VPWR_c_975_n 0.0247645f $X=5.01 $Y=3.15 $X2=0 $Y2=0
cc_438 N_A_110_82#_c_587_n N_VPWR_c_977_n 0.00564095f $X=1.5 $Y=3.15 $X2=0 $Y2=0
cc_439 N_A_110_82#_c_593_n N_VPWR_c_977_n 0.0108291f $X=0.69 $Y=2.485 $X2=0
+ $Y2=0
cc_440 N_A_110_82#_c_586_n N_VPWR_c_978_n 0.0517808f $X=3.1 $Y=3.15 $X2=0 $Y2=0
cc_441 N_A_110_82#_c_586_n N_VPWR_c_966_n 0.0327287f $X=3.1 $Y=3.15 $X2=0 $Y2=0
cc_442 N_A_110_82#_c_587_n N_VPWR_c_966_n 0.00675293f $X=1.5 $Y=3.15 $X2=0 $Y2=0
cc_443 N_A_110_82#_c_589_n N_VPWR_c_966_n 0.0507302f $X=5.01 $Y=3.15 $X2=0 $Y2=0
cc_444 N_A_110_82#_c_591_n N_VPWR_c_966_n 0.00370837f $X=3.175 $Y=3.15 $X2=0
+ $Y2=0
cc_445 N_A_110_82#_c_593_n N_VPWR_c_966_n 0.00865621f $X=0.69 $Y=2.485 $X2=0
+ $Y2=0
cc_446 N_A_110_82#_M1008_g N_A_440_463#_c_1064_n 0.00293117f $X=1.54 $Y=0.805
+ $X2=0 $Y2=0
cc_447 N_A_110_82#_M1010_g N_A_440_463#_c_1064_n 9.80664e-19 $X=2.77 $Y=0.805
+ $X2=0 $Y2=0
cc_448 N_A_110_82#_c_574_n N_A_440_463#_c_1070_n 0.00360811f $X=2.695 $Y=0.18
+ $X2=0 $Y2=0
cc_449 N_A_110_82#_M1008_g N_VGND_c_1110_n 0.0169281f $X=1.54 $Y=0.805 $X2=0
+ $Y2=0
cc_450 N_A_110_82#_c_574_n N_VGND_c_1110_n 0.0252002f $X=2.695 $Y=0.18 $X2=0
+ $Y2=0
cc_451 N_A_110_82#_M1010_g N_VGND_c_1110_n 0.00506879f $X=2.77 $Y=0.805 $X2=0
+ $Y2=0
cc_452 N_A_110_82#_c_577_n N_VGND_c_1111_n 0.0474375f $X=5.375 $Y=0.18 $X2=0
+ $Y2=0
cc_453 N_A_110_82#_c_577_n N_VGND_c_1112_n 0.00868846f $X=5.375 $Y=0.18 $X2=0
+ $Y2=0
cc_454 N_A_110_82#_c_575_n N_VGND_c_1115_n 0.0110921f $X=1.615 $Y=0.18 $X2=0
+ $Y2=0
cc_455 N_A_110_82#_c_581_n N_VGND_c_1115_n 0.00841253f $X=0.71 $Y=0.615 $X2=0
+ $Y2=0
cc_456 N_A_110_82#_c_577_n N_VGND_c_1117_n 0.0362304f $X=5.375 $Y=0.18 $X2=0
+ $Y2=0
cc_457 N_A_110_82#_c_574_n N_VGND_c_1119_n 0.0473928f $X=2.695 $Y=0.18 $X2=0
+ $Y2=0
cc_458 N_A_110_82#_c_574_n N_VGND_c_1123_n 0.0292076f $X=2.695 $Y=0.18 $X2=0
+ $Y2=0
cc_459 N_A_110_82#_c_575_n N_VGND_c_1123_n 0.0116041f $X=1.615 $Y=0.18 $X2=0
+ $Y2=0
cc_460 N_A_110_82#_c_577_n N_VGND_c_1123_n 0.0730427f $X=5.375 $Y=0.18 $X2=0
+ $Y2=0
cc_461 N_A_110_82#_c_580_n N_VGND_c_1123_n 0.00926736f $X=2.77 $Y=0.18 $X2=0
+ $Y2=0
cc_462 N_A_110_82#_c_581_n N_VGND_c_1123_n 0.00962766f $X=0.71 $Y=0.615 $X2=0
+ $Y2=0
cc_463 N_A_1149_93#_M1003_g N_A_997_119#_M1020_g 0.0124736f $X=5.97 $Y=2.105
+ $X2=0 $Y2=0
cc_464 N_A_1149_93#_c_712_n N_A_997_119#_M1020_g 0.00462776f $X=7.545 $Y=1.485
+ $X2=0 $Y2=0
cc_465 N_A_1149_93#_c_714_n N_A_997_119#_M1020_g 0.012308f $X=6.58 $Y=1.72 $X2=0
+ $Y2=0
cc_466 N_A_1149_93#_c_724_n N_A_997_119#_M1020_g 0.0118055f $X=6.725 $Y=2.04
+ $X2=0 $Y2=0
cc_467 N_A_1149_93#_c_726_n N_A_997_119#_M1020_g 0.00445369f $X=7.035 $Y=2.46
+ $X2=0 $Y2=0
cc_468 N_A_1149_93#_c_728_n N_A_997_119#_M1020_g 7.52794e-19 $X=6.06 $Y=1.57
+ $X2=0 $Y2=0
cc_469 N_A_1149_93#_c_717_n N_A_997_119#_M1020_g 0.00609966f $X=6.95 $Y=1.562
+ $X2=0 $Y2=0
cc_470 N_A_1149_93#_c_708_n N_A_997_119#_c_831_n 0.00192874f $X=5.82 $Y=1.125
+ $X2=0 $Y2=0
cc_471 N_A_1149_93#_c_709_n N_A_997_119#_c_832_n 0.0312805f $X=5.97 $Y=1.735
+ $X2=0 $Y2=0
cc_472 N_A_1149_93#_c_714_n N_A_997_119#_c_832_n 0.00979f $X=6.58 $Y=1.72 $X2=0
+ $Y2=0
cc_473 N_A_1149_93#_c_728_n N_A_997_119#_c_832_n 0.0220391f $X=6.06 $Y=1.57
+ $X2=0 $Y2=0
cc_474 N_A_1149_93#_c_709_n N_A_997_119#_c_833_n 0.00391165f $X=5.97 $Y=1.735
+ $X2=0 $Y2=0
cc_475 N_A_1149_93#_c_728_n N_A_997_119#_c_833_n 0.0114306f $X=6.06 $Y=1.57
+ $X2=0 $Y2=0
cc_476 N_A_1149_93#_c_709_n N_A_997_119#_c_834_n 0.00113672f $X=5.97 $Y=1.735
+ $X2=0 $Y2=0
cc_477 N_A_1149_93#_c_714_n N_A_997_119#_c_834_n 0.00983891f $X=6.58 $Y=1.72
+ $X2=0 $Y2=0
cc_478 N_A_1149_93#_c_715_n N_A_997_119#_c_834_n 0.00835112f $X=6.95 $Y=0.955
+ $X2=0 $Y2=0
cc_479 N_A_1149_93#_c_716_n N_A_997_119#_c_834_n 0.0137088f $X=6.95 $Y=1.32
+ $X2=0 $Y2=0
cc_480 N_A_1149_93#_c_717_n N_A_997_119#_c_834_n 0.0186552f $X=6.95 $Y=1.562
+ $X2=0 $Y2=0
cc_481 N_A_1149_93#_c_709_n N_A_997_119#_c_835_n 0.0307515f $X=5.97 $Y=1.735
+ $X2=0 $Y2=0
cc_482 N_A_1149_93#_c_712_n N_A_997_119#_c_835_n 0.00706937f $X=7.545 $Y=1.485
+ $X2=0 $Y2=0
cc_483 N_A_1149_93#_c_715_n N_A_997_119#_c_835_n 0.00302498f $X=6.95 $Y=0.955
+ $X2=0 $Y2=0
cc_484 N_A_1149_93#_c_716_n N_A_997_119#_c_835_n 0.00477293f $X=6.95 $Y=1.32
+ $X2=0 $Y2=0
cc_485 N_A_1149_93#_c_717_n N_A_997_119#_c_835_n 0.00417658f $X=6.95 $Y=1.562
+ $X2=0 $Y2=0
cc_486 N_A_1149_93#_c_708_n N_A_997_119#_c_836_n 0.011022f $X=5.82 $Y=1.125
+ $X2=0 $Y2=0
cc_487 N_A_1149_93#_c_715_n N_A_997_119#_c_836_n 0.00775648f $X=6.95 $Y=0.955
+ $X2=0 $Y2=0
cc_488 N_A_1149_93#_c_716_n N_A_997_119#_c_836_n 0.00424213f $X=6.95 $Y=1.32
+ $X2=0 $Y2=0
cc_489 N_A_1149_93#_c_725_n N_A_1401_22#_M1021_s 0.00268224f $X=8.72 $Y=2.46
+ $X2=0 $Y2=0
cc_490 N_A_1149_93#_c_710_n N_A_1401_22#_c_902_n 0.00506278f $X=7.62 $Y=1.32
+ $X2=0 $Y2=0
cc_491 N_A_1149_93#_c_710_n N_A_1401_22#_M1012_g 0.0159816f $X=7.62 $Y=1.32
+ $X2=0 $Y2=0
cc_492 N_A_1149_93#_c_713_n N_A_1401_22#_M1012_g 0.0350538f $X=7.545 $Y=1.32
+ $X2=0 $Y2=0
cc_493 N_A_1149_93#_c_725_n N_A_1401_22#_M1012_g 0.0187298f $X=8.72 $Y=2.46
+ $X2=0 $Y2=0
cc_494 N_A_1149_93#_c_727_n N_A_1401_22#_M1012_g 0.00495598f $X=8.885 $Y=1.51
+ $X2=0 $Y2=0
cc_495 N_A_1149_93#_c_718_n N_A_1401_22#_M1012_g 0.00568244f $X=9.125 $Y=1.51
+ $X2=0 $Y2=0
cc_496 N_A_1149_93#_c_710_n N_A_1401_22#_c_905_n 0.0030177f $X=7.62 $Y=1.32
+ $X2=0 $Y2=0
cc_497 N_A_1149_93#_c_715_n N_A_1401_22#_c_905_n 0.0134963f $X=6.95 $Y=0.955
+ $X2=0 $Y2=0
cc_498 N_A_1149_93#_c_710_n N_A_1401_22#_c_906_n 0.00787005f $X=7.62 $Y=1.32
+ $X2=0 $Y2=0
cc_499 N_A_1149_93#_M1021_g N_A_1401_22#_c_906_n 0.00801751f $X=7.64 $Y=2.155
+ $X2=0 $Y2=0
cc_500 N_A_1149_93#_c_712_n N_A_1401_22#_c_906_n 0.0119896f $X=7.545 $Y=1.485
+ $X2=0 $Y2=0
cc_501 N_A_1149_93#_c_713_n N_A_1401_22#_c_906_n 0.0078262f $X=7.545 $Y=1.32
+ $X2=0 $Y2=0
cc_502 N_A_1149_93#_c_724_n N_A_1401_22#_c_906_n 0.00306869f $X=6.725 $Y=2.04
+ $X2=0 $Y2=0
cc_503 N_A_1149_93#_c_716_n N_A_1401_22#_c_906_n 0.0113965f $X=6.95 $Y=1.32
+ $X2=0 $Y2=0
cc_504 N_A_1149_93#_c_717_n N_A_1401_22#_c_906_n 0.0313387f $X=6.95 $Y=1.562
+ $X2=0 $Y2=0
cc_505 N_A_1149_93#_c_715_n N_A_1401_22#_c_907_n 0.00359931f $X=6.95 $Y=0.955
+ $X2=0 $Y2=0
cc_506 N_A_1149_93#_c_715_n N_A_1401_22#_c_908_n 0.0191239f $X=6.95 $Y=0.955
+ $X2=0 $Y2=0
cc_507 N_A_1149_93#_c_710_n N_A_1401_22#_c_909_n 0.00338979f $X=7.62 $Y=1.32
+ $X2=0 $Y2=0
cc_508 N_A_1149_93#_c_712_n N_A_1401_22#_c_909_n 0.00655111f $X=7.545 $Y=1.485
+ $X2=0 $Y2=0
cc_509 N_A_1149_93#_c_715_n N_A_1401_22#_c_909_n 0.0104305f $X=6.95 $Y=0.955
+ $X2=0 $Y2=0
cc_510 N_A_1149_93#_c_716_n N_A_1401_22#_c_909_n 0.0064747f $X=6.95 $Y=1.32
+ $X2=0 $Y2=0
cc_511 N_A_1149_93#_c_717_n N_A_1401_22#_c_909_n 0.00264095f $X=6.95 $Y=1.562
+ $X2=0 $Y2=0
cc_512 N_A_1149_93#_M1021_g N_A_1401_22#_c_912_n 0.007507f $X=7.64 $Y=2.155
+ $X2=0 $Y2=0
cc_513 N_A_1149_93#_c_712_n N_A_1401_22#_c_912_n 0.00707609f $X=7.545 $Y=1.485
+ $X2=0 $Y2=0
cc_514 N_A_1149_93#_c_724_n N_A_1401_22#_c_912_n 0.0231678f $X=6.725 $Y=2.04
+ $X2=0 $Y2=0
cc_515 N_A_1149_93#_c_725_n N_A_1401_22#_c_912_n 0.0218486f $X=8.72 $Y=2.46
+ $X2=0 $Y2=0
cc_516 N_A_1149_93#_c_717_n N_A_1401_22#_c_912_n 3.22185e-19 $X=6.95 $Y=1.562
+ $X2=0 $Y2=0
cc_517 N_A_1149_93#_c_725_n N_VPWR_M1021_d 0.0122689f $X=8.72 $Y=2.46 $X2=0
+ $Y2=0
cc_518 N_A_1149_93#_c_725_n N_VPWR_M1017_s 0.00479303f $X=8.72 $Y=2.46 $X2=0
+ $Y2=0
cc_519 N_A_1149_93#_c_727_n N_VPWR_M1017_s 0.00597518f $X=8.885 $Y=1.51 $X2=0
+ $Y2=0
cc_520 N_A_1149_93#_c_709_n N_VPWR_c_971_n 8.87367e-19 $X=5.97 $Y=1.735 $X2=0
+ $Y2=0
cc_521 N_A_1149_93#_M1003_g N_VPWR_c_971_n 0.00403263f $X=5.97 $Y=2.105 $X2=0
+ $Y2=0
cc_522 N_A_1149_93#_c_714_n N_VPWR_c_971_n 0.0138236f $X=6.58 $Y=1.72 $X2=0
+ $Y2=0
cc_523 N_A_1149_93#_c_726_n N_VPWR_c_971_n 0.0157453f $X=7.035 $Y=2.46 $X2=0
+ $Y2=0
cc_524 N_A_1149_93#_c_728_n N_VPWR_c_971_n 0.0114813f $X=6.06 $Y=1.57 $X2=0
+ $Y2=0
cc_525 N_A_1149_93#_c_725_n N_VPWR_c_972_n 0.0214609f $X=8.72 $Y=2.46 $X2=0
+ $Y2=0
cc_526 N_A_1149_93#_M1017_g N_VPWR_c_974_n 0.00460896f $X=9.125 $Y=2.465 $X2=0
+ $Y2=0
cc_527 N_A_1149_93#_c_725_n N_VPWR_c_974_n 0.012083f $X=8.72 $Y=2.46 $X2=0 $Y2=0
cc_528 N_A_1149_93#_M1021_g N_VPWR_c_979_n 0.00312414f $X=7.64 $Y=2.155 $X2=0
+ $Y2=0
cc_529 N_A_1149_93#_c_726_n N_VPWR_c_979_n 0.00679071f $X=7.035 $Y=2.46 $X2=0
+ $Y2=0
cc_530 N_A_1149_93#_M1017_g N_VPWR_c_980_n 0.00585385f $X=9.125 $Y=2.465 $X2=0
+ $Y2=0
cc_531 N_A_1149_93#_M1003_g N_VPWR_c_966_n 0.00373935f $X=5.97 $Y=2.105 $X2=0
+ $Y2=0
cc_532 N_A_1149_93#_M1021_g N_VPWR_c_966_n 0.00410284f $X=7.64 $Y=2.155 $X2=0
+ $Y2=0
cc_533 N_A_1149_93#_M1017_g N_VPWR_c_966_n 0.012823f $X=9.125 $Y=2.465 $X2=0
+ $Y2=0
cc_534 N_A_1149_93#_c_725_n N_VPWR_c_966_n 0.0548512f $X=8.72 $Y=2.46 $X2=0
+ $Y2=0
cc_535 N_A_1149_93#_c_726_n N_VPWR_c_966_n 0.0159712f $X=7.035 $Y=2.46 $X2=0
+ $Y2=0
cc_536 N_A_1149_93#_c_725_n N_Q_N_M1007_d 0.00698496f $X=8.72 $Y=2.46 $X2=0
+ $Y2=0
cc_537 N_A_1149_93#_c_711_n N_Q_N_c_1084_n 0.00370208f $X=9.125 $Y=1.345 $X2=0
+ $Y2=0
cc_538 N_A_1149_93#_c_725_n N_Q_N_c_1084_n 0.0202165f $X=8.72 $Y=2.46 $X2=0
+ $Y2=0
cc_539 N_A_1149_93#_c_727_n N_Q_N_c_1084_n 0.0619811f $X=8.885 $Y=1.51 $X2=0
+ $Y2=0
cc_540 N_A_1149_93#_c_718_n N_Q_N_c_1084_n 0.00445558f $X=9.125 $Y=1.51 $X2=0
+ $Y2=0
cc_541 N_A_1149_93#_c_711_n Q 0.0255155f $X=9.125 $Y=1.345 $X2=0 $Y2=0
cc_542 N_A_1149_93#_c_727_n Q 0.0305485f $X=8.885 $Y=1.51 $X2=0 $Y2=0
cc_543 N_A_1149_93#_c_708_n N_VGND_c_1112_n 0.00905078f $X=5.82 $Y=1.125 $X2=0
+ $Y2=0
cc_544 N_A_1149_93#_c_709_n N_VGND_c_1112_n 6.32207e-19 $X=5.97 $Y=1.735 $X2=0
+ $Y2=0
cc_545 N_A_1149_93#_c_715_n N_VGND_c_1112_n 0.0239171f $X=6.95 $Y=0.955 $X2=0
+ $Y2=0
cc_546 N_A_1149_93#_c_710_n N_VGND_c_1113_n 0.00538249f $X=7.62 $Y=1.32 $X2=0
+ $Y2=0
cc_547 N_A_1149_93#_c_711_n N_VGND_c_1114_n 0.00868411f $X=9.125 $Y=1.345 $X2=0
+ $Y2=0
cc_548 N_A_1149_93#_c_727_n N_VGND_c_1114_n 0.0238909f $X=8.885 $Y=1.51 $X2=0
+ $Y2=0
cc_549 N_A_1149_93#_c_718_n N_VGND_c_1114_n 0.00687592f $X=9.125 $Y=1.51 $X2=0
+ $Y2=0
cc_550 N_A_1149_93#_c_708_n N_VGND_c_1117_n 0.00431487f $X=5.82 $Y=1.125 $X2=0
+ $Y2=0
cc_551 N_A_1149_93#_c_715_n N_VGND_c_1120_n 0.0146459f $X=6.95 $Y=0.955 $X2=0
+ $Y2=0
cc_552 N_A_1149_93#_c_711_n N_VGND_c_1122_n 0.00559701f $X=9.125 $Y=1.345 $X2=0
+ $Y2=0
cc_553 N_A_1149_93#_c_708_n N_VGND_c_1123_n 0.00477801f $X=5.82 $Y=1.125 $X2=0
+ $Y2=0
cc_554 N_A_1149_93#_c_710_n N_VGND_c_1123_n 9.67605e-19 $X=7.62 $Y=1.32 $X2=0
+ $Y2=0
cc_555 N_A_1149_93#_c_711_n N_VGND_c_1123_n 0.00537853f $X=9.125 $Y=1.345 $X2=0
+ $Y2=0
cc_556 N_A_1149_93#_c_715_n N_VGND_c_1123_n 0.0182417f $X=6.95 $Y=0.955 $X2=0
+ $Y2=0
cc_557 N_A_997_119#_c_836_n N_A_1401_22#_c_903_n 0.00594057f $X=6.6 $Y=1.125
+ $X2=0 $Y2=0
cc_558 N_A_997_119#_c_836_n N_A_1401_22#_c_908_n 5.24915e-19 $X=6.6 $Y=1.125
+ $X2=0 $Y2=0
cc_559 N_A_997_119#_M1020_g N_A_1401_22#_c_912_n 4.81011e-19 $X=6.51 $Y=2.315
+ $X2=0 $Y2=0
cc_560 N_A_997_119#_M1020_g N_VPWR_c_971_n 0.00604583f $X=6.51 $Y=2.315 $X2=0
+ $Y2=0
cc_561 N_A_997_119#_c_838_n N_VPWR_c_971_n 0.0194124f $X=5.335 $Y=2.005 $X2=0
+ $Y2=0
cc_562 N_A_997_119#_c_839_n N_VPWR_c_975_n 0.00588273f $X=5.3 $Y=2.04 $X2=0
+ $Y2=0
cc_563 N_A_997_119#_M1020_g N_VPWR_c_979_n 0.00428067f $X=6.51 $Y=2.315 $X2=0
+ $Y2=0
cc_564 N_A_997_119#_M1020_g N_VPWR_c_966_n 0.00477801f $X=6.51 $Y=2.315 $X2=0
+ $Y2=0
cc_565 N_A_997_119#_c_839_n N_VPWR_c_966_n 0.0081511f $X=5.3 $Y=2.04 $X2=0 $Y2=0
cc_566 N_A_997_119#_c_831_n N_VGND_c_1112_n 0.00902802f $X=5.365 $Y=1.295 $X2=0
+ $Y2=0
cc_567 N_A_997_119#_c_832_n N_VGND_c_1112_n 0.0269871f $X=6.435 $Y=1.21 $X2=0
+ $Y2=0
cc_568 N_A_997_119#_c_836_n N_VGND_c_1112_n 0.0103632f $X=6.6 $Y=1.125 $X2=0
+ $Y2=0
cc_569 N_A_997_119#_c_831_n N_VGND_c_1117_n 0.00699308f $X=5.365 $Y=1.295 $X2=0
+ $Y2=0
cc_570 N_A_997_119#_c_836_n N_VGND_c_1120_n 0.00418224f $X=6.6 $Y=1.125 $X2=0
+ $Y2=0
cc_571 N_A_997_119#_c_831_n N_VGND_c_1123_n 0.0108649f $X=5.365 $Y=1.295 $X2=0
+ $Y2=0
cc_572 N_A_997_119#_c_836_n N_VGND_c_1123_n 0.00544287f $X=6.6 $Y=1.125 $X2=0
+ $Y2=0
cc_573 N_A_1401_22#_M1012_g N_VPWR_c_972_n 0.0236631f $X=8.165 $Y=0.79 $X2=0
+ $Y2=0
cc_574 N_A_1401_22#_M1012_g N_VPWR_c_973_n 0.00486043f $X=8.165 $Y=0.79 $X2=0
+ $Y2=0
cc_575 N_A_1401_22#_M1012_g N_VPWR_c_974_n 0.0088953f $X=8.165 $Y=0.79 $X2=0
+ $Y2=0
cc_576 N_A_1401_22#_M1012_g N_VPWR_c_966_n 0.00590357f $X=8.165 $Y=0.79 $X2=0
+ $Y2=0
cc_577 N_A_1401_22#_M1012_g N_Q_N_c_1084_n 0.0183592f $X=8.165 $Y=0.79 $X2=0
+ $Y2=0
cc_578 N_A_1401_22#_c_906_n N_Q_N_c_1084_n 0.0165993f $X=7.52 $Y=1.875 $X2=0
+ $Y2=0
cc_579 N_A_1401_22#_c_903_n N_VGND_c_1112_n 0.0021741f $X=7.335 $Y=0.185 $X2=0
+ $Y2=0
cc_580 N_A_1401_22#_c_902_n N_VGND_c_1113_n 0.0214317f $X=8.09 $Y=0.185 $X2=0
+ $Y2=0
cc_581 N_A_1401_22#_M1012_g N_VGND_c_1113_n 0.0046248f $X=8.165 $Y=0.79 $X2=0
+ $Y2=0
cc_582 N_A_1401_22#_c_905_n N_VGND_c_1113_n 0.0102906f $X=7.3 $Y=0.83 $X2=0
+ $Y2=0
cc_583 N_A_1401_22#_c_906_n N_VGND_c_1113_n 0.0140175f $X=7.52 $Y=1.875 $X2=0
+ $Y2=0
cc_584 N_A_1401_22#_c_907_n N_VGND_c_1113_n 0.00205992f $X=7.17 $Y=0.43 $X2=0
+ $Y2=0
cc_585 N_A_1401_22#_c_908_n N_VGND_c_1113_n 0.0153293f $X=7.3 $Y=0.43 $X2=0
+ $Y2=0
cc_586 N_A_1401_22#_c_909_n N_VGND_c_1113_n 0.0163513f $X=7.52 $Y=0.935 $X2=0
+ $Y2=0
cc_587 N_A_1401_22#_c_902_n N_VGND_c_1114_n 0.00480782f $X=8.09 $Y=0.185 $X2=0
+ $Y2=0
cc_588 N_A_1401_22#_c_903_n N_VGND_c_1120_n 0.0232791f $X=7.335 $Y=0.185 $X2=0
+ $Y2=0
cc_589 N_A_1401_22#_c_908_n N_VGND_c_1120_n 0.0197838f $X=7.3 $Y=0.43 $X2=0
+ $Y2=0
cc_590 N_A_1401_22#_c_902_n N_VGND_c_1121_n 0.00595723f $X=8.09 $Y=0.185 $X2=0
+ $Y2=0
cc_591 N_A_1401_22#_c_902_n N_VGND_c_1123_n 0.0264629f $X=8.09 $Y=0.185 $X2=0
+ $Y2=0
cc_592 N_A_1401_22#_c_903_n N_VGND_c_1123_n 0.0110402f $X=7.335 $Y=0.185 $X2=0
+ $Y2=0
cc_593 N_A_1401_22#_c_908_n N_VGND_c_1123_n 0.0108415f $X=7.3 $Y=0.43 $X2=0
+ $Y2=0
cc_594 N_A_1401_22#_c_909_n N_VGND_c_1123_n 0.00674826f $X=7.52 $Y=0.935 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_966_n N_Q_N_M1007_d 0.00369895f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_596 N_VPWR_c_966_n N_Q_M1017_d 0.00336915f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_597 N_VPWR_c_980_n Q 0.0181659f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_598 N_VPWR_c_966_n Q 0.0104192f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_599 N_A_440_463#_c_1070_n N_VGND_c_1119_n 0.00688882f $X=2.555 $Y=0.8 $X2=0
+ $Y2=0
cc_600 N_A_440_463#_c_1070_n N_VGND_c_1123_n 0.0112304f $X=2.555 $Y=0.8 $X2=0
+ $Y2=0
cc_601 N_Q_N_c_1084_n N_VGND_c_1113_n 0.00270636f $X=8.38 $Y=0.52 $X2=0 $Y2=0
cc_602 N_Q_N_c_1084_n N_VGND_c_1114_n 0.0652138f $X=8.38 $Y=0.52 $X2=0 $Y2=0
cc_603 N_Q_N_c_1084_n N_VGND_c_1121_n 0.012598f $X=8.38 $Y=0.52 $X2=0 $Y2=0
cc_604 N_Q_N_c_1084_n N_VGND_c_1123_n 0.0106048f $X=8.38 $Y=0.52 $X2=0 $Y2=0
cc_605 Q N_VGND_c_1114_n 0.00255964f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_606 Q N_VGND_c_1122_n 0.0108661f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_607 Q N_VGND_c_1123_n 0.00974763f $X=9.275 $Y=0.47 $X2=0 $Y2=0
