# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o21ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o21ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.210000 3.695000 1.245000 ;
        RECT 0.125000 1.245000 1.825000 1.515000 ;
        RECT 1.420000 1.075000 3.695000 1.210000 ;
        RECT 3.445000 1.245000 3.695000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.425000 3.275000 1.760000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.905000 1.210000 5.255000 1.435000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.881600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 1.930000 4.290000 2.100000 ;
        RECT 1.840000 2.100000 2.170000 2.735000 ;
        RECT 2.700000 2.100000 3.030000 2.735000 ;
        RECT 3.445000 1.755000 5.670000 1.925000 ;
        RECT 3.445000 1.925000 4.290000 1.930000 ;
        RECT 3.865000 1.605000 5.670000 1.755000 ;
        RECT 4.080000 2.100000 4.290000 3.075000 ;
        RECT 4.100000 0.700000 5.670000 1.030000 ;
        RECT 4.960000 1.925000 5.150000 3.075000 ;
        RECT 5.425000 1.030000 5.670000 1.605000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.120000  0.255000 0.380000 0.870000 ;
      RECT 0.120000  0.870000 3.930000 0.905000 ;
      RECT 0.120000  0.905000 1.250000 1.040000 ;
      RECT 0.120000  1.815000 0.405000 3.245000 ;
      RECT 0.550000  0.085000 0.880000 0.700000 ;
      RECT 0.575000  1.755000 1.670000 1.925000 ;
      RECT 0.575000  1.925000 0.810000 3.075000 ;
      RECT 0.980000  2.095000 1.310000 3.245000 ;
      RECT 1.050000  0.255000 1.240000 0.735000 ;
      RECT 1.050000  0.735000 3.930000 0.870000 ;
      RECT 1.410000  0.085000 1.740000 0.565000 ;
      RECT 1.480000  1.925000 1.670000 2.905000 ;
      RECT 1.480000  2.905000 3.410000 3.075000 ;
      RECT 1.910000  0.255000 2.100000 0.735000 ;
      RECT 2.270000  0.085000 2.600000 0.565000 ;
      RECT 2.340000  2.270000 2.530000 2.905000 ;
      RECT 2.770000  0.255000 2.960000 0.735000 ;
      RECT 3.130000  0.085000 3.460000 0.565000 ;
      RECT 3.200000  2.270000 3.410000 2.905000 ;
      RECT 3.580000  2.270000 3.910000 3.245000 ;
      RECT 3.630000  0.255000 5.650000 0.530000 ;
      RECT 3.630000  0.530000 3.930000 0.735000 ;
      RECT 4.460000  2.095000 4.790000 3.245000 ;
      RECT 5.320000  2.105000 5.650000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__o21ai_4
END LIBRARY
