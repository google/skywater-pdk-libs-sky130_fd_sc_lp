* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_35_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_290_367# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_290_367# A2 a_35_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_35_367# A2 a_290_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND A1 a_35_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_35_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_710_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND A2 a_35_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VGND A3 a_35_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_35_47# B1 a_710_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_35_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Y A3 a_290_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_710_47# B1 a_35_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 Y C1 a_710_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_35_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VPWR A1 a_35_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
