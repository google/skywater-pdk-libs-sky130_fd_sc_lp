* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_123_480# C a_195_480# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_195_480# B a_267_480# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_267_480# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_40_480# D a_123_480# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VGND D a_40_480# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_40_480# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_40_480# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND B a_40_480# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_40_480# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR a_40_480# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
