* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfxtp_4 CLK D VGND VNB VPB VPWR Q
X0 VGND CLK a_110_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_941_379# a_110_70# a_1070_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_941_379# a_1112_93# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VPWR a_1112_93# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_684_93# a_110_70# a_941_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X5 VGND a_1112_93# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_526_413# a_217_413# a_642_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_941_379# a_1112_93# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR D a_431_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VGND D a_431_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR CLK a_110_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VGND a_526_413# a_684_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 Q a_1112_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_431_119# a_110_70# a_526_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_941_379# a_217_413# a_1116_441# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_1116_441# a_1112_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 Q a_1112_93# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_217_413# a_110_70# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VGND a_1112_93# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 Q a_1112_93# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_526_413# a_110_70# a_666_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_217_413# a_110_70# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_642_119# a_684_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_666_413# a_684_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_431_119# a_217_413# a_526_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_1070_119# a_1112_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 Q a_1112_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 a_684_93# a_217_413# a_941_379# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR a_526_413# a_684_93# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X29 VPWR a_1112_93# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
