* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 VGND a_27_114# a_196_462# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_304_533# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VPWR RESET_B a_559_533# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND a_1832_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_1417_133# a_1467_419# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_559_533# a_27_114# a_653_533# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_492_149# D a_304_533# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_695_375# a_27_114# a_1247_89# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_1832_367# a_1247_89# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_1247_89# a_196_462# a_1379_517# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1593_133# a_1247_89# a_1467_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_304_533# a_196_462# a_559_533# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VPWR a_27_114# a_196_462# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VPWR D a_304_533# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_803_149# a_695_375# a_875_149# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_695_375# a_196_462# a_1247_89# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VGND RESET_B a_492_149# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_559_533# a_695_375# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 VGND RESET_B a_1593_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_27_114# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_304_533# a_27_114# a_559_533# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_559_533# a_196_462# a_803_149# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1467_419# a_1247_89# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_27_114# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_1832_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_1832_367# a_1247_89# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1247_89# a_27_114# a_1417_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_875_149# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_653_533# a_695_375# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VPWR RESET_B a_1467_419# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 VGND a_559_533# a_695_375# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X31 a_1379_517# a_1467_419# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
