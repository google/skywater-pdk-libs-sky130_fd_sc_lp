* File: sky130_fd_sc_lp__dlclkp_4.spice
* Created: Fri Aug 28 10:25:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlclkp_4.pex.spice"
.subckt sky130_fd_sc_lp__dlclkp_4  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1022 N_VGND_M1022_d N_A_73_269#_M1022_g N_A_27_367#_M1022_s VNB NSHORT L=0.15
+ W=0.84 AD=0.22485 AS=0.2226 PD=1.84 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1009 A_253_81# N_GATE_M1009_g N_VGND_M1022_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.112425 PD=0.63 PS=0.92 NRD=14.28 NRS=74.28 M=1 R=2.8 SA=75000.9
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1001 N_A_73_269#_M1001_d N_A_295_55#_M1001_g A_253_81# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1014 A_411_81# N_A_277_367#_M1014_g N_A_73_269#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_27_367#_M1010_g A_411_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.08295 AS=0.0672 PD=0.815 PS=0.74 NRD=32.856 NRS=30 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_277_367#_M1008_d N_A_295_55#_M1008_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.08295 PD=1.37 PS=0.815 NRD=0 NRS=0 M=1 R=2.8 SA=75002.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_CLK_M1024_g N_A_295_55#_M1024_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0952 AS=0.1999 PD=0.823333 PS=1.86 NRD=49.044 NRS=34.284 M=1 R=2.8
+ SA=75000.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 A_1026_47# N_CLK_M1005_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1904 PD=1.05 PS=1.64667 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1002 N_A_1078_367#_M1002_d N_A_27_367#_M1002_g A_1026_47# VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_GCLK_M1004_d N_A_1078_367#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1013 N_GCLK_M1004_d N_A_1078_367#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1015 N_GCLK_M1015_d N_A_1078_367#_M1015_g N_VGND_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1019 N_GCLK_M1015_d N_A_1078_367#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1025 N_VPWR_M1025_d N_A_73_269#_M1025_g N_A_27_367#_M1025_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.369943 AS=0.3339 PD=2.42716 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1006 A_235_465# N_GATE_M1006_g N_VPWR_M1025_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.187907 PD=0.85 PS=1.23284 NRD=15.3857 NRS=73.4416 M=1 R=4.26667
+ SA=75000.8 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1020 N_A_73_269#_M1020_d N_A_277_367#_M1020_g A_235_465# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.134098 AS=0.0672 PD=1.24377 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.2 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1007 A_415_465# N_A_295_55#_M1007_g N_A_73_269#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0880019 PD=0.63 PS=0.816226 NRD=23.443 NRS=51.5943 M=1
+ R=2.8 SA=75001.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_27_367#_M1011_g A_415_465# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.204037 AS=0.0441 PD=1.20453 PS=0.63 NRD=56.2829 NRS=23.443 M=1 R=2.8
+ SA=75002.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 N_A_277_367#_M1021_d N_A_295_55#_M1021_g N_VPWR_M1011_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.225 AS=0.310913 PD=2.03 PS=1.83547 NRD=21.5321 NRS=93.8705
+ M=1 R=4.26667 SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_295_55#_M1012_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.176505 AS=0.27485 PD=1.16547 PS=2.21 NRD=67.9453 NRS=36.9375 M=1
+ R=4.26667 SA=75000.3 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1000 N_A_1078_367#_M1000_d N_CLK_M1000_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.347495 PD=1.54 PS=2.29453 NRD=0 NRS=14.8341 M=1 R=8.4
+ SA=75000.6 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_A_27_367#_M1017_g N_A_1078_367#_M1000_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75002 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1017_d N_A_1078_367#_M1003_g N_GCLK_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_A_1078_367#_M1016_g N_GCLK_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1016_d N_A_1078_367#_M1018_g N_GCLK_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1023 N_VPWR_M1023_d N_A_1078_367#_M1023_g N_GCLK_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.4221 AS=0.1764 PD=3.19 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75000.3 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=15.9817 P=20.94
c_87 VNB 0 1.79399e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dlclkp_4.pxi.spice"
*
.ends
*
*
