* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a311o_lp A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_257_414# B1 a_596_414# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_257_414# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VGND A3 a_294_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_596_414# C1 a_85_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 VPWR A3 a_257_414# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_372_47# A1 a_85_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_694_47# C1 a_85_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR A1 a_257_414# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_85_21# B1 a_536_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_115_47# a_85_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_294_47# A2 a_372_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_85_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 X a_85_21# a_115_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_536_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND C1 a_694_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
