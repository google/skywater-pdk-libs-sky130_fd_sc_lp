* File: sky130_fd_sc_lp__nand2_4.pxi.spice
* Created: Wed Sep  2 10:02:50 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2_4%B N_B_M1005_g N_B_M1000_g N_B_M1006_g N_B_M1001_g
+ N_B_M1013_g N_B_M1008_g N_B_M1015_g N_B_M1010_g B B B B N_B_c_68_n
+ PM_SKY130_FD_SC_LP__NAND2_4%B
x_PM_SKY130_FD_SC_LP__NAND2_4%A N_A_M1002_g N_A_M1004_g N_A_M1003_g N_A_M1007_g
+ N_A_M1009_g N_A_M1012_g N_A_M1011_g N_A_M1014_g N_A_c_142_n A A N_A_c_143_n
+ N_A_c_144_n PM_SKY130_FD_SC_LP__NAND2_4%A
x_PM_SKY130_FD_SC_LP__NAND2_4%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1010_d
+ N_VPWR_M1007_d N_VPWR_M1014_d N_VPWR_c_224_n N_VPWR_c_225_n N_VPWR_c_226_n
+ N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n N_VPWR_c_230_n N_VPWR_c_231_n
+ VPWR N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_235_n
+ N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_223_n PM_SKY130_FD_SC_LP__NAND2_4%VPWR
x_PM_SKY130_FD_SC_LP__NAND2_4%Y N_Y_M1002_s N_Y_M1009_s N_Y_M1000_s N_Y_M1008_s
+ N_Y_M1004_s N_Y_M1012_s N_Y_c_291_n N_Y_c_294_n N_Y_c_353_n N_Y_c_307_n
+ N_Y_c_295_n N_Y_c_318_n N_Y_c_290_n N_Y_c_326_n N_Y_c_330_n N_Y_c_333_n
+ N_Y_c_336_n Y Y Y Y Y Y Y N_Y_c_301_n N_Y_c_305_n N_Y_c_341_n
+ PM_SKY130_FD_SC_LP__NAND2_4%Y
x_PM_SKY130_FD_SC_LP__NAND2_4%A_63_65# N_A_63_65#_M1005_d N_A_63_65#_M1006_d
+ N_A_63_65#_M1015_d N_A_63_65#_M1003_d N_A_63_65#_M1011_d N_A_63_65#_c_377_n
+ N_A_63_65#_c_378_n N_A_63_65#_c_379_n N_A_63_65#_c_380_n N_A_63_65#_c_381_n
+ N_A_63_65#_c_382_n N_A_63_65#_c_383_n N_A_63_65#_c_416_n N_A_63_65#_c_384_n
+ N_A_63_65#_c_385_n N_A_63_65#_c_386_n N_A_63_65#_c_387_n
+ PM_SKY130_FD_SC_LP__NAND2_4%A_63_65#
x_PM_SKY130_FD_SC_LP__NAND2_4%VGND N_VGND_M1005_s N_VGND_M1013_s N_VGND_c_441_n
+ N_VGND_c_442_n VGND N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n
+ N_VGND_c_446_n N_VGND_c_447_n PM_SKY130_FD_SC_LP__NAND2_4%VGND
cc_1 VNB N_B_M1005_g 0.0259905f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.745
cc_2 VNB N_B_M1006_g 0.0190925f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.745
cc_3 VNB N_B_M1013_g 0.0190925f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.745
cc_4 VNB N_B_M1015_g 0.0193908f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.745
cc_5 VNB B 0.00384779f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_6 VNB N_B_c_68_n 0.076159f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=1.51
cc_7 VNB N_A_M1002_g 0.0194306f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.745
cc_8 VNB N_A_M1003_g 0.0204882f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.745
cc_9 VNB N_A_M1009_g 0.0208827f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.745
cc_10 VNB N_A_M1011_g 0.0268416f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.745
cc_11 VNB N_A_c_142_n 0.0280738f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_12 VNB N_A_c_143_n 0.0204866f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.51
cc_13 VNB N_A_c_144_n 0.0385524f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.51
cc_14 VNB N_VPWR_c_223_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_290_n 0.00680324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_63_65#_c_377_n 0.0311325f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.745
cc_17 VNB N_A_63_65#_c_378_n 0.00415273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_63_65#_c_379_n 0.0130877f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.675
cc_19 VNB N_A_63_65#_c_380_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_63_65#_c_381_n 0.00558452f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.745
cc_21 VNB N_A_63_65#_c_382_n 0.00273868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_63_65#_c_383_n 0.00185825f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_23 VNB N_A_63_65#_c_384_n 0.0120288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_63_65#_c_385_n 0.0327872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_63_65#_c_386_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.51
cc_26 VNB N_A_63_65#_c_387_n 0.00260516f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.51
cc_27 VNB N_VGND_c_441_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.745
cc_28 VNB N_VGND_c_442_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=2.465
cc_29 VNB N_VGND_c_443_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.745
cc_30 VNB N_VGND_c_444_n 0.0591389f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=1.675
cc_31 VNB N_VGND_c_445_n 0.25792f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=2.465
cc_32 VNB N_VGND_c_446_n 0.0275008f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_33 VNB N_VGND_c_447_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_34 VPB N_B_M1000_g 0.0249963f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.465
cc_35 VPB N_B_M1001_g 0.0178543f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=2.465
cc_36 VPB N_B_M1008_g 0.0178551f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=2.465
cc_37 VPB N_B_M1010_g 0.0179936f $X=-0.19 $Y=1.655 $X2=1.945 $Y2=2.465
cc_38 VPB B 0.010677f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.58
cc_39 VPB N_B_c_68_n 0.0130046f $X=-0.19 $Y=1.655 $X2=1.945 $Y2=1.51
cc_40 VPB N_A_M1004_g 0.0181192f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.465
cc_41 VPB N_A_M1007_g 0.019687f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=2.465
cc_42 VPB N_A_M1012_g 0.0196902f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=2.465
cc_43 VPB N_A_M1014_g 0.0252407f $X=-0.19 $Y=1.655 $X2=1.945 $Y2=2.465
cc_44 VPB N_A_c_142_n 0.00448375f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_45 VPB A 0.00676829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_c_143_n 0.00836278f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.51
cc_47 VPB N_A_c_144_n 0.00519541f $X=-0.19 $Y=1.655 $X2=1.48 $Y2=1.51
cc_48 VPB N_VPWR_c_224_n 0.0127022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_225_n 0.0648945f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=0.745
cc_50 VPB N_VPWR_c_226_n 0.0172428f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=2.465
cc_51 VPB N_VPWR_c_227_n 3.31161e-19 $X=-0.19 $Y=1.655 $X2=1.945 $Y2=0.745
cc_52 VPB N_VPWR_c_228_n 3.20114e-19 $X=-0.19 $Y=1.655 $X2=1.945 $Y2=2.465
cc_53 VPB N_VPWR_c_229_n 0.00493206f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_54 VPB N_VPWR_c_230_n 0.0109406f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.58
cc_55 VPB N_VPWR_c_231_n 0.0581494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_232_n 0.0130076f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.51
cc_57 VPB N_VPWR_c_233_n 0.0155347f $X=-0.19 $Y=1.655 $X2=1.48 $Y2=1.51
cc_58 VPB N_VPWR_c_234_n 0.0187451f $X=-0.19 $Y=1.655 $X2=1.945 $Y2=1.51
cc_59 VPB N_VPWR_c_235_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.592
cc_60 VPB N_VPWR_c_236_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.592
cc_61 VPB N_VPWR_c_237_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_223_n 0.0456494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 N_B_M1015_g N_A_M1002_g 0.0237751f $X=1.945 $Y=0.745 $X2=0 $Y2=0
cc_64 N_B_M1010_g N_A_M1004_g 0.0237751f $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_65 B N_A_c_142_n 0.00320661f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_66 N_B_c_68_n N_A_c_142_n 0.0237751f $X=1.945 $Y=1.51 $X2=0 $Y2=0
cc_67 N_B_M1000_g N_VPWR_c_225_n 0.0322235f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_68 N_B_M1000_g N_VPWR_c_226_n 0.00445288f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_69 N_B_M1001_g N_VPWR_c_226_n 0.00486043f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_70 N_B_M1000_g N_VPWR_c_227_n 5.38496e-19 $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_71 N_B_M1001_g N_VPWR_c_227_n 0.0145257f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_72 N_B_M1008_g N_VPWR_c_227_n 0.0141795f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_73 N_B_M1010_g N_VPWR_c_227_n 6.90936e-19 $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_74 N_B_M1008_g N_VPWR_c_228_n 6.90936e-19 $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_75 N_B_M1010_g N_VPWR_c_228_n 0.0140981f $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_76 N_B_M1008_g N_VPWR_c_232_n 0.00486043f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_77 N_B_M1010_g N_VPWR_c_232_n 0.00486043f $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_78 N_B_M1000_g N_VPWR_c_223_n 0.00863667f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_79 N_B_M1001_g N_VPWR_c_223_n 0.00830891f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_80 N_B_M1008_g N_VPWR_c_223_n 0.00830891f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_81 N_B_M1010_g N_VPWR_c_223_n 0.00830891f $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_82 N_B_M1000_g N_Y_c_291_n 0.00458304f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_83 B N_Y_c_291_n 0.0248473f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_84 N_B_c_68_n N_Y_c_291_n 6.37898e-19 $X=1.945 $Y=1.51 $X2=0 $Y2=0
cc_85 N_B_M1000_g N_Y_c_294_n 0.0150492f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_86 N_B_M1015_g N_Y_c_295_n 9.13036e-19 $X=1.945 $Y=0.745 $X2=0 $Y2=0
cc_87 N_B_M1010_g N_Y_c_295_n 8.31125e-19 $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_88 B N_Y_c_295_n 0.026859f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_89 N_B_c_68_n N_Y_c_295_n 2.44965e-19 $X=1.945 $Y=1.51 $X2=0 $Y2=0
cc_90 B Y 0.0154121f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_91 N_B_c_68_n Y 6.37898e-19 $X=1.945 $Y=1.51 $X2=0 $Y2=0
cc_92 N_B_M1001_g N_Y_c_301_n 0.0134574f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_93 N_B_M1008_g N_Y_c_301_n 0.0134574f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_94 B N_Y_c_301_n 0.0433781f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_95 N_B_c_68_n N_Y_c_301_n 5.73944e-19 $X=1.945 $Y=1.51 $X2=0 $Y2=0
cc_96 N_B_M1010_g N_Y_c_305_n 0.0133997f $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_97 B N_Y_c_305_n 0.0283474f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_98 N_B_M1005_g N_A_63_65#_c_377_n 0.00354503f $X=0.655 $Y=0.745 $X2=0 $Y2=0
cc_99 N_B_M1005_g N_A_63_65#_c_378_n 0.0157256f $X=0.655 $Y=0.745 $X2=0 $Y2=0
cc_100 N_B_M1006_g N_A_63_65#_c_378_n 0.0133326f $X=1.085 $Y=0.745 $X2=0 $Y2=0
cc_101 B N_A_63_65#_c_378_n 0.0419365f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_102 N_B_c_68_n N_A_63_65#_c_378_n 0.00246472f $X=1.945 $Y=1.51 $X2=0 $Y2=0
cc_103 N_B_M1006_g N_A_63_65#_c_380_n 8.28776e-19 $X=1.085 $Y=0.745 $X2=0 $Y2=0
cc_104 N_B_M1013_g N_A_63_65#_c_380_n 8.28776e-19 $X=1.515 $Y=0.745 $X2=0 $Y2=0
cc_105 N_B_M1013_g N_A_63_65#_c_381_n 0.013286f $X=1.515 $Y=0.745 $X2=0 $Y2=0
cc_106 N_B_M1015_g N_A_63_65#_c_381_n 0.0130971f $X=1.945 $Y=0.745 $X2=0 $Y2=0
cc_107 B N_A_63_65#_c_381_n 0.0653436f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_108 N_B_c_68_n N_A_63_65#_c_381_n 0.00246472f $X=1.945 $Y=1.51 $X2=0 $Y2=0
cc_109 N_B_M1015_g N_A_63_65#_c_383_n 4.90985e-19 $X=1.945 $Y=0.745 $X2=0 $Y2=0
cc_110 B N_A_63_65#_c_386_n 0.0160407f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_111 N_B_c_68_n N_A_63_65#_c_386_n 0.00256759f $X=1.945 $Y=1.51 $X2=0 $Y2=0
cc_112 N_B_M1005_g N_VGND_c_441_n 0.012533f $X=0.655 $Y=0.745 $X2=0 $Y2=0
cc_113 N_B_M1006_g N_VGND_c_441_n 0.0102222f $X=1.085 $Y=0.745 $X2=0 $Y2=0
cc_114 N_B_M1013_g N_VGND_c_441_n 5.123e-19 $X=1.515 $Y=0.745 $X2=0 $Y2=0
cc_115 N_B_M1006_g N_VGND_c_442_n 5.123e-19 $X=1.085 $Y=0.745 $X2=0 $Y2=0
cc_116 N_B_M1013_g N_VGND_c_442_n 0.0102222f $X=1.515 $Y=0.745 $X2=0 $Y2=0
cc_117 N_B_M1015_g N_VGND_c_442_n 0.0103482f $X=1.945 $Y=0.745 $X2=0 $Y2=0
cc_118 N_B_M1006_g N_VGND_c_443_n 0.00414769f $X=1.085 $Y=0.745 $X2=0 $Y2=0
cc_119 N_B_M1013_g N_VGND_c_443_n 0.00414769f $X=1.515 $Y=0.745 $X2=0 $Y2=0
cc_120 N_B_M1015_g N_VGND_c_444_n 0.00414769f $X=1.945 $Y=0.745 $X2=0 $Y2=0
cc_121 N_B_M1005_g N_VGND_c_445_n 0.00828433f $X=0.655 $Y=0.745 $X2=0 $Y2=0
cc_122 N_B_M1006_g N_VGND_c_445_n 0.00787505f $X=1.085 $Y=0.745 $X2=0 $Y2=0
cc_123 N_B_M1013_g N_VGND_c_445_n 0.00787505f $X=1.515 $Y=0.745 $X2=0 $Y2=0
cc_124 N_B_M1015_g N_VGND_c_445_n 0.0078848f $X=1.945 $Y=0.745 $X2=0 $Y2=0
cc_125 N_B_M1005_g N_VGND_c_446_n 0.00414769f $X=0.655 $Y=0.745 $X2=0 $Y2=0
cc_126 N_A_M1004_g N_VPWR_c_228_n 0.0142658f $X=2.375 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_M1007_g N_VPWR_c_228_n 5.079e-19 $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_M1007_g N_VPWR_c_229_n 0.00675679f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A_M1012_g N_VPWR_c_229_n 0.0108528f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A_M1014_g N_VPWR_c_231_n 0.00914801f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A_M1004_g N_VPWR_c_233_n 0.00486043f $X=2.375 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A_M1007_g N_VPWR_c_233_n 0.00557067f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A_M1012_g N_VPWR_c_234_n 0.00512356f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A_M1014_g N_VPWR_c_234_n 0.00557067f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_M1004_g N_VPWR_c_223_n 0.00830891f $X=2.375 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_M1007_g N_VPWR_c_223_n 0.0104944f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_M1012_g N_VPWR_c_223_n 0.00946541f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A_M1014_g N_VPWR_c_223_n 0.0109505f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_M1002_g N_Y_c_307_n 0.00497669f $X=2.375 $Y=0.745 $X2=0 $Y2=0
cc_140 N_A_M1003_g N_Y_c_307_n 0.00689779f $X=2.805 $Y=0.745 $X2=0 $Y2=0
cc_141 N_A_M1009_g N_Y_c_307_n 8.23603e-19 $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_142 N_A_M1002_g N_Y_c_295_n 0.00288853f $X=2.375 $Y=0.745 $X2=0 $Y2=0
cc_143 N_A_M1004_g N_Y_c_295_n 0.00665818f $X=2.375 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_M1003_g N_Y_c_295_n 0.00320441f $X=2.805 $Y=0.745 $X2=0 $Y2=0
cc_145 N_A_M1007_g N_Y_c_295_n 0.00706476f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_M1009_g N_Y_c_295_n 4.44951e-19 $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_147 N_A_M1012_g N_Y_c_295_n 8.23875e-19 $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_c_142_n N_Y_c_295_n 0.0254759f $X=2.88 $Y=1.51 $X2=0 $Y2=0
cc_149 A N_Y_c_295_n 0.0277198f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A_M1007_g N_Y_c_318_n 0.0112046f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_M1012_g N_Y_c_318_n 6.66723e-19 $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_M1003_g N_Y_c_290_n 0.013753f $X=2.805 $Y=0.745 $X2=0 $Y2=0
cc_153 N_A_M1009_g N_Y_c_290_n 0.0113756f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_154 N_A_M1011_g N_Y_c_290_n 0.0052413f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_155 A N_Y_c_290_n 0.065912f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_156 N_A_c_143_n N_Y_c_290_n 0.0063321f $X=3.32 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A_c_144_n N_Y_c_290_n 0.00252688f $X=3.825 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A_M1012_g N_Y_c_326_n 0.00167925f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A_M1014_g N_Y_c_326_n 0.00244933f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_160 A N_Y_c_326_n 0.0247573f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_161 N_A_c_144_n N_Y_c_326_n 6.37898e-19 $X=3.825 $Y=1.51 $X2=0 $Y2=0
cc_162 N_A_M1007_g N_Y_c_330_n 7.03279e-19 $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_M1012_g N_Y_c_330_n 0.0134008f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A_M1014_g N_Y_c_330_n 0.00983347f $X=3.825 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_M1003_g N_Y_c_333_n 8.36143e-19 $X=2.805 $Y=0.745 $X2=0 $Y2=0
cc_166 N_A_M1009_g N_Y_c_333_n 0.00740195f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_167 N_A_M1011_g N_Y_c_333_n 0.00532386f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_168 N_A_M1002_g N_Y_c_336_n 0.00266514f $X=2.375 $Y=0.745 $X2=0 $Y2=0
cc_169 N_A_M1003_g N_Y_c_336_n 0.0013353f $X=2.805 $Y=0.745 $X2=0 $Y2=0
cc_170 N_A_M1004_g Y 0.00166864f $X=2.375 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A_M1007_g Y 4.74589e-19 $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A_M1004_g N_Y_c_305_n 0.0153388f $X=2.375 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A_M1007_g N_Y_c_341_n 0.0171461f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_M1012_g N_Y_c_341_n 0.0112706f $X=3.395 $Y=2.465 $X2=0 $Y2=0
cc_175 A N_Y_c_341_n 0.0360207f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A_c_143_n N_Y_c_341_n 0.00149225f $X=3.32 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A_M1002_g N_A_63_65#_c_381_n 7.36763e-19 $X=2.375 $Y=0.745 $X2=0 $Y2=0
cc_178 N_A_M1002_g N_A_63_65#_c_382_n 0.0117986f $X=2.375 $Y=0.745 $X2=0 $Y2=0
cc_179 N_A_M1003_g N_A_63_65#_c_382_n 0.0120312f $X=2.805 $Y=0.745 $X2=0 $Y2=0
cc_180 N_A_M1009_g N_A_63_65#_c_384_n 0.0119222f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_181 N_A_M1011_g N_A_63_65#_c_384_n 0.012423f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_182 N_A_M1011_g N_A_63_65#_c_385_n 0.00354524f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_183 N_A_M1002_g N_VGND_c_442_n 5.59621e-19 $X=2.375 $Y=0.745 $X2=0 $Y2=0
cc_184 N_A_M1002_g N_VGND_c_444_n 0.0030414f $X=2.375 $Y=0.745 $X2=0 $Y2=0
cc_185 N_A_M1003_g N_VGND_c_444_n 0.0030414f $X=2.805 $Y=0.745 $X2=0 $Y2=0
cc_186 N_A_M1009_g N_VGND_c_444_n 0.0030414f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_187 N_A_M1011_g N_VGND_c_444_n 0.0030414f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_188 N_A_M1002_g N_VGND_c_445_n 0.00435814f $X=2.375 $Y=0.745 $X2=0 $Y2=0
cc_189 N_A_M1003_g N_VGND_c_445_n 0.00448682f $X=2.805 $Y=0.745 $X2=0 $Y2=0
cc_190 N_A_M1009_g N_VGND_c_445_n 0.00448682f $X=3.395 $Y=0.745 $X2=0 $Y2=0
cc_191 N_A_M1011_g N_VGND_c_445_n 0.00471417f $X=3.825 $Y=0.745 $X2=0 $Y2=0
cc_192 N_VPWR_c_223_n N_Y_M1000_s 0.00380684f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_223_n N_Y_M1008_s 0.00537116f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_c_223_n N_Y_M1004_s 0.00380684f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_223_n N_Y_M1012_s 0.00224253f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_225_n N_Y_c_291_n 0.0173425f $X=0.38 $Y=1.97 $X2=0 $Y2=0
cc_197 N_VPWR_c_225_n N_Y_c_294_n 0.0711533f $X=0.38 $Y=1.97 $X2=0 $Y2=0
cc_198 N_VPWR_c_226_n N_Y_c_294_n 0.0181313f $X=1.135 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_223_n N_Y_c_294_n 0.0121208f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_200 N_VPWR_c_232_n N_Y_c_353_n 0.0110383f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_223_n N_Y_c_353_n 0.00723852f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_c_233_n N_Y_c_318_n 0.0136146f $X=2.92 $Y=3.33 $X2=0 $Y2=0
cc_203 N_VPWR_c_223_n N_Y_c_318_n 0.00958075f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_c_229_n N_Y_c_330_n 0.0580832f $X=3.085 $Y=2.395 $X2=0 $Y2=0
cc_205 N_VPWR_c_234_n N_Y_c_330_n 0.0179976f $X=3.94 $Y=3.33 $X2=0 $Y2=0
cc_206 N_VPWR_c_223_n N_Y_c_330_n 0.012939f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_207 N_VPWR_M1001_d N_Y_c_301_n 0.00335356f $X=1.16 $Y=1.835 $X2=0 $Y2=0
cc_208 N_VPWR_c_227_n N_Y_c_301_n 0.0173266f $X=1.3 $Y=2.395 $X2=0 $Y2=0
cc_209 N_VPWR_M1010_d N_Y_c_305_n 0.00355663f $X=2.02 $Y=1.835 $X2=0 $Y2=0
cc_210 N_VPWR_c_228_n N_Y_c_305_n 0.0173266f $X=2.16 $Y=2.395 $X2=0 $Y2=0
cc_211 N_VPWR_M1007_d N_Y_c_341_n 0.00777597f $X=2.88 $Y=1.835 $X2=0 $Y2=0
cc_212 N_VPWR_c_229_n N_Y_c_341_n 0.0257501f $X=3.085 $Y=2.395 $X2=0 $Y2=0
cc_213 N_VPWR_c_225_n N_A_63_65#_c_379_n 0.00738849f $X=0.38 $Y=1.97 $X2=0 $Y2=0
cc_214 N_VPWR_c_231_n N_A_63_65#_c_385_n 0.00964856f $X=4.04 $Y=1.98 $X2=0 $Y2=0
cc_215 N_Y_c_290_n N_A_63_65#_M1003_d 0.00385954f $X=3.435 $Y=1.16 $X2=0 $Y2=0
cc_216 N_Y_c_295_n N_A_63_65#_c_381_n 8.05502e-19 $X=2.59 $Y=1.93 $X2=0 $Y2=0
cc_217 N_Y_c_336_n N_A_63_65#_c_381_n 0.0104705f $X=2.59 $Y=1.16 $X2=0 $Y2=0
cc_218 N_Y_M1002_s N_A_63_65#_c_382_n 0.00180746f $X=2.45 $Y=0.325 $X2=0 $Y2=0
cc_219 N_Y_c_307_n N_A_63_65#_c_382_n 0.015238f $X=2.59 $Y=0.7 $X2=0 $Y2=0
cc_220 N_Y_c_290_n N_A_63_65#_c_382_n 0.00280043f $X=3.435 $Y=1.16 $X2=0 $Y2=0
cc_221 N_Y_c_290_n N_A_63_65#_c_416_n 0.0263919f $X=3.435 $Y=1.16 $X2=0 $Y2=0
cc_222 N_Y_M1009_s N_A_63_65#_c_384_n 0.00176461f $X=3.47 $Y=0.325 $X2=0 $Y2=0
cc_223 N_Y_c_290_n N_A_63_65#_c_384_n 0.0025755f $X=3.435 $Y=1.16 $X2=0 $Y2=0
cc_224 N_Y_c_333_n N_A_63_65#_c_384_n 0.0166505f $X=3.61 $Y=0.69 $X2=0 $Y2=0
cc_225 N_Y_c_290_n N_A_63_65#_c_385_n 0.00539933f $X=3.435 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_63_65#_c_378_n N_VGND_M1005_s 0.00176461f $X=1.205 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_63_65#_c_381_n N_VGND_M1013_s 0.00176461f $X=2.065 $Y=1.17 $X2=0
+ $Y2=0
cc_228 N_A_63_65#_c_377_n N_VGND_c_441_n 0.0236466f $X=0.44 $Y=0.47 $X2=0 $Y2=0
cc_229 N_A_63_65#_c_378_n N_VGND_c_441_n 0.0170777f $X=1.205 $Y=1.17 $X2=0 $Y2=0
cc_230 N_A_63_65#_c_380_n N_VGND_c_441_n 0.0236157f $X=1.3 $Y=0.47 $X2=0 $Y2=0
cc_231 N_A_63_65#_c_380_n N_VGND_c_442_n 0.0236157f $X=1.3 $Y=0.47 $X2=0 $Y2=0
cc_232 N_A_63_65#_c_381_n N_VGND_c_442_n 0.0170777f $X=2.065 $Y=1.17 $X2=0 $Y2=0
cc_233 N_A_63_65#_c_383_n N_VGND_c_442_n 0.00915965f $X=2.255 $Y=0.35 $X2=0
+ $Y2=0
cc_234 N_A_63_65#_c_380_n N_VGND_c_443_n 0.0102275f $X=1.3 $Y=0.47 $X2=0 $Y2=0
cc_235 N_A_63_65#_c_382_n N_VGND_c_444_n 0.0403176f $X=2.935 $Y=0.35 $X2=0 $Y2=0
cc_236 N_A_63_65#_c_383_n N_VGND_c_444_n 0.0128106f $X=2.255 $Y=0.35 $X2=0 $Y2=0
cc_237 N_A_63_65#_c_384_n N_VGND_c_444_n 0.0578479f $X=3.945 $Y=0.35 $X2=0 $Y2=0
cc_238 N_A_63_65#_c_387_n N_VGND_c_444_n 0.0221491f $X=3.1 $Y=0.35 $X2=0 $Y2=0
cc_239 N_A_63_65#_c_377_n N_VGND_c_445_n 0.0093995f $X=0.44 $Y=0.47 $X2=0 $Y2=0
cc_240 N_A_63_65#_c_380_n N_VGND_c_445_n 0.00712543f $X=1.3 $Y=0.47 $X2=0 $Y2=0
cc_241 N_A_63_65#_c_382_n N_VGND_c_445_n 0.024032f $X=2.935 $Y=0.35 $X2=0 $Y2=0
cc_242 N_A_63_65#_c_383_n N_VGND_c_445_n 0.0073517f $X=2.255 $Y=0.35 $X2=0 $Y2=0
cc_243 N_A_63_65#_c_384_n N_VGND_c_445_n 0.0340922f $X=3.945 $Y=0.35 $X2=0 $Y2=0
cc_244 N_A_63_65#_c_387_n N_VGND_c_445_n 0.0127478f $X=3.1 $Y=0.35 $X2=0 $Y2=0
cc_245 N_A_63_65#_c_377_n N_VGND_c_446_n 0.0134916f $X=0.44 $Y=0.47 $X2=0 $Y2=0
