* File: sky130_fd_sc_lp__fahcon_1.pxi.spice
* Created: Fri Aug 28 10:35:46 2020
* 
x_PM_SKY130_FD_SC_LP__FAHCON_1%A N_A_M1030_g N_A_M1025_g A N_A_c_218_n
+ N_A_c_219_n PM_SKY130_FD_SC_LP__FAHCON_1%A
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_33_367# N_A_33_367#_M1025_s N_A_33_367#_M1005_d
+ N_A_33_367#_M1030_s N_A_33_367#_M1013_d N_A_33_367#_M1021_g
+ N_A_33_367#_c_257_n N_A_33_367#_M1003_g N_A_33_367#_c_258_n
+ N_A_33_367#_c_269_n N_A_33_367#_c_281_n N_A_33_367#_c_259_n
+ N_A_33_367#_c_260_n N_A_33_367#_c_261_n N_A_33_367#_c_262_n
+ N_A_33_367#_c_263_n N_A_33_367#_c_271_n N_A_33_367#_c_264_n
+ N_A_33_367#_c_265_n N_A_33_367#_c_266_n N_A_33_367#_c_351_p
+ N_A_33_367#_c_274_n N_A_33_367#_c_267_n PM_SKY130_FD_SC_LP__FAHCON_1%A_33_367#
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_329_269# N_A_329_269#_M1011_s
+ N_A_329_269#_M1027_s N_A_329_269#_M1022_g N_A_329_269#_M1029_g
+ N_A_329_269#_c_375_n N_A_329_269#_M1001_g N_A_329_269#_M1000_g
+ N_A_329_269#_c_378_n N_A_329_269#_c_379_n N_A_329_269#_c_380_n
+ N_A_329_269#_c_388_n N_A_329_269#_c_389_n N_A_329_269#_c_381_n
+ N_A_329_269#_c_382_n N_A_329_269#_c_383_n N_A_329_269#_c_384_n
+ N_A_329_269#_c_385_n PM_SKY130_FD_SC_LP__FAHCON_1%A_329_269#
x_PM_SKY130_FD_SC_LP__FAHCON_1%B N_B_M1005_g N_B_M1013_g N_B_c_501_n N_B_c_502_n
+ N_B_M1018_g N_B_M1031_g N_B_c_504_n N_B_c_486_n N_B_c_487_n N_B_c_488_n
+ N_B_M1027_g N_B_c_490_n N_B_c_491_n N_B_M1011_g N_B_M1024_g N_B_c_493_n
+ N_B_c_494_n N_B_M1008_g N_B_c_496_n N_B_c_497_n N_B_c_510_n N_B_c_498_n B
+ N_B_c_499_n PM_SKY130_FD_SC_LP__FAHCON_1%B
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_367_119# N_A_367_119#_M1029_d
+ N_A_367_119#_M1000_d N_A_367_119#_M1010_g N_A_367_119#_M1009_g
+ N_A_367_119#_M1019_g N_A_367_119#_M1028_g N_A_367_119#_c_628_n
+ N_A_367_119#_c_629_n N_A_367_119#_c_648_n N_A_367_119#_c_630_n
+ N_A_367_119#_c_650_n N_A_367_119#_c_651_n N_A_367_119#_c_631_n
+ N_A_367_119#_c_632_n N_A_367_119#_c_633_n N_A_367_119#_c_634_n
+ N_A_367_119#_c_635_n N_A_367_119#_c_636_n N_A_367_119#_c_664_n
+ N_A_367_119#_c_637_n N_A_367_119#_c_638_n N_A_367_119#_c_639_n
+ N_A_367_119#_c_640_n N_A_367_119#_c_641_n N_A_367_119#_c_642_n
+ N_A_367_119#_c_774_p N_A_367_119#_c_643_n N_A_367_119#_c_644_n
+ N_A_367_119#_c_645_n N_A_367_119#_c_778_p
+ PM_SKY130_FD_SC_LP__FAHCON_1%A_367_119#
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_359_367# N_A_359_367#_M1001_d
+ N_A_359_367#_M1022_d N_A_359_367#_c_876_n N_A_359_367#_M1020_g
+ N_A_359_367#_c_877_n N_A_359_367#_M1014_g N_A_359_367#_M1002_g
+ N_A_359_367#_M1006_g N_A_359_367#_c_879_n N_A_359_367#_c_880_n
+ N_A_359_367#_c_889_n N_A_359_367#_c_890_n N_A_359_367#_c_900_n
+ N_A_359_367#_c_907_n N_A_359_367#_c_891_n N_A_359_367#_c_881_n
+ N_A_359_367#_c_882_n N_A_359_367#_c_892_n N_A_359_367#_c_902_n
+ N_A_359_367#_c_893_n N_A_359_367#_c_894_n N_A_359_367#_c_895_n
+ N_A_359_367#_c_883_n N_A_359_367#_c_884_n N_A_359_367#_c_885_n
+ PM_SKY130_FD_SC_LP__FAHCON_1%A_359_367#
x_PM_SKY130_FD_SC_LP__FAHCON_1%CI N_CI_M1026_g N_CI_c_1072_n N_CI_c_1073_n
+ N_CI_M1016_g N_CI_M1023_g N_CI_c_1075_n N_CI_M1012_g CI N_CI_c_1077_n
+ N_CI_c_1078_n PM_SKY130_FD_SC_LP__FAHCON_1%CI
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_1571_367# N_A_1571_367#_M1012_d
+ N_A_1571_367#_M1023_d N_A_1571_367#_M1028_d N_A_1571_367#_M1015_g
+ N_A_1571_367#_c_1141_n N_A_1571_367#_M1007_g N_A_1571_367#_c_1142_n
+ N_A_1571_367#_c_1143_n N_A_1571_367#_c_1137_n N_A_1571_367#_c_1144_n
+ N_A_1571_367#_c_1145_n N_A_1571_367#_c_1138_n N_A_1571_367#_c_1147_n
+ N_A_1571_367#_c_1158_n N_A_1571_367#_c_1148_n N_A_1571_367#_c_1149_n
+ N_A_1571_367#_c_1139_n N_A_1571_367#_c_1140_n
+ PM_SKY130_FD_SC_LP__FAHCON_1%A_1571_367#
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_1758_87# N_A_1758_87#_M1002_d
+ N_A_1758_87#_M1006_d N_A_1758_87#_c_1258_n N_A_1758_87#_M1017_g
+ N_A_1758_87#_M1004_g N_A_1758_87#_c_1271_n N_A_1758_87#_c_1260_n
+ N_A_1758_87#_c_1261_n N_A_1758_87#_c_1262_n N_A_1758_87#_c_1263_n
+ N_A_1758_87#_c_1319_n N_A_1758_87#_c_1331_p N_A_1758_87#_c_1320_n
+ N_A_1758_87#_c_1264_n N_A_1758_87#_c_1282_n N_A_1758_87#_c_1265_n
+ N_A_1758_87#_c_1266_n PM_SKY130_FD_SC_LP__FAHCON_1%A_1758_87#
x_PM_SKY130_FD_SC_LP__FAHCON_1%VPWR N_VPWR_M1030_d N_VPWR_M1027_d N_VPWR_M1026_d
+ N_VPWR_M1007_d N_VPWR_c_1361_n N_VPWR_c_1362_n N_VPWR_c_1363_n N_VPWR_c_1364_n
+ N_VPWR_c_1365_n N_VPWR_c_1366_n VPWR N_VPWR_c_1367_n N_VPWR_c_1368_n
+ N_VPWR_c_1369_n N_VPWR_c_1360_n N_VPWR_c_1371_n N_VPWR_c_1372_n
+ N_VPWR_c_1373_n PM_SKY130_FD_SC_LP__FAHCON_1%VPWR
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_247_367# N_A_247_367#_M1003_d
+ N_A_247_367#_M1031_d N_A_247_367#_M1021_d N_A_247_367#_M1018_d
+ N_A_247_367#_c_1468_n N_A_247_367#_c_1463_n N_A_247_367#_c_1473_n
+ N_A_247_367#_c_1464_n N_A_247_367#_c_1465_n N_A_247_367#_c_1458_n
+ N_A_247_367#_c_1459_n N_A_247_367#_c_1460_n N_A_247_367#_c_1461_n
+ N_A_247_367#_c_1462_n PM_SKY130_FD_SC_LP__FAHCON_1%A_247_367#
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_1034_380# N_A_1034_380#_M1008_d
+ N_A_1034_380#_M1024_d N_A_1034_380#_c_1533_n N_A_1034_380#_c_1534_n
+ N_A_1034_380#_c_1539_n N_A_1034_380#_c_1541_n N_A_1034_380#_c_1532_n
+ N_A_1034_380#_c_1547_n PM_SKY130_FD_SC_LP__FAHCON_1%A_1034_380#
x_PM_SKY130_FD_SC_LP__FAHCON_1%COUT_N N_COUT_N_M1020_d N_COUT_N_M1010_d
+ N_COUT_N_c_1586_n N_COUT_N_c_1583_n N_COUT_N_c_1584_n N_COUT_N_c_1585_n COUT_N
+ PM_SKY130_FD_SC_LP__FAHCON_1%COUT_N
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_1340_412# N_A_1340_412#_M1009_d
+ N_A_1340_412#_M1014_d N_A_1340_412#_c_1644_n N_A_1340_412#_c_1642_n
+ N_A_1340_412#_c_1643_n PM_SKY130_FD_SC_LP__FAHCON_1%A_1340_412#
x_PM_SKY130_FD_SC_LP__FAHCON_1%A_1708_411# N_A_1708_411#_M1019_d
+ N_A_1708_411#_M1006_s N_A_1708_411#_M1007_s N_A_1708_411#_c_1690_n
+ N_A_1708_411#_c_1696_n N_A_1708_411#_c_1687_n N_A_1708_411#_c_1688_n
+ N_A_1708_411#_c_1702_n N_A_1708_411#_c_1689_n N_A_1708_411#_c_1692_n
+ PM_SKY130_FD_SC_LP__FAHCON_1%A_1708_411#
x_PM_SKY130_FD_SC_LP__FAHCON_1%SUM N_SUM_M1017_d N_SUM_M1004_d SUM SUM SUM SUM
+ SUM SUM SUM N_SUM_c_1747_n PM_SKY130_FD_SC_LP__FAHCON_1%SUM
x_PM_SKY130_FD_SC_LP__FAHCON_1%VGND N_VGND_M1025_d N_VGND_M1011_d N_VGND_M1016_d
+ N_VGND_M1015_d N_VGND_c_1759_n N_VGND_c_1760_n N_VGND_c_1761_n N_VGND_c_1762_n
+ N_VGND_c_1763_n N_VGND_c_1764_n VGND N_VGND_c_1765_n N_VGND_c_1766_n
+ N_VGND_c_1767_n N_VGND_c_1768_n N_VGND_c_1769_n N_VGND_c_1770_n
+ N_VGND_c_1771_n PM_SKY130_FD_SC_LP__FAHCON_1%VGND
cc_1 VNB A 0.00272879f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_2 VNB N_A_c_218_n 0.0257259f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.51
cc_3 VNB N_A_c_219_n 0.0219375f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.345
cc_4 VNB N_A_33_367#_c_257_n 0.0182394f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.562
cc_5 VNB N_A_33_367#_c_258_n 0.0290812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_33_367#_c_259_n 0.00364577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_33_367#_c_260_n 0.0242665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_33_367#_c_261_n 0.00353434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_33_367#_c_262_n 0.0057425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_33_367#_c_263_n 0.00748956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_33_367#_c_264_n 0.0228819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_33_367#_c_265_n 2.29632e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_33_367#_c_266_n 0.00192411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_33_367#_c_267_n 0.0353959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_329_269#_M1022_g 0.0082291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_329_269#_M1029_g 0.0286502f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.675
cc_17 VNB N_A_329_269#_c_375_n 0.0130185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_329_269#_M1001_g 0.0128528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_329_269#_M1000_g 0.00469964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_329_269#_c_378_n 0.0107892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_329_269#_c_379_n 0.0119881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_329_269#_c_380_n 0.0204328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_329_269#_c_381_n 0.0714299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_329_269#_c_382_n 0.00281934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_329_269#_c_383_n 0.00852876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_329_269#_c_384_n 0.0174649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_329_269#_c_385_n 0.0568369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_M1005_g 0.0239871f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_29 VNB N_B_M1031_g 0.0290019f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.562
cc_30 VNB N_B_c_486_n 0.00427147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B_c_487_n 0.0217914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_c_488_n 0.0100267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B_M1027_g 0.00516788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_c_490_n 0.0120411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_c_491_n 0.0220542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_M1024_g 0.00688156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_493_n 0.0279932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_B_c_494_n 0.0688041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_M1008_g 0.0207826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_B_c_496_n 0.00773258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_B_c_497_n 0.00953971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_B_c_498_n 0.00682074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_B_c_499_n 0.00586642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_367_119#_c_628_n 0.0195919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_367_119#_c_629_n 0.0256508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_367_119#_c_630_n 2.96981e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_367_119#_c_631_n 0.00464812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_367_119#_c_632_n 0.0256188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_367_119#_c_633_n 0.00160225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_367_119#_c_634_n 0.0272695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_367_119#_c_635_n 0.0113806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_367_119#_c_636_n 0.00911919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_367_119#_c_637_n 0.00245404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_367_119#_c_638_n 0.00574603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_367_119#_c_639_n 6.16417e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_367_119#_c_640_n 9.50626e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_367_119#_c_641_n 0.00322536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_367_119#_c_642_n 0.0116377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_367_119#_c_643_n 0.0382842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_367_119#_c_644_n 0.0209948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_367_119#_c_645_n 0.00240529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_359_367#_c_876_n 0.0174473f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.815
cc_63 VNB N_A_359_367#_c_877_n 0.0281288f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.51
cc_64 VNB N_A_359_367#_M1002_g 0.0214283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_359_367#_c_879_n 0.01868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_359_367#_c_880_n 0.0229056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_359_367#_c_881_n 0.00102522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_359_367#_c_882_n 0.0182089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_359_367#_c_883_n 0.00395558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_359_367#_c_884_n 0.0157147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_359_367#_c_885_n 0.00853546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_CI_M1026_g 0.00773458f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_73 VNB N_CI_c_1072_n 0.0151052f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.815
cc_74 VNB N_CI_c_1073_n 0.0193971f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.815
cc_75 VNB N_CI_M1023_g 0.00909649f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.51
cc_76 VNB N_CI_c_1075_n 0.0218467f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.675
cc_77 VNB CI 0.00480147f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.562
cc_78 VNB N_CI_c_1077_n 0.0128527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_CI_c_1078_n 0.05206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1571_367#_M1015_g 0.033158f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.51
cc_81 VNB N_A_1571_367#_c_1137_n 0.00148824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1571_367#_c_1138_n 0.00552488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1571_367#_c_1139_n 0.00237406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1571_367#_c_1140_n 0.0212339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1758_87#_c_1258_n 0.0226073f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.815
cc_86 VNB N_A_1758_87#_M1004_g 0.00935247f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.51
cc_87 VNB N_A_1758_87#_c_1260_n 0.00356084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1758_87#_c_1261_n 0.0268024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1758_87#_c_1262_n 0.00355032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1758_87#_c_1263_n 0.00598615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1758_87#_c_1264_n 0.00911686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1758_87#_c_1265_n 0.0109604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1758_87#_c_1266_n 0.0472862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VPWR_c_1360_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_247_367#_c_1458_n 0.00660112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_247_367#_c_1459_n 0.00281621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_247_367#_c_1460_n 0.00278504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_247_367#_c_1461_n 0.00354394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_247_367#_c_1462_n 0.00493883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1034_380#_c_1532_n 0.00809492f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.562
cc_101 VNB N_COUT_N_c_1583_n 0.00226751f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.675
cc_102 VNB N_COUT_N_c_1584_n 0.00502474f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.562
cc_103 VNB N_COUT_N_c_1585_n 0.00770569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1340_412#_c_1642_n 0.00731615f $X=-0.19 $Y=-0.245 $X2=0.55
+ $Y2=1.345
cc_105 VNB N_A_1340_412#_c_1643_n 0.0078f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.562
cc_106 VNB N_A_1708_411#_c_1687_n 0.00721334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1708_411#_c_1688_n 0.00281165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1708_411#_c_1689_n 0.0082397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_SUM_c_1747_n 0.0612071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1759_n 0.00969192f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.562
cc_111 VNB N_VGND_c_1760_n 0.00281759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1761_n 0.00765602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1762_n 0.00519418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1763_n 0.0631037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1764_n 0.00478085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1765_n 0.0945187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1766_n 0.0740887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1767_n 0.0202953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1768_n 0.625962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1769_n 0.0237735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1770_n 0.00370926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1771_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VPB N_A_M1030_g 0.0262075f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_124 VPB A 0.00581857f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_125 VPB N_A_c_218_n 0.00638322f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.51
cc_126 VPB N_A_33_367#_M1021_g 0.0235114f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.562
cc_127 VPB N_A_33_367#_c_269_n 0.0376809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_33_367#_c_262_n 0.00227648f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_33_367#_c_271_n 0.00781739f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_33_367#_c_264_n 0.013519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_33_367#_c_265_n 0.00391536f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_33_367#_c_274_n 5.71122e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_33_367#_c_267_n 0.0104355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_329_269#_M1022_g 0.0224792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_329_269#_M1000_g 0.0201662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_329_269#_c_388_n 0.00662768f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_329_269#_c_389_n 0.0104755f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_329_269#_c_383_n 0.00232731f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_B_M1013_g 0.0349445f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_140 VPB N_B_c_501_n 0.0631386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_B_c_502_n 0.0127165f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.51
cc_142 VPB N_B_M1018_g 0.0305044f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.675
cc_143 VPB N_B_c_504_n 0.0328344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_B_c_486_n 0.0761292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_B_M1027_g 0.0248748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_B_M1024_g 0.0291464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_B_c_496_n 0.0067025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_B_c_497_n 0.00749352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_B_c_510_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_367_119#_M1010_g 0.035928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_367_119#_M1028_g 0.0236644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_367_119#_c_648_n 0.0214923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_367_119#_c_630_n 0.00209001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_367_119#_c_650_n 7.99621e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_367_119#_c_651_n 0.00662403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_367_119#_c_631_n 0.00157915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_367_119#_c_632_n 0.0120623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_367_119#_c_633_n 0.00147179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_367_119#_c_634_n 7.58126e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_359_367#_M1014_g 0.0261183f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.675
cc_161 VPB N_A_359_367#_M1006_g 0.0218144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_359_367#_c_880_n 0.00805999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_359_367#_c_889_n 0.0382093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_359_367#_c_890_n 0.00196545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_359_367#_c_891_n 0.00598317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_359_367#_c_892_n 0.0186777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_359_367#_c_893_n 0.00964418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_359_367#_c_894_n 8.87072e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_359_367#_c_895_n 6.08529e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_359_367#_c_883_n 6.61181e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_359_367#_c_884_n 0.0332379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_359_367#_c_885_n 0.004459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_CI_M1026_g 0.0225826f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_174 VPB N_CI_M1023_g 0.0276084f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.51
cc_175 VPB N_A_1571_367#_c_1141_n 0.0214123f $X=-0.19 $Y=1.655 $X2=0.55
+ $Y2=1.675
cc_176 VPB N_A_1571_367#_c_1142_n 0.0106711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_1571_367#_c_1143_n 0.00920006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_1571_367#_c_1144_n 0.00465989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_1571_367#_c_1145_n 0.00825456f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_1571_367#_c_1138_n 0.00347804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_1571_367#_c_1147_n 0.00443044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_1571_367#_c_1148_n 0.0179501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_1571_367#_c_1149_n 0.00364849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1571_367#_c_1139_n 8.94042e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1571_367#_c_1140_n 0.0479724f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_1758_87#_M1004_g 0.0266659f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.51
cc_187 VPB N_A_1758_87#_c_1263_n 0.00774897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1361_n 0.00855338f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.562
cc_189 VPB N_VPWR_c_1362_n 0.013942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1363_n 0.00843541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1364_n 0.00589728f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1365_n 0.086913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1366_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1367_n 0.0708144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1368_n 0.0731695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1369_n 0.0191284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1360_n 0.147225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1371_n 0.0257748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1372_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1373_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_247_367#_c_1463_n 0.00484353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_247_367#_c_1464_n 0.0293475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_247_367#_c_1465_n 0.00406864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_247_367#_c_1459_n 0.0100052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_247_367#_c_1460_n 0.00254759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1034_380#_c_1533_n 0.0037499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_1034_380#_c_1534_n 0.0032424f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.51
cc_208 VPB N_A_1034_380#_c_1532_n 0.00482849f $X=-0.19 $Y=1.655 $X2=0.72
+ $Y2=1.562
cc_209 VPB N_COUT_N_c_1586_n 0.00624811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_COUT_N_c_1584_n 0.00783082f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.562
cc_211 VPB N_A_1340_412#_c_1644_n 0.00731095f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_1340_412#_c_1642_n 0.0033152f $X=-0.19 $Y=1.655 $X2=0.55
+ $Y2=1.345
cc_213 VPB N_A_1708_411#_c_1690_n 0.0292974f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.51
cc_214 VPB N_A_1708_411#_c_1689_n 0.00202312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_1708_411#_c_1692_n 0.00278628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_SUM_c_1747_n 0.0563215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 N_A_M1030_g N_A_33_367#_M1021_g 0.0222413f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_218 A N_A_33_367#_M1021_g 0.00108602f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A_c_219_n N_A_33_367#_c_257_n 0.00743123f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_220 N_A_c_219_n N_A_33_367#_c_258_n 0.0104317f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_221 N_A_M1030_g N_A_33_367#_c_269_n 0.00992971f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_222 A N_A_33_367#_c_281_n 0.0208083f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_223 N_A_c_218_n N_A_33_367#_c_281_n 0.00209843f $X=0.55 $Y=1.51 $X2=0 $Y2=0
cc_224 N_A_c_219_n N_A_33_367#_c_281_n 0.012438f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_225 N_A_c_219_n N_A_33_367#_c_259_n 0.00205798f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_226 A N_A_33_367#_c_263_n 0.00284321f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_227 N_A_c_218_n N_A_33_367#_c_263_n 0.00221147f $X=0.55 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A_c_219_n N_A_33_367#_c_263_n 7.42565e-19 $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_229 N_A_M1030_g N_A_33_367#_c_271_n 0.0023843f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_230 A N_A_33_367#_c_271_n 0.00224513f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_231 N_A_c_218_n N_A_33_367#_c_271_n 0.00115586f $X=0.55 $Y=1.51 $X2=0 $Y2=0
cc_232 N_A_M1030_g N_A_33_367#_c_264_n 0.00509804f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_233 A N_A_33_367#_c_264_n 0.0319932f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_234 N_A_c_218_n N_A_33_367#_c_264_n 0.00785554f $X=0.55 $Y=1.51 $X2=0 $Y2=0
cc_235 N_A_c_219_n N_A_33_367#_c_264_n 0.0042698f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_236 A N_A_33_367#_c_265_n 0.0244247f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_237 N_A_c_218_n N_A_33_367#_c_265_n 3.15306e-19 $X=0.55 $Y=1.51 $X2=0 $Y2=0
cc_238 N_A_c_219_n N_A_33_367#_c_266_n 0.00319923f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_239 A N_A_33_367#_c_267_n 0.00222366f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_240 N_A_c_218_n N_A_33_367#_c_267_n 0.0210693f $X=0.55 $Y=1.51 $X2=0 $Y2=0
cc_241 N_A_M1030_g N_VPWR_c_1361_n 0.0137703f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_242 A N_VPWR_c_1361_n 0.0126016f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_243 N_A_c_218_n N_VPWR_c_1361_n 3.57072e-19 $X=0.55 $Y=1.51 $X2=0 $Y2=0
cc_244 N_A_M1030_g N_VPWR_c_1360_n 0.0122769f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A_M1030_g N_VPWR_c_1371_n 0.00549284f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A_M1030_g N_A_247_367#_c_1468_n 6.70261e-19 $X=0.525 $Y=2.465 $X2=0
+ $Y2=0
cc_247 A N_A_247_367#_c_1460_n 0.00358624f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_248 N_A_c_219_n N_VGND_c_1759_n 0.00501106f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_249 N_A_c_219_n N_VGND_c_1768_n 0.00537853f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_250 N_A_c_219_n N_VGND_c_1769_n 0.00534051f $X=0.55 $Y=1.345 $X2=0 $Y2=0
cc_251 N_A_33_367#_M1021_g N_A_329_269#_M1022_g 0.0166399f $X=1.16 $Y=2.335
+ $X2=0 $Y2=0
cc_252 N_A_33_367#_c_257_n N_A_329_269#_M1029_g 0.0217243f $X=1.33 $Y=1.345
+ $X2=0 $Y2=0
cc_253 N_A_33_367#_c_259_n N_A_329_269#_M1029_g 9.95438e-19 $X=1.105 $Y=0.995
+ $X2=0 $Y2=0
cc_254 N_A_33_367#_c_260_n N_A_329_269#_M1029_g 0.017627f $X=2.455 $Y=0.35 $X2=0
+ $Y2=0
cc_255 N_A_33_367#_c_262_n N_A_329_269#_M1029_g 0.00178883f $X=2.54 $Y=0.78
+ $X2=0 $Y2=0
cc_256 N_A_33_367#_c_262_n N_A_329_269#_M1001_g 0.0169448f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_257 N_A_33_367#_c_262_n N_A_329_269#_M1000_g 0.00200213f $X=2.54 $Y=0.78
+ $X2=0 $Y2=0
cc_258 N_A_33_367#_c_274_n N_A_329_269#_M1000_g 0.0044104f $X=2.585 $Y=1.93
+ $X2=0 $Y2=0
cc_259 N_A_33_367#_c_267_n N_A_329_269#_c_378_n 0.0164405f $X=1.33 $Y=1.51 $X2=0
+ $Y2=0
cc_260 N_A_33_367#_c_262_n N_A_329_269#_c_379_n 0.00380296f $X=2.54 $Y=0.78
+ $X2=0 $Y2=0
cc_261 N_A_33_367#_c_274_n N_A_329_269#_c_379_n 8.09996e-19 $X=2.585 $Y=1.93
+ $X2=0 $Y2=0
cc_262 N_A_33_367#_c_260_n N_A_329_269#_c_381_n 0.00725032f $X=2.455 $Y=0.35
+ $X2=0 $Y2=0
cc_263 N_A_33_367#_c_262_n N_A_329_269#_c_381_n 0.00291784f $X=2.54 $Y=0.78
+ $X2=0 $Y2=0
cc_264 N_A_33_367#_c_260_n N_A_329_269#_c_382_n 0.0136575f $X=2.455 $Y=0.35
+ $X2=0 $Y2=0
cc_265 N_A_33_367#_c_262_n N_A_329_269#_c_382_n 0.00624329f $X=2.54 $Y=0.78
+ $X2=0 $Y2=0
cc_266 N_A_33_367#_c_260_n N_A_329_269#_c_385_n 0.0154834f $X=2.455 $Y=0.35
+ $X2=0 $Y2=0
cc_267 N_A_33_367#_c_260_n N_B_M1005_g 0.00293673f $X=2.455 $Y=0.35 $X2=0 $Y2=0
cc_268 N_A_33_367#_c_262_n N_B_M1005_g 0.00674406f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_269 N_A_33_367#_c_274_n N_B_M1013_g 0.00439588f $X=2.585 $Y=1.93 $X2=0 $Y2=0
cc_270 N_A_33_367#_c_262_n N_B_c_496_n 0.00295386f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_271 N_A_33_367#_M1021_g N_A_367_119#_c_630_n 3.16014e-19 $X=1.16 $Y=2.335
+ $X2=0 $Y2=0
cc_272 N_A_33_367#_c_262_n N_A_367_119#_c_630_n 0.005978f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_273 N_A_33_367#_c_274_n N_A_367_119#_c_630_n 3.18774e-19 $X=2.585 $Y=1.93
+ $X2=0 $Y2=0
cc_274 N_A_33_367#_M1013_d N_A_367_119#_c_651_n 0.00181172f $X=2.445 $Y=1.795
+ $X2=0 $Y2=0
cc_275 N_A_33_367#_c_267_n N_A_367_119#_c_635_n 2.28079e-19 $X=1.33 $Y=1.51
+ $X2=0 $Y2=0
cc_276 N_A_33_367#_M1005_d N_A_367_119#_c_636_n 0.00234379f $X=2.38 $Y=0.635
+ $X2=0 $Y2=0
cc_277 N_A_33_367#_c_260_n N_A_367_119#_c_636_n 0.00502149f $X=2.455 $Y=0.35
+ $X2=0 $Y2=0
cc_278 N_A_33_367#_c_262_n N_A_367_119#_c_636_n 0.0301483f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_279 N_A_33_367#_c_260_n N_A_367_119#_c_664_n 0.00235342f $X=2.455 $Y=0.35
+ $X2=0 $Y2=0
cc_280 N_A_33_367#_c_262_n N_A_367_119#_c_664_n 0.00232062f $X=2.54 $Y=0.78
+ $X2=0 $Y2=0
cc_281 N_A_33_367#_c_260_n N_A_367_119#_c_645_n 0.0272733f $X=2.455 $Y=0.35
+ $X2=0 $Y2=0
cc_282 N_A_33_367#_c_262_n N_A_367_119#_c_645_n 0.0694317f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_283 N_A_33_367#_c_274_n N_A_359_367#_c_890_n 0.00928848f $X=2.585 $Y=1.93
+ $X2=0 $Y2=0
cc_284 N_A_33_367#_M1013_d N_A_359_367#_c_900_n 0.00350618f $X=2.445 $Y=1.795
+ $X2=0 $Y2=0
cc_285 N_A_33_367#_c_274_n N_A_359_367#_c_900_n 0.0160901f $X=2.585 $Y=1.93
+ $X2=0 $Y2=0
cc_286 N_A_33_367#_c_274_n N_A_359_367#_c_902_n 6.10639e-19 $X=2.585 $Y=1.93
+ $X2=0 $Y2=0
cc_287 N_A_33_367#_c_262_n N_A_359_367#_c_885_n 0.0650646f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_288 N_A_33_367#_c_274_n N_A_359_367#_c_885_n 0.0094893f $X=2.585 $Y=1.93
+ $X2=0 $Y2=0
cc_289 N_A_33_367#_M1021_g N_VPWR_c_1361_n 0.00997545f $X=1.16 $Y=2.335 $X2=0
+ $Y2=0
cc_290 N_A_33_367#_c_267_n N_VPWR_c_1361_n 0.00231844f $X=1.33 $Y=1.51 $X2=0
+ $Y2=0
cc_291 N_A_33_367#_M1021_g N_VPWR_c_1365_n 0.00421151f $X=1.16 $Y=2.335 $X2=0
+ $Y2=0
cc_292 N_A_33_367#_M1030_s N_VPWR_c_1360_n 0.0023218f $X=0.165 $Y=1.835 $X2=0
+ $Y2=0
cc_293 N_A_33_367#_M1021_g N_VPWR_c_1360_n 0.00422397f $X=1.16 $Y=2.335 $X2=0
+ $Y2=0
cc_294 N_A_33_367#_c_269_n N_VPWR_c_1360_n 0.0146362f $X=0.31 $Y=2.9 $X2=0 $Y2=0
cc_295 N_A_33_367#_c_269_n N_VPWR_c_1371_n 0.0234664f $X=0.31 $Y=2.9 $X2=0 $Y2=0
cc_296 N_A_33_367#_M1021_g N_A_247_367#_c_1468_n 0.00406882f $X=1.16 $Y=2.335
+ $X2=0 $Y2=0
cc_297 N_A_33_367#_c_267_n N_A_247_367#_c_1468_n 0.00501967f $X=1.33 $Y=1.51
+ $X2=0 $Y2=0
cc_298 N_A_33_367#_M1021_g N_A_247_367#_c_1463_n 0.0151207f $X=1.16 $Y=2.335
+ $X2=0 $Y2=0
cc_299 N_A_33_367#_c_257_n N_A_247_367#_c_1473_n 0.00686873f $X=1.33 $Y=1.345
+ $X2=0 $Y2=0
cc_300 N_A_33_367#_c_259_n N_A_247_367#_c_1473_n 0.0268722f $X=1.105 $Y=0.995
+ $X2=0 $Y2=0
cc_301 N_A_33_367#_c_260_n N_A_247_367#_c_1473_n 0.0204209f $X=2.455 $Y=0.35
+ $X2=0 $Y2=0
cc_302 N_A_33_367#_c_351_p N_A_247_367#_c_1473_n 0.0134221f $X=1.105 $Y=1.08
+ $X2=0 $Y2=0
cc_303 N_A_33_367#_M1021_g N_A_247_367#_c_1465_n 0.00292293f $X=1.16 $Y=2.335
+ $X2=0 $Y2=0
cc_304 N_A_33_367#_M1021_g N_A_247_367#_c_1460_n 0.00283453f $X=1.16 $Y=2.335
+ $X2=0 $Y2=0
cc_305 N_A_33_367#_c_257_n N_A_247_367#_c_1460_n 0.00202048f $X=1.33 $Y=1.345
+ $X2=0 $Y2=0
cc_306 N_A_33_367#_c_265_n N_A_247_367#_c_1460_n 0.0170171f $X=1.09 $Y=1.51
+ $X2=0 $Y2=0
cc_307 N_A_33_367#_c_267_n N_A_247_367#_c_1460_n 0.00841818f $X=1.33 $Y=1.51
+ $X2=0 $Y2=0
cc_308 N_A_33_367#_c_257_n N_A_247_367#_c_1461_n 0.00332093f $X=1.33 $Y=1.345
+ $X2=0 $Y2=0
cc_309 N_A_33_367#_c_266_n N_A_247_367#_c_1461_n 0.0170171f $X=1.087 $Y=1.345
+ $X2=0 $Y2=0
cc_310 N_A_33_367#_c_281_n N_VGND_M1025_d 0.0176352f $X=1.02 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_311 N_A_33_367#_c_259_n N_VGND_M1025_d 0.0116406f $X=1.105 $Y=0.995 $X2=-0.19
+ $Y2=-0.245
cc_312 N_A_33_367#_c_266_n N_VGND_M1025_d 0.00155034f $X=1.087 $Y=1.345
+ $X2=-0.19 $Y2=-0.245
cc_313 N_A_33_367#_c_351_p N_VGND_M1025_d 0.00307338f $X=1.105 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_314 N_A_33_367#_c_258_n N_VGND_c_1759_n 0.0169279f $X=0.325 $Y=0.54 $X2=0
+ $Y2=0
cc_315 N_A_33_367#_c_281_n N_VGND_c_1759_n 0.0130182f $X=1.02 $Y=1.08 $X2=0
+ $Y2=0
cc_316 N_A_33_367#_c_259_n N_VGND_c_1759_n 0.0266331f $X=1.105 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A_33_367#_c_261_n N_VGND_c_1759_n 0.0137332f $X=1.19 $Y=0.35 $X2=0
+ $Y2=0
cc_318 N_A_33_367#_c_260_n N_VGND_c_1765_n 0.0921662f $X=2.455 $Y=0.35 $X2=0
+ $Y2=0
cc_319 N_A_33_367#_c_261_n N_VGND_c_1765_n 0.0114622f $X=1.19 $Y=0.35 $X2=0
+ $Y2=0
cc_320 N_A_33_367#_c_258_n N_VGND_c_1768_n 0.0144552f $X=0.325 $Y=0.54 $X2=0
+ $Y2=0
cc_321 N_A_33_367#_c_260_n N_VGND_c_1768_n 0.0525672f $X=2.455 $Y=0.35 $X2=0
+ $Y2=0
cc_322 N_A_33_367#_c_261_n N_VGND_c_1768_n 0.00657784f $X=1.19 $Y=0.35 $X2=0
+ $Y2=0
cc_323 N_A_33_367#_c_258_n N_VGND_c_1769_n 0.016068f $X=0.325 $Y=0.54 $X2=0
+ $Y2=0
cc_324 N_A_329_269#_M1022_g N_B_M1005_g 0.00448111f $X=1.72 $Y=2.255 $X2=0 $Y2=0
cc_325 N_A_329_269#_M1029_g N_B_M1005_g 0.0165002f $X=1.76 $Y=0.915 $X2=0 $Y2=0
cc_326 N_A_329_269#_c_381_n N_B_M1005_g 0.0138689f $X=3.05 $Y=0.36 $X2=0 $Y2=0
cc_327 N_A_329_269#_c_385_n N_B_M1005_g 0.00737859f $X=2.685 $Y=0.32 $X2=0 $Y2=0
cc_328 N_A_329_269#_M1022_g N_B_M1013_g 0.0182932f $X=1.72 $Y=2.255 $X2=0 $Y2=0
cc_329 N_A_329_269#_M1000_g N_B_c_501_n 0.00828781f $X=2.8 $Y=2.215 $X2=0 $Y2=0
cc_330 N_A_329_269#_M1001_g N_B_M1031_g 0.0121167f $X=2.76 $Y=0.955 $X2=0 $Y2=0
cc_331 N_A_329_269#_c_379_n N_B_M1031_g 0.0017596f $X=2.78 $Y=1.535 $X2=0 $Y2=0
cc_332 N_A_329_269#_c_380_n N_B_M1031_g 0.00481228f $X=4.095 $Y=0.35 $X2=0 $Y2=0
cc_333 N_A_329_269#_c_381_n N_B_M1031_g 0.00102597f $X=3.05 $Y=0.36 $X2=0 $Y2=0
cc_334 N_A_329_269#_c_384_n N_B_M1031_g 0.00457304f $X=4.38 $Y=0.35 $X2=0 $Y2=0
cc_335 N_A_329_269#_c_389_n N_B_c_504_n 0.00629963f $X=4.22 $Y=2.9 $X2=0 $Y2=0
cc_336 N_A_329_269#_c_388_n N_B_c_486_n 0.00629963f $X=4.22 $Y=1.94 $X2=0 $Y2=0
cc_337 N_A_329_269#_c_383_n N_B_c_486_n 0.00227357f $X=4.22 $Y=1.775 $X2=0 $Y2=0
cc_338 N_A_329_269#_c_383_n N_B_c_487_n 0.0145516f $X=4.22 $Y=1.775 $X2=0 $Y2=0
cc_339 N_A_329_269#_c_384_n N_B_c_487_n 0.00692157f $X=4.38 $Y=0.35 $X2=0 $Y2=0
cc_340 N_A_329_269#_c_388_n N_B_M1027_g 0.00313969f $X=4.22 $Y=1.94 $X2=0 $Y2=0
cc_341 N_A_329_269#_c_389_n N_B_M1027_g 0.0139784f $X=4.22 $Y=2.9 $X2=0 $Y2=0
cc_342 N_A_329_269#_c_383_n N_B_M1027_g 0.00459363f $X=4.22 $Y=1.775 $X2=0 $Y2=0
cc_343 N_A_329_269#_c_383_n N_B_c_491_n 0.00407442f $X=4.22 $Y=1.775 $X2=0 $Y2=0
cc_344 N_A_329_269#_c_384_n N_B_c_491_n 0.0139065f $X=4.38 $Y=0.35 $X2=0 $Y2=0
cc_345 N_A_329_269#_M1000_g N_B_c_496_n 0.0394161f $X=2.8 $Y=2.215 $X2=0 $Y2=0
cc_346 N_A_329_269#_M1000_g N_B_c_497_n 0.0235818f $X=2.8 $Y=2.215 $X2=0 $Y2=0
cc_347 N_A_329_269#_c_384_n N_B_c_498_n 0.00108905f $X=4.38 $Y=0.35 $X2=0 $Y2=0
cc_348 N_A_329_269#_c_383_n N_B_c_499_n 0.0267174f $X=4.22 $Y=1.775 $X2=0 $Y2=0
cc_349 N_A_329_269#_c_384_n N_B_c_499_n 0.0164739f $X=4.38 $Y=0.35 $X2=0 $Y2=0
cc_350 N_A_329_269#_M1022_g N_A_367_119#_c_630_n 0.0229257f $X=1.72 $Y=2.255
+ $X2=0 $Y2=0
cc_351 N_A_329_269#_M1022_g N_A_367_119#_c_650_n 0.00593689f $X=1.72 $Y=2.255
+ $X2=0 $Y2=0
cc_352 N_A_329_269#_M1000_g N_A_367_119#_c_651_n 0.00992149f $X=2.8 $Y=2.215
+ $X2=0 $Y2=0
cc_353 N_A_329_269#_M1022_g N_A_367_119#_c_635_n 0.00265966f $X=1.72 $Y=2.255
+ $X2=0 $Y2=0
cc_354 N_A_329_269#_c_378_n N_A_367_119#_c_635_n 0.00954111f $X=1.74 $Y=1.495
+ $X2=0 $Y2=0
cc_355 N_A_329_269#_c_379_n N_A_367_119#_c_635_n 2.47213e-19 $X=2.78 $Y=1.535
+ $X2=0 $Y2=0
cc_356 N_A_329_269#_M1011_s N_A_367_119#_c_636_n 0.00248718f $X=4.355 $Y=0.25
+ $X2=0 $Y2=0
cc_357 N_A_329_269#_M1001_g N_A_367_119#_c_636_n 0.0124054f $X=2.76 $Y=0.955
+ $X2=0 $Y2=0
cc_358 N_A_329_269#_c_379_n N_A_367_119#_c_636_n 9.79098e-19 $X=2.78 $Y=1.535
+ $X2=0 $Y2=0
cc_359 N_A_329_269#_c_380_n N_A_367_119#_c_636_n 0.0165045f $X=4.095 $Y=0.35
+ $X2=0 $Y2=0
cc_360 N_A_329_269#_c_381_n N_A_367_119#_c_636_n 0.00219154f $X=3.05 $Y=0.36
+ $X2=0 $Y2=0
cc_361 N_A_329_269#_c_382_n N_A_367_119#_c_636_n 0.00315928f $X=3.215 $Y=0.395
+ $X2=0 $Y2=0
cc_362 N_A_329_269#_c_384_n N_A_367_119#_c_636_n 0.0532457f $X=4.38 $Y=0.35
+ $X2=0 $Y2=0
cc_363 N_A_329_269#_M1029_g N_A_367_119#_c_645_n 0.00567293f $X=1.76 $Y=0.915
+ $X2=0 $Y2=0
cc_364 N_A_329_269#_M1001_g N_A_367_119#_c_645_n 2.47213e-19 $X=2.76 $Y=0.955
+ $X2=0 $Y2=0
cc_365 N_A_329_269#_M1022_g N_A_359_367#_c_890_n 0.00125332f $X=1.72 $Y=2.255
+ $X2=0 $Y2=0
cc_366 N_A_329_269#_M1000_g N_A_359_367#_c_900_n 0.0148784f $X=2.8 $Y=2.215
+ $X2=0 $Y2=0
cc_367 N_A_329_269#_M1022_g N_A_359_367#_c_907_n 6.33471e-19 $X=1.72 $Y=2.255
+ $X2=0 $Y2=0
cc_368 N_A_329_269#_c_389_n N_A_359_367#_c_892_n 0.0377876f $X=4.22 $Y=2.9 $X2=0
+ $Y2=0
cc_369 N_A_329_269#_M1001_g N_A_359_367#_c_885_n 0.0074109f $X=2.76 $Y=0.955
+ $X2=0 $Y2=0
cc_370 N_A_329_269#_c_379_n N_A_359_367#_c_885_n 0.00723923f $X=2.78 $Y=1.535
+ $X2=0 $Y2=0
cc_371 N_A_329_269#_c_380_n N_A_359_367#_c_885_n 0.00203066f $X=4.095 $Y=0.35
+ $X2=0 $Y2=0
cc_372 N_A_329_269#_c_381_n N_A_359_367#_c_885_n 0.00687214f $X=3.05 $Y=0.36
+ $X2=0 $Y2=0
cc_373 N_A_329_269#_c_382_n N_A_359_367#_c_885_n 0.0195652f $X=3.215 $Y=0.395
+ $X2=0 $Y2=0
cc_374 N_A_329_269#_c_388_n N_VPWR_c_1362_n 0.0489682f $X=4.22 $Y=1.94 $X2=0
+ $Y2=0
cc_375 N_A_329_269#_c_389_n N_VPWR_c_1365_n 0.0220321f $X=4.22 $Y=2.9 $X2=0
+ $Y2=0
cc_376 N_A_329_269#_c_389_n N_VPWR_c_1360_n 0.0125808f $X=4.22 $Y=2.9 $X2=0
+ $Y2=0
cc_377 N_A_329_269#_M1022_g N_A_247_367#_c_1468_n 0.00658209f $X=1.72 $Y=2.255
+ $X2=0 $Y2=0
cc_378 N_A_329_269#_M1029_g N_A_247_367#_c_1473_n 0.00638777f $X=1.76 $Y=0.915
+ $X2=0 $Y2=0
cc_379 N_A_329_269#_M1022_g N_A_247_367#_c_1464_n 0.00557622f $X=1.72 $Y=2.255
+ $X2=0 $Y2=0
cc_380 N_A_329_269#_M1000_g N_A_247_367#_c_1464_n 0.00105106f $X=2.8 $Y=2.215
+ $X2=0 $Y2=0
cc_381 N_A_329_269#_c_389_n N_A_247_367#_c_1464_n 0.0111807f $X=4.22 $Y=2.9
+ $X2=0 $Y2=0
cc_382 N_A_329_269#_M1001_g N_A_247_367#_c_1458_n 5.99983e-19 $X=2.76 $Y=0.955
+ $X2=0 $Y2=0
cc_383 N_A_329_269#_c_380_n N_A_247_367#_c_1458_n 0.0305372f $X=4.095 $Y=0.35
+ $X2=0 $Y2=0
cc_384 N_A_329_269#_c_384_n N_A_247_367#_c_1458_n 0.0263557f $X=4.38 $Y=0.35
+ $X2=0 $Y2=0
cc_385 N_A_329_269#_M1000_g N_A_247_367#_c_1459_n 0.00147504f $X=2.8 $Y=2.215
+ $X2=0 $Y2=0
cc_386 N_A_329_269#_c_388_n N_A_247_367#_c_1459_n 0.0691184f $X=4.22 $Y=1.94
+ $X2=0 $Y2=0
cc_387 N_A_329_269#_c_383_n N_A_247_367#_c_1459_n 0.0258892f $X=4.22 $Y=1.775
+ $X2=0 $Y2=0
cc_388 N_A_329_269#_M1029_g N_A_247_367#_c_1460_n 8.62136e-19 $X=1.76 $Y=0.915
+ $X2=0 $Y2=0
cc_389 N_A_329_269#_c_378_n N_A_247_367#_c_1460_n 0.00658209f $X=1.74 $Y=1.495
+ $X2=0 $Y2=0
cc_390 N_A_329_269#_M1029_g N_A_247_367#_c_1461_n 0.00437369f $X=1.76 $Y=0.915
+ $X2=0 $Y2=0
cc_391 N_A_329_269#_c_383_n N_A_247_367#_c_1462_n 0.0263557f $X=4.22 $Y=1.775
+ $X2=0 $Y2=0
cc_392 N_A_329_269#_c_384_n N_VGND_c_1760_n 0.0271363f $X=4.38 $Y=0.35 $X2=0
+ $Y2=0
cc_393 N_A_329_269#_c_375_n N_VGND_c_1765_n 0.0356658f $X=1.835 $Y=0.19 $X2=0
+ $Y2=0
cc_394 N_A_329_269#_c_382_n N_VGND_c_1765_n 0.0729397f $X=3.215 $Y=0.395 $X2=0
+ $Y2=0
cc_395 N_A_329_269#_c_384_n N_VGND_c_1765_n 0.0378443f $X=4.38 $Y=0.35 $X2=0
+ $Y2=0
cc_396 N_A_329_269#_c_375_n N_VGND_c_1768_n 0.00589247f $X=1.835 $Y=0.19 $X2=0
+ $Y2=0
cc_397 N_A_329_269#_c_381_n N_VGND_c_1768_n 0.0213147f $X=3.05 $Y=0.36 $X2=0
+ $Y2=0
cc_398 N_A_329_269#_c_382_n N_VGND_c_1768_n 0.0438219f $X=3.215 $Y=0.395 $X2=0
+ $Y2=0
cc_399 N_A_329_269#_c_384_n N_VGND_c_1768_n 0.0219723f $X=4.38 $Y=0.35 $X2=0
+ $Y2=0
cc_400 N_A_329_269#_c_385_n N_VGND_c_1768_n 0.0200988f $X=2.685 $Y=0.32 $X2=0
+ $Y2=0
cc_401 N_B_M1024_g N_A_367_119#_M1010_g 0.0123324f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_402 N_B_M1013_g N_A_367_119#_c_630_n 0.00471267f $X=2.37 $Y=2.215 $X2=0 $Y2=0
cc_403 N_B_c_496_n N_A_367_119#_c_630_n 8.4439e-19 $X=2.337 $Y=1.685 $X2=0 $Y2=0
cc_404 N_B_M1013_g N_A_367_119#_c_651_n 0.0114839f $X=2.37 $Y=2.215 $X2=0 $Y2=0
cc_405 N_B_c_501_n N_A_367_119#_c_651_n 0.00323622f $X=3.35 $Y=3.08 $X2=0 $Y2=0
cc_406 N_B_M1018_g N_A_367_119#_c_651_n 0.00178081f $X=3.425 $Y=2.215 $X2=0
+ $Y2=0
cc_407 N_B_c_493_n N_A_367_119#_c_631_n 0.00662549f $X=5.67 $Y=1.095 $X2=0 $Y2=0
cc_408 N_B_c_494_n N_A_367_119#_c_631_n 9.93761e-19 $X=5.38 $Y=1.095 $X2=0 $Y2=0
cc_409 N_B_c_493_n N_A_367_119#_c_632_n 0.013294f $X=5.67 $Y=1.095 $X2=0 $Y2=0
cc_410 N_B_c_494_n N_A_367_119#_c_632_n 0.0123324f $X=5.38 $Y=1.095 $X2=0 $Y2=0
cc_411 N_B_M1005_g N_A_367_119#_c_635_n 0.00325199f $X=2.305 $Y=0.955 $X2=0
+ $Y2=0
cc_412 N_B_c_496_n N_A_367_119#_c_635_n 0.00218158f $X=2.337 $Y=1.685 $X2=0
+ $Y2=0
cc_413 N_B_M1005_g N_A_367_119#_c_636_n 0.00378924f $X=2.305 $Y=0.955 $X2=0
+ $Y2=0
cc_414 N_B_M1031_g N_A_367_119#_c_636_n 0.0026373f $X=3.53 $Y=0.955 $X2=0 $Y2=0
cc_415 N_B_c_488_n N_A_367_119#_c_636_n 0.00457893f $X=4.005 $Y=1.455 $X2=0
+ $Y2=0
cc_416 N_B_c_491_n N_A_367_119#_c_636_n 0.00847661f $X=4.795 $Y=1.2 $X2=0 $Y2=0
cc_417 N_B_c_494_n N_A_367_119#_c_636_n 0.00949635f $X=5.38 $Y=1.095 $X2=0 $Y2=0
cc_418 N_B_c_496_n N_A_367_119#_c_636_n 0.00144944f $X=2.337 $Y=1.685 $X2=0
+ $Y2=0
cc_419 N_B_c_497_n N_A_367_119#_c_636_n 0.00235503f $X=3.53 $Y=1.61 $X2=0 $Y2=0
cc_420 N_B_c_499_n N_A_367_119#_c_636_n 0.0111787f $X=4.885 $Y=1.365 $X2=0 $Y2=0
cc_421 N_B_M1005_g N_A_367_119#_c_664_n 0.00238571f $X=2.305 $Y=0.955 $X2=0
+ $Y2=0
cc_422 N_B_c_493_n N_A_367_119#_c_641_n 0.00154781f $X=5.67 $Y=1.095 $X2=0 $Y2=0
cc_423 N_B_M1008_g N_A_367_119#_c_641_n 0.0104215f $X=5.745 $Y=0.57 $X2=0 $Y2=0
cc_424 N_B_M1005_g N_A_367_119#_c_645_n 0.0110308f $X=2.305 $Y=0.955 $X2=0 $Y2=0
cc_425 N_B_M1008_g N_A_359_367#_c_876_n 0.0145034f $X=5.745 $Y=0.57 $X2=0 $Y2=0
cc_426 N_B_c_493_n N_A_359_367#_c_877_n 4.3846e-19 $X=5.67 $Y=1.095 $X2=0 $Y2=0
cc_427 N_B_c_493_n N_A_359_367#_c_879_n 0.0145034f $X=5.67 $Y=1.095 $X2=0 $Y2=0
cc_428 N_B_M1013_g N_A_359_367#_c_890_n 7.412e-19 $X=2.37 $Y=2.215 $X2=0 $Y2=0
cc_429 N_B_c_496_n N_A_359_367#_c_890_n 2.71532e-19 $X=2.337 $Y=1.685 $X2=0
+ $Y2=0
cc_430 N_B_M1013_g N_A_359_367#_c_900_n 0.0135564f $X=2.37 $Y=2.215 $X2=0 $Y2=0
cc_431 N_B_M1018_g N_A_359_367#_c_900_n 0.00180201f $X=3.425 $Y=2.215 $X2=0
+ $Y2=0
cc_432 N_B_M1018_g N_A_359_367#_c_892_n 0.0109167f $X=3.425 $Y=2.215 $X2=0 $Y2=0
cc_433 N_B_c_486_n N_A_359_367#_c_892_n 0.0147591f $X=3.93 $Y=3.005 $X2=0 $Y2=0
cc_434 N_B_M1027_g N_A_359_367#_c_892_n 0.00986421f $X=4.435 $Y=2.425 $X2=0
+ $Y2=0
cc_435 N_B_M1024_g N_A_359_367#_c_892_n 0.0110341f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_436 N_B_c_494_n N_A_359_367#_c_892_n 7.43687e-19 $X=5.38 $Y=1.095 $X2=0 $Y2=0
cc_437 N_B_c_499_n N_A_359_367#_c_892_n 0.0106757f $X=4.885 $Y=1.365 $X2=0 $Y2=0
cc_438 N_B_M1018_g N_A_359_367#_c_902_n 0.00158129f $X=3.425 $Y=2.215 $X2=0
+ $Y2=0
cc_439 N_B_M1031_g N_A_359_367#_c_885_n 0.00731358f $X=3.53 $Y=0.955 $X2=0 $Y2=0
cc_440 N_B_c_497_n N_A_359_367#_c_885_n 0.00628956f $X=3.53 $Y=1.61 $X2=0 $Y2=0
cc_441 N_B_M1027_g N_VPWR_c_1362_n 0.013862f $X=4.435 $Y=2.425 $X2=0 $Y2=0
cc_442 N_B_c_490_n N_VPWR_c_1362_n 0.00673699f $X=4.72 $Y=1.455 $X2=0 $Y2=0
cc_443 N_B_M1024_g N_VPWR_c_1362_n 0.0144448f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_444 N_B_c_499_n N_VPWR_c_1362_n 0.0194035f $X=4.885 $Y=1.365 $X2=0 $Y2=0
cc_445 N_B_c_502_n N_VPWR_c_1365_n 0.035636f $X=2.445 $Y=3.08 $X2=0 $Y2=0
cc_446 N_B_M1027_g N_VPWR_c_1365_n 0.00511657f $X=4.435 $Y=2.425 $X2=0 $Y2=0
cc_447 N_B_M1024_g N_VPWR_c_1367_n 0.00510764f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_448 N_B_c_501_n N_VPWR_c_1360_n 0.0218378f $X=3.35 $Y=3.08 $X2=0 $Y2=0
cc_449 N_B_c_502_n N_VPWR_c_1360_n 0.00495874f $X=2.445 $Y=3.08 $X2=0 $Y2=0
cc_450 N_B_c_504_n N_VPWR_c_1360_n 0.0203726f $X=3.855 $Y=3.08 $X2=0 $Y2=0
cc_451 N_B_M1027_g N_VPWR_c_1360_n 0.0109276f $X=4.435 $Y=2.425 $X2=0 $Y2=0
cc_452 N_B_M1024_g N_VPWR_c_1360_n 0.00526787f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_453 N_B_c_510_n N_VPWR_c_1360_n 0.00379035f $X=3.425 $Y=3.08 $X2=0 $Y2=0
cc_454 N_B_M1013_g N_A_247_367#_c_1464_n 0.00884348f $X=2.37 $Y=2.215 $X2=0
+ $Y2=0
cc_455 N_B_c_501_n N_A_247_367#_c_1464_n 0.0219439f $X=3.35 $Y=3.08 $X2=0 $Y2=0
cc_456 N_B_c_502_n N_A_247_367#_c_1464_n 0.00342282f $X=2.445 $Y=3.08 $X2=0
+ $Y2=0
cc_457 N_B_M1018_g N_A_247_367#_c_1464_n 0.010925f $X=3.425 $Y=2.215 $X2=0 $Y2=0
cc_458 N_B_c_504_n N_A_247_367#_c_1464_n 0.00886255f $X=3.855 $Y=3.08 $X2=0
+ $Y2=0
cc_459 N_B_c_486_n N_A_247_367#_c_1464_n 0.00117892f $X=3.93 $Y=3.005 $X2=0
+ $Y2=0
cc_460 N_B_c_510_n N_A_247_367#_c_1464_n 0.00192788f $X=3.425 $Y=3.08 $X2=0
+ $Y2=0
cc_461 N_B_M1031_g N_A_247_367#_c_1458_n 0.0105199f $X=3.53 $Y=0.955 $X2=0 $Y2=0
cc_462 N_B_M1018_g N_A_247_367#_c_1459_n 0.02604f $X=3.425 $Y=2.215 $X2=0 $Y2=0
cc_463 N_B_M1031_g N_A_247_367#_c_1459_n 0.00712484f $X=3.53 $Y=0.955 $X2=0
+ $Y2=0
cc_464 N_B_c_488_n N_A_247_367#_c_1459_n 0.0147682f $X=4.005 $Y=1.455 $X2=0
+ $Y2=0
cc_465 N_B_c_497_n N_A_247_367#_c_1459_n 0.00702929f $X=3.53 $Y=1.61 $X2=0 $Y2=0
cc_466 N_B_M1031_g N_A_247_367#_c_1462_n 0.00439063f $X=3.53 $Y=0.955 $X2=0
+ $Y2=0
cc_467 N_B_c_488_n N_A_247_367#_c_1462_n 0.00284747f $X=4.005 $Y=1.455 $X2=0
+ $Y2=0
cc_468 N_B_M1024_g N_A_1034_380#_c_1533_n 0.00320884f $X=5.095 $Y=2.4 $X2=0
+ $Y2=0
cc_469 N_B_c_494_n N_A_1034_380#_c_1533_n 0.0039803f $X=5.38 $Y=1.095 $X2=0
+ $Y2=0
cc_470 N_B_M1024_g N_A_1034_380#_c_1534_n 0.0110895f $X=5.095 $Y=2.4 $X2=0 $Y2=0
cc_471 N_B_c_493_n N_A_1034_380#_c_1539_n 0.00429055f $X=5.67 $Y=1.095 $X2=0
+ $Y2=0
cc_472 N_B_M1008_g N_A_1034_380#_c_1539_n 0.009826f $X=5.745 $Y=0.57 $X2=0 $Y2=0
cc_473 N_B_c_491_n N_A_1034_380#_c_1541_n 4.57139e-19 $X=4.795 $Y=1.2 $X2=0
+ $Y2=0
cc_474 N_B_c_491_n N_A_1034_380#_c_1532_n 0.00137219f $X=4.795 $Y=1.2 $X2=0
+ $Y2=0
cc_475 N_B_c_493_n N_A_1034_380#_c_1532_n 0.00773397f $X=5.67 $Y=1.095 $X2=0
+ $Y2=0
cc_476 N_B_c_494_n N_A_1034_380#_c_1532_n 0.0235011f $X=5.38 $Y=1.095 $X2=0
+ $Y2=0
cc_477 N_B_M1008_g N_A_1034_380#_c_1532_n 0.00735521f $X=5.745 $Y=0.57 $X2=0
+ $Y2=0
cc_478 N_B_c_499_n N_A_1034_380#_c_1532_n 0.019731f $X=4.885 $Y=1.365 $X2=0
+ $Y2=0
cc_479 N_B_M1008_g N_A_1034_380#_c_1547_n 0.0099138f $X=5.745 $Y=0.57 $X2=0
+ $Y2=0
cc_480 N_B_c_491_n N_VGND_c_1760_n 0.0151743f $X=4.795 $Y=1.2 $X2=0 $Y2=0
cc_481 N_B_c_494_n N_VGND_c_1760_n 0.00322107f $X=5.38 $Y=1.095 $X2=0 $Y2=0
cc_482 N_B_M1008_g N_VGND_c_1760_n 0.00761348f $X=5.745 $Y=0.57 $X2=0 $Y2=0
cc_483 N_B_c_499_n N_VGND_c_1760_n 0.012747f $X=4.885 $Y=1.365 $X2=0 $Y2=0
cc_484 N_B_c_491_n N_VGND_c_1765_n 0.00473366f $X=4.795 $Y=1.2 $X2=0 $Y2=0
cc_485 N_B_M1008_g N_VGND_c_1766_n 0.003811f $X=5.745 $Y=0.57 $X2=0 $Y2=0
cc_486 N_B_c_491_n N_VGND_c_1768_n 0.00952851f $X=4.795 $Y=1.2 $X2=0 $Y2=0
cc_487 N_B_M1008_g N_VGND_c_1768_n 0.00670557f $X=5.745 $Y=0.57 $X2=0 $Y2=0
cc_488 N_A_367_119#_c_636_n N_A_359_367#_M1001_d 0.0115668f $X=5.855 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_489 N_A_367_119#_c_630_n N_A_359_367#_M1022_d 0.0074759f $X=1.805 $Y=2.545
+ $X2=0 $Y2=0
cc_490 N_A_367_119#_c_651_n N_A_359_367#_M1022_d 0.00949284f $X=3.095 $Y=2.63
+ $X2=0 $Y2=0
cc_491 N_A_367_119#_c_637_n N_A_359_367#_c_876_n 0.00658809f $X=6.815 $Y=0.925
+ $X2=0 $Y2=0
cc_492 N_A_367_119#_c_638_n N_A_359_367#_c_876_n 0.00149697f $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_493 N_A_367_119#_c_641_n N_A_359_367#_c_876_n 0.00355434f $X=6 $Y=0.925 $X2=0
+ $Y2=0
cc_494 N_A_367_119#_c_644_n N_A_359_367#_c_876_n 0.0134216f $X=6.82 $Y=1 $X2=0
+ $Y2=0
cc_495 N_A_367_119#_c_631_n N_A_359_367#_c_877_n 0.00176255f $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_496 N_A_367_119#_c_632_n N_A_359_367#_c_877_n 0.00947573f $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_497 N_A_367_119#_c_628_n N_A_359_367#_M1002_g 0.0110341f $X=9.54 $Y=1.185
+ $X2=0 $Y2=0
cc_498 N_A_367_119#_c_639_n N_A_359_367#_M1002_g 0.00788409f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_499 N_A_367_119#_M1028_g N_A_359_367#_M1006_g 0.020603f $X=9.445 $Y=2.475
+ $X2=0 $Y2=0
cc_500 N_A_367_119#_c_631_n N_A_359_367#_c_879_n 8.91886e-19 $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_501 N_A_367_119#_c_637_n N_A_359_367#_c_879_n 0.00160991f $X=6.815 $Y=0.925
+ $X2=0 $Y2=0
cc_502 N_A_367_119#_c_638_n N_A_359_367#_c_879_n 7.00147e-19 $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_503 N_A_367_119#_c_641_n N_A_359_367#_c_879_n 9.08539e-19 $X=6 $Y=0.925 $X2=0
+ $Y2=0
cc_504 N_A_367_119#_c_642_n N_A_359_367#_c_879_n 2.49023e-19 $X=6.96 $Y=0.925
+ $X2=0 $Y2=0
cc_505 N_A_367_119#_c_643_n N_A_359_367#_c_879_n 0.0173566f $X=6.82 $Y=1.165
+ $X2=0 $Y2=0
cc_506 N_A_367_119#_c_648_n N_A_359_367#_c_880_n 0.00305602f $X=9.56 $Y=1.855
+ $X2=0 $Y2=0
cc_507 N_A_367_119#_c_648_n N_A_359_367#_c_889_n 0.020603f $X=9.56 $Y=1.855
+ $X2=0 $Y2=0
cc_508 N_A_367_119#_c_630_n N_A_359_367#_c_890_n 0.0293101f $X=1.805 $Y=2.545
+ $X2=0 $Y2=0
cc_509 N_A_367_119#_c_635_n N_A_359_367#_c_890_n 0.0143476f $X=1.997 $Y=1.585
+ $X2=0 $Y2=0
cc_510 N_A_367_119#_M1000_d N_A_359_367#_c_900_n 0.00694341f $X=2.875 $Y=1.795
+ $X2=0 $Y2=0
cc_511 N_A_367_119#_c_651_n N_A_359_367#_c_900_n 0.0553353f $X=3.095 $Y=2.63
+ $X2=0 $Y2=0
cc_512 N_A_367_119#_c_630_n N_A_359_367#_c_907_n 0.0132519f $X=1.805 $Y=2.545
+ $X2=0 $Y2=0
cc_513 N_A_367_119#_c_651_n N_A_359_367#_c_907_n 0.0129035f $X=3.095 $Y=2.63
+ $X2=0 $Y2=0
cc_514 N_A_367_119#_c_639_n N_A_359_367#_c_881_n 0.00771398f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_515 N_A_367_119#_c_629_n N_A_359_367#_c_882_n 0.00176116f $X=9.54 $Y=1.335
+ $X2=0 $Y2=0
cc_516 N_A_367_119#_c_634_n N_A_359_367#_c_882_n 0.00305602f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_517 N_A_367_119#_c_639_n N_A_359_367#_c_882_n 4.50829e-19 $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_518 N_A_367_119#_M1000_d N_A_359_367#_c_892_n 0.00638987f $X=2.875 $Y=1.795
+ $X2=0 $Y2=0
cc_519 N_A_367_119#_M1010_g N_A_359_367#_c_892_n 0.0137722f $X=5.665 $Y=2.48
+ $X2=0 $Y2=0
cc_520 N_A_367_119#_c_631_n N_A_359_367#_c_892_n 0.00879102f $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_521 N_A_367_119#_c_632_n N_A_359_367#_c_892_n 0.00154213f $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_522 N_A_367_119#_M1000_d N_A_359_367#_c_902_n 0.00127437f $X=2.875 $Y=1.795
+ $X2=0 $Y2=0
cc_523 N_A_367_119#_c_651_n N_A_359_367#_c_902_n 0.00132944f $X=3.095 $Y=2.63
+ $X2=0 $Y2=0
cc_524 N_A_367_119#_c_637_n N_A_359_367#_c_883_n 0.00548528f $X=6.815 $Y=0.925
+ $X2=0 $Y2=0
cc_525 N_A_367_119#_M1010_g N_A_359_367#_c_884_n 0.00244376f $X=5.665 $Y=2.48
+ $X2=0 $Y2=0
cc_526 N_A_367_119#_c_642_n N_A_359_367#_c_884_n 3.32097e-19 $X=6.96 $Y=0.925
+ $X2=0 $Y2=0
cc_527 N_A_367_119#_c_643_n N_A_359_367#_c_884_n 0.0025584f $X=6.82 $Y=1.165
+ $X2=0 $Y2=0
cc_528 N_A_367_119#_M1000_d N_A_359_367#_c_885_n 0.00892671f $X=2.875 $Y=1.795
+ $X2=0 $Y2=0
cc_529 N_A_367_119#_c_636_n N_A_359_367#_c_885_n 0.0305666f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_530 N_A_367_119#_c_639_n N_CI_c_1072_n 0.00228377f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_531 N_A_367_119#_c_639_n N_CI_c_1073_n 0.0149219f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_532 N_A_367_119#_c_643_n N_CI_c_1073_n 0.00462987f $X=6.82 $Y=1.165 $X2=0
+ $Y2=0
cc_533 N_A_367_119#_c_644_n N_CI_c_1073_n 0.00863876f $X=6.82 $Y=1 $X2=0 $Y2=0
cc_534 N_A_367_119#_c_639_n N_CI_c_1075_n 0.00941657f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_535 N_A_367_119#_c_639_n CI 0.00584484f $X=9.215 $Y=0.925 $X2=0 $Y2=0
cc_536 N_A_367_119#_c_639_n N_A_1571_367#_M1012_d 0.00435947f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_537 N_A_367_119#_c_628_n N_A_1571_367#_M1015_g 0.0109986f $X=9.54 $Y=1.185
+ $X2=0 $Y2=0
cc_538 N_A_367_119#_c_629_n N_A_1571_367#_M1015_g 0.00875741f $X=9.54 $Y=1.335
+ $X2=0 $Y2=0
cc_539 N_A_367_119#_c_633_n N_A_1571_367#_M1015_g 0.00131196f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_540 N_A_367_119#_c_639_n N_A_1571_367#_c_1137_n 0.0190948f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_541 N_A_367_119#_M1028_g N_A_1571_367#_c_1144_n 0.0117331f $X=9.445 $Y=2.475
+ $X2=0 $Y2=0
cc_542 N_A_367_119#_c_639_n N_A_1571_367#_c_1158_n 0.0216944f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_543 N_A_367_119#_M1028_g N_A_1571_367#_c_1148_n 0.00887605f $X=9.445 $Y=2.475
+ $X2=0 $Y2=0
cc_544 N_A_367_119#_c_648_n N_A_1571_367#_c_1148_n 0.00477539f $X=9.56 $Y=1.855
+ $X2=0 $Y2=0
cc_545 N_A_367_119#_c_633_n N_A_1571_367#_c_1148_n 0.0150854f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_546 N_A_367_119#_M1028_g N_A_1571_367#_c_1149_n 0.00282153f $X=9.445 $Y=2.475
+ $X2=0 $Y2=0
cc_547 N_A_367_119#_c_648_n N_A_1571_367#_c_1149_n 6.26196e-19 $X=9.56 $Y=1.855
+ $X2=0 $Y2=0
cc_548 N_A_367_119#_c_633_n N_A_1571_367#_c_1149_n 0.0068797f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_549 N_A_367_119#_c_633_n N_A_1571_367#_c_1139_n 0.0241542f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_550 N_A_367_119#_c_634_n N_A_1571_367#_c_1139_n 0.00222347f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_551 N_A_367_119#_M1028_g N_A_1571_367#_c_1140_n 0.00110592f $X=9.445 $Y=2.475
+ $X2=0 $Y2=0
cc_552 N_A_367_119#_c_633_n N_A_1571_367#_c_1140_n 3.90191e-19 $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_553 N_A_367_119#_c_634_n N_A_1571_367#_c_1140_n 0.0269391f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_554 N_A_367_119#_c_639_n N_A_1758_87#_M1002_d 0.00228315f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_555 N_A_367_119#_c_774_p N_A_1758_87#_M1002_d 0.00184657f $X=9.36 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_556 N_A_367_119#_c_628_n N_A_1758_87#_c_1271_n 0.00975764f $X=9.54 $Y=1.185
+ $X2=0 $Y2=0
cc_557 N_A_367_119#_c_639_n N_A_1758_87#_c_1271_n 0.0189314f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_558 N_A_367_119#_c_774_p N_A_1758_87#_c_1271_n 0.00141363f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_559 N_A_367_119#_c_778_p N_A_1758_87#_c_1271_n 0.0111543f $X=9.585 $Y=0.925
+ $X2=0 $Y2=0
cc_560 N_A_367_119#_c_629_n N_A_1758_87#_c_1260_n 8.74235e-19 $X=9.54 $Y=1.335
+ $X2=0 $Y2=0
cc_561 N_A_367_119#_c_628_n N_A_1758_87#_c_1261_n 0.0119635f $X=9.54 $Y=1.185
+ $X2=0 $Y2=0
cc_562 N_A_367_119#_c_639_n N_A_1758_87#_c_1261_n 0.00424117f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_563 N_A_367_119#_c_774_p N_A_1758_87#_c_1261_n 0.00724804f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_564 N_A_367_119#_c_778_p N_A_1758_87#_c_1261_n 0.0111857f $X=9.585 $Y=0.925
+ $X2=0 $Y2=0
cc_565 N_A_367_119#_c_633_n N_A_1758_87#_c_1263_n 0.0319561f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_566 N_A_367_119#_c_634_n N_A_1758_87#_c_1263_n 0.00740952f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_567 N_A_367_119#_c_628_n N_A_1758_87#_c_1282_n 8.74235e-19 $X=9.54 $Y=1.185
+ $X2=0 $Y2=0
cc_568 N_A_367_119#_c_633_n N_A_1758_87#_c_1282_n 0.00656034f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_569 N_A_367_119#_c_639_n N_A_1758_87#_c_1282_n 0.0149312f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_570 N_A_367_119#_c_774_p N_A_1758_87#_c_1282_n 0.00141363f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_571 N_A_367_119#_c_629_n N_A_1758_87#_c_1265_n 0.0015305f $X=9.54 $Y=1.335
+ $X2=0 $Y2=0
cc_572 N_A_367_119#_c_633_n N_A_1758_87#_c_1265_n 0.0123954f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_573 N_A_367_119#_c_634_n N_A_1758_87#_c_1265_n 6.76053e-19 $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_574 N_A_367_119#_c_639_n N_A_1758_87#_c_1265_n 0.00589449f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_575 N_A_367_119#_c_774_p N_A_1758_87#_c_1265_n 0.0039255f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_576 N_A_367_119#_c_778_p N_A_1758_87#_c_1265_n 0.00182491f $X=9.585 $Y=0.925
+ $X2=0 $Y2=0
cc_577 N_A_367_119#_M1010_g N_VPWR_c_1367_n 0.00534427f $X=5.665 $Y=2.48 $X2=0
+ $Y2=0
cc_578 N_A_367_119#_M1028_g N_VPWR_c_1368_n 8.5177e-19 $X=9.445 $Y=2.475 $X2=0
+ $Y2=0
cc_579 N_A_367_119#_M1010_g N_VPWR_c_1360_n 0.00526787f $X=5.665 $Y=2.48 $X2=0
+ $Y2=0
cc_580 N_A_367_119#_c_630_n N_A_247_367#_c_1468_n 0.0399455f $X=1.805 $Y=2.545
+ $X2=0 $Y2=0
cc_581 N_A_367_119#_c_650_n N_A_247_367#_c_1463_n 0.0134603f $X=1.89 $Y=2.63
+ $X2=0 $Y2=0
cc_582 N_A_367_119#_c_664_n N_A_247_367#_c_1473_n 0.00122333f $X=2.305 $Y=0.925
+ $X2=0 $Y2=0
cc_583 N_A_367_119#_c_650_n N_A_247_367#_c_1464_n 0.0124675f $X=1.89 $Y=2.63
+ $X2=0 $Y2=0
cc_584 N_A_367_119#_c_651_n N_A_247_367#_c_1464_n 0.0909222f $X=3.095 $Y=2.63
+ $X2=0 $Y2=0
cc_585 N_A_367_119#_c_636_n N_A_247_367#_c_1458_n 0.0379151f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_586 N_A_367_119#_c_651_n N_A_247_367#_c_1459_n 0.0117182f $X=3.095 $Y=2.63
+ $X2=0 $Y2=0
cc_587 N_A_367_119#_c_635_n N_A_247_367#_c_1460_n 0.0399455f $X=1.997 $Y=1.585
+ $X2=0 $Y2=0
cc_588 N_A_367_119#_c_645_n N_A_247_367#_c_1460_n 0.00866185f $X=2.09 $Y=0.78
+ $X2=0 $Y2=0
cc_589 N_A_367_119#_c_638_n N_A_1034_380#_M1008_d 0.00138706f $X=6.145 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_590 N_A_367_119#_c_641_n N_A_1034_380#_M1008_d 8.29327e-19 $X=6 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_591 N_A_367_119#_M1010_g N_A_1034_380#_c_1533_n 0.00819766f $X=5.665 $Y=2.48
+ $X2=0 $Y2=0
cc_592 N_A_367_119#_c_636_n N_A_1034_380#_c_1539_n 0.00859591f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_593 N_A_367_119#_c_641_n N_A_1034_380#_c_1539_n 0.00726023f $X=6 $Y=0.925
+ $X2=0 $Y2=0
cc_594 N_A_367_119#_c_631_n N_A_1034_380#_c_1532_n 0.0489768f $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_595 N_A_367_119#_c_632_n N_A_1034_380#_c_1532_n 0.00819766f $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_596 N_A_367_119#_c_636_n N_A_1034_380#_c_1532_n 0.0181498f $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_597 N_A_367_119#_c_638_n N_A_1034_380#_c_1532_n 4.11999e-19 $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_598 N_A_367_119#_c_641_n N_A_1034_380#_c_1532_n 0.0133502f $X=6 $Y=0.925
+ $X2=0 $Y2=0
cc_599 N_A_367_119#_c_636_n N_A_1034_380#_c_1547_n 4.09611e-19 $X=5.855 $Y=0.925
+ $X2=0 $Y2=0
cc_600 N_A_367_119#_c_638_n N_A_1034_380#_c_1547_n 0.00742907f $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_601 N_A_367_119#_c_641_n N_A_1034_380#_c_1547_n 0.0142993f $X=6 $Y=0.925
+ $X2=0 $Y2=0
cc_602 N_A_367_119#_c_637_n N_COUT_N_M1020_d 0.0041739f $X=6.815 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_603 N_A_367_119#_c_642_n N_COUT_N_M1020_d 0.00249905f $X=6.96 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_604 N_A_367_119#_M1010_g N_COUT_N_c_1586_n 0.0202872f $X=5.665 $Y=2.48 $X2=0
+ $Y2=0
cc_605 N_A_367_119#_c_632_n N_COUT_N_c_1586_n 0.00134737f $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_606 N_A_367_119#_c_631_n N_COUT_N_c_1583_n 0.00629166f $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_607 N_A_367_119#_c_637_n N_COUT_N_c_1583_n 0.00966925f $X=6.815 $Y=0.925
+ $X2=0 $Y2=0
cc_608 N_A_367_119#_c_638_n N_COUT_N_c_1583_n 0.00227568f $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_609 N_A_367_119#_c_640_n N_COUT_N_c_1583_n 0.00111136f $X=7.105 $Y=0.925
+ $X2=0 $Y2=0
cc_610 N_A_367_119#_c_641_n N_COUT_N_c_1583_n 0.011582f $X=6 $Y=0.925 $X2=0
+ $Y2=0
cc_611 N_A_367_119#_c_642_n N_COUT_N_c_1583_n 0.0271091f $X=6.96 $Y=0.925 $X2=0
+ $Y2=0
cc_612 N_A_367_119#_c_643_n N_COUT_N_c_1583_n 0.0012493f $X=6.82 $Y=1.165 $X2=0
+ $Y2=0
cc_613 N_A_367_119#_c_644_n N_COUT_N_c_1583_n 0.00382895f $X=6.82 $Y=1 $X2=0
+ $Y2=0
cc_614 N_A_367_119#_M1010_g N_COUT_N_c_1584_n 0.00386934f $X=5.665 $Y=2.48 $X2=0
+ $Y2=0
cc_615 N_A_367_119#_c_631_n N_COUT_N_c_1584_n 0.024344f $X=5.755 $Y=1.575 $X2=0
+ $Y2=0
cc_616 N_A_367_119#_c_632_n N_COUT_N_c_1584_n 0.00261908f $X=5.755 $Y=1.575
+ $X2=0 $Y2=0
cc_617 N_A_367_119#_c_631_n N_COUT_N_c_1585_n 0.013301f $X=5.755 $Y=1.575 $X2=0
+ $Y2=0
cc_618 N_A_367_119#_c_637_n N_COUT_N_c_1585_n 0.00704492f $X=6.815 $Y=0.925
+ $X2=0 $Y2=0
cc_619 N_A_367_119#_c_638_n N_COUT_N_c_1585_n 0.00330148f $X=6.145 $Y=0.925
+ $X2=0 $Y2=0
cc_620 N_A_367_119#_c_641_n N_COUT_N_c_1585_n 0.00494826f $X=6 $Y=0.925 $X2=0
+ $Y2=0
cc_621 N_A_367_119#_c_642_n N_COUT_N_c_1585_n 0.00859743f $X=6.96 $Y=0.925 $X2=0
+ $Y2=0
cc_622 N_A_367_119#_c_643_n N_COUT_N_c_1585_n 6.79428e-19 $X=6.82 $Y=1.165 $X2=0
+ $Y2=0
cc_623 N_A_367_119#_c_637_n COUT_N 0.00840053f $X=6.815 $Y=0.925 $X2=0 $Y2=0
cc_624 N_A_367_119#_c_644_n COUT_N 0.00517844f $X=6.82 $Y=1 $X2=0 $Y2=0
cc_625 N_A_367_119#_c_639_n N_A_1340_412#_M1009_d 0.00972737f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_626 N_A_367_119#_c_640_n N_A_1340_412#_M1009_d 0.00634315f $X=7.105 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_627 N_A_367_119#_c_642_n N_A_1340_412#_M1009_d 8.49051e-19 $X=6.96 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_628 N_A_367_119#_c_639_n N_A_1340_412#_c_1642_n 0.0043823f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_629 N_A_367_119#_c_640_n N_A_1340_412#_c_1642_n 0.00293566f $X=7.105 $Y=0.925
+ $X2=0 $Y2=0
cc_630 N_A_367_119#_c_642_n N_A_1340_412#_c_1642_n 0.0134031f $X=6.96 $Y=0.925
+ $X2=0 $Y2=0
cc_631 N_A_367_119#_c_643_n N_A_1340_412#_c_1642_n 8.61636e-19 $X=6.82 $Y=1.165
+ $X2=0 $Y2=0
cc_632 N_A_367_119#_c_639_n N_A_1340_412#_c_1643_n 0.0253521f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_633 N_A_367_119#_c_640_n N_A_1340_412#_c_1643_n 0.00321414f $X=7.105 $Y=0.925
+ $X2=0 $Y2=0
cc_634 N_A_367_119#_c_642_n N_A_1340_412#_c_1643_n 0.0366415f $X=6.96 $Y=0.925
+ $X2=0 $Y2=0
cc_635 N_A_367_119#_c_643_n N_A_1340_412#_c_1643_n 0.001173f $X=6.82 $Y=1.165
+ $X2=0 $Y2=0
cc_636 N_A_367_119#_c_644_n N_A_1340_412#_c_1643_n 0.00920181f $X=6.82 $Y=1
+ $X2=0 $Y2=0
cc_637 N_A_367_119#_c_633_n N_A_1708_411#_M1019_d 7.33641e-19 $X=9.585 $Y=1.35
+ $X2=-0.19 $Y2=-0.245
cc_638 N_A_367_119#_c_778_p N_A_1708_411#_M1019_d 0.00477759f $X=9.585 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_639 N_A_367_119#_M1028_g N_A_1708_411#_c_1690_n 0.0107463f $X=9.445 $Y=2.475
+ $X2=0 $Y2=0
cc_640 N_A_367_119#_c_628_n N_A_1708_411#_c_1696_n 0.00424549f $X=9.54 $Y=1.185
+ $X2=0 $Y2=0
cc_641 N_A_367_119#_c_633_n N_A_1708_411#_c_1696_n 0.00241208f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_642 N_A_367_119#_c_774_p N_A_1708_411#_c_1696_n 0.00112754f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_643 N_A_367_119#_c_778_p N_A_1708_411#_c_1696_n 0.0159858f $X=9.585 $Y=0.925
+ $X2=0 $Y2=0
cc_644 N_A_367_119#_c_629_n N_A_1708_411#_c_1688_n 5.53631e-19 $X=9.54 $Y=1.335
+ $X2=0 $Y2=0
cc_645 N_A_367_119#_c_633_n N_A_1708_411#_c_1688_n 0.0136102f $X=9.585 $Y=1.35
+ $X2=0 $Y2=0
cc_646 N_A_367_119#_M1028_g N_A_1708_411#_c_1702_n 0.00348908f $X=9.445 $Y=2.475
+ $X2=0 $Y2=0
cc_647 N_A_367_119#_M1028_g N_A_1708_411#_c_1692_n 7.29384e-19 $X=9.445 $Y=2.475
+ $X2=0 $Y2=0
cc_648 N_A_367_119#_c_636_n N_VGND_M1011_d 0.0105581f $X=5.855 $Y=0.925 $X2=0
+ $Y2=0
cc_649 N_A_367_119#_c_639_n N_VGND_M1016_d 0.00828624f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_650 N_A_367_119#_c_636_n N_VGND_c_1760_n 0.0232255f $X=5.855 $Y=0.925 $X2=0
+ $Y2=0
cc_651 N_A_367_119#_c_639_n N_VGND_c_1761_n 0.02342f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_652 N_A_367_119#_c_628_n N_VGND_c_1763_n 8.5177e-19 $X=9.54 $Y=1.185 $X2=0
+ $Y2=0
cc_653 N_A_367_119#_c_644_n N_VGND_c_1766_n 0.00570116f $X=6.82 $Y=1 $X2=0 $Y2=0
cc_654 N_A_367_119#_c_641_n N_VGND_c_1768_n 3.06625e-19 $X=6 $Y=0.925 $X2=0
+ $Y2=0
cc_655 N_A_367_119#_c_642_n N_VGND_c_1768_n 0.0113144f $X=6.96 $Y=0.925 $X2=0
+ $Y2=0
cc_656 N_A_367_119#_c_644_n N_VGND_c_1768_n 0.00812063f $X=6.82 $Y=1 $X2=0 $Y2=0
cc_657 N_A_359_367#_c_893_n N_CI_M1026_g 0.00789153f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_658 N_A_359_367#_c_883_n N_CI_M1026_g 2.46678e-19 $X=6.485 $Y=1.735 $X2=0
+ $Y2=0
cc_659 N_A_359_367#_c_884_n N_CI_M1026_g 0.0235004f $X=6.625 $Y=1.735 $X2=0
+ $Y2=0
cc_660 N_A_359_367#_c_880_n N_CI_M1023_g 0.00401156f $X=8.655 $Y=1.745 $X2=0
+ $Y2=0
cc_661 N_A_359_367#_c_893_n N_CI_M1023_g 0.0078084f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_662 N_A_359_367#_M1002_g N_CI_c_1075_n 0.0137077f $X=8.715 $Y=0.755 $X2=0
+ $Y2=0
cc_663 N_A_359_367#_c_893_n CI 0.00481906f $X=8.735 $Y=2.035 $X2=0 $Y2=0
cc_664 N_A_359_367#_c_881_n N_CI_c_1078_n 2.54337e-19 $X=8.655 $Y=1.39 $X2=0
+ $Y2=0
cc_665 N_A_359_367#_c_882_n N_CI_c_1078_n 0.0147722f $X=8.655 $Y=1.39 $X2=0
+ $Y2=0
cc_666 N_A_359_367#_M1006_g N_A_1571_367#_c_1142_n 0.0104681f $X=9.015 $Y=2.475
+ $X2=0 $Y2=0
cc_667 N_A_359_367#_c_893_n N_A_1571_367#_c_1142_n 0.0306408f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_668 N_A_359_367#_c_895_n N_A_1571_367#_c_1142_n 0.00121658f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_669 N_A_359_367#_M1002_g N_A_1571_367#_c_1137_n 0.00642634f $X=8.715 $Y=0.755
+ $X2=0 $Y2=0
cc_670 N_A_359_367#_M1006_g N_A_1571_367#_c_1144_n 0.0150605f $X=9.015 $Y=2.475
+ $X2=0 $Y2=0
cc_671 N_A_359_367#_c_889_n N_A_1571_367#_c_1144_n 0.00340207f $X=9.015 $Y=1.82
+ $X2=0 $Y2=0
cc_672 N_A_359_367#_c_891_n N_A_1571_367#_c_1144_n 0.0062393f $X=8.655 $Y=1.725
+ $X2=0 $Y2=0
cc_673 N_A_359_367#_c_893_n N_A_1571_367#_c_1144_n 0.0101915f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_674 N_A_359_367#_c_895_n N_A_1571_367#_c_1144_n 0.00399037f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_675 N_A_359_367#_M1006_g N_A_1571_367#_c_1145_n 0.00109823f $X=9.015 $Y=2.475
+ $X2=0 $Y2=0
cc_676 N_A_359_367#_c_880_n N_A_1571_367#_c_1145_n 0.0032957f $X=8.655 $Y=1.745
+ $X2=0 $Y2=0
cc_677 N_A_359_367#_c_891_n N_A_1571_367#_c_1145_n 0.00841698f $X=8.655 $Y=1.725
+ $X2=0 $Y2=0
cc_678 N_A_359_367#_c_893_n N_A_1571_367#_c_1145_n 0.0272331f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_679 N_A_359_367#_c_895_n N_A_1571_367#_c_1145_n 0.00121658f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_680 N_A_359_367#_M1002_g N_A_1571_367#_c_1138_n 0.00162099f $X=8.715 $Y=0.755
+ $X2=0 $Y2=0
cc_681 N_A_359_367#_c_891_n N_A_1571_367#_c_1138_n 0.0129718f $X=8.655 $Y=1.725
+ $X2=0 $Y2=0
cc_682 N_A_359_367#_c_881_n N_A_1571_367#_c_1138_n 0.0343332f $X=8.655 $Y=1.39
+ $X2=0 $Y2=0
cc_683 N_A_359_367#_c_882_n N_A_1571_367#_c_1138_n 0.0032957f $X=8.655 $Y=1.39
+ $X2=0 $Y2=0
cc_684 N_A_359_367#_c_882_n N_A_1571_367#_c_1158_n 0.00280109f $X=8.655 $Y=1.39
+ $X2=0 $Y2=0
cc_685 N_A_359_367#_M1006_g N_A_1571_367#_c_1148_n 9.85849e-19 $X=9.015 $Y=2.475
+ $X2=0 $Y2=0
cc_686 N_A_359_367#_M1002_g N_A_1758_87#_c_1271_n 0.00644937f $X=8.715 $Y=0.755
+ $X2=0 $Y2=0
cc_687 N_A_359_367#_M1002_g N_A_1758_87#_c_1260_n 0.002211f $X=8.715 $Y=0.755
+ $X2=0 $Y2=0
cc_688 N_A_359_367#_M1002_g N_A_1758_87#_c_1262_n 0.00422714f $X=8.715 $Y=0.755
+ $X2=0 $Y2=0
cc_689 N_A_359_367#_c_880_n N_A_1758_87#_c_1263_n 0.00302898f $X=8.655 $Y=1.745
+ $X2=0 $Y2=0
cc_690 N_A_359_367#_c_889_n N_A_1758_87#_c_1263_n 0.0024353f $X=9.015 $Y=1.82
+ $X2=0 $Y2=0
cc_691 N_A_359_367#_c_891_n N_A_1758_87#_c_1263_n 0.025102f $X=8.655 $Y=1.725
+ $X2=0 $Y2=0
cc_692 N_A_359_367#_c_881_n N_A_1758_87#_c_1263_n 0.0126865f $X=8.655 $Y=1.39
+ $X2=0 $Y2=0
cc_693 N_A_359_367#_c_895_n N_A_1758_87#_c_1263_n 0.00675724f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_694 N_A_359_367#_M1002_g N_A_1758_87#_c_1282_n 0.00400097f $X=8.715 $Y=0.755
+ $X2=0 $Y2=0
cc_695 N_A_359_367#_c_889_n N_A_1758_87#_c_1282_n 5.02333e-19 $X=9.015 $Y=1.82
+ $X2=0 $Y2=0
cc_696 N_A_359_367#_c_891_n N_A_1758_87#_c_1282_n 0.00393472f $X=8.655 $Y=1.725
+ $X2=0 $Y2=0
cc_697 N_A_359_367#_c_889_n N_A_1758_87#_c_1265_n 0.00449582f $X=9.015 $Y=1.82
+ $X2=0 $Y2=0
cc_698 N_A_359_367#_c_891_n N_A_1758_87#_c_1265_n 0.00179843f $X=8.655 $Y=1.725
+ $X2=0 $Y2=0
cc_699 N_A_359_367#_c_881_n N_A_1758_87#_c_1265_n 0.0121332f $X=8.655 $Y=1.39
+ $X2=0 $Y2=0
cc_700 N_A_359_367#_c_882_n N_A_1758_87#_c_1265_n 0.00179047f $X=8.655 $Y=1.39
+ $X2=0 $Y2=0
cc_701 N_A_359_367#_c_895_n N_A_1758_87#_c_1265_n 0.00201715f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_702 N_A_359_367#_c_892_n N_VPWR_M1027_d 0.00881001f $X=6.335 $Y=2.035 $X2=0
+ $Y2=0
cc_703 N_A_359_367#_c_893_n N_VPWR_M1026_d 0.00410777f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_704 N_A_359_367#_c_892_n N_VPWR_c_1362_n 0.031153f $X=6.335 $Y=2.035 $X2=0
+ $Y2=0
cc_705 N_A_359_367#_M1014_g N_VPWR_c_1363_n 0.00196343f $X=6.625 $Y=2.48 $X2=0
+ $Y2=0
cc_706 N_A_359_367#_c_893_n N_VPWR_c_1363_n 0.0323919f $X=8.735 $Y=2.035 $X2=0
+ $Y2=0
cc_707 N_A_359_367#_M1014_g N_VPWR_c_1367_n 0.00534427f $X=6.625 $Y=2.48 $X2=0
+ $Y2=0
cc_708 N_A_359_367#_M1006_g N_VPWR_c_1368_n 8.5177e-19 $X=9.015 $Y=2.475 $X2=0
+ $Y2=0
cc_709 N_A_359_367#_M1014_g N_VPWR_c_1360_n 0.00526787f $X=6.625 $Y=2.48 $X2=0
+ $Y2=0
cc_710 N_A_359_367#_c_885_n N_A_247_367#_c_1458_n 0.0931175f $X=3.095 $Y=1 $X2=0
+ $Y2=0
cc_711 N_A_359_367#_c_900_n N_A_247_367#_c_1459_n 0.0117125f $X=2.93 $Y=2.28
+ $X2=0 $Y2=0
cc_712 N_A_359_367#_c_892_n N_A_247_367#_c_1459_n 0.0409814f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_713 N_A_359_367#_c_902_n N_A_247_367#_c_1459_n 0.0025135f $X=3.265 $Y=2.035
+ $X2=0 $Y2=0
cc_714 N_A_359_367#_c_892_n N_A_1034_380#_M1024_d 0.00441205f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_715 N_A_359_367#_c_892_n N_A_1034_380#_c_1533_n 0.0174072f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_716 N_A_359_367#_c_892_n N_A_1034_380#_c_1534_n 0.0216001f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_717 N_A_359_367#_c_876_n N_A_1034_380#_c_1547_n 0.00447965f $X=6.175 $Y=1
+ $X2=0 $Y2=0
cc_718 N_A_359_367#_c_892_n N_COUT_N_M1010_d 0.0101173f $X=6.335 $Y=2.035 $X2=0
+ $Y2=0
cc_719 N_A_359_367#_c_894_n N_COUT_N_M1010_d 0.00666521f $X=6.625 $Y=2.035 $X2=0
+ $Y2=0
cc_720 N_A_359_367#_c_883_n N_COUT_N_M1010_d 0.00228301f $X=6.485 $Y=1.735 $X2=0
+ $Y2=0
cc_721 N_A_359_367#_M1014_g N_COUT_N_c_1586_n 0.0154002f $X=6.625 $Y=2.48 $X2=0
+ $Y2=0
cc_722 N_A_359_367#_c_892_n N_COUT_N_c_1586_n 0.0253988f $X=6.335 $Y=2.035 $X2=0
+ $Y2=0
cc_723 N_A_359_367#_c_894_n N_COUT_N_c_1586_n 0.00137493f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_724 N_A_359_367#_c_876_n N_COUT_N_c_1583_n 0.00278395f $X=6.175 $Y=1 $X2=0
+ $Y2=0
cc_725 N_A_359_367#_c_877_n N_COUT_N_c_1583_n 0.00221032f $X=6.34 $Y=1.57 $X2=0
+ $Y2=0
cc_726 N_A_359_367#_c_879_n N_COUT_N_c_1583_n 0.00665297f $X=6.34 $Y=1.075 $X2=0
+ $Y2=0
cc_727 N_A_359_367#_c_877_n N_COUT_N_c_1584_n 0.00752436f $X=6.34 $Y=1.57 $X2=0
+ $Y2=0
cc_728 N_A_359_367#_M1014_g N_COUT_N_c_1584_n 0.00114064f $X=6.625 $Y=2.48 $X2=0
+ $Y2=0
cc_729 N_A_359_367#_c_892_n N_COUT_N_c_1584_n 0.00748389f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_730 N_A_359_367#_c_894_n N_COUT_N_c_1584_n 0.0013541f $X=6.625 $Y=2.035 $X2=0
+ $Y2=0
cc_731 N_A_359_367#_c_883_n N_COUT_N_c_1584_n 0.0397689f $X=6.485 $Y=1.735 $X2=0
+ $Y2=0
cc_732 N_A_359_367#_c_877_n N_COUT_N_c_1585_n 0.0108793f $X=6.34 $Y=1.57 $X2=0
+ $Y2=0
cc_733 N_A_359_367#_c_879_n N_COUT_N_c_1585_n 0.00716369f $X=6.34 $Y=1.075 $X2=0
+ $Y2=0
cc_734 N_A_359_367#_c_892_n N_COUT_N_c_1585_n 0.00414617f $X=6.335 $Y=2.035
+ $X2=0 $Y2=0
cc_735 N_A_359_367#_c_894_n N_COUT_N_c_1585_n 0.00187256f $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_736 N_A_359_367#_c_883_n N_COUT_N_c_1585_n 0.00617021f $X=6.485 $Y=1.735
+ $X2=0 $Y2=0
cc_737 N_A_359_367#_c_884_n N_COUT_N_c_1585_n 4.17737e-19 $X=6.625 $Y=1.735
+ $X2=0 $Y2=0
cc_738 N_A_359_367#_c_879_n COUT_N 3.2583e-19 $X=6.34 $Y=1.075 $X2=0 $Y2=0
cc_739 N_A_359_367#_c_893_n N_A_1340_412#_M1014_d 0.0111265f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_740 N_A_359_367#_c_893_n N_A_1340_412#_c_1644_n 0.0237014f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_741 N_A_359_367#_c_894_n N_A_1340_412#_c_1644_n 6.43861e-19 $X=6.625 $Y=2.035
+ $X2=0 $Y2=0
cc_742 N_A_359_367#_c_883_n N_A_1340_412#_c_1644_n 0.0279987f $X=6.485 $Y=1.735
+ $X2=0 $Y2=0
cc_743 N_A_359_367#_c_884_n N_A_1340_412#_c_1644_n 0.014354f $X=6.625 $Y=1.735
+ $X2=0 $Y2=0
cc_744 N_A_359_367#_c_877_n N_A_1340_412#_c_1642_n 0.00107864f $X=6.34 $Y=1.57
+ $X2=0 $Y2=0
cc_745 N_A_359_367#_c_893_n N_A_1340_412#_c_1642_n 0.00944525f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_746 N_A_359_367#_c_883_n N_A_1340_412#_c_1642_n 0.0076651f $X=6.485 $Y=1.735
+ $X2=0 $Y2=0
cc_747 N_A_359_367#_c_884_n N_A_1340_412#_c_1642_n 0.0011702f $X=6.625 $Y=1.735
+ $X2=0 $Y2=0
cc_748 N_A_359_367#_c_891_n N_A_1708_411#_M1006_s 0.00204427f $X=8.655 $Y=1.725
+ $X2=0 $Y2=0
cc_749 N_A_359_367#_c_893_n N_A_1708_411#_M1006_s 0.00233928f $X=8.735 $Y=2.035
+ $X2=0 $Y2=0
cc_750 N_A_359_367#_c_895_n N_A_1708_411#_M1006_s 0.0020856f $X=8.88 $Y=2.035
+ $X2=0 $Y2=0
cc_751 N_A_359_367#_M1006_g N_A_1708_411#_c_1690_n 0.010456f $X=9.015 $Y=2.475
+ $X2=0 $Y2=0
cc_752 N_A_359_367#_M1002_g N_VGND_c_1763_n 0.00456612f $X=8.715 $Y=0.755 $X2=0
+ $Y2=0
cc_753 N_A_359_367#_c_876_n N_VGND_c_1766_n 0.00534858f $X=6.175 $Y=1 $X2=0
+ $Y2=0
cc_754 N_A_359_367#_c_876_n N_VGND_c_1768_n 0.0104808f $X=6.175 $Y=1 $X2=0 $Y2=0
cc_755 N_A_359_367#_M1002_g N_VGND_c_1768_n 0.00437689f $X=8.715 $Y=0.755 $X2=0
+ $Y2=0
cc_756 N_CI_M1023_g N_A_1571_367#_c_1142_n 0.00628028f $X=7.78 $Y=2.465 $X2=0
+ $Y2=0
cc_757 N_CI_M1023_g N_A_1571_367#_c_1143_n 0.00390528f $X=7.78 $Y=2.465 $X2=0
+ $Y2=0
cc_758 N_CI_c_1073_n N_A_1571_367#_c_1137_n 0.00104513f $X=7.63 $Y=1.185 $X2=0
+ $Y2=0
cc_759 N_CI_c_1075_n N_A_1571_367#_c_1137_n 0.00761193f $X=8.17 $Y=1.185 $X2=0
+ $Y2=0
cc_760 N_CI_M1026_g N_A_1571_367#_c_1145_n 4.91214e-19 $X=7.27 $Y=2.335 $X2=0
+ $Y2=0
cc_761 N_CI_M1023_g N_A_1571_367#_c_1145_n 0.00375127f $X=7.78 $Y=2.465 $X2=0
+ $Y2=0
cc_762 CI N_A_1571_367#_c_1145_n 0.00996515f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_763 N_CI_c_1078_n N_A_1571_367#_c_1145_n 0.00894115f $X=8.17 $Y=1.35 $X2=0
+ $Y2=0
cc_764 N_CI_M1023_g N_A_1571_367#_c_1138_n 0.00565587f $X=7.78 $Y=2.465 $X2=0
+ $Y2=0
cc_765 N_CI_c_1075_n N_A_1571_367#_c_1138_n 0.00359083f $X=8.17 $Y=1.185 $X2=0
+ $Y2=0
cc_766 CI N_A_1571_367#_c_1138_n 0.0228396f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_767 N_CI_c_1078_n N_A_1571_367#_c_1138_n 0.00844269f $X=8.17 $Y=1.35 $X2=0
+ $Y2=0
cc_768 N_CI_M1023_g N_A_1571_367#_c_1147_n 0.00348017f $X=7.78 $Y=2.465 $X2=0
+ $Y2=0
cc_769 N_CI_c_1075_n N_A_1571_367#_c_1158_n 0.00182727f $X=8.17 $Y=1.185 $X2=0
+ $Y2=0
cc_770 N_CI_c_1075_n N_A_1758_87#_c_1271_n 2.35772e-19 $X=8.17 $Y=1.185 $X2=0
+ $Y2=0
cc_771 N_CI_M1026_g N_VPWR_c_1363_n 0.0183256f $X=7.27 $Y=2.335 $X2=0 $Y2=0
cc_772 N_CI_M1023_g N_VPWR_c_1363_n 0.0129131f $X=7.78 $Y=2.465 $X2=0 $Y2=0
cc_773 N_CI_c_1077_n N_VPWR_c_1363_n 0.00534304f $X=7.555 $Y=1.35 $X2=0 $Y2=0
cc_774 N_CI_M1026_g N_VPWR_c_1367_n 0.00407914f $X=7.27 $Y=2.335 $X2=0 $Y2=0
cc_775 N_CI_M1023_g N_VPWR_c_1368_n 0.00549284f $X=7.78 $Y=2.465 $X2=0 $Y2=0
cc_776 N_CI_M1026_g N_VPWR_c_1360_n 0.00425776f $X=7.27 $Y=2.335 $X2=0 $Y2=0
cc_777 N_CI_M1023_g N_VPWR_c_1360_n 0.0126f $X=7.78 $Y=2.465 $X2=0 $Y2=0
cc_778 N_CI_M1026_g N_A_1340_412#_c_1644_n 0.0151184f $X=7.27 $Y=2.335 $X2=0
+ $Y2=0
cc_779 N_CI_M1026_g N_A_1340_412#_c_1642_n 0.00900962f $X=7.27 $Y=2.335 $X2=0
+ $Y2=0
cc_780 N_CI_c_1072_n N_A_1340_412#_c_1642_n 0.00103376f $X=7.345 $Y=1.44 $X2=0
+ $Y2=0
cc_781 N_CI_M1023_g N_A_1340_412#_c_1642_n 0.00419545f $X=7.78 $Y=2.465 $X2=0
+ $Y2=0
cc_782 N_CI_c_1077_n N_A_1340_412#_c_1642_n 0.00115788f $X=7.555 $Y=1.35 $X2=0
+ $Y2=0
cc_783 N_CI_c_1072_n N_A_1340_412#_c_1643_n 0.0105837f $X=7.345 $Y=1.44 $X2=0
+ $Y2=0
cc_784 N_CI_c_1073_n N_A_1340_412#_c_1643_n 0.0165647f $X=7.63 $Y=1.185 $X2=0
+ $Y2=0
cc_785 N_CI_c_1075_n N_A_1340_412#_c_1643_n 3.79652e-19 $X=8.17 $Y=1.185 $X2=0
+ $Y2=0
cc_786 CI N_A_1340_412#_c_1643_n 0.0198126f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_787 N_CI_c_1077_n N_A_1340_412#_c_1643_n 0.00769627f $X=7.555 $Y=1.35 $X2=0
+ $Y2=0
cc_788 N_CI_c_1073_n N_VGND_c_1761_n 0.00687467f $X=7.63 $Y=1.185 $X2=0 $Y2=0
cc_789 N_CI_c_1075_n N_VGND_c_1761_n 0.00758746f $X=8.17 $Y=1.185 $X2=0 $Y2=0
cc_790 CI N_VGND_c_1761_n 0.0187477f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_791 N_CI_c_1078_n N_VGND_c_1761_n 0.00162178f $X=8.17 $Y=1.35 $X2=0 $Y2=0
cc_792 N_CI_c_1075_n N_VGND_c_1763_n 0.00541763f $X=8.17 $Y=1.185 $X2=0 $Y2=0
cc_793 N_CI_c_1073_n N_VGND_c_1766_n 0.00530923f $X=7.63 $Y=1.185 $X2=0 $Y2=0
cc_794 N_CI_c_1073_n N_VGND_c_1768_n 0.00525227f $X=7.63 $Y=1.185 $X2=0 $Y2=0
cc_795 N_CI_c_1075_n N_VGND_c_1768_n 0.0122211f $X=8.17 $Y=1.185 $X2=0 $Y2=0
cc_796 N_A_1571_367#_c_1144_n N_A_1758_87#_M1006_d 0.00353969f $X=9.495 $Y=2.63
+ $X2=0 $Y2=0
cc_797 N_A_1571_367#_M1015_g N_A_1758_87#_c_1258_n 0.00813478f $X=10.155
+ $Y=0.755 $X2=0 $Y2=0
cc_798 N_A_1571_367#_c_1140_n N_A_1758_87#_M1004_g 0.0285752f $X=10.155 $Y=1.665
+ $X2=0 $Y2=0
cc_799 N_A_1571_367#_c_1137_n N_A_1758_87#_c_1271_n 0.0188796f $X=8.385 $Y=0.43
+ $X2=0 $Y2=0
cc_800 N_A_1571_367#_c_1138_n N_A_1758_87#_c_1260_n 0.00574875f $X=8.107
+ $Y=1.815 $X2=0 $Y2=0
cc_801 N_A_1571_367#_M1015_g N_A_1758_87#_c_1261_n 0.0118215f $X=10.155 $Y=0.755
+ $X2=0 $Y2=0
cc_802 N_A_1571_367#_c_1137_n N_A_1758_87#_c_1262_n 0.0121486f $X=8.385 $Y=0.43
+ $X2=0 $Y2=0
cc_803 N_A_1571_367#_c_1144_n N_A_1758_87#_c_1263_n 0.0129403f $X=9.495 $Y=2.63
+ $X2=0 $Y2=0
cc_804 N_A_1571_367#_c_1148_n N_A_1758_87#_c_1263_n 0.0130013f $X=9.66 $Y=2.2
+ $X2=0 $Y2=0
cc_805 N_A_1571_367#_c_1149_n N_A_1758_87#_c_1263_n 0.00601723f $X=9.76 $Y=2.035
+ $X2=0 $Y2=0
cc_806 N_A_1571_367#_M1015_g N_A_1758_87#_c_1319_n 0.0124824f $X=10.155 $Y=0.755
+ $X2=0 $Y2=0
cc_807 N_A_1571_367#_M1015_g N_A_1758_87#_c_1320_n 0.00580117f $X=10.155
+ $Y=0.755 $X2=0 $Y2=0
cc_808 N_A_1571_367#_M1015_g N_A_1758_87#_c_1264_n 0.00327428f $X=10.155
+ $Y=0.755 $X2=0 $Y2=0
cc_809 N_A_1571_367#_c_1158_n N_A_1758_87#_c_1282_n 0.0188796f $X=8.385 $Y=0.88
+ $X2=0 $Y2=0
cc_810 N_A_1571_367#_M1015_g N_A_1758_87#_c_1266_n 0.00440228f $X=10.155
+ $Y=0.755 $X2=0 $Y2=0
cc_811 N_A_1571_367#_c_1140_n N_A_1758_87#_c_1266_n 0.00207542f $X=10.155
+ $Y=1.665 $X2=0 $Y2=0
cc_812 N_A_1571_367#_c_1145_n N_VPWR_c_1363_n 0.0277662f $X=7.995 $Y=1.98 $X2=0
+ $Y2=0
cc_813 N_A_1571_367#_c_1141_n N_VPWR_c_1364_n 0.00856616f $X=10.505 $Y=1.905
+ $X2=0 $Y2=0
cc_814 N_A_1571_367#_c_1141_n N_VPWR_c_1368_n 0.00475301f $X=10.505 $Y=1.905
+ $X2=0 $Y2=0
cc_815 N_A_1571_367#_c_1143_n N_VPWR_c_1368_n 0.019758f $X=7.995 $Y=2.9 $X2=0
+ $Y2=0
cc_816 N_A_1571_367#_c_1144_n N_VPWR_c_1368_n 0.00256113f $X=9.495 $Y=2.63 $X2=0
+ $Y2=0
cc_817 N_A_1571_367#_c_1147_n N_VPWR_c_1368_n 0.00474144f $X=8.107 $Y=2.63 $X2=0
+ $Y2=0
cc_818 N_A_1571_367#_M1023_d N_VPWR_c_1360_n 0.0023218f $X=7.855 $Y=1.835 $X2=0
+ $Y2=0
cc_819 N_A_1571_367#_c_1141_n N_VPWR_c_1360_n 0.00982677f $X=10.505 $Y=1.905
+ $X2=0 $Y2=0
cc_820 N_A_1571_367#_c_1143_n N_VPWR_c_1360_n 0.012508f $X=7.995 $Y=2.9 $X2=0
+ $Y2=0
cc_821 N_A_1571_367#_c_1144_n N_VPWR_c_1360_n 0.00589196f $X=9.495 $Y=2.63 $X2=0
+ $Y2=0
cc_822 N_A_1571_367#_c_1147_n N_VPWR_c_1360_n 0.00692171f $X=8.107 $Y=2.63 $X2=0
+ $Y2=0
cc_823 N_A_1571_367#_c_1144_n N_A_1708_411#_M1006_s 0.0107222f $X=9.495 $Y=2.63
+ $X2=0 $Y2=0
cc_824 N_A_1571_367#_c_1141_n N_A_1708_411#_c_1690_n 0.00325625f $X=10.505
+ $Y=1.905 $X2=0 $Y2=0
cc_825 N_A_1571_367#_c_1143_n N_A_1708_411#_c_1690_n 0.00882717f $X=7.995 $Y=2.9
+ $X2=0 $Y2=0
cc_826 N_A_1571_367#_c_1144_n N_A_1708_411#_c_1690_n 0.0577492f $X=9.495 $Y=2.63
+ $X2=0 $Y2=0
cc_827 N_A_1571_367#_c_1148_n N_A_1708_411#_c_1690_n 0.0370751f $X=9.66 $Y=2.2
+ $X2=0 $Y2=0
cc_828 N_A_1571_367#_M1015_g N_A_1708_411#_c_1687_n 0.0133662f $X=10.155
+ $Y=0.755 $X2=0 $Y2=0
cc_829 N_A_1571_367#_c_1139_n N_A_1708_411#_c_1687_n 0.0141552f $X=10.125
+ $Y=1.59 $X2=0 $Y2=0
cc_830 N_A_1571_367#_c_1140_n N_A_1708_411#_c_1687_n 0.00652329f $X=10.155
+ $Y=1.665 $X2=0 $Y2=0
cc_831 N_A_1571_367#_c_1139_n N_A_1708_411#_c_1688_n 0.0140843f $X=10.125
+ $Y=1.59 $X2=0 $Y2=0
cc_832 N_A_1571_367#_c_1140_n N_A_1708_411#_c_1688_n 0.00161689f $X=10.155
+ $Y=1.665 $X2=0 $Y2=0
cc_833 N_A_1571_367#_c_1141_n N_A_1708_411#_c_1702_n 0.0102083f $X=10.505
+ $Y=1.905 $X2=0 $Y2=0
cc_834 N_A_1571_367#_c_1148_n N_A_1708_411#_c_1702_n 0.0310174f $X=9.66 $Y=2.2
+ $X2=0 $Y2=0
cc_835 N_A_1571_367#_M1015_g N_A_1708_411#_c_1689_n 0.00398767f $X=10.155
+ $Y=0.755 $X2=0 $Y2=0
cc_836 N_A_1571_367#_c_1141_n N_A_1708_411#_c_1689_n 0.00115134f $X=10.505
+ $Y=1.905 $X2=0 $Y2=0
cc_837 N_A_1571_367#_c_1149_n N_A_1708_411#_c_1689_n 0.00652958f $X=9.76
+ $Y=2.035 $X2=0 $Y2=0
cc_838 N_A_1571_367#_c_1139_n N_A_1708_411#_c_1689_n 0.0239524f $X=10.125
+ $Y=1.59 $X2=0 $Y2=0
cc_839 N_A_1571_367#_c_1140_n N_A_1708_411#_c_1689_n 0.0154782f $X=10.155
+ $Y=1.665 $X2=0 $Y2=0
cc_840 N_A_1571_367#_c_1141_n N_A_1708_411#_c_1692_n 0.0124888f $X=10.505
+ $Y=1.905 $X2=0 $Y2=0
cc_841 N_A_1571_367#_c_1149_n N_A_1708_411#_c_1692_n 0.0310174f $X=9.76 $Y=2.035
+ $X2=0 $Y2=0
cc_842 N_A_1571_367#_c_1139_n N_A_1708_411#_c_1692_n 0.00193834f $X=10.125
+ $Y=1.59 $X2=0 $Y2=0
cc_843 N_A_1571_367#_c_1140_n N_A_1708_411#_c_1692_n 0.0097619f $X=10.155
+ $Y=1.665 $X2=0 $Y2=0
cc_844 N_A_1571_367#_c_1137_n N_VGND_c_1761_n 0.0521448f $X=8.385 $Y=0.43 $X2=0
+ $Y2=0
cc_845 N_A_1571_367#_M1015_g N_VGND_c_1762_n 7.86329e-19 $X=10.155 $Y=0.755
+ $X2=0 $Y2=0
cc_846 N_A_1571_367#_M1015_g N_VGND_c_1763_n 8.70381e-19 $X=10.155 $Y=0.755
+ $X2=0 $Y2=0
cc_847 N_A_1571_367#_c_1137_n N_VGND_c_1763_n 0.0200778f $X=8.385 $Y=0.43 $X2=0
+ $Y2=0
cc_848 N_A_1571_367#_M1012_d N_VGND_c_1768_n 0.0023218f $X=8.245 $Y=0.235 $X2=0
+ $Y2=0
cc_849 N_A_1571_367#_c_1137_n N_VGND_c_1768_n 0.0126785f $X=8.385 $Y=0.43 $X2=0
+ $Y2=0
cc_850 N_A_1758_87#_M1004_g N_VPWR_c_1364_n 0.00423847f $X=11.04 $Y=2.465 $X2=0
+ $Y2=0
cc_851 N_A_1758_87#_M1004_g N_VPWR_c_1369_n 0.00585385f $X=11.04 $Y=2.465 $X2=0
+ $Y2=0
cc_852 N_A_1758_87#_M1004_g N_VPWR_c_1360_n 0.0126087f $X=11.04 $Y=2.465 $X2=0
+ $Y2=0
cc_853 N_A_1758_87#_c_1261_n N_A_1708_411#_c_1696_n 0.0123205f $X=10.205 $Y=0.35
+ $X2=0 $Y2=0
cc_854 N_A_1758_87#_c_1258_n N_A_1708_411#_c_1687_n 3.64268e-19 $X=11.025
+ $Y=1.185 $X2=0 $Y2=0
cc_855 N_A_1758_87#_c_1261_n N_A_1708_411#_c_1687_n 0.00442932f $X=10.205
+ $Y=0.35 $X2=0 $Y2=0
cc_856 N_A_1758_87#_c_1331_p N_A_1708_411#_c_1687_n 0.0156651f $X=10.76 $Y=0.81
+ $X2=0 $Y2=0
cc_857 N_A_1758_87#_c_1320_n N_A_1708_411#_c_1687_n 0.010813f $X=10.375 $Y=0.81
+ $X2=0 $Y2=0
cc_858 N_A_1758_87#_c_1264_n N_A_1708_411#_c_1687_n 0.0137752f $X=10.865 $Y=1.35
+ $X2=0 $Y2=0
cc_859 N_A_1758_87#_c_1266_n N_A_1708_411#_c_1687_n 6.48798e-19 $X=11.04 $Y=1.35
+ $X2=0 $Y2=0
cc_860 N_A_1758_87#_M1004_g N_A_1708_411#_c_1702_n 9.22657e-19 $X=11.04 $Y=2.465
+ $X2=0 $Y2=0
cc_861 N_A_1758_87#_M1004_g N_A_1708_411#_c_1689_n 0.00352993f $X=11.04 $Y=2.465
+ $X2=0 $Y2=0
cc_862 N_A_1758_87#_c_1264_n N_A_1708_411#_c_1689_n 0.0187837f $X=10.865 $Y=1.35
+ $X2=0 $Y2=0
cc_863 N_A_1758_87#_c_1266_n N_A_1708_411#_c_1689_n 0.00257447f $X=11.04 $Y=1.35
+ $X2=0 $Y2=0
cc_864 N_A_1758_87#_c_1258_n N_SUM_c_1747_n 0.0045484f $X=11.025 $Y=1.185 $X2=0
+ $Y2=0
cc_865 N_A_1758_87#_c_1264_n N_SUM_c_1747_n 0.0377104f $X=10.865 $Y=1.35 $X2=0
+ $Y2=0
cc_866 N_A_1758_87#_c_1266_n N_SUM_c_1747_n 0.0210117f $X=11.04 $Y=1.35 $X2=0
+ $Y2=0
cc_867 N_A_1758_87#_c_1319_n N_VGND_M1015_d 0.00414649f $X=10.29 $Y=0.725 $X2=0
+ $Y2=0
cc_868 N_A_1758_87#_c_1331_p N_VGND_M1015_d 0.0187064f $X=10.76 $Y=0.81 $X2=0
+ $Y2=0
cc_869 N_A_1758_87#_c_1320_n N_VGND_M1015_d 9.63726e-19 $X=10.375 $Y=0.81 $X2=0
+ $Y2=0
cc_870 N_A_1758_87#_c_1264_n N_VGND_M1015_d 0.00296615f $X=10.865 $Y=1.35 $X2=0
+ $Y2=0
cc_871 N_A_1758_87#_c_1258_n N_VGND_c_1762_n 0.00932188f $X=11.025 $Y=1.185
+ $X2=0 $Y2=0
cc_872 N_A_1758_87#_c_1261_n N_VGND_c_1762_n 0.0114856f $X=10.205 $Y=0.35 $X2=0
+ $Y2=0
cc_873 N_A_1758_87#_c_1319_n N_VGND_c_1762_n 0.00644995f $X=10.29 $Y=0.725 $X2=0
+ $Y2=0
cc_874 N_A_1758_87#_c_1331_p N_VGND_c_1762_n 0.019197f $X=10.76 $Y=0.81 $X2=0
+ $Y2=0
cc_875 N_A_1758_87#_c_1266_n N_VGND_c_1762_n 4.02835e-19 $X=11.04 $Y=1.35 $X2=0
+ $Y2=0
cc_876 N_A_1758_87#_c_1261_n N_VGND_c_1763_n 0.0786461f $X=10.205 $Y=0.35 $X2=0
+ $Y2=0
cc_877 N_A_1758_87#_c_1262_n N_VGND_c_1763_n 0.0222501f $X=9.095 $Y=0.35 $X2=0
+ $Y2=0
cc_878 N_A_1758_87#_c_1331_p N_VGND_c_1763_n 0.00338075f $X=10.76 $Y=0.81 $X2=0
+ $Y2=0
cc_879 N_A_1758_87#_c_1258_n N_VGND_c_1767_n 0.00560773f $X=11.025 $Y=1.185
+ $X2=0 $Y2=0
cc_880 N_A_1758_87#_c_1331_p N_VGND_c_1767_n 0.00133214f $X=10.76 $Y=0.81 $X2=0
+ $Y2=0
cc_881 N_A_1758_87#_c_1258_n N_VGND_c_1768_n 0.0124095f $X=11.025 $Y=1.185 $X2=0
+ $Y2=0
cc_882 N_A_1758_87#_c_1261_n N_VGND_c_1768_n 0.04804f $X=10.205 $Y=0.35 $X2=0
+ $Y2=0
cc_883 N_A_1758_87#_c_1262_n N_VGND_c_1768_n 0.0127687f $X=9.095 $Y=0.35 $X2=0
+ $Y2=0
cc_884 N_A_1758_87#_c_1331_p N_VGND_c_1768_n 0.0105003f $X=10.76 $Y=0.81 $X2=0
+ $Y2=0
cc_885 N_VPWR_c_1361_n N_A_247_367#_c_1468_n 0.0585555f $X=0.82 $Y=2.125 $X2=0
+ $Y2=0
cc_886 N_VPWR_c_1365_n N_A_247_367#_c_1464_n 0.134924f $X=4.565 $Y=3.33 $X2=0
+ $Y2=0
cc_887 N_VPWR_c_1360_n N_A_247_367#_c_1464_n 0.0780561f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_888 N_VPWR_c_1361_n N_A_247_367#_c_1465_n 0.0120187f $X=0.82 $Y=2.125 $X2=0
+ $Y2=0
cc_889 N_VPWR_c_1365_n N_A_247_367#_c_1465_n 0.0222162f $X=4.565 $Y=3.33 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_1360_n N_A_247_367#_c_1465_n 0.0127633f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_891 N_VPWR_c_1362_n N_A_1034_380#_c_1533_n 0.0582556f $X=4.73 $Y=1.94 $X2=0
+ $Y2=0
cc_892 N_VPWR_c_1367_n N_A_1034_380#_c_1534_n 0.0117167f $X=7.32 $Y=3.33 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_1360_n N_A_1034_380#_c_1534_n 0.0116437f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_894 N_VPWR_c_1362_n N_A_1034_380#_c_1532_n 0.00448828f $X=4.73 $Y=1.94 $X2=0
+ $Y2=0
cc_895 N_VPWR_c_1367_n N_COUT_N_c_1586_n 0.0117826f $X=7.32 $Y=3.33 $X2=0 $Y2=0
cc_896 N_VPWR_c_1360_n N_COUT_N_c_1586_n 0.011666f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_897 N_VPWR_c_1363_n N_A_1340_412#_c_1644_n 0.0670642f $X=7.485 $Y=2.025 $X2=0
+ $Y2=0
cc_898 N_VPWR_c_1367_n N_A_1340_412#_c_1644_n 0.00890876f $X=7.32 $Y=3.33 $X2=0
+ $Y2=0
cc_899 N_VPWR_c_1360_n N_A_1340_412#_c_1644_n 0.00882062f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_900 N_VPWR_c_1363_n N_A_1340_412#_c_1642_n 0.00869681f $X=7.485 $Y=2.025
+ $X2=0 $Y2=0
cc_901 N_VPWR_c_1360_n N_A_1708_411#_M1006_s 0.00272517f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_902 N_VPWR_c_1364_n N_A_1708_411#_c_1690_n 0.0119478f $X=10.825 $Y=2.45 $X2=0
+ $Y2=0
cc_903 N_VPWR_c_1368_n N_A_1708_411#_c_1690_n 0.118614f $X=10.66 $Y=3.33 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_1360_n N_A_1708_411#_c_1690_n 0.0725277f $X=11.28 $Y=3.33 $X2=0
+ $Y2=0
cc_905 N_VPWR_c_1364_n N_A_1708_411#_c_1702_n 0.0392818f $X=10.825 $Y=2.45 $X2=0
+ $Y2=0
cc_906 N_VPWR_c_1360_n N_SUM_M1004_d 0.00358712f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_907 N_VPWR_c_1369_n N_SUM_c_1747_n 0.0169002f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_908 N_VPWR_c_1360_n N_SUM_c_1747_n 0.0101763f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_909 N_A_1034_380#_c_1533_n N_COUT_N_c_1586_n 0.0183106f $X=5.31 $Y=2.045
+ $X2=0 $Y2=0
cc_910 N_A_1034_380#_c_1534_n N_COUT_N_c_1586_n 0.0183106f $X=5.31 $Y=2.4 $X2=0
+ $Y2=0
cc_911 N_A_1034_380#_c_1532_n N_COUT_N_c_1584_n 0.00890906f $X=5.31 $Y=1.88
+ $X2=0 $Y2=0
cc_912 N_A_1034_380#_c_1539_n N_VGND_M1011_d 0.00269749f $X=5.795 $Y=0.545 $X2=0
+ $Y2=0
cc_913 N_A_1034_380#_c_1541_n N_VGND_M1011_d 0.00578475f $X=5.475 $Y=0.545 $X2=0
+ $Y2=0
cc_914 N_A_1034_380#_c_1532_n N_VGND_M1011_d 0.00706743f $X=5.31 $Y=1.88 $X2=0
+ $Y2=0
cc_915 N_A_1034_380#_c_1541_n N_VGND_c_1760_n 0.0118278f $X=5.475 $Y=0.545 $X2=0
+ $Y2=0
cc_916 N_A_1034_380#_c_1532_n N_VGND_c_1760_n 0.0225689f $X=5.31 $Y=1.88 $X2=0
+ $Y2=0
cc_917 N_A_1034_380#_c_1539_n N_VGND_c_1766_n 0.00786192f $X=5.795 $Y=0.545
+ $X2=0 $Y2=0
cc_918 N_A_1034_380#_c_1541_n N_VGND_c_1766_n 0.00506241f $X=5.475 $Y=0.545
+ $X2=0 $Y2=0
cc_919 N_A_1034_380#_c_1547_n N_VGND_c_1766_n 0.0171921f $X=5.96 $Y=0.445 $X2=0
+ $Y2=0
cc_920 N_A_1034_380#_c_1539_n N_VGND_c_1768_n 0.00983286f $X=5.795 $Y=0.545
+ $X2=0 $Y2=0
cc_921 N_A_1034_380#_c_1541_n N_VGND_c_1768_n 0.00584745f $X=5.475 $Y=0.545
+ $X2=0 $Y2=0
cc_922 N_A_1034_380#_c_1547_n N_VGND_c_1768_n 0.0122489f $X=5.96 $Y=0.445 $X2=0
+ $Y2=0
cc_923 N_COUT_N_c_1586_n N_A_1340_412#_c_1644_n 0.0218559f $X=6.04 $Y=2.205
+ $X2=0 $Y2=0
cc_924 N_COUT_N_c_1584_n N_A_1340_412#_c_1642_n 0.00190078f $X=6.04 $Y=2.04
+ $X2=0 $Y2=0
cc_925 COUT_N N_A_1340_412#_c_1643_n 0.011848f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_926 COUT_N N_VGND_c_1766_n 0.0207394f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_927 COUT_N N_VGND_c_1768_n 0.0125622f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_928 N_A_1340_412#_c_1643_n N_VGND_c_1761_n 0.0351126f $X=7.31 $Y=0.43 $X2=0
+ $Y2=0
cc_929 N_A_1340_412#_c_1643_n N_VGND_c_1766_n 0.0164235f $X=7.31 $Y=0.43 $X2=0
+ $Y2=0
cc_930 N_A_1340_412#_c_1643_n N_VGND_c_1768_n 0.0095959f $X=7.31 $Y=0.43 $X2=0
+ $Y2=0
cc_931 N_A_1708_411#_c_1689_n N_SUM_c_1747_n 0.0138846f $X=10.392 $Y=1.935 $X2=0
+ $Y2=0
cc_932 N_A_1708_411#_c_1687_n N_VGND_M1015_d 0.00193196f $X=10.41 $Y=1.16 $X2=0
+ $Y2=0
cc_933 N_SUM_c_1747_n N_VGND_c_1767_n 0.0173887f $X=11.24 $Y=0.43 $X2=0 $Y2=0
cc_934 N_SUM_M1017_d N_VGND_c_1768_n 0.0042346f $X=11.1 $Y=0.235 $X2=0 $Y2=0
cc_935 N_SUM_c_1747_n N_VGND_c_1768_n 0.0101709f $X=11.24 $Y=0.43 $X2=0 $Y2=0
