* File: sky130_fd_sc_lp__or2b_lp.spice
* Created: Wed Sep  2 10:30:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2b_lp.pex.spice"
.subckt sky130_fd_sc_lp__or2b_lp  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1006 A_117_57# N_B_N_M1006_g N_A_30_57#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B_N_M1002_g A_117_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1007 A_275_57# N_A_30_57#_M1007_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_290_409#_M1008_d N_A_30_57#_M1008_g A_275_57# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 A_439_57# N_A_M1001_g N_A_290_409#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g A_439_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1003 A_597_57# N_A_290_409#_M1003_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_290_409#_M1004_g A_597_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_B_N_M1011_g N_A_30_57#_M1011_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1005 A_397_409# N_A_30_57#_M1005_g N_A_290_409#_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g A_397_409# VPB PHIGHVT L=0.25 W=1 AD=0.2825
+ AS=0.12 PD=1.565 PS=1.24 NRD=56.145 NRS=12.7853 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1000 N_X_M1000_d N_A_290_409#_M1000_g N_VPWR_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.2825 PD=2.57 PS=1.565 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__or2b_lp.pxi.spice"
*
.ends
*
*
