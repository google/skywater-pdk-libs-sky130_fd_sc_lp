# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__buf_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__buf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.945000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.180000 0.880000 1.385000 ;
        RECT 0.095000 1.385000 1.345000 1.575000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.865000 0.305000 2.110000 1.045000 ;
        RECT 1.865000 1.045000 5.190000 1.225000 ;
        RECT 1.865000 1.745000 5.190000 1.925000 ;
        RECT 1.865000 1.925000 2.105000 2.980000 ;
        RECT 2.705000 1.925000 2.975000 2.980000 ;
        RECT 2.710000 0.305000 2.965000 1.045000 ;
        RECT 3.570000 0.305000 3.830000 1.045000 ;
        RECT 3.570000 1.925000 3.830000 2.980000 ;
        RECT 4.430000 0.305000 4.685000 1.045000 ;
        RECT 4.430000 1.925000 4.690000 2.980000 ;
        RECT 4.910000 1.225000 5.190000 1.745000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
        RECT 0.560000  0.085000 0.820000 0.670000 ;
        RECT 1.420000  0.085000 1.695000 0.875000 ;
        RECT 2.280000  0.085000 2.540000 0.875000 ;
        RECT 3.135000  0.085000 3.400000 0.875000 ;
        RECT 4.000000  0.085000 4.260000 0.875000 ;
        RECT 4.855000  0.085000 5.155000 0.875000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 5.280000 3.415000 ;
        RECT 0.560000 2.095000 0.820000 3.245000 ;
        RECT 1.420000 2.095000 1.695000 3.245000 ;
        RECT 2.275000 2.095000 2.535000 3.245000 ;
        RECT 3.145000 2.095000 3.400000 3.245000 ;
        RECT 4.000000 2.095000 4.260000 3.245000 ;
        RECT 4.860000 2.095000 5.095000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.305000 0.390000 0.840000 ;
      RECT 0.095000 0.840000 1.250000 1.010000 ;
      RECT 0.095000 1.745000 1.695000 1.925000 ;
      RECT 0.095000 1.925000 0.390000 2.980000 ;
      RECT 0.990000 0.305000 1.250000 0.840000 ;
      RECT 0.990000 1.925000 1.250000 2.980000 ;
      RECT 1.050000 1.010000 1.250000 1.045000 ;
      RECT 1.050000 1.045000 1.695000 1.215000 ;
      RECT 1.525000 1.215000 1.695000 1.395000 ;
      RECT 1.525000 1.395000 4.740000 1.575000 ;
      RECT 1.525000 1.575000 1.695000 1.745000 ;
  END
END sky130_fd_sc_lp__buf_8
