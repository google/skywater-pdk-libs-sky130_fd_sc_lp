* File: sky130_fd_sc_lp__a41o_2.pex.spice
* Created: Fri Aug 28 10:02:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41O_2%A_90_53# 1 2 3 10 12 15 17 21 24 26 27 34 37
+ 39 40 42 44 48 50 51 58
r91 46 48 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=4.385 $Y=0.995
+ $X2=4.385 $Y2=0.42
r92 45 50 5.01601 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=2.08 $Y=1.08
+ $X2=1.792 $Y2=1.08
r93 44 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.22 $Y=1.08
+ $X2=4.385 $Y2=0.995
r94 44 45 139.615 $w=1.68e-07 $l=2.14e-06 $layer=LI1_cond $X=4.22 $Y=1.08
+ $X2=2.08 $Y2=1.08
r95 40 52 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=1.945 $Y=2.01
+ $X2=1.75 $Y2=2.01
r96 40 42 34.5733 $w=2.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.945 $Y=2.1
+ $X2=1.945 $Y2=2.91
r97 39 52 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.75 $Y=1.92 $X2=1.75
+ $Y2=2.01
r98 38 51 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=1.75 $Y=1.675
+ $X2=1.67 $Y2=1.51
r99 38 39 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.75 $Y=1.675
+ $X2=1.75 $Y2=1.92
r100 37 51 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=1.345
+ $X2=1.67 $Y2=1.51
r101 36 50 2.15548 $w=4.52e-07 $l=1.58915e-07 $layer=LI1_cond $X=1.67 $Y=1.165
+ $X2=1.792 $Y2=1.08
r102 36 37 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.67 $Y=1.165
+ $X2=1.67 $Y2=1.345
r103 32 50 2.15548 $w=4.52e-07 $l=8.5e-08 $layer=LI1_cond $X=1.792 $Y=0.995
+ $X2=1.792 $Y2=1.08
r104 32 34 11.9608 $w=5.73e-07 $l=5.75e-07 $layer=LI1_cond $X=1.792 $Y=0.995
+ $X2=1.792 $Y2=0.42
r105 30 60 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.077 $Y=1.51
+ $X2=1.077 $Y2=1.675
r106 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.51 $X2=1.11 $Y2=1.51
r107 27 51 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.51
+ $X2=1.67 $Y2=1.51
r108 27 29 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=1.505 $Y=1.51
+ $X2=1.11 $Y2=1.51
r109 24 60 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.955 $Y=2.465
+ $X2=0.955 $Y2=1.675
r110 21 58 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.955 $Y=0.815
+ $X2=0.955 $Y2=1.345
r111 18 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.6 $Y=1.42
+ $X2=0.525 $Y2=1.42
r112 17 30 12.6719 $w=3.95e-07 $l=9e-08 $layer=POLY_cond $X=1.077 $Y=1.42
+ $X2=1.077 $Y2=1.51
r113 17 58 32.8921 $w=3.95e-07 $l=7.5e-08 $layer=POLY_cond $X=1.077 $Y=1.42
+ $X2=1.077 $Y2=1.345
r114 17 18 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.88 $Y=1.42
+ $X2=0.6 $Y2=1.42
r115 13 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.525 $Y=1.495
+ $X2=0.525 $Y2=1.42
r116 13 15 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.525 $Y=1.495
+ $X2=0.525 $Y2=2.465
r117 10 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.525 $Y=1.345
+ $X2=0.525 $Y2=1.42
r118 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.525 $Y=1.345
+ $X2=0.525 $Y2=0.815
r119 3 40 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.835 $X2=1.975 $Y2=2.085
r120 3 42 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.835 $X2=1.975 $Y2=2.91
r121 2 48 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=4.245
+ $Y=0.245 $X2=4.385 $Y2=0.42
r122 1 34 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=1.85
+ $Y=0.245 $X2=1.975 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_2%B1 3 7 9 12 13
r33 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.1 $Y=1.51 $X2=2.1
+ $Y2=1.675
r34 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.1 $Y=1.51 $X2=2.1
+ $Y2=1.345
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.1
+ $Y=1.51 $X2=2.1 $Y2=1.51
r36 9 13 5.95429 $w=2.98e-07 $l=1.55e-07 $layer=LI1_cond $X=2.155 $Y=1.665
+ $X2=2.155 $Y2=1.51
r37 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.19 $Y=2.465
+ $X2=2.19 $Y2=1.675
r38 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.19 $Y=0.665
+ $X2=2.19 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_2%A4 3 7 9 12 13
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=1.51
+ $X2=2.64 $Y2=1.675
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=1.51
+ $X2=2.64 $Y2=1.345
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.64
+ $Y=1.51 $X2=2.64 $Y2=1.51
r39 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.51
r40 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.73 $Y=0.665
+ $X2=2.73 $Y2=1.345
r41 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.62 $Y=2.465
+ $X2=2.62 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_2%A3 3 7 9 12 13
c36 13 0 1.93464e-19 $X=3.18 $Y=1.51
r37 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.18 $Y=1.51
+ $X2=3.18 $Y2=1.675
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.18 $Y=1.51
+ $X2=3.18 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.51 $X2=3.18 $Y2=1.51
r40 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.14 $Y=1.665
+ $X2=3.14 $Y2=1.51
r41 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.09 $Y=2.465
+ $X2=3.09 $Y2=1.675
r42 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.09 $Y=0.665
+ $X2=3.09 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_2%A2 3 7 9 10 14
c35 14 0 1.50241e-19 $X=3.72 $Y=1.51
c36 7 0 1.93464e-19 $X=3.74 $Y=2.465
r37 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=1.51
+ $X2=3.72 $Y2=1.675
r38 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=1.51
+ $X2=3.72 $Y2=1.345
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.72
+ $Y=1.51 $X2=3.72 $Y2=1.51
r40 10 15 10.2439 $w=4.03e-07 $l=3.6e-07 $layer=LI1_cond $X=4.08 $Y=1.547
+ $X2=3.72 $Y2=1.547
r41 9 15 3.41465 $w=4.03e-07 $l=1.2e-07 $layer=LI1_cond $X=3.6 $Y=1.547 $X2=3.72
+ $Y2=1.547
r42 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.74 $Y=2.465
+ $X2=3.74 $Y2=1.675
r43 3 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.63 $Y=0.665
+ $X2=3.63 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_2%A1 3 7 9 14 15
c24 15 0 1.50241e-19 $X=4.51 $Y=1.46
r25 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.51
+ $Y=1.46 $X2=4.51 $Y2=1.46
r26 11 14 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.17 $Y=1.46
+ $X2=4.51 $Y2=1.46
r27 9 15 6.47263 $w=3.63e-07 $l=2.05e-07 $layer=LI1_cond $X=4.527 $Y=1.665
+ $X2=4.527 $Y2=1.46
r28 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.17 $Y=1.625
+ $X2=4.17 $Y2=1.46
r29 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.17 $Y=1.625 $X2=4.17
+ $Y2=2.465
r30 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.17 $Y=1.295
+ $X2=4.17 $Y2=1.46
r31 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=4.17 $Y=1.295 $X2=4.17
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_2%VPWR 1 2 3 4 13 15 21 27 31 34 35 37 38 39 41
+ 57 58 64
r67 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r68 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r70 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r71 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r72 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r73 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r74 49 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r75 48 51 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r76 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r77 46 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r78 46 48 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 45 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r80 45 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r82 42 61 4.27611 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=3.33
+ $X2=0.215 $Y2=3.33
r83 42 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=3.33
+ $X2=0.72 $Y2=3.33
r84 41 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r85 41 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 39 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 39 49 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r88 37 54 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.79 $Y=3.33 $X2=3.6
+ $Y2=3.33
r89 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=3.33
+ $X2=3.955 $Y2=3.33
r90 36 57 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=3.33
+ $X2=3.955 $Y2=3.33
r92 34 51 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=3.33 $X2=2.64
+ $Y2=3.33
r93 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=2.855 $Y2=3.33
r94 33 54 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.02 $Y=3.33 $X2=3.6
+ $Y2=3.33
r95 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=2.855 $Y2=3.33
r96 29 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=3.245
+ $X2=3.955 $Y2=3.33
r97 29 31 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=3.955 $Y=3.245
+ $X2=3.955 $Y2=2.385
r98 25 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=3.245
+ $X2=2.855 $Y2=3.33
r99 25 27 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.855 $Y=3.245
+ $X2=2.855 $Y2=2.385
r100 21 24 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=1.17 $Y=2.01
+ $X2=1.17 $Y2=2.95
r101 19 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r102 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.95
r103 15 18 39.2235 $w=2.83e-07 $l=9.7e-07 $layer=LI1_cond $X=0.287 $Y=1.98
+ $X2=0.287 $Y2=2.95
r104 13 61 3.12256 $w=2.85e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.287 $Y=3.245
+ $X2=0.215 $Y2=3.33
r105 13 18 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.287 $Y=3.245
+ $X2=0.287 $Y2=2.95
r106 4 31 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=3.815
+ $Y=1.835 $X2=3.955 $Y2=2.385
r107 3 27 300 $w=1.7e-07 $l=6.249e-07 $layer=licon1_PDIFF $count=2 $X=2.695
+ $Y=1.835 $X2=2.855 $Y2=2.385
r108 2 24 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.95
r109 2 21 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.01
r110 1 18 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=2.95
r111 1 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_2%X 1 2 7 8 9 10 11 12 13
r16 13 37 5.63961 $w=2.33e-07 $l=1.15e-07 $layer=LI1_cond $X=0.717 $Y=2.775
+ $X2=0.717 $Y2=2.66
r17 12 37 12.5052 $w=2.33e-07 $l=2.55e-07 $layer=LI1_cond $X=0.717 $Y=2.405
+ $X2=0.717 $Y2=2.66
r18 11 12 20.8421 $w=2.33e-07 $l=4.25e-07 $layer=LI1_cond $X=0.717 $Y=1.98
+ $X2=0.717 $Y2=2.405
r19 10 11 15.4476 $w=2.33e-07 $l=3.15e-07 $layer=LI1_cond $X=0.717 $Y=1.665
+ $X2=0.717 $Y2=1.98
r20 9 10 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.717 $Y=1.295
+ $X2=0.717 $Y2=1.665
r21 8 9 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.717 $Y=0.925
+ $X2=0.717 $Y2=1.295
r22 7 8 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.717 $Y=0.555
+ $X2=0.717 $Y2=0.925
r23 2 37 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.74 $Y2=2.66
r24 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.74 $Y2=1.98
r25 1 7 91 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=2 $X=0.6
+ $Y=0.395 $X2=0.74 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_2%A_453_367# 1 2 3 10 12 14 18 20 22 24 29
r37 22 31 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=4.42 $Y=2.1 $X2=4.42
+ $Y2=2.01
r38 22 24 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=4.42 $Y=2.1 $X2=4.42
+ $Y2=2.91
r39 21 29 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=2.01
+ $X2=3.425 $Y2=2.01
r40 20 31 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=4.29 $Y=2.01 $X2=4.42
+ $Y2=2.01
r41 20 21 43.1313 $w=1.78e-07 $l=7e-07 $layer=LI1_cond $X=4.29 $Y=2.01 $X2=3.59
+ $Y2=2.01
r42 16 29 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.425 $Y=2.1 $X2=3.425
+ $Y2=2.01
r43 16 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.425 $Y=2.1
+ $X2=3.425 $Y2=2.47
r44 15 27 3.79804 $w=1.8e-07 $l=1.1e-07 $layer=LI1_cond $X=2.52 $Y=2.01 $X2=2.41
+ $Y2=2.01
r45 14 29 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=2.01
+ $X2=3.425 $Y2=2.01
r46 14 15 45.596 $w=1.78e-07 $l=7.4e-07 $layer=LI1_cond $X=3.26 $Y=2.01 $X2=2.52
+ $Y2=2.01
r47 10 27 3.10749 $w=2.2e-07 $l=9e-08 $layer=LI1_cond $X=2.41 $Y=2.1 $X2=2.41
+ $Y2=2.01
r48 10 12 42.4309 $w=2.18e-07 $l=8.1e-07 $layer=LI1_cond $X=2.41 $Y=2.1 $X2=2.41
+ $Y2=2.91
r49 3 31 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=1.835 $X2=4.385 $Y2=2.095
r50 3 24 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=1.835 $X2=4.385 $Y2=2.91
r51 2 29 600 $w=1.7e-07 $l=3.38231e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.835 $X2=3.425 $Y2=2.015
r52 2 18 300 $w=1.7e-07 $l=7.53873e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.835 $X2=3.425 $Y2=2.47
r53 1 27 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.265
+ $Y=1.835 $X2=2.405 $Y2=2.095
r54 1 12 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.265
+ $Y=1.835 $X2=2.405 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_2%VGND 1 2 3 10 12 16 20 23 24 25 27 40 41 47
r51 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r54 38 41 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r55 37 40 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r56 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r57 35 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r58 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r59 32 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.17
+ $Y2=0
r60 32 34 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=2.16
+ $Y2=0
r61 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r62 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r63 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r64 28 44 4.27611 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r65 28 30 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r66 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.17
+ $Y2=0
r67 27 30 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.72
+ $Y2=0
r68 25 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r69 25 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r70 23 34 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.16
+ $Y2=0
r71 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.46
+ $Y2=0
r72 22 37 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.64
+ $Y2=0
r73 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.46
+ $Y2=0
r74 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0
r75 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.46 $Y=0.085
+ $X2=2.46 $Y2=0.37
r76 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0
r77 14 16 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.54
r78 10 44 3.12256 $w=2.85e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.287 $Y=0.085
+ $X2=0.215 $Y2=0
r79 10 12 18.3987 $w=2.83e-07 $l=4.55e-07 $layer=LI1_cond $X=0.287 $Y=0.085
+ $X2=0.287 $Y2=0.54
r80 3 20 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=2.265
+ $Y=0.245 $X2=2.46 $Y2=0.37
r81 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.03
+ $Y=0.395 $X2=1.17 $Y2=0.54
r82 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.185
+ $Y=0.395 $X2=0.31 $Y2=0.54
.ends

