* NGSPICE file created from sky130_fd_sc_lp__and4_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and4_0 A B C D VGND VNB VPB VPWR X
M1000 VPWR B a_84_58# VPB phighvt w=420000u l=150000u
+  ad=5.959e+11p pd=5.52e+06u as=2.352e+11p ps=2.8e+06u
M1001 X a_84_58# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1002 a_167_58# A a_84_58# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1003 a_239_58# B a_167_58# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 VPWR D a_84_58# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_84_58# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.604e+11p ps=2.08e+06u
M1006 a_311_58# C a_239_58# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 a_84_58# C VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND D a_311_58# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_84_58# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

