* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
X0 VGND a_663_481# a_849_419# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VPWR GATE_N a_242_130# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_771_481# a_849_419# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR a_663_481# a_849_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_669_47# a_242_130# a_663_481# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_849_419# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_663_481# a_242_130# a_771_481# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_57_130# a_591_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VGND GATE_N a_242_130# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_591_481# a_349_481# a_663_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_349_481# a_242_130# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_663_481# a_349_481# a_849_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 Q a_849_419# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_849_47# a_849_419# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 Q a_849_419# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR a_849_419# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_349_481# a_242_130# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_57_130# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_57_130# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 VGND a_57_130# a_669_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
