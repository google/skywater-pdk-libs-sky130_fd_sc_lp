* File: sky130_fd_sc_lp__o2bb2ai_m.pxi.spice
* Created: Fri Aug 28 11:13:14 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2AI_M%A1_N N_A1_N_M1008_g N_A1_N_M1006_g A1_N A1_N
+ A1_N A1_N A1_N N_A1_N_c_74_n N_A1_N_c_75_n N_A1_N_c_76_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_M%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_M%A2_N N_A2_N_M1000_g N_A2_N_M1004_g
+ N_A2_N_c_105_n N_A2_N_c_106_n A2_N A2_N A2_N A2_N N_A2_N_c_108_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_M%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_M%A_110_535# N_A_110_535#_M1000_d
+ N_A_110_535#_M1008_d N_A_110_535#_M1007_g N_A_110_535#_c_151_n
+ N_A_110_535#_c_152_n N_A_110_535#_c_153_n N_A_110_535#_M1003_g
+ N_A_110_535#_c_154_n N_A_110_535#_c_159_n N_A_110_535#_c_160_n
+ N_A_110_535#_c_161_n N_A_110_535#_c_162_n N_A_110_535#_c_163_n
+ N_A_110_535#_c_155_n N_A_110_535#_c_156_n N_A_110_535#_c_165_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_M%A_110_535#
x_PM_SKY130_FD_SC_LP__O2BB2AI_M%B2 N_B2_M1002_g N_B2_M1009_g B2 B2 B2
+ N_B2_c_224_n PM_SKY130_FD_SC_LP__O2BB2AI_M%B2
x_PM_SKY130_FD_SC_LP__O2BB2AI_M%B1 N_B1_M1005_g N_B1_c_267_n N_B1_c_268_n
+ N_B1_M1001_g N_B1_c_269_n B1 B1 B1 B1 N_B1_c_265_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_M%B1
x_PM_SKY130_FD_SC_LP__O2BB2AI_M%VPWR N_VPWR_M1008_s N_VPWR_M1004_d
+ N_VPWR_M1005_d N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n
+ N_VPWR_c_304_n N_VPWR_c_305_n VPWR N_VPWR_c_306_n N_VPWR_c_307_n
+ N_VPWR_c_299_n N_VPWR_c_309_n PM_SKY130_FD_SC_LP__O2BB2AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2AI_M%Y N_Y_M1003_s N_Y_M1007_d N_Y_c_345_n
+ N_Y_c_347_n N_Y_c_350_n N_Y_c_348_n Y PM_SKY130_FD_SC_LP__O2BB2AI_M%Y
x_PM_SKY130_FD_SC_LP__O2BB2AI_M%VGND N_VGND_M1006_s N_VGND_M1009_d
+ N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n VGND N_VGND_c_393_n
+ N_VGND_c_394_n N_VGND_c_395_n N_VGND_c_396_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_M%VGND
x_PM_SKY130_FD_SC_LP__O2BB2AI_M%A_410_78# N_A_410_78#_M1003_d
+ N_A_410_78#_M1001_d N_A_410_78#_c_426_n N_A_410_78#_c_427_n
+ N_A_410_78#_c_428_n N_A_410_78#_c_429_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_M%A_410_78#
cc_1 VNB N_A1_N_M1008_g 0.0015916f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_2 VNB N_A1_N_M1006_g 0.0191936f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.615
cc_3 VNB N_A1_N_c_74_n 0.102907f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_4 VNB N_A1_N_c_75_n 0.00125626f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_5 VNB N_A1_N_c_76_n 0.00668735f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.055
cc_6 VNB N_A2_N_c_105_n 0.0201446f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB N_A2_N_c_106_n 0.040685f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB A2_N 0.01103f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_A2_N_c_108_n 0.0155379f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_10 VNB N_A_110_535#_c_151_n 0.0399299f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_11 VNB N_A_110_535#_c_152_n 0.0107331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_110_535#_c_153_n 0.0207094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_110_535#_c_154_n 0.0283527f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.12
cc_14 VNB N_A_110_535#_c_155_n 0.00834713f $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=1.665
cc_15 VNB N_A_110_535#_c_156_n 0.00984246f $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=0.925
cc_16 VNB N_B2_M1009_g 0.0373931f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.615
cc_17 VNB B2 0.00358854f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_18 VNB N_B2_c_224_n 0.0491397f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_19 VNB N_B1_M1001_g 0.0667804f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_20 VNB B1 0.0220137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_c_265_n 0.0097119f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.625
cc_22 VNB N_VPWR_c_299_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_345_n 0.00806238f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_24 VNB N_VGND_c_390_n 0.0125358f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.615
cc_25 VNB N_VGND_c_391_n 0.0228168f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_26 VNB N_VGND_c_392_n 0.00986829f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_27 VNB N_VGND_c_393_n 0.0597515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_394_n 0.0211404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_395_n 0.233731f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_30 VNB N_VGND_c_396_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_410_78#_c_426_n 8.22023e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_32 VNB N_A_410_78#_c_427_n 0.0235839f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_33 VNB N_A_410_78#_c_428_n 0.00313384f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_34 VNB N_A_410_78#_c_429_n 0.00224906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_A1_N_M1008_g 0.0743471f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_36 VPB N_A1_N_c_75_n 0.0428129f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_37 VPB N_A2_N_M1004_g 0.0535065f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.615
cc_38 VPB N_A2_N_c_106_n 0.00570137f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_39 VPB A2_N 0.00918862f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_40 VPB N_A_110_535#_M1007_g 0.0204748f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_41 VPB N_A_110_535#_c_154_n 0.00984305f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.12
cc_42 VPB N_A_110_535#_c_159_n 0.0239502f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_43 VPB N_A_110_535#_c_160_n 0.0158061f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_44 VPB N_A_110_535#_c_161_n 0.00316203f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.055
cc_45 VPB N_A_110_535#_c_162_n 0.0106325f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_46 VPB N_A_110_535#_c_163_n 0.00437533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_110_535#_c_156_n 0.00133833f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_48 VPB N_A_110_535#_c_165_n 0.0189675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B2_M1002_g 0.0448034f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_50 VPB B2 0.00387023f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_51 VPB N_B2_c_224_n 0.0456403f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_52 VPB N_B1_M1005_g 0.0333071f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_53 VPB N_B1_c_267_n 0.0595866f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.955
cc_54 VPB N_B1_c_268_n 0.00732581f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.615
cc_55 VPB N_B1_c_269_n 0.0423859f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_56 VPB B1 0.0403325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_B1_c_265_n 0.00914979f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.625
cc_58 VPB N_VPWR_c_300_n 0.0103338f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_59 VPB N_VPWR_c_301_n 0.0137479f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_60 VPB N_VPWR_c_302_n 0.00286965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_303_n 0.0128467f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_62 VPB N_VPWR_c_304_n 0.0277597f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.625
cc_63 VPB N_VPWR_c_305_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.055
cc_64 VPB N_VPWR_c_306_n 0.0138618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_307_n 0.0258507f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_299_n 0.0606342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_309_n 0.00522083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_Y_c_345_n 0.00424615f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_69 VPB N_Y_c_347_n 0.00164882f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_70 VPB N_Y_c_348_n 0.0010843f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.12
cc_71 VPB Y 0.00559339f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_72 N_A1_N_M1008_g N_A2_N_M1004_g 0.0472919f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_73 N_A1_N_M1006_g N_A2_N_c_105_n 0.0409864f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_74 N_A1_N_M1008_g N_A2_N_c_106_n 0.00603804f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_75 N_A1_N_c_74_n N_A2_N_c_106_n 0.00119031f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_76 N_A1_N_M1008_g A2_N 0.00437538f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_77 N_A1_N_M1006_g A2_N 0.00742694f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_78 N_A1_N_c_75_n A2_N 0.059016f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_79 N_A1_N_c_76_n A2_N 0.0114938f $X=0.255 $Y=1.055 $X2=0 $Y2=0
cc_80 N_A1_N_c_74_n N_A2_N_c_108_n 0.0409864f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_81 N_A1_N_c_75_n N_A2_N_c_108_n 4.02983e-19 $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_82 N_A1_N_M1008_g N_A_110_535#_c_161_n 0.00385986f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_83 N_A1_N_M1008_g N_A_110_535#_c_163_n 0.00219638f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_84 N_A1_N_c_75_n N_A_110_535#_c_163_n 0.0094365f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_85 N_A1_N_M1006_g N_A_110_535#_c_155_n 5.74079e-19 $X=0.505 $Y=0.615 $X2=0
+ $Y2=0
cc_86 N_A1_N_M1008_g N_VPWR_c_301_n 0.00930932f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_87 N_A1_N_c_75_n N_VPWR_c_301_n 0.00900898f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_88 N_A1_N_M1008_g N_VPWR_c_302_n 7.04561e-19 $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_89 N_A1_N_M1008_g N_VPWR_c_306_n 0.00486043f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_90 N_A1_N_M1008_g N_VPWR_c_299_n 0.00838234f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_91 N_A1_N_c_75_n N_VPWR_c_299_n 0.00107888f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_92 N_A1_N_M1006_g N_VGND_c_391_n 0.0106012f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_93 N_A1_N_c_74_n N_VGND_c_391_n 0.00437539f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_94 N_A1_N_c_76_n N_VGND_c_391_n 0.015936f $X=0.255 $Y=1.055 $X2=0 $Y2=0
cc_95 N_A1_N_M1006_g N_VGND_c_393_n 0.0045897f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_96 N_A1_N_M1006_g N_VGND_c_395_n 0.0044912f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_97 N_A1_N_c_76_n N_VGND_c_395_n 6.44859e-19 $X=0.255 $Y=1.055 $X2=0 $Y2=0
cc_98 N_A2_N_M1004_g N_A_110_535#_M1007_g 0.0150049f $X=0.905 $Y=2.885 $X2=0
+ $Y2=0
cc_99 N_A2_N_c_105_n N_A_110_535#_c_152_n 3.61617e-19 $X=0.955 $Y=0.935 $X2=0
+ $Y2=0
cc_100 A2_N N_A_110_535#_c_152_n 6.94276e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_101 N_A2_N_c_108_n N_A_110_535#_c_152_n 0.0166053f $X=0.955 $Y=1.1 $X2=0
+ $Y2=0
cc_102 N_A2_N_c_106_n N_A_110_535#_c_154_n 0.0234742f $X=0.955 $Y=1.44 $X2=0
+ $Y2=0
cc_103 A2_N N_A_110_535#_c_154_n 8.05472e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_104 N_A2_N_M1004_g N_A_110_535#_c_161_n 0.00395951f $X=0.905 $Y=2.885 $X2=0
+ $Y2=0
cc_105 N_A2_N_M1004_g N_A_110_535#_c_162_n 0.0112165f $X=0.905 $Y=2.885 $X2=0
+ $Y2=0
cc_106 A2_N N_A_110_535#_c_162_n 0.0156104f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_107 A2_N N_A_110_535#_c_163_n 0.0121653f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_108 N_A2_N_c_105_n N_A_110_535#_c_155_n 0.00393811f $X=0.955 $Y=0.935 $X2=0
+ $Y2=0
cc_109 A2_N N_A_110_535#_c_155_n 0.0074468f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_110 N_A2_N_c_108_n N_A_110_535#_c_155_n 0.00347149f $X=0.955 $Y=1.1 $X2=0
+ $Y2=0
cc_111 N_A2_N_M1004_g N_A_110_535#_c_156_n 0.00153064f $X=0.905 $Y=2.885 $X2=0
+ $Y2=0
cc_112 N_A2_N_c_105_n N_A_110_535#_c_156_n 0.00437259f $X=0.955 $Y=0.935 $X2=0
+ $Y2=0
cc_113 N_A2_N_c_106_n N_A_110_535#_c_156_n 7.54218e-19 $X=0.955 $Y=1.44 $X2=0
+ $Y2=0
cc_114 A2_N N_A_110_535#_c_156_n 0.0794152f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_115 N_A2_N_c_108_n N_A_110_535#_c_156_n 0.00452483f $X=0.955 $Y=1.1 $X2=0
+ $Y2=0
cc_116 N_A2_N_M1004_g N_A_110_535#_c_165_n 0.0426246f $X=0.905 $Y=2.885 $X2=0
+ $Y2=0
cc_117 A2_N N_A_110_535#_c_165_n 0.00188821f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_118 N_A2_N_M1004_g N_VPWR_c_301_n 7.38391e-19 $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_119 N_A2_N_M1004_g N_VPWR_c_302_n 0.00625883f $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_120 N_A2_N_M1004_g N_VPWR_c_306_n 0.00564095f $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_121 N_A2_N_M1004_g N_VPWR_c_299_n 0.00522858f $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_122 N_A2_N_M1004_g N_Y_c_350_n 3.81198e-19 $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_123 N_A2_N_c_105_n N_VGND_c_391_n 0.00143769f $X=0.955 $Y=0.935 $X2=0 $Y2=0
cc_124 N_A2_N_c_105_n N_VGND_c_393_n 0.00527534f $X=0.955 $Y=0.935 $X2=0 $Y2=0
cc_125 N_A2_N_c_105_n N_VGND_c_395_n 0.00534666f $X=0.955 $Y=0.935 $X2=0 $Y2=0
cc_126 A2_N N_VGND_c_395_n 0.0107437f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_127 N_A_110_535#_c_159_n N_B2_M1002_g 0.0335068f $X=1.355 $Y=2.35 $X2=0 $Y2=0
cc_128 N_A_110_535#_c_153_n N_B2_M1009_g 0.0217328f $X=1.975 $Y=0.92 $X2=0 $Y2=0
cc_129 N_A_110_535#_c_151_n N_B2_c_224_n 0.016942f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_110_535#_c_154_n N_B2_c_224_n 0.0335068f $X=1.355 $Y=1.845 $X2=0
+ $Y2=0
cc_131 N_A_110_535#_c_156_n N_B2_c_224_n 9.38875e-19 $X=1.355 $Y=2.01 $X2=0
+ $Y2=0
cc_132 N_A_110_535#_M1007_g N_VPWR_c_302_n 0.00839005f $X=1.445 $Y=2.885 $X2=0
+ $Y2=0
cc_133 N_A_110_535#_c_160_n N_VPWR_c_302_n 0.00215601f $X=1.355 $Y=2.515 $X2=0
+ $Y2=0
cc_134 N_A_110_535#_c_162_n N_VPWR_c_302_n 0.0130771f $X=1.27 $Y=2.43 $X2=0
+ $Y2=0
cc_135 N_A_110_535#_M1007_g N_VPWR_c_304_n 0.00552362f $X=1.445 $Y=2.885 $X2=0
+ $Y2=0
cc_136 N_A_110_535#_c_161_n N_VPWR_c_306_n 0.0078406f $X=0.69 $Y=2.82 $X2=0
+ $Y2=0
cc_137 N_A_110_535#_M1008_d N_VPWR_c_299_n 0.00446753f $X=0.55 $Y=2.675 $X2=0
+ $Y2=0
cc_138 N_A_110_535#_M1007_g N_VPWR_c_299_n 0.00819233f $X=1.445 $Y=2.885 $X2=0
+ $Y2=0
cc_139 N_A_110_535#_c_161_n N_VPWR_c_299_n 0.00694366f $X=0.69 $Y=2.82 $X2=0
+ $Y2=0
cc_140 N_A_110_535#_c_162_n N_VPWR_c_299_n 0.0114592f $X=1.27 $Y=2.43 $X2=0
+ $Y2=0
cc_141 N_A_110_535#_c_151_n N_Y_c_345_n 0.0156284f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_110_535#_c_153_n N_Y_c_345_n 0.00255249f $X=1.975 $Y=0.92 $X2=0 $Y2=0
cc_143 N_A_110_535#_c_154_n N_Y_c_345_n 0.0119611f $X=1.355 $Y=1.845 $X2=0 $Y2=0
cc_144 N_A_110_535#_c_155_n N_Y_c_345_n 0.0111454f $X=1.27 $Y=0.555 $X2=0 $Y2=0
cc_145 N_A_110_535#_c_156_n N_Y_c_345_n 0.101378f $X=1.355 $Y=2.01 $X2=0 $Y2=0
cc_146 N_A_110_535#_c_160_n N_Y_c_347_n 0.00434772f $X=1.355 $Y=2.515 $X2=0
+ $Y2=0
cc_147 N_A_110_535#_c_162_n N_Y_c_347_n 0.00164031f $X=1.27 $Y=2.43 $X2=0 $Y2=0
cc_148 N_A_110_535#_M1007_g N_Y_c_350_n 0.00487837f $X=1.445 $Y=2.885 $X2=0
+ $Y2=0
cc_149 N_A_110_535#_c_159_n N_Y_c_348_n 0.00138233f $X=1.355 $Y=2.35 $X2=0 $Y2=0
cc_150 N_A_110_535#_c_162_n N_Y_c_348_n 0.0106676f $X=1.27 $Y=2.43 $X2=0 $Y2=0
cc_151 N_A_110_535#_c_156_n N_Y_c_348_n 0.00164426f $X=1.355 $Y=2.01 $X2=0 $Y2=0
cc_152 N_A_110_535#_c_155_n N_VGND_c_391_n 0.00709176f $X=1.27 $Y=0.555 $X2=0
+ $Y2=0
cc_153 N_A_110_535#_c_153_n N_VGND_c_393_n 0.00563421f $X=1.975 $Y=0.92 $X2=0
+ $Y2=0
cc_154 N_A_110_535#_c_155_n N_VGND_c_393_n 0.0147613f $X=1.27 $Y=0.555 $X2=0
+ $Y2=0
cc_155 N_A_110_535#_c_153_n N_VGND_c_395_n 0.00539454f $X=1.975 $Y=0.92 $X2=0
+ $Y2=0
cc_156 N_A_110_535#_c_155_n N_VGND_c_395_n 0.0176133f $X=1.27 $Y=0.555 $X2=0
+ $Y2=0
cc_157 N_A_110_535#_c_153_n N_A_410_78#_c_426_n 4.03889e-19 $X=1.975 $Y=0.92
+ $X2=0 $Y2=0
cc_158 N_A_110_535#_c_153_n N_A_410_78#_c_428_n 0.00180793f $X=1.975 $Y=0.92
+ $X2=0 $Y2=0
cc_159 N_B2_M1002_g N_B1_c_268_n 0.0635692f $X=1.875 $Y=2.885 $X2=0 $Y2=0
cc_160 B2 N_B1_c_268_n 7.45138e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_161 N_B2_c_224_n N_B1_c_268_n 0.0207395f $X=2.405 $Y=1.645 $X2=0 $Y2=0
cc_162 N_B2_M1009_g N_B1_M1001_g 0.0317519f $X=2.405 $Y=0.6 $X2=0 $Y2=0
cc_163 B2 N_B1_M1001_g 0.00177582f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_164 B2 N_B1_c_269_n 0.00247415f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_165 N_B2_M1009_g B1 0.00319031f $X=2.405 $Y=0.6 $X2=0 $Y2=0
cc_166 B2 B1 0.0240914f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_167 N_B2_c_224_n N_B1_c_265_n 0.0317519f $X=2.405 $Y=1.645 $X2=0 $Y2=0
cc_168 N_B2_M1002_g N_VPWR_c_303_n 0.0022041f $X=1.875 $Y=2.885 $X2=0 $Y2=0
cc_169 N_B2_M1002_g N_VPWR_c_304_n 0.00552362f $X=1.875 $Y=2.885 $X2=0 $Y2=0
cc_170 N_B2_M1002_g N_VPWR_c_299_n 0.00621827f $X=1.875 $Y=2.885 $X2=0 $Y2=0
cc_171 N_B2_M1002_g N_Y_c_345_n 0.0108775f $X=1.875 $Y=2.885 $X2=0 $Y2=0
cc_172 N_B2_M1009_g N_Y_c_345_n 0.00401946f $X=2.405 $Y=0.6 $X2=0 $Y2=0
cc_173 B2 N_Y_c_345_n 0.0542345f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_174 N_B2_c_224_n N_Y_c_345_n 0.0199202f $X=2.405 $Y=1.645 $X2=0 $Y2=0
cc_175 N_B2_M1002_g N_Y_c_347_n 0.00510983f $X=1.875 $Y=2.885 $X2=0 $Y2=0
cc_176 N_B2_M1002_g N_Y_c_350_n 0.00393485f $X=1.875 $Y=2.885 $X2=0 $Y2=0
cc_177 N_B2_M1002_g N_Y_c_348_n 0.00338167f $X=1.875 $Y=2.885 $X2=0 $Y2=0
cc_178 N_B2_M1002_g Y 0.00856998f $X=1.875 $Y=2.885 $X2=0 $Y2=0
cc_179 B2 Y 0.0123255f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_180 N_B2_c_224_n Y 0.00480458f $X=2.405 $Y=1.645 $X2=0 $Y2=0
cc_181 N_B2_M1009_g N_VGND_c_392_n 0.00329204f $X=2.405 $Y=0.6 $X2=0 $Y2=0
cc_182 N_B2_M1009_g N_VGND_c_393_n 0.00563421f $X=2.405 $Y=0.6 $X2=0 $Y2=0
cc_183 N_B2_M1009_g N_VGND_c_395_n 0.00539454f $X=2.405 $Y=0.6 $X2=0 $Y2=0
cc_184 N_B2_M1009_g N_A_410_78#_c_426_n 6.71115e-19 $X=2.405 $Y=0.6 $X2=0 $Y2=0
cc_185 N_B2_M1009_g N_A_410_78#_c_427_n 0.0160784f $X=2.405 $Y=0.6 $X2=0 $Y2=0
cc_186 N_B2_c_224_n N_A_410_78#_c_427_n 0.00126371f $X=2.405 $Y=1.645 $X2=0
+ $Y2=0
cc_187 B2 N_A_410_78#_c_428_n 0.0140002f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_188 N_B2_c_224_n N_A_410_78#_c_428_n 0.00303127f $X=2.405 $Y=1.645 $X2=0
+ $Y2=0
cc_189 N_B1_M1005_g N_VPWR_c_303_n 0.0112171f $X=2.235 $Y=2.885 $X2=0 $Y2=0
cc_190 N_B1_c_267_n N_VPWR_c_303_n 0.00783066f $X=2.76 $Y=2.295 $X2=0 $Y2=0
cc_191 N_B1_M1005_g N_VPWR_c_304_n 0.00486043f $X=2.235 $Y=2.885 $X2=0 $Y2=0
cc_192 N_B1_M1005_g N_VPWR_c_299_n 0.00566698f $X=2.235 $Y=2.885 $X2=0 $Y2=0
cc_193 B1 N_VPWR_c_299_n 0.0143131f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_194 N_B1_c_268_n N_Y_c_345_n 6.33188e-19 $X=2.31 $Y=2.295 $X2=0 $Y2=0
cc_195 N_B1_M1005_g N_Y_c_347_n 0.00113725f $X=2.235 $Y=2.885 $X2=0 $Y2=0
cc_196 N_B1_M1005_g N_Y_c_350_n 8.63638e-19 $X=2.235 $Y=2.885 $X2=0 $Y2=0
cc_197 N_B1_M1005_g Y 0.00606459f $X=2.235 $Y=2.885 $X2=0 $Y2=0
cc_198 N_B1_c_268_n Y 0.00291227f $X=2.31 $Y=2.295 $X2=0 $Y2=0
cc_199 B1 Y 0.00520662f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_200 N_B1_M1001_g N_VGND_c_392_n 0.00329204f $X=2.835 $Y=0.6 $X2=0 $Y2=0
cc_201 N_B1_M1001_g N_VGND_c_394_n 0.00563421f $X=2.835 $Y=0.6 $X2=0 $Y2=0
cc_202 N_B1_M1001_g N_VGND_c_395_n 0.00539454f $X=2.835 $Y=0.6 $X2=0 $Y2=0
cc_203 N_B1_M1001_g N_A_410_78#_c_427_n 0.0156361f $X=2.835 $Y=0.6 $X2=0 $Y2=0
cc_204 B1 N_A_410_78#_c_427_n 0.0263676f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_205 N_B1_c_265_n N_A_410_78#_c_427_n 6.04532e-19 $X=2.925 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_B1_M1001_g N_A_410_78#_c_429_n 0.00143084f $X=2.835 $Y=0.6 $X2=0 $Y2=0
cc_207 N_VPWR_c_299_n N_Y_M1007_d 0.00246398f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_208 N_VPWR_c_302_n N_Y_c_350_n 0.00565391f $X=1.14 $Y=2.95 $X2=0 $Y2=0
cc_209 N_VPWR_c_303_n N_Y_c_350_n 0.0026493f $X=2.45 $Y=2.95 $X2=0 $Y2=0
cc_210 N_VPWR_c_304_n N_Y_c_350_n 0.00910408f $X=2.285 $Y=3.33 $X2=0 $Y2=0
cc_211 N_VPWR_c_299_n N_Y_c_350_n 0.0110346f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_299_n N_Y_c_348_n 0.00125261f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_299_n Y 0.0119011f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_c_299_n A_390_535# 0.00308167f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_215 N_Y_c_345_n N_VGND_c_393_n 0.00527667f $X=1.76 $Y=0.665 $X2=0 $Y2=0
cc_216 N_Y_c_345_n N_VGND_c_395_n 0.00695878f $X=1.76 $Y=0.665 $X2=0 $Y2=0
cc_217 N_Y_c_345_n N_A_410_78#_c_426_n 0.00314476f $X=1.76 $Y=0.665 $X2=0 $Y2=0
cc_218 N_Y_c_345_n N_A_410_78#_c_428_n 0.0117033f $X=1.76 $Y=0.665 $X2=0 $Y2=0
cc_219 N_VGND_c_393_n N_A_410_78#_c_426_n 0.00467386f $X=2.515 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_395_n N_A_410_78#_c_426_n 0.00677835f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_c_392_n N_A_410_78#_c_427_n 0.0142847f $X=2.62 $Y=0.515 $X2=0
+ $Y2=0
cc_222 N_VGND_c_395_n N_A_410_78#_c_427_n 0.0146356f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_394_n N_A_410_78#_c_429_n 0.00519224f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_224 N_VGND_c_395_n N_A_410_78#_c_429_n 0.00688714f $X=3.12 $Y=0 $X2=0 $Y2=0
