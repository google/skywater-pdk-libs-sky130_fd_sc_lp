# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.765000 1.450000 7.095000 2.130000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 2.320000 3.240000 2.490000 ;
        RECT 2.435000 0.655000 3.240000 0.835000 ;
        RECT 2.435000 0.835000 2.605000 2.260000 ;
        RECT 2.435000 2.260000 3.240000 2.320000 ;
        RECT 2.910000 0.255000 3.240000 0.655000 ;
        RECT 2.960000 2.490000 3.240000 3.075000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.594300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.255000 0.830000 3.075000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.345000 3.825000 1.750000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 8.305000 0.780000 8.675000 2.130000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.120000 0.085000 ;
        RECT 0.095000  0.085000 0.385000 1.095000 ;
        RECT 1.000000  0.085000 1.285000 1.095000 ;
        RECT 2.400000  0.085000 2.730000 0.465000 ;
        RECT 3.410000  0.085000 3.740000 0.835000 ;
        RECT 4.880000  0.085000 5.210000 0.970000 ;
        RECT 6.570000  0.085000 6.900000 0.930000 ;
        RECT 8.150000  0.085000 8.415000 0.610000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.120000 3.415000 ;
        RECT 0.095000 1.815000 0.385000 3.245000 ;
        RECT 1.000000 1.815000 1.290000 3.245000 ;
        RECT 2.460000 2.660000 2.790000 3.245000 ;
        RECT 3.415000 2.260000 3.745000 3.245000 ;
        RECT 4.355000 2.055000 4.685000 3.245000 ;
        RECT 6.355000 2.695000 6.695000 3.245000 ;
        RECT 8.190000 2.640000 8.520000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.000000 1.300000 2.205000 1.630000 ;
      RECT 1.875000 0.715000 2.205000 1.300000 ;
      RECT 1.920000 1.630000 2.205000 2.150000 ;
      RECT 2.775000 1.205000 3.335000 1.535000 ;
      RECT 3.165000 1.005000 4.570000 1.015000 ;
      RECT 3.165000 1.015000 4.080000 1.175000 ;
      RECT 3.165000 1.175000 3.335000 1.205000 ;
      RECT 3.165000 1.535000 3.335000 1.920000 ;
      RECT 3.165000 1.920000 4.185000 2.090000 ;
      RECT 3.910000 0.835000 4.570000 1.005000 ;
      RECT 3.925000 2.090000 4.185000 3.075000 ;
      RECT 3.995000 1.715000 5.135000 1.885000 ;
      RECT 3.995000 1.885000 4.185000 1.920000 ;
      RECT 4.240000 0.255000 4.570000 0.835000 ;
      RECT 4.250000 1.185000 5.795000 1.355000 ;
      RECT 4.250000 1.355000 4.545000 1.535000 ;
      RECT 4.805000 1.525000 5.135000 1.715000 ;
      RECT 5.115000 2.055000 5.445000 2.785000 ;
      RECT 5.115000 2.785000 6.165000 2.955000 ;
      RECT 5.625000 0.640000 6.000000 0.955000 ;
      RECT 5.625000 0.955000 5.795000 1.185000 ;
      RECT 5.625000 1.355000 5.795000 2.275000 ;
      RECT 5.625000 2.275000 5.825000 2.615000 ;
      RECT 5.965000 1.125000 6.165000 1.455000 ;
      RECT 5.995000 1.455000 6.165000 2.355000 ;
      RECT 5.995000 2.355000 7.035000 2.525000 ;
      RECT 5.995000 2.525000 6.165000 2.785000 ;
      RECT 6.335000 1.100000 7.435000 1.270000 ;
      RECT 6.335000 1.270000 6.595000 2.025000 ;
      RECT 6.865000 2.525000 7.035000 2.810000 ;
      RECT 6.865000 2.810000 8.020000 2.980000 ;
      RECT 7.070000 0.640000 7.330000 1.100000 ;
      RECT 7.205000 2.300000 7.435000 2.640000 ;
      RECT 7.265000 1.270000 7.435000 2.300000 ;
      RECT 7.615000 0.280000 7.980000 0.610000 ;
      RECT 7.615000 0.610000 7.785000 2.640000 ;
      RECT 7.615000 2.640000 8.020000 2.810000 ;
      RECT 7.955000 1.585000 8.135000 2.300000 ;
      RECT 7.955000 2.300000 9.025000 2.470000 ;
      RECT 8.585000 0.280000 9.025000 0.610000 ;
      RECT 8.690000 2.470000 9.025000 3.065000 ;
      RECT 8.845000 0.610000 9.025000 2.300000 ;
  END
END sky130_fd_sc_lp__dlrbp_2
