* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4bb_lp A B C_N D_N VGND VNB VPB VPWR Y
X0 a_782_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_302_47# a_27_409# Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_352_409# B a_788_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VGND D_N a_980_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y a_430_21# a_460_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_624_47# B Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Y A a_782_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_788_409# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 Y a_430_21# a_245_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_27_409# C_N a_144_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_27_409# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_144_47# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_27_409# a_302_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND B a_624_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_980_47# D_N a_430_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_245_409# a_27_409# a_352_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 VPWR D_N a_430_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_460_47# a_430_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
