* File: sky130_fd_sc_lp__and2_1.pex.spice
* Created: Fri Aug 28 10:04:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2_1%A 3 7 9 10 11 12
r27 12 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.7
+ $Y=1.585 $X2=0.7 $Y2=1.585
r28 11 12 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=0.24 $Y=1.62 $X2=0.7
+ $Y2=1.62
r29 9 16 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.725 $Y=1.585
+ $X2=0.7 $Y2=1.585
r30 9 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.725 $Y=1.585
+ $X2=0.8 $Y2=1.585
r31 5 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.8 $Y=1.75 $X2=0.8
+ $Y2=1.585
r32 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.8 $Y=1.75 $X2=0.8
+ $Y2=2.12
r33 1 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.8 $Y=1.42 $X2=0.8
+ $Y2=1.585
r34 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.8 $Y=1.42 $X2=0.8
+ $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_1%B 3 7 9 12
c34 9 0 1.47301e-19 $X=1.2 $Y=1.665
c35 3 0 1.77145e-19 $X=1.16 $Y=0.865
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.585
+ $X2=1.25 $Y2=1.75
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.585
+ $X2=1.25 $Y2=1.42
r38 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.585 $X2=1.25 $Y2=1.585
r39 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.34 $Y=2.12 $X2=1.34
+ $Y2=1.75
r40 3 14 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.16 $Y=0.865
+ $X2=1.16 $Y2=1.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_1%A_92_131# 1 2 7 9 12 16 18 19 20 25 27 35
c51 35 0 1.47301e-19 $X=1.925 $Y=1.35
r52 27 30 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.085 $Y=2.005
+ $X2=1.085 $Y2=2.12
r53 26 35 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.79 $Y=1.35
+ $X2=1.925 $Y2=1.35
r54 26 32 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.79 $Y=1.35 $X2=1.7
+ $Y2=1.35
r55 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.35 $X2=1.79 $Y2=1.35
r56 23 25 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=1.75 $Y=1.92
+ $X2=1.75 $Y2=1.35
r57 22 25 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=1.75 $Y=1.32 $X2=1.75
+ $Y2=1.35
r58 21 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=2.005
+ $X2=1.085 $Y2=2.005
r59 20 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.625 $Y=2.005
+ $X2=1.75 $Y2=1.92
r60 20 21 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.625 $Y=2.005
+ $X2=1.25 $Y2=2.005
r61 18 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.625 $Y=1.235
+ $X2=1.75 $Y2=1.32
r62 18 19 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.625 $Y=1.235
+ $X2=0.75 $Y2=1.235
r63 14 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.585 $Y=1.15
+ $X2=0.75 $Y2=1.235
r64 14 16 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.585 $Y=1.15
+ $X2=0.585 $Y2=0.865
r65 10 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.515
+ $X2=1.925 $Y2=1.35
r66 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.925 $Y=1.515
+ $X2=1.925 $Y2=2.465
r67 7 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.185 $X2=1.7
+ $Y2=1.35
r68 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.7 $Y=1.185 $X2=1.7
+ $Y2=0.655
r69 2 30 600 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_PDIFF $count=1 $X=0.875
+ $Y=1.91 $X2=1.085 $Y2=2.12
r70 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.46
+ $Y=0.655 $X2=0.585 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_1%VPWR 1 2 9 13 16 17 18 24 30 31 34
r25 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.71 $Y2=3.33
r29 28 30 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.71 $Y2=3.33
r31 24 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r32 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 18 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 18 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 16 21 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.42 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.42 $Y=3.33
+ $X2=0.585 $Y2=3.33
r38 15 26 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.75 $Y=3.33 $X2=1.2
+ $Y2=3.33
r39 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=3.33
+ $X2=0.585 $Y2=3.33
r40 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=3.33
r41 11 13 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=2.365
r42 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=3.245
+ $X2=0.585 $Y2=3.33
r43 7 9 39.2878 $w=3.28e-07 $l=1.125e-06 $layer=LI1_cond $X=0.585 $Y=3.245
+ $X2=0.585 $Y2=2.12
r44 2 13 300 $w=1.7e-07 $l=5.84166e-07 $layer=licon1_PDIFF $count=2 $X=1.415
+ $Y=1.91 $X2=1.71 $Y2=2.365
r45 1 9 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.46
+ $Y=1.91 $X2=0.585 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_1%X 1 2 7 8 9 10 11 12 13 39 45
c16 39 0 1.77145e-19 $X=1.915 $Y=0.38
r17 45 46 4.43927 $w=5.63e-07 $l=5.5e-08 $layer=LI1_cond $X=2.032 $Y=0.925
+ $X2=2.032 $Y2=0.98
r18 13 36 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.18 $Y=2.775
+ $X2=2.18 $Y2=2.91
r19 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.18 $Y=2.405
+ $X2=2.18 $Y2=2.775
r20 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.18 $Y=1.98
+ $X2=2.18 $Y2=2.405
r21 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.18 $Y=1.665
+ $X2=2.18 $Y2=1.98
r22 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.18 $Y=1.295
+ $X2=2.18 $Y2=1.665
r23 8 45 0.317543 $w=5.63e-07 $l=1.5e-08 $layer=LI1_cond $X=2.032 $Y=0.91
+ $X2=2.032 $Y2=0.925
r24 8 9 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=2.18 $Y=0.995 $X2=2.18
+ $Y2=1.295
r25 8 46 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.18 $Y=0.995
+ $X2=2.18 $Y2=0.98
r26 7 8 7.51518 $w=5.63e-07 $l=3.55e-07 $layer=LI1_cond $X=2.032 $Y=0.555
+ $X2=2.032 $Y2=0.91
r27 7 39 3.70467 $w=5.63e-07 $l=1.75e-07 $layer=LI1_cond $X=2.032 $Y=0.555
+ $X2=2.032 $Y2=0.38
r28 2 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.835 $X2=2.14 $Y2=2.91
r29 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.835 $X2=2.14 $Y2=1.98
r30 1 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.775
+ $Y=0.235 $X2=1.915 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_1%VGND 1 6 11 12 13 23 24
r21 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r22 16 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r23 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r24 13 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r25 13 17 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r26 13 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r27 11 20 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.21 $Y=0 $X2=1.2
+ $Y2=0
r28 11 12 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.21 $Y=0 $X2=1.395
+ $Y2=0
r29 10 23 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=2.16
+ $Y2=0
r30 10 12 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=1.395
+ $Y2=0
r31 6 8 16.0408 $w=3.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.395 $Y=0.38
+ $X2=1.395 $Y2=0.895
r32 4 12 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=0.085
+ $X2=1.395 $Y2=0
r33 4 6 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.395 $Y=0.085
+ $X2=1.395 $Y2=0.38
r34 1 8 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=1.235
+ $Y=0.655 $X2=1.375 $Y2=0.895
r35 1 6 182 $w=1.7e-07 $l=3.79967e-07 $layer=licon1_NDIFF $count=1 $X=1.235
+ $Y=0.655 $X2=1.485 $Y2=0.38
.ends

