* File: sky130_fd_sc_lp__a21boi_1.spice
* Created: Wed Sep  2 09:19:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21boi_1.pex.spice"
.subckt sky130_fd_sc_lp__a21boi_1  VNB VPB B1_N A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_B1_N_M1002_g N_A_27_508#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=27.132 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A_27_508#_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1449 AS=0.1792 PD=1.185 PS=1.62 NRD=4.284 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1005 A_380_47# N_A1_M1005_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.84 AD=0.1764
+ AS=0.1449 PD=1.26 PS=1.185 NRD=22.14 NRS=4.992 M=1 R=5.6 SA=75000.9 SB=75000.8
+ A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g A_380_47# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1764 PD=2.21 PS=1.26 NRD=0 NRS=22.14 M=1 R=5.6 SA=75001.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_B1_N_M1001_g N_A_27_508#_M1001_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_302_367#_M1000_d N_A_27_508#_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_302_367#_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2394 AS=0.1764 PD=1.64 PS=1.54 NRD=8.5892 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1003 N_A_302_367#_M1003_d N_A2_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2394 PD=3.05 PS=1.64 NRD=0 NRS=7.0329 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__a21boi_1.pxi.spice"
*
.ends
*
*
