* File: sky130_fd_sc_lp__a22oi_4.pex.spice
* Created: Fri Aug 28 09:55:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22OI_4%B2 3 5 8 10 12 15 17 19 22 24 26 29 31 32 33
+ 34 35 42 62
c87 24 0 5.31181e-20 $X=1.945 $Y=1.275
c88 17 0 9.06625e-20 $X=1.515 $Y=1.275
c89 10 0 9.06625e-20 $X=1.085 $Y=1.275
r90 60 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.985 $Y=1.44
+ $X2=2.075 $Y2=1.44
r91 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.985
+ $Y=1.44 $X2=1.985 $Y2=1.44
r92 58 60 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.945 $Y=1.44
+ $X2=1.985 $Y2=1.44
r93 56 58 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=1.645 $Y=1.44
+ $X2=1.945 $Y2=1.44
r94 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.645
+ $Y=1.44 $X2=1.645 $Y2=1.44
r95 54 56 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.515 $Y=1.44
+ $X2=1.645 $Y2=1.44
r96 53 57 12.4391 $w=3.13e-07 $l=3.4e-07 $layer=LI1_cond $X=1.305 $Y=1.367
+ $X2=1.645 $Y2=1.367
r97 52 54 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.305 $Y=1.44
+ $X2=1.515 $Y2=1.44
r98 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.305
+ $Y=1.44 $X2=1.305 $Y2=1.44
r99 50 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.215 $Y=1.44
+ $X2=1.305 $Y2=1.44
r100 49 50 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.085 $Y=1.44
+ $X2=1.215 $Y2=1.44
r101 47 49 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=0.965 $Y=1.44
+ $X2=1.085 $Y2=1.44
r102 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.44 $X2=0.965 $Y2=1.44
r103 45 47 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.785 $Y=1.44
+ $X2=0.965 $Y2=1.44
r104 44 45 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=0.655 $Y=1.44
+ $X2=0.785 $Y2=1.44
r105 42 44 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.625 $Y=1.44
+ $X2=0.655 $Y2=1.44
r106 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.625
+ $Y=1.44 $X2=0.625 $Y2=1.44
r107 35 61 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=2.16 $Y=1.367
+ $X2=1.985 $Y2=1.367
r108 34 61 11.1586 $w=3.13e-07 $l=3.05e-07 $layer=LI1_cond $X=1.68 $Y=1.367
+ $X2=1.985 $Y2=1.367
r109 34 57 1.28049 $w=3.13e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=1.367
+ $X2=1.645 $Y2=1.367
r110 33 53 3.84148 $w=3.13e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.367
+ $X2=1.305 $Y2=1.367
r111 33 48 8.59759 $w=3.13e-07 $l=2.35e-07 $layer=LI1_cond $X=1.2 $Y=1.367
+ $X2=0.965 $Y2=1.367
r112 32 48 8.96345 $w=3.13e-07 $l=2.45e-07 $layer=LI1_cond $X=0.72 $Y=1.367
+ $X2=0.965 $Y2=1.367
r113 32 43 3.47562 $w=3.13e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=1.367
+ $X2=0.625 $Y2=1.367
r114 31 43 14.0854 $w=3.13e-07 $l=3.85e-07 $layer=LI1_cond $X=0.24 $Y=1.367
+ $X2=0.625 $Y2=1.367
r115 27 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.605
+ $X2=2.075 $Y2=1.44
r116 27 29 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.075 $Y=1.605
+ $X2=2.075 $Y2=2.465
r117 24 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.945 $Y=1.275
+ $X2=1.945 $Y2=1.44
r118 24 26 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.945 $Y=1.275
+ $X2=1.945 $Y2=0.745
r119 20 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.645 $Y=1.605
+ $X2=1.645 $Y2=1.44
r120 20 22 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.645 $Y=1.605
+ $X2=1.645 $Y2=2.465
r121 17 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.275
+ $X2=1.515 $Y2=1.44
r122 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.515 $Y=1.275
+ $X2=1.515 $Y2=0.745
r123 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=1.605
+ $X2=1.215 $Y2=1.44
r124 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.215 $Y=1.605
+ $X2=1.215 $Y2=2.465
r125 10 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.275
+ $X2=1.085 $Y2=1.44
r126 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.085 $Y=1.275
+ $X2=1.085 $Y2=0.745
r127 6 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.785 $Y=1.605
+ $X2=0.785 $Y2=1.44
r128 6 8 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.785 $Y=1.605
+ $X2=0.785 $Y2=2.465
r129 3 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.275
+ $X2=0.655 $Y2=1.44
r130 3 5 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.655 $Y=1.275
+ $X2=0.655 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 51 55 69
r95 55 69 1.72325 $w=3.15e-07 $l=2.2e-08 $layer=LI1_cond $X=3.142 $Y=1.367
+ $X2=3.12 $Y2=1.367
r96 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.96
+ $Y=1.44 $X2=3.96 $Y2=1.44
r97 51 53 12.7236 $w=3.22e-07 $l=8.5e-08 $layer=POLY_cond $X=3.875 $Y=1.44
+ $X2=3.96 $Y2=1.44
r98 50 51 22.4534 $w=3.22e-07 $l=1.5e-07 $layer=POLY_cond $X=3.725 $Y=1.44
+ $X2=3.875 $Y2=1.44
r99 49 54 12.4391 $w=3.13e-07 $l=3.4e-07 $layer=LI1_cond $X=3.62 $Y=1.367
+ $X2=3.96 $Y2=1.367
r100 48 50 15.7174 $w=3.22e-07 $l=1.05e-07 $layer=POLY_cond $X=3.62 $Y=1.44
+ $X2=3.725 $Y2=1.44
r101 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.62
+ $Y=1.44 $X2=3.62 $Y2=1.44
r102 46 48 26.1957 $w=3.22e-07 $l=1.75e-07 $layer=POLY_cond $X=3.445 $Y=1.44
+ $X2=3.62 $Y2=1.44
r103 45 46 22.4534 $w=3.22e-07 $l=1.5e-07 $layer=POLY_cond $X=3.295 $Y=1.44
+ $X2=3.445 $Y2=1.44
r104 43 45 2.24534 $w=3.22e-07 $l=1.5e-08 $layer=POLY_cond $X=3.28 $Y=1.44
+ $X2=3.295 $Y2=1.44
r105 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.28
+ $Y=1.44 $X2=3.28 $Y2=1.44
r106 41 43 51.6429 $w=3.22e-07 $l=3.45e-07 $layer=POLY_cond $X=2.935 $Y=1.44
+ $X2=3.28 $Y2=1.44
r107 40 41 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=2.865 $Y=1.44
+ $X2=2.935 $Y2=1.44
r108 39 40 53.8882 $w=3.22e-07 $l=3.6e-07 $layer=POLY_cond $X=2.505 $Y=1.44
+ $X2=2.865 $Y2=1.44
r109 38 39 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=2.435 $Y=1.44
+ $X2=2.505 $Y2=1.44
r110 31 32 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.367
+ $X2=4.56 $Y2=1.367
r111 31 54 4.39026 $w=3.13e-07 $l=1.2e-07 $layer=LI1_cond $X=4.08 $Y=1.367
+ $X2=3.96 $Y2=1.367
r112 30 49 0.73171 $w=3.13e-07 $l=2e-08 $layer=LI1_cond $X=3.6 $Y=1.367 $X2=3.62
+ $Y2=1.367
r113 30 44 11.7074 $w=3.13e-07 $l=3.2e-07 $layer=LI1_cond $X=3.6 $Y=1.367
+ $X2=3.28 $Y2=1.367
r114 29 69 1.68276 $w=2.32e-07 $l=3.2e-08 $layer=LI1_cond $X=3.088 $Y=1.367
+ $X2=3.12 $Y2=1.367
r115 29 44 3.91465 $w=3.13e-07 $l=1.07e-07 $layer=LI1_cond $X=3.173 $Y=1.367
+ $X2=3.28 $Y2=1.367
r116 29 55 1.13415 $w=3.13e-07 $l=3.1e-08 $layer=LI1_cond $X=3.173 $Y=1.367
+ $X2=3.142 $Y2=1.367
r117 25 51 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.875 $Y=1.605
+ $X2=3.875 $Y2=1.44
r118 25 27 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.875 $Y=1.605
+ $X2=3.875 $Y2=2.465
r119 22 50 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.725 $Y=1.275
+ $X2=3.725 $Y2=1.44
r120 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.725 $Y=1.275
+ $X2=3.725 $Y2=0.745
r121 18 46 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.445 $Y=1.605
+ $X2=3.445 $Y2=1.44
r122 18 20 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.445 $Y=1.605
+ $X2=3.445 $Y2=2.465
r123 15 45 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.275
+ $X2=3.295 $Y2=1.44
r124 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.295 $Y=1.275
+ $X2=3.295 $Y2=0.745
r125 11 41 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.935 $Y=1.605
+ $X2=2.935 $Y2=1.44
r126 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.935 $Y=1.605
+ $X2=2.935 $Y2=2.465
r127 8 40 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.275
+ $X2=2.865 $Y2=1.44
r128 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.865 $Y=1.275
+ $X2=2.865 $Y2=0.745
r129 4 39 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=1.605
+ $X2=2.505 $Y2=1.44
r130 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.505 $Y=1.605
+ $X2=2.505 $Y2=2.465
r131 1 38 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.275
+ $X2=2.435 $Y2=1.44
r132 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.435 $Y=1.275
+ $X2=2.435 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_4%A1 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 49
r85 47 49 3.07006 $w=3.14e-07 $l=2e-08 $layer=POLY_cond $X=5.725 $Y=1.35
+ $X2=5.745 $Y2=1.35
r86 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.725
+ $Y=1.35 $X2=5.725 $Y2=1.35
r87 45 47 29.1656 $w=3.14e-07 $l=1.9e-07 $layer=POLY_cond $X=5.535 $Y=1.35
+ $X2=5.725 $Y2=1.35
r88 44 45 40.6783 $w=3.14e-07 $l=2.65e-07 $layer=POLY_cond $X=5.27 $Y=1.35
+ $X2=5.535 $Y2=1.35
r89 43 44 25.328 $w=3.14e-07 $l=1.65e-07 $layer=POLY_cond $X=5.105 $Y=1.35
+ $X2=5.27 $Y2=1.35
r90 41 43 9.21019 $w=3.14e-07 $l=6e-08 $layer=POLY_cond $X=5.045 $Y=1.35
+ $X2=5.105 $Y2=1.35
r91 39 41 31.4682 $w=3.14e-07 $l=2.05e-07 $layer=POLY_cond $X=4.84 $Y=1.35
+ $X2=5.045 $Y2=1.35
r92 38 39 25.328 $w=3.14e-07 $l=1.65e-07 $layer=POLY_cond $X=4.675 $Y=1.35
+ $X2=4.84 $Y2=1.35
r93 37 38 40.6783 $w=3.14e-07 $l=2.65e-07 $layer=POLY_cond $X=4.41 $Y=1.35
+ $X2=4.675 $Y2=1.35
r94 31 32 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6 $Y=1.322 $X2=6.48
+ $Y2=1.322
r95 31 48 14.0854 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=6 $Y=1.322
+ $X2=5.725 $Y2=1.322
r96 30 48 10.5 $w=2.23e-07 $l=2.05e-07 $layer=LI1_cond $X=5.52 $Y=1.322
+ $X2=5.725 $Y2=1.322
r97 29 30 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.322
+ $X2=5.52 $Y2=1.322
r98 29 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.045
+ $Y=1.35 $X2=5.045 $Y2=1.35
r99 26 49 33.7707 $w=3.14e-07 $l=2.91033e-07 $layer=POLY_cond $X=5.965 $Y=1.185
+ $X2=5.745 $Y2=1.35
r100 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.965 $Y=1.185
+ $X2=5.965 $Y2=0.655
r101 22 49 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.745 $Y=1.515
+ $X2=5.745 $Y2=1.35
r102 22 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.745 $Y=1.515
+ $X2=5.745 $Y2=2.465
r103 19 45 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.535 $Y=1.185
+ $X2=5.535 $Y2=1.35
r104 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.535 $Y=1.185
+ $X2=5.535 $Y2=0.655
r105 15 44 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.27 $Y=1.515
+ $X2=5.27 $Y2=1.35
r106 15 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.27 $Y=1.515
+ $X2=5.27 $Y2=2.465
r107 12 43 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.105 $Y=1.185
+ $X2=5.105 $Y2=1.35
r108 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.105 $Y=1.185
+ $X2=5.105 $Y2=0.655
r109 8 39 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.84 $Y=1.515
+ $X2=4.84 $Y2=1.35
r110 8 10 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.84 $Y=1.515
+ $X2=4.84 $Y2=2.465
r111 5 38 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.675 $Y=1.185
+ $X2=4.675 $Y2=1.35
r112 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.675 $Y=1.185
+ $X2=4.675 $Y2=0.655
r113 1 37 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=1.515
+ $X2=4.41 $Y2=1.35
r114 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.41 $Y=1.515
+ $X2=4.41 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 46
c72 13 0 1.39855e-19 $X=6.825 $Y=0.655
r73 46 48 12.4298 $w=3.49e-07 $l=9e-08 $layer=POLY_cond $X=7.595 $Y=1.535
+ $X2=7.685 $Y2=1.535
r74 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.595
+ $Y=1.51 $X2=7.595 $Y2=1.51
r75 44 46 17.9542 $w=3.49e-07 $l=1.3e-07 $layer=POLY_cond $X=7.465 $Y=1.535
+ $X2=7.595 $Y2=1.535
r76 43 44 29.0029 $w=3.49e-07 $l=2.1e-07 $layer=POLY_cond $X=7.255 $Y=1.535
+ $X2=7.465 $Y2=1.535
r77 42 43 30.384 $w=3.49e-07 $l=2.2e-07 $layer=POLY_cond $X=7.035 $Y=1.535
+ $X2=7.255 $Y2=1.535
r78 40 42 16.5731 $w=3.49e-07 $l=1.2e-07 $layer=POLY_cond $X=6.915 $Y=1.535
+ $X2=7.035 $Y2=1.535
r79 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.915
+ $Y=1.51 $X2=6.915 $Y2=1.51
r80 38 40 12.4298 $w=3.49e-07 $l=9e-08 $layer=POLY_cond $X=6.825 $Y=1.535
+ $X2=6.915 $Y2=1.535
r81 37 38 30.384 $w=3.49e-07 $l=2.2e-07 $layer=POLY_cond $X=6.605 $Y=1.535
+ $X2=6.825 $Y2=1.535
r82 36 37 29.0029 $w=3.49e-07 $l=2.1e-07 $layer=POLY_cond $X=6.395 $Y=1.535
+ $X2=6.605 $Y2=1.535
r83 31 47 11.1804 $w=3.33e-07 $l=3.25e-07 $layer=LI1_cond $X=7.92 $Y=1.592
+ $X2=7.595 $Y2=1.592
r84 30 47 5.3322 $w=3.33e-07 $l=1.55e-07 $layer=LI1_cond $X=7.44 $Y=1.592
+ $X2=7.595 $Y2=1.592
r85 29 30 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.592
+ $X2=7.44 $Y2=1.592
r86 29 41 1.54806 $w=3.33e-07 $l=4.5e-08 $layer=LI1_cond $X=6.96 $Y=1.592
+ $X2=6.915 $Y2=1.592
r87 25 48 22.56 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.685 $Y=1.345
+ $X2=7.685 $Y2=1.535
r88 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.685 $Y=1.345
+ $X2=7.685 $Y2=0.655
r89 22 44 22.56 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.465 $Y=1.725
+ $X2=7.465 $Y2=1.535
r90 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.465 $Y=1.725
+ $X2=7.465 $Y2=2.465
r91 18 43 22.56 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.255 $Y=1.345
+ $X2=7.255 $Y2=1.535
r92 18 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.255 $Y=1.345
+ $X2=7.255 $Y2=0.655
r93 15 42 22.56 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.035 $Y=1.725
+ $X2=7.035 $Y2=1.535
r94 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.035 $Y=1.725
+ $X2=7.035 $Y2=2.465
r95 11 38 22.56 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.825 $Y=1.345
+ $X2=6.825 $Y2=1.535
r96 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.825 $Y=1.345
+ $X2=6.825 $Y2=0.655
r97 8 37 22.56 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.605 $Y=1.725
+ $X2=6.605 $Y2=1.535
r98 8 10 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.605 $Y=1.725
+ $X2=6.605 $Y2=2.465
r99 4 36 22.56 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.395 $Y=1.345
+ $X2=6.395 $Y2=1.535
r100 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.395 $Y=1.345
+ $X2=6.395 $Y2=0.655
r101 1 36 30.384 $w=3.49e-07 $l=3.00333e-07 $layer=POLY_cond $X=6.175 $Y=1.725
+ $X2=6.395 $Y2=1.535
r102 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.175 $Y=1.725
+ $X2=6.175 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_4%A_89_367# 1 2 3 4 5 6 7 8 9 28 30 32 36 38
+ 42 46 50 54 57 60 61 64 68 70 72 74 78 80 82 84 89 90 91 94 100
r109 97 98 1.86463 $w=2.29e-07 $l=3.5e-08 $layer=LI1_cond $X=5.937 $Y=1.98
+ $X2=5.937 $Y2=2.015
r110 95 97 7.45852 $w=2.29e-07 $l=1.4e-07 $layer=LI1_cond $X=5.937 $Y=1.84
+ $X2=5.937 $Y2=1.98
r111 82 102 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.715 $Y=2.1
+ $X2=7.715 $Y2=2.015
r112 82 84 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=7.715 $Y=2.1
+ $X2=7.715 $Y2=2.91
r113 81 100 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.915 $Y=2.015
+ $X2=6.82 $Y2=2.015
r114 80 102 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.585 $Y=2.015
+ $X2=7.715 $Y2=2.015
r115 80 81 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.585 $Y=2.015
+ $X2=6.915 $Y2=2.015
r116 76 100 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=2.1
+ $X2=6.82 $Y2=2.015
r117 76 78 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=6.82 $Y=2.1
+ $X2=6.82 $Y2=2.91
r118 75 98 2.48377 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=6.055 $Y=2.015
+ $X2=5.937 $Y2=2.015
r119 74 100 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.725 $Y=2.015
+ $X2=6.82 $Y2=2.015
r120 74 75 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.725 $Y=2.015
+ $X2=6.055 $Y2=2.015
r121 70 98 4.41277 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=5.937 $Y=2.1
+ $X2=5.937 $Y2=2.015
r122 70 72 17.6544 $w=2.33e-07 $l=3.6e-07 $layer=LI1_cond $X=5.937 $Y=2.1
+ $X2=5.937 $Y2=2.46
r123 69 94 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.15 $Y=1.84
+ $X2=5.055 $Y2=1.84
r124 68 95 2.48377 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=5.82 $Y=1.84
+ $X2=5.937 $Y2=1.84
r125 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.82 $Y=1.84
+ $X2=5.15 $Y2=1.84
r126 64 66 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=5.055 $Y=1.98
+ $X2=5.055 $Y2=2.91
r127 62 94 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=1.925
+ $X2=5.055 $Y2=1.84
r128 62 64 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=5.055 $Y=1.925
+ $X2=5.055 $Y2=1.98
r129 60 94 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.96 $Y=1.84
+ $X2=5.055 $Y2=1.84
r130 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.96 $Y=1.84
+ $X2=4.29 $Y2=1.84
r131 57 93 2.73961 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.142 $Y=2.905
+ $X2=4.142 $Y2=2.99
r132 57 59 36.1359 $w=2.93e-07 $l=9.25e-07 $layer=LI1_cond $X=4.142 $Y=2.905
+ $X2=4.142 $Y2=1.98
r133 56 61 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=4.142 $Y=1.925
+ $X2=4.29 $Y2=1.84
r134 56 59 2.14862 $w=2.93e-07 $l=5.5e-08 $layer=LI1_cond $X=4.142 $Y=1.925
+ $X2=4.142 $Y2=1.98
r135 55 91 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.325 $Y=2.99
+ $X2=3.19 $Y2=2.99
r136 54 93 4.73791 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=3.995 $Y=2.99
+ $X2=4.142 $Y2=2.99
r137 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.995 $Y=2.99
+ $X2=3.325 $Y2=2.99
r138 50 53 29.4513 $w=2.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.19 $Y=2.21
+ $X2=3.19 $Y2=2.9
r139 48 91 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=2.905
+ $X2=3.19 $Y2=2.99
r140 48 53 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=3.19 $Y=2.905
+ $X2=3.19 $Y2=2.9
r141 47 90 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.385 $Y=2.99
+ $X2=2.29 $Y2=2.99
r142 46 91 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.055 $Y=2.99
+ $X2=3.19 $Y2=2.99
r143 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.055 $Y=2.99
+ $X2=2.385 $Y2=2.99
r144 42 45 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=2.29 $Y=2.21
+ $X2=2.29 $Y2=2.9
r145 40 90 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=2.905
+ $X2=2.29 $Y2=2.99
r146 40 45 0.291866 $w=1.88e-07 $l=5e-09 $layer=LI1_cond $X=2.29 $Y=2.905
+ $X2=2.29 $Y2=2.9
r147 39 89 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.525 $Y=2.99
+ $X2=1.43 $Y2=2.99
r148 38 90 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.195 $Y=2.99
+ $X2=2.29 $Y2=2.99
r149 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.195 $Y=2.99
+ $X2=1.525 $Y2=2.99
r150 34 89 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.43 $Y=2.905
+ $X2=1.43 $Y2=2.99
r151 34 36 40.5694 $w=1.88e-07 $l=6.95e-07 $layer=LI1_cond $X=1.43 $Y=2.905
+ $X2=1.43 $Y2=2.21
r152 33 87 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.665 $Y=2.99
+ $X2=0.535 $Y2=2.99
r153 32 89 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.335 $Y=2.99
+ $X2=1.43 $Y2=2.99
r154 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.335 $Y=2.99
+ $X2=0.665 $Y2=2.99
r155 28 87 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.535 $Y=2.905
+ $X2=0.535 $Y2=2.99
r156 28 30 40.5571 $w=2.58e-07 $l=9.15e-07 $layer=LI1_cond $X=0.535 $Y=2.905
+ $X2=0.535 $Y2=1.99
r157 9 102 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=1.835 $X2=7.68 $Y2=2.095
r158 9 84 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=1.835 $X2=7.68 $Y2=2.91
r159 8 100 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=6.68
+ $Y=1.835 $X2=6.82 $Y2=2.095
r160 8 78 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.68
+ $Y=1.835 $X2=6.82 $Y2=2.91
r161 7 97 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.835 $X2=5.96 $Y2=1.98
r162 7 72 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=5.82
+ $Y=1.835 $X2=5.96 $Y2=2.46
r163 6 66 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.915
+ $Y=1.835 $X2=5.055 $Y2=2.91
r164 6 64 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.915
+ $Y=1.835 $X2=5.055 $Y2=1.98
r165 5 93 400 $w=1.7e-07 $l=1.16614e-06 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.835 $X2=4.14 $Y2=2.91
r166 5 59 400 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.835 $X2=4.14 $Y2=1.98
r167 4 53 400 $w=1.7e-07 $l=1.1561e-06 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.835 $X2=3.2 $Y2=2.9
r168 4 50 400 $w=1.7e-07 $l=4.60299e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.835 $X2=3.2 $Y2=2.21
r169 3 45 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=2.15
+ $Y=1.835 $X2=2.29 $Y2=2.9
r170 3 42 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=2.15
+ $Y=1.835 $X2=2.29 $Y2=2.21
r171 2 89 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.29
+ $Y=1.835 $X2=1.43 $Y2=2.91
r172 2 36 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=1.29
+ $Y=1.835 $X2=1.43 $Y2=2.21
r173 1 87 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.445
+ $Y=1.835 $X2=0.57 $Y2=2.91
r174 1 30 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.445
+ $Y=1.835 $X2=0.57 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_4%Y 1 2 3 4 5 6 7 8 27 29 30 33 35 38 41 43 47
+ 49 50 52 55 57 58 59 60 61 81
c114 38 0 5.31181e-20 $X=2.51 $Y=1.705
r115 85 86 10.1738 $w=3.88e-07 $l=2.18e-07 $layer=LI1_cond $X=2.62 $Y=0.927
+ $X2=2.62 $Y2=1.145
r116 67 85 3.97128 $w=2.25e-07 $l=1.95e-07 $layer=LI1_cond $X=2.815 $Y=0.927
+ $X2=2.62 $Y2=0.927
r117 61 79 16.9025 $w=2.23e-07 $l=3.3e-07 $layer=LI1_cond $X=4.56 $Y=0.927
+ $X2=4.89 $Y2=0.927
r118 60 61 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=0.927
+ $X2=4.56 $Y2=0.927
r119 59 60 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=0.927
+ $X2=4.08 $Y2=0.927
r120 59 71 4.60977 $w=2.23e-07 $l=9e-08 $layer=LI1_cond $X=3.6 $Y=0.927 $X2=3.51
+ $Y2=0.927
r121 58 71 19.9757 $w=2.23e-07 $l=3.9e-07 $layer=LI1_cond $X=3.12 $Y=0.927
+ $X2=3.51 $Y2=0.927
r122 58 67 15.622 $w=2.23e-07 $l=3.05e-07 $layer=LI1_cond $X=3.12 $Y=0.927
+ $X2=2.815 $Y2=0.927
r123 57 85 0.0590996 $w=3.88e-07 $l=2e-09 $layer=LI1_cond $X=2.62 $Y=0.925
+ $X2=2.62 $Y2=0.927
r124 57 81 6.64871 $w=3.88e-07 $l=2.25e-07 $layer=LI1_cond $X=2.62 $Y=0.925
+ $X2=2.62 $Y2=0.7
r125 55 79 38.6709 $w=2.23e-07 $l=7.55e-07 $layer=LI1_cond $X=5.645 $Y=0.927
+ $X2=4.89 $Y2=0.927
r126 54 55 0.0152155 $w=2.25e-07 $l=1e-07 $layer=LI1_cond $X=5.745 $Y=0.927
+ $X2=5.645 $Y2=0.927
r127 52 54 3.71545 $w=1.98e-07 $l=6.7e-08 $layer=LI1_cond $X=5.745 $Y=0.86
+ $X2=5.745 $Y2=0.927
r128 45 47 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.66 $Y=1.875
+ $X2=3.66 $Y2=1.98
r129 44 50 4.30018 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.885 $Y=1.79
+ $X2=2.655 $Y2=1.79
r130 43 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.495 $Y=1.79
+ $X2=3.66 $Y2=1.875
r131 43 44 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.495 $Y=1.79
+ $X2=2.885 $Y2=1.79
r132 39 50 1.96316 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.72 $Y=1.875
+ $X2=2.655 $Y2=1.79
r133 39 41 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.72 $Y=1.875
+ $X2=2.72 $Y2=1.98
r134 38 50 1.96316 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.51 $Y=1.705
+ $X2=2.655 $Y2=1.79
r135 38 86 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.51 $Y=1.705
+ $X2=2.51 $Y2=1.145
r136 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=1.79
+ $X2=1.86 $Y2=1.79
r137 35 50 4.30018 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.425 $Y=1.79
+ $X2=2.655 $Y2=1.79
r138 35 36 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.425 $Y=1.79
+ $X2=2.025 $Y2=1.79
r139 31 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=1.875
+ $X2=1.86 $Y2=1.79
r140 31 33 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.86 $Y=1.875
+ $X2=1.86 $Y2=1.98
r141 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=1.79
+ $X2=1.86 $Y2=1.79
r142 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.695 $Y=1.79
+ $X2=1.165 $Y2=1.79
r143 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1 $Y=1.875
+ $X2=1.165 $Y2=1.79
r144 25 27 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1 $Y=1.875 $X2=1
+ $Y2=1.98
r145 8 47 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.52
+ $Y=1.835 $X2=3.66 $Y2=1.98
r146 7 41 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=1.835 $X2=2.72 $Y2=1.98
r147 6 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.72
+ $Y=1.835 $X2=1.86 $Y2=1.98
r148 5 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.86
+ $Y=1.835 $X2=1 $Y2=1.98
r149 4 52 182 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.235 $X2=5.75 $Y2=0.86
r150 3 79 182 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_NDIFF $count=1 $X=4.75
+ $Y=0.235 $X2=4.89 $Y2=0.92
r151 2 71 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.325 $X2=3.51 $Y2=0.92
r152 1 81 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=2.51
+ $Y=0.325 $X2=2.65 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_4%VPWR 1 2 3 4 15 21 27 31 34 35 37 38 39 41
+ 49 62 63 66 69
r108 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r109 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r110 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r111 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r112 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r113 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r114 57 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r115 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r116 54 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.65 $Y=3.33
+ $X2=5.485 $Y2=3.33
r117 54 56 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.65 $Y=3.33 $X2=6
+ $Y2=3.33
r118 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 53 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r120 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r121 50 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.79 $Y=3.33
+ $X2=4.625 $Y2=3.33
r122 50 52 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.79 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 49 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.32 $Y=3.33
+ $X2=5.485 $Y2=3.33
r124 49 52 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.32 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 43 47 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r126 43 44 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r127 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.625 $Y2=3.33
r128 41 47 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 39 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r130 39 44 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=0.24 $Y2=3.33
r131 39 47 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 37 59 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.085 $Y=3.33
+ $X2=6.96 $Y2=3.33
r133 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.085 $Y=3.33
+ $X2=7.25 $Y2=3.33
r134 36 62 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=7.415 $Y=3.33
+ $X2=7.92 $Y2=3.33
r135 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.415 $Y=3.33
+ $X2=7.25 $Y2=3.33
r136 34 56 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.225 $Y=3.33
+ $X2=6 $Y2=3.33
r137 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=3.33
+ $X2=6.39 $Y2=3.33
r138 33 59 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.555 $Y=3.33
+ $X2=6.96 $Y2=3.33
r139 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.555 $Y=3.33
+ $X2=6.39 $Y2=3.33
r140 29 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.25 $Y=3.245
+ $X2=7.25 $Y2=3.33
r141 29 31 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=7.25 $Y=3.245
+ $X2=7.25 $Y2=2.385
r142 25 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=3.245
+ $X2=6.39 $Y2=3.33
r143 25 27 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=6.39 $Y=3.245
+ $X2=6.39 $Y2=2.385
r144 21 24 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=5.485 $Y=2.18
+ $X2=5.485 $Y2=2.95
r145 19 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=3.245
+ $X2=5.485 $Y2=3.33
r146 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.485 $Y=3.245
+ $X2=5.485 $Y2=2.95
r147 15 18 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=4.625 $Y=2.18
+ $X2=4.625 $Y2=2.95
r148 13 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=3.33
r149 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=2.95
r150 4 31 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=7.11
+ $Y=1.835 $X2=7.25 $Y2=2.385
r151 3 27 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=6.25
+ $Y=1.835 $X2=6.39 $Y2=2.385
r152 2 24 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.345
+ $Y=1.835 $X2=5.485 $Y2=2.95
r153 2 21 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=5.345
+ $Y=1.835 $X2=5.485 $Y2=2.18
r154 1 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.835 $X2=4.625 $Y2=2.95
r155 1 15 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.835 $X2=4.625 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_4%A_63_65# 1 2 3 4 5 18 20 21 24 26 31 33 34
+ 36 38 41
c54 24 0 1.81325e-19 $X=1.3 $Y=0.48
r55 40 41 6.145 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.445
+ $X2=2.995 $Y2=0.445
r56 34 40 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.375 $Y=0.445
+ $X2=3.08 $Y2=0.445
r57 34 36 17.135 $w=3.78e-07 $l=5.65e-07 $layer=LI1_cond $X=3.375 $Y=0.445
+ $X2=3.94 $Y2=0.445
r58 33 41 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.245 $Y=0.34
+ $X2=2.995 $Y2=0.34
r59 29 31 24.6465 $w=1.78e-07 $l=4e-07 $layer=LI1_cond $X=2.155 $Y=0.87
+ $X2=2.155 $Y2=0.47
r60 28 33 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.155 $Y=0.425
+ $X2=2.245 $Y2=0.34
r61 28 31 2.77273 $w=1.78e-07 $l=4.5e-08 $layer=LI1_cond $X=2.155 $Y=0.425
+ $X2=2.155 $Y2=0.47
r62 27 38 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.395 $Y=0.955
+ $X2=1.3 $Y2=0.955
r63 26 29 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.065 $Y=0.955
+ $X2=2.155 $Y2=0.87
r64 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.065 $Y=0.955
+ $X2=1.395 $Y2=0.955
r65 22 38 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=0.87 $X2=1.3
+ $Y2=0.955
r66 22 24 22.7656 $w=1.88e-07 $l=3.9e-07 $layer=LI1_cond $X=1.3 $Y=0.87 $X2=1.3
+ $Y2=0.48
r67 20 38 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.205 $Y=0.955
+ $X2=1.3 $Y2=0.955
r68 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.205 $Y=0.955
+ $X2=0.535 $Y2=0.955
r69 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.405 $Y=0.87
+ $X2=0.535 $Y2=0.955
r70 16 18 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=0.405 $Y=0.87
+ $X2=0.405 $Y2=0.48
r71 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.8
+ $Y=0.325 $X2=3.94 $Y2=0.47
r72 4 40 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.325 $X2=3.08 $Y2=0.47
r73 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.02
+ $Y=0.325 $X2=2.16 $Y2=0.47
r74 2 24 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=1.16
+ $Y=0.325 $X2=1.3 $Y2=0.48
r75 1 18 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.315
+ $Y=0.325 $X2=0.44 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_4%VGND 1 2 3 4 17 21 25 29 31 33 38 43 50 51
+ 54 57 60 63
r97 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r98 60 61 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r99 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r100 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r101 51 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r102 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r103 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.635 $Y=0 $X2=7.47
+ $Y2=0
r104 48 50 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.635 $Y=0
+ $X2=7.92 $Y2=0
r105 47 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r106 47 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r107 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r108 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.61
+ $Y2=0
r109 44 46 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.775 $Y=0
+ $X2=6.96 $Y2=0
r110 43 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=0 $X2=7.47
+ $Y2=0
r111 43 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.305 $Y=0 $X2=6.96
+ $Y2=0
r112 42 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r113 41 42 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r114 39 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=1.73
+ $Y2=0
r115 39 41 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.895 $Y=0
+ $X2=2.16 $Y2=0
r116 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.61
+ $Y2=0
r117 38 41 279.556 $w=1.68e-07 $l=4.285e-06 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=2.16 $Y2=0
r118 37 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r119 37 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r120 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r121 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.87
+ $Y2=0
r122 34 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r123 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=1.73
+ $Y2=0
r124 33 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=1.2
+ $Y2=0
r125 31 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6.48
+ $Y2=0
r126 31 42 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.16 $Y2=0
r127 27 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=0.085
+ $X2=7.47 $Y2=0
r128 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.47 $Y=0.085
+ $X2=7.47 $Y2=0.38
r129 23 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0
r130 23 25 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0.48
r131 19 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=0.085
+ $X2=1.73 $Y2=0
r132 19 21 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.73 $Y=0.085
+ $X2=1.73 $Y2=0.575
r133 15 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=0.085
+ $X2=0.87 $Y2=0
r134 15 17 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.87 $Y=0.085
+ $X2=0.87 $Y2=0.575
r135 4 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.33
+ $Y=0.235 $X2=7.47 $Y2=0.38
r136 3 25 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=6.47
+ $Y=0.235 $X2=6.61 $Y2=0.48
r137 2 21 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.325 $X2=1.73 $Y2=0.575
r138 1 17 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.73
+ $Y=0.325 $X2=0.87 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_4%A_867_47# 1 2 3 4 5 16 22 23 24 28 30 34 40
c54 30 0 1.39855e-19 $X=7.805 $Y=1.16
r55 43 44 9.4665 $w=2.78e-07 $l=2.3e-07 $layer=LI1_cond $X=6.995 $Y=0.93
+ $X2=6.995 $Y2=1.16
r56 40 43 0.94665 $w=2.78e-07 $l=2.3e-08 $layer=LI1_cond $X=6.995 $Y=0.907
+ $X2=6.995 $Y2=0.93
r57 40 41 6.63022 $w=2.78e-07 $l=1.32e-07 $layer=LI1_cond $X=6.995 $Y=0.907
+ $X2=6.995 $Y2=0.775
r58 32 34 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=7.935 $Y=1.065
+ $X2=7.935 $Y2=0.42
r59 31 44 3.00742 $w=1.9e-07 $l=1.4e-07 $layer=LI1_cond $X=7.135 $Y=1.16
+ $X2=6.995 $Y2=1.16
r60 30 32 7.03324 $w=1.9e-07 $l=1.71026e-07 $layer=LI1_cond $X=7.805 $Y=1.16
+ $X2=7.935 $Y2=1.065
r61 30 31 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=7.805 $Y=1.16
+ $X2=7.135 $Y2=1.16
r62 28 41 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=7.04 $Y=0.42
+ $X2=7.04 $Y2=0.775
r63 25 39 3.38263 $w=2.65e-07 $l=1.3e-07 $layer=LI1_cond $X=6.275 $Y=0.907
+ $X2=6.145 $Y2=0.907
r64 24 40 1.07178 $w=2.65e-07 $l=1.4e-07 $layer=LI1_cond $X=6.855 $Y=0.907
+ $X2=6.995 $Y2=0.907
r65 24 25 25.2233 $w=2.63e-07 $l=5.8e-07 $layer=LI1_cond $X=6.855 $Y=0.907
+ $X2=6.275 $Y2=0.907
r66 23 39 3.43467 $w=2.6e-07 $l=1.32e-07 $layer=LI1_cond $X=6.145 $Y=0.775
+ $X2=6.145 $Y2=0.907
r67 22 37 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=6.145 $Y=0.525
+ $X2=6.145 $Y2=0.4
r68 22 23 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=6.145 $Y=0.525
+ $X2=6.145 $Y2=0.775
r69 18 21 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=4.46 $Y=0.4 $X2=5.32
+ $Y2=0.4
r70 16 37 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=6.015 $Y=0.4
+ $X2=6.145 $Y2=0.4
r71 16 21 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=6.015 $Y=0.4
+ $X2=5.32 $Y2=0.4
r72 5 34 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.76
+ $Y=0.235 $X2=7.9 $Y2=0.42
r73 4 43 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.235 $X2=7.04 $Y2=0.93
r74 4 28 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.9
+ $Y=0.235 $X2=7.04 $Y2=0.42
r75 3 39 182 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.235 $X2=6.18 $Y2=0.875
r76 3 37 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.235 $X2=6.18 $Y2=0.44
r77 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.18
+ $Y=0.235 $X2=5.32 $Y2=0.38
r78 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.335
+ $Y=0.235 $X2=4.46 $Y2=0.38
.ends

