* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_804_39# A2_N a_1235_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND B2 a_35_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 Y a_804_39# a_35_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_1235_65# A2_N a_804_39# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VPWR a_804_39# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_35_65# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR B1 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 Y B2 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_35_65# a_804_39# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR A1_N a_804_39# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_1235_65# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VPWR A2_N a_804_39# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_804_39# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_35_65# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VGND B2 a_35_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VGND A1_N a_1235_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VPWR B1 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_35_65# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_132_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_1235_65# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VGND B1 a_35_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_804_39# A2_N a_1235_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_804_39# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 VPWR A1_N a_804_39# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_804_39# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_132_367# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 VGND A1_N a_1235_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 VGND B1 a_35_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_1235_65# A2_N a_804_39# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 Y a_804_39# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_35_65# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 a_35_65# a_804_39# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 VPWR a_804_39# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 Y a_804_39# a_35_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 Y a_804_39# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 a_132_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 a_804_39# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 a_132_367# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 VPWR A2_N a_804_39# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 Y B2 a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
