* File: sky130_fd_sc_lp__bufinv_8.pex.spice
* Created: Wed Sep  2 09:35:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFINV_8%A_82_23# 1 2 3 4 15 19 23 27 31 35 39 43 47
+ 51 55 59 63 67 71 75 77 84 87 90 92 95 99 101 105 111 113 114 115 116
c161 84 0 1.78595e-19 $X=3.87 $Y=1.49
r162 127 128 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.065 $Y=1.49
+ $X2=3.495 $Y2=1.49
r163 126 127 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.635 $Y=1.49
+ $X2=3.065 $Y2=1.49
r164 125 126 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.205 $Y=1.49
+ $X2=2.635 $Y2=1.49
r165 124 125 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.775 $Y=1.49
+ $X2=2.205 $Y2=1.49
r166 123 124 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.345 $Y=1.49
+ $X2=1.775 $Y2=1.49
r167 119 121 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.485 $Y=1.49
+ $X2=0.915 $Y2=1.49
r168 116 128 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.57 $Y=1.49
+ $X2=3.495 $Y2=1.49
r169 109 111 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=5.1 $Y=1.055
+ $X2=5.1 $Y2=0.48
r170 105 107 40.4636 $w=2.23e-07 $l=7.9e-07 $layer=LI1_cond $X=5.082 $Y=2.05
+ $X2=5.082 $Y2=2.84
r171 103 105 6.40246 $w=2.23e-07 $l=1.25e-07 $layer=LI1_cond $X=5.082 $Y=1.925
+ $X2=5.082 $Y2=2.05
r172 102 115 2.79892 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=4.375 $Y=1.84
+ $X2=4.207 $Y2=1.84
r173 101 103 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.97 $Y=1.84
+ $X2=5.082 $Y2=1.925
r174 101 102 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.97 $Y=1.84
+ $X2=4.375 $Y2=1.84
r175 100 113 2.64776 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.335 $Y=1.14
+ $X2=4.182 $Y2=1.14
r176 99 109 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.005 $Y=1.14
+ $X2=5.1 $Y2=1.055
r177 99 100 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.005 $Y=1.14
+ $X2=4.335 $Y2=1.14
r178 95 97 27.177 $w=3.33e-07 $l=7.9e-07 $layer=LI1_cond $X=4.207 $Y=2.05
+ $X2=4.207 $Y2=2.84
r179 93 115 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=4.207 $Y=1.925
+ $X2=4.207 $Y2=1.84
r180 93 95 4.30016 $w=3.33e-07 $l=1.25e-07 $layer=LI1_cond $X=4.207 $Y=1.925
+ $X2=4.207 $Y2=2.05
r181 92 115 3.67481 $w=2.52e-07 $l=1.19143e-07 $layer=LI1_cond $X=4.125 $Y=1.755
+ $X2=4.207 $Y2=1.84
r182 91 114 5.52892 $w=1.75e-07 $l=9.74679e-08 $layer=LI1_cond $X=4.125 $Y=1.585
+ $X2=4.12 $Y2=1.49
r183 91 92 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.125 $Y=1.585
+ $X2=4.125 $Y2=1.755
r184 90 114 5.52892 $w=1.75e-07 $l=9.5e-08 $layer=LI1_cond $X=4.12 $Y=1.395
+ $X2=4.12 $Y2=1.49
r185 89 113 3.80849 $w=2.42e-07 $l=1.11781e-07 $layer=LI1_cond $X=4.12 $Y=1.225
+ $X2=4.182 $Y2=1.14
r186 89 90 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=4.12 $Y=1.225
+ $X2=4.12 $Y2=1.395
r187 85 113 3.80849 $w=2.42e-07 $l=8.5e-08 $layer=LI1_cond $X=4.182 $Y=1.055
+ $X2=4.182 $Y2=1.14
r188 85 87 21.7264 $w=3.03e-07 $l=5.75e-07 $layer=LI1_cond $X=4.182 $Y=1.055
+ $X2=4.182 $Y2=0.48
r189 84 116 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=3.87 $Y=1.49
+ $X2=3.57 $Y2=1.49
r190 83 84 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=3.87
+ $Y=1.49 $X2=3.87 $Y2=1.49
r191 80 123 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.15 $Y=1.49
+ $X2=1.345 $Y2=1.49
r192 80 121 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.15 $Y=1.49
+ $X2=0.915 $Y2=1.49
r193 79 83 158.775 $w=1.88e-07 $l=2.72e-06 $layer=LI1_cond $X=1.15 $Y=1.49
+ $X2=3.87 $Y2=1.49
r194 79 80 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=1.15
+ $Y=1.49 $X2=1.15 $Y2=1.49
r195 77 114 1.04816 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=4.03 $Y=1.49 $X2=4.12
+ $Y2=1.49
r196 77 83 9.33971 $w=1.88e-07 $l=1.6e-07 $layer=LI1_cond $X=4.03 $Y=1.49
+ $X2=3.87 $Y2=1.49
r197 73 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.655
+ $X2=3.495 $Y2=1.49
r198 73 75 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.495 $Y=1.655
+ $X2=3.495 $Y2=2.465
r199 69 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.325
+ $X2=3.495 $Y2=1.49
r200 69 71 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.495 $Y=1.325
+ $X2=3.495 $Y2=0.665
r201 65 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.655
+ $X2=3.065 $Y2=1.49
r202 65 67 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.065 $Y=1.655
+ $X2=3.065 $Y2=2.465
r203 61 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.325
+ $X2=3.065 $Y2=1.49
r204 61 63 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.065 $Y=1.325
+ $X2=3.065 $Y2=0.665
r205 57 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.655
+ $X2=2.635 $Y2=1.49
r206 57 59 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.635 $Y=1.655
+ $X2=2.635 $Y2=2.465
r207 53 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.325
+ $X2=2.635 $Y2=1.49
r208 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.635 $Y=1.325
+ $X2=2.635 $Y2=0.665
r209 49 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.655
+ $X2=2.205 $Y2=1.49
r210 49 51 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.205 $Y=1.655
+ $X2=2.205 $Y2=2.465
r211 45 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.325
+ $X2=2.205 $Y2=1.49
r212 45 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.205 $Y=1.325
+ $X2=2.205 $Y2=0.665
r213 41 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.655
+ $X2=1.775 $Y2=1.49
r214 41 43 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.775 $Y=1.655
+ $X2=1.775 $Y2=2.465
r215 37 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.325
+ $X2=1.775 $Y2=1.49
r216 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.775 $Y=1.325
+ $X2=1.775 $Y2=0.665
r217 33 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.655
+ $X2=1.345 $Y2=1.49
r218 33 35 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.345 $Y=1.655
+ $X2=1.345 $Y2=2.465
r219 29 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.325
+ $X2=1.345 $Y2=1.49
r220 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.345 $Y=1.325
+ $X2=1.345 $Y2=0.665
r221 25 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.655
+ $X2=0.915 $Y2=1.49
r222 25 27 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.915 $Y=1.655
+ $X2=0.915 $Y2=2.465
r223 21 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.325
+ $X2=0.915 $Y2=1.49
r224 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.915 $Y=1.325
+ $X2=0.915 $Y2=0.665
r225 17 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.655
+ $X2=0.485 $Y2=1.49
r226 17 19 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.485 $Y=1.655
+ $X2=0.485 $Y2=2.465
r227 13 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=1.49
r228 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.485 $Y=1.325
+ $X2=0.485 $Y2=0.665
r229 4 107 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=1.835 $X2=5.1 $Y2=2.84
r230 4 105 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=1.835 $X2=5.1 $Y2=2.05
r231 3 97 400 $w=1.7e-07 $l=1.06567e-06 $layer=licon1_PDIFF $count=1 $X=4.115
+ $Y=1.835 $X2=4.24 $Y2=2.84
r232 3 95 400 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=4.115
+ $Y=1.835 $X2=4.24 $Y2=2.05
r233 2 111 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.96
+ $Y=0.245 $X2=5.1 $Y2=0.48
r234 1 87 91 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=2 $X=4.105
+ $Y=0.245 $X2=4.23 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_8%A_876_23# 1 2 9 13 17 21 25 29 31 40 42 43
+ 44 45 46 49 51 53 55 63
c90 31 0 1.78595e-19 $X=5.385 $Y=1.49
r91 51 57 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.995 $Y=2.14
+ $X2=5.995 $Y2=2.055
r92 51 53 29.9192 $w=2.58e-07 $l=6.75e-07 $layer=LI1_cond $X=5.995 $Y=2.14
+ $X2=5.995 $Y2=2.815
r93 47 49 16.0519 $w=2.78e-07 $l=3.9e-07 $layer=LI1_cond $X=6.005 $Y=0.87
+ $X2=6.005 $Y2=0.48
r94 45 57 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.865 $Y=2.055
+ $X2=5.995 $Y2=2.055
r95 45 46 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.865 $Y=2.055
+ $X2=5.555 $Y2=2.055
r96 43 47 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=5.865 $Y=0.955
+ $X2=6.005 $Y2=0.87
r97 43 44 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.865 $Y=0.955
+ $X2=5.555 $Y2=0.955
r98 42 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.47 $Y=1.97
+ $X2=5.555 $Y2=2.055
r99 41 55 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.47 $Y=1.585
+ $X2=5.47 $Y2=1.49
r100 41 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.47 $Y=1.585
+ $X2=5.47 $Y2=1.97
r101 40 55 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.47 $Y=1.395
+ $X2=5.47 $Y2=1.49
r102 39 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.47 $Y=1.04
+ $X2=5.555 $Y2=0.955
r103 39 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.47 $Y=1.04
+ $X2=5.47 $Y2=1.395
r104 38 63 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.225 $Y=1.49
+ $X2=5.315 $Y2=1.49
r105 38 61 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.225 $Y=1.49
+ $X2=4.885 $Y2=1.49
r106 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.225
+ $Y=1.49 $X2=5.225 $Y2=1.49
r107 34 61 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.545 $Y=1.49
+ $X2=4.885 $Y2=1.49
r108 34 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.545 $Y=1.49
+ $X2=4.455 $Y2=1.49
r109 33 37 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=4.545 $Y=1.49
+ $X2=5.225 $Y2=1.49
r110 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.545
+ $Y=1.49 $X2=4.545 $Y2=1.49
r111 31 55 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=1.49
+ $X2=5.47 $Y2=1.49
r112 31 37 9.33971 $w=1.88e-07 $l=1.6e-07 $layer=LI1_cond $X=5.385 $Y=1.49
+ $X2=5.225 $Y2=1.49
r113 27 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.315 $Y=1.655
+ $X2=5.315 $Y2=1.49
r114 27 29 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.315 $Y=1.655
+ $X2=5.315 $Y2=2.465
r115 23 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.315 $Y=1.325
+ $X2=5.315 $Y2=1.49
r116 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.315 $Y=1.325
+ $X2=5.315 $Y2=0.665
r117 19 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.885 $Y=1.655
+ $X2=4.885 $Y2=1.49
r118 19 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.885 $Y=1.655
+ $X2=4.885 $Y2=2.465
r119 15 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.885 $Y=1.325
+ $X2=4.885 $Y2=1.49
r120 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.885 $Y=1.325
+ $X2=4.885 $Y2=0.665
r121 11 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=1.655
+ $X2=4.455 $Y2=1.49
r122 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.455 $Y=1.655
+ $X2=4.455 $Y2=2.465
r123 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=1.325
+ $X2=4.455 $Y2=1.49
r124 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.455 $Y=1.325
+ $X2=4.455 $Y2=0.665
r125 2 57 400 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.835 $X2=5.96 $Y2=2.135
r126 2 53 400 $w=1.7e-07 $l=1.04766e-06 $layer=licon1_PDIFF $count=1 $X=5.82
+ $Y=1.835 $X2=5.96 $Y2=2.815
r127 1 49 91 $w=1.7e-07 $l=3.04672e-07 $layer=licon1_NDIFF $count=2 $X=5.82
+ $Y=0.245 $X2=5.98 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_8%A 3 6 8 9 13 15
r29 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.835 $Y=1.375
+ $X2=5.835 $Y2=1.54
r30 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.835 $Y=1.375
+ $X2=5.835 $Y2=1.21
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.835
+ $Y=1.375 $X2=5.835 $Y2=1.375
r32 9 14 8.25206 $w=4.03e-07 $l=2.9e-07 $layer=LI1_cond $X=5.952 $Y=1.665
+ $X2=5.952 $Y2=1.375
r33 8 14 2.27643 $w=4.03e-07 $l=8e-08 $layer=LI1_cond $X=5.952 $Y=1.295
+ $X2=5.952 $Y2=1.375
r34 6 16 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=5.745 $Y=2.465
+ $X2=5.745 $Y2=1.54
r35 3 15 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.745 $Y=0.665
+ $X2=5.745 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_8%VPWR 1 2 3 4 5 6 7 22 24 30 36 42 46 50 54
+ 58 64 67 68 70 71 72 73 74 86 93 94 100 103 106
r101 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r102 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r104 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r106 94 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r107 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r108 91 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.695 $Y=3.33
+ $X2=5.53 $Y2=3.33
r109 91 93 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.695 $Y=3.33
+ $X2=6 $Y2=3.33
r110 90 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r111 90 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r113 87 103 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.8 $Y=3.33
+ $X2=4.672 $Y2=3.33
r114 87 89 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r115 86 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=3.33
+ $X2=5.53 $Y2=3.33
r116 86 89 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.365 $Y=3.33
+ $X2=5.04 $Y2=3.33
r117 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r121 79 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r122 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 76 97 4.4377 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.2
+ $Y2=3.33
r124 76 78 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.72
+ $Y2=3.33
r125 74 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r126 74 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r127 72 84 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.72 $Y=3.33 $X2=2.64
+ $Y2=3.33
r128 72 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.72 $Y=3.33
+ $X2=2.85 $Y2=3.33
r129 70 81 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.86 $Y=3.33
+ $X2=1.68 $Y2=3.33
r130 70 71 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.86 $Y=3.33
+ $X2=1.99 $Y2=3.33
r131 69 84 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r132 69 71 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.12 $Y=3.33
+ $X2=1.99 $Y2=3.33
r133 67 78 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r134 67 68 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=1.13
+ $Y2=3.33
r135 66 81 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.26 $Y=3.33
+ $X2=1.68 $Y2=3.33
r136 66 68 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.26 $Y=3.33
+ $X2=1.13 $Y2=3.33
r137 62 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=3.33
r138 62 64 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=2.435
r139 58 61 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=4.672 $Y=2.26
+ $X2=4.672 $Y2=2.94
r140 56 103 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.672 $Y=3.245
+ $X2=4.672 $Y2=3.33
r141 56 61 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=4.672 $Y=3.245
+ $X2=4.672 $Y2=2.94
r142 55 100 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.87 $Y=3.33
+ $X2=3.725 $Y2=3.33
r143 54 103 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=4.672 $Y2=3.33
r144 54 55 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=3.87 $Y2=3.33
r145 50 53 31.3941 $w=2.88e-07 $l=7.9e-07 $layer=LI1_cond $X=3.725 $Y=2.05
+ $X2=3.725 $Y2=2.84
r146 48 100 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=3.245
+ $X2=3.725 $Y2=3.33
r147 48 53 16.0945 $w=2.88e-07 $l=4.05e-07 $layer=LI1_cond $X=3.725 $Y=3.245
+ $X2=3.725 $Y2=2.84
r148 47 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.98 $Y=3.33
+ $X2=2.85 $Y2=3.33
r149 46 100 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.58 $Y=3.33
+ $X2=3.725 $Y2=3.33
r150 46 47 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.58 $Y=3.33 $X2=2.98
+ $Y2=3.33
r151 42 45 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=2.85 $Y=2.26
+ $X2=2.85 $Y2=2.94
r152 40 73 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=3.33
r153 40 45 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=2.94
r154 36 39 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.99 $Y=2.26
+ $X2=1.99 $Y2=2.94
r155 34 71 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=3.33
r156 34 39 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=2.94
r157 30 33 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.13 $Y=2.26
+ $X2=1.13 $Y2=2.94
r158 28 68 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=3.245
+ $X2=1.13 $Y2=3.33
r159 28 33 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.13 $Y=3.245
+ $X2=1.13 $Y2=2.94
r160 24 27 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.252 $Y=2.26
+ $X2=0.252 $Y2=2.94
r161 22 97 3.03982 $w=2.95e-07 $l=1.07912e-07 $layer=LI1_cond $X=0.252 $Y=3.245
+ $X2=0.2 $Y2=3.33
r162 22 27 11.9151 $w=2.93e-07 $l=3.05e-07 $layer=LI1_cond $X=0.252 $Y=3.245
+ $X2=0.252 $Y2=2.94
r163 7 64 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=5.39
+ $Y=1.835 $X2=5.53 $Y2=2.435
r164 6 61 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=4.53
+ $Y=1.835 $X2=4.67 $Y2=2.94
r165 6 58 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=4.53
+ $Y=1.835 $X2=4.67 $Y2=2.26
r166 5 53 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=1.835 $X2=3.71 $Y2=2.84
r167 5 50 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=1.835 $X2=3.71 $Y2=2.05
r168 4 45 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.835 $X2=2.85 $Y2=2.94
r169 4 42 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.835 $X2=2.85 $Y2=2.26
r170 3 39 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.835 $X2=1.99 $Y2=2.94
r171 3 36 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.835 $X2=1.99 $Y2=2.26
r172 2 33 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=2.94
r173 2 30 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=2.26
r174 1 27 400 $w=1.7e-07 $l=1.16583e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.94
r175 1 24 400 $w=1.7e-07 $l=4.83477e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_8%Y 1 2 3 4 5 6 7 8 27 29 31 35 37 41 45 49
+ 51 55 59 63 65 69 73 77 78 79 80 81 82
r93 82 96 3.19611 $w=6.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.462 $Y=1.665
+ $X2=0.462 $Y2=1.84
r94 81 82 6.75748 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.462 $Y=1.295
+ $X2=0.462 $Y2=1.665
r95 73 75 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=3.28 $Y=2.05
+ $X2=3.28 $Y2=2.84
r96 71 73 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=3.28 $Y=1.925
+ $X2=3.28 $Y2=2.05
r97 67 69 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=3.28 $Y=1.055
+ $X2=3.28 $Y2=0.48
r98 66 80 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.55 $Y=1.84 $X2=2.42
+ $Y2=1.84
r99 65 71 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.15 $Y=1.84
+ $X2=3.28 $Y2=1.925
r100 65 66 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.15 $Y=1.84 $X2=2.55
+ $Y2=1.84
r101 64 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.55 $Y=1.14
+ $X2=2.42 $Y2=1.14
r102 63 67 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.15 $Y=1.14
+ $X2=3.28 $Y2=1.055
r103 63 64 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.15 $Y=1.14 $X2=2.55
+ $Y2=1.14
r104 59 61 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=2.42 $Y=2.05
+ $X2=2.42 $Y2=2.84
r105 57 80 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=1.925
+ $X2=2.42 $Y2=1.84
r106 57 59 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=2.42 $Y=1.925
+ $X2=2.42 $Y2=2.05
r107 53 79 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=1.055
+ $X2=2.42 $Y2=1.14
r108 53 55 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=2.42 $Y=1.055
+ $X2=2.42 $Y2=0.48
r109 52 78 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.69 $Y=1.84
+ $X2=1.56 $Y2=1.84
r110 51 80 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.29 $Y=1.84
+ $X2=2.42 $Y2=1.84
r111 51 52 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.29 $Y=1.84 $X2=1.69
+ $Y2=1.84
r112 50 77 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.69 $Y=1.14
+ $X2=1.56 $Y2=1.14
r113 49 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.29 $Y=1.14
+ $X2=2.42 $Y2=1.14
r114 49 50 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.29 $Y=1.14 $X2=1.69
+ $Y2=1.14
r115 45 47 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=1.56 $Y=2.05
+ $X2=1.56 $Y2=2.84
r116 43 78 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=1.925
+ $X2=1.56 $Y2=1.84
r117 43 45 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=1.56 $Y=1.925
+ $X2=1.56 $Y2=2.05
r118 39 77 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=1.055
+ $X2=1.56 $Y2=1.14
r119 39 41 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=1.56 $Y=1.055
+ $X2=1.56 $Y2=0.48
r120 38 96 9.01427 $w=1.7e-07 $l=3.68e-07 $layer=LI1_cond $X=0.83 $Y=1.84
+ $X2=0.462 $Y2=1.84
r121 37 78 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.43 $Y=1.84
+ $X2=1.56 $Y2=1.84
r122 37 38 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.43 $Y=1.84 $X2=0.83
+ $Y2=1.84
r123 36 81 2.83084 $w=6.68e-07 $l=4.38707e-07 $layer=LI1_cond $X=0.83 $Y=1.14
+ $X2=0.462 $Y2=1.295
r124 35 77 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.43 $Y=1.14
+ $X2=1.56 $Y2=1.14
r125 35 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.43 $Y=1.14 $X2=0.83
+ $Y2=1.14
r126 31 33 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=0.7 $Y=2.05 $X2=0.7
+ $Y2=2.84
r127 29 96 6.27933 $w=6.68e-07 $l=2.77262e-07 $layer=LI1_cond $X=0.7 $Y=1.925
+ $X2=0.462 $Y2=1.84
r128 29 31 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.7 $Y=1.925
+ $X2=0.7 $Y2=2.05
r129 25 36 6.27933 $w=6.68e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.7 $Y=1.055
+ $X2=0.83 $Y2=1.14
r130 25 27 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=0.7 $Y=1.055
+ $X2=0.7 $Y2=0.48
r131 8 75 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.835 $X2=3.28 $Y2=2.84
r132 8 73 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.835 $X2=3.28 $Y2=2.05
r133 7 61 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=2.84
r134 7 59 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=2.05
r135 6 47 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.835 $X2=1.56 $Y2=2.84
r136 6 45 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.835 $X2=1.56 $Y2=2.05
r137 5 33 400 $w=1.7e-07 $l=1.07272e-06 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=2.84
r138 5 31 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=2.05
r139 4 69 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=3.14
+ $Y=0.245 $X2=3.28 $Y2=0.48
r140 3 55 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=2.28
+ $Y=0.245 $X2=2.42 $Y2=0.48
r141 2 41 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=1.42
+ $Y=0.245 $X2=1.56 $Y2=0.48
r142 1 27 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.245 $X2=0.7 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__BUFINV_8%VGND 1 2 3 4 5 6 7 22 24 28 32 36 38 42 44
+ 48 52 55 56 58 59 60 61 62 74 81 82 88 91 94
r100 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r101 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r102 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r103 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r104 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r105 82 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r106 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r107 79 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.695 $Y=0 $X2=5.53
+ $Y2=0
r108 79 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.695 $Y=0 $X2=6
+ $Y2=0
r109 78 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r110 78 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r111 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r112 75 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=4.67
+ $Y2=0
r113 75 77 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=5.04 $Y2=0
r114 74 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=0 $X2=5.53
+ $Y2=0
r115 74 77 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.365 $Y=0
+ $X2=5.04 $Y2=0
r116 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r117 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r118 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r119 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r120 67 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r121 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r122 64 85 4.4377 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.2 $Y2=0
r123 64 66 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.72
+ $Y2=0
r124 62 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r125 62 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r126 60 72 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.64
+ $Y2=0
r127 60 61 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.85
+ $Y2=0
r128 58 69 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.68
+ $Y2=0
r129 58 59 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.99
+ $Y2=0
r130 57 72 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.64
+ $Y2=0
r131 57 59 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=1.99
+ $Y2=0
r132 55 66 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.72
+ $Y2=0
r133 55 56 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1 $Y=0 $X2=1.13
+ $Y2=0
r134 54 69 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.68
+ $Y2=0
r135 54 56 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.13
+ $Y2=0
r136 50 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=0.085
+ $X2=5.53 $Y2=0
r137 50 52 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.53 $Y=0.085
+ $X2=5.53 $Y2=0.535
r138 46 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.67 $Y2=0
r139 46 48 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.67 $Y=0.085
+ $X2=4.67 $Y2=0.42
r140 45 88 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.86 $Y=0 $X2=3.72
+ $Y2=0
r141 44 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.505 $Y=0 $X2=4.67
+ $Y2=0
r142 44 45 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.505 $Y=0
+ $X2=3.86 $Y2=0
r143 40 88 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0
r144 40 42 16.2577 $w=2.78e-07 $l=3.95e-07 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0.48
r145 39 61 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.98 $Y=0 $X2=2.85
+ $Y2=0
r146 38 88 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=3.72
+ $Y2=0
r147 38 39 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=2.98
+ $Y2=0
r148 34 61 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=0.085
+ $X2=2.85 $Y2=0
r149 34 36 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=2.85 $Y=0.085
+ $X2=2.85 $Y2=0.37
r150 30 59 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0
r151 30 32 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0.37
r152 26 56 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.13 $Y2=0
r153 26 28 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.13 $Y2=0.37
r154 22 85 3.03982 $w=2.95e-07 $l=1.07912e-07 $layer=LI1_cond $X=0.252 $Y=0.085
+ $X2=0.2 $Y2=0
r155 22 24 15.6263 $w=2.93e-07 $l=4e-07 $layer=LI1_cond $X=0.252 $Y=0.085
+ $X2=0.252 $Y2=0.485
r156 7 52 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=5.39
+ $Y=0.245 $X2=5.53 $Y2=0.535
r157 6 48 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=4.53
+ $Y=0.245 $X2=4.67 $Y2=0.42
r158 5 42 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=3.57
+ $Y=0.245 $X2=3.71 $Y2=0.48
r159 4 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.71
+ $Y=0.245 $X2=2.85 $Y2=0.37
r160 3 32 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.85
+ $Y=0.245 $X2=1.99 $Y2=0.37
r161 2 28 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.99
+ $Y=0.245 $X2=1.13 $Y2=0.37
r162 1 24 91 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.245 $X2=0.27 $Y2=0.485
.ends

