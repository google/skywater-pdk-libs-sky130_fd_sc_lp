* File: sky130_fd_sc_lp__nor4_m.pxi.spice
* Created: Wed Sep  2 10:10:47 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4_M%A N_A_M1003_g N_A_c_65_n N_A_M1002_g N_A_c_62_n
+ N_A_c_68_n N_A_c_69_n A A N_A_c_64_n PM_SKY130_FD_SC_LP__NOR4_M%A
x_PM_SKY130_FD_SC_LP__NOR4_M%B N_B_M1004_g N_B_M1005_g N_B_c_101_n N_B_c_106_n B
+ B N_B_c_103_n PM_SKY130_FD_SC_LP__NOR4_M%B
x_PM_SKY130_FD_SC_LP__NOR4_M%C N_C_M1000_g N_C_M1006_g N_C_c_139_n N_C_c_144_n C
+ C N_C_c_141_n PM_SKY130_FD_SC_LP__NOR4_M%C
x_PM_SKY130_FD_SC_LP__NOR4_M%D N_D_M1001_g N_D_M1007_g N_D_c_175_n N_D_c_181_n D
+ D D N_D_c_177_n N_D_c_178_n PM_SKY130_FD_SC_LP__NOR4_M%D
x_PM_SKY130_FD_SC_LP__NOR4_M%VPWR N_VPWR_M1002_s N_VPWR_c_210_n N_VPWR_c_211_n
+ N_VPWR_c_212_n VPWR N_VPWR_c_213_n N_VPWR_c_209_n
+ PM_SKY130_FD_SC_LP__NOR4_M%VPWR
x_PM_SKY130_FD_SC_LP__NOR4_M%Y N_Y_M1003_d N_Y_M1006_d N_Y_M1001_d N_Y_c_228_n
+ N_Y_c_235_n N_Y_c_236_n N_Y_c_229_n N_Y_c_237_n N_Y_c_230_n N_Y_c_231_n Y Y Y
+ N_Y_c_233_n PM_SKY130_FD_SC_LP__NOR4_M%Y
x_PM_SKY130_FD_SC_LP__NOR4_M%VGND N_VGND_M1003_s N_VGND_M1004_d N_VGND_M1007_d
+ N_VGND_c_287_n N_VGND_c_288_n N_VGND_c_289_n N_VGND_c_290_n N_VGND_c_291_n
+ N_VGND_c_292_n VGND N_VGND_c_293_n N_VGND_c_294_n N_VGND_c_295_n
+ N_VGND_c_296_n PM_SKY130_FD_SC_LP__NOR4_M%VGND
cc_1 VNB N_A_M1003_g 0.0383435f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.56
cc_2 VNB N_A_c_62_n 0.0209276f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.695
cc_3 VNB A 0.00498258f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_c_64_n 0.0164912f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_5 VNB N_B_M1004_g 0.035968f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.56
cc_6 VNB N_B_c_101_n 0.0192517f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_7 VNB B 0.00503411f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.695
cc_8 VNB N_B_c_103_n 0.0156645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C_M1006_g 0.0367492f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.25
cc_10 VNB N_C_c_139_n 0.0211789f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_11 VNB C 5.64814e-19 $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.695
cc_12 VNB N_C_c_141_n 0.0165486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D_c_175_n 0.00582141f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.625
cc_14 VNB D 0.0373555f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.86
cc_15 VNB N_D_c_177_n 0.102718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_D_c_178_n 0.0205615f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_17 VNB N_VPWR_c_209_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_228_n 0.0307677f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_19 VNB N_Y_c_229_n 0.0014249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_230_n 0.0113044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_231_n 0.0288592f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_22 VNB Y 0.014688f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_23 VNB N_Y_c_233_n 6.59409e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_287_n 0.0140554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_288_n 0.0101417f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.19
cc_26 VNB N_VGND_c_289_n 0.00580139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_290_n 0.0107763f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_28 VNB N_VGND_c_291_n 0.0244031f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_29 VNB N_VGND_c_292_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_30 VNB N_VGND_c_293_n 0.0187737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_294_n 0.0153494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_295_n 0.185801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_296_n 0.00601391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_A_c_65_n 0.0151477f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.1
cc_35 VPB N_A_M1002_g 0.0242967f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.625
cc_36 VPB N_A_c_62_n 0.00272969f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.695
cc_37 VPB N_A_c_68_n 0.0165105f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.86
cc_38 VPB N_A_c_69_n 0.0226514f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.175
cc_39 VPB A 0.00302965f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_40 VPB N_B_M1005_g 0.038722f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.25
cc_41 VPB N_B_c_101_n 0.00251109f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.355
cc_42 VPB N_B_c_106_n 0.0155932f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.19
cc_43 VPB B 0.00273855f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.695
cc_44 VPB N_C_M1000_g 0.0387014f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.56
cc_45 VPB N_C_c_139_n 0.00276247f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.355
cc_46 VPB N_C_c_144_n 0.0166881f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.19
cc_47 VPB C 0.00112272f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.695
cc_48 VPB N_D_M1001_g 0.0234165f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.56
cc_49 VPB N_D_c_175_n 0.0339174f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.625
cc_50 VPB N_D_c_181_n 0.0224131f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.19
cc_51 VPB D 0.01745f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.86
cc_52 VPB N_VPWR_c_210_n 0.0233609f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.1
cc_53 VPB N_VPWR_c_211_n 0.0172587f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.625
cc_54 VPB N_VPWR_c_212_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_213_n 0.0707465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_209_n 0.125398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_228_n 0.0194385f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.355
cc_58 VPB N_Y_c_235_n 0.0701733f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.19
cc_59 VPB N_Y_c_236_n 0.0148348f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.695
cc_60 VPB N_Y_c_237_n 0.0109251f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_61 N_A_M1003_g N_B_M1004_g 0.0285099f $X=0.615 $Y=0.56 $X2=0 $Y2=0
cc_62 N_A_c_65_n N_B_M1005_g 0.00797626f $X=0.615 $Y=2.1 $X2=0 $Y2=0
cc_63 N_A_c_69_n N_B_M1005_g 0.0476886f $X=0.795 $Y=2.175 $X2=0 $Y2=0
cc_64 N_A_c_62_n N_B_c_101_n 0.0116511f $X=0.525 $Y=1.695 $X2=0 $Y2=0
cc_65 N_A_c_68_n N_B_c_106_n 0.0116511f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_66 A B 0.0458013f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A_c_64_n B 6.16665e-19 $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_68 A N_B_c_103_n 0.00481894f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_c_64_n N_B_c_103_n 0.0116511f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_70 N_A_M1002_g N_VPWR_c_210_n 0.00624048f $X=0.795 $Y=2.625 $X2=0 $Y2=0
cc_71 N_A_c_69_n N_VPWR_c_210_n 0.0040175f $X=0.795 $Y=2.175 $X2=0 $Y2=0
cc_72 N_A_M1002_g N_VPWR_c_213_n 0.00490845f $X=0.795 $Y=2.625 $X2=0 $Y2=0
cc_73 N_A_M1002_g N_VPWR_c_209_n 0.00506877f $X=0.795 $Y=2.625 $X2=0 $Y2=0
cc_74 N_A_M1003_g N_Y_c_228_n 0.00544769f $X=0.615 $Y=0.56 $X2=0 $Y2=0
cc_75 N_A_c_65_n N_Y_c_228_n 0.0059042f $X=0.615 $Y=2.1 $X2=0 $Y2=0
cc_76 A N_Y_c_228_n 0.0485272f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_64_n N_Y_c_228_n 0.0163648f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_78 N_A_c_65_n N_Y_c_235_n 0.00443396f $X=0.615 $Y=2.1 $X2=0 $Y2=0
cc_79 N_A_c_68_n N_Y_c_235_n 0.00391136f $X=0.525 $Y=1.86 $X2=0 $Y2=0
cc_80 N_A_c_69_n N_Y_c_235_n 0.019341f $X=0.795 $Y=2.175 $X2=0 $Y2=0
cc_81 A N_Y_c_235_n 0.0260653f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_M1003_g Y 0.0123502f $X=0.615 $Y=0.56 $X2=0 $Y2=0
cc_83 A Y 0.0288881f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_84 N_A_c_64_n Y 0.00397544f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_Y_c_233_n 0.0121552f $X=0.615 $Y=0.56 $X2=0 $Y2=0
cc_86 N_A_M1003_g N_VGND_c_288_n 0.00495038f $X=0.615 $Y=0.56 $X2=0 $Y2=0
cc_87 N_A_M1003_g N_VGND_c_289_n 6.63511e-19 $X=0.615 $Y=0.56 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_VGND_c_293_n 0.00420318f $X=0.615 $Y=0.56 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VGND_c_295_n 0.00485886f $X=0.615 $Y=0.56 $X2=0 $Y2=0
cc_90 N_B_M1005_g N_C_M1000_g 0.024831f $X=1.185 $Y=2.625 $X2=0 $Y2=0
cc_91 N_B_M1004_g N_C_M1006_g 0.0178636f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_92 N_B_c_101_n N_C_c_139_n 0.024831f $X=1.095 $Y=1.695 $X2=0 $Y2=0
cc_93 N_B_c_106_n N_C_c_144_n 0.024831f $X=1.095 $Y=1.86 $X2=0 $Y2=0
cc_94 B C 0.0332503f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_95 N_B_c_103_n C 7.33711e-19 $X=1.095 $Y=1.355 $X2=0 $Y2=0
cc_96 B N_C_c_141_n 0.00460798f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_97 N_B_c_103_n N_C_c_141_n 0.024831f $X=1.095 $Y=1.355 $X2=0 $Y2=0
cc_98 N_B_M1005_g N_VPWR_c_213_n 0.00490845f $X=1.185 $Y=2.625 $X2=0 $Y2=0
cc_99 N_B_M1005_g N_VPWR_c_209_n 0.00506877f $X=1.185 $Y=2.625 $X2=0 $Y2=0
cc_100 N_B_M1005_g N_Y_c_235_n 0.0148742f $X=1.185 $Y=2.625 $X2=0 $Y2=0
cc_101 N_B_c_106_n N_Y_c_235_n 0.00392628f $X=1.095 $Y=1.86 $X2=0 $Y2=0
cc_102 B N_Y_c_235_n 0.0191767f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B_M1004_g N_Y_c_231_n 0.0140215f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_104 B N_Y_c_231_n 0.0205626f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B_c_103_n N_Y_c_231_n 0.00236831f $X=1.095 $Y=1.355 $X2=0 $Y2=0
cc_106 N_B_c_103_n Y 2.31676e-19 $X=1.095 $Y=1.355 $X2=0 $Y2=0
cc_107 N_B_M1004_g N_Y_c_233_n 0.00186443f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_VGND_c_289_n 0.00743985f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_109 N_B_M1004_g N_VGND_c_293_n 0.00460631f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_110 N_B_M1004_g N_VGND_c_295_n 0.00460842f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_111 N_C_M1000_g N_D_c_175_n 0.00799385f $X=1.575 $Y=2.625 $X2=0 $Y2=0
cc_112 N_C_c_139_n N_D_c_175_n 0.0189157f $X=1.665 $Y=1.695 $X2=0 $Y2=0
cc_113 N_C_M1000_g N_D_c_181_n 0.0474257f $X=1.575 $Y=2.625 $X2=0 $Y2=0
cc_114 N_C_M1006_g D 6.87217e-19 $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_115 C D 0.0139304f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_116 N_C_c_141_n D 8.16289e-19 $X=1.665 $Y=1.355 $X2=0 $Y2=0
cc_117 C N_D_c_177_n 0.00286186f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_118 N_C_c_141_n N_D_c_177_n 0.0189157f $X=1.665 $Y=1.355 $X2=0 $Y2=0
cc_119 N_C_M1006_g N_D_c_178_n 0.0284996f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_120 N_C_M1000_g N_VPWR_c_213_n 0.00490845f $X=1.575 $Y=2.625 $X2=0 $Y2=0
cc_121 N_C_M1000_g N_VPWR_c_209_n 0.00506877f $X=1.575 $Y=2.625 $X2=0 $Y2=0
cc_122 N_C_M1000_g N_Y_c_235_n 0.0172693f $X=1.575 $Y=2.625 $X2=0 $Y2=0
cc_123 N_C_c_144_n N_Y_c_235_n 0.00342161f $X=1.665 $Y=1.86 $X2=0 $Y2=0
cc_124 C N_Y_c_235_n 0.0129003f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_C_M1006_g N_Y_c_229_n 0.0017418f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_126 N_C_M1006_g N_Y_c_231_n 0.0133464f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_127 C N_Y_c_231_n 0.0135179f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_128 N_C_c_141_n N_Y_c_231_n 0.00536932f $X=1.665 $Y=1.355 $X2=0 $Y2=0
cc_129 N_C_M1006_g N_VGND_c_289_n 0.00730912f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_130 N_C_M1006_g N_VGND_c_291_n 0.00478016f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_131 N_C_M1006_g N_VGND_c_295_n 0.00510824f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_132 N_D_M1001_g N_VPWR_c_213_n 0.00490845f $X=1.965 $Y=2.625 $X2=0 $Y2=0
cc_133 N_D_M1001_g N_VPWR_c_209_n 0.00506877f $X=1.965 $Y=2.625 $X2=0 $Y2=0
cc_134 N_D_c_175_n N_Y_c_235_n 0.00948571f $X=2.145 $Y=2.1 $X2=0 $Y2=0
cc_135 N_D_c_181_n N_Y_c_235_n 0.017621f $X=2.145 $Y=2.175 $X2=0 $Y2=0
cc_136 N_D_c_177_n N_Y_c_235_n 0.0021957f $X=2.495 $Y=1.045 $X2=0 $Y2=0
cc_137 N_D_c_178_n N_Y_c_229_n 0.0017418f $X=2.365 $Y=0.88 $X2=0 $Y2=0
cc_138 N_D_M1001_g N_Y_c_237_n 0.0076447f $X=1.965 $Y=2.625 $X2=0 $Y2=0
cc_139 N_D_c_181_n N_Y_c_237_n 0.00442092f $X=2.145 $Y=2.175 $X2=0 $Y2=0
cc_140 D N_Y_c_231_n 0.00808349f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_141 N_D_c_178_n N_Y_c_231_n 0.00233f $X=2.365 $Y=0.88 $X2=0 $Y2=0
cc_142 D N_VGND_c_290_n 0.00453639f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_143 N_D_c_177_n N_VGND_c_290_n 0.00693862f $X=2.495 $Y=1.045 $X2=0 $Y2=0
cc_144 N_D_c_178_n N_VGND_c_290_n 0.00512127f $X=2.365 $Y=0.88 $X2=0 $Y2=0
cc_145 N_D_c_178_n N_VGND_c_291_n 0.00478016f $X=2.365 $Y=0.88 $X2=0 $Y2=0
cc_146 D N_VGND_c_295_n 0.0104502f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_147 N_D_c_177_n N_VGND_c_295_n 8.89559e-19 $X=2.495 $Y=1.045 $X2=0 $Y2=0
cc_148 N_D_c_178_n N_VGND_c_295_n 0.00960025f $X=2.365 $Y=0.88 $X2=0 $Y2=0
cc_149 N_VPWR_c_210_n N_Y_c_235_n 0.0163208f $X=0.58 $Y=2.63 $X2=0 $Y2=0
cc_150 N_VPWR_c_213_n N_Y_c_237_n 0.00598543f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_151 N_VPWR_c_209_n N_Y_c_237_n 0.00703216f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_152 N_Y_c_230_n N_VGND_c_288_n 0.00119831f $X=0.26 $Y=0.925 $X2=0 $Y2=0
cc_153 Y N_VGND_c_288_n 0.0149451f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_154 N_Y_c_233_n N_VGND_c_288_n 0.0142489f $X=0.83 $Y=0.625 $X2=0 $Y2=0
cc_155 N_Y_c_231_n N_VGND_c_289_n 0.0179657f $X=1.825 $Y=0.925 $X2=0 $Y2=0
cc_156 N_Y_c_229_n N_VGND_c_291_n 0.00554182f $X=1.93 $Y=0.625 $X2=0 $Y2=0
cc_157 N_Y_c_233_n N_VGND_c_293_n 0.00760797f $X=0.83 $Y=0.625 $X2=0 $Y2=0
cc_158 N_Y_c_229_n N_VGND_c_295_n 0.00709428f $X=1.93 $Y=0.625 $X2=0 $Y2=0
cc_159 N_Y_c_230_n N_VGND_c_295_n 0.00620348f $X=0.26 $Y=0.925 $X2=0 $Y2=0
cc_160 N_Y_c_231_n N_VGND_c_295_n 0.0184947f $X=1.825 $Y=0.925 $X2=0 $Y2=0
cc_161 Y N_VGND_c_295_n 0.00619742f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_162 N_Y_c_233_n N_VGND_c_295_n 0.00988127f $X=0.83 $Y=0.625 $X2=0 $Y2=0
