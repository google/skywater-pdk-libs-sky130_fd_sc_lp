* File: sky130_fd_sc_lp__nand3_1.pxi.spice
* Created: Wed Sep  2 10:04:09 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3_1%C N_C_M1005_g N_C_M1000_g C C N_C_c_36_n
+ N_C_c_37_n PM_SKY130_FD_SC_LP__NAND3_1%C
x_PM_SKY130_FD_SC_LP__NAND3_1%B N_B_M1004_g N_B_M1002_g B B B B N_B_c_64_n
+ N_B_c_65_n PM_SKY130_FD_SC_LP__NAND3_1%B
x_PM_SKY130_FD_SC_LP__NAND3_1%A N_A_M1003_g N_A_M1001_g A A A A N_A_c_100_n
+ N_A_c_101_n PM_SKY130_FD_SC_LP__NAND3_1%A
x_PM_SKY130_FD_SC_LP__NAND3_1%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_c_131_n
+ N_VPWR_c_132_n N_VPWR_c_133_n N_VPWR_c_134_n VPWR N_VPWR_c_135_n
+ N_VPWR_c_130_n N_VPWR_c_137_n PM_SKY130_FD_SC_LP__NAND3_1%VPWR
x_PM_SKY130_FD_SC_LP__NAND3_1%Y N_Y_M1003_d N_Y_M1000_d N_Y_M1001_d N_Y_c_159_n
+ Y Y Y N_Y_c_167_n N_Y_c_165_n N_Y_c_162_n PM_SKY130_FD_SC_LP__NAND3_1%Y
x_PM_SKY130_FD_SC_LP__NAND3_1%VGND N_VGND_M1005_s N_VGND_c_193_n N_VGND_c_194_n
+ VGND N_VGND_c_195_n N_VGND_c_196_n PM_SKY130_FD_SC_LP__NAND3_1%VGND
cc_1 VNB C 0.029426f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_2 VNB N_C_c_36_n 0.0295893f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.495
cc_3 VNB N_C_c_37_n 0.0180641f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.33
cc_4 VNB B 0.00264738f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_B_c_64_n 0.0260631f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.495
cc_6 VNB N_B_c_65_n 0.0169729f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.33
cc_7 VNB A 0.00380079f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_A_c_100_n 0.0296845f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.495
cc_9 VNB N_A_c_101_n 0.0215435f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.33
cc_10 VNB N_VPWR_c_130_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_Y_c_159_n 0.0658098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_193_n 0.0164093f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.66
cc_13 VNB N_VGND_c_194_n 0.036195f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.465
cc_14 VNB N_VGND_c_195_n 0.0535523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_196_n 0.190065f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.495
cc_16 VPB N_C_M1000_g 0.0255266f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_17 VPB C 0.017288f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_18 VPB N_C_c_36_n 0.00552203f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.495
cc_19 VPB N_B_M1002_g 0.0207635f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_20 VPB B 0.00249382f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_21 VPB N_B_c_64_n 0.00543356f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.495
cc_22 VPB N_A_M1001_g 0.0246051f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.465
cc_23 VPB A 0.00239288f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_24 VPB N_A_c_100_n 0.00525405f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.495
cc_25 VPB N_VPWR_c_131_n 0.0138386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_VPWR_c_132_n 0.0493047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_133_n 0.0186115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_134_n 0.00557173f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.495
cc_29 VPB N_VPWR_c_135_n 0.024782f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_130_n 0.0514474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_137_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_Y_c_159_n 0.01619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB Y 0.0111971f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.495
cc_34 VPB N_Y_c_162_n 0.0549716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 N_C_M1000_g N_B_M1002_g 0.0200852f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_36 C N_B_M1002_g 6.12626e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_37 C B 0.0451321f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_38 N_C_c_37_n B 0.00315199f $X=0.54 $Y=1.33 $X2=0 $Y2=0
cc_39 N_C_c_36_n N_B_c_64_n 0.0356066f $X=0.54 $Y=1.495 $X2=0 $Y2=0
cc_40 C N_B_c_65_n 0.00336484f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_41 N_C_c_37_n N_B_c_65_n 0.0356066f $X=0.54 $Y=1.33 $X2=0 $Y2=0
cc_42 N_C_M1000_g N_VPWR_c_132_n 0.00935083f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_43 C N_VPWR_c_132_n 0.0223692f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_44 N_C_c_36_n N_VPWR_c_132_n 5.61224e-19 $X=0.54 $Y=1.495 $X2=0 $Y2=0
cc_45 N_C_M1000_g N_VPWR_c_133_n 0.00480635f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_46 N_C_M1000_g N_VPWR_c_130_n 0.00929616f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_47 N_C_M1000_g Y 0.0037434f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_48 C Y 0.0166818f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_49 N_C_M1000_g N_Y_c_165_n 0.0150994f $X=0.63 $Y=2.465 $X2=0 $Y2=0
cc_50 C N_VGND_M1005_s 0.00234692f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_51 C N_VGND_c_194_n 0.0228747f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_52 N_C_c_36_n N_VGND_c_194_n 9.19692e-19 $X=0.54 $Y=1.495 $X2=0 $Y2=0
cc_53 N_C_c_37_n N_VGND_c_194_n 0.0168001f $X=0.54 $Y=1.33 $X2=0 $Y2=0
cc_54 N_C_c_37_n N_VGND_c_195_n 0.0047441f $X=0.54 $Y=1.33 $X2=0 $Y2=0
cc_55 N_C_c_37_n N_VGND_c_196_n 0.00455844f $X=0.54 $Y=1.33 $X2=0 $Y2=0
cc_56 C A_141_76# 0.00415592f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_57 N_B_M1002_g N_A_M1001_g 0.0257814f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_58 N_B_M1002_g A 2.04582e-19 $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_59 B A 0.0729499f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_60 N_B_c_64_n A 9.1409e-19 $X=1.11 $Y=1.495 $X2=0 $Y2=0
cc_61 N_B_c_65_n A 7.11459e-19 $X=1.11 $Y=1.33 $X2=0 $Y2=0
cc_62 N_B_c_64_n N_A_c_100_n 0.0181513f $X=1.11 $Y=1.495 $X2=0 $Y2=0
cc_63 B N_A_c_101_n 0.00476121f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_64 N_B_c_65_n N_A_c_101_n 0.0297886f $X=1.11 $Y=1.33 $X2=0 $Y2=0
cc_65 N_B_M1002_g N_VPWR_c_133_n 0.00571722f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_66 N_B_M1002_g N_VPWR_c_134_n 0.00412705f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_67 N_B_M1002_g N_VPWR_c_130_n 0.0105533f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_68 N_B_M1002_g Y 6.36733e-19 $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_69 N_B_M1002_g N_Y_c_167_n 0.0146313f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_70 B N_Y_c_167_n 0.0234085f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_71 N_B_c_64_n N_Y_c_167_n 6.81338e-19 $X=1.11 $Y=1.495 $X2=0 $Y2=0
cc_72 N_B_M1002_g N_Y_c_165_n 0.0120157f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_73 B N_VGND_c_194_n 0.019207f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_74 N_B_c_65_n N_VGND_c_194_n 0.00263969f $X=1.11 $Y=1.33 $X2=0 $Y2=0
cc_75 B N_VGND_c_195_n 0.00818334f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_76 N_B_c_65_n N_VGND_c_195_n 0.00500936f $X=1.11 $Y=1.33 $X2=0 $Y2=0
cc_77 B N_VGND_c_196_n 0.010622f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_78 N_B_c_65_n N_VGND_c_196_n 0.00542671f $X=1.11 $Y=1.33 $X2=0 $Y2=0
cc_79 B A_219_76# 0.0113912f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_80 N_A_M1001_g N_VPWR_c_134_n 0.00420957f $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_81 N_A_M1001_g N_VPWR_c_135_n 0.00585385f $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A_M1001_g N_VPWR_c_130_n 0.0120969f $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_83 A N_Y_M1003_d 0.00870458f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_84 N_A_M1001_g N_Y_c_159_n 0.00498464f $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_85 A N_Y_c_159_n 0.102103f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_86 N_A_c_100_n N_Y_c_159_n 0.00830671f $X=1.68 $Y=1.495 $X2=0 $Y2=0
cc_87 N_A_c_101_n N_Y_c_159_n 0.00879565f $X=1.68 $Y=1.33 $X2=0 $Y2=0
cc_88 A Y 0.0065314f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_89 N_A_c_100_n Y 0.00374652f $X=1.68 $Y=1.495 $X2=0 $Y2=0
cc_90 N_A_M1001_g N_Y_c_167_n 0.0144661f $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_91 A N_Y_c_167_n 0.0117073f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_92 N_A_M1001_g N_Y_c_165_n 4.85002e-19 $X=1.59 $Y=2.465 $X2=0 $Y2=0
cc_93 A N_VGND_c_195_n 0.00627065f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_94 N_A_c_101_n N_VGND_c_195_n 0.00418753f $X=1.68 $Y=1.33 $X2=0 $Y2=0
cc_95 A N_VGND_c_196_n 0.00848957f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_96 N_A_c_101_n N_VGND_c_196_n 0.00542671f $X=1.68 $Y=1.33 $X2=0 $Y2=0
cc_97 N_VPWR_c_130_n N_Y_M1000_d 0.00223559f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_98 N_VPWR_c_130_n N_Y_M1001_d 0.00215158f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_99 N_VPWR_c_132_n Y 0.0161534f $X=0.38 $Y=2.085 $X2=0 $Y2=0
cc_100 N_VPWR_M1002_d N_Y_c_167_n 0.00909596f $X=1.135 $Y=1.835 $X2=0 $Y2=0
cc_101 N_VPWR_c_134_n N_Y_c_167_n 0.0218807f $X=1.33 $Y=2.4 $X2=0 $Y2=0
cc_102 N_VPWR_c_132_n N_Y_c_165_n 0.0730185f $X=0.38 $Y=2.085 $X2=0 $Y2=0
cc_103 N_VPWR_c_133_n N_Y_c_165_n 0.0209688f $X=1.165 $Y=3.33 $X2=0 $Y2=0
cc_104 N_VPWR_c_130_n N_Y_c_165_n 0.013415f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_105 N_VPWR_c_135_n N_Y_c_162_n 0.0441397f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_106 N_VPWR_c_130_n N_Y_c_162_n 0.0251927f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_107 N_Y_c_159_n N_VGND_c_195_n 0.0162156f $X=2.02 $Y=0.525 $X2=0 $Y2=0
cc_108 N_Y_c_159_n N_VGND_c_196_n 0.0138765f $X=2.02 $Y=0.525 $X2=0 $Y2=0
