* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__srsdfrtp_1 CLK D RESET_B SCD SCE SLEEP_B KAPWR VGND VNB VPB
+ VPWR Q
X0 a_220_136# SCE a_332_136# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1098_271# CLK a_3335_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_1128_424# a_1176_349# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_462_136# a_27_110# a_534_136# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_3063_390# RESET_B a_2176_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_929_152# a_1176_349# a_1343_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_3335_97# SLEEP_B a_3407_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR RESET_B a_999_424# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND RESET_B a_534_136# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_2069_397# a_1098_271# a_1176_349# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 a_1931_125# a_969_318# a_1982_397# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_2472_119# a_1982_397# a_2544_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR SCE a_313_466# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_332_136# a_27_110# a_552_466# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_332_136# a_969_318# a_999_424# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_332_136# D a_462_136# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_27_110# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 KAPWR CLK a_1098_271# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 VPWR a_1098_271# a_969_318# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_2176_99# a_1982_397# a_2472_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1176_349# a_999_424# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_3751_367# a_1982_397# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_3694_73# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_999_424# a_1098_271# a_1128_424# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_1343_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_1982_397# a_3751_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_929_152# a_969_318# a_999_424# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 KAPWR a_2586_249# a_3063_390# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X28 a_2544_119# a_2586_249# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1982_397# a_1098_271# a_2134_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_1982_397# a_969_318# a_2836_390# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X31 KAPWR SLEEP_B a_2586_249# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X32 a_552_466# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 a_1176_349# a_999_424# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X34 a_2206_125# a_2176_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_2836_390# a_2176_99# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X36 a_999_424# a_1098_271# a_332_136# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VGND a_1098_271# a_969_318# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_3407_97# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VGND a_3751_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X40 a_2586_249# SLEEP_B a_3694_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 VGND RESET_B a_2544_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_313_466# D a_332_136# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X43 a_2134_125# a_2176_99# a_2206_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_534_136# SCD a_220_136# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 a_2176_99# a_1982_397# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X46 VPWR a_3751_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X47 VPWR RESET_B a_332_136# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X48 a_1982_397# a_1098_271# a_2069_397# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X49 a_1176_349# a_969_318# a_1931_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X50 a_1098_271# SLEEP_B KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X51 a_27_110# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
