* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__srdlstp_1 D GATE SET_B SLEEP_B KAPWR VGND VNB VPB VPWR Q
X0 a_217_130# a_27_400# a_300_130# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_1294_315# SLEEP_B a_2144_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_700_451# a_404_353# a_844_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_667_47# a_434_405# a_700_451# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_988_47# a_1294_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_830_419# a_878_357# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_844_47# a_878_357# a_916_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_217_130# a_404_353# a_628_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 VGND SET_B a_988_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 KAPWR SLEEP_B a_1294_315# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_1455_127# a_700_451# a_878_357# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_700_451# SET_B a_1246_341# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_404_353# SLEEP_B KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_700_451# a_434_405# a_830_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 a_2144_131# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VPWR a_27_400# a_217_130# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 VGND a_700_451# a_1455_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_404_353# GATE a_1798_174# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1246_341# a_1294_315# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X19 a_217_130# a_434_405# a_667_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_1876_174# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_628_451# a_404_353# a_700_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 KAPWR a_700_451# a_878_357# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X23 a_2266_367# a_700_451# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 VGND a_700_451# a_2266_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_1798_174# SLEEP_B a_1876_174# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND D a_27_400# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VPWR a_404_353# a_434_405# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 VPWR a_2266_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_300_130# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 a_916_47# a_878_357# a_988_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 KAPWR GATE a_404_353# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 VGND a_2266_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 a_27_400# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X34 VGND a_404_353# a_434_405# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
