* File: sky130_fd_sc_lp__sdfbbp_1.spice
* Created: Wed Sep  2 10:33:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfbbp_1.pex.spice"
.subckt sky130_fd_sc_lp__sdfbbp_1  VNB VPB SCD D SCE CLK SET_B RESET_B VPWR Q_N
+ Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* CLK	CLK
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1033 A_126_119# N_SCD_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1013 N_A_204_119#_M1013_d N_SCE_M1013_g A_126_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1019 A_290_119# N_D_M1019_g N_A_204_119#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_332_93#_M1003_g A_290_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.0441 PD=0.97 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1034 N_A_332_93#_M1034_d N_SCE_M1034_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1155 PD=1.41 PS=0.97 NRD=0 NRS=77.136 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_A_755_106#_M1015_d N_CLK_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1764 AS=0.1764 PD=1.68 PS=1.68 NRD=38.568 NRS=38.568 M=1 R=2.8
+ SA=75000.3 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_755_106#_M1022_g N_A_893_101#_M1022_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.3123 AS=0.1197 PD=2.28 PS=1.41 NRD=78.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1004 N_A_1216_457#_M1004_d N_A_755_106#_M1004_g N_A_204_119#_M1004_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1023 A_1318_47# N_A_893_101#_M1023_g N_A_1216_457#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1297_290#_M1010_g A_1318_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0847528 AS=0.0441 PD=0.792453 PS=0.63 NRD=22.848 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1026 N_A_1492_47#_M1026_d N_SET_B_M1026_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.129147 PD=0.92 PS=1.20755 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_1297_290#_M1001_d N_A_1216_457#_M1001_g N_A_1492_47#_M1026_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1152 AS=0.0896 PD=1 PS=0.92 NRD=14.988 NRS=0 M=1
+ R=4.26667 SA=75001.5 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1007 N_A_1492_47#_M1007_d N_A_1650_21#_M1007_g N_A_1297_290#_M1001_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1824 AS=0.1152 PD=1.85 PS=1 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75002 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 A_1880_57# N_A_1297_290#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.1888 PD=0.91 PS=1.87 NRD=15 NRS=1.872 M=1 R=4.26667 SA=75000.2
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1018 N_A_1861_431#_M1018_d N_A_893_101#_M1018_g A_1880_57# VNB NSHORT L=0.15
+ W=0.64 AD=0.129147 AS=0.0864 PD=1.20755 PS=0.91 NRD=0 NRS=15 M=1 R=4.26667
+ SA=75000.6 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1027 A_2066_101# N_A_755_106#_M1027_g N_A_1861_431#_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75001.1 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_2064_453#_M1009_g A_2066_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.119185 AS=0.0504 PD=0.923208 PS=0.66 NRD=48.564 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 N_A_2279_57#_M1011_d N_SET_B_M1011_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.181615 PD=0.92 PS=1.40679 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75001.6 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1028 N_A_2064_453#_M1028_d N_A_1861_431#_M1028_g N_A_2279_57#_M1011_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.23975 AS=0.0896 PD=1.73 PS=0.92 NRD=59.916 NRS=0 M=1
+ R=4.26667 SA=75002 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1047 N_A_2279_57#_M1047_d N_A_1650_21#_M1047_g N_A_2064_453#_M1028_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1696 AS=0.23975 PD=1.81 PS=1.73 NRD=0 NRS=59.916 M=1
+ R=4.26667 SA=75002.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1002_d N_RESET_B_M1002_g N_A_1650_21#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1036 N_Q_N_M1036_d N_A_2064_453#_M1036_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1806 PD=2.25 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1039 N_VGND_M1039_d N_A_2064_453#_M1039_g N_A_2892_137#_M1039_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1030 N_Q_M1030_d N_A_2892_137#_M1030_g N_VGND_M1039_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1806 PD=2.25 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1037 N_VPWR_M1037_d N_SCD_M1037_g N_A_27_481#_M1037_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.128 AS=0.1824 PD=1.04 PS=1.85 NRD=24.6053 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1032 A_224_481# N_SCE_M1032_g N_VPWR_M1037_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.128 PD=0.88 PS=1.04 NRD=19.9955 NRS=12.2928 M=1 R=4.26667
+ SA=75000.8 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 N_A_204_119#_M1005_d N_D_M1005_g A_224_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1041 N_A_27_481#_M1041_d N_A_332_93#_M1041_g N_A_204_119#_M1005_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2336 AS=0.0896 PD=2.01 PS=0.92 NRD=24.6053 NRS=0 M=1
+ R=4.26667 SA=75001.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1038 N_A_332_93#_M1038_d N_SCE_M1038_g N_VPWR_M1038_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_755_106#_M1006_d N_CLK_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1042 N_VPWR_M1042_d N_A_755_106#_M1042_g N_A_893_101#_M1042_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2336 AS=0.1824 PD=2.01 PS=1.85 NRD=24.6053 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1012 N_A_1216_457#_M1012_d N_A_893_101#_M1012_g N_A_204_119#_M1012_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1043 A_1302_457# N_A_755_106#_M1043_g N_A_1216_457#_M1012_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75004 A=0.063 P=1.14 MULT=1
MM1016 N_VPWR_M1016_d N_A_1297_290#_M1016_g A_1302_457# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.14025 AS=0.0504 PD=1.04333 PS=0.66 NRD=130.828 NRS=30.4759 M=1
+ R=2.8 SA=75001 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1040 N_A_1297_290#_M1040_d N_SET_B_M1040_g N_VPWR_M1016_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1176 AS=0.2805 PD=1.12 PS=2.08667 NRD=0 NRS=65.404 M=1 R=5.6
+ SA=75001 SB=75002.3 A=0.126 P=1.98 MULT=1
MM1024 A_1584_373# N_A_1216_457#_M1024_g N_A_1297_290#_M1040_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1386 AS=0.1176 PD=1.17 PS=1.12 NRD=25.7873 NRS=0 M=1 R=5.6
+ SA=75001.4 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1046 N_VPWR_M1046_d N_A_1650_21#_M1046_g A_1584_373# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1176 AS=0.1386 PD=1.12 PS=1.17 NRD=0 NRS=25.7873 M=1 R=5.6 SA=75001.9
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1031 A_1766_373# N_A_1297_290#_M1031_g N_VPWR_M1046_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.161875 AS=0.1176 PD=1.455 PS=1.12 NRD=32.2883 NRS=0 M=1 R=5.6
+ SA=75002.3 SB=75001 A=0.126 P=1.98 MULT=1
MM1035 N_A_1861_431#_M1035_d N_A_755_106#_M1035_g A_1766_373# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1806 AS=0.161875 PD=1.6 PS=1.455 NRD=0 NRS=32.2883 M=1 R=5.6
+ SA=75002.1 SB=75001.8 A=0.126 P=1.98 MULT=1
MM1029 A_1963_515# N_A_893_101#_M1029_g N_A_1861_431#_M1035_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.10605 AS=0.0903 PD=0.925 PS=0.8 NRD=92.6294 NRS=37.5088 M=1 R=2.8
+ SA=75001.7 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_A_2064_453#_M1017_g A_1963_515# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1582 AS=0.10605 PD=1.12333 PS=0.925 NRD=265.004 NRS=92.6294 M=1
+ R=2.8 SA=75002.3 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1020 N_A_2064_453#_M1020_d N_SET_B_M1020_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1512 AS=0.3164 PD=1.2 PS=2.24667 NRD=18.7544 NRS=0 M=1 R=5.6
+ SA=75001.8 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1021 A_2395_451# N_A_1861_431#_M1021_g N_A_2064_453#_M1020_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1134 AS=0.1512 PD=1.11 PS=1.2 NRD=18.7544 NRS=0 M=1 R=5.6
+ SA=75002.3 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1014 N_VPWR_M1014_d N_A_1650_21#_M1014_g A_2395_451# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2394 AS=0.1134 PD=2.25 PS=1.11 NRD=0 NRS=18.7544 M=1 R=5.6 SA=75002.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_RESET_B_M1000_g N_A_1650_21#_M1000_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.137128 AS=0.1824 PD=1.09137 PS=1.85 NRD=49.0136 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1045 N_Q_N_M1045_d N_A_2064_453#_M1045_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.269972 PD=3.09 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1025_d N_A_2064_453#_M1025_g N_A_2892_137#_M1025_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.137128 AS=0.1824 PD=1.09137 PS=1.85 NRD=25.3933 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1044 N_Q_M1044_d N_A_2892_137#_M1044_g N_VPWR_M1025_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.269972 PD=3.09 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX48_noxref VNB VPB NWDIODE A=29.8059 P=37.11
c_194 VNB 0 3.33237e-19 $X=0 $Y=0
c_2198 A_224_481# 0 2.49076e-20 $X=1.12 $Y=2.405
*
.include "sky130_fd_sc_lp__sdfbbp_1.pxi.spice"
*
.ends
*
*
