* NGSPICE file created from sky130_fd_sc_lp__a2bb2o_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2bb2o_lp A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_742_74# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.549e+11p ps=4.21e+06u
M1001 a_900_74# A2_N a_284_31# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1002 a_43_408# B1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.9e+11p pd=5.18e+06u as=7.2e+11p ps=5.44e+06u
M1003 VPWR a_63_57# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1004 VGND A2_N a_900_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_63_57# a_284_31# a_43_408# VPB phighvt w=1e+06u l=250000u
+  ad=5.9e+11p pd=3.18e+06u as=0p ps=0u
M1006 a_794_409# A1_N VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1007 VGND B1 a_150_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 VPWR B2 a_43_408# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_150_57# B2 a_63_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.82e+06u
M1010 a_584_74# a_63_57# X VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1011 VGND a_63_57# a_584_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_314_57# a_284_31# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1013 a_284_31# A1_N a_742_74# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_63_57# a_284_31# a_314_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_284_31# A2_N a_794_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends

