* File: sky130_fd_sc_lp__a41o_1.spice
* Created: Wed Sep  2 09:28:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41o_1.pex.spice"
.subckt sky130_fd_sc_lp__a41o_1  VNB VPB B1 A1 A2 A3 A4 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_113_237#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.3255 AS=0.2226 PD=1.615 PS=2.21 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1010 N_A_113_237#_M1010_d N_B1_M1010_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2352 AS=0.3255 PD=1.4 PS=1.615 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1002 A_478_47# N_A1_M1002_g N_A_113_237#_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2352 PD=1.05 PS=1.4 NRD=7.14 NRS=39.996 M=1 R=5.6 SA=75001.8
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1000 A_550_47# N_A2_M1000_g A_478_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75002.2 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1004 A_658_47# N_A3_M1004_g A_550_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.1638 PD=1.23 PS=1.23 NRD=19.992 NRS=19.992 M=1 R=5.6 SA=75002.7
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A4_M1007_g A_658_47# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6 SA=75003.3 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A_113_237#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1011 N_A_346_367#_M1011_d N_B1_M1011_g N_A_113_237#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_346_367#_M1011_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3906 AS=0.1764 PD=1.88 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_A_346_367#_M1003_d N_A2_M1003_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3906 PD=1.54 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75001.4
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A3_M1009_g N_A_346_367#_M1003_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75001.8 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1006 N_A_346_367#_M1006_d N_A4_M1006_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2016 PD=3.05 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75002.3 SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__a41o_1.pxi.spice"
*
.ends
*
*
