* File: sky130_fd_sc_lp__or4bb_1.spice
* Created: Fri Aug 28 11:26:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4bb_1.pex.spice"
.subckt sky130_fd_sc_lp__or4bb_1  VNB VPB C_N D_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C_N_M1008_g N_A_27_535#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_196_535#_M1009_d N_D_N_M1009_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_332_391#_M1010_d N_A_196_535#_M1010_g N_VGND_M1010_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_27_535#_M1004_g N_A_332_391#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1013 N_A_332_391#_M1013_d N_B_M1013_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001.1
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_332_391#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.098 AS=0.0588 PD=0.85 PS=0.7 NRD=34.284 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1012 N_X_M1012_d N_A_332_391#_M1012_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.196 PD=2.21 PS=1.7 NRD=0 NRS=2.496 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_VPWR_M1011_d N_C_N_M1011_g N_A_27_535#_M1011_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_196_535#_M1003_d N_D_N_M1003_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_415_391# N_A_196_535#_M1000_g N_A_332_391#_M1000_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1002 A_487_391# N_A_27_535#_M1002_g A_415_391# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=65.6601 NRS=23.443 M=1 R=2.8
+ SA=75000.6 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1005 A_595_391# N_B_M1005_g A_487_391# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=65.6601 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_595_391# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0441 PD=0.8175 PS=0.63 NRD=46.886 NRS=23.443 M=1 R=2.8
+ SA=75001.4 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_332_391#_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__or4bb_1.pxi.spice"
*
.ends
*
*
