* File: sky130_fd_sc_lp__nor2_0.spice
* Created: Wed Sep  2 10:07:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor2_0.pex.spice"
.subckt sky130_fd_sc_lp__nor2_0  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_B_M1000_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1001 A_120_483# N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.1696 PD=0.88 PS=1.81 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g A_120_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.1696
+ AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
c_96 A_120_483# 0 1.06273e-19 $X=0.6 $Y=2.415
*
.include "sky130_fd_sc_lp__nor2_0.pxi.spice"
*
.ends
*
*
