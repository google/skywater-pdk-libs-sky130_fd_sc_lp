* File: sky130_fd_sc_lp__and4_2.spice
* Created: Fri Aug 28 10:07:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4_2.pex.spice"
.subckt sky130_fd_sc_lp__and4_2  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1010 A_155_49# N_A_M1010_g N_A_72_49#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1007 A_227_49# N_B_M1007_g A_155_49# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1001 A_335_49# N_C_M1001_g A_227_49# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=39.996 M=1 R=2.8 SA=75001.1
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_D_M1006_g A_335_49# VNB NSHORT L=0.15 W=0.42 AD=0.1232
+ AS=0.0819 PD=0.97 PS=0.81 NRD=48.564 NRS=39.996 M=1 R=2.8 SA=75001.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_72_49#_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2464 PD=1.12 PS=1.94 NRD=0 NRS=23.568 M=1 R=5.6 SA=75001.3
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1002_d N_A_72_49#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_A_72_49#_M1009_d N_A_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.8
+ A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_A_72_49#_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.105 AS=0.0588 PD=0.92 PS=0.7 NRD=46.886 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1005 N_A_72_49#_M1005_d N_C_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.105 PD=0.7 PS=0.92 NRD=0 NRS=56.2829 M=1 R=2.8 SA=75001.3
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_72_49#_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.112875 AS=0.0588 PD=0.9025 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_72_49#_M1004_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.338625 PD=1.54 PS=2.7075 NRD=0 NRS=13.8097 M=1 R=8.4 SA=75000.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1011 N_X_M1004_d N_A_72_49#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_66 VPB 0 1.0248e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__and4_2.pxi.spice"
*
.ends
*
*
