* File: sky130_fd_sc_lp__o41ai_4.pxi.spice
* Created: Fri Aug 28 11:20:35 2020
* 
x_PM_SKY130_FD_SC_LP__O41AI_4%B1 N_B1_M1004_g N_B1_M1010_g N_B1_M1006_g
+ N_B1_M1014_g N_B1_M1018_g N_B1_M1026_g N_B1_M1033_g N_B1_M1029_g B1 B1 B1 B1
+ B1 B1 N_B1_c_171_n N_B1_c_172_n N_B1_c_173_n PM_SKY130_FD_SC_LP__O41AI_4%B1
x_PM_SKY130_FD_SC_LP__O41AI_4%A4 N_A4_c_253_n N_A4_M1007_g N_A4_M1013_g
+ N_A4_M1021_g N_A4_c_256_n N_A4_M1008_g N_A4_M1024_g N_A4_c_258_n N_A4_M1037_g
+ N_A4_M1035_g N_A4_c_260_n N_A4_M1038_g N_A4_c_300_p A4 A4 N_A4_c_261_n
+ N_A4_c_262_n N_A4_c_263_n PM_SKY130_FD_SC_LP__O41AI_4%A4
x_PM_SKY130_FD_SC_LP__O41AI_4%A3 N_A3_c_356_n N_A3_M1002_g N_A3_M1015_g
+ N_A3_c_357_n N_A3_M1016_g N_A3_M1030_g N_A3_c_358_n N_A3_M1022_g N_A3_M1034_g
+ N_A3_c_359_n N_A3_M1027_g N_A3_M1039_g A3 A3 A3 A3 N_A3_c_355_n
+ PM_SKY130_FD_SC_LP__O41AI_4%A3
x_PM_SKY130_FD_SC_LP__O41AI_4%A2 N_A2_M1009_g N_A2_M1000_g N_A2_M1012_g
+ N_A2_M1011_g N_A2_M1028_g N_A2_M1020_g N_A2_M1032_g N_A2_M1025_g N_A2_c_458_n
+ A2 N_A2_c_459_n N_A2_c_460_n PM_SKY130_FD_SC_LP__O41AI_4%A2
x_PM_SKY130_FD_SC_LP__O41AI_4%A1 N_A1_c_551_n N_A1_M1001_g N_A1_M1005_g
+ N_A1_c_553_n N_A1_M1003_g N_A1_M1017_g N_A1_c_555_n N_A1_M1019_g N_A1_M1023_g
+ N_A1_c_557_n N_A1_M1031_g N_A1_M1036_g A1 A1 N_A1_c_560_n
+ PM_SKY130_FD_SC_LP__O41AI_4%A1
x_PM_SKY130_FD_SC_LP__O41AI_4%VPWR N_VPWR_M1004_d N_VPWR_M1006_d N_VPWR_M1033_d
+ N_VPWR_M1005_d N_VPWR_M1023_d N_VPWR_c_621_n N_VPWR_c_622_n N_VPWR_c_623_n
+ N_VPWR_c_624_n N_VPWR_c_625_n N_VPWR_c_626_n N_VPWR_c_627_n N_VPWR_c_628_n
+ N_VPWR_c_629_n VPWR N_VPWR_c_630_n N_VPWR_c_631_n N_VPWR_c_632_n
+ N_VPWR_c_633_n N_VPWR_c_620_n N_VPWR_c_635_n N_VPWR_c_636_n N_VPWR_c_637_n
+ PM_SKY130_FD_SC_LP__O41AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O41AI_4%Y N_Y_M1010_d N_Y_M1026_d N_Y_M1004_s N_Y_M1018_s
+ N_Y_M1013_d N_Y_M1024_d N_Y_c_757_n N_Y_c_819_n N_Y_c_759_n N_Y_c_842_p
+ N_Y_c_749_n N_Y_c_750_n N_Y_c_823_n N_Y_c_754_n N_Y_c_846_p N_Y_c_751_n
+ N_Y_c_788_n N_Y_c_793_n N_Y_c_776_n N_Y_c_752_n N_Y_c_796_n Y Y N_Y_c_756_n Y
+ PM_SKY130_FD_SC_LP__O41AI_4%Y
x_PM_SKY130_FD_SC_LP__O41AI_4%A_554_361# N_A_554_361#_M1013_s
+ N_A_554_361#_M1021_s N_A_554_361#_M1035_s N_A_554_361#_M1016_d
+ N_A_554_361#_M1027_d N_A_554_361#_c_858_n N_A_554_361#_c_859_n
+ N_A_554_361#_c_860_n N_A_554_361#_c_903_n N_A_554_361#_c_861_n
+ N_A_554_361#_c_862_n N_A_554_361#_c_872_n N_A_554_361#_c_871_n
+ N_A_554_361#_c_914_p N_A_554_361#_c_877_n N_A_554_361#_c_863_n
+ N_A_554_361#_c_864_n N_A_554_361#_c_865_n N_A_554_361#_c_883_n
+ PM_SKY130_FD_SC_LP__O41AI_4%A_554_361#
x_PM_SKY130_FD_SC_LP__O41AI_4%A_981_361# N_A_981_361#_M1002_s
+ N_A_981_361#_M1022_s N_A_981_361#_M1000_s N_A_981_361#_M1020_s
+ N_A_981_361#_c_928_n N_A_981_361#_c_924_n N_A_981_361#_c_925_n
+ N_A_981_361#_c_935_n N_A_981_361#_c_926_n N_A_981_361#_c_942_n
+ N_A_981_361#_c_945_n N_A_981_361#_c_947_n N_A_981_361#_c_948_n
+ N_A_981_361#_c_927_n N_A_981_361#_c_949_n
+ PM_SKY130_FD_SC_LP__O41AI_4%A_981_361#
x_PM_SKY130_FD_SC_LP__O41AI_4%A_1346_367# N_A_1346_367#_M1000_d
+ N_A_1346_367#_M1011_d N_A_1346_367#_M1025_d N_A_1346_367#_M1017_s
+ N_A_1346_367#_M1036_s N_A_1346_367#_c_990_n N_A_1346_367#_c_991_n
+ N_A_1346_367#_c_1002_n N_A_1346_367#_c_1007_n N_A_1346_367#_c_992_n
+ N_A_1346_367#_c_1034_n N_A_1346_367#_c_993_n N_A_1346_367#_c_1038_n
+ N_A_1346_367#_c_994_n N_A_1346_367#_c_995_n N_A_1346_367#_c_996_n
+ N_A_1346_367#_c_997_n N_A_1346_367#_c_998_n
+ PM_SKY130_FD_SC_LP__O41AI_4%A_1346_367#
x_PM_SKY130_FD_SC_LP__O41AI_4%A_192_47# N_A_192_47#_M1010_s N_A_192_47#_M1014_s
+ N_A_192_47#_M1029_s N_A_192_47#_M1008_d N_A_192_47#_M1038_d
+ N_A_192_47#_M1030_s N_A_192_47#_M1039_s N_A_192_47#_M1012_s
+ N_A_192_47#_M1032_s N_A_192_47#_M1003_d N_A_192_47#_M1031_d
+ N_A_192_47#_c_1060_n N_A_192_47#_c_1076_n N_A_192_47#_c_1061_n
+ N_A_192_47#_c_1078_n N_A_192_47#_c_1080_n N_A_192_47#_c_1081_n
+ N_A_192_47#_c_1088_n N_A_192_47#_c_1083_n N_A_192_47#_c_1090_n
+ N_A_192_47#_c_1094_n N_A_192_47#_c_1100_n N_A_192_47#_c_1096_n
+ N_A_192_47#_c_1062_n N_A_192_47#_c_1063_n N_A_192_47#_c_1199_p
+ N_A_192_47#_c_1064_n N_A_192_47#_c_1182_p N_A_192_47#_c_1065_n
+ N_A_192_47#_c_1123_n N_A_192_47#_c_1066_n N_A_192_47#_c_1129_n
+ N_A_192_47#_c_1138_n N_A_192_47#_c_1201_p N_A_192_47#_c_1067_n
+ N_A_192_47#_c_1068_n N_A_192_47#_c_1084_n N_A_192_47#_c_1098_n
+ N_A_192_47#_c_1114_n N_A_192_47#_c_1069_n N_A_192_47#_c_1070_n
+ N_A_192_47#_c_1071_n N_A_192_47#_c_1072_n N_A_192_47#_c_1147_n
+ PM_SKY130_FD_SC_LP__O41AI_4%A_192_47#
x_PM_SKY130_FD_SC_LP__O41AI_4%VGND N_VGND_M1007_s N_VGND_M1037_s N_VGND_M1015_d
+ N_VGND_M1034_d N_VGND_M1009_d N_VGND_M1028_d N_VGND_M1001_s N_VGND_M1019_s
+ N_VGND_c_1229_n N_VGND_c_1230_n N_VGND_c_1231_n N_VGND_c_1232_n
+ N_VGND_c_1233_n N_VGND_c_1234_n N_VGND_c_1235_n N_VGND_c_1236_n
+ N_VGND_c_1237_n N_VGND_c_1238_n N_VGND_c_1239_n N_VGND_c_1240_n
+ N_VGND_c_1241_n N_VGND_c_1242_n N_VGND_c_1243_n N_VGND_c_1244_n
+ N_VGND_c_1245_n N_VGND_c_1246_n VGND N_VGND_c_1247_n N_VGND_c_1248_n
+ N_VGND_c_1249_n N_VGND_c_1250_n N_VGND_c_1251_n N_VGND_c_1252_n
+ N_VGND_c_1253_n N_VGND_c_1254_n PM_SKY130_FD_SC_LP__O41AI_4%VGND
cc_1 VNB N_B1_M1004_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.465
cc_2 VNB N_B1_M1010_g 0.0303789f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.655
cc_3 VNB N_B1_M1006_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.465
cc_4 VNB N_B1_M1014_g 0.0208457f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=0.655
cc_5 VNB N_B1_M1018_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.465
cc_6 VNB N_B1_M1026_g 0.0208457f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=0.655
cc_7 VNB N_B1_M1033_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=2.465
cc_8 VNB N_B1_M1029_g 0.0221179f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.655
cc_9 VNB N_B1_c_171_n 0.0905758f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.46
cc_10 VNB N_B1_c_172_n 0.119106f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.46
cc_11 VNB N_B1_c_173_n 0.0136787f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.46
cc_12 VNB N_A4_c_253_n 0.0165325f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.625
cc_13 VNB N_A4_M1013_g 7.5798e-19 $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.655
cc_14 VNB N_A4_M1021_g 8.07393e-19 $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.465
cc_15 VNB N_A4_c_256_n 0.0159768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A4_M1024_g 9.60681e-19 $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.625
cc_17 VNB N_A4_c_258_n 0.0160583f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.465
cc_18 VNB N_A4_M1035_g 8.87946e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A4_c_260_n 0.016586f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=2.465
cc_20 VNB N_A4_c_261_n 0.104348f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_21 VNB N_A4_c_262_n 0.00212684f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.46
cc_22 VNB N_A4_c_263_n 2.34925e-19 $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.46
cc_23 VNB N_A3_M1015_g 0.0242964f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.655
cc_24 VNB N_A3_M1030_g 0.0228993f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.295
cc_25 VNB N_A3_M1034_g 0.0217473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A3_M1039_g 0.0219843f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=2.465
cc_27 VNB A3 0.00346044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A3_c_355_n 0.0827594f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_29 VNB N_A2_M1009_g 0.0199433f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.465
cc_30 VNB N_A2_M1000_g 0.00237454f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.655
cc_31 VNB N_A2_M1012_g 0.0197131f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.465
cc_32 VNB N_A2_M1011_g 0.00247727f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=0.655
cc_33 VNB N_A2_M1028_g 0.0215227f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=2.465
cc_34 VNB N_A2_M1020_g 0.0024903f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=0.655
cc_35 VNB N_A2_M1032_g 0.0218108f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=2.465
cc_36 VNB N_A2_M1025_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.655
cc_37 VNB N_A2_c_458_n 0.00140263f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_38 VNB N_A2_c_459_n 0.0965304f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.46
cc_39 VNB N_A2_c_460_n 0.00246341f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.46
cc_40 VNB N_A1_c_551_n 0.0164412f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.625
cc_41 VNB N_A1_M1005_g 0.0072706f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.655
cc_42 VNB N_A1_c_553_n 0.0162013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A1_M1017_g 0.00700214f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.295
cc_44 VNB N_A1_c_555_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=0.655
cc_45 VNB N_A1_M1023_g 0.00700214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A1_c_557_n 0.0218799f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=0.655
cc_47 VNB N_A1_M1036_g 0.0110049f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=2.465
cc_48 VNB A1 0.0246677f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.655
cc_49 VNB N_A1_c_560_n 0.116685f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_50 VNB N_VPWR_c_620_n 0.442315f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.567
cc_51 VNB N_Y_c_749_n 0.00316451f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=1.295
cc_52 VNB N_Y_c_750_n 0.00325523f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.655
cc_53 VNB N_Y_c_751_n 0.0157768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_Y_c_752_n 0.00147586f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.46
cc_55 VNB Y 0.00347744f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.46
cc_56 VNB N_A_192_47#_c_1060_n 0.0280113f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_57 VNB N_A_192_47#_c_1061_n 0.00746637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_192_47#_c_1062_n 0.00312562f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.46
cc_59 VNB N_A_192_47#_c_1063_n 0.00147353f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.46
cc_60 VNB N_A_192_47#_c_1064_n 0.00295761f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.46
cc_61 VNB N_A_192_47#_c_1065_n 0.00287687f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.567
cc_62 VNB N_A_192_47#_c_1066_n 0.00320439f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.567
cc_63 VNB N_A_192_47#_c_1067_n 0.00740486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_192_47#_c_1068_n 0.0235964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_192_47#_c_1069_n 0.00145145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_192_47#_c_1070_n 0.00695479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_192_47#_c_1071_n 0.00186571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_192_47#_c_1072_n 0.00380767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1229_n 0.002833f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=2.465
cc_70 VNB N_VGND_c_1230_n 0.00288811f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=0.655
cc_71 VNB N_VGND_c_1231_n 0.00272739f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_72 VNB N_VGND_c_1232_n 3.10008e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1233_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1234_n 3.20903e-19 $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.46
cc_75 VNB N_VGND_c_1235_n 0.0154314f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.46
cc_76 VNB N_VGND_c_1236_n 0.00434038f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.46
cc_77 VNB N_VGND_c_1237_n 0.00410954f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.46
cc_78 VNB N_VGND_c_1238_n 0.00204381f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.46
cc_79 VNB N_VGND_c_1239_n 0.080764f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.46
cc_80 VNB N_VGND_c_1240_n 0.00510363f $X=-0.19 $Y=-0.245 $X2=2.59 $Y2=1.46
cc_81 VNB N_VGND_c_1241_n 0.0170844f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.46
cc_82 VNB N_VGND_c_1242_n 0.00516281f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.46
cc_83 VNB N_VGND_c_1243_n 0.0166818f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.567
cc_84 VNB N_VGND_c_1244_n 0.00516057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1245_n 0.0130989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1246_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.567
cc_87 VNB N_VGND_c_1247_n 0.0170402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1248_n 0.0162758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1249_n 0.0182108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1250_n 0.525441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1251_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1252_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1253_n 0.00528956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1254_n 0.00429093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VPB N_B1_M1004_g 0.0245754f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=2.465
cc_96 VPB N_B1_M1006_g 0.0187475f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.465
cc_97 VPB N_B1_M1018_g 0.0187475f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.465
cc_98 VPB N_B1_M1033_g 0.0245754f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=2.465
cc_99 VPB N_B1_c_172_n 0.00642874f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=1.46
cc_100 VPB N_B1_c_173_n 0.0378364f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=1.46
cc_101 VPB N_A4_M1013_g 0.0246398f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=0.655
cc_102 VPB N_A4_M1021_g 0.0187364f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.465
cc_103 VPB N_A4_M1024_g 0.0193914f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.625
cc_104 VPB N_A4_M1035_g 0.0187098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A4_c_262_n 0.00432863f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.46
cc_106 VPB N_A4_c_263_n 0.00201984f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=1.46
cc_107 VPB N_A3_c_356_n 0.0163121f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.625
cc_108 VPB N_A3_c_357_n 0.0158001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A3_c_358_n 0.0158022f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=0.655
cc_110 VPB N_A3_c_359_n 0.0209633f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=0.655
cc_111 VPB A3 0.0144031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A3_c_355_n 0.0341576f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_113 VPB N_A2_M1000_g 0.0252886f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=0.655
cc_114 VPB N_A2_M1011_g 0.0197262f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=0.655
cc_115 VPB N_A2_M1020_g 0.0186059f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=0.655
cc_116 VPB N_A2_M1025_g 0.0187442f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=0.655
cc_117 VPB N_A2_c_460_n 0.00555451f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.46
cc_118 VPB N_A1_M1005_g 0.0185451f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=0.655
cc_119 VPB N_A1_M1017_g 0.0184123f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.295
cc_120 VPB N_A1_M1023_g 0.0184123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A1_M1036_g 0.0243928f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=2.465
cc_122 VPB N_VPWR_c_621_n 0.0478673f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.465
cc_123 VPB N_VPWR_c_622_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_623_n 0.010528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_624_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_625_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.58
cc_127 VPB N_VPWR_c_626_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_627_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_628_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_130 VPB N_VPWR_c_629_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_131 VPB N_VPWR_c_630_n 0.0177361f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.46
cc_132 VPB N_VPWR_c_631_n 0.145154f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.46
cc_133 VPB N_VPWR_c_632_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=1.46
cc_134 VPB N_VPWR_c_633_n 0.015535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_620_n 0.0915257f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.567
cc_136 VPB N_VPWR_c_635_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=1.567
cc_137 VPB N_VPWR_c_636_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.97 $Y2=1.567
cc_138 VPB N_VPWR_c_637_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=1.567
cc_139 VPB N_Y_c_754_n 0.0107298f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_140 VPB Y 4.91169e-19 $X=-0.19 $Y=1.655 $X2=1.97 $Y2=1.46
cc_141 VPB N_Y_c_756_n 0.00346786f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=1.46
cc_142 VPB N_A_554_361#_c_858_n 0.0058574f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.465
cc_143 VPB N_A_554_361#_c_859_n 0.00262279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_554_361#_c_860_n 0.00355243f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.295
cc_145 VPB N_A_554_361#_c_861_n 0.00262279f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=2.465
cc_146 VPB N_A_554_361#_c_862_n 0.00145278f $X=-0.19 $Y=1.655 $X2=2.59 $Y2=1.295
cc_147 VPB N_A_554_361#_c_863_n 0.00299384f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.58
cc_148 VPB N_A_554_361#_c_864_n 0.00441432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_554_361#_c_865_n 0.00138314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_981_361#_c_924_n 0.00200254f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.625
cc_151 VPB N_A_981_361#_c_925_n 0.00203831f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=2.465
cc_152 VPB N_A_981_361#_c_926_n 0.0135584f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=0.655
cc_153 VPB N_A_981_361#_c_927_n 0.00203831f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_154 VPB N_A_1346_367#_c_990_n 0.00324748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_1346_367#_c_991_n 0.00551768f $X=-0.19 $Y=1.655 $X2=1.73
+ $Y2=2.465
cc_156 VPB N_A_1346_367#_c_992_n 0.00288963f $X=-0.19 $Y=1.655 $X2=2.16
+ $Y2=2.465
cc_157 VPB N_A_1346_367#_c_993_n 0.00309865f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.58
cc_158 VPB N_A_1346_367#_c_994_n 0.0125869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_1346_367#_c_995_n 0.0454116f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.46
cc_160 VPB N_A_1346_367#_c_996_n 0.0031124f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.46
cc_161 VPB N_A_1346_367#_c_997_n 0.0028792f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=1.46
cc_162 VPB N_A_1346_367#_c_998_n 0.00146192f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.46
cc_163 N_B1_M1029_g N_A4_c_253_n 0.0276984f $X=2.59 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_164 N_B1_c_172_n N_A4_M1013_g 0.00119454f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_165 N_B1_c_173_n N_A4_M1013_g 9.61013e-19 $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_166 N_B1_c_172_n N_A4_c_261_n 0.0214095f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_167 N_B1_c_173_n N_A4_c_261_n 2.58749e-19 $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_168 N_B1_c_172_n N_A4_c_262_n 0.0014926f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_169 N_B1_c_173_n N_A4_c_262_n 0.0348009f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_170 N_B1_M1004_g N_VPWR_c_621_n 0.0200737f $X=0.87 $Y=2.465 $X2=0 $Y2=0
cc_171 N_B1_M1006_g N_VPWR_c_621_n 7.26038e-19 $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_172 N_B1_c_171_n N_VPWR_c_621_n 0.00159857f $X=0.795 $Y=1.46 $X2=0 $Y2=0
cc_173 N_B1_c_173_n N_VPWR_c_621_n 0.0260594f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_174 N_B1_M1004_g N_VPWR_c_622_n 6.77662e-19 $X=0.87 $Y=2.465 $X2=0 $Y2=0
cc_175 N_B1_M1006_g N_VPWR_c_622_n 0.0144369f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_176 N_B1_M1018_g N_VPWR_c_622_n 0.0146218f $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_177 N_B1_M1033_g N_VPWR_c_622_n 6.90148e-19 $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_178 N_B1_M1018_g N_VPWR_c_623_n 6.77662e-19 $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_179 N_B1_M1033_g N_VPWR_c_623_n 0.0168606f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_180 N_B1_M1004_g N_VPWR_c_626_n 0.00486043f $X=0.87 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B1_M1006_g N_VPWR_c_626_n 0.00486043f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B1_M1018_g N_VPWR_c_628_n 0.00486043f $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B1_M1033_g N_VPWR_c_628_n 0.00486043f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_184 N_B1_M1004_g N_VPWR_c_620_n 0.00824727f $X=0.87 $Y=2.465 $X2=0 $Y2=0
cc_185 N_B1_M1006_g N_VPWR_c_620_n 0.00824727f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B1_M1018_g N_VPWR_c_620_n 0.00824727f $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_187 N_B1_M1033_g N_VPWR_c_620_n 0.00824727f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_188 N_B1_c_172_n N_Y_c_757_n 5.70981e-19 $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_189 N_B1_c_173_n N_Y_c_757_n 0.0155814f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_190 N_B1_M1006_g N_Y_c_759_n 0.0122595f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B1_M1018_g N_Y_c_759_n 0.0122129f $X=1.73 $Y=2.465 $X2=0 $Y2=0
cc_192 N_B1_c_172_n N_Y_c_759_n 5.04482e-19 $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_193 N_B1_c_173_n N_Y_c_759_n 0.0438476f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_194 N_B1_M1014_g N_Y_c_749_n 0.0119277f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_195 N_B1_M1026_g N_Y_c_749_n 0.012224f $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_196 N_B1_c_172_n N_Y_c_749_n 0.00243312f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_197 N_B1_c_173_n N_Y_c_749_n 0.0456563f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_198 N_B1_M1010_g N_Y_c_750_n 0.00346282f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_199 N_B1_c_172_n N_Y_c_750_n 0.00252548f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_200 N_B1_c_173_n N_Y_c_750_n 0.0174368f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_201 N_B1_M1033_g N_Y_c_754_n 0.0143f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B1_c_172_n N_Y_c_754_n 0.00280821f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_203 N_B1_c_173_n N_Y_c_754_n 0.0568f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_204 N_B1_M1029_g N_Y_c_751_n 0.0126655f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_205 N_B1_c_172_n N_Y_c_751_n 0.00364968f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_206 N_B1_c_173_n N_Y_c_751_n 0.0235251f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_207 N_B1_c_172_n N_Y_c_776_n 5.70981e-19 $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_208 N_B1_c_173_n N_Y_c_776_n 0.0151534f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_209 N_B1_c_172_n N_Y_c_752_n 0.00252548f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_210 N_B1_c_173_n N_Y_c_752_n 0.0147242f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_211 N_B1_M1033_g N_A_554_361#_c_858_n 0.00130567f $X=2.16 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_B1_M1010_g N_A_192_47#_c_1060_n 0.00248138f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_213 N_B1_c_172_n N_A_192_47#_c_1060_n 0.00780822f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_214 N_B1_c_173_n N_A_192_47#_c_1060_n 0.0172135f $X=2.65 $Y=1.46 $X2=0 $Y2=0
cc_215 N_B1_M1010_g N_A_192_47#_c_1076_n 0.012237f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_216 N_B1_M1014_g N_A_192_47#_c_1076_n 0.0083908f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_217 N_B1_M1026_g N_A_192_47#_c_1078_n 0.0083908f $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_218 N_B1_M1029_g N_A_192_47#_c_1078_n 0.0083908f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_219 N_B1_M1029_g N_A_192_47#_c_1080_n 5.89773e-19 $X=2.59 $Y=0.655 $X2=0
+ $Y2=0
cc_220 N_B1_M1026_g N_A_192_47#_c_1081_n 4.572e-19 $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_221 N_B1_M1029_g N_A_192_47#_c_1081_n 0.00374699f $X=2.59 $Y=0.655 $X2=0
+ $Y2=0
cc_222 N_B1_M1029_g N_A_192_47#_c_1083_n 0.00207134f $X=2.59 $Y=0.655 $X2=0
+ $Y2=0
cc_223 N_B1_M1010_g N_A_192_47#_c_1084_n 5.12807e-19 $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_224 N_B1_M1014_g N_A_192_47#_c_1084_n 0.00648278f $X=1.73 $Y=0.655 $X2=0
+ $Y2=0
cc_225 N_B1_M1026_g N_A_192_47#_c_1084_n 0.00638749f $X=2.16 $Y=0.655 $X2=0
+ $Y2=0
cc_226 N_B1_M1029_g N_A_192_47#_c_1084_n 5.05577e-19 $X=2.59 $Y=0.655 $X2=0
+ $Y2=0
cc_227 N_B1_M1029_g N_VGND_c_1229_n 9.77997e-19 $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_228 N_B1_M1010_g N_VGND_c_1239_n 0.00357877f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_229 N_B1_M1014_g N_VGND_c_1239_n 0.00357842f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_230 N_B1_M1026_g N_VGND_c_1239_n 0.00357842f $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_231 N_B1_M1029_g N_VGND_c_1239_n 0.00357842f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_232 N_B1_M1010_g N_VGND_c_1250_n 0.00681251f $X=1.3 $Y=0.655 $X2=0 $Y2=0
cc_233 N_B1_M1014_g N_VGND_c_1250_n 0.00535118f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_234 N_B1_M1026_g N_VGND_c_1250_n 0.00535118f $X=2.16 $Y=0.655 $X2=0 $Y2=0
cc_235 N_B1_M1029_g N_VGND_c_1250_n 0.00555736f $X=2.59 $Y=0.655 $X2=0 $Y2=0
cc_236 N_A4_M1035_g N_A3_c_356_n 0.0131056f $X=4.4 $Y=2.435 $X2=-0.19 $Y2=-0.245
cc_237 N_A4_c_260_n N_A3_M1015_g 0.0267347f $X=4.56 $Y=1.185 $X2=0 $Y2=0
cc_238 N_A4_c_261_n A3 3.47954e-19 $X=4.4 $Y=1.395 $X2=0 $Y2=0
cc_239 N_A4_c_261_n N_A3_c_355_n 0.0210491f $X=4.4 $Y=1.395 $X2=0 $Y2=0
cc_240 N_A4_M1013_g N_VPWR_c_623_n 0.00232792f $X=3.11 $Y=2.435 $X2=0 $Y2=0
cc_241 N_A4_M1013_g N_VPWR_c_631_n 0.00338313f $X=3.11 $Y=2.435 $X2=0 $Y2=0
cc_242 N_A4_M1021_g N_VPWR_c_631_n 0.00338313f $X=3.54 $Y=2.435 $X2=0 $Y2=0
cc_243 N_A4_M1024_g N_VPWR_c_631_n 0.00338313f $X=3.97 $Y=2.435 $X2=0 $Y2=0
cc_244 N_A4_M1035_g N_VPWR_c_631_n 0.00338313f $X=4.4 $Y=2.435 $X2=0 $Y2=0
cc_245 N_A4_M1013_g N_VPWR_c_620_n 0.00619097f $X=3.11 $Y=2.435 $X2=0 $Y2=0
cc_246 N_A4_M1021_g N_VPWR_c_620_n 0.00509124f $X=3.54 $Y=2.435 $X2=0 $Y2=0
cc_247 N_A4_M1024_g N_VPWR_c_620_n 0.00509124f $X=3.97 $Y=2.435 $X2=0 $Y2=0
cc_248 N_A4_M1035_g N_VPWR_c_620_n 0.00511267f $X=4.4 $Y=2.435 $X2=0 $Y2=0
cc_249 N_A4_M1013_g N_Y_c_754_n 0.0131906f $X=3.11 $Y=2.435 $X2=0 $Y2=0
cc_250 N_A4_c_262_n N_Y_c_754_n 0.0111892f $X=3.483 $Y=1.557 $X2=0 $Y2=0
cc_251 N_A4_c_253_n N_Y_c_751_n 0.0113175f $X=3.1 $Y=1.185 $X2=0 $Y2=0
cc_252 N_A4_c_256_n N_Y_c_751_n 0.0109352f $X=3.61 $Y=1.185 $X2=0 $Y2=0
cc_253 N_A4_c_258_n N_Y_c_751_n 0.0109203f $X=4.04 $Y=1.185 $X2=0 $Y2=0
cc_254 N_A4_c_260_n N_Y_c_751_n 0.00804944f $X=4.56 $Y=1.185 $X2=0 $Y2=0
cc_255 N_A4_c_261_n N_Y_c_751_n 0.0153117f $X=4.4 $Y=1.395 $X2=0 $Y2=0
cc_256 N_A4_c_262_n N_Y_c_751_n 0.0926304f $X=3.483 $Y=1.557 $X2=0 $Y2=0
cc_257 N_A4_M1021_g N_Y_c_788_n 0.01115f $X=3.54 $Y=2.435 $X2=0 $Y2=0
cc_258 N_A4_M1024_g N_Y_c_788_n 0.0121857f $X=3.97 $Y=2.435 $X2=0 $Y2=0
cc_259 N_A4_c_300_p N_Y_c_788_n 0.0106412f $X=4.09 $Y=1.44 $X2=0 $Y2=0
cc_260 N_A4_c_261_n N_Y_c_788_n 0.00233422f $X=4.4 $Y=1.395 $X2=0 $Y2=0
cc_261 N_A4_c_263_n N_Y_c_788_n 0.0125202f $X=3.685 $Y=1.557 $X2=0 $Y2=0
cc_262 N_A4_M1021_g N_Y_c_793_n 5.63573e-19 $X=3.54 $Y=2.435 $X2=0 $Y2=0
cc_263 N_A4_M1024_g N_Y_c_793_n 0.00787502f $X=3.97 $Y=2.435 $X2=0 $Y2=0
cc_264 N_A4_M1035_g N_Y_c_793_n 0.00663117f $X=4.4 $Y=2.435 $X2=0 $Y2=0
cc_265 N_A4_M1013_g N_Y_c_796_n 0.0153389f $X=3.11 $Y=2.435 $X2=0 $Y2=0
cc_266 N_A4_M1021_g N_Y_c_796_n 0.0107138f $X=3.54 $Y=2.435 $X2=0 $Y2=0
cc_267 N_A4_M1024_g N_Y_c_796_n 5.63573e-19 $X=3.97 $Y=2.435 $X2=0 $Y2=0
cc_268 N_A4_c_261_n N_Y_c_796_n 5.45588e-19 $X=4.4 $Y=1.395 $X2=0 $Y2=0
cc_269 N_A4_c_262_n N_Y_c_796_n 0.0234531f $X=3.483 $Y=1.557 $X2=0 $Y2=0
cc_270 N_A4_M1024_g Y 5.05234e-19 $X=3.97 $Y=2.435 $X2=0 $Y2=0
cc_271 N_A4_M1035_g Y 0.00277097f $X=4.4 $Y=2.435 $X2=0 $Y2=0
cc_272 N_A4_c_300_p Y 0.0131467f $X=4.09 $Y=1.44 $X2=0 $Y2=0
cc_273 N_A4_c_261_n Y 0.0252721f $X=4.4 $Y=1.395 $X2=0 $Y2=0
cc_274 N_A4_M1021_g N_Y_c_756_n 8.82418e-19 $X=3.54 $Y=2.435 $X2=0 $Y2=0
cc_275 N_A4_M1024_g N_Y_c_756_n 0.00596223f $X=3.97 $Y=2.435 $X2=0 $Y2=0
cc_276 N_A4_M1035_g N_Y_c_756_n 0.0167512f $X=4.4 $Y=2.435 $X2=0 $Y2=0
cc_277 N_A4_c_300_p N_Y_c_756_n 0.0180518f $X=4.09 $Y=1.44 $X2=0 $Y2=0
cc_278 N_A4_c_261_n N_Y_c_756_n 0.0028902f $X=4.4 $Y=1.395 $X2=0 $Y2=0
cc_279 N_A4_c_263_n N_Y_c_756_n 0.00289276f $X=3.685 $Y=1.557 $X2=0 $Y2=0
cc_280 N_A4_M1013_g N_A_554_361#_c_859_n 0.0118654f $X=3.11 $Y=2.435 $X2=0 $Y2=0
cc_281 N_A4_M1021_g N_A_554_361#_c_859_n 0.0117993f $X=3.54 $Y=2.435 $X2=0 $Y2=0
cc_282 N_A4_M1024_g N_A_554_361#_c_861_n 0.0117499f $X=3.97 $Y=2.435 $X2=0 $Y2=0
cc_283 N_A4_M1035_g N_A_554_361#_c_861_n 0.0117779f $X=4.4 $Y=2.435 $X2=0 $Y2=0
cc_284 N_A4_M1035_g N_A_554_361#_c_871_n 3.18291e-19 $X=4.4 $Y=2.435 $X2=0 $Y2=0
cc_285 N_A4_c_253_n N_A_192_47#_c_1088_n 0.0125885f $X=3.1 $Y=1.185 $X2=0 $Y2=0
cc_286 N_A4_c_256_n N_A_192_47#_c_1088_n 0.00908486f $X=3.61 $Y=1.185 $X2=0
+ $Y2=0
cc_287 N_A4_c_253_n N_A_192_47#_c_1090_n 6.31797e-19 $X=3.1 $Y=1.185 $X2=0 $Y2=0
cc_288 N_A4_c_256_n N_A_192_47#_c_1090_n 0.00610136f $X=3.61 $Y=1.185 $X2=0
+ $Y2=0
cc_289 N_A4_c_258_n N_A_192_47#_c_1090_n 0.00613052f $X=4.04 $Y=1.185 $X2=0
+ $Y2=0
cc_290 N_A4_c_260_n N_A_192_47#_c_1090_n 6.26692e-19 $X=4.56 $Y=1.185 $X2=0
+ $Y2=0
cc_291 N_A4_c_258_n N_A_192_47#_c_1094_n 0.00913391f $X=4.04 $Y=1.185 $X2=0
+ $Y2=0
cc_292 N_A4_c_260_n N_A_192_47#_c_1094_n 0.0126874f $X=4.56 $Y=1.185 $X2=0 $Y2=0
cc_293 N_A4_c_260_n N_A_192_47#_c_1096_n 0.00322681f $X=4.56 $Y=1.185 $X2=0
+ $Y2=0
cc_294 N_A4_c_260_n N_A_192_47#_c_1063_n 8.80962e-19 $X=4.56 $Y=1.185 $X2=0
+ $Y2=0
cc_295 N_A4_c_256_n N_A_192_47#_c_1098_n 7.15561e-19 $X=3.61 $Y=1.185 $X2=0
+ $Y2=0
cc_296 N_A4_c_258_n N_A_192_47#_c_1098_n 7.15561e-19 $X=4.04 $Y=1.185 $X2=0
+ $Y2=0
cc_297 N_A4_c_253_n N_VGND_c_1229_n 0.00816542f $X=3.1 $Y=1.185 $X2=0 $Y2=0
cc_298 N_A4_c_256_n N_VGND_c_1229_n 0.00443027f $X=3.61 $Y=1.185 $X2=0 $Y2=0
cc_299 N_A4_c_258_n N_VGND_c_1230_n 0.00447699f $X=4.04 $Y=1.185 $X2=0 $Y2=0
cc_300 N_A4_c_260_n N_VGND_c_1230_n 0.00759674f $X=4.56 $Y=1.185 $X2=0 $Y2=0
cc_301 N_A4_c_253_n N_VGND_c_1239_n 0.00358332f $X=3.1 $Y=1.185 $X2=0 $Y2=0
cc_302 N_A4_c_256_n N_VGND_c_1241_n 0.00420209f $X=3.61 $Y=1.185 $X2=0 $Y2=0
cc_303 N_A4_c_258_n N_VGND_c_1241_n 0.00420209f $X=4.04 $Y=1.185 $X2=0 $Y2=0
cc_304 N_A4_c_260_n N_VGND_c_1243_n 0.00387059f $X=4.56 $Y=1.185 $X2=0 $Y2=0
cc_305 N_A4_c_253_n N_VGND_c_1250_n 0.00449581f $X=3.1 $Y=1.185 $X2=0 $Y2=0
cc_306 N_A4_c_256_n N_VGND_c_1250_n 0.00601396f $X=3.61 $Y=1.185 $X2=0 $Y2=0
cc_307 N_A4_c_258_n N_VGND_c_1250_n 0.00603785f $X=4.04 $Y=1.185 $X2=0 $Y2=0
cc_308 N_A4_c_260_n N_VGND_c_1250_n 0.0047669f $X=4.56 $Y=1.185 $X2=0 $Y2=0
cc_309 N_A3_M1039_g N_A2_M1009_g 0.0202924f $X=6.43 $Y=0.655 $X2=0 $Y2=0
cc_310 A3 N_A2_M1000_g 4.78828e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_311 N_A3_c_355_n N_A2_M1000_g 0.00200098f $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_312 N_A3_M1039_g N_A2_c_459_n 0.00261992f $X=6.43 $Y=0.655 $X2=0 $Y2=0
cc_313 A3 N_A2_c_459_n 9.73923e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_314 N_A3_c_355_n N_A2_c_459_n 0.0195329f $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_315 A3 N_A2_c_460_n 0.036367f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_316 N_A3_c_355_n N_A2_c_460_n 6.45364e-19 $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_317 N_A3_c_356_n N_VPWR_c_631_n 0.00519058f $X=4.83 $Y=1.695 $X2=0 $Y2=0
cc_318 N_A3_c_357_n N_VPWR_c_631_n 0.0033828f $X=5.26 $Y=1.695 $X2=0 $Y2=0
cc_319 N_A3_c_358_n N_VPWR_c_631_n 0.0033828f $X=5.69 $Y=1.695 $X2=0 $Y2=0
cc_320 N_A3_c_359_n N_VPWR_c_631_n 0.0033828f $X=6.12 $Y=1.695 $X2=0 $Y2=0
cc_321 N_A3_c_356_n N_VPWR_c_620_n 0.00974507f $X=4.83 $Y=1.695 $X2=0 $Y2=0
cc_322 N_A3_c_357_n N_VPWR_c_620_n 0.00509122f $X=5.26 $Y=1.695 $X2=0 $Y2=0
cc_323 N_A3_c_358_n N_VPWR_c_620_n 0.00509122f $X=5.69 $Y=1.695 $X2=0 $Y2=0
cc_324 N_A3_c_359_n N_VPWR_c_620_n 0.00619096f $X=6.12 $Y=1.695 $X2=0 $Y2=0
cc_325 N_A3_M1015_g N_Y_c_751_n 5.85447e-19 $X=5.06 $Y=0.655 $X2=0 $Y2=0
cc_326 N_A3_M1015_g Y 0.00250897f $X=5.06 $Y=0.655 $X2=0 $Y2=0
cc_327 A3 Y 0.0294244f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_328 N_A3_c_355_n Y 0.00279179f $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_329 N_A3_c_356_n N_Y_c_756_n 0.00464426f $X=4.83 $Y=1.695 $X2=0 $Y2=0
cc_330 A3 N_Y_c_756_n 0.00391078f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_331 N_A3_c_357_n N_A_554_361#_c_872_n 0.0138154f $X=5.26 $Y=1.695 $X2=0 $Y2=0
cc_332 A3 N_A_554_361#_c_872_n 0.0264899f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_333 N_A3_c_355_n N_A_554_361#_c_872_n 6.13168e-19 $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_334 N_A3_c_356_n N_A_554_361#_c_871_n 0.0191776f $X=4.83 $Y=1.695 $X2=0 $Y2=0
cc_335 A3 N_A_554_361#_c_871_n 0.0099333f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_336 N_A3_c_358_n N_A_554_361#_c_877_n 0.013865f $X=5.69 $Y=1.695 $X2=0 $Y2=0
cc_337 N_A3_c_359_n N_A_554_361#_c_877_n 0.0143809f $X=6.12 $Y=1.695 $X2=0 $Y2=0
cc_338 A3 N_A_554_361#_c_877_n 0.0451315f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_339 N_A3_c_355_n N_A_554_361#_c_877_n 6.2798e-19 $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_340 A3 N_A_554_361#_c_863_n 0.0224129f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_341 N_A3_c_355_n N_A_554_361#_c_863_n 0.00172984f $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_342 A3 N_A_554_361#_c_883_n 0.0156438f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_343 N_A3_c_355_n N_A_554_361#_c_883_n 6.77318e-19 $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_344 N_A3_c_356_n N_A_981_361#_c_928_n 0.00581317f $X=4.83 $Y=1.695 $X2=0
+ $Y2=0
cc_345 N_A3_c_357_n N_A_981_361#_c_928_n 0.00705518f $X=5.26 $Y=1.695 $X2=0
+ $Y2=0
cc_346 N_A3_c_358_n N_A_981_361#_c_928_n 5.16893e-19 $X=5.69 $Y=1.695 $X2=0
+ $Y2=0
cc_347 N_A3_c_357_n N_A_981_361#_c_924_n 0.00964216f $X=5.26 $Y=1.695 $X2=0
+ $Y2=0
cc_348 N_A3_c_358_n N_A_981_361#_c_924_n 0.00964216f $X=5.69 $Y=1.695 $X2=0
+ $Y2=0
cc_349 N_A3_c_356_n N_A_981_361#_c_925_n 0.00251022f $X=4.83 $Y=1.695 $X2=0
+ $Y2=0
cc_350 N_A3_c_357_n N_A_981_361#_c_925_n 7.94187e-19 $X=5.26 $Y=1.695 $X2=0
+ $Y2=0
cc_351 N_A3_c_357_n N_A_981_361#_c_935_n 5.16893e-19 $X=5.26 $Y=1.695 $X2=0
+ $Y2=0
cc_352 N_A3_c_358_n N_A_981_361#_c_935_n 0.00705518f $X=5.69 $Y=1.695 $X2=0
+ $Y2=0
cc_353 N_A3_c_359_n N_A_981_361#_c_935_n 0.0115899f $X=6.12 $Y=1.695 $X2=0 $Y2=0
cc_354 N_A3_c_359_n N_A_981_361#_c_926_n 0.01229f $X=6.12 $Y=1.695 $X2=0 $Y2=0
cc_355 N_A3_c_358_n N_A_981_361#_c_927_n 7.94187e-19 $X=5.69 $Y=1.695 $X2=0
+ $Y2=0
cc_356 N_A3_c_359_n N_A_981_361#_c_927_n 7.94187e-19 $X=6.12 $Y=1.695 $X2=0
+ $Y2=0
cc_357 N_A3_c_359_n N_A_1346_367#_c_991_n 9.27273e-19 $X=6.12 $Y=1.695 $X2=0
+ $Y2=0
cc_358 N_A3_M1015_g N_A_192_47#_c_1100_n 0.00467055f $X=5.06 $Y=0.655 $X2=0
+ $Y2=0
cc_359 N_A3_M1015_g N_A_192_47#_c_1096_n 0.00374685f $X=5.06 $Y=0.655 $X2=0
+ $Y2=0
cc_360 N_A3_M1030_g N_A_192_47#_c_1096_n 3.41721e-19 $X=5.57 $Y=0.655 $X2=0
+ $Y2=0
cc_361 N_A3_M1015_g N_A_192_47#_c_1062_n 0.011225f $X=5.06 $Y=0.655 $X2=0 $Y2=0
cc_362 N_A3_M1030_g N_A_192_47#_c_1062_n 0.0139872f $X=5.57 $Y=0.655 $X2=0 $Y2=0
cc_363 A3 N_A_192_47#_c_1062_n 0.0504576f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_364 N_A3_c_355_n N_A_192_47#_c_1062_n 0.00491309f $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_365 N_A3_M1015_g N_A_192_47#_c_1063_n 0.00239327f $X=5.06 $Y=0.655 $X2=0
+ $Y2=0
cc_366 A3 N_A_192_47#_c_1063_n 0.0144049f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_367 N_A3_c_355_n N_A_192_47#_c_1063_n 0.00395198f $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_368 N_A3_M1034_g N_A_192_47#_c_1064_n 0.013453f $X=6 $Y=0.655 $X2=0 $Y2=0
cc_369 N_A3_M1039_g N_A_192_47#_c_1064_n 0.0134258f $X=6.43 $Y=0.655 $X2=0 $Y2=0
cc_370 A3 N_A_192_47#_c_1064_n 0.0500236f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A3_c_355_n N_A_192_47#_c_1064_n 0.00320968f $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_372 N_A3_M1015_g N_A_192_47#_c_1114_n 0.00190401f $X=5.06 $Y=0.655 $X2=0
+ $Y2=0
cc_373 N_A3_c_355_n N_A_192_47#_c_1114_n 0.0024702f $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_374 A3 N_A_192_47#_c_1069_n 0.0162528f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_375 N_A3_c_355_n N_A_192_47#_c_1069_n 0.00282284f $X=6.37 $Y=1.48 $X2=0 $Y2=0
cc_376 A3 N_A_192_47#_c_1070_n 0.00224441f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_377 N_A3_M1015_g N_VGND_c_1230_n 9.73119e-19 $X=5.06 $Y=0.655 $X2=0 $Y2=0
cc_378 N_A3_M1015_g N_VGND_c_1231_n 0.0062184f $X=5.06 $Y=0.655 $X2=0 $Y2=0
cc_379 N_A3_M1030_g N_VGND_c_1231_n 0.00988398f $X=5.57 $Y=0.655 $X2=0 $Y2=0
cc_380 N_A3_M1034_g N_VGND_c_1231_n 6.12742e-19 $X=6 $Y=0.655 $X2=0 $Y2=0
cc_381 N_A3_M1030_g N_VGND_c_1232_n 6.16059e-19 $X=5.57 $Y=0.655 $X2=0 $Y2=0
cc_382 N_A3_M1034_g N_VGND_c_1232_n 0.0101887f $X=6 $Y=0.655 $X2=0 $Y2=0
cc_383 N_A3_M1039_g N_VGND_c_1232_n 0.010177f $X=6.43 $Y=0.655 $X2=0 $Y2=0
cc_384 N_A3_M1039_g N_VGND_c_1233_n 0.00486043f $X=6.43 $Y=0.655 $X2=0 $Y2=0
cc_385 N_A3_M1039_g N_VGND_c_1234_n 6.14008e-19 $X=6.43 $Y=0.655 $X2=0 $Y2=0
cc_386 N_A3_M1015_g N_VGND_c_1243_n 0.00541359f $X=5.06 $Y=0.655 $X2=0 $Y2=0
cc_387 N_A3_M1030_g N_VGND_c_1245_n 0.00505556f $X=5.57 $Y=0.655 $X2=0 $Y2=0
cc_388 N_A3_M1034_g N_VGND_c_1245_n 0.00486043f $X=6 $Y=0.655 $X2=0 $Y2=0
cc_389 N_A3_M1015_g N_VGND_c_1250_n 0.010095f $X=5.06 $Y=0.655 $X2=0 $Y2=0
cc_390 N_A3_M1030_g N_VGND_c_1250_n 0.00855618f $X=5.57 $Y=0.655 $X2=0 $Y2=0
cc_391 N_A3_M1034_g N_VGND_c_1250_n 0.00824727f $X=6 $Y=0.655 $X2=0 $Y2=0
cc_392 N_A3_M1039_g N_VGND_c_1250_n 0.0082726f $X=6.43 $Y=0.655 $X2=0 $Y2=0
cc_393 N_A2_M1032_g N_A1_c_551_n 0.0202195f $X=8.285 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_394 N_A2_c_459_n N_A1_M1005_g 0.0276558f $X=8.36 $Y=1.44 $X2=0 $Y2=0
cc_395 N_A2_M1032_g A1 3.09326e-19 $X=8.285 $Y=0.655 $X2=0 $Y2=0
cc_396 N_A2_c_458_n A1 0.00879175f $X=8.27 $Y=1.44 $X2=0 $Y2=0
cc_397 N_A2_c_459_n A1 6.00143e-19 $X=8.36 $Y=1.44 $X2=0 $Y2=0
cc_398 N_A2_c_458_n N_A1_c_560_n 7.33669e-19 $X=8.27 $Y=1.44 $X2=0 $Y2=0
cc_399 N_A2_c_459_n N_A1_c_560_n 0.0168297f $X=8.36 $Y=1.44 $X2=0 $Y2=0
cc_400 N_A2_M1025_g N_VPWR_c_624_n 0.00138364f $X=8.36 $Y=2.465 $X2=0 $Y2=0
cc_401 N_A2_M1000_g N_VPWR_c_631_n 0.00357842f $X=7.07 $Y=2.465 $X2=0 $Y2=0
cc_402 N_A2_M1011_g N_VPWR_c_631_n 0.00357842f $X=7.5 $Y=2.465 $X2=0 $Y2=0
cc_403 N_A2_M1020_g N_VPWR_c_631_n 0.00357877f $X=7.93 $Y=2.465 $X2=0 $Y2=0
cc_404 N_A2_M1025_g N_VPWR_c_631_n 0.00547432f $X=8.36 $Y=2.465 $X2=0 $Y2=0
cc_405 N_A2_M1000_g N_VPWR_c_620_n 0.00675085f $X=7.07 $Y=2.465 $X2=0 $Y2=0
cc_406 N_A2_M1011_g N_VPWR_c_620_n 0.00535118f $X=7.5 $Y=2.465 $X2=0 $Y2=0
cc_407 N_A2_M1020_g N_VPWR_c_620_n 0.0053512f $X=7.93 $Y=2.465 $X2=0 $Y2=0
cc_408 N_A2_M1025_g N_VPWR_c_620_n 0.00990114f $X=8.36 $Y=2.465 $X2=0 $Y2=0
cc_409 N_A2_M1000_g N_A_981_361#_c_926_n 0.0145156f $X=7.07 $Y=2.465 $X2=0 $Y2=0
cc_410 N_A2_M1000_g N_A_981_361#_c_942_n 0.00874385f $X=7.07 $Y=2.465 $X2=0
+ $Y2=0
cc_411 N_A2_M1011_g N_A_981_361#_c_942_n 0.00894822f $X=7.5 $Y=2.465 $X2=0 $Y2=0
cc_412 N_A2_M1020_g N_A_981_361#_c_942_n 6.76282e-19 $X=7.93 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_A2_M1011_g N_A_981_361#_c_945_n 0.0126509f $X=7.5 $Y=2.465 $X2=0 $Y2=0
cc_414 N_A2_M1020_g N_A_981_361#_c_945_n 0.0164629f $X=7.93 $Y=2.465 $X2=0 $Y2=0
cc_415 N_A2_M1025_g N_A_981_361#_c_947_n 0.00365671f $X=8.36 $Y=2.465 $X2=0
+ $Y2=0
cc_416 N_A2_M1025_g N_A_981_361#_c_948_n 0.00729561f $X=8.36 $Y=2.465 $X2=0
+ $Y2=0
cc_417 N_A2_M1000_g N_A_981_361#_c_949_n 0.00635181f $X=7.07 $Y=2.465 $X2=0
+ $Y2=0
cc_418 N_A2_M1011_g N_A_981_361#_c_949_n 9.73964e-19 $X=7.5 $Y=2.465 $X2=0 $Y2=0
cc_419 N_A2_c_459_n N_A_1346_367#_c_990_n 0.0011079f $X=8.36 $Y=1.44 $X2=0 $Y2=0
cc_420 N_A2_c_460_n N_A_1346_367#_c_990_n 0.0175025f $X=7.335 $Y=1.547 $X2=0
+ $Y2=0
cc_421 N_A2_M1000_g N_A_1346_367#_c_1002_n 0.0125125f $X=7.07 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A2_M1011_g N_A_1346_367#_c_1002_n 0.0116927f $X=7.5 $Y=2.465 $X2=0
+ $Y2=0
cc_423 N_A2_c_458_n N_A_1346_367#_c_1002_n 0.008158f $X=8.27 $Y=1.44 $X2=0 $Y2=0
cc_424 N_A2_c_459_n N_A_1346_367#_c_1002_n 4.89658e-19 $X=8.36 $Y=1.44 $X2=0
+ $Y2=0
cc_425 N_A2_c_460_n N_A_1346_367#_c_1002_n 0.0258654f $X=7.335 $Y=1.547 $X2=0
+ $Y2=0
cc_426 N_A2_M1020_g N_A_1346_367#_c_1007_n 0.00433465f $X=7.93 $Y=2.465 $X2=0
+ $Y2=0
cc_427 N_A2_M1020_g N_A_1346_367#_c_992_n 0.0125355f $X=7.93 $Y=2.465 $X2=0
+ $Y2=0
cc_428 N_A2_M1025_g N_A_1346_367#_c_992_n 0.0141987f $X=8.36 $Y=2.465 $X2=0
+ $Y2=0
cc_429 N_A2_c_458_n N_A_1346_367#_c_992_n 0.0390092f $X=8.27 $Y=1.44 $X2=0 $Y2=0
cc_430 N_A2_c_459_n N_A_1346_367#_c_992_n 0.00279051f $X=8.36 $Y=1.44 $X2=0
+ $Y2=0
cc_431 N_A2_M1011_g N_A_1346_367#_c_996_n 0.0027321f $X=7.5 $Y=2.465 $X2=0 $Y2=0
cc_432 N_A2_M1020_g N_A_1346_367#_c_996_n 0.00628286f $X=7.93 $Y=2.465 $X2=0
+ $Y2=0
cc_433 N_A2_M1025_g N_A_1346_367#_c_996_n 5.36938e-19 $X=8.36 $Y=2.465 $X2=0
+ $Y2=0
cc_434 N_A2_c_458_n N_A_1346_367#_c_996_n 0.0207876f $X=8.27 $Y=1.44 $X2=0 $Y2=0
cc_435 N_A2_c_459_n N_A_1346_367#_c_996_n 0.00299787f $X=8.36 $Y=1.44 $X2=0
+ $Y2=0
cc_436 N_A2_c_460_n N_A_1346_367#_c_996_n 0.00323096f $X=7.335 $Y=1.547 $X2=0
+ $Y2=0
cc_437 N_A2_M1009_g N_A_192_47#_c_1065_n 0.0134258f $X=6.86 $Y=0.655 $X2=0 $Y2=0
cc_438 N_A2_M1012_g N_A_192_47#_c_1065_n 0.013453f $X=7.29 $Y=0.655 $X2=0 $Y2=0
cc_439 N_A2_c_459_n N_A_192_47#_c_1065_n 0.00383472f $X=8.36 $Y=1.44 $X2=0 $Y2=0
cc_440 N_A2_c_460_n N_A_192_47#_c_1065_n 0.0492415f $X=7.335 $Y=1.547 $X2=0
+ $Y2=0
cc_441 N_A2_M1028_g N_A_192_47#_c_1123_n 0.0107314f $X=7.72 $Y=0.655 $X2=0 $Y2=0
cc_442 N_A2_M1032_g N_A_192_47#_c_1123_n 6.49735e-19 $X=8.285 $Y=0.655 $X2=0
+ $Y2=0
cc_443 N_A2_M1028_g N_A_192_47#_c_1066_n 0.0118478f $X=7.72 $Y=0.655 $X2=0 $Y2=0
cc_444 N_A2_M1032_g N_A_192_47#_c_1066_n 0.0122165f $X=8.285 $Y=0.655 $X2=0
+ $Y2=0
cc_445 N_A2_c_458_n N_A_192_47#_c_1066_n 0.0471008f $X=8.27 $Y=1.44 $X2=0 $Y2=0
cc_446 N_A2_c_459_n N_A_192_47#_c_1066_n 0.00661602f $X=8.36 $Y=1.44 $X2=0 $Y2=0
cc_447 N_A2_M1028_g N_A_192_47#_c_1129_n 2.23836e-19 $X=7.72 $Y=0.655 $X2=0
+ $Y2=0
cc_448 N_A2_M1032_g N_A_192_47#_c_1129_n 0.00781498f $X=8.285 $Y=0.655 $X2=0
+ $Y2=0
cc_449 N_A2_M1028_g N_A_192_47#_c_1071_n 0.00193846f $X=7.72 $Y=0.655 $X2=0
+ $Y2=0
cc_450 N_A2_c_458_n N_A_192_47#_c_1071_n 0.0209452f $X=8.27 $Y=1.44 $X2=0 $Y2=0
cc_451 N_A2_c_459_n N_A_192_47#_c_1071_n 0.00296179f $X=8.36 $Y=1.44 $X2=0 $Y2=0
cc_452 N_A2_M1028_g N_A_192_47#_c_1072_n 4.179e-19 $X=7.72 $Y=0.655 $X2=0 $Y2=0
cc_453 N_A2_M1032_g N_A_192_47#_c_1072_n 0.00422018f $X=8.285 $Y=0.655 $X2=0
+ $Y2=0
cc_454 N_A2_c_458_n N_A_192_47#_c_1072_n 0.00760276f $X=8.27 $Y=1.44 $X2=0 $Y2=0
cc_455 N_A2_c_459_n N_A_192_47#_c_1072_n 0.00222134f $X=8.36 $Y=1.44 $X2=0 $Y2=0
cc_456 N_A2_M1009_g N_VGND_c_1232_n 6.14008e-19 $X=6.86 $Y=0.655 $X2=0 $Y2=0
cc_457 N_A2_M1009_g N_VGND_c_1233_n 0.00486043f $X=6.86 $Y=0.655 $X2=0 $Y2=0
cc_458 N_A2_M1009_g N_VGND_c_1234_n 0.010177f $X=6.86 $Y=0.655 $X2=0 $Y2=0
cc_459 N_A2_M1012_g N_VGND_c_1234_n 0.0103352f $X=7.29 $Y=0.655 $X2=0 $Y2=0
cc_460 N_A2_M1028_g N_VGND_c_1234_n 6.96622e-19 $X=7.72 $Y=0.655 $X2=0 $Y2=0
cc_461 N_A2_M1012_g N_VGND_c_1235_n 0.00486043f $X=7.29 $Y=0.655 $X2=0 $Y2=0
cc_462 N_A2_M1028_g N_VGND_c_1235_n 0.0054895f $X=7.72 $Y=0.655 $X2=0 $Y2=0
cc_463 N_A2_M1028_g N_VGND_c_1236_n 0.00531244f $X=7.72 $Y=0.655 $X2=0 $Y2=0
cc_464 N_A2_M1032_g N_VGND_c_1236_n 0.00540437f $X=8.285 $Y=0.655 $X2=0 $Y2=0
cc_465 N_A2_M1032_g N_VGND_c_1247_n 0.0055654f $X=8.285 $Y=0.655 $X2=0 $Y2=0
cc_466 N_A2_M1009_g N_VGND_c_1250_n 0.0082726f $X=6.86 $Y=0.655 $X2=0 $Y2=0
cc_467 N_A2_M1012_g N_VGND_c_1250_n 0.00824727f $X=7.29 $Y=0.655 $X2=0 $Y2=0
cc_468 N_A2_M1028_g N_VGND_c_1250_n 0.0102076f $X=7.72 $Y=0.655 $X2=0 $Y2=0
cc_469 N_A2_M1032_g N_VGND_c_1250_n 0.0104167f $X=8.285 $Y=0.655 $X2=0 $Y2=0
cc_470 N_A1_M1005_g N_VPWR_c_624_n 0.0163983f $X=8.79 $Y=2.465 $X2=0 $Y2=0
cc_471 N_A1_M1017_g N_VPWR_c_624_n 0.0152057f $X=9.22 $Y=2.465 $X2=0 $Y2=0
cc_472 N_A1_M1023_g N_VPWR_c_624_n 7.41316e-19 $X=9.65 $Y=2.465 $X2=0 $Y2=0
cc_473 N_A1_M1017_g N_VPWR_c_625_n 7.41316e-19 $X=9.22 $Y=2.465 $X2=0 $Y2=0
cc_474 N_A1_M1023_g N_VPWR_c_625_n 0.0152057f $X=9.65 $Y=2.465 $X2=0 $Y2=0
cc_475 N_A1_M1036_g N_VPWR_c_625_n 0.0172133f $X=10.08 $Y=2.465 $X2=0 $Y2=0
cc_476 N_A1_M1005_g N_VPWR_c_631_n 0.00486043f $X=8.79 $Y=2.465 $X2=0 $Y2=0
cc_477 N_A1_M1017_g N_VPWR_c_632_n 0.00486043f $X=9.22 $Y=2.465 $X2=0 $Y2=0
cc_478 N_A1_M1023_g N_VPWR_c_632_n 0.00486043f $X=9.65 $Y=2.465 $X2=0 $Y2=0
cc_479 N_A1_M1036_g N_VPWR_c_633_n 0.00486043f $X=10.08 $Y=2.465 $X2=0 $Y2=0
cc_480 N_A1_M1005_g N_VPWR_c_620_n 0.0082726f $X=8.79 $Y=2.465 $X2=0 $Y2=0
cc_481 N_A1_M1017_g N_VPWR_c_620_n 0.00824727f $X=9.22 $Y=2.465 $X2=0 $Y2=0
cc_482 N_A1_M1023_g N_VPWR_c_620_n 0.00824727f $X=9.65 $Y=2.465 $X2=0 $Y2=0
cc_483 N_A1_M1036_g N_VPWR_c_620_n 0.00918457f $X=10.08 $Y=2.465 $X2=0 $Y2=0
cc_484 N_A1_M1005_g N_A_1346_367#_c_993_n 0.014944f $X=8.79 $Y=2.465 $X2=0 $Y2=0
cc_485 N_A1_M1017_g N_A_1346_367#_c_993_n 0.014237f $X=9.22 $Y=2.465 $X2=0 $Y2=0
cc_486 A1 N_A_1346_367#_c_993_n 0.0436016f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_487 N_A1_c_560_n N_A_1346_367#_c_993_n 0.00206437f $X=10.29 $Y=1.35 $X2=0
+ $Y2=0
cc_488 N_A1_M1023_g N_A_1346_367#_c_994_n 0.014237f $X=9.65 $Y=2.465 $X2=0 $Y2=0
cc_489 N_A1_M1036_g N_A_1346_367#_c_994_n 0.0153768f $X=10.08 $Y=2.465 $X2=0
+ $Y2=0
cc_490 A1 N_A_1346_367#_c_994_n 0.0736238f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_491 N_A1_c_560_n N_A_1346_367#_c_994_n 0.00295582f $X=10.29 $Y=1.35 $X2=0
+ $Y2=0
cc_492 N_A1_c_560_n N_A_1346_367#_c_997_n 8.37869e-19 $X=10.29 $Y=1.35 $X2=0
+ $Y2=0
cc_493 A1 N_A_1346_367#_c_998_n 0.0167501f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_494 N_A1_c_560_n N_A_1346_367#_c_998_n 7.64548e-19 $X=10.29 $Y=1.35 $X2=0
+ $Y2=0
cc_495 N_A1_c_551_n N_A_192_47#_c_1138_n 0.0145448f $X=8.72 $Y=1.185 $X2=0 $Y2=0
cc_496 N_A1_c_553_n N_A_192_47#_c_1138_n 0.0129934f $X=9.15 $Y=1.185 $X2=0 $Y2=0
cc_497 A1 N_A_192_47#_c_1138_n 0.0297913f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_498 N_A1_c_560_n N_A_192_47#_c_1138_n 0.0025922f $X=10.29 $Y=1.35 $X2=0 $Y2=0
cc_499 N_A1_c_555_n N_A_192_47#_c_1067_n 0.0129934f $X=9.58 $Y=1.185 $X2=0 $Y2=0
cc_500 N_A1_c_557_n N_A_192_47#_c_1067_n 0.0127618f $X=10.01 $Y=1.185 $X2=0
+ $Y2=0
cc_501 A1 N_A_192_47#_c_1067_n 0.0609078f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_502 N_A1_c_560_n N_A_192_47#_c_1067_n 0.00939432f $X=10.29 $Y=1.35 $X2=0
+ $Y2=0
cc_503 N_A1_c_551_n N_A_192_47#_c_1072_n 0.00410617f $X=8.72 $Y=1.185 $X2=0
+ $Y2=0
cc_504 A1 N_A_192_47#_c_1147_n 0.0168084f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_505 N_A1_c_560_n N_A_192_47#_c_1147_n 0.00268449f $X=10.29 $Y=1.35 $X2=0
+ $Y2=0
cc_506 N_A1_c_551_n N_VGND_c_1237_n 0.0022121f $X=8.72 $Y=1.185 $X2=0 $Y2=0
cc_507 N_A1_c_553_n N_VGND_c_1237_n 0.00213564f $X=9.15 $Y=1.185 $X2=0 $Y2=0
cc_508 N_A1_c_555_n N_VGND_c_1238_n 0.00213812f $X=9.58 $Y=1.185 $X2=0 $Y2=0
cc_509 N_A1_c_557_n N_VGND_c_1238_n 0.00968522f $X=10.01 $Y=1.185 $X2=0 $Y2=0
cc_510 N_A1_c_551_n N_VGND_c_1247_n 0.00583607f $X=8.72 $Y=1.185 $X2=0 $Y2=0
cc_511 N_A1_c_553_n N_VGND_c_1248_n 0.00585385f $X=9.15 $Y=1.185 $X2=0 $Y2=0
cc_512 N_A1_c_555_n N_VGND_c_1248_n 0.00585385f $X=9.58 $Y=1.185 $X2=0 $Y2=0
cc_513 N_A1_c_557_n N_VGND_c_1249_n 0.00564095f $X=10.01 $Y=1.185 $X2=0 $Y2=0
cc_514 N_A1_c_551_n N_VGND_c_1250_n 0.0106398f $X=8.72 $Y=1.185 $X2=0 $Y2=0
cc_515 N_A1_c_553_n N_VGND_c_1250_n 0.0106161f $X=9.15 $Y=1.185 $X2=0 $Y2=0
cc_516 N_A1_c_555_n N_VGND_c_1250_n 0.0106161f $X=9.58 $Y=1.185 $X2=0 $Y2=0
cc_517 N_A1_c_557_n N_VGND_c_1250_n 0.0104791f $X=10.01 $Y=1.185 $X2=0 $Y2=0
cc_518 N_VPWR_c_620_n N_Y_M1004_s 0.00536646f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_519 N_VPWR_c_620_n N_Y_M1018_s 0.00571434f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_520 N_VPWR_c_626_n N_Y_c_819_n 0.0124525f $X=1.35 $Y=3.33 $X2=0 $Y2=0
cc_521 N_VPWR_c_620_n N_Y_c_819_n 0.00730901f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_522 N_VPWR_M1006_d N_Y_c_759_n 0.00334931f $X=1.375 $Y=1.835 $X2=0 $Y2=0
cc_523 N_VPWR_c_622_n N_Y_c_759_n 0.0170777f $X=1.515 $Y=2.395 $X2=0 $Y2=0
cc_524 N_VPWR_c_628_n N_Y_c_823_n 0.0120977f $X=2.21 $Y=3.33 $X2=0 $Y2=0
cc_525 N_VPWR_c_620_n N_Y_c_823_n 0.00691495f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_526 N_VPWR_M1033_d N_Y_c_754_n 0.00483478f $X=2.235 $Y=1.835 $X2=0 $Y2=0
cc_527 N_VPWR_c_623_n N_Y_c_754_n 0.0220026f $X=2.375 $Y=2.395 $X2=0 $Y2=0
cc_528 N_VPWR_c_623_n N_A_554_361#_c_858_n 0.0472363f $X=2.375 $Y=2.395 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_631_n N_A_554_361#_c_859_n 0.0423919f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_620_n N_A_554_361#_c_859_n 0.0238473f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_623_n N_A_554_361#_c_860_n 0.0147176f $X=2.375 $Y=2.395 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_631_n N_A_554_361#_c_860_n 0.0186386f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_620_n N_A_554_361#_c_860_n 0.0101082f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_631_n N_A_554_361#_c_861_n 0.0423919f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_620_n N_A_554_361#_c_861_n 0.0238473f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_631_n N_A_554_361#_c_862_n 0.0136205f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_620_n N_A_554_361#_c_862_n 0.00738676f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_631_n N_A_554_361#_c_865_n 0.0136205f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_620_n N_A_554_361#_c_865_n 0.00738676f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_620_n N_A_981_361#_M1000_s 0.00223559f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_620_n N_A_981_361#_M1020_s 0.00223562f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_631_n N_A_981_361#_c_924_n 0.0339507f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_620_n N_A_981_361#_c_924_n 0.0188912f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_631_n N_A_981_361#_c_925_n 0.0234809f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_620_n N_A_981_361#_c_925_n 0.0126009f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_631_n N_A_981_361#_c_926_n 0.0660993f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_620_n N_A_981_361#_c_926_n 0.0385512f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_631_n N_A_981_361#_c_945_n 0.0343061f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_620_n N_A_981_361#_c_945_n 0.0215747f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_631_n N_A_981_361#_c_947_n 0.0157917f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_620_n N_A_981_361#_c_947_n 0.00992063f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_631_n N_A_981_361#_c_927_n 0.0234809f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_620_n N_A_981_361#_c_927_n 0.0126009f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_631_n N_A_981_361#_c_949_n 0.01906f $X=8.84 $Y=3.33 $X2=0 $Y2=0
cc_555 N_VPWR_c_620_n N_A_981_361#_c_949_n 0.0124545f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_620_n N_A_1346_367#_M1000_d 0.0021598f $X=10.32 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_557 N_VPWR_c_620_n N_A_1346_367#_M1011_d 0.00225186f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_620_n N_A_1346_367#_M1025_d 0.00536646f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_620_n N_A_1346_367#_M1017_s 0.00536646f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_620_n N_A_1346_367#_M1036_s 0.00371702f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_631_n N_A_1346_367#_c_1034_n 0.0124525f $X=8.84 $Y=3.33 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_620_n N_A_1346_367#_c_1034_n 0.00730901f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_563 N_VPWR_M1005_d N_A_1346_367#_c_993_n 0.00176773f $X=8.865 $Y=1.835 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_624_n N_A_1346_367#_c_993_n 0.0171443f $X=9.005 $Y=2.13 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_632_n N_A_1346_367#_c_1038_n 0.0124525f $X=9.7 $Y=3.33 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_620_n N_A_1346_367#_c_1038_n 0.00730901f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_567 N_VPWR_M1023_d N_A_1346_367#_c_994_n 0.00176773f $X=9.725 $Y=1.835 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_625_n N_A_1346_367#_c_994_n 0.0171443f $X=9.865 $Y=2.13 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_633_n N_A_1346_367#_c_995_n 0.0178111f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_620_n N_A_1346_367#_c_995_n 0.0100304f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_571 N_Y_c_754_n N_A_554_361#_M1013_s 0.00961746f $X=3.16 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_572 N_Y_c_788_n N_A_554_361#_M1021_s 0.00404356f $X=4.02 $Y=2.015 $X2=0 $Y2=0
cc_573 N_Y_c_756_n N_A_554_361#_M1035_s 0.00252733f $X=4.55 $Y=1.705 $X2=0 $Y2=0
cc_574 N_Y_c_754_n N_A_554_361#_c_858_n 0.0202165f $X=3.16 $Y=2.015 $X2=0 $Y2=0
cc_575 N_Y_M1013_d N_A_554_361#_c_859_n 0.00176773f $X=3.185 $Y=1.805 $X2=0
+ $Y2=0
cc_576 N_Y_c_796_n N_A_554_361#_c_859_n 0.0160814f $X=3.325 $Y=2.045 $X2=0 $Y2=0
cc_577 N_Y_c_788_n N_A_554_361#_c_903_n 0.0135055f $X=4.02 $Y=2.015 $X2=0 $Y2=0
cc_578 N_Y_M1024_d N_A_554_361#_c_861_n 0.00176773f $X=4.045 $Y=1.805 $X2=0
+ $Y2=0
cc_579 N_Y_c_793_n N_A_554_361#_c_861_n 0.0160814f $X=4.185 $Y=2.64 $X2=0 $Y2=0
cc_580 N_Y_c_756_n N_A_554_361#_c_871_n 0.0172763f $X=4.55 $Y=1.705 $X2=0 $Y2=0
cc_581 N_Y_c_749_n N_A_192_47#_M1014_s 0.00176461f $X=2.28 $Y=1.1 $X2=0 $Y2=0
cc_582 N_Y_c_751_n N_A_192_47#_M1029_s 0.00261503f $X=4.425 $Y=1.1 $X2=0 $Y2=0
cc_583 N_Y_c_751_n N_A_192_47#_M1008_d 0.00176461f $X=4.425 $Y=1.1 $X2=0 $Y2=0
cc_584 N_Y_c_750_n N_A_192_47#_c_1060_n 0.00166618f $X=1.61 $Y=1.1 $X2=0 $Y2=0
cc_585 N_Y_M1010_d N_A_192_47#_c_1076_n 0.00332344f $X=1.375 $Y=0.235 $X2=0
+ $Y2=0
cc_586 N_Y_c_842_p N_A_192_47#_c_1076_n 0.0124977f $X=1.515 $Y=0.76 $X2=0 $Y2=0
cc_587 N_Y_c_749_n N_A_192_47#_c_1076_n 0.00301993f $X=2.28 $Y=1.1 $X2=0 $Y2=0
cc_588 N_Y_M1026_d N_A_192_47#_c_1078_n 0.00332344f $X=2.235 $Y=0.235 $X2=0
+ $Y2=0
cc_589 N_Y_c_749_n N_A_192_47#_c_1078_n 0.00301993f $X=2.28 $Y=1.1 $X2=0 $Y2=0
cc_590 N_Y_c_846_p N_A_192_47#_c_1078_n 0.0124977f $X=2.375 $Y=0.76 $X2=0 $Y2=0
cc_591 N_Y_c_751_n N_A_192_47#_c_1078_n 0.00301993f $X=4.425 $Y=1.1 $X2=0 $Y2=0
cc_592 N_Y_c_751_n N_A_192_47#_c_1088_n 0.0364735f $X=4.425 $Y=1.1 $X2=0 $Y2=0
cc_593 N_Y_c_751_n N_A_192_47#_c_1083_n 0.0216248f $X=4.425 $Y=1.1 $X2=0 $Y2=0
cc_594 N_Y_c_751_n N_A_192_47#_c_1094_n 0.0384489f $X=4.425 $Y=1.1 $X2=0 $Y2=0
cc_595 N_Y_c_751_n N_A_192_47#_c_1063_n 0.0120256f $X=4.425 $Y=1.1 $X2=0 $Y2=0
cc_596 N_Y_c_749_n N_A_192_47#_c_1084_n 0.016881f $X=2.28 $Y=1.1 $X2=0 $Y2=0
cc_597 N_Y_c_751_n N_A_192_47#_c_1098_n 0.0170334f $X=4.425 $Y=1.1 $X2=0 $Y2=0
cc_598 N_Y_c_751_n N_VGND_M1007_s 0.0026214f $X=4.425 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_599 N_Y_c_751_n N_VGND_M1037_s 0.00268534f $X=4.425 $Y=1.1 $X2=0 $Y2=0
cc_600 N_Y_M1010_d N_VGND_c_1250_n 0.00225186f $X=1.375 $Y=0.235 $X2=0 $Y2=0
cc_601 N_Y_M1026_d N_VGND_c_1250_n 0.00225186f $X=2.235 $Y=0.235 $X2=0 $Y2=0
cc_602 N_A_554_361#_c_872_n N_A_981_361#_M1002_s 0.00260826f $X=5.38 $Y=2.072
+ $X2=-0.19 $Y2=1.655
cc_603 N_A_554_361#_c_871_n N_A_981_361#_M1002_s 7.5685e-19 $X=4.997 $Y=2.072
+ $X2=-0.19 $Y2=1.655
cc_604 N_A_554_361#_c_877_n N_A_981_361#_M1022_s 0.00338201f $X=6.24 $Y=2.072
+ $X2=0 $Y2=0
cc_605 N_A_554_361#_c_872_n N_A_981_361#_c_928_n 0.0129178f $X=5.38 $Y=2.072
+ $X2=0 $Y2=0
cc_606 N_A_554_361#_c_871_n N_A_981_361#_c_928_n 0.00485138f $X=4.997 $Y=2.072
+ $X2=0 $Y2=0
cc_607 N_A_554_361#_M1016_d N_A_981_361#_c_924_n 0.00177869f $X=5.335 $Y=1.805
+ $X2=0 $Y2=0
cc_608 N_A_554_361#_c_872_n N_A_981_361#_c_924_n 0.00302081f $X=5.38 $Y=2.072
+ $X2=0 $Y2=0
cc_609 N_A_554_361#_c_914_p N_A_981_361#_c_924_n 0.0130042f $X=5.475 $Y=2.52
+ $X2=0 $Y2=0
cc_610 N_A_554_361#_c_877_n N_A_981_361#_c_924_n 0.00302081f $X=6.24 $Y=2.072
+ $X2=0 $Y2=0
cc_611 N_A_554_361#_c_862_n N_A_981_361#_c_925_n 0.00803992f $X=4.615 $Y=2.895
+ $X2=0 $Y2=0
cc_612 N_A_554_361#_c_877_n N_A_981_361#_c_935_n 0.0177847f $X=6.24 $Y=2.072
+ $X2=0 $Y2=0
cc_613 N_A_554_361#_M1027_d N_A_981_361#_c_926_n 0.00321202f $X=6.195 $Y=1.805
+ $X2=0 $Y2=0
cc_614 N_A_554_361#_c_877_n N_A_981_361#_c_926_n 0.00303329f $X=6.24 $Y=2.072
+ $X2=0 $Y2=0
cc_615 N_A_554_361#_c_864_n N_A_981_361#_c_926_n 0.0194666f $X=6.335 $Y=2.52
+ $X2=0 $Y2=0
cc_616 N_A_554_361#_c_863_n N_A_1346_367#_c_990_n 0.0155813f $X=6.37 $Y=2.225
+ $X2=0 $Y2=0
cc_617 N_A_554_361#_c_863_n N_A_1346_367#_c_991_n 0.0100121f $X=6.37 $Y=2.225
+ $X2=0 $Y2=0
cc_618 N_A_554_361#_c_864_n N_A_1346_367#_c_991_n 0.0341283f $X=6.335 $Y=2.52
+ $X2=0 $Y2=0
cc_619 N_A_981_361#_c_926_n N_A_1346_367#_M1000_d 0.00522319f $X=7.12 $Y=2.965
+ $X2=-0.19 $Y2=1.655
cc_620 N_A_981_361#_c_945_n N_A_1346_367#_M1011_d 0.00371525f $X=8.05 $Y=2.905
+ $X2=0 $Y2=0
cc_621 N_A_981_361#_c_926_n N_A_1346_367#_c_991_n 0.0194666f $X=7.12 $Y=2.965
+ $X2=0 $Y2=0
cc_622 N_A_981_361#_M1000_s N_A_1346_367#_c_1002_n 0.00353346f $X=7.145 $Y=1.835
+ $X2=0 $Y2=0
cc_623 N_A_981_361#_c_942_n N_A_1346_367#_c_1002_n 0.0171443f $X=7.285 $Y=2.355
+ $X2=0 $Y2=0
cc_624 N_A_981_361#_c_945_n N_A_1346_367#_c_1002_n 0.00297991f $X=8.05 $Y=2.905
+ $X2=0 $Y2=0
cc_625 N_A_981_361#_c_945_n N_A_1346_367#_c_1007_n 0.011418f $X=8.05 $Y=2.905
+ $X2=0 $Y2=0
cc_626 N_A_981_361#_M1020_s N_A_1346_367#_c_992_n 0.00176773f $X=8.005 $Y=1.835
+ $X2=0 $Y2=0
cc_627 N_A_981_361#_c_948_n N_A_1346_367#_c_992_n 0.015351f $X=8.145 $Y=2.21
+ $X2=0 $Y2=0
cc_628 N_A_1346_367#_c_993_n N_A_192_47#_c_1138_n 0.00224249f $X=9.34 $Y=1.785
+ $X2=0 $Y2=0
cc_629 N_A_1346_367#_c_997_n N_A_192_47#_c_1138_n 0.00107422f $X=8.575 $Y=1.785
+ $X2=0 $Y2=0
cc_630 N_A_1346_367#_c_992_n N_A_192_47#_c_1072_n 0.00173699f $X=8.48 $Y=1.785
+ $X2=0 $Y2=0
cc_631 N_A_1346_367#_c_997_n N_A_192_47#_c_1072_n 0.00528662f $X=8.575 $Y=1.785
+ $X2=0 $Y2=0
cc_632 N_A_192_47#_c_1088_n N_VGND_M1007_s 0.00484349f $X=3.66 $Y=0.76 $X2=-0.19
+ $Y2=-0.245
cc_633 N_A_192_47#_c_1094_n N_VGND_M1037_s 0.00509679f $X=4.68 $Y=0.76 $X2=0
+ $Y2=0
cc_634 N_A_192_47#_c_1062_n N_VGND_M1015_d 0.00261503f $X=5.69 $Y=1.09 $X2=0
+ $Y2=0
cc_635 N_A_192_47#_c_1064_n N_VGND_M1034_d 0.00176461f $X=6.55 $Y=1.09 $X2=0
+ $Y2=0
cc_636 N_A_192_47#_c_1065_n N_VGND_M1009_d 0.00176461f $X=7.41 $Y=1.09 $X2=0
+ $Y2=0
cc_637 N_A_192_47#_c_1066_n N_VGND_M1028_d 0.00340974f $X=8.34 $Y=1.09 $X2=0
+ $Y2=0
cc_638 N_A_192_47#_c_1138_n N_VGND_M1001_s 0.00329816f $X=9.24 $Y=0.955 $X2=0
+ $Y2=0
cc_639 N_A_192_47#_c_1067_n N_VGND_M1019_s 0.00329816f $X=10.11 $Y=0.955 $X2=0
+ $Y2=0
cc_640 N_A_192_47#_c_1088_n N_VGND_c_1229_n 0.0206746f $X=3.66 $Y=0.76 $X2=0
+ $Y2=0
cc_641 N_A_192_47#_c_1094_n N_VGND_c_1230_n 0.0207239f $X=4.68 $Y=0.76 $X2=0
+ $Y2=0
cc_642 N_A_192_47#_c_1062_n N_VGND_c_1231_n 0.0214194f $X=5.69 $Y=1.09 $X2=0
+ $Y2=0
cc_643 N_A_192_47#_c_1064_n N_VGND_c_1232_n 0.0170777f $X=6.55 $Y=1.09 $X2=0
+ $Y2=0
cc_644 N_A_192_47#_c_1182_p N_VGND_c_1233_n 0.0124525f $X=6.645 $Y=0.42 $X2=0
+ $Y2=0
cc_645 N_A_192_47#_c_1065_n N_VGND_c_1234_n 0.0170777f $X=7.41 $Y=1.09 $X2=0
+ $Y2=0
cc_646 N_A_192_47#_c_1123_n N_VGND_c_1235_n 0.015688f $X=7.505 $Y=0.42 $X2=0
+ $Y2=0
cc_647 N_A_192_47#_c_1066_n N_VGND_c_1236_n 0.0244889f $X=8.34 $Y=1.09 $X2=0
+ $Y2=0
cc_648 N_A_192_47#_c_1138_n N_VGND_c_1237_n 0.0135055f $X=9.24 $Y=0.955 $X2=0
+ $Y2=0
cc_649 N_A_192_47#_c_1067_n N_VGND_c_1238_n 0.0137681f $X=10.11 $Y=0.955 $X2=0
+ $Y2=0
cc_650 N_A_192_47#_c_1076_n N_VGND_c_1239_n 0.0317578f $X=1.78 $Y=0.34 $X2=0
+ $Y2=0
cc_651 N_A_192_47#_c_1061_n N_VGND_c_1239_n 0.0191601f $X=1.215 $Y=0.34 $X2=0
+ $Y2=0
cc_652 N_A_192_47#_c_1078_n N_VGND_c_1239_n 0.0298674f $X=2.64 $Y=0.34 $X2=0
+ $Y2=0
cc_653 N_A_192_47#_c_1080_n N_VGND_c_1239_n 0.0208666f $X=2.805 $Y=0.425 $X2=0
+ $Y2=0
cc_654 N_A_192_47#_c_1088_n N_VGND_c_1239_n 0.00233949f $X=3.66 $Y=0.76 $X2=0
+ $Y2=0
cc_655 N_A_192_47#_c_1084_n N_VGND_c_1239_n 0.0189074f $X=1.945 $Y=0.38 $X2=0
+ $Y2=0
cc_656 N_A_192_47#_c_1088_n N_VGND_c_1241_n 0.0023334f $X=3.66 $Y=0.76 $X2=0
+ $Y2=0
cc_657 N_A_192_47#_c_1090_n N_VGND_c_1241_n 0.018771f $X=3.825 $Y=0.38 $X2=0
+ $Y2=0
cc_658 N_A_192_47#_c_1094_n N_VGND_c_1241_n 0.0023334f $X=4.68 $Y=0.76 $X2=0
+ $Y2=0
cc_659 N_A_192_47#_c_1094_n N_VGND_c_1243_n 0.0024004f $X=4.68 $Y=0.76 $X2=0
+ $Y2=0
cc_660 N_A_192_47#_c_1100_n N_VGND_c_1243_n 0.0208397f $X=4.845 $Y=0.38 $X2=0
+ $Y2=0
cc_661 N_A_192_47#_c_1199_p N_VGND_c_1245_n 0.0124525f $X=5.785 $Y=0.42 $X2=0
+ $Y2=0
cc_662 N_A_192_47#_c_1129_n N_VGND_c_1247_n 0.0165858f $X=8.5 $Y=0.42 $X2=0
+ $Y2=0
cc_663 N_A_192_47#_c_1201_p N_VGND_c_1248_n 0.0145813f $X=9.365 $Y=0.42 $X2=0
+ $Y2=0
cc_664 N_A_192_47#_c_1068_n N_VGND_c_1249_n 0.0185207f $X=10.225 $Y=0.42 $X2=0
+ $Y2=0
cc_665 N_A_192_47#_M1010_s N_VGND_c_1250_n 0.00215159f $X=0.96 $Y=0.235 $X2=0
+ $Y2=0
cc_666 N_A_192_47#_M1014_s N_VGND_c_1250_n 0.00223559f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_667 N_A_192_47#_M1029_s N_VGND_c_1250_n 0.00311628f $X=2.665 $Y=0.235 $X2=0
+ $Y2=0
cc_668 N_A_192_47#_M1008_d N_VGND_c_1250_n 0.00223559f $X=3.685 $Y=0.235 $X2=0
+ $Y2=0
cc_669 N_A_192_47#_M1038_d N_VGND_c_1250_n 0.00298613f $X=4.635 $Y=0.235 $X2=0
+ $Y2=0
cc_670 N_A_192_47#_M1030_s N_VGND_c_1250_n 0.00536646f $X=5.645 $Y=0.235 $X2=0
+ $Y2=0
cc_671 N_A_192_47#_M1039_s N_VGND_c_1250_n 0.00536646f $X=6.505 $Y=0.235 $X2=0
+ $Y2=0
cc_672 N_A_192_47#_M1012_s N_VGND_c_1250_n 0.00380103f $X=7.365 $Y=0.235 $X2=0
+ $Y2=0
cc_673 N_A_192_47#_M1032_s N_VGND_c_1250_n 0.00297155f $X=8.36 $Y=0.235 $X2=0
+ $Y2=0
cc_674 N_A_192_47#_M1003_d N_VGND_c_1250_n 0.00327921f $X=9.225 $Y=0.235 $X2=0
+ $Y2=0
cc_675 N_A_192_47#_M1031_d N_VGND_c_1250_n 0.00302127f $X=10.085 $Y=0.235 $X2=0
+ $Y2=0
cc_676 N_A_192_47#_c_1076_n N_VGND_c_1250_n 0.0199132f $X=1.78 $Y=0.34 $X2=0
+ $Y2=0
cc_677 N_A_192_47#_c_1061_n N_VGND_c_1250_n 0.0114689f $X=1.215 $Y=0.34 $X2=0
+ $Y2=0
cc_678 N_A_192_47#_c_1078_n N_VGND_c_1250_n 0.0187823f $X=2.64 $Y=0.34 $X2=0
+ $Y2=0
cc_679 N_A_192_47#_c_1080_n N_VGND_c_1250_n 0.0125846f $X=2.805 $Y=0.425 $X2=0
+ $Y2=0
cc_680 N_A_192_47#_c_1088_n N_VGND_c_1250_n 0.0100982f $X=3.66 $Y=0.76 $X2=0
+ $Y2=0
cc_681 N_A_192_47#_c_1090_n N_VGND_c_1250_n 0.0123393f $X=3.825 $Y=0.38 $X2=0
+ $Y2=0
cc_682 N_A_192_47#_c_1094_n N_VGND_c_1250_n 0.0100517f $X=4.68 $Y=0.76 $X2=0
+ $Y2=0
cc_683 N_A_192_47#_c_1100_n N_VGND_c_1250_n 0.0127168f $X=4.845 $Y=0.38 $X2=0
+ $Y2=0
cc_684 N_A_192_47#_c_1199_p N_VGND_c_1250_n 0.00730901f $X=5.785 $Y=0.42 $X2=0
+ $Y2=0
cc_685 N_A_192_47#_c_1182_p N_VGND_c_1250_n 0.00730901f $X=6.645 $Y=0.42 $X2=0
+ $Y2=0
cc_686 N_A_192_47#_c_1123_n N_VGND_c_1250_n 0.00984745f $X=7.505 $Y=0.42 $X2=0
+ $Y2=0
cc_687 N_A_192_47#_c_1129_n N_VGND_c_1250_n 0.0108423f $X=8.5 $Y=0.42 $X2=0
+ $Y2=0
cc_688 N_A_192_47#_c_1201_p N_VGND_c_1250_n 0.00964167f $X=9.365 $Y=0.42 $X2=0
+ $Y2=0
cc_689 N_A_192_47#_c_1068_n N_VGND_c_1250_n 0.010808f $X=10.225 $Y=0.42 $X2=0
+ $Y2=0
cc_690 N_A_192_47#_c_1084_n N_VGND_c_1250_n 0.0124079f $X=1.945 $Y=0.38 $X2=0
+ $Y2=0
