* File: sky130_fd_sc_lp__mux4_0.pex.spice
* Created: Wed Sep  2 10:01:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX4_0%A2 2 3 5 9 13 15 19
c50 13 0 4.79205e-19 $X=1.275 $Y=1.625
c51 3 0 6.26605e-20 $X=1.035 $Y=2.305
r52 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.945
+ $Y=2.08 $X2=0.945 $Y2=2.08
r53 15 19 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=0.72 $Y=2.06
+ $X2=0.945 $Y2=2.06
r54 11 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.035 $Y=1.625
+ $X2=1.275 $Y2=1.625
r55 7 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.275 $Y=1.55
+ $X2=1.275 $Y2=1.625
r56 7 9 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=1.275 $Y=1.55
+ $X2=1.275 $Y2=0.805
r57 3 18 47.986 $w=3.06e-07 $l=2.66224e-07 $layer=POLY_cond $X=1.035 $Y=2.305
+ $X2=0.945 $Y2=2.08
r58 3 5 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.035 $Y=2.305
+ $X2=1.035 $Y2=2.74
r59 2 18 38.535 $w=3.06e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.035 $Y=1.915
+ $X2=0.945 $Y2=2.08
r60 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.035 $Y=1.7
+ $X2=1.035 $Y2=1.625
r61 1 2 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.035 $Y=1.7
+ $X2=1.035 $Y2=1.915
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%S0 2 3 5 10 11 12 13 15 19 21 24 26 27 31 35
+ 37 40 44 47 48 55
c161 44 0 1.67278e-19 $X=1.515 $Y=2.105
c162 40 0 6.26605e-20 $X=1.375 $Y=1.94
c163 24 0 4.04258e-21 $X=3.495 $Y=1.125
c164 19 0 1.18057e-19 $X=2.135 $Y=0.805
c165 13 0 1.87965e-19 $X=1.395 $Y=2.305
r166 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.555
+ $Y=1.54 $X2=0.555 $Y2=1.54
r167 48 55 4.03357 $w=3.85e-07 $l=1.02e-07 $layer=LI1_cond $X=1.2 $Y=1.567
+ $X2=1.098 $Y2=1.567
r168 47 55 11.3149 $w=3.83e-07 $l=3.78e-07 $layer=LI1_cond $X=0.72 $Y=1.567
+ $X2=1.098 $Y2=1.567
r169 47 53 4.93904 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=1.567
+ $X2=0.555 $Y2=1.567
r170 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.515
+ $Y=2.105 $X2=1.515 $Y2=2.105
r171 41 44 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=1.375 $Y=2.065
+ $X2=1.515 $Y2=2.065
r172 40 41 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.375 $Y=1.94
+ $X2=1.375 $Y2=2.065
r173 39 48 7.41319 $w=2.88e-07 $l=2.66503e-07 $layer=LI1_cond $X=1.375 $Y=1.76
+ $X2=1.2 $Y2=1.567
r174 39 40 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.375 $Y=1.76
+ $X2=1.375 $Y2=1.94
r175 29 31 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=3.89 $Y=1.535
+ $X2=3.89 $Y2=2.73
r176 28 38 4.37345 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.6 $Y=1.46 $X2=3.51
+ $Y2=1.46
r177 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.815 $Y=1.46
+ $X2=3.89 $Y2=1.535
r178 27 28 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.815 $Y=1.46
+ $X2=3.6 $Y2=1.46
r179 24 38 101.17 $w=1.6e-07 $l=3.42418e-07 $layer=POLY_cond $X=3.495 $Y=1.125
+ $X2=3.51 $Y2=1.46
r180 24 26 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.495 $Y=1.125
+ $X2=3.495 $Y2=0.805
r181 23 26 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.495 $Y=0.255
+ $X2=3.495 $Y2=0.805
r182 22 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.21 $Y=0.18
+ $X2=2.135 $Y2=0.18
r183 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.42 $Y=0.18
+ $X2=3.495 $Y2=0.255
r184 21 22 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=3.42 $Y=0.18
+ $X2=2.21 $Y2=0.18
r185 17 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.135 $Y=0.255
+ $X2=2.135 $Y2=0.18
r186 17 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.135 $Y=0.255
+ $X2=2.135 $Y2=0.805
r187 13 45 43.6313 $w=3.42e-07 $l=2.46982e-07 $layer=POLY_cond $X=1.395 $Y=2.305
+ $X2=1.5 $Y2=2.105
r188 13 15 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.395 $Y=2.305
+ $X2=1.395 $Y2=2.74
r189 11 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.06 $Y=0.18
+ $X2=2.135 $Y2=0.18
r190 11 12 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=2.06 $Y=0.18
+ $X2=0.92 $Y2=0.18
r191 8 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=1.19
+ $X2=0.845 $Y2=1.265
r192 8 10 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.845 $Y=1.19
+ $X2=0.845 $Y2=0.805
r193 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.845 $Y=0.255
+ $X2=0.92 $Y2=0.18
r194 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.845 $Y=0.255
+ $X2=0.845 $Y2=0.805
r195 3 52 80.7642 $w=2.46e-07 $l=4.03887e-07 $layer=POLY_cond $X=0.495 $Y=1.915
+ $X2=0.555 $Y2=1.54
r196 3 5 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=0.495 $Y=1.915
+ $X2=0.495 $Y2=2.74
r197 2 52 3.22709 $w=3.3e-07 $l=8.75758e-08 $layer=POLY_cond $X=0.555 $Y=1.54
+ $X2=0.555 $Y2=1.54
r198 1 35 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.555 $Y=1.265
+ $X2=0.845 $Y2=1.265
r199 1 2 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.555 $Y=1.34 $X2=0.555
+ $Y2=1.54
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%A_31_506# 1 2 9 13 17 21 23 24 26 28 31 33 37
+ 39 43 44 47 51 52 53 57 58 59 61 67 68 73 80
c193 61 0 1.83003e-19 $X=4.735 $Y=2.075
c194 47 0 2.82839e-19 $X=1.725 $Y=1.52
c195 42 0 9.03317e-20 $X=1.22 $Y=2.905
c196 39 0 1.53137e-19 $X=1.485 $Y=1.12
c197 26 0 3.36516e-20 $X=4.83 $Y=1.91
c198 13 0 1.85747e-19 $X=2.055 $Y=2.73
r199 62 80 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=4.735 $Y=2.075
+ $X2=4.83 $Y2=2.075
r200 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.735
+ $Y=2.075 $X2=4.735 $Y2=2.075
r201 59 61 60.1275 $w=2.28e-07 $l=1.2e-06 $layer=LI1_cond $X=3.535 $Y=2.045
+ $X2=4.735 $Y2=2.045
r202 58 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=2.195
+ $X2=3.44 $Y2=2.36
r203 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=2.195 $X2=3.44 $Y2=2.195
r204 55 57 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=3.405 $Y=2.3
+ $X2=3.405 $Y2=2.195
r205 54 59 6.84978 $w=2.3e-07 $l=1.78466e-07 $layer=LI1_cond $X=3.405 $Y=2.16
+ $X2=3.535 $Y2=2.045
r206 54 57 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=3.405 $Y=2.16
+ $X2=3.405 $Y2=2.195
r207 52 55 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.275 $Y=2.385
+ $X2=3.405 $Y2=2.3
r208 52 53 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.275 $Y=2.385
+ $X2=2.5 $Y2=2.385
r209 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.415 $Y=2.47
+ $X2=2.5 $Y2=2.385
r210 50 51 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.415 $Y=2.47
+ $X2=2.415 $Y2=2.905
r211 48 73 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.725 $Y=1.52
+ $X2=2.055 $Y2=1.52
r212 48 70 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.725 $Y=1.52
+ $X2=1.635 $Y2=1.52
r213 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.52 $X2=1.725 $Y2=1.52
r214 45 69 2.36997 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=1.365
+ $X2=1.725 $Y2=1.2
r215 45 47 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.725 $Y=1.365
+ $X2=1.725 $Y2=1.52
r216 43 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.33 $Y=2.99
+ $X2=2.415 $Y2=2.905
r217 43 44 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.33 $Y=2.99
+ $X2=1.305 $Y2=2.99
r218 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=2.905
+ $X2=1.305 $Y2=2.99
r219 41 42 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.22 $Y=2.53
+ $X2=1.22 $Y2=2.905
r220 39 69 12.9425 $w=2.51e-07 $l=2.77128e-07 $layer=LI1_cond $X=1.485 $Y=1.12
+ $X2=1.725 $Y2=1.2
r221 39 67 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.485 $Y=1.12
+ $X2=0.725 $Y2=1.12
r222 35 67 8.05689 $w=1.78e-07 $l=1.3e-07 $layer=LI1_cond $X=0.595 $Y=1.115
+ $X2=0.725 $Y2=1.115
r223 35 64 23.9071 $w=1.78e-07 $l=3.88e-07 $layer=LI1_cond $X=0.595 $Y=1.115
+ $X2=0.207 $Y2=1.115
r224 35 37 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.595 $Y=1.025
+ $X2=0.595 $Y2=0.805
r225 34 68 2.87242 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.445
+ $X2=0.28 $Y2=2.445
r226 33 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.135 $Y=2.445
+ $X2=1.22 $Y2=2.53
r227 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.135 $Y=2.445
+ $X2=0.445 $Y2=2.445
r228 29 68 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.53
+ $X2=0.28 $Y2=2.445
r229 29 31 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.28 $Y=2.53
+ $X2=0.28 $Y2=2.74
r230 28 68 3.6114 $w=2.57e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.207 $Y=2.36
+ $X2=0.28 $Y2=2.445
r231 27 64 0.5826 $w=1.85e-07 $l=9e-08 $layer=LI1_cond $X=0.207 $Y=1.205
+ $X2=0.207 $Y2=1.115
r232 27 28 69.2432 $w=1.83e-07 $l=1.155e-06 $layer=LI1_cond $X=0.207 $Y=1.205
+ $X2=0.207 $Y2=2.36
r233 26 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.83 $Y=1.91
+ $X2=4.83 $Y2=2.075
r234 25 26 848.628 $w=1.5e-07 $l=1.655e-06 $layer=POLY_cond $X=4.83 $Y=0.255
+ $X2=4.83 $Y2=1.91
r235 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.755 $Y=0.18
+ $X2=4.83 $Y2=0.255
r236 23 24 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=4.755 $Y=0.18
+ $X2=4 $Y2=0.18
r237 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.925 $Y=0.255
+ $X2=4 $Y2=0.18
r238 19 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.925 $Y=0.255
+ $X2=3.925 $Y2=0.805
r239 17 77 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.35 $Y=2.73
+ $X2=3.35 $Y2=2.36
r240 11 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.055 $Y=1.685
+ $X2=2.055 $Y2=1.52
r241 11 13 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=2.055 $Y=1.685
+ $X2=2.055 $Y2=2.73
r242 7 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.355
+ $X2=1.635 $Y2=1.52
r243 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.635 $Y=1.355
+ $X2=1.635 $Y2=0.805
r244 2 31 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=2.53 $X2=0.28 $Y2=2.74
r245 1 37 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.505
+ $Y=0.595 $X2=0.63 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%A3 3 7 9 12
r42 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=2.035
+ $X2=2.505 $Y2=2.2
r43 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=2.035
+ $X2=2.505 $Y2=1.87
r44 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.505
+ $Y=2.035 $X2=2.505 $Y2=2.035
r45 9 13 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=2.64 $Y=2.03
+ $X2=2.505 $Y2=2.03
r46 7 14 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=2.495 $Y=0.805
+ $X2=2.495 $Y2=1.87
r47 3 15 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.415 $Y=2.73
+ $X2=2.415 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%A1 3 7 11 12 14 16 25
c52 11 0 1.82378e-19 $X=3.045 $Y=1.655
r53 14 16 10.7939 $w=6.13e-07 $l=5.55e-07 $layer=LI1_cond $X=3.045 $Y=1.452
+ $X2=3.6 $Y2=1.452
r54 14 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.045
+ $Y=1.315 $X2=3.045 $Y2=1.315
r55 12 14 7.87661 $w=6.13e-07 $l=4.05e-07 $layer=LI1_cond $X=2.64 $Y=1.452
+ $X2=3.045 $Y2=1.452
r56 11 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.045 $Y=1.655
+ $X2=3.045 $Y2=1.315
r57 10 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.045 $Y=1.15
+ $X2=3.045 $Y2=1.315
r58 7 10 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=3.135 $Y=0.805
+ $X2=3.135 $Y2=1.15
r59 1 11 71.2267 $w=2.47e-07 $l=3.91535e-07 $layer=POLY_cond $X=2.99 $Y=2.02
+ $X2=3.045 $Y2=1.655
r60 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.99 $Y=2.02 $X2=2.99
+ $Y2=2.73
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%A0 1 3 5 7 8
c38 8 0 4.04258e-21 $X=4.56 $Y=1.295
c39 1 0 1.83003e-19 $X=4.25 $Y=1.61
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.38
+ $Y=1.295 $X2=4.38 $Y2=1.295
r41 8 12 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=4.56 $Y=1.265
+ $X2=4.38 $Y2=1.265
r42 5 11 38.6342 $w=2.88e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.285 $Y=1.13
+ $X2=4.36 $Y2=1.295
r43 5 7 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=4.285 $Y=1.13
+ $X2=4.285 $Y2=0.805
r44 1 11 63.7384 $w=2.88e-07 $l=3.65889e-07 $layer=POLY_cond $X=4.25 $Y=1.61
+ $X2=4.36 $Y2=1.295
r45 1 3 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=4.25 $Y=1.61 $X2=4.25
+ $Y2=2.73
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%A_1029_37# 1 2 9 12 14 15 19 24 27 30 33 34
+ 37 39 43
c91 30 0 3.3992e-20 $X=6.4 $Y=1.69
r92 36 39 5.19411 $w=3.53e-07 $l=1.6e-07 $layer=LI1_cond $X=6.4 $Y=0.432
+ $X2=6.56 $Y2=0.432
r93 36 37 4.03829 $w=3.53e-07 $l=9e-08 $layer=LI1_cond $X=6.4 $Y=0.432 $X2=6.31
+ $Y2=0.432
r94 33 34 7.81899 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.465 $Y=2.225
+ $X2=6.465 $Y2=2.06
r95 29 30 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=6.395 $Y=1.69 $X2=6.4
+ $Y2=1.69
r96 27 46 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.215 $Y=1.69
+ $X2=6.215 $Y2=1.85
r97 26 29 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=6.215 $Y=1.69
+ $X2=6.395 $Y2=1.69
r98 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=1.69 $X2=6.215 $Y2=1.69
r99 24 30 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.4 $Y=1.525 $X2=6.4
+ $Y2=1.69
r100 23 36 4.71797 $w=1.8e-07 $l=1.78e-07 $layer=LI1_cond $X=6.4 $Y=0.61 $X2=6.4
+ $Y2=0.432
r101 23 24 56.3788 $w=1.78e-07 $l=9.15e-07 $layer=LI1_cond $X=6.4 $Y=0.61
+ $X2=6.4 $Y2=1.525
r102 21 29 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=1.855
+ $X2=6.395 $Y2=1.69
r103 21 34 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=6.395 $Y=1.855
+ $X2=6.395 $Y2=2.06
r104 19 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=0.35
+ $X2=5.31 $Y2=0.515
r105 18 37 47.0385 $w=2.43e-07 $l=1e-06 $layer=LI1_cond $X=5.31 $Y=0.377
+ $X2=6.31 $Y2=0.377
r106 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.31
+ $Y=0.35 $X2=5.31 $Y2=0.35
r107 14 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.05 $Y=1.85
+ $X2=6.215 $Y2=1.85
r108 14 15 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=6.05 $Y=1.85
+ $X2=5.805 $Y2=1.85
r109 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.73 $Y=1.925
+ $X2=5.805 $Y2=1.85
r110 10 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.73 $Y=1.925
+ $X2=5.73 $Y2=2.675
r111 9 43 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.33 $Y=0.835
+ $X2=5.33 $Y2=0.515
r112 2 33 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=6.34
+ $Y=2.015 $X2=6.465 $Y2=2.225
r113 1 39 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=6.435
+ $Y=0.235 $X2=6.56 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%S1 3 5 6 7 9 10 14 18 20 23 25 26 27 28 33
c98 33 0 1.4009e-19 $X=6.755 $Y=1.32
c99 23 0 1.42172e-19 $X=6.755 $Y=1.23
c100 20 0 3.3992e-20 $X=5.747 $Y=1.23
c101 14 0 2.90591e-20 $X=6.68 $Y=2.225
c102 10 0 1.42075e-19 $X=6.59 $Y=1.23
c103 6 0 1.38929e-19 $X=5.375 $Y=1.49
r104 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.755
+ $Y=1.32 $X2=6.755 $Y2=1.32
r105 28 34 9.06917 $w=4.53e-07 $l=3.45e-07 $layer=LI1_cond $X=6.887 $Y=1.665
+ $X2=6.887 $Y2=1.32
r106 27 34 0.657186 $w=4.53e-07 $l=2.5e-08 $layer=LI1_cond $X=6.887 $Y=1.295
+ $X2=6.887 $Y2=1.32
r107 26 27 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=6.887 $Y=0.925
+ $X2=6.887 $Y2=1.295
r108 24 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.755 $Y=1.66
+ $X2=6.755 $Y2=1.32
r109 24 25 43.7316 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.755 $Y=1.66
+ $X2=6.755 $Y2=1.825
r110 22 33 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.755 $Y=1.305
+ $X2=6.755 $Y2=1.32
r111 22 23 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=6.755 $Y=1.305
+ $X2=6.755 $Y2=1.23
r112 20 21 78.8176 $w=1.59e-07 $l=2.6e-07 $layer=POLY_cond $X=5.747 $Y=1.23
+ $X2=5.747 $Y2=1.49
r113 16 23 13.5877 $w=2.4e-07 $l=8.44097e-08 $layer=POLY_cond $X=6.775 $Y=1.155
+ $X2=6.755 $Y2=1.23
r114 16 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.775 $Y=1.155
+ $X2=6.775 $Y2=0.445
r115 14 25 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=6.68 $Y=2.225
+ $X2=6.68 $Y2=1.825
r116 11 20 4.22461 $w=1.5e-07 $l=8.8e-08 $layer=POLY_cond $X=5.835 $Y=1.23
+ $X2=5.747 $Y2=1.23
r117 10 23 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.59 $Y=1.23
+ $X2=6.755 $Y2=1.23
r118 10 11 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=6.59 $Y=1.23
+ $X2=5.835 $Y2=1.23
r119 7 20 22.9461 $w=1.59e-07 $l=8.12404e-08 $layer=POLY_cond $X=5.76 $Y=1.155
+ $X2=5.747 $Y2=1.23
r120 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.76 $Y=1.155
+ $X2=5.76 $Y2=0.835
r121 5 21 4.22461 $w=1.5e-07 $l=8.7e-08 $layer=POLY_cond $X=5.66 $Y=1.49
+ $X2=5.747 $Y2=1.49
r122 5 6 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.66 $Y=1.49
+ $X2=5.375 $Y2=1.49
r123 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.3 $Y=1.565
+ $X2=5.375 $Y2=1.49
r124 1 3 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=5.3 $Y=1.565 $X2=5.3
+ $Y2=2.675
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%A_1075_493# 1 2 7 11 15 18 19 20 21 25 27 29
+ 33 35 37
c75 25 0 3.36516e-20 $X=5.515 $Y=2.74
c76 19 0 3.32533e-19 $X=7.22 $Y=0.915
r77 34 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.58 $Y=2.945 $X2=6.58
+ $Y2=2.855
r78 33 35 8.49766 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=6.58 $Y=2.927
+ $X2=6.415 $Y2=2.927
r79 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.58
+ $Y=2.945 $X2=6.58 $Y2=2.945
r80 29 31 9.15117 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=5.53 $Y=0.835
+ $X2=5.53 $Y2=1.005
r81 27 35 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=5.61 $Y=2.99
+ $X2=6.415 $Y2=2.99
r82 25 31 101.278 $w=1.88e-07 $l=1.735e-06 $layer=LI1_cond $X=5.515 $Y=2.74
+ $X2=5.515 $Y2=1.005
r83 23 27 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.515 $Y=2.905
+ $X2=5.61 $Y2=2.99
r84 23 25 9.63158 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.515 $Y=2.905
+ $X2=5.515 $Y2=2.74
r85 20 21 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=7.22 $Y=1.755
+ $X2=7.22 $Y2=1.905
r86 19 20 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=7.235 $Y=0.915
+ $X2=7.235 $Y2=1.755
r87 18 19 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=7.22 $Y=0.765
+ $X2=7.22 $Y2=0.915
r88 15 21 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.205 $Y=2.335
+ $X2=7.205 $Y2=1.905
r89 13 15 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.205 $Y=2.78
+ $X2=7.205 $Y2=2.335
r90 11 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.205 $Y=0.445
+ $X2=7.205 $Y2=0.765
r91 8 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.745 $Y=2.855
+ $X2=6.58 $Y2=2.855
r92 7 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.13 $Y=2.855
+ $X2=7.205 $Y2=2.78
r93 7 8 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.13 $Y=2.855
+ $X2=6.745 $Y2=2.855
r94 2 25 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=5.375
+ $Y=2.465 $X2=5.515 $Y2=2.74
r95 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.625 $X2=5.545 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%VPWR 1 2 3 4 15 19 23 25 27 29 32 34 35 36 38
+ 50 59 60 63 66 69
r89 69 70 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r90 67 70 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.96 $Y2=3.33
r91 66 67 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r92 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r93 60 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r94 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r95 57 69 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.095 $Y=3.33 $X2=7.005
+ $Y2=3.33
r96 57 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.095 $Y=3.33
+ $X2=7.44 $Y2=3.33
r97 56 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r98 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r99 52 55 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33 $X2=4.08
+ $Y2=3.33
r100 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 50 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=3.33
+ $X2=4.465 $Y2=3.33
r102 50 55 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.3 $Y=3.33
+ $X2=4.08 $Y2=3.33
r103 49 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r104 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 46 49 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 46 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 45 48 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r108 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 43 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r110 43 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 41 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 38 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r114 38 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r115 36 56 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r116 36 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.12 $Y2=3.33
r117 34 48 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=3.33 $X2=2.64
+ $Y2=3.33
r118 34 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.795 $Y2=3.33
r119 33 52 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.92 $Y=3.33 $X2=3.12
+ $Y2=3.33
r120 33 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.92 $Y=3.33
+ $X2=2.795 $Y2=3.33
r121 32 69 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.005 $Y=3.245
+ $X2=7.005 $Y2=3.33
r122 31 32 35.1212 $w=1.78e-07 $l=5.7e-07 $layer=LI1_cond $X=7.005 $Y=2.675
+ $X2=7.005 $Y2=3.245
r123 27 31 9.31882 $w=2.71e-07 $l=2.34211e-07 $layer=LI1_cond $X=6.947 $Y=2.468
+ $X2=7.005 $Y2=2.675
r124 27 29 12.0323 $w=2.93e-07 $l=3.08e-07 $layer=LI1_cond $X=6.947 $Y=2.468
+ $X2=6.947 $Y2=2.16
r125 26 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=3.33
+ $X2=4.465 $Y2=3.33
r126 25 69 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=6.915 $Y=3.33
+ $X2=7.005 $Y2=3.33
r127 25 26 149.075 $w=1.68e-07 $l=2.285e-06 $layer=LI1_cond $X=6.915 $Y=3.33
+ $X2=4.63 $Y2=3.33
r128 21 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=3.245
+ $X2=4.465 $Y2=3.33
r129 21 23 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=4.465 $Y=3.245
+ $X2=4.465 $Y2=2.775
r130 17 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=3.245
+ $X2=2.795 $Y2=3.33
r131 17 19 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=2.795 $Y=3.245
+ $X2=2.795 $Y2=2.805
r132 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r133 13 15 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.805
r134 4 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.755
+ $Y=2.015 $X2=6.895 $Y2=2.16
r135 3 23 600 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=2.52 $X2=4.465 $Y2=2.775
r136 2 19 600 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=1 $X=2.49
+ $Y=2.52 $X2=2.755 $Y2=2.805
r137 1 15 600 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.53 $X2=0.78 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%A_294_506# 1 2 3 4 13 18 23 25 26 28 29 35 39
+ 43
c119 35 0 1.42075e-19 $X=6 $Y=0.925
c120 29 0 3.50795e-20 $X=2.305 $Y=0.925
c121 26 0 2.90591e-20 $X=5.945 $Y=2.46
c122 18 0 3.13049e-20 $X=2.075 $Y=2.475
r123 42 43 5.25278 $w=3.6e-07 $l=1.55e-07 $layer=LI1_cond $X=1.92 $Y=0.827
+ $X2=2.075 $Y2=0.827
r124 35 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0.925 $X2=6
+ $Y2=0.925
r125 32 43 2.88056 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.827
+ $X2=2.075 $Y2=0.827
r126 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=0.925
r127 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=0.925
+ $X2=2.16 $Y2=0.925
r128 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.855 $Y=0.925
+ $X2=6 $Y2=0.925
r129 28 29 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=5.855 $Y=0.925
+ $X2=2.305 $Y2=0.925
r130 25 26 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.945 $Y=2.625
+ $X2=5.945 $Y2=2.46
r131 23 26 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.865 $Y=1.345
+ $X2=5.865 $Y2=2.46
r132 22 39 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.975 $Y=1.175
+ $X2=5.975 $Y2=0.835
r133 22 23 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.96 $Y=1.175
+ $X2=5.96 $Y2=1.345
r134 17 43 5.14255 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=2.075 $Y=1.015
+ $X2=2.075 $Y2=0.827
r135 17 18 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.075 $Y=1.015
+ $X2=2.075 $Y2=2.475
r136 13 18 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.99 $Y=2.605
+ $X2=2.075 $Y2=2.475
r137 13 15 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=1.99 $Y=2.605
+ $X2=1.725 $Y2=2.605
r138 4 25 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=2.465 $X2=5.945 $Y2=2.625
r139 3 15 600 $w=1.7e-07 $l=3.05082e-07 $layer=licon1_PDIFF $count=1 $X=1.47
+ $Y=2.53 $X2=1.725 $Y2=2.64
r140 2 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.835
+ $Y=0.625 $X2=5.975 $Y2=0.835
r141 1 42 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=1.71
+ $Y=0.595 $X2=1.92 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%A_685_504# 1 2 3 4 14 16 17 18 19 20 23 27 30
+ 34 39 41 42
c90 42 0 1.38929e-19 $X=5.1 $Y=1.645
c91 20 0 1.09665e-19 $X=4.035 $Y=1.645
c92 16 0 7.27131e-20 $X=3.95 $Y=1.56
c93 14 0 1.9902e-19 $X=3.79 $Y=2.64
r94 37 39 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.71 $Y=0.805
+ $X2=3.95 $Y2=0.805
r95 32 34 6.99698 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=3.62 $Y=2.78
+ $X2=3.79 $Y2=2.78
r96 30 41 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.165 $Y=2.33
+ $X2=5.085 $Y2=2.415
r97 29 42 3.91525 $w=2.35e-07 $l=1.12916e-07 $layer=LI1_cond $X=5.165 $Y=1.73
+ $X2=5.1 $Y2=1.645
r98 29 30 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.165 $Y=1.73
+ $X2=5.165 $Y2=2.33
r99 25 42 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=1.56 $X2=5.1
+ $Y2=1.645
r100 25 27 27.8507 $w=2.98e-07 $l=7.25e-07 $layer=LI1_cond $X=5.1 $Y=1.56
+ $X2=5.1 $Y2=0.835
r101 21 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=2.5
+ $X2=5.085 $Y2=2.415
r102 21 23 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=5.085 $Y=2.5
+ $X2=5.085 $Y2=2.675
r103 19 42 2.53056 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.95 $Y=1.645
+ $X2=5.1 $Y2=1.645
r104 19 20 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=4.95 $Y=1.645
+ $X2=4.035 $Y2=1.645
r105 17 41 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.92 $Y=2.415
+ $X2=5.085 $Y2=2.415
r106 17 18 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=4.92 $Y=2.415
+ $X2=3.875 $Y2=2.415
r107 16 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.95 $Y=1.56
+ $X2=4.035 $Y2=1.645
r108 15 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.95 $Y=0.97
+ $X2=3.95 $Y2=0.805
r109 15 16 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.95 $Y=0.97
+ $X2=3.95 $Y2=1.56
r110 14 34 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.79 $Y=2.64
+ $X2=3.79 $Y2=2.78
r111 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.79 $Y=2.5
+ $X2=3.875 $Y2=2.415
r112 13 14 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.79 $Y=2.5
+ $X2=3.79 $Y2=2.64
r113 4 23 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=2.465 $X2=5.085 $Y2=2.675
r114 3 32 600 $w=1.7e-07 $l=3.17884e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=2.52 $X2=3.62 $Y2=2.755
r115 2 27 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=4.99
+ $Y=0.625 $X2=5.115 $Y2=0.835
r116 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.595 $X2=3.71 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%X 1 2 7 8 9 10 11 18
r18 11 31 4.80185 $w=2.98e-07 $l=1.25e-07 $layer=LI1_cond $X=7.435 $Y=2.035
+ $X2=7.435 $Y2=2.16
r19 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=7.435 $Y=1.665
+ $X2=7.435 $Y2=2.035
r20 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=7.435 $Y=1.295
+ $X2=7.435 $Y2=1.665
r21 8 9 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=7.435 $Y=0.925
+ $X2=7.435 $Y2=1.295
r22 7 8 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=7.435 $Y=0.555
+ $X2=7.435 $Y2=0.925
r23 7 18 4.22562 $w=2.98e-07 $l=1.1e-07 $layer=LI1_cond $X=7.435 $Y=0.555
+ $X2=7.435 $Y2=0.445
r24 2 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.28
+ $Y=2.015 $X2=7.42 $Y2=2.16
r25 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.28
+ $Y=0.235 $X2=7.42 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_0%VGND 1 2 3 4 15 19 23 27 30 31 32 34 43 50 60
+ 61 64 67 70
c86 61 0 1.6034e-19 $X=7.44 $Y=0
c87 60 0 1.72194e-19 $X=7.44 $Y=0
c88 27 0 1.42172e-19 $X=6.99 $Y=0.445
r89 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r90 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r91 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 61 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r93 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r94 58 70 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=7.115 $Y=0 $X2=6.987
+ $Y2=0
r95 58 60 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.115 $Y=0 $X2=7.44
+ $Y2=0
r96 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r97 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r98 54 57 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r99 54 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r100 53 56 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r101 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r102 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=0 $X2=4.5
+ $Y2=0
r103 51 53 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.665 $Y=0
+ $X2=5.04 $Y2=0
r104 50 70 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=6.86 $Y=0 $X2=6.987
+ $Y2=0
r105 50 56 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.86 $Y=0 $X2=6.48
+ $Y2=0
r106 49 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r107 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r108 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r109 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r110 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.5
+ $Y2=0
r111 43 48 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=4.08 $Y2=0
r112 42 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r113 42 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.2
+ $Y2=0
r114 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r115 39 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.06
+ $Y2=0
r116 39 41 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=1.225 $Y=0
+ $X2=2.64 $Y2=0
r117 37 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r118 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r119 34 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.06
+ $Y2=0
r120 34 36 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.72 $Y2=0
r121 32 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r122 32 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.12
+ $Y2=0
r123 30 41 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.655 $Y=0 $X2=2.64
+ $Y2=0
r124 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=0 $X2=2.82
+ $Y2=0
r125 29 45 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.985 $Y=0
+ $X2=3.12 $Y2=0
r126 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=2.82
+ $Y2=0
r127 25 70 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=6.987 $Y=0.085
+ $X2=6.987 $Y2=0
r128 25 27 16.2698 $w=2.53e-07 $l=3.6e-07 $layer=LI1_cond $X=6.987 $Y=0.085
+ $X2=6.987 $Y2=0.445
r129 21 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=0.085 $X2=4.5
+ $Y2=0
r130 21 23 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=4.5 $Y=0.085
+ $X2=4.5 $Y2=0.805
r131 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=0.085
+ $X2=2.82 $Y2=0
r132 17 19 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=2.82 $Y=0.085
+ $X2=2.82 $Y2=0.805
r133 13 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=0.085
+ $X2=1.06 $Y2=0
r134 13 15 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=1.06 $Y=0.085
+ $X2=1.06 $Y2=0.755
r135 4 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.85
+ $Y=0.235 $X2=6.99 $Y2=0.445
r136 3 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.36
+ $Y=0.595 $X2=4.5 $Y2=0.805
r137 2 19 182 $w=1.7e-07 $l=3.39116e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.595 $X2=2.82 $Y2=0.805
r138 1 15 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=0.92
+ $Y=0.595 $X2=1.06 $Y2=0.755
.ends

