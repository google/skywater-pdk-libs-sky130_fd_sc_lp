* File: sky130_fd_sc_lp__o22ai_m.spice
* Created: Wed Sep  2 10:21:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22ai_m.pex.spice"
.subckt sky130_fd_sc_lp__o22ai_m  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_85_82#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1449 PD=0.7 PS=1.53 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.3
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_85_82#_M1006_d N_B2_M1006_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_85_82#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.0756 PD=0.72 PS=0.78 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_85_82#_M1003_d N_A1_M1003_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.063 PD=1.37 PS=0.72 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 A_198_535# N_B1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g A_198_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1007 A_356_535# N_A2_M1007_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g A_356_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
c_32 VNB 0 1.54761e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o22ai_m.pxi.spice"
*
.ends
*
*
