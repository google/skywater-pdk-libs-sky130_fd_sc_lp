* File: sky130_fd_sc_lp__dlygate4s15_1.pxi.spice
* Created: Wed Sep  2 09:49:58 2020
* 
x_PM_SKY130_FD_SC_LP__DLYGATE4S15_1%A N_A_M1005_g N_A_M1004_g N_A_c_69_n
+ N_A_c_74_n A A N_A_c_71_n PM_SKY130_FD_SC_LP__DLYGATE4S15_1%A
x_PM_SKY130_FD_SC_LP__DLYGATE4S15_1%A_27_52# N_A_27_52#_M1005_s
+ N_A_27_52#_M1004_s N_A_27_52#_c_103_n N_A_27_52#_M1002_g N_A_27_52#_M1000_g
+ N_A_27_52#_c_105_n N_A_27_52#_c_111_n N_A_27_52#_c_112_n N_A_27_52#_c_113_n
+ N_A_27_52#_c_106_n N_A_27_52#_c_107_n N_A_27_52#_c_114_n N_A_27_52#_c_108_n
+ N_A_27_52#_c_115_n PM_SKY130_FD_SC_LP__DLYGATE4S15_1%A_27_52#
x_PM_SKY130_FD_SC_LP__DLYGATE4S15_1%A_288_52# N_A_288_52#_M1002_d
+ N_A_288_52#_M1000_d N_A_288_52#_M1006_g N_A_288_52#_M1007_g
+ N_A_288_52#_c_162_n N_A_288_52#_c_163_n N_A_288_52#_c_164_n
+ N_A_288_52#_c_165_n N_A_288_52#_c_166_n N_A_288_52#_c_171_n
+ N_A_288_52#_c_172_n N_A_288_52#_c_167_n
+ PM_SKY130_FD_SC_LP__DLYGATE4S15_1%A_288_52#
x_PM_SKY130_FD_SC_LP__DLYGATE4S15_1%A_405_136# N_A_405_136#_M1006_s
+ N_A_405_136#_M1007_s N_A_405_136#_M1001_g N_A_405_136#_M1003_g
+ N_A_405_136#_c_222_n N_A_405_136#_c_227_n N_A_405_136#_c_223_n
+ N_A_405_136#_c_228_n N_A_405_136#_c_224_n N_A_405_136#_c_229_n
+ N_A_405_136#_c_225_n PM_SKY130_FD_SC_LP__DLYGATE4S15_1%A_405_136#
x_PM_SKY130_FD_SC_LP__DLYGATE4S15_1%VPWR N_VPWR_M1004_d N_VPWR_M1007_d
+ N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_288_n VPWR
+ N_VPWR_c_289_n N_VPWR_c_290_n N_VPWR_c_284_n N_VPWR_c_292_n
+ PM_SKY130_FD_SC_LP__DLYGATE4S15_1%VPWR
x_PM_SKY130_FD_SC_LP__DLYGATE4S15_1%X N_X_M1001_d N_X_M1003_d X X X X X X X
+ N_X_c_317_n X X N_X_c_321_n PM_SKY130_FD_SC_LP__DLYGATE4S15_1%X
x_PM_SKY130_FD_SC_LP__DLYGATE4S15_1%VGND N_VGND_M1005_d N_VGND_M1006_d
+ N_VGND_c_338_n N_VGND_c_339_n N_VGND_c_340_n N_VGND_c_341_n VGND
+ N_VGND_c_342_n N_VGND_c_343_n N_VGND_c_344_n N_VGND_c_345_n
+ PM_SKY130_FD_SC_LP__DLYGATE4S15_1%VGND
cc_1 VNB N_A_M1005_g 0.0567674f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.47
cc_2 VNB N_A_c_69_n 0.0239894f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.695
cc_3 VNB A 0.0252844f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A_c_71_n 0.0183476f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_5 VNB N_A_27_52#_c_103_n 0.0471722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_52#_M1002_g 0.0343363f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.695
cc_7 VNB N_A_27_52#_c_105_n 0.0205357f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_8 VNB N_A_27_52#_c_106_n 0.0195126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_52#_c_107_n 0.0120797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_52#_c_108_n 0.0345386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_288_52#_M1006_g 0.0321707f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_12 VNB N_A_288_52#_c_162_n 0.0246818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_288_52#_c_163_n 0.0177778f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_14 VNB N_A_288_52#_c_164_n 0.0225004f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.355
cc_15 VNB N_A_288_52#_c_165_n 0.0251362f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.665
cc_16 VNB N_A_288_52#_c_166_n 0.0105713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_288_52#_c_167_n 0.00394989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_405_136#_M1001_g 0.0283569f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_19 VNB N_A_405_136#_M1003_g 0.00154623f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB N_A_405_136#_c_222_n 0.00473003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_405_136#_c_223_n 0.00359467f $X=-0.19 $Y=-0.245 $X2=0.565
+ $Y2=1.355
cc_22 VNB N_A_405_136#_c_224_n 0.00807403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_405_136#_c_225_n 0.0357919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_284_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB X 0.0283845f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_26 VNB N_X_c_317_n 0.0329417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.014713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_338_n 0.00648778f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_29 VNB N_VGND_c_339_n 0.0170107f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_VGND_c_340_n 0.0569179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_341_n 0.00532387f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.355
cc_32 VNB N_VGND_c_342_n 0.0179296f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.295
cc_33 VNB N_VGND_c_343_n 0.0191738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_344_n 0.256015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_345_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_A_M1004_g 0.0539905f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.545
cc_37 VPB N_A_c_69_n 0.00312906f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.695
cc_38 VPB N_A_c_74_n 0.0183476f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.86
cc_39 VPB A 0.0136529f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_40 VPB N_A_27_52#_c_103_n 0.00226073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_27_52#_M1000_g 0.0449968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_27_52#_c_111_n 0.0220524f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.355
cc_43 VPB N_A_27_52#_c_112_n 0.0293341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_27_52#_c_113_n 0.0109405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_27_52#_c_114_n 0.00128612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_27_52#_c_115_n 0.0338046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_288_52#_M1007_g 0.0301174f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_48 VPB N_A_288_52#_c_162_n 0.0066533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_288_52#_c_165_n 0.00952145f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.665
cc_50 VPB N_A_288_52#_c_171_n 0.0125296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_288_52#_c_172_n 0.0183511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_405_136#_M1003_g 0.0272364f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_53 VPB N_A_405_136#_c_227_n 0.00392555f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_54 VPB N_A_405_136#_c_228_n 0.00216151f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.295
cc_55 VPB N_A_405_136#_c_229_n 0.00724414f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_285_n 0.0278295f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_57 VPB N_VPWR_c_286_n 0.0319012f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_58 VPB N_VPWR_c_287_n 0.059762f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_59 VPB N_VPWR_c_288_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_60 VPB N_VPWR_c_289_n 0.0188373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_290_n 0.0190092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_284_n 0.120263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_292_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB X 0.00847673f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.355
cc_65 VPB X 0.0492827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_X_c_321_n 0.0147363f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 A N_A_27_52#_c_103_n 0.00257472f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A_c_71_n N_A_27_52#_c_103_n 0.0211578f $X=0.565 $Y=1.355 $X2=0 $Y2=0
cc_69 N_A_M1005_g N_A_27_52#_c_105_n 0.013604f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_70 N_A_M1004_g N_A_27_52#_c_111_n 0.00631563f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_A_27_52#_c_112_n 0.0152432f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_72 N_A_c_74_n N_A_27_52#_c_112_n 0.00124917f $X=0.565 $Y=1.86 $X2=0 $Y2=0
cc_73 A N_A_27_52#_c_112_n 0.0257186f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_M1004_g N_A_27_52#_c_113_n 0.00349519f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_75 A N_A_27_52#_c_113_n 0.0280303f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_M1005_g N_A_27_52#_c_106_n 0.0117266f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_77 A N_A_27_52#_c_106_n 0.0251942f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A_c_71_n N_A_27_52#_c_106_n 0.00126146f $X=0.565 $Y=1.355 $X2=0 $Y2=0
cc_79 N_A_M1005_g N_A_27_52#_c_107_n 0.00435937f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_80 A N_A_27_52#_c_107_n 0.028939f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_M1005_g N_A_27_52#_c_114_n 9.13906e-19 $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_82 N_A_M1004_g N_A_27_52#_c_114_n 0.0031951f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_83 A N_A_27_52#_c_114_n 0.0394078f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_84 N_A_c_71_n N_A_27_52#_c_114_n 0.00220877f $X=0.565 $Y=1.355 $X2=0 $Y2=0
cc_85 N_A_M1005_g N_A_27_52#_c_108_n 0.00890898f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_A_27_52#_c_115_n 0.00247485f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_87 N_A_c_69_n N_A_27_52#_c_115_n 0.0211578f $X=0.565 $Y=1.695 $X2=0 $Y2=0
cc_88 N_A_M1004_g N_VPWR_c_285_n 0.00595698f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_89 N_A_M1004_g N_VPWR_c_289_n 0.00442668f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_90 N_A_M1004_g N_VPWR_c_284_n 0.0048347f $X=0.475 $Y=2.545 $X2=0 $Y2=0
cc_91 N_A_M1005_g N_VGND_c_338_n 0.00508082f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_92 N_A_M1005_g N_VGND_c_342_n 0.00547602f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_93 N_A_M1005_g N_VGND_c_344_n 0.00791561f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_94 N_A_27_52#_c_103_n N_A_288_52#_c_162_n 0.00405527f $X=1.19 $Y=1.68 $X2=0
+ $Y2=0
cc_95 N_A_27_52#_M1002_g N_A_288_52#_c_163_n 0.0211634f $X=1.365 $Y=0.47 $X2=0
+ $Y2=0
cc_96 N_A_27_52#_c_106_n N_A_288_52#_c_163_n 0.01637f $X=0.975 $Y=0.92 $X2=0
+ $Y2=0
cc_97 N_A_27_52#_c_114_n N_A_288_52#_c_163_n 0.0280969f $X=1.14 $Y=1.085 $X2=0
+ $Y2=0
cc_98 N_A_27_52#_M1002_g N_A_288_52#_c_166_n 0.00758366f $X=1.365 $Y=0.47 $X2=0
+ $Y2=0
cc_99 N_A_27_52#_M1000_g N_A_288_52#_c_171_n 0.00781162f $X=1.365 $Y=2.545 $X2=0
+ $Y2=0
cc_100 N_A_27_52#_c_103_n N_A_288_52#_c_172_n 0.0198174f $X=1.19 $Y=1.68 $X2=0
+ $Y2=0
cc_101 N_A_27_52#_c_112_n N_A_288_52#_c_172_n 0.0143606f $X=0.975 $Y=2.117 $X2=0
+ $Y2=0
cc_102 N_A_27_52#_c_114_n N_A_288_52#_c_172_n 0.0288323f $X=1.14 $Y=1.085 $X2=0
+ $Y2=0
cc_103 N_A_27_52#_c_103_n N_A_288_52#_c_167_n 0.00411974f $X=1.19 $Y=1.68 $X2=0
+ $Y2=0
cc_104 N_A_27_52#_c_114_n N_A_288_52#_c_167_n 0.0227663f $X=1.14 $Y=1.085 $X2=0
+ $Y2=0
cc_105 N_A_27_52#_M1000_g N_VPWR_c_285_n 0.0108947f $X=1.365 $Y=2.545 $X2=0
+ $Y2=0
cc_106 N_A_27_52#_c_112_n N_VPWR_c_285_n 0.0250261f $X=0.975 $Y=2.117 $X2=0
+ $Y2=0
cc_107 N_A_27_52#_M1000_g N_VPWR_c_287_n 0.00426083f $X=1.365 $Y=2.545 $X2=0
+ $Y2=0
cc_108 N_A_27_52#_c_111_n N_VPWR_c_289_n 0.00572829f $X=0.26 $Y=2.56 $X2=0 $Y2=0
cc_109 N_A_27_52#_M1000_g N_VPWR_c_284_n 0.0048347f $X=1.365 $Y=2.545 $X2=0
+ $Y2=0
cc_110 N_A_27_52#_c_111_n N_VPWR_c_284_n 0.00940928f $X=0.26 $Y=2.56 $X2=0 $Y2=0
cc_111 N_A_27_52#_M1002_g N_VGND_c_338_n 0.0102701f $X=1.365 $Y=0.47 $X2=0 $Y2=0
cc_112 N_A_27_52#_c_106_n N_VGND_c_338_n 0.0255952f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_113 N_A_27_52#_M1002_g N_VGND_c_340_n 0.00526675f $X=1.365 $Y=0.47 $X2=0
+ $Y2=0
cc_114 N_A_27_52#_c_105_n N_VGND_c_342_n 0.0152237f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_115 N_A_27_52#_M1002_g N_VGND_c_344_n 0.0116684f $X=1.365 $Y=0.47 $X2=0 $Y2=0
cc_116 N_A_27_52#_c_105_n N_VGND_c_344_n 0.0118277f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_117 N_A_27_52#_c_106_n N_VGND_c_344_n 0.0216353f $X=0.975 $Y=0.92 $X2=0 $Y2=0
cc_118 N_A_288_52#_M1006_g N_A_405_136#_M1001_g 0.00712749f $X=2.365 $Y=0.89
+ $X2=0 $Y2=0
cc_119 N_A_288_52#_M1007_g N_A_405_136#_M1003_g 0.00716311f $X=2.365 $Y=2.045
+ $X2=0 $Y2=0
cc_120 N_A_288_52#_c_165_n N_A_405_136#_M1003_g 0.00170317f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_121 N_A_288_52#_M1006_g N_A_405_136#_c_222_n 0.0107484f $X=2.365 $Y=0.89
+ $X2=0 $Y2=0
cc_122 N_A_288_52#_c_164_n N_A_405_136#_c_222_n 0.0288449f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_123 N_A_288_52#_c_165_n N_A_405_136#_c_222_n 0.00844207f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_124 N_A_288_52#_M1007_g N_A_405_136#_c_227_n 0.0106675f $X=2.365 $Y=2.045
+ $X2=0 $Y2=0
cc_125 N_A_288_52#_c_164_n N_A_405_136#_c_227_n 0.0288455f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_126 N_A_288_52#_c_165_n N_A_405_136#_c_227_n 0.00824234f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_127 N_A_288_52#_M1006_g N_A_405_136#_c_223_n 0.00237499f $X=2.365 $Y=0.89
+ $X2=0 $Y2=0
cc_128 N_A_288_52#_c_164_n N_A_405_136#_c_223_n 0.0203279f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_129 N_A_288_52#_c_165_n N_A_405_136#_c_223_n 0.00272912f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_130 N_A_288_52#_M1007_g N_A_405_136#_c_228_n 0.0026795f $X=2.365 $Y=2.045
+ $X2=0 $Y2=0
cc_131 N_A_288_52#_c_164_n N_A_405_136#_c_228_n 0.00234001f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_132 N_A_288_52#_c_165_n N_A_405_136#_c_228_n 8.04366e-19 $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_133 N_A_288_52#_M1006_g N_A_405_136#_c_224_n 0.0173794f $X=2.365 $Y=0.89
+ $X2=0 $Y2=0
cc_134 N_A_288_52#_c_162_n N_A_405_136#_c_224_n 0.00532229f $X=2.255 $Y=1.51
+ $X2=0 $Y2=0
cc_135 N_A_288_52#_c_163_n N_A_405_136#_c_224_n 0.0304038f $X=1.597 $Y=1.385
+ $X2=0 $Y2=0
cc_136 N_A_288_52#_c_164_n N_A_405_136#_c_224_n 0.0291548f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_137 N_A_288_52#_M1007_g N_A_405_136#_c_229_n 0.0129818f $X=2.365 $Y=2.045
+ $X2=0 $Y2=0
cc_138 N_A_288_52#_c_162_n N_A_405_136#_c_229_n 0.00514979f $X=2.255 $Y=1.51
+ $X2=0 $Y2=0
cc_139 N_A_288_52#_c_164_n N_A_405_136#_c_229_n 0.0284046f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_140 N_A_288_52#_c_172_n N_A_405_136#_c_229_n 0.021975f $X=1.567 $Y=2.395
+ $X2=0 $Y2=0
cc_141 N_A_288_52#_M1006_g N_A_405_136#_c_225_n 7.71641e-19 $X=2.365 $Y=0.89
+ $X2=0 $Y2=0
cc_142 N_A_288_52#_c_164_n N_A_405_136#_c_225_n 2.28029e-19 $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_143 N_A_288_52#_c_165_n N_A_405_136#_c_225_n 0.0184236f $X=2.575 $Y=1.51
+ $X2=0 $Y2=0
cc_144 N_A_288_52#_c_171_n N_VPWR_c_285_n 0.0107593f $X=1.58 $Y=2.56 $X2=0 $Y2=0
cc_145 N_A_288_52#_M1007_g N_VPWR_c_286_n 0.00431362f $X=2.365 $Y=2.045 $X2=0
+ $Y2=0
cc_146 N_A_288_52#_c_171_n N_VPWR_c_287_n 0.0056234f $X=1.58 $Y=2.56 $X2=0 $Y2=0
cc_147 N_A_288_52#_c_171_n N_VPWR_c_284_n 0.00929046f $X=1.58 $Y=2.56 $X2=0
+ $Y2=0
cc_148 N_A_288_52#_c_166_n N_VGND_c_338_n 0.0109344f $X=1.58 $Y=0.47 $X2=0 $Y2=0
cc_149 N_A_288_52#_M1006_g N_VGND_c_339_n 0.00486675f $X=2.365 $Y=0.89 $X2=0
+ $Y2=0
cc_150 N_A_288_52#_M1006_g N_VGND_c_340_n 0.00357582f $X=2.365 $Y=0.89 $X2=0
+ $Y2=0
cc_151 N_A_288_52#_c_166_n N_VGND_c_340_n 0.0145253f $X=1.58 $Y=0.47 $X2=0 $Y2=0
cc_152 N_A_288_52#_M1006_g N_VGND_c_344_n 0.00454494f $X=2.365 $Y=0.89 $X2=0
+ $Y2=0
cc_153 N_A_288_52#_c_166_n N_VGND_c_344_n 0.0113149f $X=1.58 $Y=0.47 $X2=0 $Y2=0
cc_154 N_A_405_136#_c_227_n N_VPWR_M1007_d 0.0181369f $X=2.91 $Y=1.91 $X2=0
+ $Y2=0
cc_155 N_A_405_136#_M1003_g N_VPWR_c_286_n 0.016516f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_405_136#_c_227_n N_VPWR_c_286_n 0.0234833f $X=2.91 $Y=1.91 $X2=0
+ $Y2=0
cc_157 N_A_405_136#_c_229_n N_VPWR_c_286_n 8.73769e-19 $X=2.165 $Y=1.91 $X2=0
+ $Y2=0
cc_158 N_A_405_136#_c_225_n N_VPWR_c_286_n 3.8937e-19 $X=3.165 $Y=1.46 $X2=0
+ $Y2=0
cc_159 N_A_405_136#_M1003_g N_VPWR_c_290_n 0.00486043f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_405_136#_M1003_g N_VPWR_c_284_n 0.00930006f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_405_136#_M1001_g X 0.00260428f $X=3.205 $Y=0.68 $X2=0 $Y2=0
cc_162 N_A_405_136#_M1003_g X 0.00292053f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_405_136#_c_223_n X 0.0327253f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_164 N_A_405_136#_c_228_n X 0.00710015f $X=3.032 $Y=1.825 $X2=0 $Y2=0
cc_165 N_A_405_136#_c_225_n X 0.00794767f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_166 N_A_405_136#_M1001_g N_X_c_317_n 0.00337221f $X=3.205 $Y=0.68 $X2=0 $Y2=0
cc_167 N_A_405_136#_c_223_n X 0.00398111f $X=3.032 $Y=1.625 $X2=0 $Y2=0
cc_168 N_A_405_136#_M1003_g N_X_c_321_n 0.00335846f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_405_136#_c_227_n N_X_c_321_n 0.00755038f $X=2.91 $Y=1.91 $X2=0 $Y2=0
cc_170 N_A_405_136#_c_228_n N_X_c_321_n 7.53353e-19 $X=3.032 $Y=1.825 $X2=0
+ $Y2=0
cc_171 N_A_405_136#_c_222_n N_VGND_M1006_d 0.0142993f $X=2.91 $Y=1.13 $X2=0
+ $Y2=0
cc_172 N_A_405_136#_c_223_n N_VGND_M1006_d 0.00192557f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_173 N_A_405_136#_M1001_g N_VGND_c_339_n 0.012902f $X=3.205 $Y=0.68 $X2=0
+ $Y2=0
cc_174 N_A_405_136#_c_222_n N_VGND_c_339_n 0.00679764f $X=2.91 $Y=1.13 $X2=0
+ $Y2=0
cc_175 N_A_405_136#_c_223_n N_VGND_c_339_n 0.0166857f $X=3.032 $Y=1.625 $X2=0
+ $Y2=0
cc_176 N_A_405_136#_c_224_n N_VGND_c_339_n 0.00576687f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_177 N_A_405_136#_c_225_n N_VGND_c_339_n 4.81801e-19 $X=3.165 $Y=1.46 $X2=0
+ $Y2=0
cc_178 N_A_405_136#_c_224_n N_VGND_c_340_n 0.00527907f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_179 N_A_405_136#_M1001_g N_VGND_c_343_n 0.00465098f $X=3.205 $Y=0.68 $X2=0
+ $Y2=0
cc_180 N_A_405_136#_M1001_g N_VGND_c_344_n 0.0091589f $X=3.205 $Y=0.68 $X2=0
+ $Y2=0
cc_181 N_A_405_136#_c_224_n N_VGND_c_344_n 0.0100519f $X=2.15 $Y=0.875 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_284_n N_X_M1003_d 0.00371702f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_290_n X 0.0289225f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_284_n X 0.0160565f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_185 N_X_c_317_n N_VGND_c_339_n 0.0234362f $X=3.42 $Y=0.42 $X2=0 $Y2=0
cc_186 N_X_c_317_n N_VGND_c_343_n 0.0296066f $X=3.42 $Y=0.42 $X2=0 $Y2=0
cc_187 N_X_c_317_n N_VGND_c_344_n 0.0160565f $X=3.42 $Y=0.42 $X2=0 $Y2=0
