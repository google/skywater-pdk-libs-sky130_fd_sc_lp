* File: sky130_fd_sc_lp__a22oi_m.pex.spice
* Created: Fri Aug 28 09:55:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22OI_M%B2 2 5 9 14 17 20 22 23 24 25 26 33
r37 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.085 $X2=0.27 $Y2=1.085
r38 25 26 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r39 24 25 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r40 23 24 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r41 23 34 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.085
r42 22 34 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.085
r43 18 20 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.36 $Y=1.825
+ $X2=0.635 $Y2=1.825
r44 16 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.425
+ $X2=0.27 $Y2=1.085
r45 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.425
+ $X2=0.27 $Y2=1.59
r46 12 33 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.07
+ $X2=0.27 $Y2=1.085
r47 12 14 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.27 $Y=0.995
+ $X2=0.59 $Y2=0.995
r48 7 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.635 $Y=1.9
+ $X2=0.635 $Y2=1.825
r49 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.635 $Y=1.9 $X2=0.635
+ $Y2=2.69
r50 3 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.59 $Y=0.92 $X2=0.59
+ $Y2=0.995
r51 3 5 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=0.59 $Y=0.92 $X2=0.59
+ $Y2=0.445
r52 2 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=1.75 $X2=0.36
+ $Y2=1.825
r53 2 17 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.36 $Y=1.75 $X2=0.36
+ $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_M%B1 3 6 9 11 12 13 14 15 21
c39 9 0 1.72493e-19 $X=1.065 $Y=2.69
r40 21 23 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.042 $Y=1.005
+ $X2=1.042 $Y2=0.84
r41 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.045
+ $Y=1.005 $X2=1.045 $Y2=1.005
r42 14 15 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.122 $Y=1.665
+ $X2=1.122 $Y2=2.035
r43 13 14 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.122 $Y=1.295
+ $X2=1.122 $Y2=1.665
r44 13 22 10.2833 $w=3.23e-07 $l=2.9e-07 $layer=LI1_cond $X=1.122 $Y=1.295
+ $X2=1.122 $Y2=1.005
r45 12 22 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=1.122 $Y=0.925
+ $X2=1.122 $Y2=1.005
r46 9 11 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.065 $Y=2.69
+ $X2=1.065 $Y2=1.51
r47 6 11 38.9802 $w=3.35e-07 $l=1.67e-07 $layer=POLY_cond $X=1.042 $Y=1.343
+ $X2=1.042 $Y2=1.51
r48 5 21 0.344503 $w=3.35e-07 $l=2e-09 $layer=POLY_cond $X=1.042 $Y=1.007
+ $X2=1.042 $Y2=1.005
r49 5 6 57.8765 $w=3.35e-07 $l=3.36e-07 $layer=POLY_cond $X=1.042 $Y=1.007
+ $X2=1.042 $Y2=1.343
r50 3 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.95 $Y=0.445
+ $X2=0.95 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_M%A1 3 6 9 11 12 13 14 15 16 23
c45 9 0 2.51603e-19 $X=1.495 $Y=2.69
r46 23 25 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.587 $Y=1.475
+ $X2=1.587 $Y2=1.31
r47 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.59
+ $Y=1.475 $X2=1.59 $Y2=1.475
r48 15 16 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.635 $Y=1.665
+ $X2=1.635 $Y2=2.035
r49 15 24 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=1.635 $Y=1.665
+ $X2=1.635 $Y2=1.475
r50 14 24 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=1.635 $Y=1.295
+ $X2=1.635 $Y2=1.475
r51 13 14 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.635 $Y=0.925
+ $X2=1.635 $Y2=1.295
r52 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.635 $Y=0.555
+ $X2=1.635 $Y2=0.925
r53 9 11 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.495 $Y=2.69
+ $X2=1.495 $Y2=1.98
r54 6 11 46.5995 $w=3.35e-07 $l=1.67e-07 $layer=POLY_cond $X=1.587 $Y=1.813
+ $X2=1.587 $Y2=1.98
r55 5 23 0.344503 $w=3.35e-07 $l=2e-09 $layer=POLY_cond $X=1.587 $Y=1.477
+ $X2=1.587 $Y2=1.475
r56 5 6 57.8765 $w=3.35e-07 $l=3.36e-07 $layer=POLY_cond $X=1.587 $Y=1.477
+ $X2=1.587 $Y2=1.813
r57 3 25 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=1.495 $Y=0.445
+ $X2=1.495 $Y2=1.31
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_M%A2 3 5 7 9 13 17 20 21 22 23 24 30
c35 21 0 1.29722e-19 $X=2.16 $Y=0.925
r36 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.13
+ $Y=1.085 $X2=2.13 $Y2=1.085
r37 23 24 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.145 $Y=1.665
+ $X2=2.145 $Y2=2.035
r38 22 23 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.145 $Y=1.295
+ $X2=2.145 $Y2=1.665
r39 22 31 11.6455 $w=1.98e-07 $l=2.1e-07 $layer=LI1_cond $X=2.145 $Y=1.295
+ $X2=2.145 $Y2=1.085
r40 21 31 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.145 $Y=0.925
+ $X2=2.145 $Y2=1.085
r41 19 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.13 $Y=1.425
+ $X2=2.13 $Y2=1.085
r42 19 20 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.425
+ $X2=2.13 $Y2=1.59
r43 15 17 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.925 $Y=2.295
+ $X2=2.07 $Y2=2.295
r44 13 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.13 $Y=1.07
+ $X2=2.13 $Y2=1.085
r45 10 13 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=1.855 $Y=0.995
+ $X2=2.13 $Y2=0.995
r46 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.07 $Y=2.22 $X2=2.07
+ $Y2=2.295
r47 9 20 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.07 $Y=2.22 $X2=2.07
+ $Y2=1.59
r48 5 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=2.37
+ $X2=1.925 $Y2=2.295
r49 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.925 $Y=2.37
+ $X2=1.925 $Y2=2.69
r50 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.855 $Y=0.92
+ $X2=1.855 $Y2=0.995
r51 1 3 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.855 $Y=0.92
+ $X2=1.855 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_M%A_39_496# 1 2 3 10 16 17 20 23
r31 23 25 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.34 $Y=2.775 $X2=0.34
+ $Y2=2.975
r32 18 20 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=2.15 $Y=2.49
+ $X2=2.15 $Y2=2.625
r33 16 18 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.055 $Y=2.405
+ $X2=2.15 $Y2=2.49
r34 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.055 $Y=2.405
+ $X2=1.365 $Y2=2.405
r35 13 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.28 $Y=2.89
+ $X2=1.28 $Y2=2.605
r36 12 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.28 $Y=2.49
+ $X2=1.365 $Y2=2.405
r37 12 15 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.28 $Y=2.49
+ $X2=1.28 $Y2=2.605
r38 11 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.505 $Y=2.975
+ $X2=0.34 $Y2=2.975
r39 10 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.195 $Y=2.975
+ $X2=1.28 $Y2=2.89
r40 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.195 $Y=2.975
+ $X2=0.505 $Y2=2.975
r41 3 20 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2 $Y=2.48
+ $X2=2.14 $Y2=2.625
r42 2 15 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=2.48 $X2=1.28 $Y2=2.605
r43 1 23 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=2.48 $X2=0.34 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_M%Y 1 2 7 9 12
c29 12 0 1.21881e-19 $X=0.72 $Y=2.405
r30 12 21 4.54441 $w=3.49e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=2.515
+ $X2=0.85 $Y2=2.515
r31 12 17 0.873926 $w=3.49e-07 $l=2.5e-08 $layer=LI1_cond $X=0.72 $Y=2.515
+ $X2=0.695 $Y2=2.515
r32 12 17 4.95691 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.695 $Y=2.32
+ $X2=0.695 $Y2=2.515
r33 11 12 62.0593 $w=3.13e-07 $l=1.66e-06 $layer=LI1_cond $X=0.695 $Y=0.66
+ $X2=0.695 $Y2=2.32
r34 7 11 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=0.495
+ $X2=0.695 $Y2=0.66
r35 7 9 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.78 $Y=0.495
+ $X2=1.165 $Y2=0.495
r36 2 21 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=2.48 $X2=0.85 $Y2=2.605
r37 1 9 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.165 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_M%VPWR 1 6 8 10 20 21 24
c25 6 0 1.72493e-19 $X=1.71 $Y=2.775
r26 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r28 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.71 $Y2=3.33
r30 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 12 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.71 $Y2=3.33
r34 10 16 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r35 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r36 8 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.24
+ $Y2=3.33
r37 8 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=3.245 $X2=1.71
+ $Y2=3.33
r39 4 6 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.71 $Y=3.245 $X2=1.71
+ $Y2=2.775
r40 1 6 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=2.48 $X2=1.71 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_M%VGND 1 2 7 9 11 13 15 17 30
r33 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r36 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r37 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r38 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r39 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 18 26 3.50342 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r41 18 20 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r42 17 29 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.172
+ $Y2=0
r43 17 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.68
+ $Y2=0
r44 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r45 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r46 11 29 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.172 $Y2=0
r47 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.38
r48 7 26 3.34047 $w=1.9e-07 $l=1.56844e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.215 $Y2=0
r49 7 9 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.38
r50 2 13 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.235 $X2=2.11 $Y2=0.38
r51 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.22
+ $Y=0.235 $X2=0.345 $Y2=0.38
.ends

