* File: sky130_fd_sc_lp__o2111a_lp.pex.spice
* Created: Fri Aug 28 11:00:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111A_LP%A1 3 7 10 11 12 15 16
r31 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.505
+ $Y=1.39 $X2=0.505 $Y2=1.39
r32 12 16 4.73076 $w=6.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.24 $Y=1.56
+ $X2=0.505 $Y2=1.56
r33 10 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.505 $Y=1.73
+ $X2=0.505 $Y2=1.39
r34 10 11 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.73
+ $X2=0.505 $Y2=1.895
r35 5 15 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.225
+ $X2=0.505 $Y2=1.39
r36 5 7 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.505 $Y=1.225
+ $X2=0.505 $Y2=0.465
r37 3 11 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.545 $Y=2.595
+ $X2=0.545 $Y2=1.895
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_LP%A2 3 7 11 12 13 16
r38 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.075
+ $Y=1.39 $X2=1.075 $Y2=1.39
r39 13 17 2.23149 $w=6.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=1.56
+ $X2=1.075 $Y2=1.56
r40 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.075 $Y=1.73
+ $X2=1.075 $Y2=1.39
r41 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.73
+ $X2=1.075 $Y2=1.895
r42 10 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.225
+ $X2=1.075 $Y2=1.39
r43 7 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.015 $Y=0.465
+ $X2=1.015 $Y2=1.225
r44 3 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.035 $Y=2.595
+ $X2=1.035 $Y2=1.895
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_LP%B1 3 7 9 10 11 12 18
c44 3 0 1.93746e-19 $X=1.555 $Y=0.465
r45 18 21 32.0725 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.652 $Y=1.73
+ $X2=1.652 $Y2=1.895
r46 18 20 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.652 $Y=1.73
+ $X2=1.652 $Y2=1.565
r47 12 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=1.73 $X2=1.66 $Y2=1.73
r48 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=1.295
+ $X2=1.66 $Y2=1.665
r49 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=0.925
+ $X2=1.66 $Y2=1.295
r50 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=0.555
+ $X2=1.66 $Y2=0.925
r51 7 21 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.605 $Y=2.595
+ $X2=1.605 $Y2=1.895
r52 3 20 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=1.555 $Y=0.465
+ $X2=1.555 $Y2=1.565
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_LP%C1 3 6 9 12 13 16 17
c53 17 0 3.84897e-20 $X=2.23 $Y=1.77
r54 16 18 31.3435 $w=5.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.322 $Y=1.77
+ $X2=2.322 $Y2=1.935
r55 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.77 $X2=2.23 $Y2=1.77
r56 13 17 8.72564 $w=3.48e-07 $l=2.65e-07 $layer=LI1_cond $X=2.22 $Y=2.035
+ $X2=2.22 $Y2=1.77
r57 11 12 45.4127 $w=5.15e-07 $l=1.5e-07 $layer=POLY_cond $X=2.225 $Y=1.175
+ $X2=2.225 $Y2=1.325
r58 9 18 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.455 $Y=2.595
+ $X2=2.455 $Y2=1.935
r59 6 16 9.55781 $w=5.15e-07 $l=9.2e-08 $layer=POLY_cond $X=2.322 $Y=1.678
+ $X2=2.322 $Y2=1.77
r60 6 12 36.6729 $w=5.15e-07 $l=3.53e-07 $layer=POLY_cond $X=2.322 $Y=1.678
+ $X2=2.322 $Y2=1.325
r61 3 11 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.945 $Y=0.465
+ $X2=1.945 $Y2=1.175
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_LP%D1 1 3 4 5 8 10 11 14
c51 5 0 3.84897e-20 $X=2.41 $Y=0.84
r52 17 19 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.985 $Y=0.93
+ $X2=2.985 $Y2=1.095
r53 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.985
+ $Y=0.93 $X2=2.985 $Y2=0.93
r54 14 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.985 $Y=0.84
+ $X2=2.985 $Y2=0.93
r55 11 18 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=3.12 $Y=0.925
+ $X2=2.985 $Y2=0.925
r56 10 18 12.4248 $w=3.18e-07 $l=3.45e-07 $layer=LI1_cond $X=2.64 $Y=0.925
+ $X2=2.985 $Y2=0.925
r57 8 19 372.68 $w=2.5e-07 $l=1.5e-06 $layer=POLY_cond $X=3.005 $Y=2.595
+ $X2=3.005 $Y2=1.095
r58 4 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.82 $Y=0.84
+ $X2=2.985 $Y2=0.84
r59 4 5 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.82 $Y=0.84 $X2=2.41
+ $Y2=0.84
r60 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.335 $Y=0.765
+ $X2=2.41 $Y2=0.84
r61 1 3 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.335 $Y=0.765 $X2=2.335
+ $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_LP%A_232_419# 1 2 3 12 16 20 24 26 29 32 33
+ 35 37 38 40 44 47 51 52 55 57 58 59
c120 38 0 1.33735e-19 $X=2.345 $Y=1.35
c121 32 0 6.00116e-20 $X=2.26 $Y=1.265
r122 55 57 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.34 $Y=2.24
+ $X2=1.34 $Y2=2.415
r123 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.58
+ $Y=1.38 $X2=3.58 $Y2=1.38
r124 49 51 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.58 $Y=1.715
+ $X2=3.58 $Y2=1.38
r125 48 58 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=1.8
+ $X2=2.74 $Y2=1.8
r126 47 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.415 $Y=1.8
+ $X2=3.58 $Y2=1.715
r127 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.415 $Y=1.8
+ $X2=2.905 $Y2=1.8
r128 42 59 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=2.33
+ $X2=2.74 $Y2=2.415
r129 42 44 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.74 $Y=2.33 $X2=2.74
+ $Y2=2.24
r130 41 58 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=1.885
+ $X2=2.74 $Y2=1.8
r131 41 44 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.74 $Y=1.885
+ $X2=2.74 $Y2=2.24
r132 40 58 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.66 $Y=1.715
+ $X2=2.74 $Y2=1.8
r133 39 40 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.66 $Y=1.435
+ $X2=2.66 $Y2=1.715
r134 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=1.35
+ $X2=2.66 $Y2=1.435
r135 37 38 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.575 $Y=1.35
+ $X2=2.345 $Y2=1.35
r136 33 35 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.345 $Y=0.45
+ $X2=2.55 $Y2=0.45
r137 32 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.26 $Y=1.265
+ $X2=2.345 $Y2=1.35
r138 31 33 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.26 $Y=0.585
+ $X2=2.345 $Y2=0.45
r139 31 32 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.26 $Y=0.585
+ $X2=2.26 $Y2=1.265
r140 30 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=2.415
+ $X2=1.34 $Y2=2.415
r141 29 59 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=2.415
+ $X2=2.74 $Y2=2.415
r142 29 30 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=2.575 $Y=2.415
+ $X2=1.505 $Y2=2.415
r143 25 52 53.3155 $w=3.55e-07 $l=3.28e-07 $layer=POLY_cond $X=3.567 $Y=1.708
+ $X2=3.567 $Y2=1.38
r144 25 26 32.478 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=3.567 $Y=1.708
+ $X2=3.567 $Y2=1.885
r145 24 52 2.43821 $w=3.55e-07 $l=1.5e-08 $layer=POLY_cond $X=3.567 $Y=1.365
+ $X2=3.567 $Y2=1.38
r146 16 26 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.535 $Y=2.595
+ $X2=3.535 $Y2=1.885
r147 10 24 25.9344 $w=3.55e-07 $l=1.5e-07 $layer=POLY_cond $X=3.645 $Y=1.215
+ $X2=3.645 $Y2=1.365
r148 10 20 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.825 $Y=1.215
+ $X2=3.825 $Y2=0.445
r149 10 12 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.465 $Y=1.215
+ $X2=3.465 $Y2=0.445
r150 3 44 300 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=2.095 $X2=2.74 $Y2=2.24
r151 2 55 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=1.16
+ $Y=2.095 $X2=1.34 $Y2=2.24
r152 1 35 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.41
+ $Y=0.255 $X2=2.55 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_LP%VPWR 1 2 3 10 12 18 22 27 28 29 38 44 45
+ 51
r54 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 45 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 42 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=3.33
+ $X2=3.27 $Y2=3.33
r59 42 44 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.435 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=3.27 $Y2=3.33
r61 38 40 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 34 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r65 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r66 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 31 48 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r68 31 33 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 29 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 29 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 27 36 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.87 $Y2=3.33
r74 26 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.87 $Y2=3.33
r76 22 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.27 $Y=2.24 $X2=3.27
+ $Y2=2.95
r77 20 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=3.245
+ $X2=3.27 $Y2=3.33
r78 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.27 $Y=3.245
+ $X2=3.27 $Y2=2.95
r79 16 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=3.33
r80 16 18 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=2.895
r81 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.24 $X2=0.28
+ $Y2=2.95
r82 10 48 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r83 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.95
r84 3 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.095 $X2=3.27 $Y2=2.95
r85 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.095 $X2=3.27 $Y2=2.24
r86 2 18 600 $w=1.7e-07 $l=8.67179e-07 $layer=licon1_PDIFF $count=1 $X=1.73
+ $Y=2.095 $X2=1.87 $Y2=2.895
r87 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.95
r88 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_LP%X 1 2 7 8 9 10 11 12 13 33 36
r26 34 36 0.944272 $w=5.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.92 $Y=2.36
+ $X2=3.92 $Y2=2.405
r27 33 47 1.92074 $w=2.38e-07 $l=4e-08 $layer=LI1_cond $X=4.085 $Y=2.035
+ $X2=4.085 $Y2=2.075
r28 12 34 0.419677 $w=5.68e-07 $l=2e-08 $layer=LI1_cond $X=3.92 $Y=2.34 $X2=3.92
+ $Y2=2.36
r29 12 49 2.09838 $w=5.68e-07 $l=1e-07 $layer=LI1_cond $X=3.92 $Y=2.34 $X2=3.92
+ $Y2=2.24
r30 12 13 7.34434 $w=5.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.92 $Y=2.425
+ $X2=3.92 $Y2=2.775
r31 12 36 0.419677 $w=5.68e-07 $l=2e-08 $layer=LI1_cond $X=3.92 $Y=2.425
+ $X2=3.92 $Y2=2.405
r32 11 49 3.00069 $w=5.68e-07 $l=1.43e-07 $layer=LI1_cond $X=3.92 $Y=2.097
+ $X2=3.92 $Y2=2.24
r33 11 47 4.56511 $w=5.68e-07 $l=2.2e-08 $layer=LI1_cond $X=3.92 $Y=2.097
+ $X2=3.92 $Y2=2.075
r34 11 33 1.10442 $w=2.38e-07 $l=2.3e-08 $layer=LI1_cond $X=4.085 $Y=2.012
+ $X2=4.085 $Y2=2.035
r35 10 11 16.6624 $w=2.38e-07 $l=3.47e-07 $layer=LI1_cond $X=4.085 $Y=1.665
+ $X2=4.085 $Y2=2.012
r36 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.085 $Y=1.295
+ $X2=4.085 $Y2=1.665
r37 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.085 $Y=0.925
+ $X2=4.085 $Y2=1.295
r38 8 45 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=4.085 $Y=0.925
+ $X2=4.085 $Y2=0.675
r39 7 45 8.03684 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.04 $Y=0.47
+ $X2=4.04 $Y2=0.675
r40 2 49 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.66
+ $Y=2.095 $X2=3.8 $Y2=2.24
r41 1 7 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_LP%A_29_51# 1 2 9 11 12 15
r26 13 15 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=1.19 $Y=0.875
+ $X2=1.19 $Y2=0.48
r27 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.065 $Y=0.96
+ $X2=1.19 $Y2=0.875
r28 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.065 $Y=0.96
+ $X2=0.375 $Y2=0.96
r29 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.25 $Y=0.875
+ $X2=0.375 $Y2=0.96
r30 7 9 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=0.25 $Y=0.875
+ $X2=0.25 $Y2=0.48
r31 2 15 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.255 $X2=1.23 $Y2=0.48
r32 1 9 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.255 $X2=0.29 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r51 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r52 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r54 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r55 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.25
+ $Y2=0
r56 27 29 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=4.08
+ $Y2=0
r57 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r58 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.72
+ $Y2=0
r60 23 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.2
+ $Y2=0
r61 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.25
+ $Y2=0
r62 22 25 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=3.085 $Y=0 $X2=1.2
+ $Y2=0
r63 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r64 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.72
+ $Y2=0
r66 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.24
+ $Y2=0
r67 15 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r68 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r69 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0
r70 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0.4
r71 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085 $X2=0.72
+ $Y2=0
r72 7 9 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.72 $Y=0.085 $X2=0.72
+ $Y2=0.465
r73 2 13 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=3.105
+ $Y=0.235 $X2=3.25 $Y2=0.4
r74 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.58
+ $Y=0.255 $X2=0.72 $Y2=0.465
.ends

