* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o22a_0 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_80_313# B2 a_286_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR B1 a_372_489# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 VGND A1 a_286_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_536_489# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_286_125# B1 a_80_313# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_80_313# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_80_313# A2 a_536_489# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_372_489# B2 a_80_313# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 X a_80_313# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_286_125# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
