* File: sky130_fd_sc_lp__dlrtp_4.spice
* Created: Wed Sep  2 09:47:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrtp_4.pex.spice"
.subckt sky130_fd_sc_lp__dlrtp_4  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_D_M1001_g N_A_49_70#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.1113 PD=0.97 PS=1.37 NRD=77.136 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1025 N_A_267_464#_M1025_d N_GATE_M1025_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1155 PD=1.37 PS=0.97 NRD=0 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_267_464#_M1002_g N_A_414_47#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.1113 PD=0.78 PS=1.37 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1012 A_599_47# N_A_49_70#_M1012_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0756 PD=0.63 PS=0.78 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_671_47#_M1009_d N_A_414_47#_M1009_g A_599_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1017 A_779_47# N_A_267_464#_M1017_g N_A_671_47#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_857_21#_M1024_g A_779_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 A_1083_73# N_A_671_47#_M1013_g N_A_857_21#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1512 AS=0.2226 PD=1.2 PS=2.21 NRD=17.856 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1021 N_VGND_M1021_d N_RESET_B_M1021_g A_1083_73# VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=17.856 M=1 R=5.6 SA=75000.7
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1003 N_Q_M1003_d N_A_857_21#_M1003_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1005 N_Q_M1003_d N_A_857_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1011 N_Q_M1011_d N_A_857_21#_M1011_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1019 N_Q_M1011_d N_A_857_21#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_D_M1006_g N_A_49_70#_M1006_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.168 AS=0.1696 PD=1.165 PS=1.81 NRD=3.0732 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1022 N_A_267_464#_M1022_d N_GATE_M1022_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1856 AS=0.168 PD=1.86 PS=1.165 NRD=7.683 NRS=72.3187 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_267_464#_M1000_g N_A_414_47#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1984 AS=0.1696 PD=1.26 PS=1.81 NRD=93.8705 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75004 A=0.096 P=1.58 MULT=1
MM1004 A_651_469# N_A_49_70#_M1004_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1984 PD=0.85 PS=1.26 NRD=15.3857 NRS=10.7562 M=1 R=4.26667
+ SA=75001 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1020 N_A_671_47#_M1020_d N_A_267_464#_M1020_g A_651_469# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.130294 AS=0.0672 PD=1.22566 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.3 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1016 A_828_469# N_A_414_47#_M1016_g N_A_671_47#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.04725 AS=0.0855057 PD=0.645 PS=0.80434 NRD=26.9693 NRS=44.5417 M=1
+ R=2.8 SA=75001.8 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_857_21#_M1010_g A_828_469# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1344 AS=0.04725 PD=1.005 PS=0.645 NRD=222.787 NRS=26.9693 M=1 R=2.8
+ SA=75002.2 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1014 N_A_857_21#_M1014_d N_A_671_47#_M1014_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.4032 PD=1.54 PS=3.015 NRD=0 NRS=0 M=1 R=8.4 SA=75001.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_RESET_B_M1007_g N_A_857_21#_M1014_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.22365 AS=0.1764 PD=1.615 PS=1.54 NRD=4.6886 NRS=0 M=1 R=8.4
+ SA=75001.6 SB=75002 A=0.189 P=2.82 MULT=1
MM1008 N_Q_M1008_d N_A_857_21#_M1008_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.22365 PD=1.54 PS=1.615 NRD=0 NRS=7.0329 M=1 R=8.4 SA=75002.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1015 N_Q_M1008_d N_A_857_21#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1018 N_Q_M1018_d N_A_857_21#_M1018_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1023 N_Q_M1018_d N_A_857_21#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=15.9271 P=20.81
c_103 VNB 0 1.59482e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dlrtp_4.pxi.spice"
*
.ends
*
*
