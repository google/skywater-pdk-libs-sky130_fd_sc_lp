* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor3_lp A B C VGND VNB VPB VPWR X
X0 a_763_347# a_647_367# a_27_109# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1860_132# a_1348_111# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_265_409# B a_763_347# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_265_409# B a_803_81# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_1318_85# C a_1634_89# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1634_89# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_763_347# a_647_367# a_265_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_1348_111# C a_803_81# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VGND a_1348_111# a_1860_132# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_27_109# B a_803_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_803_81# a_1318_85# a_1348_111# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_27_109# a_265_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_114_109# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR a_1348_111# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VPWR B a_647_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_27_109# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_27_109# A a_114_109# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_272_109# a_27_109# a_265_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_570_101# B a_647_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1348_111# C a_763_347# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_803_81# a_647_367# a_265_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_763_347# a_1318_85# a_1348_111# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_27_109# B a_763_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X23 a_1318_85# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X24 VGND a_27_109# a_272_109# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND B a_570_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_803_81# a_647_367# a_27_109# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
