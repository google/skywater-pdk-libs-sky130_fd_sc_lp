* File: sky130_fd_sc_lp__dlxbp_1.spice
* Created: Wed Sep  2 09:48:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxbp_1.pex.spice"
.subckt sky130_fd_sc_lp__dlxbp_1  VNB VPB D GATE VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_D_M1021_g N_A_46_62#_M1021_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1020 N_A_215_62#_M1020_d N_GATE_M1020_g N_VGND_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_215_62#_M1013_g N_A_367_491#_M1013_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0777 AS=0.1113 PD=0.79 PS=1.37 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1007 A_568_47# N_A_46_62#_M1007_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0777 PD=0.63 PS=0.79 NRD=14.28 NRS=12.852 M=1 R=2.8 SA=75000.7
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1003 N_A_608_491#_M1003_d N_A_367_491#_M1003_g A_568_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1015 A_748_47# N_A_215_62#_M1015_g N_A_608_491#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=17.136 M=1 R=2.8
+ SA=75001.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_758_359#_M1001_g A_748_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0938 AS=0.0441 PD=0.83 PS=0.63 NRD=18.564 NRS=14.28 M=1 R=2.8 SA=75002
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1018 N_A_758_359#_M1018_d N_A_608_491#_M1018_g N_VGND_M1001_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2394 AS=0.1876 PD=2.25 PS=1.66 NRD=2.856 NRS=8.928 M=1
+ R=5.6 SA=75001.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_758_359#_M1004_g N_Q_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1792 AS=0.2226 PD=1.62 PS=2.21 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.5 A=0.126 P=1.98 MULT=1
MM1016 N_A_1266_147#_M1016_d N_A_758_359#_M1016_g N_VGND_M1004_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0896 PD=1.37 PS=0.81 NRD=0 NRS=15.708 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_Q_N_M1014_d N_A_1266_147#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_D_M1002_g N_A_46_62#_M1002_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_215_62#_M1008_d N_GATE_M1008_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1010_d N_A_215_62#_M1010_g N_A_367_491#_M1010_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1005 A_536_491# N_A_46_62#_M1005_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1019 N_A_608_491#_M1019_d N_A_215_62#_M1019_g A_536_491# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.130294 AS=0.0672 PD=1.22566 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1011 A_713_491# N_A_367_491#_M1011_g N_A_608_491#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.04725 AS=0.0855057 PD=0.645 PS=0.80434 NRD=26.9693 NRS=46.886 M=1
+ R=2.8 SA=75001.5 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_758_359#_M1006_g A_713_491# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.135975 AS=0.04725 PD=1.0125 PS=0.645 NRD=229.82 NRS=26.9693 M=1 R=2.8
+ SA=75001.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_A_758_359#_M1009_d N_A_608_491#_M1009_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.407925 PD=3.05 PS=3.0375 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_A_758_359#_M1017_g N_Q_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.268115 AS=0.3339 PD=2.16853 PS=3.05 NRD=2.6004 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.5 A=0.189 P=2.82 MULT=1
MM1012 N_A_1266_147#_M1012_d N_A_758_359#_M1012_g N_VPWR_M1017_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.136185 PD=1.81 PS=1.10147 NRD=0 NRS=22.3004 M=1
+ R=4.26667 SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_Q_N_M1000_d N_A_1266_147#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.1159 P=19.97
c_150 VPB 0 9.24665e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlxbp_1.pxi.spice"
*
.ends
*
*
