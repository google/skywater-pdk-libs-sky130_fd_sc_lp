* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or3_lp A B C VGND VNB VPB VPWR X
X0 a_454_57# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND C a_612_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_108_31# a_138_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND A a_296_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_541_409# C a_108_31# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VPWR A a_443_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_612_57# C a_108_31# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_443_409# B a_541_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_296_57# A a_108_31# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_108_31# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_108_31# B a_454_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_138_57# a_108_31# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
