* File: sky130_fd_sc_lp__nand2_m.pex.spice
* Created: Fri Aug 28 10:47:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2_M%B 2 5 9 11 12 13 14 15 21
r32 21 23 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.005
+ $X2=0.402 $Y2=0.84
r33 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.35
+ $Y=1.005 $X2=0.35 $Y2=1.005
r34 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.295 $Y=1.665
+ $X2=0.295 $Y2=2.035
r35 13 14 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.295 $Y=1.295
+ $X2=0.295 $Y2=1.665
r36 13 22 11.936 $w=2.78e-07 $l=2.9e-07 $layer=LI1_cond $X=0.295 $Y=1.295
+ $X2=0.295 $Y2=1.005
r37 12 22 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=0.295 $Y=0.925
+ $X2=0.295 $Y2=1.005
r38 9 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.545 $Y=0.445
+ $X2=0.545 $Y2=0.84
r39 5 11 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.505 $Y=2.52
+ $X2=0.505 $Y2=1.51
r40 2 11 47.7177 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=0.402 $Y=1.293
+ $X2=0.402 $Y2=1.51
r41 1 21 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=0.402 $Y=1.057
+ $X2=0.402 $Y2=1.005
r42 1 2 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=0.402 $Y=1.057
+ $X2=0.402 $Y2=1.293
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_M%A 3 6 9 11 12 13 14 15 21
r26 21 23 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.047 $Y=1.005
+ $X2=1.047 $Y2=0.84
r27 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.07
+ $Y=1.005 $X2=1.07 $Y2=1.005
r28 14 15 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=1.665
+ $X2=1.135 $Y2=2.035
r29 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=1.295
+ $X2=1.135 $Y2=1.665
r30 13 22 11.1403 $w=2.98e-07 $l=2.9e-07 $layer=LI1_cond $X=1.135 $Y=1.295
+ $X2=1.135 $Y2=1.005
r31 12 22 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=1.135 $Y=0.925
+ $X2=1.135 $Y2=1.005
r32 9 11 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.935 $Y=2.52
+ $X2=0.935 $Y2=1.51
r33 6 11 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=1.047 $Y=1.323
+ $X2=1.047 $Y2=1.51
r34 5 21 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=1.047 $Y=1.027
+ $X2=1.047 $Y2=1.005
r35 5 6 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=1.047 $Y=1.027
+ $X2=1.047 $Y2=1.323
r36 3 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.935 $Y=0.445
+ $X2=0.935 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_M%VPWR 1 2 7 9 11 13 15 17 27
r19 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r20 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r21 18 23 3.64151 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.197 $Y2=3.33
r22 18 20 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.72 $Y2=3.33
r23 17 26 3.64249 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=1.242 $Y2=3.33
r24 17 20 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r26 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 11 26 3.2727 $w=2.1e-07 $l=1.27609e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.242 $Y2=3.33
r29 11 13 38.026 $w=2.08e-07 $l=7.2e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=2.525
r30 7 23 3.27368 $w=2.1e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.197 $Y2=3.33
r31 7 9 38.026 $w=2.08e-07 $l=7.2e-07 $layer=LI1_cond $X=0.29 $Y=3.245 $X2=0.29
+ $Y2=2.525
r32 2 13 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=2.31 $X2=1.15 $Y2=2.525
r33 1 9 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.31 $X2=0.29 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_M%Y 1 2 7 8 9 10 11 12 13 22 40
r25 13 34 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=0.71 $Y=2.775
+ $X2=0.71 $Y2=2.525
r26 12 34 7.00478 $w=1.88e-07 $l=1.2e-07 $layer=LI1_cond $X=0.71 $Y=2.405
+ $X2=0.71 $Y2=2.525
r27 11 12 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=2.035
+ $X2=0.71 $Y2=2.405
r28 10 11 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=1.665
+ $X2=0.71 $Y2=2.035
r29 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=1.295
+ $X2=0.71 $Y2=1.665
r30 8 9 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=0.925 $X2=0.71
+ $Y2=1.295
r31 8 22 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=0.71 $Y=0.925
+ $X2=0.71 $Y2=0.66
r32 7 22 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=0.495
+ $X2=0.71 $Y2=0.66
r33 7 40 9.63663 $w=4.98e-07 $l=3.45e-07 $layer=LI1_cond $X=0.805 $Y=0.495
+ $X2=1.15 $Y2=0.495
r34 2 34 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=2.31 $X2=0.72 $Y2=2.525
r35 1 40 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.235 $X2=1.15 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_M%VGND 1 4 6 8 12 13
r20 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r21 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r22 10 16 3.62383 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r23 10 12 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=1.2
+ $Y2=0
r24 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r25 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r26 4 16 3.29137 $w=2.1e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.217 $Y2=0
r27 4 6 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.33 $Y2=0.38
r28 1 6 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.235 $X2=0.33 $Y2=0.38
.ends

