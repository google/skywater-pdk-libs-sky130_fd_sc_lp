* File: sky130_fd_sc_lp__o2111ai_1.pxi.spice
* Created: Fri Aug 28 11:00:55 2020
* 
x_PM_SKY130_FD_SC_LP__O2111AI_1%D1 N_D1_M1002_g N_D1_M1009_g D1 D1 N_D1_c_55_n
+ N_D1_c_56_n PM_SKY130_FD_SC_LP__O2111AI_1%D1
x_PM_SKY130_FD_SC_LP__O2111AI_1%C1 N_C1_M1003_g N_C1_M1005_g C1 C1 C1
+ N_C1_c_84_n N_C1_c_85_n PM_SKY130_FD_SC_LP__O2111AI_1%C1
x_PM_SKY130_FD_SC_LP__O2111AI_1%B1 N_B1_M1007_g N_B1_M1006_g B1 N_B1_c_119_n
+ N_B1_c_120_n PM_SKY130_FD_SC_LP__O2111AI_1%B1
x_PM_SKY130_FD_SC_LP__O2111AI_1%A2 N_A2_M1001_g N_A2_M1000_g A2 A2 N_A2_c_152_n
+ PM_SKY130_FD_SC_LP__O2111AI_1%A2
x_PM_SKY130_FD_SC_LP__O2111AI_1%A1 N_A1_M1008_g N_A1_M1004_g A1 N_A1_c_183_n
+ N_A1_c_184_n PM_SKY130_FD_SC_LP__O2111AI_1%A1
x_PM_SKY130_FD_SC_LP__O2111AI_1%VPWR N_VPWR_M1009_s N_VPWR_M1005_d
+ N_VPWR_M1004_d N_VPWR_c_206_n N_VPWR_c_207_n N_VPWR_c_208_n N_VPWR_c_209_n
+ N_VPWR_c_210_n N_VPWR_c_211_n VPWR N_VPWR_c_212_n N_VPWR_c_213_n
+ N_VPWR_c_214_n N_VPWR_c_205_n PM_SKY130_FD_SC_LP__O2111AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O2111AI_1%Y N_Y_M1002_s N_Y_M1009_d N_Y_M1006_d
+ N_Y_c_246_n N_Y_c_249_n N_Y_c_250_n N_Y_c_266_n N_Y_c_274_n N_Y_c_283_n
+ N_Y_c_247_n Y Y Y Y PM_SKY130_FD_SC_LP__O2111AI_1%Y
x_PM_SKY130_FD_SC_LP__O2111AI_1%A_361_47# N_A_361_47#_M1007_d
+ N_A_361_47#_M1008_d N_A_361_47#_c_312_p N_A_361_47#_c_294_n
+ N_A_361_47#_c_295_n N_A_361_47#_c_296_n
+ PM_SKY130_FD_SC_LP__O2111AI_1%A_361_47#
x_PM_SKY130_FD_SC_LP__O2111AI_1%VGND N_VGND_M1001_d N_VGND_c_318_n VGND
+ N_VGND_c_319_n N_VGND_c_320_n N_VGND_c_321_n N_VGND_c_322_n
+ PM_SKY130_FD_SC_LP__O2111AI_1%VGND
cc_1 VNB N_D1_M1009_g 0.00883768f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=2.465
cc_2 VNB D1 0.00237101f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_3 VNB N_D1_c_55_n 0.0368578f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_4 VNB N_D1_c_56_n 0.0203263f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.185
cc_5 VNB N_C1_M1005_g 0.0076702f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=2.465
cc_6 VNB C1 0.00593f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_7 VNB N_C1_c_84_n 0.0328343f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.185
cc_8 VNB N_C1_c_85_n 0.0157478f $X=-0.19 $Y=-0.245 $X2=0.747 $Y2=0.925
cc_9 VNB N_B1_M1007_g 0.026784f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=0.655
cc_10 VNB N_B1_c_119_n 0.00892103f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.185
cc_11 VNB N_B1_c_120_n 0.0246601f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.515
cc_12 VNB N_A2_M1001_g 0.0278022f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=0.655
cc_13 VNB A2 0.00645726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_152_n 0.0235062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_M1008_g 0.0305761f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=0.655
cc_16 VNB N_A1_M1004_g 0.00176076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_183_n 0.0557027f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_18 VNB N_A1_c_184_n 0.00111806f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.185
cc_19 VNB N_VPWR_c_205_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_246_n 0.0485875f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_21 VNB N_Y_c_247_n 0.0178017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_361_47#_c_294_n 0.0139876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_361_47#_c_295_n 0.00703825f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.35
cc_24 VNB N_A_361_47#_c_296_n 0.0292785f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.185
cc_25 VNB N_VGND_c_318_n 0.00557321f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=2.465
cc_26 VNB N_VGND_c_319_n 0.0667536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_320_n 0.0189813f $X=-0.19 $Y=-0.245 $X2=0.747 $Y2=1.295
cc_28 VNB N_VGND_c_321_n 0.191001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_322_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_D1_M1009_g 0.0241095f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=2.465
cc_31 VPB N_C1_M1005_g 0.0219367f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=2.465
cc_32 VPB N_B1_M1006_g 0.0214782f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_B1_c_119_n 0.00361801f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.185
cc_34 VPB N_B1_c_120_n 0.0065661f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.515
cc_35 VPB N_A2_M1000_g 0.0189326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB A2 0.0123408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A2_c_152_n 0.00716719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A1_M1004_g 0.0245277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A1_c_184_n 0.00674287f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.185
cc_40 VPB N_VPWR_c_206_n 0.0429753f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.35
cc_41 VPB N_VPWR_c_207_n 0.00561626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_208_n 0.0113538f $X=-0.19 $Y=1.655 $X2=0.747 $Y2=1.295
cc_43 VPB N_VPWR_c_209_n 0.0481497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_210_n 0.0158267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_211_n 0.00549311f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_212_n 0.0180322f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_213_n 0.0304898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_214_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_205_n 0.0589629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_Y_c_246_n 0.00176411f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.35
cc_51 VPB N_Y_c_249_n 0.0151126f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.35
cc_52 VPB N_Y_c_250_n 0.0258084f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.185
cc_53 N_D1_M1009_g N_C1_M1005_g 0.0176165f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_54 D1 C1 0.0520683f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_55 N_D1_c_56_n C1 0.00826145f $X=0.73 $Y=1.185 $X2=0 $Y2=0
cc_56 D1 N_C1_c_84_n 3.54126e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_57 N_D1_c_55_n N_C1_c_84_n 0.0206581f $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_58 D1 N_C1_c_85_n 3.40042e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_59 N_D1_c_56_n N_C1_c_85_n 0.0437987f $X=0.73 $Y=1.185 $X2=0 $Y2=0
cc_60 N_D1_M1009_g N_VPWR_c_206_n 0.0169041f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_61 N_D1_M1009_g N_VPWR_c_212_n 0.00486043f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_62 N_D1_M1009_g N_VPWR_c_205_n 0.00851476f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_63 D1 N_Y_M1002_s 0.00349333f $X=0.635 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_64 N_D1_M1009_g N_Y_c_246_n 0.00537056f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_65 D1 N_Y_c_246_n 0.0534037f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_66 N_D1_c_55_n N_Y_c_246_n 0.0081237f $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_67 N_D1_c_56_n N_Y_c_246_n 0.00486224f $X=0.73 $Y=1.185 $X2=0 $Y2=0
cc_68 N_D1_M1009_g N_Y_c_249_n 0.0192218f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_69 D1 N_Y_c_249_n 0.0218533f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_70 N_D1_c_55_n N_Y_c_249_n 0.00322512f $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_71 D1 N_Y_c_247_n 0.00927291f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_72 N_D1_c_55_n N_Y_c_247_n 0.00206326f $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_73 N_D1_c_56_n N_Y_c_247_n 0.00793105f $X=0.73 $Y=1.185 $X2=0 $Y2=0
cc_74 N_D1_c_56_n N_VGND_c_319_n 0.00547467f $X=0.73 $Y=1.185 $X2=0 $Y2=0
cc_75 D1 N_VGND_c_321_n 0.00359928f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_76 N_D1_c_56_n N_VGND_c_321_n 0.00842204f $X=0.73 $Y=1.185 $X2=0 $Y2=0
cc_77 C1 N_B1_M1007_g 0.00389578f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_78 N_C1_c_84_n N_B1_M1007_g 0.0151227f $X=1.28 $Y=1.35 $X2=0 $Y2=0
cc_79 N_C1_c_85_n N_B1_M1007_g 0.0411969f $X=1.28 $Y=1.185 $X2=0 $Y2=0
cc_80 N_C1_M1005_g N_B1_M1006_g 0.0380601f $X=1.37 $Y=2.465 $X2=0 $Y2=0
cc_81 C1 N_B1_c_119_n 0.0135149f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_82 N_C1_c_84_n N_B1_c_119_n 0.00615108f $X=1.28 $Y=1.35 $X2=0 $Y2=0
cc_83 N_C1_M1005_g N_B1_c_120_n 0.0151227f $X=1.37 $Y=2.465 $X2=0 $Y2=0
cc_84 N_C1_M1005_g N_VPWR_c_206_n 0.00114941f $X=1.37 $Y=2.465 $X2=0 $Y2=0
cc_85 N_C1_M1005_g N_VPWR_c_207_n 0.00810561f $X=1.37 $Y=2.465 $X2=0 $Y2=0
cc_86 N_C1_M1005_g N_VPWR_c_212_n 0.00585385f $X=1.37 $Y=2.465 $X2=0 $Y2=0
cc_87 N_C1_M1005_g N_VPWR_c_205_n 0.0112749f $X=1.37 $Y=2.465 $X2=0 $Y2=0
cc_88 C1 N_Y_c_246_n 0.00515484f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_89 N_C1_M1005_g N_Y_c_249_n 0.0129737f $X=1.37 $Y=2.465 $X2=0 $Y2=0
cc_90 C1 N_Y_c_249_n 0.027172f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_91 N_C1_c_84_n N_Y_c_249_n 0.00141163f $X=1.28 $Y=1.35 $X2=0 $Y2=0
cc_92 N_C1_M1005_g N_Y_c_266_n 0.0114241f $X=1.37 $Y=2.465 $X2=0 $Y2=0
cc_93 C1 N_Y_c_247_n 0.0163343f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_94 N_C1_c_85_n N_Y_c_247_n 8.51421e-19 $X=1.28 $Y=1.185 $X2=0 $Y2=0
cc_95 C1 A_181_47# 0.00844828f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_96 C1 N_A_361_47#_c_295_n 0.00424545f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_97 C1 N_VGND_c_319_n 0.0102788f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_98 N_C1_c_85_n N_VGND_c_319_n 0.00382445f $X=1.28 $Y=1.185 $X2=0 $Y2=0
cc_99 C1 N_VGND_c_321_n 0.0104349f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_100 N_C1_c_85_n N_VGND_c_321_n 0.00566996f $X=1.28 $Y=1.185 $X2=0 $Y2=0
cc_101 N_B1_M1007_g N_A2_M1001_g 0.0306531f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_102 N_B1_M1006_g N_A2_M1000_g 0.0348873f $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_103 N_B1_c_119_n A2 0.0349758f $X=1.82 $Y=1.51 $X2=0 $Y2=0
cc_104 N_B1_c_120_n A2 0.0031801f $X=1.92 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B1_c_119_n N_A2_c_152_n 2.77051e-19 $X=1.82 $Y=1.51 $X2=0 $Y2=0
cc_106 N_B1_c_120_n N_A2_c_152_n 0.0204734f $X=1.92 $Y=1.51 $X2=0 $Y2=0
cc_107 N_B1_M1006_g N_VPWR_c_207_n 0.00810561f $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_108 N_B1_M1006_g N_VPWR_c_213_n 0.00585385f $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_109 N_B1_M1006_g N_VPWR_c_205_n 0.0114658f $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_110 N_B1_M1006_g N_Y_c_249_n 9.92087e-19 $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_111 N_B1_c_119_n N_Y_c_249_n 0.00608971f $X=1.82 $Y=1.51 $X2=0 $Y2=0
cc_112 N_B1_M1006_g N_Y_c_266_n 0.0186366f $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B1_c_119_n N_Y_c_266_n 0.0268906f $X=1.82 $Y=1.51 $X2=0 $Y2=0
cc_114 N_B1_c_120_n N_Y_c_266_n 9.54588e-19 $X=1.92 $Y=1.51 $X2=0 $Y2=0
cc_115 N_B1_M1007_g N_A_361_47#_c_295_n 0.00198729f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_116 N_B1_c_119_n N_A_361_47#_c_295_n 0.00550979f $X=1.82 $Y=1.51 $X2=0 $Y2=0
cc_117 N_B1_c_120_n N_A_361_47#_c_295_n 0.00490405f $X=1.92 $Y=1.51 $X2=0 $Y2=0
cc_118 N_B1_M1007_g N_VGND_c_319_n 0.00585385f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_119 N_B1_M1007_g N_VGND_c_321_n 0.0113938f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_120 N_A2_M1001_g N_A1_M1008_g 0.0306173f $X=2.28 $Y=0.655 $X2=0 $Y2=0
cc_121 N_A2_M1000_g N_A1_M1004_g 0.0563522f $X=2.49 $Y=2.465 $X2=0 $Y2=0
cc_122 A2 N_A1_c_183_n 0.00336663f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_123 N_A2_c_152_n N_A1_c_183_n 0.0563522f $X=2.49 $Y=1.51 $X2=0 $Y2=0
cc_124 A2 N_A1_c_184_n 0.0343638f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A2_c_152_n N_A1_c_184_n 3.0539e-19 $X=2.49 $Y=1.51 $X2=0 $Y2=0
cc_126 N_A2_M1000_g N_VPWR_c_209_n 0.00450323f $X=2.49 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A2_M1000_g N_VPWR_c_213_n 0.00585385f $X=2.49 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A2_M1000_g N_VPWR_c_205_n 0.0111635f $X=2.49 $Y=2.465 $X2=0 $Y2=0
cc_129 A2 N_Y_c_274_n 0.0252535f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A2_c_152_n N_Y_c_274_n 9.9155e-19 $X=2.49 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A2_M1001_g N_A_361_47#_c_294_n 0.0160427f $X=2.28 $Y=0.655 $X2=0 $Y2=0
cc_132 A2 N_A_361_47#_c_294_n 0.0434936f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A2_c_152_n N_A_361_47#_c_294_n 0.0052993f $X=2.49 $Y=1.51 $X2=0 $Y2=0
cc_134 A2 N_A_361_47#_c_295_n 0.00854387f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A2_M1001_g N_A_361_47#_c_296_n 0.00101994f $X=2.28 $Y=0.655 $X2=0 $Y2=0
cc_136 N_A2_M1001_g N_VGND_c_318_n 0.00662084f $X=2.28 $Y=0.655 $X2=0 $Y2=0
cc_137 N_A2_M1001_g N_VGND_c_319_n 0.00585385f $X=2.28 $Y=0.655 $X2=0 $Y2=0
cc_138 N_A2_M1001_g N_VGND_c_321_n 0.0114931f $X=2.28 $Y=0.655 $X2=0 $Y2=0
cc_139 N_A1_M1004_g N_VPWR_c_209_n 0.0297269f $X=2.85 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A1_c_183_n N_VPWR_c_209_n 0.00161609f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_141 N_A1_c_184_n N_VPWR_c_209_n 0.0259088f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_142 N_A1_M1004_g N_VPWR_c_213_n 0.00486043f $X=2.85 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A1_M1004_g N_VPWR_c_205_n 0.00818711f $X=2.85 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A1_M1008_g N_A_361_47#_c_294_n 0.0185653f $X=2.85 $Y=0.655 $X2=0 $Y2=0
cc_145 N_A1_c_183_n N_A_361_47#_c_294_n 0.00754271f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_146 N_A1_c_184_n N_A_361_47#_c_294_n 0.0277825f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_147 N_A1_M1008_g N_A_361_47#_c_296_n 0.0123544f $X=2.85 $Y=0.655 $X2=0 $Y2=0
cc_148 N_A1_M1008_g N_VGND_c_318_n 0.00662084f $X=2.85 $Y=0.655 $X2=0 $Y2=0
cc_149 N_A1_M1008_g N_VGND_c_320_n 0.0054895f $X=2.85 $Y=0.655 $X2=0 $Y2=0
cc_150 N_A1_M1008_g N_VGND_c_321_n 0.0111877f $X=2.85 $Y=0.655 $X2=0 $Y2=0
cc_151 N_VPWR_c_205_n N_Y_M1009_d 0.00504357f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_152 N_VPWR_c_205_n N_Y_M1006_d 0.00659813f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_153 N_VPWR_M1009_s N_Y_c_249_n 0.00265343f $X=0.49 $Y=1.835 $X2=0 $Y2=0
cc_154 N_VPWR_c_206_n N_Y_c_249_n 0.0234402f $X=0.615 $Y=2.18 $X2=0 $Y2=0
cc_155 N_VPWR_c_206_n N_Y_c_250_n 7.9643e-19 $X=0.615 $Y=2.18 $X2=0 $Y2=0
cc_156 N_VPWR_M1005_d N_Y_c_266_n 0.00712086f $X=1.445 $Y=1.835 $X2=0 $Y2=0
cc_157 N_VPWR_c_207_n N_Y_c_266_n 0.0232685f $X=1.645 $Y=2.435 $X2=0 $Y2=0
cc_158 N_VPWR_c_213_n N_Y_c_283_n 0.0222962f $X=2.9 $Y=3.33 $X2=0 $Y2=0
cc_159 N_VPWR_c_205_n N_Y_c_283_n 0.0127519f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_c_212_n Y 0.0214287f $X=1.48 $Y=3.33 $X2=0 $Y2=0
cc_161 N_VPWR_c_205_n Y 0.0129463f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_162 N_VPWR_c_205_n A_513_367# 0.00899413f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_163 N_Y_c_247_n N_VGND_c_319_n 0.0433241f $X=0.275 $Y=0.42 $X2=0 $Y2=0
cc_164 N_Y_M1002_s N_VGND_c_321_n 0.0050085f $X=0.15 $Y=0.235 $X2=0 $Y2=0
cc_165 N_Y_c_247_n N_VGND_c_321_n 0.0255934f $X=0.275 $Y=0.42 $X2=0 $Y2=0
cc_166 A_181_47# N_VGND_c_321_n 0.00766031f $X=0.905 $Y=0.235 $X2=0 $Y2=0
cc_167 A_269_47# N_VGND_c_321_n 0.0126264f $X=1.345 $Y=0.235 $X2=3.12 $Y2=0
cc_168 N_A_361_47#_c_294_n N_VGND_M1001_d 0.00371685f $X=2.9 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_361_47#_c_294_n N_VGND_c_318_n 0.0220556f $X=2.9 $Y=1.09 $X2=0 $Y2=0
cc_170 N_A_361_47#_c_312_p N_VGND_c_319_n 0.0215996f $X=2.005 $Y=0.42 $X2=0
+ $Y2=0
cc_171 N_A_361_47#_c_296_n N_VGND_c_320_n 0.0210467f $X=3.065 $Y=0.42 $X2=0
+ $Y2=0
cc_172 N_A_361_47#_M1007_d N_VGND_c_321_n 0.00573482f $X=1.805 $Y=0.235 $X2=0
+ $Y2=0
cc_173 N_A_361_47#_M1008_d N_VGND_c_321_n 0.00215158f $X=2.925 $Y=0.235 $X2=0
+ $Y2=0
cc_174 N_A_361_47#_c_312_p N_VGND_c_321_n 0.0127519f $X=2.005 $Y=0.42 $X2=0
+ $Y2=0
cc_175 N_A_361_47#_c_296_n N_VGND_c_321_n 0.0125689f $X=3.065 $Y=0.42 $X2=0
+ $Y2=0
