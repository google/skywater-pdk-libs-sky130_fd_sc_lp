* File: sky130_fd_sc_lp__a32oi_0.pex.spice
* Created: Fri Aug 28 10:01:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32OI_0%B2 3 7 11 13 14 15 16 21
c30 7 0 1.82199e-19 $X=0.63 $Y=0.445
c31 3 0 1.81942e-19 $X=0.525 $Y=2.305
r32 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.33
+ $Y=1.005 $X2=0.33 $Y2=1.005
r33 15 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.665
r34 15 22 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.005
r35 14 22 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=0.27 $Y=0.925 $X2=0.27
+ $Y2=1.005
r36 12 21 36.8212 $w=4.35e-07 $l=2.88e-07 $layer=POLY_cond $X=0.382 $Y=1.293
+ $X2=0.382 $Y2=1.005
r37 12 13 53.1843 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=0.382 $Y=1.293
+ $X2=0.382 $Y2=1.51
r38 11 21 1.91777 $w=4.35e-07 $l=1.5e-08 $layer=POLY_cond $X=0.382 $Y=0.99
+ $X2=0.382 $Y2=1.005
r39 10 11 44.6182 $w=4.35e-07 $l=1.5e-07 $layer=POLY_cond $X=0.435 $Y=0.84
+ $X2=0.435 $Y2=0.99
r40 7 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.63 $Y=0.445
+ $X2=0.63 $Y2=0.84
r41 3 13 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.525 $Y=2.305
+ $X2=0.525 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_0%B1 3 7 9 10 12 13 14 18
c38 13 0 1.82199e-19 $X=1.2 $Y=0.925
c39 3 0 1.81942e-19 $X=0.955 $Y=2.305
r40 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.11
+ $Y=0.94 $X2=1.11 $Y2=0.94
r41 14 19 12.2125 $w=3.33e-07 $l=3.55e-07 $layer=LI1_cond $X=1.192 $Y=1.295
+ $X2=1.192 $Y2=0.94
r42 13 19 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=1.192 $Y=0.925
+ $X2=1.192 $Y2=0.94
r43 12 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=0.775
+ $X2=1.11 $Y2=0.94
r44 9 18 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.11 $Y=1.295
+ $X2=1.11 $Y2=0.94
r45 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.077 $Y=1.295
+ $X2=1.077 $Y2=1.445
r46 7 12 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.02 $Y=0.445 $X2=1.02
+ $Y2=0.775
r47 3 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.955 $Y=2.305
+ $X2=0.955 $Y2=1.445
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_0%A1 3 7 9 12 15 16 17 18 19 20 25
c50 9 0 2.54468e-20 $X=1.59 $Y=1.685
r51 19 20 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.925
+ $X2=1.69 $Y2=1.295
r52 19 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=0.93 $X2=1.68 $Y2=0.93
r53 18 19 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.555
+ $X2=1.69 $Y2=0.925
r54 16 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.68 $Y=1.27
+ $X2=1.68 $Y2=0.93
r55 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.27
+ $X2=1.68 $Y2=1.435
r56 15 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=0.765
+ $X2=1.68 $Y2=0.93
r57 10 12 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=1.385 $Y=1.76
+ $X2=1.59 $Y2=1.76
r58 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.59 $Y=1.685
+ $X2=1.59 $Y2=1.76
r59 9 17 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.59 $Y=1.685
+ $X2=1.59 $Y2=1.435
r60 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.59 $Y=0.445
+ $X2=1.59 $Y2=0.765
r61 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.385 $Y=1.835
+ $X2=1.385 $Y2=1.76
r62 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.385 $Y=1.835 $X2=1.385
+ $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_0%A2 3 7 10 11 13 14 15 16 17 18 23
c50 23 0 2.64121e-20 $X=2.25 $Y=0.93
c51 16 0 1.1034e-19 $X=2.16 $Y=0.555
r52 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.25
+ $Y=0.93 $X2=2.25 $Y2=0.93
r53 18 24 10.6492 $w=3.93e-07 $l=3.65e-07 $layer=LI1_cond $X=2.217 $Y=1.295
+ $X2=2.217 $Y2=0.93
r54 17 24 0.145879 $w=3.93e-07 $l=5e-09 $layer=LI1_cond $X=2.217 $Y=0.925
+ $X2=2.217 $Y2=0.93
r55 16 17 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.217 $Y=0.555
+ $X2=2.217 $Y2=0.925
r56 14 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.25 $Y=1.27
+ $X2=2.25 $Y2=0.93
r57 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.27
+ $X2=2.25 $Y2=1.435
r58 13 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=0.765
+ $X2=2.25 $Y2=0.93
r59 10 11 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=2.157 $Y=1.675
+ $X2=2.157 $Y2=1.825
r60 10 15 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.16 $Y=1.675
+ $X2=2.16 $Y2=1.435
r61 7 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.16 $Y=0.445
+ $X2=2.16 $Y2=0.765
r62 3 11 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.155 $Y=2.305
+ $X2=2.155 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_0%A3 3 7 10 12 17 18 19 20 25
c35 17 0 8.48931e-20 $X=2.805 $Y=1.51
r36 25 27 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.005
+ $X2=2.805 $Y2=0.84
r37 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.82
+ $Y=1.005 $X2=2.82 $Y2=1.005
r38 19 20 7.19592 $w=6.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.967 $Y=1.295
+ $X2=2.967 $Y2=1.665
r39 19 26 5.64004 $w=6.13e-07 $l=2.9e-07 $layer=LI1_cond $X=2.967 $Y=1.295
+ $X2=2.967 $Y2=1.005
r40 18 26 1.55587 $w=6.13e-07 $l=8e-08 $layer=LI1_cond $X=2.967 $Y=0.925
+ $X2=2.967 $Y2=1.005
r41 12 13 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=2.715 $Y=1.75
+ $X2=2.585 $Y2=1.75
r42 12 17 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.675
+ $X2=2.715 $Y2=1.51
r43 10 17 43.2685 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=2.805 $Y=1.33
+ $X2=2.805 $Y2=1.51
r44 9 25 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=2.805 $Y=1.02
+ $X2=2.805 $Y2=1.005
r45 9 10 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=2.805 $Y=1.02
+ $X2=2.805 $Y2=1.33
r46 7 27 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.7 $Y=0.445 $X2=2.7
+ $Y2=0.84
r47 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.585 $Y=1.825
+ $X2=2.585 $Y2=1.75
r48 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.585 $Y=1.825
+ $X2=2.585 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_0%A_37_397# 1 2 3 12 14 15 19 20 21 24
r49 22 24 15.7579 $w=2.43e-07 $l=3.35e-07 $layer=LI1_cond $X=2.367 $Y=1.795
+ $X2=2.367 $Y2=2.13
r50 20 22 7.02594 $w=1.8e-07 $l=1.60823e-07 $layer=LI1_cond $X=2.245 $Y=1.705
+ $X2=2.367 $Y2=1.795
r51 20 21 58.2273 $w=1.78e-07 $l=9.45e-07 $layer=LI1_cond $X=2.245 $Y=1.705
+ $X2=1.3 $Y2=1.705
r52 17 19 28.7063 $w=2.73e-07 $l=6.85e-07 $layer=LI1_cond $X=1.162 $Y=2.815
+ $X2=1.162 $Y2=2.13
r53 16 21 7.21025 $w=1.8e-07 $l=1.77381e-07 $layer=LI1_cond $X=1.162 $Y=1.795
+ $X2=1.3 $Y2=1.705
r54 16 19 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=1.162 $Y=1.795
+ $X2=1.162 $Y2=2.13
r55 14 17 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=1.025 $Y=2.9
+ $X2=1.162 $Y2=2.815
r56 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.025 $Y=2.9
+ $X2=0.455 $Y2=2.9
r57 10 15 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.3 $Y=2.815
+ $X2=0.455 $Y2=2.9
r58 10 12 25.4653 $w=3.08e-07 $l=6.85e-07 $layer=LI1_cond $X=0.3 $Y=2.815
+ $X2=0.3 $Y2=2.13
r59 3 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.23
+ $Y=1.985 $X2=2.37 $Y2=2.13
r60 2 19 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=1.985 $X2=1.17 $Y2=2.13
r61 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=1.985 $X2=0.31 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_0%Y 1 2 9 11 12 13 14 15 16 24
r30 16 35 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.74 $Y=2.405
+ $X2=0.74 $Y2=2.13
r31 15 35 4.76009 $w=2.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.74 $Y=2.035
+ $X2=0.74 $Y2=2.13
r32 14 15 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=1.665
+ $X2=0.74 $Y2=2.035
r33 13 14 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=1.295
+ $X2=0.74 $Y2=1.665
r34 12 13 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=0.925
+ $X2=0.74 $Y2=1.295
r35 11 24 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.74 $Y=0.43
+ $X2=0.74 $Y2=0.595
r36 11 12 15.4327 $w=2.28e-07 $l=3.08e-07 $layer=LI1_cond $X=0.74 $Y=0.617
+ $X2=0.74 $Y2=0.925
r37 11 24 1.10234 $w=2.28e-07 $l=2.2e-08 $layer=LI1_cond $X=0.74 $Y=0.617
+ $X2=0.74 $Y2=0.595
r38 7 11 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=0.855 $Y=0.43
+ $X2=0.74 $Y2=0.43
r39 7 9 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.855 $Y=0.43
+ $X2=1.26 $Y2=0.43
r40 2 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.985 $X2=0.74 $Y2=2.13
r41 1 9 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.235 $X2=1.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_0%VPWR 1 2 9 13 16 17 18 20 33 34 37
c33 20 0 3.63885e-19 $X=1.47 $Y=3.33
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 28 37 12.6176 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=2.075 $Y=3.33
+ $X2=1.772 $Y2=3.33
r38 28 30 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.075 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 23 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 22 26 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 20 37 12.6176 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=1.47 $Y=3.33
+ $X2=1.772 $Y2=3.33
r44 20 26 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.47 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 18 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 18 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 16 30 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.66 $Y=3.33 $X2=2.64
+ $Y2=3.33
r49 16 17 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.66 $Y=3.33
+ $X2=2.812 $Y2=3.33
r50 15 33 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 15 17 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.812 $Y2=3.33
r52 11 17 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.812 $Y=3.245
+ $X2=2.812 $Y2=3.33
r53 11 13 42.1303 $w=3.03e-07 $l=1.115e-06 $layer=LI1_cond $X=2.812 $Y=3.245
+ $X2=2.812 $Y2=2.13
r54 7 37 2.53987 $w=6.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.772 $Y=3.245
+ $X2=1.772 $Y2=3.33
r55 7 9 22.0434 $w=6.03e-07 $l=1.115e-06 $layer=LI1_cond $X=1.772 $Y=3.245
+ $X2=1.772 $Y2=2.13
r56 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.66
+ $Y=1.985 $X2=2.8 $Y2=2.13
r57 1 9 150 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=4 $X=1.46
+ $Y=1.985 $X2=1.94 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_0%VGND 1 2 7 9 13 15 16 17 18 29
c44 29 0 2.64121e-20 $X=3.12 $Y=0
r45 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 26 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r48 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r49 23 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r50 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r51 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 20 31 3.6162 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r53 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r54 18 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r55 18 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r56 16 25 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.64
+ $Y2=0
r57 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.915
+ $Y2=0
r58 15 28 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.12
+ $Y2=0
r59 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.915
+ $Y2=0
r60 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0
r61 11 13 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.445
r62 7 31 3.29899 $w=2.1e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.35 $Y=0.085
+ $X2=0.227 $Y2=0
r63 7 9 19.013 $w=2.08e-07 $l=3.6e-07 $layer=LI1_cond $X=0.35 $Y=0.085 $X2=0.35
+ $Y2=0.445
r64 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.235 $X2=2.915 $Y2=0.445
r65 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.235 $X2=0.35 $Y2=0.445
.ends

