* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__iso0p_lp2 A SLEEP KAPWR VGND VNB VPB VPWR X
X0 KAPWR a_342_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VGND a_342_417# a_602_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_27_93# SLEEP KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_112_93# SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 KAPWR a_27_93# a_342_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_27_93# SLEEP a_112_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_27_93# a_340_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_340_93# A a_342_417# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_342_417# A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_602_93# a_342_417# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
