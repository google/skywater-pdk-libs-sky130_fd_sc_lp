* File: sky130_fd_sc_lp__or2_2.pxi.spice
* Created: Fri Aug 28 11:21:28 2020
* 
x_PM_SKY130_FD_SC_LP__OR2_2%B N_B_c_56_n N_B_M1004_g N_B_c_63_n N_B_M1000_g
+ N_B_c_58_n N_B_c_59_n N_B_c_64_n B B N_B_c_61_n PM_SKY130_FD_SC_LP__OR2_2%B
x_PM_SKY130_FD_SC_LP__OR2_2%A N_A_M1003_g N_A_M1006_g A N_A_c_99_n N_A_c_100_n
+ PM_SKY130_FD_SC_LP__OR2_2%A
x_PM_SKY130_FD_SC_LP__OR2_2%A_48_390# N_A_48_390#_M1004_d N_A_48_390#_M1000_s
+ N_A_48_390#_M1002_g N_A_48_390#_M1001_g N_A_48_390#_M1007_g
+ N_A_48_390#_M1005_g N_A_48_390#_c_149_n N_A_48_390#_c_139_n
+ N_A_48_390#_c_140_n N_A_48_390#_c_141_n N_A_48_390#_c_142_n
+ N_A_48_390#_c_143_n N_A_48_390#_c_144_n N_A_48_390#_c_145_n
+ N_A_48_390#_c_146_n PM_SKY130_FD_SC_LP__OR2_2%A_48_390#
x_PM_SKY130_FD_SC_LP__OR2_2%VPWR N_VPWR_M1006_d N_VPWR_M1005_d N_VPWR_c_222_n
+ N_VPWR_c_223_n N_VPWR_c_224_n N_VPWR_c_225_n VPWR N_VPWR_c_226_n
+ N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_221_n PM_SKY130_FD_SC_LP__OR2_2%VPWR
x_PM_SKY130_FD_SC_LP__OR2_2%X N_X_M1002_s N_X_M1001_s N_X_c_271_p N_X_c_249_n
+ N_X_c_252_n N_X_c_250_n X X X PM_SKY130_FD_SC_LP__OR2_2%X
x_PM_SKY130_FD_SC_LP__OR2_2%VGND N_VGND_M1004_s N_VGND_M1003_d N_VGND_M1007_d
+ N_VGND_c_274_n N_VGND_c_275_n N_VGND_c_276_n N_VGND_c_277_n N_VGND_c_278_n
+ N_VGND_c_279_n VGND N_VGND_c_280_n N_VGND_c_281_n N_VGND_c_282_n
+ N_VGND_c_283_n PM_SKY130_FD_SC_LP__OR2_2%VGND
cc_1 VNB N_B_c_56_n 0.0161914f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.69
cc_2 VNB N_B_M1004_g 0.0243261f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.445
cc_3 VNB N_B_c_58_n 0.029961f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.94
cc_4 VNB N_B_c_59_n 0.0183495f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_5 VNB B 0.0355109f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_B_c_61_n 0.03004f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.955
cc_7 VNB N_A_M1003_g 0.0382194f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.79
cc_8 VNB N_A_M1006_g 0.00983652f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.84
cc_9 VNB N_A_c_99_n 0.0334894f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.94
cc_10 VNB N_A_c_100_n 0.00317185f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_11 VNB N_A_48_390#_M1002_g 0.0210764f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.16
cc_12 VNB N_A_48_390#_M1001_g 0.0026975f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_A_48_390#_M1007_g 0.0278741f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.765
cc_14 VNB N_A_48_390#_M1005_g 0.00392723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_48_390#_c_139_n 0.00931001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_48_390#_c_140_n 0.00176558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_48_390#_c_141_n 8.89968e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_48_390#_c_142_n 0.00484773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_48_390#_c_143_n 0.00412654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_48_390#_c_144_n 0.00156696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_48_390#_c_145_n 0.00387775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_48_390#_c_146_n 0.062606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_221_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_249_n 0.00286337f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_25 VNB N_X_c_250_n 0.0018296f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.765
cc_26 VNB N_VGND_c_274_n 0.0119006f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.94
cc_27 VNB N_VGND_c_275_n 0.0191247f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.94
cc_28 VNB N_VGND_c_276_n 0.0043455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_277_n 0.0113226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_278_n 0.028433f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_31 VNB N_VGND_c_279_n 0.0193203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_280_n 0.0162793f $X=-0.19 $Y=-0.245 $X2=0.245 $Y2=0.925
cc_33 VNB N_VGND_c_281_n 0.0152549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_282_n 0.0063162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_283_n 0.148723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_B_c_56_n 0.00214245f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.69
cc_37 VPB N_B_c_63_n 0.0224907f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.84
cc_38 VPB N_B_c_64_n 0.0249685f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.765
cc_39 VPB N_A_M1006_g 0.0266898f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.84
cc_40 VPB N_A_48_390#_M1001_g 0.0232385f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_41 VPB N_A_48_390#_M1005_g 0.0263513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_48_390#_c_149_n 0.00626523f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.955
cc_43 VPB N_A_48_390#_c_139_n 0.00876374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_48_390#_c_140_n 0.00590548f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_48_390#_c_145_n 0.00283244f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_222_n 0.0305226f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.16
cc_47 VPB N_VPWR_c_223_n 0.0291968f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_48 VPB N_VPWR_c_224_n 0.0112967f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_49 VPB N_VPWR_c_225_n 0.0348039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_226_n 0.0326924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_227_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0.245 $Y2=0.925
cc_52 VPB N_VPWR_c_228_n 0.00795653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_221_n 0.0751077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_X_c_249_n 0.00172475f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_55 VPB N_X_c_252_n 0.00399743f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.765
cc_56 N_B_M1004_g N_A_M1003_g 0.0201614f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_57 B N_A_M1003_g 0.00138253f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_58 N_B_c_61_n N_A_M1003_g 0.00645674f $X=0.27 $Y=0.955 $X2=0 $Y2=0
cc_59 N_B_c_56_n N_A_M1006_g 0.00662377f $X=0.36 $Y=1.69 $X2=0 $Y2=0
cc_60 N_B_c_64_n N_A_M1006_g 0.0489386f $X=0.58 $Y=1.765 $X2=0 $Y2=0
cc_61 N_B_c_64_n N_A_c_99_n 6.25947e-19 $X=0.58 $Y=1.765 $X2=0 $Y2=0
cc_62 B N_A_c_99_n 3.16581e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_63 N_B_c_61_n N_A_c_99_n 0.0206847f $X=0.27 $Y=0.955 $X2=0 $Y2=0
cc_64 N_B_c_58_n N_A_c_100_n 4.22191e-19 $X=0.345 $Y=0.94 $X2=0 $Y2=0
cc_65 N_B_c_64_n N_A_c_100_n 4.45351e-19 $X=0.58 $Y=1.765 $X2=0 $Y2=0
cc_66 B N_A_c_100_n 0.0247801f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_67 N_B_c_61_n N_A_c_100_n 0.00187742f $X=0.27 $Y=0.955 $X2=0 $Y2=0
cc_68 N_B_c_63_n N_A_48_390#_c_149_n 0.00443413f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_69 N_B_c_64_n N_A_48_390#_c_149_n 0.00583408f $X=0.58 $Y=1.765 $X2=0 $Y2=0
cc_70 N_B_c_58_n N_A_48_390#_c_139_n 0.00255178f $X=0.345 $Y=0.94 $X2=0 $Y2=0
cc_71 N_B_c_64_n N_A_48_390#_c_139_n 0.0134561f $X=0.58 $Y=1.765 $X2=0 $Y2=0
cc_72 N_B_c_56_n N_A_48_390#_c_140_n 0.0059382f $X=0.36 $Y=1.69 $X2=0 $Y2=0
cc_73 N_B_c_58_n N_A_48_390#_c_140_n 9.77567e-19 $X=0.345 $Y=0.94 $X2=0 $Y2=0
cc_74 N_B_c_64_n N_A_48_390#_c_140_n 0.00403333f $X=0.58 $Y=1.765 $X2=0 $Y2=0
cc_75 B N_A_48_390#_c_140_n 0.0122176f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_76 N_B_M1004_g N_A_48_390#_c_141_n 0.00209872f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_77 N_B_M1004_g N_A_48_390#_c_143_n 0.00331263f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_78 B N_A_48_390#_c_143_n 0.00828995f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_79 N_B_c_63_n N_VPWR_c_222_n 0.00213306f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_80 N_B_c_63_n N_VPWR_c_221_n 0.00386017f $X=0.58 $Y=1.84 $X2=0 $Y2=0
cc_81 N_B_M1004_g N_VGND_c_275_n 0.00370449f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_82 N_B_c_58_n N_VGND_c_275_n 0.00203332f $X=0.345 $Y=0.94 $X2=0 $Y2=0
cc_83 B N_VGND_c_275_n 0.0210248f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_84 N_B_M1004_g N_VGND_c_280_n 0.00585385f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_85 N_B_M1004_g N_VGND_c_283_n 0.011707f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_86 N_B_c_58_n N_VGND_c_283_n 3.96635e-19 $X=0.345 $Y=0.94 $X2=0 $Y2=0
cc_87 B N_VGND_c_283_n 0.00274317f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_A_48_390#_M1002_g 0.0232588f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_M1006_g N_A_48_390#_M1001_g 0.0172089f $X=0.94 $Y=2.16 $X2=0 $Y2=0
cc_90 N_A_M1006_g N_A_48_390#_c_139_n 0.014791f $X=0.94 $Y=2.16 $X2=0 $Y2=0
cc_91 N_A_c_99_n N_A_48_390#_c_139_n 0.00487498f $X=0.81 $Y=1.315 $X2=0 $Y2=0
cc_92 N_A_c_100_n N_A_48_390#_c_139_n 0.0297931f $X=0.81 $Y=1.315 $X2=0 $Y2=0
cc_93 N_A_M1003_g N_A_48_390#_c_141_n 0.0067791f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_M1003_g N_A_48_390#_c_142_n 0.0119209f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_c_100_n N_A_48_390#_c_142_n 0.00537189f $X=0.81 $Y=1.315 $X2=0 $Y2=0
cc_96 N_A_M1003_g N_A_48_390#_c_143_n 0.00177814f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_c_99_n N_A_48_390#_c_143_n 0.00486942f $X=0.81 $Y=1.315 $X2=0 $Y2=0
cc_98 N_A_c_100_n N_A_48_390#_c_143_n 0.0175007f $X=0.81 $Y=1.315 $X2=0 $Y2=0
cc_99 N_A_M1003_g N_A_48_390#_c_144_n 0.00684931f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_c_100_n N_A_48_390#_c_144_n 0.00825735f $X=0.81 $Y=1.315 $X2=0 $Y2=0
cc_101 N_A_c_99_n N_A_48_390#_c_145_n 0.00494493f $X=0.81 $Y=1.315 $X2=0 $Y2=0
cc_102 N_A_c_100_n N_A_48_390#_c_145_n 0.0125792f $X=0.81 $Y=1.315 $X2=0 $Y2=0
cc_103 N_A_c_99_n N_A_48_390#_c_146_n 0.0203712f $X=0.81 $Y=1.315 $X2=0 $Y2=0
cc_104 N_A_M1006_g N_VPWR_c_222_n 0.0145489f $X=0.94 $Y=2.16 $X2=0 $Y2=0
cc_105 N_A_M1006_g N_VPWR_c_221_n 0.00247051f $X=0.94 $Y=2.16 $X2=0 $Y2=0
cc_106 N_A_M1003_g N_VGND_c_276_n 0.00177437f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_M1003_g N_VGND_c_280_n 0.00436698f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_M1003_g N_VGND_c_283_n 0.00609604f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_48_390#_M1001_g N_VPWR_c_222_n 0.00622366f $X=1.465 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_48_390#_c_139_n N_VPWR_c_222_n 0.0155325f $X=1.185 $Y=1.715 $X2=0
+ $Y2=0
cc_111 N_A_48_390#_c_145_n N_VPWR_c_222_n 0.0155264f $X=1.39 $Y=1.44 $X2=0 $Y2=0
cc_112 N_A_48_390#_c_146_n N_VPWR_c_222_n 6.65145e-19 $X=1.895 $Y=1.44 $X2=0
+ $Y2=0
cc_113 N_A_48_390#_M1005_g N_VPWR_c_223_n 0.00511185f $X=1.895 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_48_390#_M1001_g N_VPWR_c_225_n 6.96433e-19 $X=1.465 $Y=2.465 $X2=0
+ $Y2=0
cc_115 N_A_48_390#_M1005_g N_VPWR_c_225_n 0.0154728f $X=1.895 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_48_390#_M1001_g N_VPWR_c_227_n 0.00585385f $X=1.465 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_48_390#_M1005_g N_VPWR_c_227_n 0.00486043f $X=1.895 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_48_390#_M1001_g N_VPWR_c_221_n 0.0118358f $X=1.465 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_A_48_390#_M1005_g N_VPWR_c_221_n 0.00824727f $X=1.895 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_48_390#_M1002_g N_X_c_249_n 9.50605e-19 $X=1.465 $Y=0.655 $X2=0 $Y2=0
cc_121 N_A_48_390#_M1001_g N_X_c_249_n 0.00120642f $X=1.465 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_48_390#_M1005_g N_X_c_249_n 0.00559377f $X=1.895 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_48_390#_c_144_n N_X_c_249_n 0.00781615f $X=1.3 $Y=1.275 $X2=0 $Y2=0
cc_124 N_A_48_390#_c_145_n N_X_c_249_n 0.0330347f $X=1.39 $Y=1.44 $X2=0 $Y2=0
cc_125 N_A_48_390#_c_146_n N_X_c_249_n 0.0264224f $X=1.895 $Y=1.44 $X2=0 $Y2=0
cc_126 N_A_48_390#_M1001_g N_X_c_252_n 0.00193384f $X=1.465 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_48_390#_c_145_n N_X_c_252_n 0.00305014f $X=1.39 $Y=1.44 $X2=0 $Y2=0
cc_128 N_A_48_390#_c_146_n N_X_c_252_n 4.50677e-19 $X=1.895 $Y=1.44 $X2=0 $Y2=0
cc_129 N_A_48_390#_M1002_g N_X_c_250_n 9.89688e-19 $X=1.465 $Y=0.655 $X2=0 $Y2=0
cc_130 N_A_48_390#_M1007_g N_X_c_250_n 0.00477868f $X=1.895 $Y=0.655 $X2=0 $Y2=0
cc_131 N_A_48_390#_c_144_n N_X_c_250_n 0.0111836f $X=1.3 $Y=1.275 $X2=0 $Y2=0
cc_132 N_A_48_390#_c_146_n N_X_c_250_n 4.65933e-19 $X=1.895 $Y=1.44 $X2=0 $Y2=0
cc_133 N_A_48_390#_c_142_n N_VGND_M1003_d 0.00460078f $X=1.185 $Y=0.81 $X2=0
+ $Y2=0
cc_134 N_A_48_390#_c_144_n N_VGND_M1003_d 0.00230255f $X=1.3 $Y=1.275 $X2=0
+ $Y2=0
cc_135 N_A_48_390#_M1002_g N_VGND_c_276_n 0.00173608f $X=1.465 $Y=0.655 $X2=0
+ $Y2=0
cc_136 N_A_48_390#_c_142_n N_VGND_c_276_n 0.0227452f $X=1.185 $Y=0.81 $X2=0
+ $Y2=0
cc_137 N_A_48_390#_M1007_g N_VGND_c_278_n 0.00465399f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_138 N_A_48_390#_M1002_g N_VGND_c_279_n 5.85269e-19 $X=1.465 $Y=0.655 $X2=0
+ $Y2=0
cc_139 N_A_48_390#_M1007_g N_VGND_c_279_n 0.0112393f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_140 N_A_48_390#_c_141_n N_VGND_c_280_n 0.0156912f $X=0.725 $Y=0.42 $X2=0
+ $Y2=0
cc_141 N_A_48_390#_c_142_n N_VGND_c_280_n 0.00230424f $X=1.185 $Y=0.81 $X2=0
+ $Y2=0
cc_142 N_A_48_390#_M1002_g N_VGND_c_281_n 0.00560773f $X=1.465 $Y=0.655 $X2=0
+ $Y2=0
cc_143 N_A_48_390#_M1007_g N_VGND_c_281_n 0.00486043f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_144 N_A_48_390#_c_142_n N_VGND_c_281_n 5.15771e-19 $X=1.185 $Y=0.81 $X2=0
+ $Y2=0
cc_145 N_A_48_390#_M1004_d N_VGND_c_283_n 0.00240953f $X=0.585 $Y=0.235 $X2=0
+ $Y2=0
cc_146 N_A_48_390#_M1002_g N_VGND_c_283_n 0.010029f $X=1.465 $Y=0.655 $X2=0
+ $Y2=0
cc_147 N_A_48_390#_M1007_g N_VGND_c_283_n 0.00824727f $X=1.895 $Y=0.655 $X2=0
+ $Y2=0
cc_148 N_A_48_390#_c_141_n N_VGND_c_283_n 0.0106994f $X=0.725 $Y=0.42 $X2=0
+ $Y2=0
cc_149 N_A_48_390#_c_142_n N_VGND_c_283_n 0.00622123f $X=1.185 $Y=0.81 $X2=0
+ $Y2=0
cc_150 N_VPWR_c_221_n N_X_M1001_s 0.00397496f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_151 N_VPWR_c_223_n N_X_c_252_n 0.00154926f $X=2.11 $Y=2.26 $X2=0 $Y2=0
cc_152 N_VPWR_c_227_n X 0.0138717f $X=1.945 $Y=3.33 $X2=0 $Y2=0
cc_153 N_VPWR_c_221_n X 0.00886411f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_154 N_X_c_250_n N_VGND_c_278_n 0.00153077f $X=1.7 $Y=1.14 $X2=0 $Y2=0
cc_155 N_X_c_271_p N_VGND_c_281_n 0.0124525f $X=1.68 $Y=0.42 $X2=0 $Y2=0
cc_156 N_X_M1002_s N_VGND_c_283_n 0.00536646f $X=1.54 $Y=0.235 $X2=0 $Y2=0
cc_157 N_X_c_271_p N_VGND_c_283_n 0.00730901f $X=1.68 $Y=0.42 $X2=0 $Y2=0
