* File: sky130_fd_sc_lp__clkbuf_1.pxi.spice
* Created: Fri Aug 28 10:14:48 2020
* 
x_PM_SKY130_FD_SC_LP__CLKBUF_1%A_69_161# N_A_69_161#_M1002_d N_A_69_161#_M1000_d
+ N_A_69_161#_M1001_g N_A_69_161#_M1003_g N_A_69_161#_c_35_n N_A_69_161#_c_36_n
+ N_A_69_161#_c_41_n N_A_69_161#_c_37_n N_A_69_161#_c_42_n N_A_69_161#_c_38_n
+ N_A_69_161#_c_39_n PM_SKY130_FD_SC_LP__CLKBUF_1%A_69_161#
x_PM_SKY130_FD_SC_LP__CLKBUF_1%A N_A_M1000_g N_A_M1002_g A N_A_c_86_n N_A_c_87_n
+ A PM_SKY130_FD_SC_LP__CLKBUF_1%A
x_PM_SKY130_FD_SC_LP__CLKBUF_1%X N_X_M1001_s N_X_M1003_s N_X_c_118_n X X X X
+ N_X_c_120_n X PM_SKY130_FD_SC_LP__CLKBUF_1%X
x_PM_SKY130_FD_SC_LP__CLKBUF_1%VPWR N_VPWR_M1003_d N_VPWR_c_139_n VPWR
+ N_VPWR_c_140_n N_VPWR_c_141_n N_VPWR_c_138_n N_VPWR_c_143_n
+ PM_SKY130_FD_SC_LP__CLKBUF_1%VPWR
x_PM_SKY130_FD_SC_LP__CLKBUF_1%VGND N_VGND_M1001_d N_VGND_c_158_n VGND
+ N_VGND_c_159_n N_VGND_c_160_n N_VGND_c_161_n N_VGND_c_162_n
+ PM_SKY130_FD_SC_LP__CLKBUF_1%VGND
cc_1 VNB N_A_69_161#_M1001_g 0.0213921f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.465
cc_2 VNB N_A_69_161#_M1003_g 0.0289756f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_3 VNB N_A_69_161#_c_35_n 0.003896f $X=-0.19 $Y=-0.245 $X2=1.045 $Y2=0.97
cc_4 VNB N_A_69_161#_c_36_n 0.0346228f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.97
cc_5 VNB N_A_69_161#_c_37_n 0.0217203f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=0.465
cc_6 VNB N_A_69_161#_c_38_n 0.0243778f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.92
cc_7 VNB N_A_69_161#_c_39_n 0.0193996f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.97
cc_8 VNB N_A_M1002_g 0.0529541f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.805
cc_9 VNB N_A_c_86_n 0.025799f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_10 VNB N_A_c_87_n 0.00342117f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_11 VNB N_X_c_118_n 0.013747f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.465
cc_12 VNB X 0.0114707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_X_c_120_n 0.0422583f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.135
cc_14 VNB N_VPWR_c_138_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=2.1
cc_15 VNB N_VGND_c_158_n 0.00592013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_159_n 0.0182657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_160_n 0.0174691f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.97
cc_18 VNB N_VGND_c_161_n 0.112498f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.97
cc_19 VNB N_VGND_c_162_n 0.00526527f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=2.905
cc_20 VPB N_A_69_161#_M1003_g 0.023346f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_21 VPB N_A_69_161#_c_41_n 0.0411921f $X=-0.19 $Y=1.655 $X2=1.125 $Y2=2.905
cc_22 VPB N_A_69_161#_c_42_n 0.00747259f $X=-0.19 $Y=1.655 $X2=1.125 $Y2=2.085
cc_23 VPB N_A_69_161#_c_38_n 0.012168f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=1.92
cc_24 VPB N_A_M1000_g 0.0213969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 VPB N_A_c_86_n 0.00764657f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_26 VPB N_A_c_87_n 0.00389708f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_27 VPB X 0.0588167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_139_n 0.00522139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_140_n 0.0172252f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.465
cc_30 VPB N_VPWR_c_141_n 0.0183459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_138_n 0.04424f $X=-0.19 $Y=1.655 $X2=1.175 $Y2=2.1
cc_32 VPB N_VPWR_c_143_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 N_A_69_161#_M1003_g N_A_M1000_g 0.0161582f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_34 N_A_69_161#_c_38_n N_A_M1000_g 0.0043607f $X=1.175 $Y=1.92 $X2=0 $Y2=0
cc_35 N_A_69_161#_M1001_g N_A_M1002_g 0.0107736f $X=0.48 $Y=0.465 $X2=0 $Y2=0
cc_36 N_A_69_161#_M1003_g N_A_M1002_g 0.00773538f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_37 N_A_69_161#_c_35_n N_A_M1002_g 0.0210085f $X=1.045 $Y=0.97 $X2=0 $Y2=0
cc_38 N_A_69_161#_c_36_n N_A_M1002_g 0.0213328f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_39 N_A_69_161#_c_37_n N_A_M1002_g 0.00595534f $X=1.175 $Y=0.465 $X2=0 $Y2=0
cc_40 N_A_69_161#_c_38_n N_A_M1002_g 0.00558047f $X=1.175 $Y=1.92 $X2=0 $Y2=0
cc_41 N_A_69_161#_M1003_g N_A_c_86_n 0.0204969f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_42 N_A_69_161#_c_35_n N_A_c_86_n 0.00324655f $X=1.045 $Y=0.97 $X2=0 $Y2=0
cc_43 N_A_69_161#_c_42_n N_A_c_86_n 0.00282521f $X=1.125 $Y=2.085 $X2=0 $Y2=0
cc_44 N_A_69_161#_c_38_n N_A_c_86_n 0.00863799f $X=1.175 $Y=1.92 $X2=0 $Y2=0
cc_45 N_A_69_161#_c_39_n N_A_c_86_n 0.00214147f $X=1.2 $Y=0.97 $X2=0 $Y2=0
cc_46 N_A_69_161#_M1003_g N_A_c_87_n 0.00342332f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_47 N_A_69_161#_c_35_n N_A_c_87_n 0.025912f $X=1.045 $Y=0.97 $X2=0 $Y2=0
cc_48 N_A_69_161#_c_36_n N_A_c_87_n 8.95202e-19 $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_49 N_A_69_161#_c_38_n N_A_c_87_n 0.0309912f $X=1.175 $Y=1.92 $X2=0 $Y2=0
cc_50 N_A_69_161#_M1001_g N_X_c_118_n 0.00463188f $X=0.48 $Y=0.465 $X2=0 $Y2=0
cc_51 N_A_69_161#_c_35_n N_X_c_118_n 3.65009e-19 $X=1.045 $Y=0.97 $X2=0 $Y2=0
cc_52 N_A_69_161#_c_36_n N_X_c_118_n 0.00127441f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_53 N_A_69_161#_M1003_g X 0.0113345f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_54 N_A_69_161#_c_36_n X 0.00172472f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_55 N_A_69_161#_M1001_g N_X_c_120_n 0.00549866f $X=0.48 $Y=0.465 $X2=0 $Y2=0
cc_56 N_A_69_161#_M1003_g N_X_c_120_n 0.0112861f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_57 N_A_69_161#_c_35_n N_X_c_120_n 0.0262099f $X=1.045 $Y=0.97 $X2=0 $Y2=0
cc_58 N_A_69_161#_c_36_n N_X_c_120_n 0.00816168f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_59 N_A_69_161#_M1003_g N_VPWR_c_139_n 0.00328234f $X=0.48 $Y=2.465 $X2=0
+ $Y2=0
cc_60 N_A_69_161#_M1003_g N_VPWR_c_140_n 0.00585385f $X=0.48 $Y=2.465 $X2=0
+ $Y2=0
cc_61 N_A_69_161#_c_41_n N_VPWR_c_141_n 0.0237126f $X=1.125 $Y=2.905 $X2=0 $Y2=0
cc_62 N_A_69_161#_M1000_d N_VPWR_c_138_n 0.00249946f $X=0.985 $Y=1.835 $X2=0
+ $Y2=0
cc_63 N_A_69_161#_M1003_g N_VPWR_c_138_n 0.011485f $X=0.48 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A_69_161#_c_41_n N_VPWR_c_138_n 0.0139182f $X=1.125 $Y=2.905 $X2=0 $Y2=0
cc_65 N_A_69_161#_M1001_g N_VGND_c_158_n 0.00300513f $X=0.48 $Y=0.465 $X2=0
+ $Y2=0
cc_66 N_A_69_161#_c_35_n N_VGND_c_158_n 0.0202667f $X=1.045 $Y=0.97 $X2=0 $Y2=0
cc_67 N_A_69_161#_c_36_n N_VGND_c_158_n 0.00169036f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_68 N_A_69_161#_M1001_g N_VGND_c_159_n 0.0052984f $X=0.48 $Y=0.465 $X2=0 $Y2=0
cc_69 N_A_69_161#_c_37_n N_VGND_c_160_n 0.0156318f $X=1.175 $Y=0.465 $X2=0 $Y2=0
cc_70 N_A_69_161#_M1001_g N_VGND_c_161_n 0.0069061f $X=0.48 $Y=0.465 $X2=0 $Y2=0
cc_71 N_A_69_161#_c_35_n N_VGND_c_161_n 0.0116632f $X=1.045 $Y=0.97 $X2=0 $Y2=0
cc_72 N_A_69_161#_c_36_n N_VGND_c_161_n 0.00106485f $X=0.51 $Y=0.97 $X2=0 $Y2=0
cc_73 N_A_69_161#_c_37_n N_VGND_c_161_n 0.0117053f $X=1.175 $Y=0.465 $X2=0 $Y2=0
cc_74 N_A_c_87_n X 0.0147469f $X=0.93 $Y=1.51 $X2=0 $Y2=0
cc_75 N_A_c_87_n N_X_c_120_n 0.00819403f $X=0.93 $Y=1.51 $X2=0 $Y2=0
cc_76 N_A_M1000_g N_VPWR_c_139_n 0.00328234f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A_c_86_n N_VPWR_c_139_n 2.78168e-19 $X=0.93 $Y=1.51 $X2=0 $Y2=0
cc_78 N_A_c_87_n N_VPWR_c_139_n 0.0145685f $X=0.93 $Y=1.51 $X2=0 $Y2=0
cc_79 N_A_M1000_g N_VPWR_c_141_n 0.00585385f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A_M1000_g N_VPWR_c_138_n 0.0115284f $X=0.91 $Y=2.465 $X2=0 $Y2=0
cc_81 N_A_M1002_g N_VGND_c_158_n 0.0032119f $X=0.96 $Y=0.465 $X2=0 $Y2=0
cc_82 N_A_M1002_g N_VGND_c_160_n 0.00565115f $X=0.96 $Y=0.465 $X2=0 $Y2=0
cc_83 N_A_M1002_g N_VGND_c_161_n 0.00697852f $X=0.96 $Y=0.465 $X2=0 $Y2=0
cc_84 X N_VPWR_c_140_n 0.0201282f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_85 N_X_M1003_s N_VPWR_c_138_n 0.00249946f $X=0.14 $Y=1.835 $X2=0 $Y2=0
cc_86 X N_VPWR_c_138_n 0.0119743f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_87 N_X_c_118_n N_VGND_c_159_n 0.0164381f $X=0.265 $Y=0.465 $X2=0 $Y2=0
cc_88 N_X_c_118_n N_VGND_c_161_n 0.0127105f $X=0.265 $Y=0.465 $X2=0 $Y2=0
