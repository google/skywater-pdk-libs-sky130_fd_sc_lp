* File: sky130_fd_sc_lp__and3b_1.pxi.spice
* Created: Wed Sep  2 09:32:06 2020
* 
x_PM_SKY130_FD_SC_LP__AND3B_1%A_N N_A_N_c_69_n N_A_N_M1003_g N_A_N_M1006_g
+ N_A_N_c_72_n A_N A_N A_N A_N N_A_N_c_74_n PM_SKY130_FD_SC_LP__AND3B_1%A_N
x_PM_SKY130_FD_SC_LP__AND3B_1%A_110_47# N_A_110_47#_M1003_d N_A_110_47#_M1006_d
+ N_A_110_47#_c_96_n N_A_110_47#_c_97_n N_A_110_47#_M1004_g N_A_110_47#_c_99_n
+ N_A_110_47#_M1007_g N_A_110_47#_c_100_n N_A_110_47#_c_101_n
+ N_A_110_47#_c_102_n N_A_110_47#_c_103_n N_A_110_47#_c_106_n
+ N_A_110_47#_c_104_n PM_SKY130_FD_SC_LP__AND3B_1%A_110_47#
x_PM_SKY130_FD_SC_LP__AND3B_1%B N_B_M1002_g N_B_M1008_g B B B N_B_c_157_n
+ PM_SKY130_FD_SC_LP__AND3B_1%B
x_PM_SKY130_FD_SC_LP__AND3B_1%C N_C_M1009_g N_C_M1001_g N_C_c_192_n N_C_c_193_n
+ N_C_c_194_n C C C N_C_c_196_n PM_SKY130_FD_SC_LP__AND3B_1%C
x_PM_SKY130_FD_SC_LP__AND3B_1%A_185_367# N_A_185_367#_M1007_s
+ N_A_185_367#_M1004_s N_A_185_367#_M1002_d N_A_185_367#_M1000_g
+ N_A_185_367#_M1005_g N_A_185_367#_c_244_n N_A_185_367#_c_232_n
+ N_A_185_367#_c_238_n N_A_185_367#_c_239_n N_A_185_367#_c_240_n
+ N_A_185_367#_c_233_n N_A_185_367#_c_241_n N_A_185_367#_c_234_n
+ N_A_185_367#_c_235_n PM_SKY130_FD_SC_LP__AND3B_1%A_185_367#
x_PM_SKY130_FD_SC_LP__AND3B_1%VPWR N_VPWR_M1006_s N_VPWR_M1004_d N_VPWR_M1001_d
+ N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_315_n
+ N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n VPWR N_VPWR_c_319_n
+ N_VPWR_c_310_n PM_SKY130_FD_SC_LP__AND3B_1%VPWR
x_PM_SKY130_FD_SC_LP__AND3B_1%X N_X_M1005_d N_X_M1000_d N_X_c_345_n N_X_c_346_n
+ X X X N_X_c_347_n X PM_SKY130_FD_SC_LP__AND3B_1%X
x_PM_SKY130_FD_SC_LP__AND3B_1%VGND N_VGND_M1003_s N_VGND_M1009_d N_VGND_c_363_n
+ N_VGND_c_364_n N_VGND_c_365_n VGND N_VGND_c_366_n N_VGND_c_367_n
+ N_VGND_c_368_n N_VGND_c_369_n PM_SKY130_FD_SC_LP__AND3B_1%VGND
cc_1 VNB N_A_N_c_69_n 0.0209464f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.288
cc_2 VNB N_A_N_M1003_g 0.0304076f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_3 VNB N_A_N_M1006_g 0.0094104f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_4 VNB N_A_N_c_72_n 0.0302281f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_5 VNB A_N 0.0352546f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A_N_c_74_n 0.0292967f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_7 VNB N_A_110_47#_c_96_n 0.0279074f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_8 VNB N_A_110_47#_c_97_n 0.0163812f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_9 VNB N_A_110_47#_M1004_g 0.0132677f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_10 VNB N_A_110_47#_c_99_n 0.0195604f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A_110_47#_c_100_n 0.0270399f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.005
cc_12 VNB N_A_110_47#_c_101_n 0.00599842f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.925
cc_13 VNB N_A_110_47#_c_102_n 0.0169397f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_14 VNB N_A_110_47#_c_103_n 0.0224012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_110_47#_c_104_n 0.00396954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_M1002_g 0.0098643f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.84
cc_17 VNB N_B_M1008_g 0.0345641f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_18 VNB B 0.00475756f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_19 VNB N_B_c_157_n 0.0340613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_M1001_g 0.0123005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C_c_192_n 0.016615f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_22 VNB N_C_c_193_n 0.0229855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_c_194_n 0.0156706f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_24 VNB C 0.0071558f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_25 VNB N_C_c_196_n 0.0169877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_185_367#_M1005_g 0.0298752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_185_367#_c_232_n 0.00906157f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=0.84
cc_28 VNB N_A_185_367#_c_233_n 0.00352778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_185_367#_c_234_n 0.00576014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_185_367#_c_235_n 0.0280315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_310_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_345_n 0.0276295f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_33 VNB N_X_c_346_n 0.00861101f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_X_c_347_n 0.0281863f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.035
cc_35 VNB N_VGND_c_363_n 0.0109765f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_36 VNB N_VGND_c_364_n 0.0198639f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.77
cc_37 VNB N_VGND_c_365_n 0.00818742f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_38 VNB N_VGND_c_366_n 0.0572704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_367_n 0.015618f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_40 VNB N_VGND_c_368_n 0.191187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_369_n 0.00474961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_A_N_M1006_g 0.0828131f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.77
cc_43 VPB A_N 0.0342825f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_44 VPB N_A_110_47#_M1004_g 0.0270468f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.51
cc_45 VPB N_A_110_47#_c_106_n 0.00712513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_110_47#_c_104_n 0.0212985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B_M1002_g 0.0244724f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.84
cc_48 VPB N_C_M1001_g 0.0232145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_185_367#_M1000_g 0.0250005f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_50 VPB N_A_185_367#_c_232_n 3.70161e-19 $X=-0.19 $Y=1.655 $X2=0.327 $Y2=0.84
cc_51 VPB N_A_185_367#_c_238_n 0.00634603f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=0.925
cc_52 VPB N_A_185_367#_c_239_n 0.00409329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_185_367#_c_240_n 0.00466398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_185_367#_c_241_n 0.00707384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_185_367#_c_234_n 0.00163954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_185_367#_c_235_n 0.00604755f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_311_n 0.0109759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_312_n 0.0267403f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_59 VPB N_VPWR_c_313_n 0.0417022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_314_n 0.017962f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.005
cc_61 VPB N_VPWR_c_315_n 0.0283745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_316_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_317_n 0.0193478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_318_n 0.00699479f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.665
cc_65 VPB N_VPWR_c_319_n 0.0207215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_310_n 0.0938625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB X 0.0552502f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_68 VPB N_X_c_347_n 0.00970872f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.035
cc_69 N_A_N_M1003_g N_A_110_47#_c_97_n 0.0117265f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_70 A_N N_A_110_47#_c_97_n 4.05374e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_71 N_A_N_c_72_n N_A_110_47#_M1004_g 0.00788602f $X=0.327 $Y=1.51 $X2=0 $Y2=0
cc_72 N_A_N_c_69_n N_A_110_47#_c_100_n 0.0117265f $X=0.327 $Y=1.288 $X2=0 $Y2=0
cc_73 N_A_N_M1003_g N_A_110_47#_c_101_n 0.0113632f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_74 A_N N_A_110_47#_c_102_n 0.112486f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_75 N_A_N_c_74_n N_A_110_47#_c_102_n 0.0113632f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_76 N_A_N_c_74_n N_A_110_47#_c_103_n 0.0117265f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_77 N_A_N_c_72_n N_A_110_47#_c_104_n 0.0113632f $X=0.327 $Y=1.51 $X2=0 $Y2=0
cc_78 N_A_N_M1006_g N_VPWR_c_312_n 0.00583068f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_79 A_N N_VPWR_c_312_n 0.0139182f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 N_A_N_M1006_g N_VPWR_c_315_n 0.00478016f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_81 N_A_N_M1006_g N_VPWR_c_310_n 0.00977894f $X=0.475 $Y=2.77 $X2=0 $Y2=0
cc_82 N_A_N_M1003_g N_VGND_c_364_n 0.00525416f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_83 A_N N_VGND_c_364_n 0.0213581f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A_N_c_74_n N_VGND_c_364_n 0.001893f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_85 N_A_N_M1003_g N_VGND_c_366_n 0.00585385f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A_N_M1003_g N_VGND_c_368_n 0.0131279f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_87 A_N N_VGND_c_368_n 0.00163474f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A_110_47#_M1004_g N_B_M1002_g 0.0166634f $X=1.265 $Y=2.045 $X2=0 $Y2=0
cc_89 N_A_110_47#_c_99_n N_B_M1008_g 0.0502741f $X=1.445 $Y=0.765 $X2=0 $Y2=0
cc_90 N_A_110_47#_c_103_n N_B_M1008_g 0.00185604f $X=0.955 $Y=0.93 $X2=0 $Y2=0
cc_91 N_A_110_47#_c_99_n B 0.00280601f $X=1.445 $Y=0.765 $X2=0 $Y2=0
cc_92 N_A_110_47#_c_100_n B 2.17247e-19 $X=1.265 $Y=1.36 $X2=0 $Y2=0
cc_93 N_A_110_47#_c_100_n N_B_c_157_n 0.0124557f $X=1.265 $Y=1.36 $X2=0 $Y2=0
cc_94 N_A_110_47#_c_103_n N_B_c_157_n 8.44703e-19 $X=0.955 $Y=0.93 $X2=0 $Y2=0
cc_95 N_A_110_47#_c_104_n N_A_185_367#_c_244_n 0.0281027f $X=0.71 $Y=2.605 $X2=0
+ $Y2=0
cc_96 N_A_110_47#_c_96_n N_A_185_367#_c_232_n 0.0113399f $X=1.37 $Y=0.84 $X2=0
+ $Y2=0
cc_97 N_A_110_47#_M1004_g N_A_185_367#_c_232_n 0.00744811f $X=1.265 $Y=2.045
+ $X2=0 $Y2=0
cc_98 N_A_110_47#_c_99_n N_A_185_367#_c_232_n 0.00408881f $X=1.445 $Y=0.765
+ $X2=0 $Y2=0
cc_99 N_A_110_47#_c_100_n N_A_185_367#_c_232_n 0.00589716f $X=1.265 $Y=1.36
+ $X2=0 $Y2=0
cc_100 N_A_110_47#_c_101_n N_A_185_367#_c_232_n 0.00821767f $X=0.69 $Y=0.445
+ $X2=0 $Y2=0
cc_101 N_A_110_47#_c_102_n N_A_185_367#_c_232_n 0.0507858f $X=0.955 $Y=0.93
+ $X2=0 $Y2=0
cc_102 N_A_110_47#_c_103_n N_A_185_367#_c_232_n 0.00206713f $X=0.955 $Y=0.93
+ $X2=0 $Y2=0
cc_103 N_A_110_47#_c_104_n N_A_185_367#_c_232_n 0.00815481f $X=0.71 $Y=2.605
+ $X2=0 $Y2=0
cc_104 N_A_110_47#_M1004_g N_A_185_367#_c_239_n 0.0153773f $X=1.265 $Y=2.045
+ $X2=0 $Y2=0
cc_105 N_A_110_47#_c_100_n N_A_185_367#_c_239_n 0.00573485f $X=1.265 $Y=1.36
+ $X2=0 $Y2=0
cc_106 N_A_110_47#_c_102_n N_A_185_367#_c_239_n 0.00762972f $X=0.955 $Y=0.93
+ $X2=0 $Y2=0
cc_107 N_A_110_47#_c_104_n N_A_185_367#_c_239_n 0.014281f $X=0.71 $Y=2.605 $X2=0
+ $Y2=0
cc_108 N_A_110_47#_c_96_n N_A_185_367#_c_233_n 7.11899e-19 $X=1.37 $Y=0.84 $X2=0
+ $Y2=0
cc_109 N_A_110_47#_c_97_n N_A_185_367#_c_233_n 0.00602633f $X=1.12 $Y=0.84 $X2=0
+ $Y2=0
cc_110 N_A_110_47#_c_99_n N_A_185_367#_c_233_n 0.00410776f $X=1.445 $Y=0.765
+ $X2=0 $Y2=0
cc_111 N_A_110_47#_c_101_n N_A_185_367#_c_233_n 0.0216288f $X=0.69 $Y=0.445
+ $X2=0 $Y2=0
cc_112 N_A_110_47#_M1004_g N_VPWR_c_313_n 0.00206718f $X=1.265 $Y=2.045 $X2=0
+ $Y2=0
cc_113 N_A_110_47#_c_106_n N_VPWR_c_313_n 0.0129013f $X=0.69 $Y=2.77 $X2=0 $Y2=0
cc_114 N_A_110_47#_c_104_n N_VPWR_c_313_n 0.0122104f $X=0.71 $Y=2.605 $X2=0
+ $Y2=0
cc_115 N_A_110_47#_c_106_n N_VPWR_c_315_n 0.00971925f $X=0.69 $Y=2.77 $X2=0
+ $Y2=0
cc_116 N_A_110_47#_c_106_n N_VPWR_c_310_n 0.0102543f $X=0.69 $Y=2.77 $X2=0 $Y2=0
cc_117 N_A_110_47#_c_97_n N_VGND_c_366_n 0.00195006f $X=1.12 $Y=0.84 $X2=0 $Y2=0
cc_118 N_A_110_47#_c_99_n N_VGND_c_366_n 0.0054833f $X=1.445 $Y=0.765 $X2=0
+ $Y2=0
cc_119 N_A_110_47#_c_101_n N_VGND_c_366_n 0.0162773f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_120 N_A_110_47#_M1003_d N_VGND_c_368_n 0.00272496f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_121 N_A_110_47#_c_97_n N_VGND_c_368_n 4.35162e-19 $X=1.12 $Y=0.84 $X2=0 $Y2=0
cc_122 N_A_110_47#_c_99_n N_VGND_c_368_n 0.011278f $X=1.445 $Y=0.765 $X2=0 $Y2=0
cc_123 N_A_110_47#_c_101_n N_VGND_c_368_n 0.0110608f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_124 N_A_110_47#_c_102_n N_VGND_c_368_n 0.00739482f $X=0.955 $Y=0.93 $X2=0
+ $Y2=0
cc_125 N_B_M1002_g N_C_M1001_g 0.0199035f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_126 N_B_c_157_n N_C_M1001_g 0.00210398f $X=1.715 $Y=1.32 $X2=0 $Y2=0
cc_127 N_B_M1008_g N_C_c_192_n 0.0405405f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_128 B N_C_c_192_n 0.00112803f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_129 N_B_c_157_n N_C_c_193_n 0.0405405f $X=1.715 $Y=1.32 $X2=0 $Y2=0
cc_130 N_B_M1008_g C 0.005709f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_131 B C 0.0815721f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_132 N_B_M1002_g N_A_185_367#_c_232_n 0.00346998f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_133 N_B_M1008_g N_A_185_367#_c_232_n 0.00109083f $X=1.805 $Y=0.445 $X2=0
+ $Y2=0
cc_134 B N_A_185_367#_c_232_n 0.0653386f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_135 N_B_c_157_n N_A_185_367#_c_232_n 0.00347462f $X=1.715 $Y=1.32 $X2=0 $Y2=0
cc_136 N_B_M1002_g N_A_185_367#_c_238_n 0.0131907f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_137 B N_A_185_367#_c_238_n 0.0206242f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_138 N_B_c_157_n N_A_185_367#_c_238_n 0.00154486f $X=1.715 $Y=1.32 $X2=0 $Y2=0
cc_139 N_B_M1008_g N_A_185_367#_c_233_n 6.75732e-19 $X=1.805 $Y=0.445 $X2=0
+ $Y2=0
cc_140 N_B_M1002_g N_A_185_367#_c_241_n 0.00218396f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_141 N_B_c_157_n N_A_185_367#_c_241_n 9.61836e-19 $X=1.715 $Y=1.32 $X2=0 $Y2=0
cc_142 B N_A_185_367#_c_234_n 0.00138433f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_143 N_B_M1002_g N_VPWR_c_313_n 0.00206274f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_144 N_B_M1002_g N_VPWR_c_314_n 5.18629e-19 $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_145 N_B_M1008_g N_VGND_c_366_n 0.00411659f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_146 B N_VGND_c_366_n 0.00970031f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_147 N_B_M1008_g N_VGND_c_368_n 0.00594837f $X=1.805 $Y=0.445 $X2=0 $Y2=0
cc_148 B N_VGND_c_368_n 0.00995888f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_149 B A_304_47# 0.00121399f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_150 N_C_M1001_g N_A_185_367#_M1000_g 0.0146661f $X=2.245 $Y=2.045 $X2=0 $Y2=0
cc_151 N_C_c_192_n N_A_185_367#_M1005_g 0.010454f $X=2.255 $Y=0.765 $X2=0 $Y2=0
cc_152 C N_A_185_367#_M1005_g 0.00214272f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_153 N_C_c_196_n N_A_185_367#_M1005_g 0.0121654f $X=2.255 $Y=0.93 $X2=0 $Y2=0
cc_154 N_C_M1001_g N_A_185_367#_c_240_n 0.015078f $X=2.245 $Y=2.045 $X2=0 $Y2=0
cc_155 N_C_c_194_n N_A_185_367#_c_240_n 0.00350111f $X=2.255 $Y=1.435 $X2=0
+ $Y2=0
cc_156 C N_A_185_367#_c_240_n 0.0125751f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_157 N_C_c_194_n N_A_185_367#_c_241_n 2.54824e-19 $X=2.255 $Y=1.435 $X2=0
+ $Y2=0
cc_158 C N_A_185_367#_c_241_n 0.00662052f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_159 N_C_M1001_g N_A_185_367#_c_234_n 0.00495113f $X=2.245 $Y=2.045 $X2=0
+ $Y2=0
cc_160 N_C_c_194_n N_A_185_367#_c_234_n 6.39891e-19 $X=2.255 $Y=1.435 $X2=0
+ $Y2=0
cc_161 C N_A_185_367#_c_234_n 0.00696351f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_162 N_C_M1001_g N_A_185_367#_c_235_n 0.00840202f $X=2.245 $Y=2.045 $X2=0
+ $Y2=0
cc_163 N_C_c_194_n N_A_185_367#_c_235_n 0.00589162f $X=2.255 $Y=1.435 $X2=0
+ $Y2=0
cc_164 N_C_M1001_g N_VPWR_c_314_n 0.00791814f $X=2.245 $Y=2.045 $X2=0 $Y2=0
cc_165 C N_VGND_M1009_d 0.00309749f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_166 N_C_c_192_n N_VGND_c_365_n 0.00669601f $X=2.255 $Y=0.765 $X2=0 $Y2=0
cc_167 C N_VGND_c_365_n 0.0563567f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_168 N_C_c_196_n N_VGND_c_365_n 0.00296605f $X=2.255 $Y=0.93 $X2=0 $Y2=0
cc_169 N_C_c_192_n N_VGND_c_366_n 0.00383378f $X=2.255 $Y=0.765 $X2=0 $Y2=0
cc_170 C N_VGND_c_366_n 0.00938312f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_171 N_C_c_196_n N_VGND_c_366_n 0.00183476f $X=2.255 $Y=0.93 $X2=0 $Y2=0
cc_172 N_C_c_192_n N_VGND_c_368_n 0.00594508f $X=2.255 $Y=0.765 $X2=0 $Y2=0
cc_173 C N_VGND_c_368_n 0.0103847f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_174 N_C_c_196_n N_VGND_c_368_n 0.00213938f $X=2.255 $Y=0.93 $X2=0 $Y2=0
cc_175 C A_376_47# 0.00227854f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_176 N_A_185_367#_c_238_n N_VPWR_M1004_d 0.00266818f $X=1.855 $Y=1.76 $X2=0
+ $Y2=0
cc_177 N_A_185_367#_c_240_n N_VPWR_M1001_d 0.00161579f $X=2.53 $Y=1.76 $X2=0
+ $Y2=0
cc_178 N_A_185_367#_c_234_n N_VPWR_M1001_d 0.00118436f $X=2.795 $Y=1.505 $X2=0
+ $Y2=0
cc_179 N_A_185_367#_c_238_n N_VPWR_c_313_n 0.020421f $X=1.855 $Y=1.76 $X2=0
+ $Y2=0
cc_180 N_A_185_367#_M1000_g N_VPWR_c_314_n 0.00675249f $X=2.77 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_185_367#_c_240_n N_VPWR_c_314_n 0.0141975f $X=2.53 $Y=1.76 $X2=0
+ $Y2=0
cc_182 N_A_185_367#_c_234_n N_VPWR_c_314_n 0.00952729f $X=2.795 $Y=1.505 $X2=0
+ $Y2=0
cc_183 N_A_185_367#_M1000_g N_VPWR_c_319_n 0.00585385f $X=2.77 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_185_367#_M1000_g N_VPWR_c_310_n 0.0129151f $X=2.77 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A_185_367#_M1005_g N_X_c_346_n 0.00277214f $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_186 N_A_185_367#_c_235_n X 0.00300488f $X=2.795 $Y=1.505 $X2=0 $Y2=0
cc_187 N_A_185_367#_M1000_g N_X_c_347_n 0.00343652f $X=2.77 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_185_367#_M1005_g N_X_c_347_n 0.00911749f $X=2.87 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A_185_367#_c_234_n N_X_c_347_n 0.0335744f $X=2.795 $Y=1.505 $X2=0 $Y2=0
cc_190 N_A_185_367#_c_235_n N_X_c_347_n 0.00807855f $X=2.795 $Y=1.505 $X2=0
+ $Y2=0
cc_191 N_A_185_367#_M1005_g N_VGND_c_365_n 0.0229989f $X=2.87 $Y=0.655 $X2=0
+ $Y2=0
cc_192 N_A_185_367#_c_240_n N_VGND_c_365_n 6.66316e-19 $X=2.53 $Y=1.76 $X2=0
+ $Y2=0
cc_193 N_A_185_367#_c_234_n N_VGND_c_365_n 0.0192802f $X=2.795 $Y=1.505 $X2=0
+ $Y2=0
cc_194 N_A_185_367#_c_235_n N_VGND_c_365_n 0.00124152f $X=2.795 $Y=1.505 $X2=0
+ $Y2=0
cc_195 N_A_185_367#_c_233_n N_VGND_c_366_n 0.0172608f $X=1.307 $Y=0.432 $X2=0
+ $Y2=0
cc_196 N_A_185_367#_M1005_g N_VGND_c_367_n 0.00486043f $X=2.87 $Y=0.655 $X2=0
+ $Y2=0
cc_197 N_A_185_367#_M1007_s N_VGND_c_368_n 0.0021695f $X=1.105 $Y=0.235 $X2=0
+ $Y2=0
cc_198 N_A_185_367#_M1005_g N_VGND_c_368_n 0.00919377f $X=2.87 $Y=0.655 $X2=0
+ $Y2=0
cc_199 N_A_185_367#_c_233_n N_VGND_c_368_n 0.0122689f $X=1.307 $Y=0.432 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_310_n N_X_M1000_d 0.00336915f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_319_n X 0.0271267f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_c_310_n X 0.0152789f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_203 N_X_c_346_n N_VGND_c_365_n 0.0319916f $X=3.132 $Y=1.095 $X2=0 $Y2=0
cc_204 N_X_c_345_n N_VGND_c_367_n 0.0196033f $X=3.085 $Y=0.42 $X2=0 $Y2=0
cc_205 N_X_M1005_d N_VGND_c_368_n 0.00371702f $X=2.945 $Y=0.235 $X2=0 $Y2=0
cc_206 N_X_c_345_n N_VGND_c_368_n 0.0110024f $X=3.085 $Y=0.42 $X2=0 $Y2=0
cc_207 N_VGND_c_368_n A_304_47# 0.00338427f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_208 N_VGND_c_368_n A_376_47# 0.00697595f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
