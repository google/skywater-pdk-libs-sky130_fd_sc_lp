* File: sky130_fd_sc_lp__or3b_2.spice
* Created: Fri Aug 28 11:24:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or3b_2.pex.spice"
.subckt sky130_fd_sc_lp__or3b_2  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_C_N_M1004_g N_A_33_131#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0952 AS=0.1113 PD=0.823333 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_195_21#_M1001_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1904 PD=1.12 PS=1.64667 NRD=0 NRS=9.636 M=1 R=5.6 SA=75000.5
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1001_d N_A_195_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=6.78 M=1 R=5.6 SA=75000.9
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1011 N_A_195_21#_M1011_d N_A_M1011_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0896 PD=0.7 PS=0.81 NRD=0 NRS=0 M=1 R=2.8 SA=75001.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g N_A_195_21#_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.0588 PD=0.72 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_195_21#_M1005_d N_A_33_131#_M1005_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.063 PD=1.37 PS=0.72 NRD=0 NRS=5.712 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_C_N_M1002_g N_A_33_131#_M1002_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=80.3169 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1002_d N_A_195_21#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75001 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_A_195_21#_M1010_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2898 AS=0.1764 PD=2.475 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 A_448_385# N_A_M1000_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0966 PD=0.63 PS=0.825 NRD=23.443 NRS=82.0702 M=1 R=2.8 SA=75001.6
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1008 A_520_385# N_B_M1008_g A_448_385# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_195_21#_M1009_d N_A_33_131#_M1009_g A_520_385# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75002.3 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_74 VPB 0 9.29714e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__or3b_2.pxi.spice"
*
.ends
*
*
