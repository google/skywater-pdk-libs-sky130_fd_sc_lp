* File: sky130_fd_sc_lp__nand4_m.spice
* Created: Fri Aug 28 10:51:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4_m.pex.spice"
.subckt sky130_fd_sc_lp__nand4_m  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1004 A_159_47# N_D_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1113 PD=0.66 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1005 A_237_47# N_C_M1005_g A_159_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=44.28 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1007 A_351_47# N_B_M1007_g A_237_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0882 PD=0.84 PS=0.84 NRD=44.28 NRS=44.28 M=1 R=2.8 SA=75001.1 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_351_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0882 PD=1.41 PS=0.84 NRD=5.712 NRS=44.28 M=1 R=2.8 SA=75001.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_D_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1806 AS=0.0588 PD=1.7 PS=0.7 NRD=77.3816 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.4 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__nand4_m.pxi.spice"
*
.ends
*
*
