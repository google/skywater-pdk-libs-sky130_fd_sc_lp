* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfsbp_lp CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 a_904_125# a_946_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1441_419# a_263_409# a_1519_125# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_531_113# a_263_409# a_476_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_2628_57# a_2383_57# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_263_409# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_1519_125# a_263_409# a_1621_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1621_125# a_1686_40# a_1716_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_712_419# a_946_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VPWR D a_145_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VPWR a_712_419# a_1441_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_712_419# a_476_409# a_904_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_2383_57# a_1519_125# a_2470_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_2200_57# a_1519_125# Q_N VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1249_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_2383_57# a_1519_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_1686_40# a_1519_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_373_113# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_884_419# a_946_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X18 VGND a_712_419# a_1441_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1686_40# a_1519_125# a_2042_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_263_409# a_476_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 a_263_409# CLK a_373_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_946_99# a_712_419# a_1249_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_145_409# a_476_409# a_712_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X24 a_2042_57# a_1519_125# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_2383_57# a_2628_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR SET_B a_1519_125# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 VGND a_1519_125# a_2200_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_946_99# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X29 VGND a_263_409# a_531_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VPWR a_1519_125# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X31 a_145_409# a_263_409# a_712_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_1441_125# a_476_409# a_1519_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_1716_66# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1719_419# a_1686_40# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X35 VPWR a_2383_57# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X36 a_712_419# a_263_409# a_884_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X37 a_2470_57# a_1519_125# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_1519_125# a_476_409# a_1719_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X39 a_110_57# D a_145_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VGND D a_110_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
