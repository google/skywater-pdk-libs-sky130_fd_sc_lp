* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfrbp_lp CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_2388_115# RESET_B a_2719_518# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_342_261# a_29_47# a_506_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_911_219# a_967_193# a_342_261# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_342_491# D a_342_261# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_2081_439# a_2388_115# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_2682_141# a_2168_439# a_2388_115# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_2340_141# a_2388_115# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_3684_53# a_3416_137# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_255_261# SCE a_342_261# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1303_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_2168_439# a_3233_357# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_3075_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VGND a_2168_439# a_3233_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VPWR RESET_B a_735_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VPWR a_2168_439# a_2523_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_2719_518# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_824_219# a_876_93# a_911_219# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_3233_47# a_2168_439# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_735_491# RESET_B a_342_261# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_2168_439# a_967_193# a_1147_490# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 a_1661_87# a_911_219# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_911_219# a_967_193# a_1020_491# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_116_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_3503_137# a_2168_439# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_342_261# a_876_93# a_911_219# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_1020_491# a_1147_490# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_342_261# D a_428_261# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_29_47# SCE a_116_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_2523_397# a_2168_439# a_2388_115# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_1147_490# a_911_219# a_1661_87# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 a_1147_490# a_876_93# a_2168_439# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X31 VGND a_3416_137# a_3684_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 a_967_193# CLK a_3075_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 a_500_261# SCD a_255_261# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_125_491# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 a_506_491# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 a_3416_137# a_2168_439# a_3503_137# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_1880_47# a_967_193# a_876_93# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 VPWR a_3416_137# a_3684_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 a_3684_367# a_3416_137# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X40 a_1147_490# a_911_219# a_1673_375# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X41 a_1673_375# a_911_219# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X42 a_3233_357# a_2168_439# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X43 a_3416_137# a_2168_439# a_3503_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X44 a_3503_367# a_2168_439# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X45 a_29_47# SCE a_125_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X46 VGND a_967_193# a_1880_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X47 a_428_261# a_29_47# a_500_261# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X48 VPWR RESET_B a_1375_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X49 a_1375_535# RESET_B a_911_219# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X50 VGND RESET_B a_2682_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X51 a_2081_439# a_876_93# a_2168_439# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X52 a_967_193# CLK a_3075_357# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X53 a_3075_357# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X54 a_2168_439# a_967_193# a_2340_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X55 VPWR a_967_193# a_1870_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X56 VGND RESET_B a_500_261# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X57 a_824_219# a_1147_490# a_1303_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X58 VPWR SCE a_342_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X59 a_1870_367# a_967_193# a_876_93# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
