* File: sky130_fd_sc_lp__xnor2_2.spice
* Created: Fri Aug 28 11:35:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xnor2_2.pex.spice"
.subckt sky130_fd_sc_lp__xnor2_2  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_27_47#_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2436 AS=0.2226 PD=1.42 PS=2.21 NRD=4.284 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1007_d N_A_M1011_g N_A_27_47#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2436 AS=0.1176 PD=1.42 PS=1.12 NRD=38.568 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1002 N_A_27_47#_M1011_s N_B_M1002_g N_A_162_367#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.3
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1018 N_A_27_47#_M1018_d N_B_M1018_g N_A_162_367#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2814 AS=0.1176 PD=2.35 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6
+ SA=75001.8 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A_M1008_g N_A_555_65#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1008_d N_A_M1009_g N_A_555_65#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1016 N_A_555_65#_M1009_s N_B_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2982 PD=1.12 PS=1.55 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1 SB=75002
+ A=0.126 P=1.98 MULT=1
MM1017 N_A_555_65#_M1017_d N_B_M1017_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2982 PD=1.12 PS=1.55 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_162_367#_M1003_g N_A_555_65#_M1017_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1012 N_Y_M1003_d N_A_162_367#_M1012_g N_A_555_65#_M1012_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2814 PD=1.12 PS=2.35 NRD=0 NRS=9.996 M=1 R=5.6
+ SA=75002.8 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_A_162_367#_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4788 AS=0.1764 PD=3.28 PS=1.54 NRD=4.9447 NRS=0 M=1 R=8.4 SA=75000.3
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1019_d N_A_M1019_g N_A_162_367#_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75000.7
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1005 N_A_162_367#_M1005_d N_B_M1005_g N_VPWR_M1019_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75001.2
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1015 N_A_162_367#_M1005_d N_B_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.27405 PD=1.54 PS=1.695 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75001.6
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1015_s N_A_M1000_g N_A_545_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.27405 AS=0.1764 PD=1.695 PS=1.54 NRD=11.7215 NRS=0 M=1 R=8.4 SA=75002.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g N_A_545_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_A_545_367#_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_B_M1006_g N_A_545_367#_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1006_d N_A_162_367#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_Y_M1013_d N_A_162_367#_M1013_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3463 P=16.97
*
.include "sky130_fd_sc_lp__xnor2_2.pxi.spice"
*
.ends
*
*
