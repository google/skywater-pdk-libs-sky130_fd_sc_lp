# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__isolatch_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__isolatch_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.255000 0.835000 1.780000 ;
        RECT 0.125000 1.780000 0.295000 2.185000 ;
        RECT 0.125000 2.185000 0.585000 2.515000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.459700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.450000 0.440000 7.085000 2.955000 ;
    END
  END Q
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.675000 7.130000 2.945000 ;
    END
  END KAPWR
  PIN SLEEP_B
    ANTENNAGATEAREA  0.222000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.355000 1.450000 4.685000 1.780000 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.130000  2.685000 0.460000 3.245000 ;
      RECT 0.160000  0.345000 0.410000 0.915000 ;
      RECT 0.160000  0.915000 1.355000 1.085000 ;
      RECT 0.590000  0.085000 0.920000 0.745000 ;
      RECT 1.155000  1.950000 1.515000 2.120000 ;
      RECT 1.155000  2.120000 1.325000 2.905000 ;
      RECT 1.155000  2.905000 2.345000 3.075000 ;
      RECT 1.185000  1.085000 1.355000 1.670000 ;
      RECT 1.185000  1.670000 1.515000 1.950000 ;
      RECT 1.495000  2.290000 1.855000 2.735000 ;
      RECT 1.575000  0.345000 1.970000 0.555000 ;
      RECT 1.575000  0.555000 2.585000 0.725000 ;
      RECT 1.575000  0.725000 1.745000 1.330000 ;
      RECT 1.575000  1.330000 1.855000 1.500000 ;
      RECT 1.685000  1.500000 1.855000 2.290000 ;
      RECT 1.915000  0.895000 2.245000 1.160000 ;
      RECT 2.075000  1.160000 2.245000 1.285000 ;
      RECT 2.075000  1.285000 3.980000 1.445000 ;
      RECT 2.075000  1.445000 4.185000 1.615000 ;
      RECT 2.175000  1.785000 3.295000 1.955000 ;
      RECT 2.175000  1.955000 2.345000 2.905000 ;
      RECT 2.415000  0.725000 2.585000 0.945000 ;
      RECT 2.415000  0.945000 3.560000 1.115000 ;
      RECT 2.515000  2.125000 2.845000 3.075000 ;
      RECT 2.970000  0.085000 3.220000 0.775000 ;
      RECT 3.045000  1.955000 3.295000 3.075000 ;
      RECT 3.390000  0.255000 4.320000 0.425000 ;
      RECT 3.390000  0.425000 3.560000 0.945000 ;
      RECT 3.515000  1.785000 3.845000 2.905000 ;
      RECT 3.515000  2.905000 4.605000 3.075000 ;
      RECT 3.730000  0.595000 3.980000 1.285000 ;
      RECT 4.015000  1.615000 4.185000 2.055000 ;
      RECT 4.015000  2.055000 4.265000 2.735000 ;
      RECT 4.150000  0.425000 4.320000 1.075000 ;
      RECT 4.150000  1.075000 5.225000 1.245000 ;
      RECT 4.435000  1.950000 5.665000 2.120000 ;
      RECT 4.435000  2.120000 4.605000 2.905000 ;
      RECT 4.600000  0.085000 4.850000 0.905000 ;
      RECT 4.775000  2.290000 5.155000 2.905000 ;
      RECT 4.895000  1.245000 5.225000 1.745000 ;
      RECT 5.335000  1.915000 5.665000 1.950000 ;
      RECT 5.335000  2.120000 5.665000 2.955000 ;
      RECT 5.460000  0.445000 5.665000 0.775000 ;
      RECT 5.495000  0.775000 5.665000 1.915000 ;
      RECT 5.865000  1.915000 6.195000 2.955000 ;
      RECT 5.950000  0.085000 6.280000 1.325000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  2.735000 2.725000 2.905000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  2.735000 5.125000 2.905000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  2.735000 6.085000 2.905000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_lp__isolatch_lp
END LIBRARY
