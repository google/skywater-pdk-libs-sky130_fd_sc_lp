* File: sky130_fd_sc_lp__dfstp_1.pxi.spice
* Created: Wed Sep  2 09:44:20 2020
* 
x_PM_SKY130_FD_SC_LP__DFSTP_1%CLK N_CLK_c_216_n N_CLK_c_221_n N_CLK_M1012_g
+ N_CLK_c_217_n N_CLK_M1017_g N_CLK_c_222_n CLK CLK N_CLK_c_219_n
+ PM_SKY130_FD_SC_LP__DFSTP_1%CLK
x_PM_SKY130_FD_SC_LP__DFSTP_1%D N_D_c_261_n N_D_M1005_g N_D_c_264_n N_D_M1009_g
+ N_D_c_262_n N_D_c_265_n D N_D_c_263_n PM_SKY130_FD_SC_LP__DFSTP_1%D
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_202_463# N_A_202_463#_M1018_d
+ N_A_202_463#_M1024_d N_A_202_463#_M1001_g N_A_202_463#_c_309_n
+ N_A_202_463#_M1030_g N_A_202_463#_M1013_g N_A_202_463#_M1031_g
+ N_A_202_463#_c_312_n N_A_202_463#_c_313_n N_A_202_463#_c_314_n
+ N_A_202_463#_c_315_n N_A_202_463#_c_330_n N_A_202_463#_c_316_n
+ N_A_202_463#_c_317_n N_A_202_463#_c_318_n N_A_202_463#_c_319_n
+ N_A_202_463#_c_334_n N_A_202_463#_c_320_n N_A_202_463#_c_321_n
+ N_A_202_463#_c_322_n PM_SKY130_FD_SC_LP__DFSTP_1%A_202_463#
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_614_93# N_A_614_93#_M1027_s N_A_614_93#_M1003_d
+ N_A_614_93#_M1022_g N_A_614_93#_M1023_g N_A_614_93#_c_486_n
+ N_A_614_93#_c_487_n N_A_614_93#_c_479_n N_A_614_93#_c_488_n
+ N_A_614_93#_c_480_n N_A_614_93#_c_481_n N_A_614_93#_c_482_n
+ N_A_614_93#_c_500_p N_A_614_93#_c_483_n N_A_614_93#_c_484_n
+ PM_SKY130_FD_SC_LP__DFSTP_1%A_614_93#
x_PM_SKY130_FD_SC_LP__DFSTP_1%SET_B N_SET_B_M1025_g N_SET_B_M1016_g
+ N_SET_B_M1008_g N_SET_B_M1021_g N_SET_B_c_566_n N_SET_B_c_567_n
+ N_SET_B_c_568_n N_SET_B_c_569_n N_SET_B_c_577_n N_SET_B_c_578_n SET_B SET_B
+ SET_B SET_B N_SET_B_c_571_n N_SET_B_c_572_n N_SET_B_c_581_n SET_B
+ N_SET_B_c_573_n PM_SKY130_FD_SC_LP__DFSTP_1%SET_B
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_486_119# N_A_486_119#_M1028_d
+ N_A_486_119#_M1001_d N_A_486_119#_M1003_g N_A_486_119#_M1027_g
+ N_A_486_119#_c_696_n N_A_486_119#_c_697_n N_A_486_119#_M1007_g
+ N_A_486_119#_c_699_n N_A_486_119#_c_700_n N_A_486_119#_c_701_n
+ N_A_486_119#_c_702_n N_A_486_119#_M1029_g N_A_486_119#_c_703_n
+ N_A_486_119#_c_730_n N_A_486_119#_c_704_n N_A_486_119#_c_709_n
+ N_A_486_119#_c_705_n N_A_486_119#_c_739_n N_A_486_119#_c_711_n
+ N_A_486_119#_c_706_n PM_SKY130_FD_SC_LP__DFSTP_1%A_486_119#
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_33_463# N_A_33_463#_M1017_s N_A_33_463#_M1012_s
+ N_A_33_463#_M1024_g N_A_33_463#_M1018_g N_A_33_463#_c_854_n
+ N_A_33_463#_c_855_n N_A_33_463#_c_844_n N_A_33_463#_c_845_n
+ N_A_33_463#_M1028_g N_A_33_463#_M1020_g N_A_33_463#_c_857_n
+ N_A_33_463#_M1004_g N_A_33_463#_M1014_g N_A_33_463#_c_860_n
+ N_A_33_463#_c_861_n N_A_33_463#_c_848_n N_A_33_463#_c_862_n
+ N_A_33_463#_c_849_n N_A_33_463#_c_850_n N_A_33_463#_c_851_n
+ N_A_33_463#_c_852_n PM_SKY130_FD_SC_LP__DFSTP_1%A_33_463#
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_1329_65# N_A_1329_65#_M1019_d
+ N_A_1329_65#_M1010_d N_A_1329_65#_M1015_g N_A_1329_65#_c_985_n
+ N_A_1329_65#_c_986_n N_A_1329_65#_c_987_n N_A_1329_65#_M1002_g
+ N_A_1329_65#_c_989_n N_A_1329_65#_c_990_n N_A_1329_65#_c_991_n
+ N_A_1329_65#_c_981_n N_A_1329_65#_c_982_n N_A_1329_65#_c_993_n
+ N_A_1329_65#_c_983_n PM_SKY130_FD_SC_LP__DFSTP_1%A_1329_65#
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_1175_417# N_A_1175_417#_M1031_d
+ N_A_1175_417#_M1013_d N_A_1175_417#_M1021_d N_A_1175_417#_c_1069_n
+ N_A_1175_417#_M1019_g N_A_1175_417#_c_1070_n N_A_1175_417#_c_1071_n
+ N_A_1175_417#_M1010_g N_A_1175_417#_c_1073_n N_A_1175_417#_c_1074_n
+ N_A_1175_417#_M1011_g N_A_1175_417#_M1026_g N_A_1175_417#_c_1076_n
+ N_A_1175_417#_c_1077_n N_A_1175_417#_c_1078_n N_A_1175_417#_c_1079_n
+ N_A_1175_417#_c_1080_n N_A_1175_417#_c_1086_n N_A_1175_417#_c_1081_n
+ N_A_1175_417#_c_1088_n N_A_1175_417#_c_1106_n N_A_1175_417#_c_1108_n
+ N_A_1175_417#_c_1082_n N_A_1175_417#_c_1083_n N_A_1175_417#_c_1089_n
+ PM_SKY130_FD_SC_LP__DFSTP_1%A_1175_417#
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_1832_131# N_A_1832_131#_M1011_s
+ N_A_1832_131#_M1026_s N_A_1832_131#_M1000_g N_A_1832_131#_M1006_g
+ N_A_1832_131#_c_1188_n N_A_1832_131#_c_1193_n N_A_1832_131#_c_1189_n
+ N_A_1832_131#_c_1190_n N_A_1832_131#_c_1191_n
+ PM_SKY130_FD_SC_LP__DFSTP_1%A_1832_131#
x_PM_SKY130_FD_SC_LP__DFSTP_1%VPWR N_VPWR_M1012_d N_VPWR_M1009_s N_VPWR_M1023_d
+ N_VPWR_M1025_d N_VPWR_M1002_d N_VPWR_M1010_s N_VPWR_M1026_d N_VPWR_c_1229_n
+ N_VPWR_c_1230_n N_VPWR_c_1231_n N_VPWR_c_1232_n N_VPWR_c_1233_n
+ N_VPWR_c_1234_n N_VPWR_c_1235_n N_VPWR_c_1236_n N_VPWR_c_1237_n
+ N_VPWR_c_1238_n N_VPWR_c_1239_n N_VPWR_c_1240_n N_VPWR_c_1241_n VPWR
+ N_VPWR_c_1242_n N_VPWR_c_1243_n N_VPWR_c_1244_n N_VPWR_c_1245_n
+ N_VPWR_c_1246_n N_VPWR_c_1247_n N_VPWR_c_1228_n N_VPWR_c_1249_n
+ N_VPWR_c_1250_n N_VPWR_c_1251_n N_VPWR_c_1252_n N_VPWR_c_1253_n
+ PM_SKY130_FD_SC_LP__DFSTP_1%VPWR
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_400_119# N_A_400_119#_M1005_d
+ N_A_400_119#_M1009_d N_A_400_119#_c_1363_n N_A_400_119#_c_1366_n
+ N_A_400_119#_c_1364_n N_A_400_119#_c_1365_n N_A_400_119#_c_1368_n
+ PM_SKY130_FD_SC_LP__DFSTP_1%A_400_119#
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_985_379# N_A_985_379#_M1007_d
+ N_A_985_379#_M1004_d N_A_985_379#_c_1414_n N_A_985_379#_c_1415_n
+ N_A_985_379#_c_1416_n PM_SKY130_FD_SC_LP__DFSTP_1%A_985_379#
x_PM_SKY130_FD_SC_LP__DFSTP_1%A_1092_417# N_A_1092_417#_M1013_s
+ N_A_1092_417#_M1002_s N_A_1092_417#_c_1440_n N_A_1092_417#_c_1441_n
+ N_A_1092_417#_c_1442_n N_A_1092_417#_c_1443_n
+ PM_SKY130_FD_SC_LP__DFSTP_1%A_1092_417#
x_PM_SKY130_FD_SC_LP__DFSTP_1%Q N_Q_M1000_d N_Q_M1006_d N_Q_c_1466_n
+ N_Q_c_1467_n Q Q Q Q Q PM_SKY130_FD_SC_LP__DFSTP_1%Q
x_PM_SKY130_FD_SC_LP__DFSTP_1%VGND N_VGND_M1017_d N_VGND_M1005_s N_VGND_M1022_d
+ N_VGND_M1016_d N_VGND_M1008_d N_VGND_M1011_d N_VGND_c_1483_n N_VGND_c_1484_n
+ N_VGND_c_1485_n N_VGND_c_1486_n N_VGND_c_1487_n VGND N_VGND_c_1488_n
+ N_VGND_c_1489_n N_VGND_c_1490_n N_VGND_c_1491_n N_VGND_c_1492_n
+ N_VGND_c_1493_n N_VGND_c_1494_n N_VGND_c_1495_n N_VGND_c_1496_n
+ N_VGND_c_1497_n N_VGND_c_1498_n N_VGND_c_1499_n N_VGND_c_1500_n
+ PM_SKY130_FD_SC_LP__DFSTP_1%VGND
cc_1 VNB N_CLK_c_216_n 0.0252316f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=2.05
cc_2 VNB N_CLK_c_217_n 0.0225381f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.91
cc_3 VNB CLK 0.0108088f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_4 VNB N_CLK_c_219_n 0.0510096f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.075
cc_5 VNB N_D_c_261_n 0.0167208f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=1.24
cc_6 VNB N_D_c_262_n 0.0375567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_D_c_263_n 0.0271126f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.075
cc_8 VNB N_A_202_463#_c_309_n 0.01393f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.125
cc_9 VNB N_A_202_463#_M1030_g 0.0368011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_202_463#_M1031_g 0.0393882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_202_463#_c_312_n 0.0160388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_202_463#_c_313_n 0.00580056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_202_463#_c_314_n 0.0237866f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.075
cc_14 VNB N_A_202_463#_c_315_n 0.0147454f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.295
cc_15 VNB N_A_202_463#_c_316_n 0.00182506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_202_463#_c_317_n 2.79276e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_202_463#_c_318_n 0.00173158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_202_463#_c_319_n 0.0344449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_202_463#_c_320_n 0.00830897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_202_463#_c_321_n 0.00980386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_202_463#_c_322_n 0.0134342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_614_93#_c_479_n 0.0151301f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.075
cc_23 VNB N_A_614_93#_c_480_n 0.0125424f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.075
cc_24 VNB N_A_614_93#_c_481_n 5.59107e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_614_93#_c_482_n 0.0353664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_614_93#_c_483_n 0.0181071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_614_93#_c_484_n 0.0102077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_SET_B_M1008_g 0.030722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_SET_B_c_566_n 0.00873866f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=1.075
cc_30 VNB N_SET_B_c_567_n 0.00522014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_SET_B_c_568_n 0.00402841f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.075
cc_32 VNB N_SET_B_c_569_n 0.0322542f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.075
cc_33 VNB SET_B 0.0066768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_SET_B_c_571_n 0.0185953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_SET_B_c_572_n 0.072208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_SET_B_c_573_n 0.00260165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_486_119#_M1003_g 0.00241197f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=2.125
cc_38 VNB N_A_486_119#_M1027_g 0.0496073f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_39 VNB N_A_486_119#_c_696_n 0.0271047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_486_119#_c_697_n 0.0559669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_486_119#_M1007_g 0.0111163f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.075
cc_42 VNB N_A_486_119#_c_699_n 0.0145785f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.075
cc_43 VNB N_A_486_119#_c_700_n 0.0230123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_486_119#_c_701_n 0.00946809f $X=-0.19 $Y=-0.245 $X2=0.657
+ $Y2=0.925
cc_45 VNB N_A_486_119#_c_702_n 0.0186994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_486_119#_c_703_n 0.019743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_486_119#_c_704_n 0.0035226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_486_119#_c_705_n 0.0050692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_486_119#_c_706_n 0.0014183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_33_463#_M1018_g 0.0475271f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_51 VNB N_A_33_463#_c_844_n 0.102594f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=1.075
cc_52 VNB N_A_33_463#_c_845_n 0.012349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_33_463#_M1028_g 0.0362599f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.075
cc_54 VNB N_A_33_463#_M1014_g 0.0463511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_33_463#_c_848_n 0.0320258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_33_463#_c_849_n 0.00112671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_33_463#_c_850_n 0.0131264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_33_463#_c_851_n 0.00515535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_33_463#_c_852_n 0.0257213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1329_65#_M1015_g 0.0437087f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=2.125
cc_61 VNB N_A_1329_65#_c_981_n 0.0165747f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.075
cc_62 VNB N_A_1329_65#_c_982_n 0.0178958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1329_65#_c_983_n 0.00279198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1175_417#_c_1069_n 0.015011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1175_417#_c_1070_n 0.0552969f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=0.84
cc_66 VNB N_A_1175_417#_c_1071_n 0.0116398f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_67 VNB N_A_1175_417#_M1010_g 0.00578958f $X=-0.19 $Y=-0.245 $X2=0.22
+ $Y2=1.075
cc_68 VNB N_A_1175_417#_c_1073_n 0.0584899f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.075
cc_69 VNB N_A_1175_417#_c_1074_n 0.0187521f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.075
cc_70 VNB N_A_1175_417#_M1026_g 0.0174971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1175_417#_c_1076_n 0.0231177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1175_417#_c_1077_n 0.00558097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1175_417#_c_1078_n 0.0025412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1175_417#_c_1079_n 0.0282884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1175_417#_c_1080_n 0.00361575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1175_417#_c_1081_n 9.94938e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1175_417#_c_1082_n 0.0217566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1175_417#_c_1083_n 0.0725222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1832_131#_M1000_g 0.0301963f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=2.125
cc_80 VNB N_A_1832_131#_M1006_g 5.54595e-19 $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=0.84
cc_81 VNB N_A_1832_131#_c_1188_n 0.00584082f $X=-0.19 $Y=-0.245 $X2=0.22
+ $Y2=1.075
cc_82 VNB N_A_1832_131#_c_1189_n 0.00538894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1832_131#_c_1190_n 0.0361397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1832_131#_c_1191_n 0.00294665f $X=-0.19 $Y=-0.245 $X2=0.657
+ $Y2=1.295
cc_85 VNB N_VPWR_c_1228_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_400_119#_c_1363_n 0.0045616f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=2.125
cc_87 VNB N_A_400_119#_c_1364_n 0.00340127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_400_119#_c_1365_n 0.0128375f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.075
cc_89 VNB N_Q_c_1466_n 0.0284879f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=2.125
cc_90 VNB N_Q_c_1467_n 0.0109607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB Q 0.0298675f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_92 VNB N_VGND_c_1483_n 0.00839338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1484_n 0.0133554f $X=-0.19 $Y=-0.245 $X2=0.657 $Y2=1.075
cc_94 VNB N_VGND_c_1485_n 0.0238047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1486_n 0.0107514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1487_n 0.015784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1488_n 0.0183897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1489_n 0.0415939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1490_n 0.0276682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1491_n 0.0494317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1492_n 0.0554222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1493_n 0.0187942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1494_n 0.564601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1495_n 0.024227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1496_n 0.00399507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1497_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1498_n 0.0178816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1499_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1500_n 0.00682834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VPB N_CLK_c_216_n 0.0225386f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=2.05
cc_111 VPB N_CLK_c_221_n 0.0209835f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.2
cc_112 VPB N_CLK_c_222_n 0.0303237f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.125
cc_113 VPB N_D_c_264_n 0.0170364f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.635
cc_114 VPB N_D_c_265_n 0.0391555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB D 0.0049849f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.075
cc_116 VPB N_D_c_263_n 0.0278923f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.075
cc_117 VPB N_A_202_463#_M1001_g 0.0372381f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=2.125
cc_118 VPB N_A_202_463#_c_309_n 0.0113748f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.125
cc_119 VPB N_A_202_463#_M1013_g 0.0417121f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.075
cc_120 VPB N_A_202_463#_c_312_n 0.0186533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_202_463#_c_313_n 0.00714039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_202_463#_c_314_n 0.00938642f $X=-0.19 $Y=1.655 $X2=0.657
+ $Y2=1.075
cc_123 VPB N_A_202_463#_c_315_n 7.94824e-19 $X=-0.19 $Y=1.655 $X2=0.657
+ $Y2=1.295
cc_124 VPB N_A_202_463#_c_330_n 0.016474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_202_463#_c_316_n 0.00476375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_202_463#_c_317_n 0.00428027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_202_463#_c_318_n 0.00258928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_614_93#_M1023_g 0.0187654f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_129 VPB N_A_614_93#_c_486_n 0.0103283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_614_93#_c_487_n 0.0321733f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.075
cc_131 VPB N_A_614_93#_c_488_n 0.00145834f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=0.925
cc_132 VPB N_A_614_93#_c_484_n 0.0105138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_SET_B_M1025_g 0.0202843f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.2
cc_134 VPB N_SET_B_M1021_g 0.0400975f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_135 VPB N_SET_B_c_566_n 0.00230808f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.075
cc_136 VPB N_SET_B_c_577_n 0.00472475f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=0.925
cc_137 VPB N_SET_B_c_578_n 0.0347167f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=1.075
cc_138 VPB SET_B 0.0069238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_SET_B_c_572_n 0.0393116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_SET_B_c_581_n 0.0204928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_SET_B_c_573_n 0.0032204f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_486_119#_M1003_g 0.0419852f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=2.125
cc_143 VPB N_A_486_119#_M1007_g 0.0294797f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.075
cc_144 VPB N_A_486_119#_c_709_n 0.00997659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_486_119#_c_705_n 0.00971681f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_486_119#_c_711_n 3.95607e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_486_119#_c_706_n 0.00187711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_33_463#_M1024_g 0.0381516f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_33_463#_c_854_n 0.132012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_33_463#_c_855_n 0.0115084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_33_463#_M1020_g 0.0338551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_33_463#_c_857_n 0.254061f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=1.075
cc_153 VPB N_A_33_463#_M1004_g 0.015989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_33_463#_M1014_g 0.00743671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_33_463#_c_860_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_33_463#_c_861_n 0.00959926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_33_463#_c_862_n 0.0508794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_33_463#_c_849_n 0.00147517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_33_463#_c_851_n 0.00631276f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_33_463#_c_852_n 0.0226968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_1329_65#_M1015_g 0.00935737f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=2.125
cc_162 VPB N_A_1329_65#_c_985_n 0.0638342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_1329_65#_c_986_n 0.0210735f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_164 VPB N_A_1329_65#_c_987_n 0.0104278f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_165 VPB N_A_1329_65#_M1002_g 0.027265f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.075
cc_166 VPB N_A_1329_65#_c_989_n 0.102795f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.075
cc_167 VPB N_A_1329_65#_c_990_n 0.0232702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_1329_65#_c_991_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_1329_65#_c_982_n 0.0250014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_1329_65#_c_993_n 0.0700811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_1175_417#_M1010_g 0.0255919f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.075
cc_172 VPB N_A_1175_417#_M1026_g 0.0242343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_1175_417#_c_1086_n 0.0159526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_1175_417#_c_1081_n 0.00554859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_1175_417#_c_1088_n 5.51325e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_1175_417#_c_1089_n 0.00534719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_1832_131#_M1006_g 0.0261028f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_178 VPB N_A_1832_131#_c_1193_n 0.0157411f $X=-0.19 $Y=1.655 $X2=0.525
+ $Y2=1.075
cc_179 VPB N_VPWR_c_1229_n 0.00535543f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=0.925
cc_180 VPB N_VPWR_c_1230_n 0.0194684f $X=-0.19 $Y=1.655 $X2=0.657 $Y2=1.295
cc_181 VPB N_VPWR_c_1231_n 0.014895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1232_n 0.00235552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1233_n 0.0151625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1234_n 0.00854941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1235_n 0.0192756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1236_n 0.0156651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1237_n 0.0393344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1238_n 0.00376942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1239_n 0.0666457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1240_n 0.00223798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1241_n 0.00194187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1242_n 0.0176864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1243_n 0.019164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1244_n 0.0186716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1245_n 0.016117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1246_n 0.0306926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1247_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1228_n 0.0679329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1249_n 0.00469783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1250_n 0.00396918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1251_n 0.00590013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1252_n 0.00223798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1253_n 0.00789746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_400_119#_c_1366_n 0.00313824f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=0.84
cc_205 VPB N_A_400_119#_c_1364_n 0.00286824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_400_119#_c_1368_n 0.00815972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_985_379#_c_1414_n 0.0124106f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=2.125
cc_208 VPB N_A_985_379#_c_1415_n 0.00329908f $X=-0.19 $Y=1.655 $X2=0.505
+ $Y2=2.125
cc_209 VPB N_A_985_379#_c_1416_n 0.027781f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_210 VPB N_A_1092_417#_c_1440_n 0.00358247f $X=-0.19 $Y=1.655 $X2=0.22
+ $Y2=2.125
cc_211 VPB N_A_1092_417#_c_1441_n 0.00411073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_1092_417#_c_1442_n 0.00148549f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.21
cc_213 VPB N_A_1092_417#_c_1443_n 0.00364126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB Q 0.0576472f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_215 CLK N_A_202_463#_c_334_n 0.00163262f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_216 N_CLK_c_217_n N_A_202_463#_c_322_n 8.59152e-19 $X=0.545 $Y=0.91 $X2=0
+ $Y2=0
cc_217 CLK N_A_202_463#_c_322_n 0.0426089f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_218 N_CLK_c_219_n N_A_202_463#_c_322_n 2.35324e-19 $X=0.545 $Y=1.075 $X2=0
+ $Y2=0
cc_219 N_CLK_c_216_n N_A_33_463#_M1024_g 0.00228702f $X=0.22 $Y=2.05 $X2=0 $Y2=0
cc_220 N_CLK_c_222_n N_A_33_463#_M1024_g 0.00870166f $X=0.505 $Y=2.125 $X2=0
+ $Y2=0
cc_221 N_CLK_c_216_n N_A_33_463#_M1018_g 0.00244705f $X=0.22 $Y=2.05 $X2=0 $Y2=0
cc_222 CLK N_A_33_463#_M1018_g 0.00576717f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_223 N_CLK_c_219_n N_A_33_463#_M1018_g 0.0193178f $X=0.545 $Y=1.075 $X2=0
+ $Y2=0
cc_224 N_CLK_c_221_n N_A_33_463#_c_855_n 0.00870166f $X=0.505 $Y=2.2 $X2=0 $Y2=0
cc_225 N_CLK_c_217_n N_A_33_463#_c_845_n 0.0133852f $X=0.545 $Y=0.91 $X2=0 $Y2=0
cc_226 N_CLK_c_216_n N_A_33_463#_c_848_n 0.012404f $X=0.22 $Y=2.05 $X2=0 $Y2=0
cc_227 N_CLK_c_217_n N_A_33_463#_c_848_n 0.00473144f $X=0.545 $Y=0.91 $X2=0
+ $Y2=0
cc_228 CLK N_A_33_463#_c_848_n 0.0395466f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_229 N_CLK_c_219_n N_A_33_463#_c_848_n 0.0152336f $X=0.545 $Y=1.075 $X2=0
+ $Y2=0
cc_230 N_CLK_c_216_n N_A_33_463#_c_862_n 0.00862274f $X=0.22 $Y=2.05 $X2=0 $Y2=0
cc_231 N_CLK_c_221_n N_A_33_463#_c_862_n 0.0035646f $X=0.505 $Y=2.2 $X2=0 $Y2=0
cc_232 N_CLK_c_222_n N_A_33_463#_c_862_n 0.0169562f $X=0.505 $Y=2.125 $X2=0
+ $Y2=0
cc_233 N_CLK_c_222_n N_A_33_463#_c_849_n 0.00564902f $X=0.505 $Y=2.125 $X2=0
+ $Y2=0
cc_234 CLK N_A_33_463#_c_849_n 0.034841f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_235 N_CLK_c_219_n N_A_33_463#_c_849_n 0.00211969f $X=0.545 $Y=1.075 $X2=0
+ $Y2=0
cc_236 N_CLK_c_217_n N_A_33_463#_c_850_n 0.0034398f $X=0.545 $Y=0.91 $X2=0 $Y2=0
cc_237 CLK N_A_33_463#_c_850_n 0.00309811f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_238 N_CLK_c_219_n N_A_33_463#_c_850_n 0.00676674f $X=0.545 $Y=1.075 $X2=0
+ $Y2=0
cc_239 N_CLK_c_216_n N_A_33_463#_c_851_n 0.0116095f $X=0.22 $Y=2.05 $X2=0 $Y2=0
cc_240 N_CLK_c_219_n N_A_33_463#_c_851_n 0.00378702f $X=0.545 $Y=1.075 $X2=0
+ $Y2=0
cc_241 N_CLK_c_216_n N_A_33_463#_c_852_n 0.0183218f $X=0.22 $Y=2.05 $X2=0 $Y2=0
cc_242 N_CLK_c_222_n N_A_33_463#_c_852_n 0.00273223f $X=0.505 $Y=2.125 $X2=0
+ $Y2=0
cc_243 CLK N_A_33_463#_c_852_n 0.00609563f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_244 N_CLK_c_219_n N_A_33_463#_c_852_n 0.00809438f $X=0.545 $Y=1.075 $X2=0
+ $Y2=0
cc_245 N_CLK_c_221_n N_VPWR_c_1229_n 0.0137999f $X=0.505 $Y=2.2 $X2=0 $Y2=0
cc_246 N_CLK_c_221_n N_VPWR_c_1242_n 0.00410286f $X=0.505 $Y=2.2 $X2=0 $Y2=0
cc_247 N_CLK_c_221_n N_VPWR_c_1228_n 0.00493487f $X=0.505 $Y=2.2 $X2=0 $Y2=0
cc_248 N_CLK_c_217_n N_VGND_c_1483_n 0.00320103f $X=0.545 $Y=0.91 $X2=0 $Y2=0
cc_249 CLK N_VGND_c_1483_n 0.0160352f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_250 N_CLK_c_217_n N_VGND_c_1494_n 0.00450325f $X=0.545 $Y=0.91 $X2=0 $Y2=0
cc_251 CLK N_VGND_c_1494_n 0.00682803f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_252 N_CLK_c_217_n N_VGND_c_1495_n 0.00434051f $X=0.545 $Y=0.91 $X2=0 $Y2=0
cc_253 N_D_c_265_n N_A_202_463#_M1001_g 0.0175102f $X=1.975 $Y=2.13 $X2=0 $Y2=0
cc_254 D N_A_202_463#_M1001_g 0.00196012f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_255 N_D_c_263_n N_A_202_463#_M1001_g 0.00192756f $X=1.6 $Y=1.99 $X2=0 $Y2=0
cc_256 N_D_c_262_n N_A_202_463#_M1030_g 0.00150115f $X=1.925 $Y=1.2 $X2=0 $Y2=0
cc_257 N_D_c_262_n N_A_202_463#_c_312_n 0.00155301f $X=1.925 $Y=1.2 $X2=0 $Y2=0
cc_258 N_D_c_265_n N_A_202_463#_c_312_n 0.00521921f $X=1.975 $Y=2.13 $X2=0 $Y2=0
cc_259 N_D_c_263_n N_A_202_463#_c_312_n 0.0223588f $X=1.6 $Y=1.99 $X2=0 $Y2=0
cc_260 N_D_c_264_n N_A_202_463#_c_330_n 0.00395451f $X=1.975 $Y=2.205 $X2=0
+ $Y2=0
cc_261 N_D_c_265_n N_A_202_463#_c_330_n 3.92145e-19 $X=1.975 $Y=2.13 $X2=0 $Y2=0
cc_262 D N_A_202_463#_c_330_n 0.0247977f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_263 N_D_c_263_n N_A_202_463#_c_330_n 0.00524982f $X=1.6 $Y=1.99 $X2=0 $Y2=0
cc_264 N_D_c_262_n N_A_202_463#_c_316_n 0.00550011f $X=1.925 $Y=1.2 $X2=0 $Y2=0
cc_265 N_D_c_265_n N_A_202_463#_c_316_n 0.00426427f $X=1.975 $Y=2.13 $X2=0 $Y2=0
cc_266 D N_A_202_463#_c_316_n 0.028026f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_267 N_D_c_263_n N_A_202_463#_c_316_n 0.0197212f $X=1.6 $Y=1.99 $X2=0 $Y2=0
cc_268 N_D_c_265_n N_A_202_463#_c_318_n 3.39184e-19 $X=1.975 $Y=2.13 $X2=0 $Y2=0
cc_269 N_D_c_263_n N_A_202_463#_c_318_n 0.00116834f $X=1.6 $Y=1.99 $X2=0 $Y2=0
cc_270 N_D_c_262_n N_A_202_463#_c_319_n 0.016825f $X=1.925 $Y=1.2 $X2=0 $Y2=0
cc_271 N_D_c_263_n N_A_202_463#_c_319_n 0.00462151f $X=1.6 $Y=1.99 $X2=0 $Y2=0
cc_272 N_D_c_261_n N_A_202_463#_c_322_n 0.00298049f $X=1.925 $Y=1.125 $X2=0
+ $Y2=0
cc_273 N_D_c_262_n N_A_202_463#_c_322_n 0.00789225f $X=1.925 $Y=1.2 $X2=0 $Y2=0
cc_274 N_D_c_265_n N_A_33_463#_M1024_g 0.00633326f $X=1.975 $Y=2.13 $X2=0 $Y2=0
cc_275 N_D_c_262_n N_A_33_463#_M1018_g 0.0074267f $X=1.925 $Y=1.2 $X2=0 $Y2=0
cc_276 N_D_c_264_n N_A_33_463#_c_854_n 0.0104164f $X=1.975 $Y=2.205 $X2=0 $Y2=0
cc_277 N_D_c_261_n N_A_33_463#_c_844_n 0.0104164f $X=1.925 $Y=1.125 $X2=0 $Y2=0
cc_278 N_D_c_261_n N_A_33_463#_M1028_g 0.0117695f $X=1.925 $Y=1.125 $X2=0 $Y2=0
cc_279 N_D_c_263_n N_A_33_463#_c_852_n 0.01376f $X=1.6 $Y=1.99 $X2=0 $Y2=0
cc_280 N_D_c_264_n N_VPWR_c_1230_n 0.00598921f $X=1.975 $Y=2.205 $X2=0 $Y2=0
cc_281 N_D_c_265_n N_VPWR_c_1230_n 0.00720581f $X=1.975 $Y=2.13 $X2=0 $Y2=0
cc_282 D N_VPWR_c_1230_n 0.0198258f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_283 N_D_c_264_n N_VPWR_c_1228_n 9.39239e-19 $X=1.975 $Y=2.205 $X2=0 $Y2=0
cc_284 N_D_c_261_n N_A_400_119#_c_1363_n 0.00267292f $X=1.925 $Y=1.125 $X2=0
+ $Y2=0
cc_285 N_D_c_265_n N_A_400_119#_c_1366_n 0.00350618f $X=1.975 $Y=2.13 $X2=0
+ $Y2=0
cc_286 D N_A_400_119#_c_1364_n 0.00493741f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_287 N_D_c_263_n N_A_400_119#_c_1364_n 0.00365197f $X=1.6 $Y=1.99 $X2=0 $Y2=0
cc_288 N_D_c_262_n N_A_400_119#_c_1365_n 0.00222981f $X=1.925 $Y=1.2 $X2=0 $Y2=0
cc_289 N_D_c_265_n N_A_400_119#_c_1368_n 0.0014731f $X=1.975 $Y=2.13 $X2=0 $Y2=0
cc_290 D N_A_400_119#_c_1368_n 0.0113899f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_291 N_D_c_261_n N_VGND_c_1484_n 0.00598921f $X=1.925 $Y=1.125 $X2=0 $Y2=0
cc_292 N_D_c_262_n N_VGND_c_1484_n 0.00889024f $X=1.925 $Y=1.2 $X2=0 $Y2=0
cc_293 N_D_c_261_n N_VGND_c_1494_n 9.39239e-19 $X=1.925 $Y=1.125 $X2=0 $Y2=0
cc_294 N_A_202_463#_c_319_n N_A_614_93#_c_486_n 9.75623e-19 $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_295 N_A_202_463#_M1001_g N_A_614_93#_c_487_n 0.00301598f $X=2.405 $Y=2.525
+ $X2=0 $Y2=0
cc_296 N_A_202_463#_c_319_n N_A_614_93#_c_479_n 0.0229961f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_297 N_A_202_463#_M1030_g N_A_614_93#_c_481_n 5.5359e-19 $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_298 N_A_202_463#_c_319_n N_A_614_93#_c_481_n 0.0236301f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_299 N_A_202_463#_c_319_n N_A_614_93#_c_482_n 0.00358296f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_300 N_A_202_463#_M1030_g N_A_614_93#_c_483_n 0.0606885f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_301 N_A_202_463#_M1030_g N_A_614_93#_c_484_n 0.00995233f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_302 N_A_202_463#_c_313_n N_A_614_93#_c_484_n 0.00301598f $X=2.405 $Y=1.68
+ $X2=0 $Y2=0
cc_303 N_A_202_463#_c_319_n N_SET_B_c_566_n 0.0256069f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_304 N_A_202_463#_c_319_n N_SET_B_c_568_n 0.0119359f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_305 N_A_202_463#_c_319_n N_SET_B_c_569_n 0.00446679f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_306 N_A_202_463#_c_319_n N_SET_B_c_577_n 0.00649093f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_307 N_A_202_463#_c_319_n N_SET_B_c_578_n 3.45956e-19 $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_308 N_A_202_463#_M1013_g N_SET_B_c_581_n 0.019011f $X=5.8 $Y=2.295 $X2=0
+ $Y2=0
cc_309 N_A_202_463#_c_314_n N_SET_B_c_581_n 0.00892654f $X=5.725 $Y=1.51 $X2=0
+ $Y2=0
cc_310 N_A_202_463#_c_315_n N_SET_B_c_581_n 3.57318e-19 $X=5.725 $Y=1.345 $X2=0
+ $Y2=0
cc_311 N_A_202_463#_c_319_n N_SET_B_c_581_n 0.026533f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_312 N_A_202_463#_c_320_n N_SET_B_c_581_n 0.00142993f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_313 N_A_202_463#_c_321_n N_SET_B_c_581_n 0.0237638f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_314 N_A_202_463#_M1031_g N_SET_B_c_573_n 0.00284962f $X=5.835 $Y=0.555 $X2=0
+ $Y2=0
cc_315 N_A_202_463#_c_315_n N_SET_B_c_573_n 0.0127778f $X=5.725 $Y=1.345 $X2=0
+ $Y2=0
cc_316 N_A_202_463#_c_320_n N_SET_B_c_573_n 0.00113103f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_317 N_A_202_463#_c_321_n N_SET_B_c_573_n 0.026186f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_318 N_A_202_463#_c_319_n N_A_486_119#_M1027_g 0.00794791f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_319 N_A_202_463#_c_319_n N_A_486_119#_c_696_n 0.00433769f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_320 N_A_202_463#_c_319_n N_A_486_119#_c_697_n 0.0125111f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_321 N_A_202_463#_c_314_n N_A_486_119#_M1007_g 0.00534963f $X=5.725 $Y=1.51
+ $X2=0 $Y2=0
cc_322 N_A_202_463#_c_321_n N_A_486_119#_M1007_g 6.0798e-19 $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_323 N_A_202_463#_M1031_g N_A_486_119#_c_699_n 0.0036183f $X=5.835 $Y=0.555
+ $X2=0 $Y2=0
cc_324 N_A_202_463#_c_319_n N_A_486_119#_c_699_n 0.00502906f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_325 N_A_202_463#_c_320_n N_A_486_119#_c_699_n 7.47463e-19 $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_326 N_A_202_463#_c_321_n N_A_486_119#_c_699_n 0.00219474f $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_327 N_A_202_463#_c_314_n N_A_486_119#_c_700_n 0.0115306f $X=5.725 $Y=1.51
+ $X2=0 $Y2=0
cc_328 N_A_202_463#_c_319_n N_A_486_119#_c_700_n 0.00464229f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_329 N_A_202_463#_c_320_n N_A_486_119#_c_700_n 0.00283145f $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_330 N_A_202_463#_c_321_n N_A_486_119#_c_700_n 0.00294218f $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_331 N_A_202_463#_M1031_g N_A_486_119#_c_702_n 0.0626345f $X=5.835 $Y=0.555
+ $X2=0 $Y2=0
cc_332 N_A_202_463#_c_314_n N_A_486_119#_c_703_n 0.00953349f $X=5.725 $Y=1.51
+ $X2=0 $Y2=0
cc_333 N_A_202_463#_c_319_n N_A_486_119#_c_703_n 0.0061641f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_334 N_A_202_463#_c_321_n N_A_486_119#_c_703_n 0.00131332f $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_335 N_A_202_463#_c_309_n N_A_486_119#_c_730_n 0.00262201f $X=2.71 $Y=1.59
+ $X2=0 $Y2=0
cc_336 N_A_202_463#_M1030_g N_A_486_119#_c_730_n 0.00917911f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_337 N_A_202_463#_c_319_n N_A_486_119#_c_730_n 0.0088717f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_338 N_A_202_463#_c_309_n N_A_486_119#_c_704_n 0.00110908f $X=2.71 $Y=1.59
+ $X2=0 $Y2=0
cc_339 N_A_202_463#_M1030_g N_A_486_119#_c_704_n 0.011312f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_340 N_A_202_463#_c_319_n N_A_486_119#_c_704_n 0.0234185f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_341 N_A_202_463#_M1001_g N_A_486_119#_c_709_n 0.00151667f $X=2.405 $Y=2.525
+ $X2=0 $Y2=0
cc_342 N_A_202_463#_c_313_n N_A_486_119#_c_709_n 9.29497e-19 $X=2.405 $Y=1.68
+ $X2=0 $Y2=0
cc_343 N_A_202_463#_c_319_n N_A_486_119#_c_705_n 0.0166916f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_344 N_A_202_463#_M1001_g N_A_486_119#_c_739_n 0.00402094f $X=2.405 $Y=2.525
+ $X2=0 $Y2=0
cc_345 N_A_202_463#_c_309_n N_A_486_119#_c_739_n 0.00352831f $X=2.71 $Y=1.59
+ $X2=0 $Y2=0
cc_346 N_A_202_463#_c_309_n N_A_486_119#_c_711_n 0.00593159f $X=2.71 $Y=1.59
+ $X2=0 $Y2=0
cc_347 N_A_202_463#_c_313_n N_A_486_119#_c_711_n 2.3586e-19 $X=2.405 $Y=1.68
+ $X2=0 $Y2=0
cc_348 N_A_202_463#_c_319_n N_A_486_119#_c_706_n 0.0102366f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_349 N_A_202_463#_c_322_n N_A_33_463#_M1018_g 0.0253985f $X=1.19 $Y=0.575
+ $X2=0 $Y2=0
cc_350 N_A_202_463#_M1001_g N_A_33_463#_c_854_n 0.0103135f $X=2.405 $Y=2.525
+ $X2=0 $Y2=0
cc_351 N_A_202_463#_c_330_n N_A_33_463#_c_854_n 0.00361319f $X=1.15 $Y=2.46
+ $X2=0 $Y2=0
cc_352 N_A_202_463#_c_322_n N_A_33_463#_c_844_n 0.00488572f $X=1.19 $Y=0.575
+ $X2=0 $Y2=0
cc_353 N_A_202_463#_M1030_g N_A_33_463#_M1028_g 0.0132634f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_354 N_A_202_463#_c_312_n N_A_33_463#_M1028_g 0.00439319f $X=2.33 $Y=1.68
+ $X2=0 $Y2=0
cc_355 N_A_202_463#_M1001_g N_A_33_463#_M1020_g 0.0134264f $X=2.405 $Y=2.525
+ $X2=0 $Y2=0
cc_356 N_A_202_463#_c_309_n N_A_33_463#_M1020_g 0.00181966f $X=2.71 $Y=1.59
+ $X2=0 $Y2=0
cc_357 N_A_202_463#_M1013_g N_A_33_463#_c_857_n 0.00313337f $X=5.8 $Y=2.295
+ $X2=0 $Y2=0
cc_358 N_A_202_463#_M1031_g N_A_33_463#_M1014_g 0.0233111f $X=5.835 $Y=0.555
+ $X2=0 $Y2=0
cc_359 N_A_202_463#_c_315_n N_A_33_463#_M1014_g 0.00817844f $X=5.725 $Y=1.345
+ $X2=0 $Y2=0
cc_360 N_A_202_463#_M1013_g N_A_33_463#_c_861_n 0.0205863f $X=5.8 $Y=2.295 $X2=0
+ $Y2=0
cc_361 N_A_202_463#_c_330_n N_A_33_463#_c_862_n 0.0147212f $X=1.15 $Y=2.46 $X2=0
+ $Y2=0
cc_362 N_A_202_463#_c_330_n N_A_33_463#_c_849_n 0.0095956f $X=1.15 $Y=2.46 $X2=0
+ $Y2=0
cc_363 N_A_202_463#_c_317_n N_A_33_463#_c_849_n 0.0102702f $X=1.2 $Y=1.6 $X2=0
+ $Y2=0
cc_364 N_A_202_463#_c_330_n N_A_33_463#_c_852_n 0.01096f $X=1.15 $Y=2.46 $X2=0
+ $Y2=0
cc_365 N_A_202_463#_c_317_n N_A_33_463#_c_852_n 0.00588528f $X=1.2 $Y=1.6 $X2=0
+ $Y2=0
cc_366 N_A_202_463#_c_322_n N_A_33_463#_c_852_n 0.00195277f $X=1.19 $Y=0.575
+ $X2=0 $Y2=0
cc_367 N_A_202_463#_M1031_g N_A_1175_417#_c_1078_n 0.0105184f $X=5.835 $Y=0.555
+ $X2=0 $Y2=0
cc_368 N_A_202_463#_M1031_g N_A_1175_417#_c_1080_n 0.00604642f $X=5.835 $Y=0.555
+ $X2=0 $Y2=0
cc_369 N_A_202_463#_c_330_n N_VPWR_c_1229_n 0.0252281f $X=1.15 $Y=2.46 $X2=0
+ $Y2=0
cc_370 N_A_202_463#_c_330_n N_VPWR_c_1230_n 0.0290117f $X=1.15 $Y=2.46 $X2=0
+ $Y2=0
cc_371 N_A_202_463#_c_316_n N_VPWR_c_1230_n 9.68106e-19 $X=2.005 $Y=1.6 $X2=0
+ $Y2=0
cc_372 N_A_202_463#_c_330_n N_VPWR_c_1243_n 0.00874746f $X=1.15 $Y=2.46 $X2=0
+ $Y2=0
cc_373 N_A_202_463#_M1001_g N_VPWR_c_1228_n 9.39239e-19 $X=2.405 $Y=2.525 $X2=0
+ $Y2=0
cc_374 N_A_202_463#_c_330_n N_VPWR_c_1228_n 0.00677813f $X=1.15 $Y=2.46 $X2=0
+ $Y2=0
cc_375 N_A_202_463#_M1030_g N_A_400_119#_c_1363_n 5.0512e-19 $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_376 N_A_202_463#_c_319_n N_A_400_119#_c_1363_n 0.00232109f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_377 N_A_202_463#_c_322_n N_A_400_119#_c_1363_n 0.00562089f $X=1.19 $Y=0.575
+ $X2=0 $Y2=0
cc_378 N_A_202_463#_M1001_g N_A_400_119#_c_1366_n 0.00156129f $X=2.405 $Y=2.525
+ $X2=0 $Y2=0
cc_379 N_A_202_463#_M1001_g N_A_400_119#_c_1364_n 0.0061702f $X=2.405 $Y=2.525
+ $X2=0 $Y2=0
cc_380 N_A_202_463#_c_309_n N_A_400_119#_c_1364_n 0.00691721f $X=2.71 $Y=1.59
+ $X2=0 $Y2=0
cc_381 N_A_202_463#_M1030_g N_A_400_119#_c_1364_n 0.00331333f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_382 N_A_202_463#_c_313_n N_A_400_119#_c_1364_n 0.00995053f $X=2.405 $Y=1.68
+ $X2=0 $Y2=0
cc_383 N_A_202_463#_c_318_n N_A_400_119#_c_1364_n 0.0228995f $X=2.12 $Y=1.6
+ $X2=0 $Y2=0
cc_384 N_A_202_463#_c_319_n N_A_400_119#_c_1364_n 0.00564604f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_385 N_A_202_463#_M1030_g N_A_400_119#_c_1365_n 0.00211719f $X=2.785 $Y=0.805
+ $X2=0 $Y2=0
cc_386 N_A_202_463#_c_312_n N_A_400_119#_c_1365_n 0.00404983f $X=2.33 $Y=1.68
+ $X2=0 $Y2=0
cc_387 N_A_202_463#_c_313_n N_A_400_119#_c_1365_n 7.311e-19 $X=2.405 $Y=1.68
+ $X2=0 $Y2=0
cc_388 N_A_202_463#_c_318_n N_A_400_119#_c_1365_n 0.0144231f $X=2.12 $Y=1.6
+ $X2=0 $Y2=0
cc_389 N_A_202_463#_c_319_n N_A_400_119#_c_1365_n 0.0230827f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_390 N_A_202_463#_c_322_n N_A_400_119#_c_1365_n 0.00341899f $X=1.19 $Y=0.575
+ $X2=0 $Y2=0
cc_391 N_A_202_463#_M1001_g N_A_400_119#_c_1368_n 0.0144857f $X=2.405 $Y=2.525
+ $X2=0 $Y2=0
cc_392 N_A_202_463#_c_309_n N_A_400_119#_c_1368_n 2.88929e-19 $X=2.71 $Y=1.59
+ $X2=0 $Y2=0
cc_393 N_A_202_463#_c_312_n N_A_400_119#_c_1368_n 0.00379625f $X=2.33 $Y=1.68
+ $X2=0 $Y2=0
cc_394 N_A_202_463#_c_318_n N_A_400_119#_c_1368_n 0.0127641f $X=2.12 $Y=1.6
+ $X2=0 $Y2=0
cc_395 N_A_202_463#_M1013_g N_A_985_379#_c_1414_n 0.00115351f $X=5.8 $Y=2.295
+ $X2=0 $Y2=0
cc_396 N_A_202_463#_M1013_g N_A_985_379#_c_1416_n 5.2646e-19 $X=5.8 $Y=2.295
+ $X2=0 $Y2=0
cc_397 N_A_202_463#_M1013_g N_A_1092_417#_c_1440_n 0.00591332f $X=5.8 $Y=2.295
+ $X2=0 $Y2=0
cc_398 N_A_202_463#_M1013_g N_A_1092_417#_c_1441_n 0.00333555f $X=5.8 $Y=2.295
+ $X2=0 $Y2=0
cc_399 N_A_202_463#_M1013_g N_A_1092_417#_c_1443_n 0.007797f $X=5.8 $Y=2.295
+ $X2=0 $Y2=0
cc_400 N_A_202_463#_c_316_n N_VGND_c_1484_n 0.00375685f $X=2.005 $Y=1.6 $X2=0
+ $Y2=0
cc_401 N_A_202_463#_c_319_n N_VGND_c_1484_n 0.00775753f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_402 N_A_202_463#_c_322_n N_VGND_c_1484_n 0.0426097f $X=1.19 $Y=0.575 $X2=0
+ $Y2=0
cc_403 N_A_202_463#_c_319_n N_VGND_c_1485_n 6.72865e-19 $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_404 N_A_202_463#_c_322_n N_VGND_c_1488_n 0.0098177f $X=1.19 $Y=0.575 $X2=0
+ $Y2=0
cc_405 N_A_202_463#_M1030_g N_VGND_c_1489_n 0.00333474f $X=2.785 $Y=0.805 $X2=0
+ $Y2=0
cc_406 N_A_202_463#_M1031_g N_VGND_c_1491_n 0.00549943f $X=5.835 $Y=0.555 $X2=0
+ $Y2=0
cc_407 N_A_202_463#_M1030_g N_VGND_c_1494_n 0.00477801f $X=2.785 $Y=0.805 $X2=0
+ $Y2=0
cc_408 N_A_202_463#_M1031_g N_VGND_c_1494_n 0.0111536f $X=5.835 $Y=0.555 $X2=0
+ $Y2=0
cc_409 N_A_202_463#_c_322_n N_VGND_c_1494_n 0.00967822f $X=1.19 $Y=0.575 $X2=0
+ $Y2=0
cc_410 N_A_202_463#_M1031_g N_VGND_c_1498_n 0.00308692f $X=5.835 $Y=0.555 $X2=0
+ $Y2=0
cc_411 N_A_202_463#_c_319_n N_VGND_c_1498_n 0.0228091f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_412 N_A_202_463#_c_320_n N_VGND_c_1498_n 0.00145022f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_413 N_A_202_463#_c_321_n N_VGND_c_1498_n 8.88587e-19 $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_414 N_A_614_93#_c_488_n N_SET_B_M1025_g 0.00181625f $X=3.835 $Y=2.36 $X2=0
+ $Y2=0
cc_415 N_A_614_93#_c_500_p N_SET_B_M1025_g 0.00418347f $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_416 N_A_614_93#_c_479_n N_SET_B_c_566_n 7.41974e-19 $X=3.81 $Y=1.02 $X2=0
+ $Y2=0
cc_417 N_A_614_93#_c_479_n N_SET_B_c_567_n 0.0135397f $X=3.81 $Y=1.02 $X2=0
+ $Y2=0
cc_418 N_A_614_93#_c_480_n N_SET_B_c_567_n 0.00707492f $X=3.975 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_614_93#_c_486_n N_SET_B_c_577_n 0.0216534f $X=3.75 $Y=2.025 $X2=0
+ $Y2=0
cc_420 N_A_614_93#_c_500_p N_SET_B_c_577_n 0.00161064f $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_421 N_A_614_93#_c_486_n N_SET_B_c_578_n 0.00183212f $X=3.75 $Y=2.025 $X2=0
+ $Y2=0
cc_422 N_A_614_93#_c_500_p N_SET_B_c_578_n 0.00161634f $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_423 N_A_614_93#_M1023_g N_A_486_119#_M1003_g 0.0131453f $X=3.195 $Y=2.525
+ $X2=0 $Y2=0
cc_424 N_A_614_93#_c_486_n N_A_486_119#_M1003_g 0.0132855f $X=3.75 $Y=2.025
+ $X2=0 $Y2=0
cc_425 N_A_614_93#_c_487_n N_A_486_119#_M1003_g 0.0215558f $X=3.285 $Y=1.99
+ $X2=0 $Y2=0
cc_426 N_A_614_93#_c_488_n N_A_486_119#_M1003_g 0.00579968f $X=3.835 $Y=2.36
+ $X2=0 $Y2=0
cc_427 N_A_614_93#_c_500_p N_A_486_119#_M1003_g 0.00527628f $X=3.95 $Y=2.525
+ $X2=0 $Y2=0
cc_428 N_A_614_93#_c_479_n N_A_486_119#_M1027_g 0.00406888f $X=3.81 $Y=1.02
+ $X2=0 $Y2=0
cc_429 N_A_614_93#_c_480_n N_A_486_119#_M1027_g 0.0103177f $X=3.975 $Y=0.445
+ $X2=0 $Y2=0
cc_430 N_A_614_93#_c_481_n N_A_486_119#_M1027_g 0.00126311f $X=3.27 $Y=1.02
+ $X2=0 $Y2=0
cc_431 N_A_614_93#_c_482_n N_A_486_119#_M1027_g 0.00288132f $X=3.27 $Y=1.29
+ $X2=0 $Y2=0
cc_432 N_A_614_93#_c_486_n N_A_486_119#_c_697_n 6.3026e-19 $X=3.75 $Y=2.025
+ $X2=0 $Y2=0
cc_433 N_A_614_93#_c_479_n N_A_486_119#_c_697_n 0.00800195f $X=3.81 $Y=1.02
+ $X2=0 $Y2=0
cc_434 N_A_614_93#_c_481_n N_A_486_119#_c_697_n 3.7339e-19 $X=3.27 $Y=1.02 $X2=0
+ $Y2=0
cc_435 N_A_614_93#_c_482_n N_A_486_119#_c_697_n 0.0112512f $X=3.27 $Y=1.29 $X2=0
+ $Y2=0
cc_436 N_A_614_93#_c_484_n N_A_486_119#_c_697_n 0.0120902f $X=3.285 $Y=1.825
+ $X2=0 $Y2=0
cc_437 N_A_614_93#_c_481_n N_A_486_119#_c_730_n 0.00309468f $X=3.27 $Y=1.02
+ $X2=0 $Y2=0
cc_438 N_A_614_93#_c_483_n N_A_486_119#_c_730_n 0.00565171f $X=3.252 $Y=1.125
+ $X2=0 $Y2=0
cc_439 N_A_614_93#_c_481_n N_A_486_119#_c_704_n 0.0282623f $X=3.27 $Y=1.02 $X2=0
+ $Y2=0
cc_440 N_A_614_93#_c_483_n N_A_486_119#_c_704_n 0.00354763f $X=3.252 $Y=1.125
+ $X2=0 $Y2=0
cc_441 N_A_614_93#_c_484_n N_A_486_119#_c_704_n 0.00196561f $X=3.285 $Y=1.825
+ $X2=0 $Y2=0
cc_442 N_A_614_93#_c_486_n N_A_486_119#_c_709_n 0.0185796f $X=3.75 $Y=2.025
+ $X2=0 $Y2=0
cc_443 N_A_614_93#_c_487_n N_A_486_119#_c_709_n 0.00436738f $X=3.285 $Y=1.99
+ $X2=0 $Y2=0
cc_444 N_A_614_93#_c_484_n N_A_486_119#_c_709_n 0.0040441f $X=3.285 $Y=1.825
+ $X2=0 $Y2=0
cc_445 N_A_614_93#_c_486_n N_A_486_119#_c_705_n 0.0388424f $X=3.75 $Y=2.025
+ $X2=0 $Y2=0
cc_446 N_A_614_93#_c_487_n N_A_486_119#_c_705_n 0.00174871f $X=3.285 $Y=1.99
+ $X2=0 $Y2=0
cc_447 N_A_614_93#_c_479_n N_A_486_119#_c_705_n 0.00401656f $X=3.81 $Y=1.02
+ $X2=0 $Y2=0
cc_448 N_A_614_93#_c_481_n N_A_486_119#_c_705_n 0.0226805f $X=3.27 $Y=1.02 $X2=0
+ $Y2=0
cc_449 N_A_614_93#_c_482_n N_A_486_119#_c_705_n 0.00340995f $X=3.27 $Y=1.29
+ $X2=0 $Y2=0
cc_450 N_A_614_93#_c_484_n N_A_486_119#_c_705_n 0.0111361f $X=3.285 $Y=1.825
+ $X2=0 $Y2=0
cc_451 N_A_614_93#_c_486_n N_A_486_119#_c_706_n 0.0204436f $X=3.75 $Y=2.025
+ $X2=0 $Y2=0
cc_452 N_A_614_93#_c_479_n N_A_486_119#_c_706_n 0.0159748f $X=3.81 $Y=1.02 $X2=0
+ $Y2=0
cc_453 N_A_614_93#_c_481_n N_A_486_119#_c_706_n 0.00499564f $X=3.27 $Y=1.02
+ $X2=0 $Y2=0
cc_454 N_A_614_93#_c_482_n N_A_486_119#_c_706_n 8.49171e-19 $X=3.27 $Y=1.29
+ $X2=0 $Y2=0
cc_455 N_A_614_93#_c_484_n N_A_486_119#_c_706_n 6.90045e-19 $X=3.285 $Y=1.825
+ $X2=0 $Y2=0
cc_456 N_A_614_93#_M1023_g N_A_33_463#_M1020_g 0.0406737f $X=3.195 $Y=2.525
+ $X2=0 $Y2=0
cc_457 N_A_614_93#_M1023_g N_A_33_463#_c_857_n 0.0104164f $X=3.195 $Y=2.525
+ $X2=0 $Y2=0
cc_458 N_A_614_93#_c_500_p N_A_33_463#_c_857_n 0.00479477f $X=3.95 $Y=2.525
+ $X2=0 $Y2=0
cc_459 N_A_614_93#_M1023_g N_VPWR_c_1231_n 0.00381479f $X=3.195 $Y=2.525 $X2=0
+ $Y2=0
cc_460 N_A_614_93#_c_486_n N_VPWR_c_1231_n 0.0192115f $X=3.75 $Y=2.025 $X2=0
+ $Y2=0
cc_461 N_A_614_93#_c_487_n N_VPWR_c_1231_n 0.00341875f $X=3.285 $Y=1.99 $X2=0
+ $Y2=0
cc_462 N_A_614_93#_c_500_p N_VPWR_c_1231_n 0.0254941f $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_463 N_A_614_93#_c_488_n N_VPWR_c_1232_n 0.00671235f $X=3.835 $Y=2.36 $X2=0
+ $Y2=0
cc_464 N_A_614_93#_c_500_p N_VPWR_c_1244_n 0.00551488f $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_465 N_A_614_93#_M1023_g N_VPWR_c_1228_n 9.39239e-19 $X=3.195 $Y=2.525 $X2=0
+ $Y2=0
cc_466 N_A_614_93#_c_500_p N_VPWR_c_1228_n 0.009118f $X=3.95 $Y=2.525 $X2=0
+ $Y2=0
cc_467 N_A_614_93#_c_484_n N_A_400_119#_c_1364_n 3.77668e-19 $X=3.285 $Y=1.825
+ $X2=0 $Y2=0
cc_468 N_A_614_93#_c_479_n N_VGND_M1022_d 0.0018073f $X=3.81 $Y=1.02 $X2=0 $Y2=0
cc_469 N_A_614_93#_c_481_n N_VGND_M1022_d 0.00240407f $X=3.27 $Y=1.02 $X2=0
+ $Y2=0
cc_470 N_A_614_93#_c_479_n N_VGND_c_1485_n 0.0144186f $X=3.81 $Y=1.02 $X2=0
+ $Y2=0
cc_471 N_A_614_93#_c_480_n N_VGND_c_1485_n 0.0367878f $X=3.975 $Y=0.445 $X2=0
+ $Y2=0
cc_472 N_A_614_93#_c_481_n N_VGND_c_1485_n 0.0119973f $X=3.27 $Y=1.02 $X2=0
+ $Y2=0
cc_473 N_A_614_93#_c_482_n N_VGND_c_1485_n 7.27774e-19 $X=3.27 $Y=1.29 $X2=0
+ $Y2=0
cc_474 N_A_614_93#_c_483_n N_VGND_c_1485_n 0.010445f $X=3.252 $Y=1.125 $X2=0
+ $Y2=0
cc_475 N_A_614_93#_c_483_n N_VGND_c_1489_n 0.00431487f $X=3.252 $Y=1.125 $X2=0
+ $Y2=0
cc_476 N_A_614_93#_c_480_n N_VGND_c_1490_n 0.0156583f $X=3.975 $Y=0.445 $X2=0
+ $Y2=0
cc_477 N_A_614_93#_M1027_s N_VGND_c_1494_n 0.00342001f $X=3.85 $Y=0.235 $X2=0
+ $Y2=0
cc_478 N_A_614_93#_c_480_n N_VGND_c_1494_n 0.0102927f $X=3.975 $Y=0.445 $X2=0
+ $Y2=0
cc_479 N_A_614_93#_c_483_n N_VGND_c_1494_n 0.00477801f $X=3.252 $Y=1.125 $X2=0
+ $Y2=0
cc_480 N_SET_B_M1025_g N_A_486_119#_M1003_g 0.0131801f $X=4.165 $Y=2.525 $X2=0
+ $Y2=0
cc_481 N_SET_B_c_566_n N_A_486_119#_M1003_g 0.00154126f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_482 N_SET_B_c_577_n N_A_486_119#_M1003_g 0.00282069f $X=4.44 $Y=1.85 $X2=0
+ $Y2=0
cc_483 N_SET_B_c_578_n N_A_486_119#_M1003_g 0.0205812f $X=4.185 $Y=1.99 $X2=0
+ $Y2=0
cc_484 N_SET_B_c_566_n N_A_486_119#_M1027_g 0.00863616f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_485 N_SET_B_c_567_n N_A_486_119#_M1027_g 0.00201521f $X=4.44 $Y=0.97 $X2=0
+ $Y2=0
cc_486 N_SET_B_c_571_n N_A_486_119#_M1027_g 0.0601159f $X=4.64 $Y=0.765 $X2=0
+ $Y2=0
cc_487 N_SET_B_c_566_n N_A_486_119#_c_696_n 0.0162146f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_488 N_SET_B_c_568_n N_A_486_119#_c_696_n 0.00180668f $X=4.64 $Y=0.93 $X2=0
+ $Y2=0
cc_489 N_SET_B_c_569_n N_A_486_119#_c_696_n 0.0203848f $X=4.64 $Y=0.93 $X2=0
+ $Y2=0
cc_490 N_SET_B_c_581_n N_A_486_119#_c_696_n 0.00697048f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_491 N_SET_B_c_566_n N_A_486_119#_c_697_n 0.0027806f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_492 N_SET_B_c_577_n N_A_486_119#_c_697_n 0.00416284f $X=4.44 $Y=1.85 $X2=0
+ $Y2=0
cc_493 N_SET_B_c_578_n N_A_486_119#_c_697_n 0.0122738f $X=4.185 $Y=1.99 $X2=0
+ $Y2=0
cc_494 N_SET_B_M1025_g N_A_486_119#_M1007_g 0.00503758f $X=4.165 $Y=2.525 $X2=0
+ $Y2=0
cc_495 N_SET_B_c_566_n N_A_486_119#_M1007_g 0.00801263f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_496 N_SET_B_c_577_n N_A_486_119#_M1007_g 8.1252e-19 $X=4.44 $Y=1.85 $X2=0
+ $Y2=0
cc_497 N_SET_B_c_578_n N_A_486_119#_M1007_g 0.00830787f $X=4.185 $Y=1.99 $X2=0
+ $Y2=0
cc_498 N_SET_B_c_581_n N_A_486_119#_M1007_g 0.0183571f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_499 N_SET_B_c_581_n N_A_486_119#_c_700_n 0.00445615f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_500 N_SET_B_c_566_n N_A_486_119#_c_701_n 0.00450057f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_501 N_SET_B_c_568_n N_A_486_119#_c_701_n 8.1028e-19 $X=4.64 $Y=0.93 $X2=0
+ $Y2=0
cc_502 N_SET_B_c_569_n N_A_486_119#_c_701_n 0.0071852f $X=4.64 $Y=0.93 $X2=0
+ $Y2=0
cc_503 N_SET_B_c_568_n N_A_486_119#_c_702_n 5.11372e-19 $X=4.64 $Y=0.93 $X2=0
+ $Y2=0
cc_504 N_SET_B_c_569_n N_A_486_119#_c_702_n 0.00234103f $X=4.64 $Y=0.93 $X2=0
+ $Y2=0
cc_505 N_SET_B_c_581_n N_A_486_119#_c_703_n 0.00859788f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_506 N_SET_B_c_566_n N_A_486_119#_c_706_n 0.017879f $X=4.355 $Y=1.765 $X2=0
+ $Y2=0
cc_507 N_SET_B_M1025_g N_A_33_463#_c_857_n 0.0103123f $X=4.165 $Y=2.525 $X2=0
+ $Y2=0
cc_508 SET_B N_A_33_463#_M1014_g 0.0239759f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_509 SET_B N_A_33_463#_c_861_n 0.00695453f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_510 N_SET_B_c_573_n N_A_33_463#_c_861_n 5.29598e-19 $X=6.055 $Y=1.59 $X2=0
+ $Y2=0
cc_511 N_SET_B_M1008_g N_A_1329_65#_M1015_g 0.0682058f $X=7.08 $Y=0.665 $X2=0
+ $Y2=0
cc_512 SET_B N_A_1329_65#_M1015_g 0.0256264f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_513 N_SET_B_c_572_n N_A_1329_65#_M1015_g 0.00965721f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_514 N_SET_B_M1021_g N_A_1329_65#_M1002_g 0.0145372f $X=7.83 $Y=2.525 $X2=0
+ $Y2=0
cc_515 N_SET_B_c_572_n N_A_1329_65#_M1002_g 0.00718355f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_516 N_SET_B_M1021_g N_A_1329_65#_c_989_n 0.0103162f $X=7.83 $Y=2.525 $X2=0
+ $Y2=0
cc_517 SET_B N_A_1329_65#_c_990_n 0.0110687f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_518 N_SET_B_c_572_n N_A_1329_65#_c_990_n 0.00241035f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_519 N_SET_B_M1021_g N_A_1329_65#_c_993_n 0.00310094f $X=7.83 $Y=2.525 $X2=0
+ $Y2=0
cc_520 N_SET_B_c_572_n N_A_1329_65#_c_983_n 4.72116e-19 $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_521 N_SET_B_c_572_n N_A_1175_417#_c_1069_n 0.00836355f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_522 N_SET_B_M1008_g N_A_1175_417#_c_1071_n 0.0154854f $X=7.08 $Y=0.665 $X2=0
+ $Y2=0
cc_523 N_SET_B_c_572_n N_A_1175_417#_M1010_g 0.00969809f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_524 N_SET_B_c_572_n N_A_1175_417#_c_1076_n 0.00499022f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_525 N_SET_B_M1008_g N_A_1175_417#_c_1079_n 0.014662f $X=7.08 $Y=0.665 $X2=0
+ $Y2=0
cc_526 SET_B N_A_1175_417#_c_1079_n 0.103542f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_527 N_SET_B_c_572_n N_A_1175_417#_c_1079_n 0.0148871f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_528 N_SET_B_c_573_n N_A_1175_417#_c_1080_n 0.0386748f $X=6.055 $Y=1.59 $X2=0
+ $Y2=0
cc_529 N_SET_B_M1021_g N_A_1175_417#_c_1086_n 0.00501345f $X=7.83 $Y=2.525 $X2=0
+ $Y2=0
cc_530 N_SET_B_c_572_n N_A_1175_417#_c_1086_n 0.0117511f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_531 N_SET_B_M1021_g N_A_1175_417#_c_1081_n 0.0112855f $X=7.83 $Y=2.525 $X2=0
+ $Y2=0
cc_532 SET_B N_A_1175_417#_c_1081_n 0.0455806f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_533 N_SET_B_c_572_n N_A_1175_417#_c_1081_n 0.0222612f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_534 N_SET_B_M1021_g N_A_1175_417#_c_1088_n 0.00722671f $X=7.83 $Y=2.525 $X2=0
+ $Y2=0
cc_535 SET_B N_A_1175_417#_c_1106_n 0.0124662f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_536 N_SET_B_c_573_n N_A_1175_417#_c_1106_n 0.0109259f $X=6.055 $Y=1.59 $X2=0
+ $Y2=0
cc_537 SET_B N_A_1175_417#_c_1108_n 0.102648f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_538 N_SET_B_M1008_g N_A_1175_417#_c_1082_n 0.00435706f $X=7.08 $Y=0.665 $X2=0
+ $Y2=0
cc_539 SET_B N_A_1175_417#_c_1082_n 0.00755058f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_540 N_SET_B_c_572_n N_A_1175_417#_c_1082_n 0.00602152f $X=7.44 $Y=1.41 $X2=0
+ $Y2=0
cc_541 N_SET_B_M1021_g N_A_1175_417#_c_1089_n 0.0101885f $X=7.83 $Y=2.525 $X2=0
+ $Y2=0
cc_542 N_SET_B_c_581_n N_VPWR_M1025_d 0.00235139f $X=5.885 $Y=1.59 $X2=0 $Y2=0
cc_543 N_SET_B_M1025_g N_VPWR_c_1232_n 0.00224459f $X=4.165 $Y=2.525 $X2=0 $Y2=0
cc_544 N_SET_B_c_577_n N_VPWR_c_1232_n 0.0109302f $X=4.44 $Y=1.85 $X2=0 $Y2=0
cc_545 N_SET_B_c_578_n N_VPWR_c_1232_n 0.00182828f $X=4.185 $Y=1.99 $X2=0 $Y2=0
cc_546 N_SET_B_c_581_n N_VPWR_c_1232_n 0.0215763f $X=5.885 $Y=1.59 $X2=0 $Y2=0
cc_547 N_SET_B_M1025_g N_VPWR_c_1233_n 0.00415721f $X=4.165 $Y=2.525 $X2=0 $Y2=0
cc_548 N_SET_B_M1021_g N_VPWR_c_1234_n 0.0016085f $X=7.83 $Y=2.525 $X2=0 $Y2=0
cc_549 N_SET_B_M1021_g N_VPWR_c_1235_n 0.00331863f $X=7.83 $Y=2.525 $X2=0 $Y2=0
cc_550 N_SET_B_c_572_n N_VPWR_c_1241_n 9.83618e-19 $X=7.44 $Y=1.41 $X2=0 $Y2=0
cc_551 N_SET_B_M1025_g N_VPWR_c_1228_n 9.39239e-19 $X=4.165 $Y=2.525 $X2=0 $Y2=0
cc_552 N_SET_B_M1021_g N_VPWR_c_1228_n 9.39239e-19 $X=7.83 $Y=2.525 $X2=0 $Y2=0
cc_553 N_SET_B_c_581_n N_A_985_379#_M1007_d 0.00239457f $X=5.885 $Y=1.59
+ $X2=-0.19 $Y2=-0.245
cc_554 N_SET_B_c_581_n N_A_985_379#_c_1414_n 0.0220026f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_555 N_SET_B_c_581_n N_A_1092_417#_c_1440_n 0.0221533f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_556 N_SET_B_c_581_n N_A_1092_417#_c_1443_n 0.00402723f $X=5.885 $Y=1.59 $X2=0
+ $Y2=0
cc_557 N_SET_B_M1008_g N_VGND_c_1486_n 0.00952745f $X=7.08 $Y=0.665 $X2=0 $Y2=0
cc_558 N_SET_B_c_571_n N_VGND_c_1490_n 0.00486043f $X=4.64 $Y=0.765 $X2=0 $Y2=0
cc_559 N_SET_B_M1008_g N_VGND_c_1491_n 0.00429764f $X=7.08 $Y=0.665 $X2=0 $Y2=0
cc_560 N_SET_B_M1008_g N_VGND_c_1494_n 0.00435987f $X=7.08 $Y=0.665 $X2=0 $Y2=0
cc_561 N_SET_B_c_567_n N_VGND_c_1494_n 0.00667388f $X=4.44 $Y=0.97 $X2=0 $Y2=0
cc_562 N_SET_B_c_568_n N_VGND_c_1494_n 0.0054653f $X=4.64 $Y=0.93 $X2=0 $Y2=0
cc_563 N_SET_B_c_571_n N_VGND_c_1494_n 0.00444257f $X=4.64 $Y=0.765 $X2=0 $Y2=0
cc_564 N_SET_B_c_568_n N_VGND_c_1498_n 0.011981f $X=4.64 $Y=0.93 $X2=0 $Y2=0
cc_565 N_SET_B_c_569_n N_VGND_c_1498_n 0.00643657f $X=4.64 $Y=0.93 $X2=0 $Y2=0
cc_566 N_SET_B_c_571_n N_VGND_c_1498_n 0.0176324f $X=4.64 $Y=0.765 $X2=0 $Y2=0
cc_567 N_A_486_119#_c_739_n N_A_33_463#_c_854_n 0.00325473f $X=2.84 $Y=2.52
+ $X2=0 $Y2=0
cc_568 N_A_486_119#_c_730_n N_A_33_463#_M1028_g 0.00407425f $X=2.755 $Y=0.81
+ $X2=0 $Y2=0
cc_569 N_A_486_119#_c_704_n N_A_33_463#_M1028_g 5.14308e-19 $X=2.84 $Y=1.555
+ $X2=0 $Y2=0
cc_570 N_A_486_119#_c_709_n N_A_33_463#_M1020_g 0.00664889f $X=2.84 $Y=2.355
+ $X2=0 $Y2=0
cc_571 N_A_486_119#_c_739_n N_A_33_463#_M1020_g 0.00904011f $X=2.84 $Y=2.52
+ $X2=0 $Y2=0
cc_572 N_A_486_119#_M1003_g N_A_33_463#_c_857_n 0.0101666f $X=3.735 $Y=2.525
+ $X2=0 $Y2=0
cc_573 N_A_486_119#_M1007_g N_A_33_463#_c_857_n 0.0103024f $X=4.85 $Y=2.315
+ $X2=0 $Y2=0
cc_574 N_A_486_119#_c_702_n N_A_1175_417#_c_1078_n 0.00172593f $X=5.475 $Y=0.985
+ $X2=0 $Y2=0
cc_575 N_A_486_119#_c_702_n N_A_1175_417#_c_1080_n 8.99128e-19 $X=5.475 $Y=0.985
+ $X2=0 $Y2=0
cc_576 N_A_486_119#_M1003_g N_VPWR_c_1231_n 0.00746904f $X=3.735 $Y=2.525 $X2=0
+ $Y2=0
cc_577 N_A_486_119#_M1007_g N_VPWR_c_1233_n 0.00258018f $X=4.85 $Y=2.315 $X2=0
+ $Y2=0
cc_578 N_A_486_119#_c_739_n N_VPWR_c_1237_n 0.00709383f $X=2.84 $Y=2.52 $X2=0
+ $Y2=0
cc_579 N_A_486_119#_M1003_g N_VPWR_c_1228_n 9.39239e-19 $X=3.735 $Y=2.525 $X2=0
+ $Y2=0
cc_580 N_A_486_119#_M1007_g N_VPWR_c_1228_n 7.82699e-19 $X=4.85 $Y=2.315 $X2=0
+ $Y2=0
cc_581 N_A_486_119#_c_739_n N_VPWR_c_1228_n 0.0115646f $X=2.84 $Y=2.52 $X2=0
+ $Y2=0
cc_582 N_A_486_119#_c_704_n N_A_400_119#_c_1363_n 0.00554507f $X=2.84 $Y=1.555
+ $X2=0 $Y2=0
cc_583 N_A_486_119#_c_709_n N_A_400_119#_c_1366_n 0.00487418f $X=2.84 $Y=2.355
+ $X2=0 $Y2=0
cc_584 N_A_486_119#_c_704_n N_A_400_119#_c_1364_n 0.0140774f $X=2.84 $Y=1.555
+ $X2=0 $Y2=0
cc_585 N_A_486_119#_c_709_n N_A_400_119#_c_1364_n 0.0209364f $X=2.84 $Y=2.355
+ $X2=0 $Y2=0
cc_586 N_A_486_119#_c_711_n N_A_400_119#_c_1364_n 0.0128674f $X=2.84 $Y=1.64
+ $X2=0 $Y2=0
cc_587 N_A_486_119#_c_730_n N_A_400_119#_c_1365_n 0.00881685f $X=2.755 $Y=0.81
+ $X2=0 $Y2=0
cc_588 N_A_486_119#_c_704_n N_A_400_119#_c_1365_n 0.0115092f $X=2.84 $Y=1.555
+ $X2=0 $Y2=0
cc_589 N_A_486_119#_c_709_n N_A_400_119#_c_1368_n 0.0133057f $X=2.84 $Y=2.355
+ $X2=0 $Y2=0
cc_590 N_A_486_119#_c_739_n N_A_400_119#_c_1368_n 0.00684858f $X=2.84 $Y=2.52
+ $X2=0 $Y2=0
cc_591 N_A_486_119#_M1007_g N_A_985_379#_c_1414_n 0.00990962f $X=4.85 $Y=2.315
+ $X2=0 $Y2=0
cc_592 N_A_486_119#_M1007_g N_A_985_379#_c_1415_n 0.0012693f $X=4.85 $Y=2.315
+ $X2=0 $Y2=0
cc_593 N_A_486_119#_M1027_g N_VGND_c_1485_n 0.00354944f $X=4.19 $Y=0.445 $X2=0
+ $Y2=0
cc_594 N_A_486_119#_c_730_n N_VGND_c_1485_n 0.00568777f $X=2.755 $Y=0.81 $X2=0
+ $Y2=0
cc_595 N_A_486_119#_c_730_n N_VGND_c_1489_n 0.00773276f $X=2.755 $Y=0.81 $X2=0
+ $Y2=0
cc_596 N_A_486_119#_M1027_g N_VGND_c_1490_n 0.00585385f $X=4.19 $Y=0.445 $X2=0
+ $Y2=0
cc_597 N_A_486_119#_c_702_n N_VGND_c_1491_n 0.00486043f $X=5.475 $Y=0.985 $X2=0
+ $Y2=0
cc_598 N_A_486_119#_M1027_g N_VGND_c_1494_n 0.0122126f $X=4.19 $Y=0.445 $X2=0
+ $Y2=0
cc_599 N_A_486_119#_c_702_n N_VGND_c_1494_n 0.00813827f $X=5.475 $Y=0.985 $X2=0
+ $Y2=0
cc_600 N_A_486_119#_c_730_n N_VGND_c_1494_n 0.0149813f $X=2.755 $Y=0.81 $X2=0
+ $Y2=0
cc_601 N_A_486_119#_M1027_g N_VGND_c_1498_n 0.00235615f $X=4.19 $Y=0.445 $X2=0
+ $Y2=0
cc_602 N_A_486_119#_c_701_n N_VGND_c_1498_n 0.0168315f $X=5.165 $Y=1.06 $X2=0
+ $Y2=0
cc_603 N_A_486_119#_c_702_n N_VGND_c_1498_n 0.0174752f $X=5.475 $Y=0.985 $X2=0
+ $Y2=0
cc_604 N_A_486_119#_c_730_n A_572_119# 0.004104f $X=2.755 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_605 N_A_486_119#_c_704_n A_572_119# 3.3084e-19 $X=2.84 $Y=1.555 $X2=-0.19
+ $Y2=-0.245
cc_606 N_A_33_463#_M1014_g N_A_1329_65#_M1015_g 0.052164f $X=6.36 $Y=0.665 $X2=0
+ $Y2=0
cc_607 N_A_33_463#_M1004_g N_A_1329_65#_c_985_n 0.0169034f $X=6.325 $Y=2.505
+ $X2=0 $Y2=0
cc_608 N_A_33_463#_c_857_n N_A_1329_65#_c_987_n 0.0169034f $X=6.25 $Y=3.15 $X2=0
+ $Y2=0
cc_609 N_A_33_463#_M1004_g N_A_1329_65#_c_990_n 0.00210997f $X=6.325 $Y=2.505
+ $X2=0 $Y2=0
cc_610 N_A_33_463#_c_861_n N_A_1329_65#_c_990_n 0.052164f $X=6.342 $Y=1.975
+ $X2=0 $Y2=0
cc_611 N_A_33_463#_M1014_g N_A_1175_417#_c_1078_n 0.0138293f $X=6.36 $Y=0.665
+ $X2=0 $Y2=0
cc_612 N_A_33_463#_M1014_g N_A_1175_417#_c_1079_n 0.0107724f $X=6.36 $Y=0.665
+ $X2=0 $Y2=0
cc_613 N_A_33_463#_M1014_g N_A_1175_417#_c_1080_n 0.00308349f $X=6.36 $Y=0.665
+ $X2=0 $Y2=0
cc_614 N_A_33_463#_M1004_g N_A_1175_417#_c_1108_n 0.0104863f $X=6.325 $Y=2.505
+ $X2=0 $Y2=0
cc_615 N_A_33_463#_M1024_g N_VPWR_c_1229_n 0.0132707f $X=0.935 $Y=2.635 $X2=0
+ $Y2=0
cc_616 N_A_33_463#_c_855_n N_VPWR_c_1229_n 0.00720415f $X=1.01 $Y=3.15 $X2=0
+ $Y2=0
cc_617 N_A_33_463#_c_862_n N_VPWR_c_1229_n 0.0252688f $X=0.29 $Y=2.46 $X2=0
+ $Y2=0
cc_618 N_A_33_463#_c_849_n N_VPWR_c_1229_n 0.0110562f $X=0.7 $Y=1.645 $X2=0
+ $Y2=0
cc_619 N_A_33_463#_c_852_n N_VPWR_c_1229_n 0.0053015f $X=0.935 $Y=1.645 $X2=0
+ $Y2=0
cc_620 N_A_33_463#_M1024_g N_VPWR_c_1230_n 0.00396098f $X=0.935 $Y=2.635 $X2=0
+ $Y2=0
cc_621 N_A_33_463#_c_854_n N_VPWR_c_1230_n 0.0243917f $X=2.76 $Y=3.15 $X2=0
+ $Y2=0
cc_622 N_A_33_463#_M1020_g N_VPWR_c_1231_n 0.0063877f $X=2.835 $Y=2.525 $X2=0
+ $Y2=0
cc_623 N_A_33_463#_c_857_n N_VPWR_c_1231_n 0.0235458f $X=6.25 $Y=3.15 $X2=0
+ $Y2=0
cc_624 N_A_33_463#_c_857_n N_VPWR_c_1233_n 0.0326657f $X=6.25 $Y=3.15 $X2=0
+ $Y2=0
cc_625 N_A_33_463#_c_854_n N_VPWR_c_1237_n 0.0432727f $X=2.76 $Y=3.15 $X2=0
+ $Y2=0
cc_626 N_A_33_463#_c_857_n N_VPWR_c_1239_n 0.037049f $X=6.25 $Y=3.15 $X2=0 $Y2=0
cc_627 N_A_33_463#_c_862_n N_VPWR_c_1242_n 0.0127518f $X=0.29 $Y=2.46 $X2=0
+ $Y2=0
cc_628 N_A_33_463#_c_855_n N_VPWR_c_1243_n 0.0233436f $X=1.01 $Y=3.15 $X2=0
+ $Y2=0
cc_629 N_A_33_463#_c_857_n N_VPWR_c_1244_n 0.0209676f $X=6.25 $Y=3.15 $X2=0
+ $Y2=0
cc_630 N_A_33_463#_c_854_n N_VPWR_c_1228_n 0.0521499f $X=2.76 $Y=3.15 $X2=0
+ $Y2=0
cc_631 N_A_33_463#_c_855_n N_VPWR_c_1228_n 0.00811614f $X=1.01 $Y=3.15 $X2=0
+ $Y2=0
cc_632 N_A_33_463#_c_857_n N_VPWR_c_1228_n 0.0836396f $X=6.25 $Y=3.15 $X2=0
+ $Y2=0
cc_633 N_A_33_463#_c_860_n N_VPWR_c_1228_n 0.00433536f $X=2.835 $Y=3.15 $X2=0
+ $Y2=0
cc_634 N_A_33_463#_c_862_n N_VPWR_c_1228_n 0.0110892f $X=0.29 $Y=2.46 $X2=0
+ $Y2=0
cc_635 N_A_33_463#_c_844_n N_A_400_119#_c_1363_n 0.00306975f $X=2.28 $Y=0.18
+ $X2=0 $Y2=0
cc_636 N_A_33_463#_M1028_g N_A_400_119#_c_1363_n 0.00163937f $X=2.355 $Y=0.805
+ $X2=0 $Y2=0
cc_637 N_A_33_463#_c_854_n N_A_400_119#_c_1366_n 0.00383069f $X=2.76 $Y=3.15
+ $X2=0 $Y2=0
cc_638 N_A_33_463#_M1028_g N_A_400_119#_c_1365_n 0.00381956f $X=2.355 $Y=0.805
+ $X2=0 $Y2=0
cc_639 N_A_33_463#_c_857_n N_A_985_379#_c_1415_n 0.00774103f $X=6.25 $Y=3.15
+ $X2=0 $Y2=0
cc_640 N_A_33_463#_c_857_n N_A_985_379#_c_1416_n 0.0200606f $X=6.25 $Y=3.15
+ $X2=0 $Y2=0
cc_641 N_A_33_463#_M1004_g N_A_985_379#_c_1416_n 0.0160197f $X=6.325 $Y=2.505
+ $X2=0 $Y2=0
cc_642 N_A_33_463#_M1004_g N_A_1092_417#_c_1440_n 5.54749e-19 $X=6.325 $Y=2.505
+ $X2=0 $Y2=0
cc_643 N_A_33_463#_M1004_g N_A_1092_417#_c_1443_n 0.0119077f $X=6.325 $Y=2.505
+ $X2=0 $Y2=0
cc_644 N_A_33_463#_c_845_n N_VGND_c_1483_n 0.00844007f $X=1.05 $Y=0.18 $X2=0
+ $Y2=0
cc_645 N_A_33_463#_M1018_g N_VGND_c_1484_n 0.0049891f $X=0.975 $Y=0.58 $X2=0
+ $Y2=0
cc_646 N_A_33_463#_c_844_n N_VGND_c_1484_n 0.0241897f $X=2.28 $Y=0.18 $X2=0
+ $Y2=0
cc_647 N_A_33_463#_M1028_g N_VGND_c_1484_n 0.00610494f $X=2.355 $Y=0.805 $X2=0
+ $Y2=0
cc_648 N_A_33_463#_c_845_n N_VGND_c_1488_n 0.0195697f $X=1.05 $Y=0.18 $X2=0
+ $Y2=0
cc_649 N_A_33_463#_c_844_n N_VGND_c_1489_n 0.0189195f $X=2.28 $Y=0.18 $X2=0
+ $Y2=0
cc_650 N_A_33_463#_M1014_g N_VGND_c_1491_n 0.00462152f $X=6.36 $Y=0.665 $X2=0
+ $Y2=0
cc_651 N_A_33_463#_c_844_n N_VGND_c_1494_n 0.0429268f $X=2.28 $Y=0.18 $X2=0
+ $Y2=0
cc_652 N_A_33_463#_c_845_n N_VGND_c_1494_n 0.0111932f $X=1.05 $Y=0.18 $X2=0
+ $Y2=0
cc_653 N_A_33_463#_M1014_g N_VGND_c_1494_n 0.00453288f $X=6.36 $Y=0.665 $X2=0
+ $Y2=0
cc_654 N_A_33_463#_c_850_n N_VGND_c_1494_n 0.0140092f $X=0.33 $Y=0.555 $X2=0
+ $Y2=0
cc_655 N_A_33_463#_c_850_n N_VGND_c_1495_n 0.0133721f $X=0.33 $Y=0.555 $X2=0
+ $Y2=0
cc_656 N_A_1329_65#_c_983_n N_A_1175_417#_c_1069_n 0.00530795f $X=7.825 $Y=0.4
+ $X2=0 $Y2=0
cc_657 N_A_1329_65#_c_981_n N_A_1175_417#_c_1070_n 0.00776126f $X=8.65 $Y=0.4
+ $X2=0 $Y2=0
cc_658 N_A_1329_65#_c_983_n N_A_1175_417#_c_1070_n 0.00899666f $X=7.825 $Y=0.4
+ $X2=0 $Y2=0
cc_659 N_A_1329_65#_c_983_n N_A_1175_417#_c_1071_n 2.83293e-19 $X=7.825 $Y=0.4
+ $X2=0 $Y2=0
cc_660 N_A_1329_65#_c_982_n N_A_1175_417#_M1010_g 0.0123917f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_661 N_A_1329_65#_c_993_n N_A_1175_417#_M1010_g 0.00333207f $X=8.745 $Y=2.56
+ $X2=0 $Y2=0
cc_662 N_A_1329_65#_c_982_n N_A_1175_417#_c_1073_n 0.0201771f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_663 N_A_1329_65#_c_982_n N_A_1175_417#_c_1074_n 0.00323914f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_664 N_A_1329_65#_c_982_n N_A_1175_417#_M1026_g 0.00335744f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_665 N_A_1329_65#_c_993_n N_A_1175_417#_M1026_g 0.00307517f $X=8.745 $Y=2.56
+ $X2=0 $Y2=0
cc_666 N_A_1329_65#_M1015_g N_A_1175_417#_c_1078_n 0.00286555f $X=6.72 $Y=0.665
+ $X2=0 $Y2=0
cc_667 N_A_1329_65#_M1015_g N_A_1175_417#_c_1079_n 0.013786f $X=6.72 $Y=0.665
+ $X2=0 $Y2=0
cc_668 N_A_1329_65#_c_983_n N_A_1175_417#_c_1079_n 0.00658936f $X=7.825 $Y=0.4
+ $X2=0 $Y2=0
cc_669 N_A_1329_65#_c_985_n N_A_1175_417#_c_1086_n 0.0128608f $X=6.91 $Y=3.075
+ $X2=0 $Y2=0
cc_670 N_A_1329_65#_M1002_g N_A_1175_417#_c_1086_n 0.00984479f $X=7.4 $Y=2.525
+ $X2=0 $Y2=0
cc_671 N_A_1329_65#_c_990_n N_A_1175_417#_c_1086_n 0.00523991f $X=6.91 $Y=1.935
+ $X2=0 $Y2=0
cc_672 N_A_1329_65#_c_982_n N_A_1175_417#_c_1081_n 0.00833685f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_673 N_A_1329_65#_M1002_g N_A_1175_417#_c_1088_n 8.40754e-19 $X=7.4 $Y=2.525
+ $X2=0 $Y2=0
cc_674 N_A_1329_65#_c_989_n N_A_1175_417#_c_1088_n 0.00422438f $X=8.58 $Y=3.15
+ $X2=0 $Y2=0
cc_675 N_A_1329_65#_c_981_n N_A_1175_417#_c_1082_n 0.0289092f $X=8.65 $Y=0.4
+ $X2=0 $Y2=0
cc_676 N_A_1329_65#_c_982_n N_A_1175_417#_c_1082_n 0.0526375f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_677 N_A_1329_65#_c_983_n N_A_1175_417#_c_1082_n 0.0246181f $X=7.825 $Y=0.4
+ $X2=0 $Y2=0
cc_678 N_A_1329_65#_c_981_n N_A_1175_417#_c_1083_n 0.0136718f $X=8.65 $Y=0.4
+ $X2=0 $Y2=0
cc_679 N_A_1329_65#_c_982_n N_A_1175_417#_c_1083_n 0.00879973f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_680 N_A_1329_65#_c_983_n N_A_1175_417#_c_1083_n 0.0035906f $X=7.825 $Y=0.4
+ $X2=0 $Y2=0
cc_681 N_A_1329_65#_c_982_n N_A_1832_131#_c_1188_n 0.0449741f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_682 N_A_1329_65#_c_982_n N_A_1832_131#_c_1193_n 0.0628816f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_683 N_A_1329_65#_c_993_n N_A_1832_131#_c_1193_n 3.49476e-19 $X=8.745 $Y=2.56
+ $X2=0 $Y2=0
cc_684 N_A_1329_65#_c_982_n N_A_1832_131#_c_1191_n 0.0264953f $X=8.765 $Y=1.75
+ $X2=0 $Y2=0
cc_685 N_A_1329_65#_M1002_g N_VPWR_c_1234_n 0.0112141f $X=7.4 $Y=2.525 $X2=0
+ $Y2=0
cc_686 N_A_1329_65#_c_989_n N_VPWR_c_1234_n 0.0153703f $X=8.58 $Y=3.15 $X2=0
+ $Y2=0
cc_687 N_A_1329_65#_c_989_n N_VPWR_c_1235_n 0.0158587f $X=8.58 $Y=3.15 $X2=0
+ $Y2=0
cc_688 N_A_1329_65#_c_993_n N_VPWR_c_1235_n 0.0108989f $X=8.745 $Y=2.56 $X2=0
+ $Y2=0
cc_689 N_A_1329_65#_c_982_n N_VPWR_c_1236_n 0.0191763f $X=8.765 $Y=1.75 $X2=0
+ $Y2=0
cc_690 N_A_1329_65#_c_993_n N_VPWR_c_1236_n 0.00514956f $X=8.745 $Y=2.56 $X2=0
+ $Y2=0
cc_691 N_A_1329_65#_c_987_n N_VPWR_c_1239_n 0.0210917f $X=6.985 $Y=3.15 $X2=0
+ $Y2=0
cc_692 N_A_1329_65#_c_982_n N_VPWR_c_1241_n 0.0945019f $X=8.765 $Y=1.75 $X2=0
+ $Y2=0
cc_693 N_A_1329_65#_c_989_n N_VPWR_c_1245_n 0.0187498f $X=8.58 $Y=3.15 $X2=0
+ $Y2=0
cc_694 N_A_1329_65#_c_989_n N_VPWR_c_1246_n 0.0128089f $X=8.58 $Y=3.15 $X2=0
+ $Y2=0
cc_695 N_A_1329_65#_c_982_n N_VPWR_c_1246_n 0.0178471f $X=8.765 $Y=1.75 $X2=0
+ $Y2=0
cc_696 N_A_1329_65#_c_986_n N_VPWR_c_1228_n 0.00953891f $X=7.325 $Y=3.15 $X2=0
+ $Y2=0
cc_697 N_A_1329_65#_c_987_n N_VPWR_c_1228_n 0.00564429f $X=6.985 $Y=3.15 $X2=0
+ $Y2=0
cc_698 N_A_1329_65#_c_989_n N_VPWR_c_1228_n 0.0450714f $X=8.58 $Y=3.15 $X2=0
+ $Y2=0
cc_699 N_A_1329_65#_c_991_n N_VPWR_c_1228_n 0.00833318f $X=7.4 $Y=3.15 $X2=0
+ $Y2=0
cc_700 N_A_1329_65#_c_982_n N_VPWR_c_1228_n 0.00956371f $X=8.765 $Y=1.75 $X2=0
+ $Y2=0
cc_701 N_A_1329_65#_c_985_n N_A_985_379#_c_1416_n 0.00819404f $X=6.91 $Y=3.075
+ $X2=0 $Y2=0
cc_702 N_A_1329_65#_c_985_n N_A_1092_417#_c_1442_n 0.00169146f $X=6.91 $Y=3.075
+ $X2=0 $Y2=0
cc_703 N_A_1329_65#_c_986_n N_A_1092_417#_c_1442_n 0.00281234f $X=7.325 $Y=3.15
+ $X2=0 $Y2=0
cc_704 N_A_1329_65#_M1002_g N_A_1092_417#_c_1442_n 0.00325423f $X=7.4 $Y=2.525
+ $X2=0 $Y2=0
cc_705 N_A_1329_65#_c_985_n N_A_1092_417#_c_1443_n 0.0134041f $X=6.91 $Y=3.075
+ $X2=0 $Y2=0
cc_706 N_A_1329_65#_M1015_g N_VGND_c_1486_n 0.00205641f $X=6.72 $Y=0.665 $X2=0
+ $Y2=0
cc_707 N_A_1329_65#_c_983_n N_VGND_c_1486_n 0.0189622f $X=7.825 $Y=0.4 $X2=0
+ $Y2=0
cc_708 N_A_1329_65#_c_981_n N_VGND_c_1487_n 0.00598222f $X=8.65 $Y=0.4 $X2=0
+ $Y2=0
cc_709 N_A_1329_65#_c_982_n N_VGND_c_1487_n 0.00631443f $X=8.765 $Y=1.75 $X2=0
+ $Y2=0
cc_710 N_A_1329_65#_M1015_g N_VGND_c_1491_n 0.00517164f $X=6.72 $Y=0.665 $X2=0
+ $Y2=0
cc_711 N_A_1329_65#_c_981_n N_VGND_c_1492_n 0.0441249f $X=8.65 $Y=0.4 $X2=0
+ $Y2=0
cc_712 N_A_1329_65#_c_983_n N_VGND_c_1492_n 0.0154368f $X=7.825 $Y=0.4 $X2=0
+ $Y2=0
cc_713 N_A_1329_65#_M1015_g N_VGND_c_1494_n 0.00519032f $X=6.72 $Y=0.665 $X2=0
+ $Y2=0
cc_714 N_A_1329_65#_c_981_n N_VGND_c_1494_n 0.0321349f $X=8.65 $Y=0.4 $X2=0
+ $Y2=0
cc_715 N_A_1329_65#_c_983_n N_VGND_c_1494_n 0.0105988f $X=7.825 $Y=0.4 $X2=0
+ $Y2=0
cc_716 N_A_1175_417#_c_1074_n N_A_1832_131#_M1000_g 0.0173766f $X=9.5 $Y=1.185
+ $X2=0 $Y2=0
cc_717 N_A_1175_417#_M1026_g N_A_1832_131#_M1006_g 0.0195898f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_718 N_A_1175_417#_c_1073_n N_A_1832_131#_c_1188_n 0.0122892f $X=9.425 $Y=1.26
+ $X2=0 $Y2=0
cc_719 N_A_1175_417#_c_1074_n N_A_1832_131#_c_1188_n 0.00450458f $X=9.5 $Y=1.185
+ $X2=0 $Y2=0
cc_720 N_A_1175_417#_M1026_g N_A_1832_131#_c_1193_n 0.00785299f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_721 N_A_1175_417#_c_1073_n N_A_1832_131#_c_1189_n 0.00163492f $X=9.425
+ $Y=1.26 $X2=0 $Y2=0
cc_722 N_A_1175_417#_M1026_g N_A_1832_131#_c_1189_n 0.020029f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_723 N_A_1175_417#_c_1077_n N_A_1832_131#_c_1189_n 0.00741485f $X=9.5 $Y=1.26
+ $X2=0 $Y2=0
cc_724 N_A_1175_417#_c_1077_n N_A_1832_131#_c_1190_n 0.0213342f $X=9.5 $Y=1.26
+ $X2=0 $Y2=0
cc_725 N_A_1175_417#_c_1073_n N_A_1832_131#_c_1191_n 0.00599512f $X=9.425
+ $Y=1.26 $X2=0 $Y2=0
cc_726 N_A_1175_417#_c_1086_n N_VPWR_c_1234_n 0.0138021f $X=7.775 $Y=2.18 $X2=0
+ $Y2=0
cc_727 N_A_1175_417#_M1010_g N_VPWR_c_1235_n 0.0047141f $X=8.55 $Y=1.815 $X2=0
+ $Y2=0
cc_728 N_A_1175_417#_c_1081_n N_VPWR_c_1235_n 0.00968185f $X=7.912 $Y=2.095
+ $X2=0 $Y2=0
cc_729 N_A_1175_417#_c_1088_n N_VPWR_c_1235_n 0.0324819f $X=8.045 $Y=2.525 $X2=0
+ $Y2=0
cc_730 N_A_1175_417#_c_1089_n N_VPWR_c_1235_n 0.0143577f $X=7.957 $Y=2.18 $X2=0
+ $Y2=0
cc_731 N_A_1175_417#_M1026_g N_VPWR_c_1236_n 0.0221348f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_732 N_A_1175_417#_M1010_g N_VPWR_c_1241_n 0.00342887f $X=8.55 $Y=1.815 $X2=0
+ $Y2=0
cc_733 N_A_1175_417#_c_1076_n N_VPWR_c_1241_n 0.00177848f $X=8.385 $Y=1.26 $X2=0
+ $Y2=0
cc_734 N_A_1175_417#_c_1081_n N_VPWR_c_1241_n 0.025793f $X=7.912 $Y=2.095 $X2=0
+ $Y2=0
cc_735 N_A_1175_417#_c_1082_n N_VPWR_c_1241_n 0.0159768f $X=7.912 $Y=1 $X2=0
+ $Y2=0
cc_736 N_A_1175_417#_c_1088_n N_VPWR_c_1245_n 0.00432583f $X=8.045 $Y=2.525
+ $X2=0 $Y2=0
cc_737 N_A_1175_417#_M1026_g N_VPWR_c_1246_n 0.00280576f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_738 N_A_1175_417#_M1026_g N_VPWR_c_1228_n 0.00371991f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_739 N_A_1175_417#_c_1088_n N_VPWR_c_1228_n 0.00672715f $X=8.045 $Y=2.525
+ $X2=0 $Y2=0
cc_740 N_A_1175_417#_c_1086_n N_A_985_379#_M1004_d 0.00739738f $X=7.775 $Y=2.18
+ $X2=0 $Y2=0
cc_741 N_A_1175_417#_M1013_d N_A_985_379#_c_1416_n 0.00265888f $X=5.875 $Y=2.085
+ $X2=0 $Y2=0
cc_742 N_A_1175_417#_c_1086_n N_A_1092_417#_c_1442_n 0.0226634f $X=7.775 $Y=2.18
+ $X2=0 $Y2=0
cc_743 N_A_1175_417#_M1013_d N_A_1092_417#_c_1443_n 0.00481321f $X=5.875
+ $Y=2.085 $X2=0 $Y2=0
cc_744 N_A_1175_417#_c_1086_n N_A_1092_417#_c_1443_n 0.0322666f $X=7.775 $Y=2.18
+ $X2=0 $Y2=0
cc_745 N_A_1175_417#_c_1106_n N_A_1092_417#_c_1443_n 0.0297041f $X=6.235 $Y=2.21
+ $X2=0 $Y2=0
cc_746 N_A_1175_417#_c_1071_n N_VGND_c_1486_n 0.00840698f $X=7.665 $Y=0.27 $X2=0
+ $Y2=0
cc_747 N_A_1175_417#_c_1079_n N_VGND_c_1486_n 0.0243206f $X=7.775 $Y=0.99 $X2=0
+ $Y2=0
cc_748 N_A_1175_417#_c_1074_n N_VGND_c_1487_n 0.0102915f $X=9.5 $Y=1.185 $X2=0
+ $Y2=0
cc_749 N_A_1175_417#_c_1078_n N_VGND_c_1491_n 0.0230821f $X=6.05 $Y=0.39 $X2=0
+ $Y2=0
cc_750 N_A_1175_417#_c_1071_n N_VGND_c_1492_n 0.0208194f $X=7.665 $Y=0.27 $X2=0
+ $Y2=0
cc_751 N_A_1175_417#_c_1074_n N_VGND_c_1492_n 0.00385681f $X=9.5 $Y=1.185 $X2=0
+ $Y2=0
cc_752 N_A_1175_417#_M1031_d N_VGND_c_1494_n 0.00216391f $X=5.91 $Y=0.235 $X2=0
+ $Y2=0
cc_753 N_A_1175_417#_c_1070_n N_VGND_c_1494_n 0.0206743f $X=8.145 $Y=0.27 $X2=0
+ $Y2=0
cc_754 N_A_1175_417#_c_1071_n N_VGND_c_1494_n 0.00984503f $X=7.665 $Y=0.27 $X2=0
+ $Y2=0
cc_755 N_A_1175_417#_c_1074_n N_VGND_c_1494_n 0.0044892f $X=9.5 $Y=1.185 $X2=0
+ $Y2=0
cc_756 N_A_1175_417#_c_1078_n N_VGND_c_1494_n 0.0158284f $X=6.05 $Y=0.39 $X2=0
+ $Y2=0
cc_757 N_A_1175_417#_c_1078_n N_VGND_c_1498_n 0.0211948f $X=6.05 $Y=0.39 $X2=0
+ $Y2=0
cc_758 N_A_1832_131#_M1006_g N_VPWR_c_1236_n 0.0296406f $X=10.085 $Y=2.465 $X2=0
+ $Y2=0
cc_759 N_A_1832_131#_c_1193_n N_VPWR_c_1236_n 0.02691f $X=9.285 $Y=1.98 $X2=0
+ $Y2=0
cc_760 N_A_1832_131#_c_1189_n N_VPWR_c_1236_n 0.0389112f $X=9.95 $Y=1.48 $X2=0
+ $Y2=0
cc_761 N_A_1832_131#_c_1190_n N_VPWR_c_1236_n 0.00550832f $X=9.95 $Y=1.48 $X2=0
+ $Y2=0
cc_762 N_A_1832_131#_M1006_g N_VPWR_c_1247_n 0.00486043f $X=10.085 $Y=2.465
+ $X2=0 $Y2=0
cc_763 N_A_1832_131#_M1006_g N_VPWR_c_1228_n 0.00917987f $X=10.085 $Y=2.465
+ $X2=0 $Y2=0
cc_764 N_A_1832_131#_c_1193_n N_VPWR_c_1228_n 0.0105212f $X=9.285 $Y=1.98 $X2=0
+ $Y2=0
cc_765 N_A_1832_131#_M1000_g N_Q_c_1467_n 0.0028883f $X=10.01 $Y=0.655 $X2=0
+ $Y2=0
cc_766 N_A_1832_131#_c_1190_n N_Q_c_1467_n 0.00293445f $X=9.95 $Y=1.48 $X2=0
+ $Y2=0
cc_767 N_A_1832_131#_M1000_g Q 0.00836651f $X=10.01 $Y=0.655 $X2=0 $Y2=0
cc_768 N_A_1832_131#_c_1189_n Q 0.0271104f $X=9.95 $Y=1.48 $X2=0 $Y2=0
cc_769 N_A_1832_131#_c_1190_n Q 0.0188468f $X=9.95 $Y=1.48 $X2=0 $Y2=0
cc_770 N_A_1832_131#_M1000_g N_VGND_c_1487_n 0.00800888f $X=10.01 $Y=0.655 $X2=0
+ $Y2=0
cc_771 N_A_1832_131#_c_1188_n N_VGND_c_1487_n 0.0150529f $X=9.285 $Y=0.865 $X2=0
+ $Y2=0
cc_772 N_A_1832_131#_c_1189_n N_VGND_c_1487_n 0.0254204f $X=9.95 $Y=1.48 $X2=0
+ $Y2=0
cc_773 N_A_1832_131#_c_1190_n N_VGND_c_1487_n 0.00315416f $X=9.95 $Y=1.48 $X2=0
+ $Y2=0
cc_774 N_A_1832_131#_c_1188_n N_VGND_c_1492_n 0.00436993f $X=9.285 $Y=0.865
+ $X2=0 $Y2=0
cc_775 N_A_1832_131#_M1000_g N_VGND_c_1493_n 0.00585385f $X=10.01 $Y=0.655 $X2=0
+ $Y2=0
cc_776 N_A_1832_131#_M1000_g N_VGND_c_1494_n 0.0128183f $X=10.01 $Y=0.655 $X2=0
+ $Y2=0
cc_777 N_A_1832_131#_c_1188_n N_VGND_c_1494_n 0.00775106f $X=9.285 $Y=0.865
+ $X2=0 $Y2=0
cc_778 N_VPWR_c_1237_n N_A_400_119#_c_1366_n 0.00359983f $X=3.295 $Y=3.33 $X2=0
+ $Y2=0
cc_779 N_VPWR_c_1228_n N_A_400_119#_c_1366_n 0.00564431f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_780 N_VPWR_c_1233_n N_A_985_379#_c_1414_n 0.0139526f $X=4.507 $Y=3.245 $X2=0
+ $Y2=0
cc_781 N_VPWR_c_1233_n N_A_985_379#_c_1415_n 0.0215578f $X=4.507 $Y=3.245 $X2=0
+ $Y2=0
cc_782 N_VPWR_c_1239_n N_A_985_379#_c_1415_n 0.0224969f $X=7.53 $Y=3.33 $X2=0
+ $Y2=0
cc_783 N_VPWR_c_1228_n N_A_985_379#_c_1415_n 0.0113197f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_784 N_VPWR_c_1239_n N_A_985_379#_c_1416_n 0.10281f $X=7.53 $Y=3.33 $X2=0
+ $Y2=0
cc_785 N_VPWR_c_1228_n N_A_985_379#_c_1416_n 0.0546904f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_786 N_VPWR_c_1239_n N_A_1092_417#_c_1443_n 0.00854806f $X=7.53 $Y=3.33 $X2=0
+ $Y2=0
cc_787 N_VPWR_c_1228_n N_A_1092_417#_c_1443_n 0.0151104f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_788 N_VPWR_c_1228_n N_Q_M1006_d 0.00371702f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_789 N_VPWR_c_1236_n Q 0.0499532f $X=9.775 $Y=2.02 $X2=0 $Y2=0
cc_790 N_VPWR_c_1247_n Q 0.018528f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_791 N_VPWR_c_1228_n Q 0.0104192f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_792 N_A_400_119#_c_1363_n N_VGND_c_1489_n 0.00361302f $X=2.14 $Y=0.805 $X2=0
+ $Y2=0
cc_793 N_A_400_119#_c_1363_n N_VGND_c_1494_n 0.00566138f $X=2.14 $Y=0.805 $X2=0
+ $Y2=0
cc_794 N_A_985_379#_c_1414_n N_A_1092_417#_c_1440_n 0.0284524f $X=5.065 $Y=2.22
+ $X2=0 $Y2=0
cc_795 N_A_985_379#_c_1414_n N_A_1092_417#_c_1441_n 0.0139f $X=5.065 $Y=2.22
+ $X2=0 $Y2=0
cc_796 N_A_985_379#_c_1416_n N_A_1092_417#_c_1441_n 0.0266401f $X=6.635 $Y=2.93
+ $X2=0 $Y2=0
cc_797 N_A_985_379#_M1004_d N_A_1092_417#_c_1443_n 0.00733131f $X=6.4 $Y=2.085
+ $X2=0 $Y2=0
cc_798 N_A_985_379#_c_1416_n N_A_1092_417#_c_1443_n 0.0665834f $X=6.635 $Y=2.93
+ $X2=0 $Y2=0
cc_799 N_Q_c_1467_n N_VGND_c_1487_n 0.00160678f $X=10.285 $Y=1.095 $X2=0 $Y2=0
cc_800 N_Q_c_1466_n N_VGND_c_1493_n 0.0251463f $X=10.225 $Y=0.42 $X2=0 $Y2=0
cc_801 N_Q_M1000_d N_VGND_c_1494_n 0.00249946f $X=10.085 $Y=0.235 $X2=0 $Y2=0
cc_802 N_Q_c_1466_n N_VGND_c_1494_n 0.0146958f $X=10.225 $Y=0.42 $X2=0 $Y2=0
cc_803 N_VGND_c_1494_n A_853_47# 0.00323522f $X=10.32 $Y=0 $X2=-0.19 $Y2=-0.245
cc_804 N_VGND_c_1494_n A_1110_47# 0.00899413f $X=10.32 $Y=0 $X2=-0.19 $Y2=-0.245
