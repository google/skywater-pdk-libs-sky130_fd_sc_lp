* File: sky130_fd_sc_lp__a21o_1.pex.spice
* Created: Wed Sep  2 09:19:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21O_1%A_80_237# 1 2 9 11 13 14 15 16 18 20 24 29
c54 14 0 1.87876e-19 $X=0.8 $Y=1.515
r55 35 37 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.475 $Y=1.35
+ $X2=0.48 $Y2=1.35
r56 29 37 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.69 $Y=1.35
+ $X2=0.48 $Y2=1.35
r57 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.35 $X2=0.69 $Y2=1.35
r58 22 24 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=1.555 $Y=0.985
+ $X2=1.555 $Y2=0.42
r59 18 30 23.4141 $w=1.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.18 $Y=2.01 $X2=0.8
+ $Y2=2.01
r60 18 20 34.5733 $w=2.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.18 $Y=2.1 $X2=1.18
+ $Y2=2.91
r61 17 28 11.8611 $w=2.88e-07 $l=3.58887e-07 $layer=LI1_cond $X=0.885 $Y=1.07
+ $X2=0.705 $Y2=1.35
r62 16 22 24.0951 $w=8e-08 $l=2.03101e-07 $layer=LI1_cond $X=1.39 $Y=1.07
+ $X2=1.555 $Y2=0.985
r63 16 17 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.39 $Y=1.07
+ $X2=0.885 $Y2=1.07
r64 15 30 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.8 $Y=1.92 $X2=0.8
+ $Y2=2.01
r65 14 28 9.02084 $w=2.88e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.8 $Y=1.515
+ $X2=0.705 $Y2=1.35
r66 14 15 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.8 $Y=1.515
+ $X2=0.8 $Y2=1.92
r67 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.185
+ $X2=0.48 $Y2=1.35
r68 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.48 $Y=1.185
+ $X2=0.48 $Y2=0.655
r69 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=1.35
r70 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=2.465
r71 2 18 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.21 $Y2=2.085
r72 2 20 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.21 $Y2=2.91
r73 1 24 91 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=2 $X=1.345
+ $Y=0.235 $X2=1.555 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_1%B1 3 7 9 12 13
c36 13 0 1.82227e-19 $X=1.29 $Y=1.51
c37 12 0 1.87876e-19 $X=1.29 $Y=1.51
r38 12 15 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.312 $Y=1.51
+ $X2=1.312 $Y2=1.675
r39 12 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.312 $Y=1.51
+ $X2=1.312 $Y2=1.345
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.29
+ $Y=1.51 $X2=1.29 $Y2=1.51
r41 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.51
r42 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.425 $Y=2.465
+ $X2=1.425 $Y2=1.675
r43 3 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.27 $Y=0.655
+ $X2=1.27 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_1%A1 3 6 8 9 10 15 17
c36 15 0 3.18426e-19 $X=1.905 $Y=1.35
r37 19 27 1.01705 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=2.097 $Y=1.185
+ $X2=2.097 $Y2=1.35
r38 16 27 6.70512 $w=3.28e-07 $l=1.92e-07 $layer=LI1_cond $X=1.905 $Y=1.35
+ $X2=2.097 $Y2=1.35
r39 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.35
+ $X2=1.905 $Y2=1.515
r40 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.35
+ $X2=1.905 $Y2=1.185
r41 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.905
+ $Y=1.35 $X2=1.905 $Y2=1.35
r42 10 27 2.20012 $w=3.28e-07 $l=6.3e-08 $layer=LI1_cond $X=2.16 $Y=1.35
+ $X2=2.097 $Y2=1.35
r43 9 19 9.51223 $w=3.13e-07 $l=2.6e-07 $layer=LI1_cond $X=2.097 $Y=0.925
+ $X2=2.097 $Y2=1.185
r44 8 9 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.097 $Y=0.555
+ $X2=2.097 $Y2=0.925
r45 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.855 $Y=2.465
+ $X2=1.855 $Y2=1.515
r46 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.815 $Y=0.655
+ $X2=1.815 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_1%A2 3 6 8 11 13
r23 11 14 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.492 $Y=1.35
+ $X2=2.492 $Y2=1.515
r24 11 13 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.492 $Y=1.35
+ $X2=2.492 $Y2=1.185
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.35 $X2=2.51 $Y2=1.35
r26 8 12 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=1.35 $X2=2.51
+ $Y2=1.35
r27 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.385 $Y=2.465
+ $X2=2.385 $Y2=1.515
r28 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.385 $Y=0.655
+ $X2=2.385 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_1%X 1 2 7 8 9 10 11 12 13 22
r12 13 40 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.225 $Y=2.775
+ $X2=0.225 $Y2=2.91
r13 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=2.405
+ $X2=0.225 $Y2=2.775
r14 11 12 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=0.225 $Y=1.98
+ $X2=0.225 $Y2=2.405
r15 10 11 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=1.98
r16 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r17 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r18 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.555
+ $X2=0.225 $Y2=0.925
r19 7 22 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.225 $Y=0.555
+ $X2=0.225 $Y2=0.42
r20 2 40 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r21 2 11 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
r22 1 22 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_1%VPWR 1 2 9 13 17 19 24 31 32 35 38
r39 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=2.125 $Y2=3.33
r44 29 31 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.29 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 25 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r48 25 27 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.96 $Y=3.33
+ $X2=2.125 $Y2=3.33
r50 24 27 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 19 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r54 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 17 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 17 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 13 16 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.125 $Y=2.11
+ $X2=2.125 $Y2=2.95
r58 11 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=3.33
r59 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=2.95
r60 7 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r61 7 9 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.355
r62 2 16 400 $w=1.7e-07 $l=1.20857e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.835 $X2=2.125 $Y2=2.95
r63 2 13 400 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.835 $X2=2.125 $Y2=2.11
r64 1 9 300 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_1%A_300_367# 1 2 9 13 14 17
c22 14 0 1.36199e-19 $X=1.745 $Y=1.77
r23 17 19 35.1401 $w=3.03e-07 $l=9.3e-07 $layer=LI1_cond $X=2.612 $Y=1.98
+ $X2=2.612 $Y2=2.91
r24 15 17 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=2.612 $Y=1.855
+ $X2=2.612 $Y2=1.98
r25 13 15 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=2.46 $Y=1.77
+ $X2=2.612 $Y2=1.855
r26 13 14 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.46 $Y=1.77
+ $X2=1.745 $Y2=1.77
r27 9 11 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.65 $Y=1.98 $X2=1.65
+ $Y2=2.91
r28 7 14 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.65 $Y=1.855
+ $X2=1.745 $Y2=1.77
r29 7 9 7.29665 $w=1.88e-07 $l=1.25e-07 $layer=LI1_cond $X=1.65 $Y=1.855
+ $X2=1.65 $Y2=1.98
r30 2 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.835 $X2=2.6 $Y2=2.91
r31 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.835 $X2=2.6 $Y2=1.98
r32 1 11 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=2.91
r33 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_1%VGND 1 2 9 11 13 15 17 22 28 34
r36 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r37 29 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r38 28 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r40 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r41 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 23 28 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=0.875
+ $Y2=0
r43 23 25 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=2.16
+ $Y2=0
r44 22 33 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.435 $Y=0 $X2=2.657
+ $Y2=0
r45 22 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.435 $Y=0 $X2=2.16
+ $Y2=0
r46 20 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 17 28 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.875
+ $Y2=0
r49 17 19 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.24
+ $Y2=0
r50 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r51 15 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r52 11 33 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.6 $Y=0.085
+ $X2=2.657 $Y2=0
r53 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.6 $Y=0.085
+ $X2=2.6 $Y2=0.38
r54 7 28 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=0.085
+ $X2=0.875 $Y2=0
r55 7 9 4.76698 $w=6.88e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=0.085
+ $X2=0.875 $Y2=0.36
r56 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.46
+ $Y=0.235 $X2=2.6 $Y2=0.38
r57 1 9 45.5 $w=1.7e-07 $l=5.59017e-07 $layer=licon1_NDIFF $count=4 $X=0.555
+ $Y=0.235 $X2=1.055 $Y2=0.36
.ends

