* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 a_113_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND A2 a_113_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_113_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_457_367# A2 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VGND A3 a_113_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_113_47# B1 a_1166_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND A2 a_113_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_113_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VGND A1 a_113_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_113_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR A1 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_113_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_1166_65# C1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 Y C1 a_1166_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VGND A3 a_113_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_30_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 Y A3 a_457_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_30_367# A2 a_457_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_30_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 Y A3 a_457_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_1166_65# B1 a_113_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 a_1166_65# C1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_457_367# A2 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_457_367# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 VPWR A1 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 a_30_367# A2 a_457_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 a_457_367# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 Y C1 a_1166_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 a_113_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X37 a_1166_65# B1 a_113_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 VGND A1 a_113_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 a_113_47# B1 a_1166_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
