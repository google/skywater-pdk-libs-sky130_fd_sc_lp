* File: sky130_fd_sc_lp__nor4b_1.pex.spice
* Created: Fri Aug 28 10:58:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4B_1%D_N 3 7 9 10 11 15
r29 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.51 $X2=0.43 $Y2=1.51
r30 11 15 6.53624 $w=3.33e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.592
+ $X2=0.43 $Y2=1.592
r31 9 14 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.665 $Y=1.51
+ $X2=0.43 $Y2=1.51
r32 9 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.665 $Y=1.51
+ $X2=0.74 $Y2=1.51
r33 5 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.74 $Y=1.675
+ $X2=0.74 $Y2=1.51
r34 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.74 $Y=1.675 $X2=0.74
+ $Y2=2.045
r35 1 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.74 $Y=1.345
+ $X2=0.74 $Y2=1.51
r36 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.74 $Y=1.345 $X2=0.74
+ $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_1%A 3 6 8 9 13 15
c38 8 0 1.59179e-19 $X=1.2 $Y=1.295
r39 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.35
+ $X2=1.19 $Y2=1.515
r40 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.35
+ $X2=1.19 $Y2=1.185
r41 8 9 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.665
r42 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=1.35 $X2=1.19 $Y2=1.35
r43 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.28 $Y=2.465
+ $X2=1.28 $Y2=1.515
r44 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.28 $Y=0.655
+ $X2=1.28 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_1%B 3 7 8 11 12 13
c38 13 0 1.89639e-19 $X=1.73 $Y=1.185
c39 12 0 5.79604e-20 $X=1.73 $Y=1.42
r40 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.42
+ $X2=1.73 $Y2=1.585
r41 11 13 58.4518 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.73 $Y=1.42
+ $X2=1.73 $Y2=1.185
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.42 $X2=1.73 $Y2=1.42
r43 8 12 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.73 $Y=1.665
+ $X2=1.73 $Y2=1.42
r44 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.755 $Y=0.655
+ $X2=1.755 $Y2=1.185
r45 3 14 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.64 $Y=2.465
+ $X2=1.64 $Y2=1.585
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_1%C 3 6 8 11 12 14
c40 6 0 5.79604e-20 $X=2.29 $Y=0.655
r41 11 14 54.9546 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.27 $Y=1.51
+ $X2=2.27 $Y2=1.725
r42 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.51
+ $X2=2.27 $Y2=1.345
r43 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.27
+ $Y=1.51 $X2=2.27 $Y2=1.51
r44 8 12 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.21 $Y=1.665
+ $X2=2.21 $Y2=1.51
r45 6 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.29 $Y=0.655
+ $X2=2.29 $Y2=1.345
r46 3 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.18 $Y=2.465
+ $X2=2.18 $Y2=1.725
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_1%A_80_131# 1 2 9 13 17 19 24 25 28 31 33 37
+ 38
r82 38 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.51
+ $X2=2.81 $Y2=1.675
r83 38 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.51
+ $X2=2.81 $Y2=1.345
r84 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=1.51 $X2=2.81 $Y2=1.51
r85 34 37 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.61 $Y=1.51 $X2=2.81
+ $Y2=1.51
r86 27 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=1.675
+ $X2=2.61 $Y2=1.51
r87 27 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.61 $Y=1.675
+ $X2=2.61 $Y2=1.97
r88 26 33 4.70473 $w=1.9e-07 $l=9.44722e-08 $layer=LI1_cond $X=0.935 $Y=2.055
+ $X2=0.85 $Y2=2.035
r89 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.525 $Y=2.055
+ $X2=2.61 $Y2=1.97
r90 25 26 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=2.525 $Y=2.055
+ $X2=0.935 $Y2=2.055
r91 24 33 1.74598 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.85 $Y=1.93
+ $X2=0.85 $Y2=2.035
r92 23 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=1.255
+ $X2=0.85 $Y2=1.17
r93 23 24 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.85 $Y=1.255
+ $X2=0.85 $Y2=1.93
r94 19 33 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.035
+ $X2=0.85 $Y2=2.035
r95 19 21 12.6753 $w=2.08e-07 $l=2.4e-07 $layer=LI1_cond $X=0.765 $Y=2.035
+ $X2=0.525 $Y2=2.035
r96 15 31 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.49 $Y=1.17
+ $X2=0.85 $Y2=1.17
r97 15 17 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.49 $Y=1.085
+ $X2=0.49 $Y2=0.865
r98 13 42 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.72 $Y=2.465
+ $X2=2.72 $Y2=1.675
r99 9 41 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.72 $Y=0.655
+ $X2=2.72 $Y2=1.345
r100 2 21 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.4
+ $Y=1.835 $X2=0.525 $Y2=2.035
r101 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.4
+ $Y=0.655 $X2=0.525 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_1%VPWR 1 6 8 10 17 18 21
r28 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r29 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r30 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=3.33
+ $X2=1.065 $Y2=3.33
r31 15 17 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=1.23 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=1.065 $Y2=3.33
r35 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=0.72
+ $Y2=3.33
r36 8 18 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 8 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=3.245
+ $X2=1.065 $Y2=3.33
r39 4 6 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=1.065 $Y=3.245
+ $X2=1.065 $Y2=2.425
r40 1 6 300 $w=1.7e-07 $l=7.03989e-07 $layer=licon1_PDIFF $count=2 $X=0.815
+ $Y=1.835 $X2=1.065 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_1%Y 1 2 3 12 14 15 18 20 24 25 26 27 42 46
c54 24 0 3.04599e-20 $X=2.477 $Y=1.075
r55 44 46 0.702709 $w=4.08e-07 $l=2.5e-08 $layer=LI1_cond $X=3.07 $Y=2.01
+ $X2=3.07 $Y2=2.035
r56 32 46 0.421625 $w=4.08e-07 $l=1.5e-08 $layer=LI1_cond $X=3.07 $Y=2.05
+ $X2=3.07 $Y2=2.035
r57 27 39 3.79463 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=3.07 $Y=2.775
+ $X2=3.07 $Y2=2.91
r58 26 27 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=3.07 $Y=2.405
+ $X2=3.07 $Y2=2.775
r59 25 44 0.281084 $w=4.08e-07 $l=1e-08 $layer=LI1_cond $X=3.07 $Y=2 $X2=3.07
+ $Y2=2.01
r60 25 42 7.09111 $w=4.08e-07 $l=1.55e-07 $layer=LI1_cond $X=3.07 $Y=2 $X2=3.07
+ $Y2=1.845
r61 25 26 8.99468 $w=4.08e-07 $l=3.2e-07 $layer=LI1_cond $X=3.07 $Y=2.085
+ $X2=3.07 $Y2=2.405
r62 25 32 0.983793 $w=4.08e-07 $l=3.5e-08 $layer=LI1_cond $X=3.07 $Y=2.085
+ $X2=3.07 $Y2=2.05
r63 22 42 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=3.17 $Y=1.165
+ $X2=3.17 $Y2=1.845
r64 21 24 6.76825 $w=1.75e-07 $l=1.23e-07 $layer=LI1_cond $X=2.6 $Y=1.075
+ $X2=2.477 $Y2=1.075
r65 20 22 6.86909 $w=1.8e-07 $l=1.43091e-07 $layer=LI1_cond $X=3.065 $Y=1.075
+ $X2=3.17 $Y2=1.165
r66 20 21 28.6515 $w=1.78e-07 $l=4.65e-07 $layer=LI1_cond $X=3.065 $Y=1.075
+ $X2=2.6 $Y2=1.075
r67 16 24 0.164012 $w=2.45e-07 $l=9e-08 $layer=LI1_cond $X=2.477 $Y=0.985
+ $X2=2.477 $Y2=1.075
r68 16 18 26.5767 $w=2.43e-07 $l=5.65e-07 $layer=LI1_cond $X=2.477 $Y=0.985
+ $X2=2.477 $Y2=0.42
r69 14 24 6.76825 $w=1.75e-07 $l=1.24475e-07 $layer=LI1_cond $X=2.355 $Y=1.08
+ $X2=2.477 $Y2=1.075
r70 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.355 $Y=1.08
+ $X2=1.685 $Y2=1.08
r71 10 15 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.57 $Y=0.995
+ $X2=1.685 $Y2=1.08
r72 10 12 28.8111 $w=2.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.57 $Y=0.995
+ $X2=1.57 $Y2=0.42
r73 3 44 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=1.835 $X2=2.97 $Y2=2.01
r74 3 39 400 $w=1.7e-07 $l=1.1592e-06 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=1.835 $X2=2.97 $Y2=2.91
r75 2 18 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.365
+ $Y=0.235 $X2=2.505 $Y2=0.42
r76 1 12 91 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=2 $X=1.355
+ $Y=0.235 $X2=1.54 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_1%VGND 1 2 3 12 18 20 22 25 26 28 29 30 39 45
r43 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r44 42 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r45 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 39 44 4.4922 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.77 $Y=0 $X2=3.065
+ $Y2=0
r47 39 41 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.77 $Y=0 $X2=2.64
+ $Y2=0
r48 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r49 30 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 30 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r51 30 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 28 37 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.68
+ $Y2=0
r53 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.02
+ $Y2=0
r54 27 41 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.64
+ $Y2=0
r55 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.02
+ $Y2=0
r56 25 33 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.72
+ $Y2=0
r57 25 26 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=1.015
+ $Y2=0
r58 24 37 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.68
+ $Y2=0
r59 24 26 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.015
+ $Y2=0
r60 20 44 3.27398 $w=3.3e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.935 $Y=0.085
+ $X2=3.065 $Y2=0
r61 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=0.085
+ $X2=2.935 $Y2=0.38
r62 16 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r63 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.38
r64 12 14 11.8279 $w=4.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.015 $Y=0.38
+ $X2=1.015 $Y2=0.825
r65 10 26 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.085
+ $X2=1.015 $Y2=0
r66 10 12 7.84096 $w=4.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=0.085
+ $X2=1.015 $Y2=0.38
r67 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.795
+ $Y=0.235 $X2=2.935 $Y2=0.38
r68 2 18 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=1.83
+ $Y=0.235 $X2=2.02 $Y2=0.38
r69 1 14 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=0.815
+ $Y=0.655 $X2=0.955 $Y2=0.825
r70 1 12 182 $w=1.7e-07 $l=3.79967e-07 $layer=licon1_NDIFF $count=1 $X=0.815
+ $Y=0.655 $X2=1.065 $Y2=0.38
.ends

