* File: sky130_fd_sc_lp__nor3b_lp.pxi.spice
* Created: Wed Sep  2 10:09:56 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3B_LP%A N_A_c_70_n N_A_M1001_g N_A_c_71_n N_A_c_72_n
+ N_A_M1010_g N_A_c_73_n N_A_M1011_g N_A_c_74_n N_A_c_75_n A A N_A_c_77_n
+ N_A_c_78_n PM_SKY130_FD_SC_LP__NOR3B_LP%A
x_PM_SKY130_FD_SC_LP__NOR3B_LP%B N_B_M1003_g N_B_c_113_n N_B_M1002_g N_B_c_114_n
+ N_B_c_115_n N_B_M1004_g N_B_c_116_n N_B_c_117_n N_B_c_123_n N_B_c_118_n B B B
+ B B N_B_c_120_n PM_SKY130_FD_SC_LP__NOR3B_LP%B
x_PM_SKY130_FD_SC_LP__NOR3B_LP%A_350_269# N_A_350_269#_M1009_d
+ N_A_350_269#_M1006_d N_A_350_269#_M1000_g N_A_350_269#_c_177_n
+ N_A_350_269#_M1007_g N_A_350_269#_c_178_n N_A_350_269#_M1005_g
+ N_A_350_269#_c_179_n N_A_350_269#_c_180_n N_A_350_269#_c_186_n
+ N_A_350_269#_c_187_n N_A_350_269#_c_181_n N_A_350_269#_c_182_n
+ N_A_350_269#_c_183_n N_A_350_269#_c_184_n
+ PM_SKY130_FD_SC_LP__NOR3B_LP%A_350_269#
x_PM_SKY130_FD_SC_LP__NOR3B_LP%C_N N_C_N_M1008_g N_C_N_M1006_g N_C_N_M1009_g C_N
+ C_N N_C_N_c_246_n PM_SKY130_FD_SC_LP__NOR3B_LP%C_N
x_PM_SKY130_FD_SC_LP__NOR3B_LP%VPWR N_VPWR_M1010_s N_VPWR_M1006_s N_VPWR_c_278_n
+ N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n
+ VPWR N_VPWR_c_284_n N_VPWR_c_277_n PM_SKY130_FD_SC_LP__NOR3B_LP%VPWR
x_PM_SKY130_FD_SC_LP__NOR3B_LP%Y N_Y_M1001_s N_Y_M1004_d N_Y_M1000_d N_Y_c_312_n
+ N_Y_c_313_n N_Y_c_317_n N_Y_c_318_n N_Y_c_314_n N_Y_c_315_n Y
+ PM_SKY130_FD_SC_LP__NOR3B_LP%Y
x_PM_SKY130_FD_SC_LP__NOR3B_LP%VGND N_VGND_M1011_d N_VGND_M1005_d N_VGND_c_371_n
+ N_VGND_c_372_n VGND N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n
+ N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n PM_SKY130_FD_SC_LP__NOR3B_LP%VGND
cc_1 VNB N_A_c_70_n 0.0171842f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.78
cc_2 VNB N_A_c_71_n 0.023214f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.64
cc_3 VNB N_A_c_72_n 0.0147293f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=0.855
cc_4 VNB N_A_c_73_n 0.013881f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.78
cc_5 VNB N_A_c_74_n 0.00667205f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.855
cc_6 VNB N_A_c_75_n 0.00134965f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.845
cc_7 VNB A 0.0273716f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_A_c_77_n 0.0225549f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.34
cc_9 VNB N_A_c_78_n 0.0170168f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.175
cc_10 VNB N_B_c_113_n 0.0138865f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.175
cc_11 VNB N_B_c_114_n 0.0173512f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.845
cc_12 VNB N_B_c_115_n 0.0137713f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=2.545
cc_13 VNB N_B_c_116_n 0.0200912f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.495
cc_14 VNB N_B_c_117_n 0.01799f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.855
cc_15 VNB N_B_c_118_n 0.00466383f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB B 0.00866304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_c_120_n 0.015832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_350_269#_M1000_g 0.0106128f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.855
cc_19 VNB N_A_350_269#_c_177_n 0.0157362f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=2.545
cc_20 VNB N_A_350_269#_c_178_n 0.0161154f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.78
cc_21 VNB N_A_350_269#_c_179_n 0.0166304f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_A_350_269#_c_180_n 0.0240181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_350_269#_c_181_n 0.0142454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_350_269#_c_182_n 0.0999297f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.51
cc_25 VNB N_A_350_269#_c_183_n 0.0132078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_350_269#_c_184_n 0.0314522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C_N_M1008_g 0.0311565f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.495
cc_28 VNB N_C_N_M1009_g 0.0400902f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=2.545
cc_29 VNB C_N 2.87194e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_N_c_246_n 0.053128f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.845
cc_31 VNB N_VPWR_c_277_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_312_n 0.0130915f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.845
cc_33 VNB N_Y_c_313_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.78
cc_34 VNB N_Y_c_314_n 0.00224806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_315_n 0.00905013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB Y 0.0425197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_371_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.855
cc_38 VNB N_VGND_c_372_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_373_n 0.027925f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.855
cc_40 VNB N_VGND_c_374_n 0.0351604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_375_n 0.0275168f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.34
cc_42 VNB N_VGND_c_376_n 0.22915f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.175
cc_43 VNB N_VGND_c_377_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_378_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A_M1010_g 0.0354954f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=2.545
cc_46 VPB N_A_c_75_n 0.0212745f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.845
cc_47 VPB A 0.0212557f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_48 VPB N_B_M1003_g 0.0262177f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.495
cc_49 VPB N_B_c_117_n 0.00168838f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.855
cc_50 VPB N_B_c_123_n 0.0118896f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.845
cc_51 VPB B 0.00345404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_350_269#_M1000_g 0.0453489f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.855
cc_53 VPB N_A_350_269#_c_186_n 0.0118411f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.34
cc_54 VPB N_A_350_269#_c_187_n 0.035517f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.34
cc_55 VPB N_A_350_269#_c_184_n 0.0175873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_C_N_M1006_g 0.0407534f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.64
cc_57 VPB C_N 0.00242689f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_C_N_c_246_n 0.0325415f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.845
cc_59 VPB N_VPWR_c_278_n 0.0465298f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.855
cc_60 VPB N_VPWR_c_279_n 0.0248819f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=0.495
cc_61 VPB N_VPWR_c_280_n 0.0143948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_281_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_63 VPB N_VPWR_c_282_n 0.059657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_283_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_284_n 0.0192431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_277_n 0.0936149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_Y_c_317_n 0.00522059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_Y_c_318_n 0.016426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_Y_c_315_n 0.0126765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 N_A_M1010_g N_B_M1003_g 0.0264724f $X=0.815 $Y=2.545 $X2=0 $Y2=0
cc_71 N_A_c_73_n N_B_c_113_n 0.00957171f $X=0.965 $Y=0.78 $X2=0 $Y2=0
cc_72 N_A_c_78_n N_B_c_116_n 0.00153974f $X=0.735 $Y=1.175 $X2=0 $Y2=0
cc_73 N_A_c_71_n N_B_c_117_n 0.0264724f $X=0.735 $Y=1.64 $X2=0 $Y2=0
cc_74 N_A_c_75_n N_B_c_123_n 0.0264724f $X=0.735 $Y=1.845 $X2=0 $Y2=0
cc_75 N_A_c_72_n N_B_c_118_n 0.00957171f $X=0.89 $Y=0.855 $X2=0 $Y2=0
cc_76 A B 0.04783f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_77_n B 0.0188855f $X=0.695 $Y=1.34 $X2=0 $Y2=0
cc_78 A N_B_c_120_n 6.29825e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A_c_77_n N_B_c_120_n 0.0264724f $X=0.695 $Y=1.34 $X2=0 $Y2=0
cc_80 N_A_M1010_g N_VPWR_c_278_n 0.0242186f $X=0.815 $Y=2.545 $X2=0 $Y2=0
cc_81 N_A_c_75_n N_VPWR_c_278_n 0.00432933f $X=0.735 $Y=1.845 $X2=0 $Y2=0
cc_82 A N_VPWR_c_278_n 0.0283965f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A_M1010_g N_VPWR_c_282_n 0.00802402f $X=0.815 $Y=2.545 $X2=0 $Y2=0
cc_84 N_A_M1010_g N_VPWR_c_277_n 0.0142664f $X=0.815 $Y=2.545 $X2=0 $Y2=0
cc_85 N_A_c_72_n N_Y_c_312_n 0.00969118f $X=0.89 $Y=0.855 $X2=0 $Y2=0
cc_86 A N_Y_c_312_n 0.00186599f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A_c_77_n N_Y_c_312_n 0.00186276f $X=0.695 $Y=1.34 $X2=0 $Y2=0
cc_88 N_A_c_70_n Y 0.01433f $X=0.605 $Y=0.78 $X2=0 $Y2=0
cc_89 N_A_c_72_n Y 0.00431495f $X=0.89 $Y=0.855 $X2=0 $Y2=0
cc_90 N_A_c_73_n Y 0.00360399f $X=0.965 $Y=0.78 $X2=0 $Y2=0
cc_91 N_A_c_74_n Y 0.00535129f $X=0.605 $Y=0.855 $X2=0 $Y2=0
cc_92 A Y 0.0610875f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A_c_77_n Y 0.00110439f $X=0.695 $Y=1.34 $X2=0 $Y2=0
cc_94 N_A_c_78_n Y 0.00450674f $X=0.735 $Y=1.175 $X2=0 $Y2=0
cc_95 N_A_c_70_n N_VGND_c_371_n 0.00149712f $X=0.605 $Y=0.78 $X2=0 $Y2=0
cc_96 N_A_c_73_n N_VGND_c_371_n 0.00946538f $X=0.965 $Y=0.78 $X2=0 $Y2=0
cc_97 N_A_c_70_n N_VGND_c_373_n 0.00352123f $X=0.605 $Y=0.78 $X2=0 $Y2=0
cc_98 N_A_c_73_n N_VGND_c_373_n 0.00445056f $X=0.965 $Y=0.78 $X2=0 $Y2=0
cc_99 N_A_c_70_n N_VGND_c_376_n 0.005602f $X=0.605 $Y=0.78 $X2=0 $Y2=0
cc_100 N_A_c_73_n N_VGND_c_376_n 0.0041956f $X=0.965 $Y=0.78 $X2=0 $Y2=0
cc_101 N_B_M1003_g N_A_350_269#_M1000_g 0.0521984f $X=1.305 $Y=2.545 $X2=0 $Y2=0
cc_102 N_B_c_123_n N_A_350_269#_M1000_g 0.0138499f $X=1.345 $Y=1.85 $X2=0 $Y2=0
cc_103 B N_A_350_269#_M1000_g 0.0446403f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B_c_115_n N_A_350_269#_c_177_n 0.00898095f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_105 N_B_c_114_n N_A_350_269#_c_182_n 0.0111524f $X=1.68 $Y=0.855 $X2=0 $Y2=0
cc_106 N_B_c_116_n N_A_350_269#_c_182_n 0.00306982f $X=1.345 $Y=1.18 $X2=0 $Y2=0
cc_107 N_B_c_117_n N_A_350_269#_c_182_n 0.0138499f $X=1.345 $Y=1.685 $X2=0 $Y2=0
cc_108 B N_A_350_269#_c_182_n 0.00548186f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B_c_120_n N_A_350_269#_c_182_n 0.00226032f $X=1.345 $Y=1.345 $X2=0
+ $Y2=0
cc_110 N_B_M1003_g N_VPWR_c_278_n 0.00216731f $X=1.305 $Y=2.545 $X2=0 $Y2=0
cc_111 B N_VPWR_c_278_n 0.0393372f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B_M1003_g N_VPWR_c_282_n 0.00595064f $X=1.305 $Y=2.545 $X2=0 $Y2=0
cc_113 B N_VPWR_c_282_n 0.0194157f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B_M1003_g N_VPWR_c_277_n 0.00772137f $X=1.305 $Y=2.545 $X2=0 $Y2=0
cc_115 B N_VPWR_c_277_n 0.0232206f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_116 B A_188_409# 0.0106484f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_117 B A_286_409# 0.00286113f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_118 N_B_c_114_n N_Y_c_312_n 0.0151974f $X=1.68 $Y=0.855 $X2=0 $Y2=0
cc_119 N_B_c_116_n N_Y_c_312_n 0.00579982f $X=1.345 $Y=1.18 $X2=0 $Y2=0
cc_120 N_B_c_118_n N_Y_c_312_n 0.00594488f $X=1.395 $Y=0.855 $X2=0 $Y2=0
cc_121 B N_Y_c_312_n 0.0542287f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B_c_120_n N_Y_c_312_n 0.00108014f $X=1.345 $Y=1.345 $X2=0 $Y2=0
cc_123 N_B_c_113_n N_Y_c_313_n 0.00170583f $X=1.395 $Y=0.78 $X2=0 $Y2=0
cc_124 N_B_c_114_n N_Y_c_313_n 0.00260361f $X=1.68 $Y=0.855 $X2=0 $Y2=0
cc_125 N_B_c_115_n N_Y_c_313_n 0.0100197f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_126 N_B_M1003_g N_Y_c_318_n 7.47128e-19 $X=1.305 $Y=2.545 $X2=0 $Y2=0
cc_127 N_B_c_114_n N_Y_c_314_n 0.00169138f $X=1.68 $Y=0.855 $X2=0 $Y2=0
cc_128 N_B_M1003_g N_Y_c_315_n 5.89775e-19 $X=1.305 $Y=2.545 $X2=0 $Y2=0
cc_129 N_B_c_116_n N_Y_c_315_n 0.00293654f $X=1.345 $Y=1.18 $X2=0 $Y2=0
cc_130 N_B_c_117_n N_Y_c_315_n 2.97019e-19 $X=1.345 $Y=1.685 $X2=0 $Y2=0
cc_131 B N_Y_c_315_n 0.128502f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B_c_120_n N_Y_c_315_n 3.43325e-19 $X=1.345 $Y=1.345 $X2=0 $Y2=0
cc_133 N_B_c_118_n Y 2.15578e-19 $X=1.395 $Y=0.855 $X2=0 $Y2=0
cc_134 N_B_c_113_n N_VGND_c_371_n 0.0106455f $X=1.395 $Y=0.78 $X2=0 $Y2=0
cc_135 N_B_c_115_n N_VGND_c_371_n 0.00189426f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_136 N_B_c_113_n N_VGND_c_374_n 0.00445056f $X=1.395 $Y=0.78 $X2=0 $Y2=0
cc_137 N_B_c_114_n N_VGND_c_374_n 4.57848e-19 $X=1.68 $Y=0.855 $X2=0 $Y2=0
cc_138 N_B_c_115_n N_VGND_c_374_n 0.00502664f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_139 N_B_c_113_n N_VGND_c_376_n 0.0041956f $X=1.395 $Y=0.78 $X2=0 $Y2=0
cc_140 N_B_c_114_n N_VGND_c_376_n 6.33118e-19 $X=1.68 $Y=0.855 $X2=0 $Y2=0
cc_141 N_B_c_115_n N_VGND_c_376_n 0.00563733f $X=1.755 $Y=0.78 $X2=0 $Y2=0
cc_142 N_A_350_269#_c_178_n N_C_N_M1008_g 0.0147173f $X=2.545 $Y=0.825 $X2=0
+ $Y2=0
cc_143 N_A_350_269#_c_179_n N_C_N_M1008_g 0.0111491f $X=3.385 $Y=0.91 $X2=0
+ $Y2=0
cc_144 N_A_350_269#_c_180_n N_C_N_M1008_g 0.00193397f $X=3.55 $Y=0.495 $X2=0
+ $Y2=0
cc_145 N_A_350_269#_c_181_n N_C_N_M1008_g 0.00244844f $X=2.49 $Y=0.99 $X2=0
+ $Y2=0
cc_146 N_A_350_269#_c_182_n N_C_N_M1008_g 0.0369189f $X=2.49 $Y=0.99 $X2=0 $Y2=0
cc_147 N_A_350_269#_c_186_n N_C_N_M1006_g 0.00451956f $X=3.55 $Y=2.19 $X2=0
+ $Y2=0
cc_148 N_A_350_269#_c_187_n N_C_N_M1006_g 0.015872f $X=3.55 $Y=2.9 $X2=0 $Y2=0
cc_149 N_A_350_269#_c_179_n N_C_N_M1009_g 0.0118348f $X=3.385 $Y=0.91 $X2=0
+ $Y2=0
cc_150 N_A_350_269#_c_180_n N_C_N_M1009_g 0.01276f $X=3.55 $Y=0.495 $X2=0 $Y2=0
cc_151 N_A_350_269#_c_183_n N_C_N_M1009_g 0.00513266f $X=3.55 $Y=0.91 $X2=0
+ $Y2=0
cc_152 N_A_350_269#_c_184_n N_C_N_M1009_g 0.0277429f $X=3.55 $Y=2.025 $X2=0
+ $Y2=0
cc_153 N_A_350_269#_c_179_n C_N 0.0245266f $X=3.385 $Y=0.91 $X2=0 $Y2=0
cc_154 N_A_350_269#_c_181_n C_N 0.0176462f $X=2.49 $Y=0.99 $X2=0 $Y2=0
cc_155 N_A_350_269#_c_182_n C_N 0.00132975f $X=2.49 $Y=0.99 $X2=0 $Y2=0
cc_156 N_A_350_269#_c_184_n C_N 0.0321436f $X=3.55 $Y=2.025 $X2=0 $Y2=0
cc_157 N_A_350_269#_c_179_n N_C_N_c_246_n 2.06304e-19 $X=3.385 $Y=0.91 $X2=0
+ $Y2=0
cc_158 N_A_350_269#_c_186_n N_VPWR_c_279_n 0.0684934f $X=3.55 $Y=2.19 $X2=0
+ $Y2=0
cc_159 N_A_350_269#_M1000_g N_VPWR_c_282_n 0.00807509f $X=1.875 $Y=2.545 $X2=0
+ $Y2=0
cc_160 N_A_350_269#_c_187_n N_VPWR_c_284_n 0.0220321f $X=3.55 $Y=2.9 $X2=0 $Y2=0
cc_161 N_A_350_269#_M1000_g N_VPWR_c_277_n 0.0151816f $X=1.875 $Y=2.545 $X2=0
+ $Y2=0
cc_162 N_A_350_269#_c_187_n N_VPWR_c_277_n 0.0125808f $X=3.55 $Y=2.9 $X2=0 $Y2=0
cc_163 N_A_350_269#_c_182_n N_Y_c_312_n 3.01841e-19 $X=2.49 $Y=0.99 $X2=0 $Y2=0
cc_164 N_A_350_269#_c_177_n N_Y_c_313_n 0.0117349f $X=2.185 $Y=0.825 $X2=0 $Y2=0
cc_165 N_A_350_269#_c_178_n N_Y_c_313_n 0.00196674f $X=2.545 $Y=0.825 $X2=0
+ $Y2=0
cc_166 N_A_350_269#_M1000_g N_Y_c_317_n 0.00303908f $X=1.875 $Y=2.545 $X2=0
+ $Y2=0
cc_167 N_A_350_269#_c_182_n N_Y_c_317_n 0.00527997f $X=2.49 $Y=0.99 $X2=0 $Y2=0
cc_168 N_A_350_269#_M1000_g N_Y_c_318_n 0.0154719f $X=1.875 $Y=2.545 $X2=0 $Y2=0
cc_169 N_A_350_269#_c_181_n N_Y_c_314_n 0.0137383f $X=2.49 $Y=0.99 $X2=0 $Y2=0
cc_170 N_A_350_269#_c_182_n N_Y_c_314_n 0.0120765f $X=2.49 $Y=0.99 $X2=0 $Y2=0
cc_171 N_A_350_269#_M1000_g N_Y_c_315_n 0.0173651f $X=1.875 $Y=2.545 $X2=0 $Y2=0
cc_172 N_A_350_269#_c_181_n N_Y_c_315_n 0.0340384f $X=2.49 $Y=0.99 $X2=0 $Y2=0
cc_173 N_A_350_269#_c_182_n N_Y_c_315_n 0.02374f $X=2.49 $Y=0.99 $X2=0 $Y2=0
cc_174 N_A_350_269#_c_177_n N_VGND_c_372_n 0.00188833f $X=2.185 $Y=0.825 $X2=0
+ $Y2=0
cc_175 N_A_350_269#_c_178_n N_VGND_c_372_n 0.0105779f $X=2.545 $Y=0.825 $X2=0
+ $Y2=0
cc_176 N_A_350_269#_c_179_n N_VGND_c_372_n 0.0171154f $X=3.385 $Y=0.91 $X2=0
+ $Y2=0
cc_177 N_A_350_269#_c_180_n N_VGND_c_372_n 0.0127138f $X=3.55 $Y=0.495 $X2=0
+ $Y2=0
cc_178 N_A_350_269#_c_181_n N_VGND_c_372_n 0.00316485f $X=2.49 $Y=0.99 $X2=0
+ $Y2=0
cc_179 N_A_350_269#_c_177_n N_VGND_c_374_n 0.00488765f $X=2.185 $Y=0.825 $X2=0
+ $Y2=0
cc_180 N_A_350_269#_c_178_n N_VGND_c_374_n 0.00445056f $X=2.545 $Y=0.825 $X2=0
+ $Y2=0
cc_181 N_A_350_269#_c_180_n N_VGND_c_375_n 0.0220321f $X=3.55 $Y=0.495 $X2=0
+ $Y2=0
cc_182 N_A_350_269#_c_177_n N_VGND_c_376_n 0.00905024f $X=2.185 $Y=0.825 $X2=0
+ $Y2=0
cc_183 N_A_350_269#_c_178_n N_VGND_c_376_n 0.0041935f $X=2.545 $Y=0.825 $X2=0
+ $Y2=0
cc_184 N_A_350_269#_c_179_n N_VGND_c_376_n 0.0152176f $X=3.385 $Y=0.91 $X2=0
+ $Y2=0
cc_185 N_A_350_269#_c_180_n N_VGND_c_376_n 0.0125808f $X=3.55 $Y=0.495 $X2=0
+ $Y2=0
cc_186 N_A_350_269#_c_181_n N_VGND_c_376_n 0.00947285f $X=2.49 $Y=0.99 $X2=0
+ $Y2=0
cc_187 N_C_N_M1006_g N_VPWR_c_279_n 0.0249766f $X=3.285 $Y=2.545 $X2=0 $Y2=0
cc_188 C_N N_VPWR_c_279_n 0.0235964f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_189 N_C_N_c_246_n N_VPWR_c_279_n 0.00225955f $X=3.07 $Y=1.34 $X2=0 $Y2=0
cc_190 N_C_N_M1006_g N_VPWR_c_284_n 0.00769046f $X=3.285 $Y=2.545 $X2=0 $Y2=0
cc_191 N_C_N_M1006_g N_VPWR_c_277_n 0.0140911f $X=3.285 $Y=2.545 $X2=0 $Y2=0
cc_192 N_C_N_M1008_g N_VGND_c_372_n 0.0106455f $X=2.975 $Y=0.495 $X2=0 $Y2=0
cc_193 N_C_N_M1009_g N_VGND_c_372_n 0.00189426f $X=3.335 $Y=0.495 $X2=0 $Y2=0
cc_194 N_C_N_M1008_g N_VGND_c_375_n 0.00445056f $X=2.975 $Y=0.495 $X2=0 $Y2=0
cc_195 N_C_N_M1009_g N_VGND_c_375_n 0.00502664f $X=3.335 $Y=0.495 $X2=0 $Y2=0
cc_196 N_C_N_M1008_g N_VGND_c_376_n 0.0041956f $X=2.975 $Y=0.495 $X2=0 $Y2=0
cc_197 N_C_N_M1009_g N_VGND_c_376_n 0.00628426f $X=3.335 $Y=0.495 $X2=0 $Y2=0
cc_198 N_VPWR_c_279_n N_Y_c_317_n 0.038352f $X=3.02 $Y=2.19 $X2=0 $Y2=0
cc_199 N_VPWR_c_282_n N_Y_c_318_n 0.0220321f $X=2.855 $Y=3.33 $X2=0 $Y2=0
cc_200 N_VPWR_c_277_n N_Y_c_318_n 0.0125808f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_201 Y A_136_57# 0.00132459f $X=0.155 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_202 N_Y_c_312_n N_VGND_c_371_n 0.0200008f $X=1.805 $Y=0.91 $X2=0 $Y2=0
cc_203 N_Y_c_313_n N_VGND_c_371_n 0.0127429f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_204 Y N_VGND_c_371_n 0.00598935f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_205 N_Y_c_313_n N_VGND_c_372_n 0.0129849f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_206 Y N_VGND_c_373_n 0.0366057f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_207 N_Y_c_313_n N_VGND_c_374_n 0.0225886f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_208 N_Y_c_312_n N_VGND_c_376_n 0.0198925f $X=1.805 $Y=0.91 $X2=0 $Y2=0
cc_209 N_Y_c_313_n N_VGND_c_376_n 0.0128111f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_210 Y N_VGND_c_376_n 0.0255735f $X=0.155 $Y=0.47 $X2=0 $Y2=0
