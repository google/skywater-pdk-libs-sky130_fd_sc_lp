* File: sky130_fd_sc_lp__and4bb_m.pxi.spice
* Created: Fri Aug 28 10:09:42 2020
* 
x_PM_SKY130_FD_SC_LP__AND4BB_M%A_N N_A_N_M1000_g N_A_N_M1010_g N_A_N_c_94_n
+ N_A_N_c_95_n N_A_N_c_96_n A_N A_N N_A_N_c_98_n
+ PM_SKY130_FD_SC_LP__AND4BB_M%A_N
x_PM_SKY130_FD_SC_LP__AND4BB_M%B_N N_B_N_M1001_g N_B_N_M1012_g N_B_N_c_128_n
+ N_B_N_c_129_n N_B_N_c_130_n B_N B_N N_B_N_c_132_n
+ PM_SKY130_FD_SC_LP__AND4BB_M%B_N
x_PM_SKY130_FD_SC_LP__AND4BB_M%A_54_55# N_A_54_55#_M1000_s N_A_54_55#_M1010_s
+ N_A_54_55#_M1008_g N_A_54_55#_c_167_n N_A_54_55#_M1004_g N_A_54_55#_c_168_n
+ N_A_54_55#_c_174_n N_A_54_55#_c_175_n N_A_54_55#_c_176_n N_A_54_55#_c_169_n
+ N_A_54_55#_c_177_n N_A_54_55#_c_178_n N_A_54_55#_c_170_n N_A_54_55#_c_171_n
+ N_A_54_55#_c_172_n N_A_54_55#_c_173_n PM_SKY130_FD_SC_LP__AND4BB_M%A_54_55#
x_PM_SKY130_FD_SC_LP__AND4BB_M%A_223_55# N_A_223_55#_M1001_d N_A_223_55#_M1012_d
+ N_A_223_55#_M1003_g N_A_223_55#_M1013_g N_A_223_55#_c_247_n
+ N_A_223_55#_c_248_n N_A_223_55#_c_242_n N_A_223_55#_c_243_n
+ N_A_223_55#_c_249_n N_A_223_55#_c_267_n N_A_223_55#_c_244_n
+ N_A_223_55#_c_245_n N_A_223_55#_c_274_n PM_SKY130_FD_SC_LP__AND4BB_M%A_223_55#
x_PM_SKY130_FD_SC_LP__AND4BB_M%C N_C_M1011_g N_C_M1006_g C C N_C_c_315_n
+ N_C_c_316_n N_C_c_317_n PM_SKY130_FD_SC_LP__AND4BB_M%C
x_PM_SKY130_FD_SC_LP__AND4BB_M%D N_D_M1007_g N_D_M1002_g D N_D_c_365_n
+ PM_SKY130_FD_SC_LP__AND4BB_M%D
x_PM_SKY130_FD_SC_LP__AND4BB_M%A_332_125# N_A_332_125#_M1004_s
+ N_A_332_125#_M1008_d N_A_332_125#_M1011_d N_A_332_125#_c_411_n
+ N_A_332_125#_M1005_g N_A_332_125#_M1009_g N_A_332_125#_c_413_n
+ N_A_332_125#_c_424_n N_A_332_125#_c_414_n N_A_332_125#_c_415_n
+ N_A_332_125#_c_416_n N_A_332_125#_c_417_n N_A_332_125#_c_406_n
+ N_A_332_125#_c_446_n N_A_332_125#_c_419_n N_A_332_125#_c_420_n
+ N_A_332_125#_c_407_n N_A_332_125#_c_408_n N_A_332_125#_c_482_n
+ N_A_332_125#_c_409_n N_A_332_125#_c_410_n
+ PM_SKY130_FD_SC_LP__AND4BB_M%A_332_125#
x_PM_SKY130_FD_SC_LP__AND4BB_M%VPWR N_VPWR_M1010_d N_VPWR_M1008_s N_VPWR_M1003_d
+ N_VPWR_M1007_d N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n
+ N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n
+ N_VPWR_c_532_n VPWR N_VPWR_c_533_n N_VPWR_c_522_n N_VPWR_c_535_n
+ PM_SKY130_FD_SC_LP__AND4BB_M%VPWR
x_PM_SKY130_FD_SC_LP__AND4BB_M%X N_X_M1009_d N_X_M1005_d N_X_c_573_n X X X X
+ PM_SKY130_FD_SC_LP__AND4BB_M%X
x_PM_SKY130_FD_SC_LP__AND4BB_M%VGND N_VGND_M1000_d N_VGND_M1002_d N_VGND_c_588_n
+ N_VGND_c_589_n VGND N_VGND_c_590_n N_VGND_c_591_n N_VGND_c_592_n
+ N_VGND_c_593_n N_VGND_c_594_n PM_SKY130_FD_SC_LP__AND4BB_M%VGND
cc_1 VNB N_A_N_M1010_g 0.0104537f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.195
cc_2 VNB N_A_N_c_94_n 0.0202581f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.805
cc_3 VNB N_A_N_c_95_n 0.0236573f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.31
cc_4 VNB N_A_N_c_96_n 0.0164899f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.475
cc_5 VNB A_N 0.00857592f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_A_N_c_98_n 0.0164912f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.97
cc_7 VNB N_B_N_M1012_g 0.0105631f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.195
cc_8 VNB N_B_N_c_128_n 0.0206692f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.805
cc_9 VNB N_B_N_c_129_n 0.0261581f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.31
cc_10 VNB N_B_N_c_130_n 0.0167786f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.475
cc_11 VNB B_N 0.00359178f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_12 VNB N_B_N_c_132_n 0.0187731f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.97
cc_13 VNB N_A_54_55#_c_167_n 0.0190697f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_14 VNB N_A_54_55#_c_168_n 0.0370505f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.97
cc_15 VNB N_A_54_55#_c_169_n 0.0489707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_54_55#_c_170_n 0.00359747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_54_55#_c_171_n 0.0274159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_54_55#_c_172_n 0.0157146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_54_55#_c_173_n 0.00510731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_223_55#_M1013_g 0.0299576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_223_55#_c_242_n 0.0338096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_223_55#_c_243_n 0.049737f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.97
cc_23 VNB N_A_223_55#_c_244_n 0.0129429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_223_55#_c_245_n 0.00168036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C_M1011_g 0.00892365f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.485
cc_26 VNB N_C_c_315_n 0.0292245f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_27 VNB N_C_c_316_n 0.0151807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C_c_317_n 0.0177382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_D_M1002_g 0.0429735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_332_125#_M1009_g 0.0457411f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.97
cc_31 VNB N_A_332_125#_c_406_n 0.00352653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_332_125#_c_407_n 0.00467597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_332_125#_c_408_n 0.00651897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_332_125#_c_409_n 0.00377759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_332_125#_c_410_n 0.0121826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_522_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB X 0.0405401f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_38 VNB N_VGND_c_588_n 0.00603613f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.475
cc_39 VNB N_VGND_c_589_n 0.0273835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_590_n 0.0652968f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.925
cc_41 VNB N_VGND_c_591_n 0.0202355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_592_n 0.27046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_593_n 0.0258079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_594_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A_N_M1010_g 0.0357248f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.195
cc_46 VPB N_B_N_M1012_g 0.0328871f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.195
cc_47 VPB N_A_54_55#_c_174_n 0.0166433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_54_55#_c_175_n 0.0354032f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.97
cc_49 VPB N_A_54_55#_c_176_n 0.0377905f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.295
cc_50 VPB N_A_54_55#_c_177_n 0.0281918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_54_55#_c_178_n 0.0281602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_54_55#_c_173_n 0.0134772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_223_55#_M1003_g 0.0346759f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=0.805
cc_54 VPB N_A_223_55#_c_247_n 0.0230851f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=0.97
cc_55 VPB N_A_223_55#_c_248_n 0.014625f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=0.97
cc_56 VPB N_A_223_55#_c_249_n 0.0240066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_223_55#_c_244_n 0.00312871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_C_M1011_g 0.0577162f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.485
cc_59 VPB N_D_M1007_g 0.0368983f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.485
cc_60 VPB N_D_M1002_g 0.0106064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB D 0.00229918f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=0.805
cc_62 VPB N_D_c_365_n 0.0314523f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_63 VPB N_A_332_125#_c_411_n 0.023491f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.475
cc_64 VPB N_A_332_125#_M1005_g 0.0385842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_332_125#_c_413_n 0.0218957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_332_125#_c_414_n 0.00136805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_332_125#_c_415_n 0.0112322f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_332_125#_c_416_n 0.0042372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_332_125#_c_417_n 0.0063613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_332_125#_c_406_n 0.00717241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_332_125#_c_419_n 0.00984692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_332_125#_c_420_n 0.00195925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_332_125#_c_408_n 0.00721425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_332_125#_c_409_n 0.00227797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_332_125#_c_410_n 0.00869902f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_523_n 0.0447948f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=0.97
cc_77 VPB N_VPWR_c_524_n 0.00381618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_525_n 0.00380657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_526_n 4.12476e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_527_n 0.0193478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_528_n 0.00401177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_529_n 0.0181538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_530_n 0.00401177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_531_n 0.0158304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_532_n 0.00436274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_533_n 0.0221696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_522_n 0.091729f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_535_n 0.0290685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_X_c_573_n 0.0220189f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.31
cc_90 VPB X 0.0500603f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_91 N_A_N_M1010_g N_B_N_M1012_g 0.031561f $X=0.61 $Y=2.195 $X2=0 $Y2=0
cc_92 N_A_N_c_94_n N_B_N_c_128_n 0.0151035f $X=0.56 $Y=0.805 $X2=0 $Y2=0
cc_93 N_A_N_c_95_n N_B_N_c_129_n 0.0117125f $X=0.56 $Y=1.31 $X2=0 $Y2=0
cc_94 N_A_N_c_96_n N_B_N_c_130_n 0.0117125f $X=0.56 $Y=1.475 $X2=0 $Y2=0
cc_95 A_N B_N 0.0400301f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_96 N_A_N_c_98_n B_N 6.6259e-19 $X=0.56 $Y=0.97 $X2=0 $Y2=0
cc_97 A_N N_B_N_c_132_n 0.00476259f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_98 N_A_N_c_98_n N_B_N_c_132_n 0.0117125f $X=0.56 $Y=0.97 $X2=0 $Y2=0
cc_99 N_A_N_M1010_g N_A_54_55#_c_169_n 0.00568449f $X=0.61 $Y=2.195 $X2=0 $Y2=0
cc_100 N_A_N_c_94_n N_A_54_55#_c_169_n 0.00523038f $X=0.56 $Y=0.805 $X2=0 $Y2=0
cc_101 A_N N_A_54_55#_c_169_n 0.0481549f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_102 N_A_N_c_98_n N_A_54_55#_c_169_n 0.0163648f $X=0.56 $Y=0.97 $X2=0 $Y2=0
cc_103 N_A_N_M1010_g N_A_54_55#_c_177_n 0.00694169f $X=0.61 $Y=2.195 $X2=0 $Y2=0
cc_104 N_A_N_M1010_g N_A_54_55#_c_178_n 0.0167061f $X=0.61 $Y=2.195 $X2=0 $Y2=0
cc_105 N_A_N_c_96_n N_A_54_55#_c_178_n 5.13711e-19 $X=0.56 $Y=1.475 $X2=0 $Y2=0
cc_106 A_N N_A_54_55#_c_178_n 0.0229928f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_107 A_N N_A_54_55#_c_172_n 9.77165e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_108 N_A_N_c_98_n N_A_54_55#_c_172_n 0.0036397f $X=0.56 $Y=0.97 $X2=0 $Y2=0
cc_109 N_A_N_c_96_n N_A_54_55#_c_173_n 0.00397881f $X=0.56 $Y=1.475 $X2=0 $Y2=0
cc_110 A_N N_A_54_55#_c_173_n 0.00203714f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_111 N_A_N_M1010_g N_VPWR_c_523_n 0.00329204f $X=0.61 $Y=2.195 $X2=0 $Y2=0
cc_112 N_A_N_M1010_g N_VPWR_c_522_n 0.00393927f $X=0.61 $Y=2.195 $X2=0 $Y2=0
cc_113 N_A_N_c_94_n N_VGND_c_588_n 0.00290284f $X=0.56 $Y=0.805 $X2=0 $Y2=0
cc_114 A_N N_VGND_c_588_n 0.00517229f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_115 N_A_N_c_94_n N_VGND_c_592_n 0.00664473f $X=0.56 $Y=0.805 $X2=0 $Y2=0
cc_116 A_N N_VGND_c_592_n 0.00793156f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_117 N_A_N_c_94_n N_VGND_c_593_n 0.00545548f $X=0.56 $Y=0.805 $X2=0 $Y2=0
cc_118 B_N N_A_54_55#_c_167_n 7.76146e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_119 N_B_N_c_132_n N_A_54_55#_c_167_n 0.00466496f $X=1.13 $Y=0.97 $X2=0 $Y2=0
cc_120 N_B_N_c_129_n N_A_54_55#_c_168_n 0.00856803f $X=1.13 $Y=1.31 $X2=0 $Y2=0
cc_121 B_N N_A_54_55#_c_168_n 0.00126963f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_122 N_B_N_M1012_g N_A_54_55#_c_175_n 0.0111877f $X=1.04 $Y=2.195 $X2=0 $Y2=0
cc_123 N_B_N_M1012_g N_A_54_55#_c_178_n 0.0181748f $X=1.04 $Y=2.195 $X2=0 $Y2=0
cc_124 N_B_N_c_130_n N_A_54_55#_c_178_n 0.00161003f $X=1.13 $Y=1.475 $X2=0 $Y2=0
cc_125 B_N N_A_54_55#_c_178_n 0.0179287f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_126 N_B_N_M1012_g N_A_54_55#_c_170_n 8.87838e-19 $X=1.04 $Y=2.195 $X2=0 $Y2=0
cc_127 N_B_N_c_129_n N_A_54_55#_c_170_n 0.00104878f $X=1.13 $Y=1.31 $X2=0 $Y2=0
cc_128 B_N N_A_54_55#_c_170_n 0.0130555f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_129 N_B_N_M1012_g N_A_54_55#_c_171_n 0.010142f $X=1.04 $Y=2.195 $X2=0 $Y2=0
cc_130 N_B_N_c_130_n N_A_54_55#_c_171_n 0.00856803f $X=1.13 $Y=1.475 $X2=0 $Y2=0
cc_131 N_B_N_c_128_n N_A_223_55#_c_245_n 2.30416e-19 $X=1.13 $Y=0.805 $X2=0
+ $Y2=0
cc_132 B_N N_A_223_55#_c_245_n 0.0081533f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_133 N_B_N_c_132_n N_A_223_55#_c_245_n 0.00134549f $X=1.13 $Y=0.97 $X2=0 $Y2=0
cc_134 N_B_N_c_128_n N_A_332_125#_c_424_n 0.00431971f $X=1.13 $Y=0.805 $X2=0
+ $Y2=0
cc_135 B_N N_A_332_125#_c_424_n 0.00711855f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_136 N_B_N_c_132_n N_A_332_125#_c_424_n 0.0016497f $X=1.13 $Y=0.97 $X2=0 $Y2=0
cc_137 N_B_N_M1012_g N_VPWR_c_523_n 0.00329204f $X=1.04 $Y=2.195 $X2=0 $Y2=0
cc_138 N_B_N_M1012_g N_VPWR_c_522_n 0.00393927f $X=1.04 $Y=2.195 $X2=0 $Y2=0
cc_139 N_B_N_c_128_n N_VGND_c_588_n 0.00274755f $X=1.13 $Y=0.805 $X2=0 $Y2=0
cc_140 N_B_N_c_128_n N_VGND_c_590_n 0.00545548f $X=1.13 $Y=0.805 $X2=0 $Y2=0
cc_141 N_B_N_c_128_n N_VGND_c_592_n 0.00929637f $X=1.13 $Y=0.805 $X2=0 $Y2=0
cc_142 B_N N_VGND_c_592_n 0.00384164f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_143 N_A_54_55#_c_175_n N_A_223_55#_M1003_g 0.00867821f $X=1.825 $Y=2.415
+ $X2=0 $Y2=0
cc_144 N_A_54_55#_c_176_n N_A_223_55#_M1003_g 0.0203532f $X=1.825 $Y=2.565 $X2=0
+ $Y2=0
cc_145 N_A_54_55#_c_168_n N_A_223_55#_M1013_g 0.0265151f $X=2 $Y=1.23 $X2=0
+ $Y2=0
cc_146 N_A_54_55#_c_170_n N_A_223_55#_M1013_g 0.00100273f $X=1.7 $Y=1.32 $X2=0
+ $Y2=0
cc_147 N_A_54_55#_c_171_n N_A_223_55#_M1013_g 0.00656987f $X=1.7 $Y=1.32 $X2=0
+ $Y2=0
cc_148 N_A_54_55#_c_174_n N_A_223_55#_c_247_n 0.0123224f $X=1.7 $Y=1.825 $X2=0
+ $Y2=0
cc_149 N_A_54_55#_c_175_n N_A_223_55#_c_248_n 0.0123224f $X=1.825 $Y=2.415 $X2=0
+ $Y2=0
cc_150 N_A_54_55#_c_167_n N_A_223_55#_c_242_n 0.00458653f $X=2 $Y=1.155 $X2=0
+ $Y2=0
cc_151 N_A_54_55#_c_167_n N_A_223_55#_c_243_n 0.0265151f $X=2 $Y=1.155 $X2=0
+ $Y2=0
cc_152 N_A_54_55#_c_174_n N_A_223_55#_c_249_n 0.00275075f $X=1.7 $Y=1.825 $X2=0
+ $Y2=0
cc_153 N_A_54_55#_c_175_n N_A_223_55#_c_249_n 0.0172143f $X=1.825 $Y=2.415 $X2=0
+ $Y2=0
cc_154 N_A_54_55#_c_176_n N_A_223_55#_c_249_n 0.002695f $X=1.825 $Y=2.565 $X2=0
+ $Y2=0
cc_155 N_A_54_55#_c_178_n N_A_223_55#_c_249_n 0.0308076f $X=1.615 $Y=1.74 $X2=0
+ $Y2=0
cc_156 N_A_54_55#_c_178_n N_A_223_55#_c_267_n 0.00811233f $X=1.615 $Y=1.74 $X2=0
+ $Y2=0
cc_157 N_A_54_55#_c_170_n N_A_223_55#_c_267_n 0.00170109f $X=1.7 $Y=1.32 $X2=0
+ $Y2=0
cc_158 N_A_54_55#_c_171_n N_A_223_55#_c_267_n 0.00196832f $X=1.7 $Y=1.32 $X2=0
+ $Y2=0
cc_159 N_A_54_55#_c_178_n N_A_223_55#_c_244_n 5.49453e-19 $X=1.615 $Y=1.74 $X2=0
+ $Y2=0
cc_160 N_A_54_55#_c_170_n N_A_223_55#_c_244_n 6.0318e-19 $X=1.7 $Y=1.32 $X2=0
+ $Y2=0
cc_161 N_A_54_55#_c_171_n N_A_223_55#_c_244_n 0.0123224f $X=1.7 $Y=1.32 $X2=0
+ $Y2=0
cc_162 N_A_54_55#_c_167_n N_A_223_55#_c_245_n 0.00232609f $X=2 $Y=1.155 $X2=0
+ $Y2=0
cc_163 N_A_54_55#_c_175_n N_A_223_55#_c_274_n 0.00331521f $X=1.825 $Y=2.415
+ $X2=0 $Y2=0
cc_164 N_A_54_55#_c_178_n N_A_223_55#_c_274_n 0.0147756f $X=1.615 $Y=1.74 $X2=0
+ $Y2=0
cc_165 N_A_54_55#_c_168_n N_C_c_316_n 0.00111972f $X=2 $Y=1.23 $X2=0 $Y2=0
cc_166 N_A_54_55#_c_170_n N_C_c_316_n 0.0100146f $X=1.7 $Y=1.32 $X2=0 $Y2=0
cc_167 N_A_54_55#_c_171_n N_C_c_316_n 9.71899e-19 $X=1.7 $Y=1.32 $X2=0 $Y2=0
cc_168 N_A_54_55#_c_167_n N_A_332_125#_c_424_n 0.0155139f $X=2 $Y=1.155 $X2=0
+ $Y2=0
cc_169 N_A_54_55#_c_168_n N_A_332_125#_c_424_n 0.00537146f $X=2 $Y=1.23 $X2=0
+ $Y2=0
cc_170 N_A_54_55#_c_170_n N_A_332_125#_c_424_n 0.00818786f $X=1.7 $Y=1.32 $X2=0
+ $Y2=0
cc_171 N_A_54_55#_c_176_n N_A_332_125#_c_414_n 0.0017418f $X=1.825 $Y=2.565
+ $X2=0 $Y2=0
cc_172 N_A_54_55#_c_176_n N_A_332_125#_c_416_n 0.00556162f $X=1.825 $Y=2.565
+ $X2=0 $Y2=0
cc_173 N_A_54_55#_c_178_n N_VPWR_c_523_n 0.0109835f $X=1.615 $Y=1.74 $X2=0 $Y2=0
cc_174 N_A_54_55#_c_176_n N_VPWR_c_524_n 0.00417089f $X=1.825 $Y=2.565 $X2=0
+ $Y2=0
cc_175 N_A_54_55#_c_176_n N_VPWR_c_529_n 0.0065431f $X=1.825 $Y=2.565 $X2=0
+ $Y2=0
cc_176 N_A_54_55#_c_176_n N_VPWR_c_522_n 0.0129498f $X=1.825 $Y=2.565 $X2=0
+ $Y2=0
cc_177 N_A_54_55#_c_172_n N_VGND_c_592_n 0.0139896f $X=0.395 $Y=0.46 $X2=0 $Y2=0
cc_178 N_A_54_55#_c_172_n N_VGND_c_593_n 0.0194396f $X=0.395 $Y=0.46 $X2=0 $Y2=0
cc_179 N_A_223_55#_M1003_g N_C_M1011_g 0.0306565f $X=2.29 $Y=2.885 $X2=0 $Y2=0
cc_180 N_A_223_55#_c_247_n N_C_M1011_g 0.0325757f $X=2.27 $Y=2.04 $X2=0 $Y2=0
cc_181 N_A_223_55#_c_249_n N_C_M1011_g 5.15001e-19 $X=2.105 $Y=2.09 $X2=0 $Y2=0
cc_182 N_A_223_55#_c_267_n N_C_M1011_g 0.00118458f $X=2.27 $Y=1.7 $X2=0 $Y2=0
cc_183 N_A_223_55#_M1013_g N_C_c_315_n 0.0325757f $X=2.36 $Y=0.835 $X2=0 $Y2=0
cc_184 N_A_223_55#_M1013_g N_C_c_316_n 0.0111861f $X=2.36 $Y=0.835 $X2=0 $Y2=0
cc_185 N_A_223_55#_c_249_n N_C_c_316_n 9.34281e-19 $X=2.105 $Y=2.09 $X2=0 $Y2=0
cc_186 N_A_223_55#_c_267_n N_C_c_316_n 0.0216387f $X=2.27 $Y=1.7 $X2=0 $Y2=0
cc_187 N_A_223_55#_c_244_n N_C_c_316_n 0.00504688f $X=2.27 $Y=1.7 $X2=0 $Y2=0
cc_188 N_A_223_55#_M1013_g N_C_c_317_n 0.0211267f $X=2.36 $Y=0.835 $X2=0 $Y2=0
cc_189 N_A_223_55#_c_243_n N_C_c_317_n 0.00140261f $X=2.45 $Y=0.35 $X2=0 $Y2=0
cc_190 N_A_223_55#_M1013_g N_A_332_125#_c_424_n 0.0173274f $X=2.36 $Y=0.835
+ $X2=0 $Y2=0
cc_191 N_A_223_55#_c_242_n N_A_332_125#_c_424_n 0.0488888f $X=2.45 $Y=0.35 $X2=0
+ $Y2=0
cc_192 N_A_223_55#_c_243_n N_A_332_125#_c_424_n 0.00421546f $X=2.45 $Y=0.35
+ $X2=0 $Y2=0
cc_193 N_A_223_55#_M1003_g N_A_332_125#_c_414_n 9.4709e-19 $X=2.29 $Y=2.885
+ $X2=0 $Y2=0
cc_194 N_A_223_55#_M1003_g N_A_332_125#_c_415_n 0.0122928f $X=2.29 $Y=2.885
+ $X2=0 $Y2=0
cc_195 N_A_223_55#_c_248_n N_A_332_125#_c_415_n 0.00266408f $X=2.27 $Y=2.205
+ $X2=0 $Y2=0
cc_196 N_A_223_55#_c_249_n N_A_332_125#_c_415_n 0.0139658f $X=2.105 $Y=2.09
+ $X2=0 $Y2=0
cc_197 N_A_223_55#_c_248_n N_A_332_125#_c_416_n 0.00195486f $X=2.27 $Y=2.205
+ $X2=0 $Y2=0
cc_198 N_A_223_55#_c_249_n N_A_332_125#_c_416_n 0.0130089f $X=2.105 $Y=2.09
+ $X2=0 $Y2=0
cc_199 N_A_223_55#_M1003_g N_A_332_125#_c_417_n 0.00142142f $X=2.29 $Y=2.885
+ $X2=0 $Y2=0
cc_200 N_A_223_55#_c_247_n N_A_332_125#_c_417_n 0.00107243f $X=2.27 $Y=2.04
+ $X2=0 $Y2=0
cc_201 N_A_223_55#_c_248_n N_A_332_125#_c_417_n 2.10863e-19 $X=2.27 $Y=2.205
+ $X2=0 $Y2=0
cc_202 N_A_223_55#_c_249_n N_A_332_125#_c_417_n 0.0104916f $X=2.105 $Y=2.09
+ $X2=0 $Y2=0
cc_203 N_A_223_55#_c_267_n N_A_332_125#_c_417_n 0.0144692f $X=2.27 $Y=1.7 $X2=0
+ $Y2=0
cc_204 N_A_223_55#_c_267_n N_A_332_125#_c_446_n 0.00905294f $X=2.27 $Y=1.7 $X2=0
+ $Y2=0
cc_205 N_A_223_55#_c_244_n N_A_332_125#_c_446_n 6.83399e-19 $X=2.27 $Y=1.7 $X2=0
+ $Y2=0
cc_206 N_A_223_55#_c_249_n N_VPWR_c_524_n 0.00627621f $X=2.105 $Y=2.09 $X2=0
+ $Y2=0
cc_207 N_A_223_55#_M1003_g N_VPWR_c_525_n 0.00156327f $X=2.29 $Y=2.885 $X2=0
+ $Y2=0
cc_208 N_A_223_55#_M1003_g N_VPWR_c_529_n 0.00437852f $X=2.29 $Y=2.885 $X2=0
+ $Y2=0
cc_209 N_A_223_55#_M1003_g N_VPWR_c_522_n 0.00604796f $X=2.29 $Y=2.885 $X2=0
+ $Y2=0
cc_210 N_A_223_55#_c_245_n N_VGND_c_588_n 5.83564e-19 $X=1.255 $Y=0.35 $X2=0
+ $Y2=0
cc_211 N_A_223_55#_c_242_n N_VGND_c_590_n 0.0751512f $X=2.45 $Y=0.35 $X2=0 $Y2=0
cc_212 N_A_223_55#_c_243_n N_VGND_c_590_n 0.00651318f $X=2.45 $Y=0.35 $X2=0
+ $Y2=0
cc_213 N_A_223_55#_c_245_n N_VGND_c_590_n 0.0132975f $X=1.255 $Y=0.35 $X2=0
+ $Y2=0
cc_214 N_A_223_55#_c_242_n N_VGND_c_592_n 0.0453925f $X=2.45 $Y=0.35 $X2=0 $Y2=0
cc_215 N_A_223_55#_c_243_n N_VGND_c_592_n 0.0101042f $X=2.45 $Y=0.35 $X2=0 $Y2=0
cc_216 N_A_223_55#_c_245_n N_VGND_c_592_n 0.00789949f $X=1.255 $Y=0.35 $X2=0
+ $Y2=0
cc_217 N_C_M1011_g N_D_M1007_g 0.0288522f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_218 N_C_M1011_g N_D_M1002_g 0.0106306f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_219 N_C_c_316_n N_D_M1002_g 2.28806e-19 $X=2.81 $Y=1.32 $X2=0 $Y2=0
cc_220 N_C_c_317_n N_D_M1002_g 0.0623038f $X=2.81 $Y=1.155 $X2=0 $Y2=0
cc_221 N_C_M1011_g D 2.00959e-19 $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_222 N_C_M1011_g N_D_c_365_n 0.0209571f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_223 N_C_c_315_n N_A_332_125#_c_424_n 0.00460062f $X=2.81 $Y=1.32 $X2=0 $Y2=0
cc_224 N_C_c_316_n N_A_332_125#_c_424_n 0.0461452f $X=2.81 $Y=1.32 $X2=0 $Y2=0
cc_225 N_C_c_317_n N_A_332_125#_c_424_n 0.0176752f $X=2.81 $Y=1.155 $X2=0 $Y2=0
cc_226 N_C_M1011_g N_A_332_125#_c_415_n 0.00272839f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_227 N_C_M1011_g N_A_332_125#_c_417_n 0.0173416f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_228 N_C_c_315_n N_A_332_125#_c_406_n 0.00430857f $X=2.81 $Y=1.32 $X2=0 $Y2=0
cc_229 N_C_c_316_n N_A_332_125#_c_406_n 0.010344f $X=2.81 $Y=1.32 $X2=0 $Y2=0
cc_230 N_C_M1011_g N_A_332_125#_c_446_n 0.00810562f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_231 N_C_c_315_n N_A_332_125#_c_446_n 7.66562e-19 $X=2.81 $Y=1.32 $X2=0 $Y2=0
cc_232 N_C_c_316_n N_A_332_125#_c_446_n 0.0126204f $X=2.81 $Y=1.32 $X2=0 $Y2=0
cc_233 N_C_M1011_g N_A_332_125#_c_419_n 0.00778708f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_234 N_C_M1011_g N_A_332_125#_c_420_n 9.56501e-19 $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_235 N_C_M1011_g N_A_332_125#_c_407_n 0.00171438f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_236 N_C_c_315_n N_A_332_125#_c_407_n 0.00220635f $X=2.81 $Y=1.32 $X2=0 $Y2=0
cc_237 N_C_c_316_n N_A_332_125#_c_407_n 0.0147674f $X=2.81 $Y=1.32 $X2=0 $Y2=0
cc_238 N_C_c_317_n N_A_332_125#_c_407_n 0.00345085f $X=2.81 $Y=1.155 $X2=0 $Y2=0
cc_239 N_C_M1011_g N_VPWR_c_525_n 0.00151442f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_240 N_C_M1011_g N_VPWR_c_526_n 7.33522e-19 $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_241 N_C_M1011_g N_VPWR_c_531_n 0.00437852f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_242 N_C_M1011_g N_VPWR_c_522_n 0.00604796f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_243 N_C_c_317_n N_VGND_c_590_n 0.00321586f $X=2.81 $Y=1.155 $X2=0 $Y2=0
cc_244 N_C_c_317_n N_VGND_c_592_n 0.00469432f $X=2.81 $Y=1.155 $X2=0 $Y2=0
cc_245 D N_A_332_125#_c_411_n 6.33438e-19 $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_246 N_D_c_365_n N_A_332_125#_c_411_n 0.020174f $X=3.17 $Y=2.035 $X2=0 $Y2=0
cc_247 N_D_M1002_g N_A_332_125#_M1009_g 0.0203835f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_248 N_D_M1007_g N_A_332_125#_c_413_n 0.0277747f $X=3.15 $Y=2.885 $X2=0 $Y2=0
cc_249 N_D_M1002_g N_A_332_125#_c_424_n 0.0118161f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_250 N_D_M1007_g N_A_332_125#_c_417_n 0.00440992f $X=3.15 $Y=2.885 $X2=0 $Y2=0
cc_251 N_D_M1002_g N_A_332_125#_c_417_n 0.00197413f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_252 D N_A_332_125#_c_417_n 0.0121504f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_253 N_D_c_365_n N_A_332_125#_c_417_n 0.00376619f $X=3.17 $Y=2.035 $X2=0 $Y2=0
cc_254 D N_A_332_125#_c_406_n 0.00964495f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_255 N_D_c_365_n N_A_332_125#_c_406_n 0.00396944f $X=3.17 $Y=2.035 $X2=0 $Y2=0
cc_256 N_D_M1007_g N_A_332_125#_c_419_n 0.00544896f $X=3.15 $Y=2.885 $X2=0 $Y2=0
cc_257 D N_A_332_125#_c_419_n 0.00158244f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_258 N_D_c_365_n N_A_332_125#_c_419_n 7.78442e-19 $X=3.17 $Y=2.035 $X2=0 $Y2=0
cc_259 N_D_M1007_g N_A_332_125#_c_420_n 0.0017629f $X=3.15 $Y=2.885 $X2=0 $Y2=0
cc_260 N_D_M1002_g N_A_332_125#_c_407_n 0.018533f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_261 N_D_M1002_g N_A_332_125#_c_408_n 0.00217759f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_262 D N_A_332_125#_c_408_n 5.76918e-19 $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_263 N_D_M1002_g N_A_332_125#_c_482_n 0.00697856f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_264 D N_A_332_125#_c_482_n 0.0117328f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_265 N_D_c_365_n N_A_332_125#_c_482_n 8.86366e-19 $X=3.17 $Y=2.035 $X2=0 $Y2=0
cc_266 N_D_M1007_g N_A_332_125#_c_409_n 2.86238e-19 $X=3.15 $Y=2.885 $X2=0 $Y2=0
cc_267 N_D_M1002_g N_A_332_125#_c_409_n 0.00111624f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_268 D N_A_332_125#_c_409_n 0.00783131f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_269 N_D_c_365_n N_A_332_125#_c_409_n 6.7367e-19 $X=3.17 $Y=2.035 $X2=0 $Y2=0
cc_270 N_D_M1002_g N_A_332_125#_c_410_n 0.020174f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_271 N_D_M1007_g N_VPWR_c_526_n 0.00646024f $X=3.15 $Y=2.885 $X2=0 $Y2=0
cc_272 N_D_c_365_n N_VPWR_c_526_n 0.00237303f $X=3.17 $Y=2.035 $X2=0 $Y2=0
cc_273 N_D_M1007_g N_VPWR_c_531_n 0.00564095f $X=3.15 $Y=2.885 $X2=0 $Y2=0
cc_274 N_D_M1007_g N_VPWR_c_522_n 0.00961799f $X=3.15 $Y=2.885 $X2=0 $Y2=0
cc_275 N_D_M1002_g N_VGND_c_589_n 0.00558541f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_276 N_D_M1002_g N_VGND_c_590_n 0.0032778f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_277 N_D_M1002_g N_VGND_c_592_n 0.00469432f $X=3.26 $Y=0.835 $X2=0 $Y2=0
cc_278 N_A_332_125#_c_415_n N_VPWR_c_525_n 0.0139569f $X=2.655 $Y=2.52 $X2=0
+ $Y2=0
cc_279 N_A_332_125#_M1005_g N_VPWR_c_526_n 0.0100105f $X=3.62 $Y=2.885 $X2=0
+ $Y2=0
cc_280 N_A_332_125#_c_414_n N_VPWR_c_529_n 0.008231f $X=2.075 $Y=2.82 $X2=0
+ $Y2=0
cc_281 N_A_332_125#_c_415_n N_VPWR_c_529_n 0.00305343f $X=2.655 $Y=2.52 $X2=0
+ $Y2=0
cc_282 N_A_332_125#_c_415_n N_VPWR_c_531_n 0.00308568f $X=2.655 $Y=2.52 $X2=0
+ $Y2=0
cc_283 N_A_332_125#_c_420_n N_VPWR_c_531_n 0.00805099f $X=2.935 $Y=2.82 $X2=0
+ $Y2=0
cc_284 N_A_332_125#_M1005_g N_VPWR_c_533_n 0.00564095f $X=3.62 $Y=2.885 $X2=0
+ $Y2=0
cc_285 N_A_332_125#_M1008_d N_VPWR_c_522_n 0.00373063f $X=1.935 $Y=2.675 $X2=0
+ $Y2=0
cc_286 N_A_332_125#_M1011_d N_VPWR_c_522_n 0.00370075f $X=2.795 $Y=2.675 $X2=0
+ $Y2=0
cc_287 N_A_332_125#_M1005_g N_VPWR_c_522_n 0.0107615f $X=3.62 $Y=2.885 $X2=0
+ $Y2=0
cc_288 N_A_332_125#_c_414_n N_VPWR_c_522_n 0.00765087f $X=2.075 $Y=2.82 $X2=0
+ $Y2=0
cc_289 N_A_332_125#_c_415_n N_VPWR_c_522_n 0.0110027f $X=2.655 $Y=2.52 $X2=0
+ $Y2=0
cc_290 N_A_332_125#_c_420_n N_VPWR_c_522_n 0.00756149f $X=2.935 $Y=2.82 $X2=0
+ $Y2=0
cc_291 N_A_332_125#_M1005_g N_X_c_573_n 8.22342e-19 $X=3.62 $Y=2.885 $X2=0 $Y2=0
cc_292 N_A_332_125#_c_413_n N_X_c_573_n 0.00478426f $X=3.732 $Y=2.255 $X2=0
+ $Y2=0
cc_293 N_A_332_125#_c_409_n N_X_c_573_n 0.00282308f $X=3.71 $Y=1.75 $X2=0 $Y2=0
cc_294 N_A_332_125#_M1005_g X 0.0123188f $X=3.62 $Y=2.885 $X2=0 $Y2=0
cc_295 N_A_332_125#_M1009_g X 0.0374362f $X=3.845 $Y=0.835 $X2=0 $Y2=0
cc_296 N_A_332_125#_c_407_n X 0.0146696f $X=3.24 $Y=1.585 $X2=0 $Y2=0
cc_297 N_A_332_125#_c_409_n X 0.0475752f $X=3.71 $Y=1.75 $X2=0 $Y2=0
cc_298 N_A_332_125#_M1009_g N_VGND_c_589_n 0.00134801f $X=3.845 $Y=0.835 $X2=0
+ $Y2=0
cc_299 N_A_332_125#_c_424_n N_VGND_c_589_n 0.0221267f $X=3.155 $Y=0.81 $X2=0
+ $Y2=0
cc_300 N_A_332_125#_c_408_n N_VGND_c_589_n 0.00339649f $X=3.625 $Y=1.67 $X2=0
+ $Y2=0
cc_301 N_A_332_125#_c_409_n N_VGND_c_589_n 0.0026595f $X=3.71 $Y=1.75 $X2=0
+ $Y2=0
cc_302 N_A_332_125#_c_410_n N_VGND_c_589_n 0.0020631f $X=3.71 $Y=1.75 $X2=0
+ $Y2=0
cc_303 N_A_332_125#_c_424_n N_VGND_c_590_n 0.0110309f $X=3.155 $Y=0.81 $X2=0
+ $Y2=0
cc_304 N_A_332_125#_M1009_g N_VGND_c_591_n 0.00415323f $X=3.845 $Y=0.835 $X2=0
+ $Y2=0
cc_305 N_A_332_125#_M1009_g N_VGND_c_592_n 0.00469432f $X=3.845 $Y=0.835 $X2=0
+ $Y2=0
cc_306 N_A_332_125#_c_424_n N_VGND_c_592_n 0.0228564f $X=3.155 $Y=0.81 $X2=0
+ $Y2=0
cc_307 N_A_332_125#_c_424_n A_415_125# 0.00217728f $X=3.155 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_308 N_A_332_125#_c_424_n A_487_125# 0.00750127f $X=3.155 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_309 N_A_332_125#_c_424_n A_595_125# 0.00354526f $X=3.155 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_310 N_VPWR_c_522_n N_X_M1005_d 0.00344799f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_311 N_VPWR_c_533_n N_X_c_573_n 0.0180548f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_312 N_VPWR_c_522_n N_X_c_573_n 0.0157272f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_313 X N_VGND_c_589_n 0.00882845f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_314 X N_VGND_c_591_n 0.00563668f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_315 X N_VGND_c_592_n 0.00642236f $X=3.995 $Y=0.47 $X2=0 $Y2=0
