* File: sky130_fd_sc_lp__or4bb_lp.spice
* Created: Wed Sep  2 10:33:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4bb_lp.pex.spice"
.subckt sky130_fd_sc_lp__or4bb_lp  VNB VPB C_N B A D_N X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* D_N	D_N
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1012 A_116_47# N_A_86_21#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_86_21#_M1002_g A_116_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1015 A_274_47# N_C_N_M1015_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1017 N_A_318_409#_M1017_d N_C_N_M1017_g A_274_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_86_21#_M1013_d N_A_M1013_g N_A_476_125#_M1013_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.2664 PD=0.7 PS=2.35 NRD=0 NRS=165.504 M=1 R=2.8
+ SA=75000.3 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1016 A_665_125# N_A_318_409#_M1016_g N_A_86_21#_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_318_409#_M1008_g A_665_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1010 A_823_125# N_A_654_355#_M1010_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_86_21#_M1004_d N_A_654_355#_M1004_g A_823_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1007 A_981_125# N_B_M1007_g N_A_86_21#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_B_M1005_g A_981_125# VNB NSHORT L=0.15 W=0.42 AD=0.1359
+ AS=0.0441 PD=1.16 PS=0.63 NRD=22.848 NRS=14.28 M=1 R=2.8 SA=75002.7 SB=75000.4
+ A=0.063 P=1.14 MULT=1
MM1018 N_A_476_125#_M1018_d N_A_M1018_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1359 PD=1.41 PS=1.16 NRD=0 NRS=22.848 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_1284_47# N_D_N_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_654_355#_M1006_d N_D_N_M1006_g A_1284_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_86_21#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1000 N_A_318_409#_M1000_d N_C_N_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1014 A_612_400# N_A_318_409#_M1014_g N_A_505_400#_M1014_s VPB PHIGHVT L=0.25
+ W=1 AD=0.105 AS=0.285 PD=1.21 PS=2.57 NRD=9.8303 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1019 N_A_86_21#_M1019_d N_A_654_355#_M1019_g A_612_400# VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.105 PD=2.57 PS=1.21 NRD=0 NRS=9.8303 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1011 A_1076_419# N_B_M1011_g N_A_505_400#_M1011_s VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g A_1076_419# VPB PHIGHVT L=0.25 W=1 AD=0.15
+ AS=0.12 PD=1.3 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1001 N_A_654_355#_M1001_d N_D_N_M1001_g N_VPWR_M1020_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.15 PD=2.57 PS=1.3 NRD=0 NRS=3.9203 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX21_noxref VNB VPB NWDIODE A=13.214 P=19.41
c_96 VNB 0 6.61614e-20 $X=0 $Y=0
c_155 VPB 0 9.45599e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__or4bb_lp.pxi.spice"
*
.ends
*
*
