* File: sky130_fd_sc_lp__o31a_lp.spice
* Created: Fri Aug 28 11:15:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o31a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o31a_lp  VNB VPB B1 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_A_140_57#_M1009_d N_B1_M1009_g N_A_37_57#_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0651 AS=0.1533 PD=0.73 PS=1.57 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75000.3 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A3_M1004_g N_A_140_57#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0861 AS=0.0651 PD=0.83 PS=0.73 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75000.7
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1005 N_A_140_57#_M1005_d N_A2_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0861 PD=0.7 PS=0.83 NRD=0 NRS=22.848 M=1 R=2.8 SA=75001.3
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A1_M1008_g N_A_140_57#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1000 A_516_57# N_A_37_57#_M1000_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_37_57#_M1001_g A_516_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_37_57#_M1010_d N_B1_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1006 A_256_410# N_A3_M1006_g N_A_37_57#_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.135 AS=0.14 PD=1.27 PS=1.28 NRD=15.7403 NRS=0 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1002 A_360_410# N_A2_M1002_g A_256_410# VPB PHIGHVT L=0.25 W=1 AD=0.145
+ AS=0.135 PD=1.29 PS=1.27 NRD=17.7103 NRS=15.7403 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g A_360_410# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.145 PD=1.28 PS=1.29 NRD=0 NRS=17.7103 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1003 N_X_M1003_d N_A_37_57#_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX11_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o31a_lp.pxi.spice"
*
.ends
*
*
