* File: sky130_fd_sc_lp__a21oi_0.pxi.spice
* Created: Wed Sep  2 09:20:26 2020
* 
x_PM_SKY130_FD_SC_LP__A21OI_0%A2 N_A2_c_47_n N_A2_M1005_g N_A2_c_48_n
+ N_A2_M1000_g N_A2_c_49_n N_A2_c_50_n N_A2_c_55_n A2 A2 A2 N_A2_c_52_n
+ PM_SKY130_FD_SC_LP__A21OI_0%A2
x_PM_SKY130_FD_SC_LP__A21OI_0%A1 N_A1_c_92_n N_A1_M1003_g N_A1_M1002_g
+ N_A1_c_94_n A1 A1 A1 A1 N_A1_c_95_n A1 PM_SKY130_FD_SC_LP__A21OI_0%A1
x_PM_SKY130_FD_SC_LP__A21OI_0%B1 N_B1_M1001_g N_B1_M1004_g B1 B1 N_B1_c_144_n
+ PM_SKY130_FD_SC_LP__A21OI_0%B1
x_PM_SKY130_FD_SC_LP__A21OI_0%A_45_473# N_A_45_473#_M1005_s N_A_45_473#_M1002_d
+ N_A_45_473#_c_169_n N_A_45_473#_c_170_n N_A_45_473#_c_171_n
+ N_A_45_473#_c_172_n PM_SKY130_FD_SC_LP__A21OI_0%A_45_473#
x_PM_SKY130_FD_SC_LP__A21OI_0%VPWR N_VPWR_M1005_d N_VPWR_c_198_n VPWR
+ N_VPWR_c_199_n N_VPWR_c_197_n N_VPWR_c_201_n PM_SKY130_FD_SC_LP__A21OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A21OI_0%Y N_Y_M1003_d N_Y_M1004_d N_Y_c_219_n N_Y_c_220_n
+ N_Y_c_221_n N_Y_c_246_p Y Y Y Y PM_SKY130_FD_SC_LP__A21OI_0%Y
x_PM_SKY130_FD_SC_LP__A21OI_0%VGND N_VGND_M1000_s N_VGND_M1001_d N_VGND_c_249_n
+ N_VGND_c_250_n N_VGND_c_251_n N_VGND_c_252_n VGND N_VGND_c_253_n
+ N_VGND_c_254_n PM_SKY130_FD_SC_LP__A21OI_0%VGND
cc_1 VNB N_A2_c_47_n 0.00891899f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.035
cc_2 VNB N_A2_c_48_n 0.0212525f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.765
cc_3 VNB N_A2_c_49_n 0.0377727f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.84
cc_4 VNB N_A2_c_50_n 0.0185653f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_5 VNB A2 0.0327919f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A2_c_52_n 0.0344417f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_7 VNB N_A1_c_92_n 0.0199627f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.035
cc_8 VNB N_A1_M1003_g 0.0363349f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.685
cc_9 VNB N_A1_c_94_n 0.00196713f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.915
cc_10 VNB N_A1_c_95_n 0.0212611f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB A1 0.00470727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_M1001_g 0.0441286f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.185
cc_13 VNB N_B1_M1004_g 0.0157741f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.765
cc_14 VNB B1 0.0277515f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.445
cc_15 VNB N_B1_c_144_n 0.0469163f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_16 VNB N_VPWR_c_197_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_17 VNB N_Y_c_219_n 0.0166173f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.445
cc_18 VNB N_Y_c_220_n 0.00227481f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.445
cc_19 VNB N_Y_c_221_n 7.50231e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.84
cc_20 VNB Y 0.00643894f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_21 VNB N_VGND_c_249_n 0.0135235f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.765
cc_22 VNB N_VGND_c_250_n 0.0192286f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.445
cc_23 VNB N_VGND_c_251_n 0.0115183f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.915
cc_24 VNB N_VGND_c_252_n 0.0198437f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.84
cc_25 VNB N_VGND_c_253_n 0.0289699f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.11
cc_26 VNB N_VGND_c_254_n 0.128659f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_27 VPB N_A2_c_47_n 0.0265833f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.035
cc_28 VPB N_A2_M1005_g 0.0243568f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.685
cc_29 VPB N_A2_c_55_n 0.0239374f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.11
cc_30 VPB A2 0.0117413f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_31 VPB N_A1_M1002_g 0.0416532f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.445
cc_32 VPB N_A1_c_94_n 0.0194013f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.915
cc_33 VPB A1 0.0041384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_B1_M1004_g 0.0542542f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.765
cc_35 VPB N_A_45_473#_c_169_n 0.0360932f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.445
cc_36 VPB N_A_45_473#_c_170_n 0.0141727f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.915
cc_37 VPB N_A_45_473#_c_171_n 0.0092819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_45_473#_c_172_n 0.00567993f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_39 VPB N_VPWR_c_198_n 0.0101805f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.445
cc_40 VPB N_VPWR_c_199_n 0.0291462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_197_n 0.0561069f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_42 VPB N_VPWR_c_201_n 0.0253276f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_Y_c_220_n 0.00123566f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.445
cc_44 VPB N_Y_c_221_n 0.00286468f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.84
cc_45 VPB Y 0.00441374f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_46 VPB Y 0.0626631f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.51
cc_47 N_A2_c_50_n N_A1_c_92_n 0.0113859f $X=0.27 $Y=1.51 $X2=0 $Y2=0
cc_48 N_A2_c_48_n N_A1_M1003_g 0.0443938f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_49 A2 N_A1_M1003_g 4.13112e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_50 N_A2_c_52_n N_A1_M1003_g 0.00282005f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_51 N_A2_c_47_n N_A1_M1002_g 0.003558f $X=0.36 $Y=2.035 $X2=0 $Y2=0
cc_52 N_A2_c_55_n N_A1_M1002_g 0.019345f $X=0.565 $Y=2.11 $X2=0 $Y2=0
cc_53 N_A2_c_47_n N_A1_c_94_n 0.0113859f $X=0.36 $Y=2.035 $X2=0 $Y2=0
cc_54 N_A2_c_48_n A1 0.0128912f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_55 N_A2_c_48_n A1 0.00284572f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_56 N_A2_c_49_n A1 0.00834966f $X=0.605 $Y=0.84 $X2=0 $Y2=0
cc_57 A2 A1 0.0829008f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_58 N_A2_c_49_n N_A1_c_95_n 2.77132e-19 $X=0.605 $Y=0.84 $X2=0 $Y2=0
cc_59 A2 N_A1_c_95_n 6.55052e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_60 N_A2_c_52_n N_A1_c_95_n 0.0113859f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_61 N_A2_c_55_n A1 4.97996e-19 $X=0.565 $Y=2.11 $X2=0 $Y2=0
cc_62 N_A2_c_52_n A1 0.00569836f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_63 N_A2_M1005_g N_A_45_473#_c_169_n 0.00572322f $X=0.565 $Y=2.685 $X2=0 $Y2=0
cc_64 N_A2_c_55_n N_A_45_473#_c_169_n 0.00517434f $X=0.565 $Y=2.11 $X2=0 $Y2=0
cc_65 N_A2_c_55_n N_A_45_473#_c_170_n 0.0133131f $X=0.565 $Y=2.11 $X2=0 $Y2=0
cc_66 N_A2_c_47_n N_A_45_473#_c_171_n 0.00439715f $X=0.36 $Y=2.035 $X2=0 $Y2=0
cc_67 N_A2_c_50_n N_A_45_473#_c_171_n 3.91957e-19 $X=0.27 $Y=1.51 $X2=0 $Y2=0
cc_68 N_A2_c_55_n N_A_45_473#_c_171_n 0.00535942f $X=0.565 $Y=2.11 $X2=0 $Y2=0
cc_69 A2 N_A_45_473#_c_171_n 0.0190199f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_70 N_A2_M1005_g N_VPWR_c_198_n 0.00315881f $X=0.565 $Y=2.685 $X2=0 $Y2=0
cc_71 N_A2_M1005_g N_VPWR_c_197_n 0.0100922f $X=0.565 $Y=2.685 $X2=0 $Y2=0
cc_72 N_A2_M1005_g N_VPWR_c_201_n 0.00499542f $X=0.565 $Y=2.685 $X2=0 $Y2=0
cc_73 N_A2_c_49_n N_VGND_c_249_n 0.00198834f $X=0.605 $Y=0.84 $X2=0 $Y2=0
cc_74 N_A2_c_48_n N_VGND_c_250_n 0.00708294f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_75 N_A2_c_49_n N_VGND_c_250_n 0.00789683f $X=0.605 $Y=0.84 $X2=0 $Y2=0
cc_76 A2 N_VGND_c_250_n 0.0164715f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_77 N_A2_c_48_n N_VGND_c_253_n 0.00460899f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_78 N_A2_c_49_n N_VGND_c_253_n 0.00116078f $X=0.605 $Y=0.84 $X2=0 $Y2=0
cc_79 N_A2_c_48_n N_VGND_c_254_n 0.00824889f $X=0.605 $Y=0.765 $X2=0 $Y2=0
cc_80 N_A2_c_49_n N_VGND_c_254_n 0.00431698f $X=0.605 $Y=0.84 $X2=0 $Y2=0
cc_81 A2 N_VGND_c_254_n 0.00528744f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_82 N_A1_M1003_g N_B1_M1001_g 0.0267943f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A1_c_94_n N_B1_M1004_g 0.0267943f $X=0.872 $Y=1.825 $X2=0 $Y2=0
cc_84 A1 N_B1_M1004_g 3.14862e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_85 A1 N_B1_M1004_g 3.74626e-19 $X=0.72 $Y=0.925 $X2=0 $Y2=0
cc_86 N_A1_c_95_n N_B1_c_144_n 0.0267943f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_87 N_A1_M1002_g N_A_45_473#_c_170_n 0.019272f $X=0.995 $Y=2.685 $X2=0 $Y2=0
cc_88 N_A1_c_94_n N_A_45_473#_c_170_n 0.00165695f $X=0.872 $Y=1.825 $X2=0 $Y2=0
cc_89 A1 N_A_45_473#_c_170_n 0.0297766f $X=0.72 $Y=0.925 $X2=0 $Y2=0
cc_90 N_A1_M1002_g N_A_45_473#_c_172_n 0.0027375f $X=0.995 $Y=2.685 $X2=0 $Y2=0
cc_91 N_A1_M1002_g N_VPWR_c_198_n 0.00315881f $X=0.995 $Y=2.685 $X2=0 $Y2=0
cc_92 N_A1_M1002_g N_VPWR_c_199_n 0.00499542f $X=0.995 $Y=2.685 $X2=0 $Y2=0
cc_93 N_A1_M1002_g N_VPWR_c_197_n 0.00971452f $X=0.995 $Y=2.685 $X2=0 $Y2=0
cc_94 N_A1_M1003_g N_Y_c_219_n 0.00734857f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_95 A1 N_Y_c_219_n 0.0786549f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_96 N_A1_c_92_n N_Y_c_221_n 0.0017918f $X=0.872 $Y=1.628 $X2=0 $Y2=0
cc_97 A1 N_Y_c_221_n 0.0156394f $X=0.72 $Y=0.925 $X2=0 $Y2=0
cc_98 A1 Y 0.0026042f $X=0.72 $Y=0.925 $X2=0 $Y2=0
cc_99 A1 N_VGND_c_250_n 0.0162222f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_100 N_A1_M1003_g N_VGND_c_253_n 0.00580047f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_101 A1 N_VGND_c_253_n 0.00887562f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_102 A1 N_VGND_c_253_n 7.70547e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_103 N_A1_M1003_g N_VGND_c_254_n 0.0107423f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_104 A1 N_VGND_c_254_n 0.0104175f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_105 A1 N_VGND_c_254_n 0.00123759f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_106 A1 A_136_47# 0.00162168f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_107 N_B1_M1004_g N_A_45_473#_c_170_n 0.00151072f $X=1.425 $Y=2.685 $X2=0
+ $Y2=0
cc_108 N_B1_M1004_g N_A_45_473#_c_172_n 0.00166677f $X=1.425 $Y=2.685 $X2=0
+ $Y2=0
cc_109 N_B1_M1004_g N_VPWR_c_199_n 0.00499542f $X=1.425 $Y=2.685 $X2=0 $Y2=0
cc_110 N_B1_M1004_g N_VPWR_c_197_n 0.0102811f $X=1.425 $Y=2.685 $X2=0 $Y2=0
cc_111 N_B1_M1001_g N_Y_c_219_n 0.0126379f $X=1.425 $Y=0.445 $X2=0 $Y2=0
cc_112 B1 N_Y_c_219_n 0.0470278f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_113 N_B1_M1004_g N_Y_c_220_n 0.0201638f $X=1.425 $Y=2.685 $X2=0 $Y2=0
cc_114 B1 N_Y_c_220_n 0.00410256f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_115 N_B1_c_144_n N_Y_c_220_n 2.32935e-19 $X=1.62 $Y=1.27 $X2=0 $Y2=0
cc_116 B1 Y 0.0284313f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_117 N_B1_c_144_n Y 0.00671852f $X=1.62 $Y=1.27 $X2=0 $Y2=0
cc_118 N_B1_M1004_g Y 0.0190484f $X=1.425 $Y=2.685 $X2=0 $Y2=0
cc_119 N_B1_M1001_g N_VGND_c_252_n 0.00520298f $X=1.425 $Y=0.445 $X2=0 $Y2=0
cc_120 B1 N_VGND_c_252_n 0.0239432f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_121 N_B1_c_144_n N_VGND_c_252_n 0.00100672f $X=1.62 $Y=1.27 $X2=0 $Y2=0
cc_122 N_B1_M1001_g N_VGND_c_253_n 0.00585385f $X=1.425 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B1_M1001_g N_VGND_c_254_n 0.0104397f $X=1.425 $Y=0.445 $X2=0 $Y2=0
cc_124 B1 N_VGND_c_254_n 0.00406817f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_125 N_A_45_473#_c_169_n N_VPWR_c_198_n 0.00308399f $X=0.35 $Y=2.51 $X2=0
+ $Y2=0
cc_126 N_A_45_473#_c_170_n N_VPWR_c_198_n 0.0226353f $X=1.085 $Y=2.09 $X2=0
+ $Y2=0
cc_127 N_A_45_473#_c_172_n N_VPWR_c_198_n 0.00305408f $X=1.21 $Y=2.51 $X2=0
+ $Y2=0
cc_128 N_A_45_473#_c_172_n N_VPWR_c_199_n 0.0137636f $X=1.21 $Y=2.51 $X2=0 $Y2=0
cc_129 N_A_45_473#_c_169_n N_VPWR_c_197_n 0.0109155f $X=0.35 $Y=2.51 $X2=0 $Y2=0
cc_130 N_A_45_473#_c_172_n N_VPWR_c_197_n 0.00958901f $X=1.21 $Y=2.51 $X2=0
+ $Y2=0
cc_131 N_A_45_473#_c_169_n N_VPWR_c_201_n 0.0156677f $X=0.35 $Y=2.51 $X2=0 $Y2=0
cc_132 N_A_45_473#_c_170_n N_Y_c_220_n 0.00348911f $X=1.085 $Y=2.09 $X2=0 $Y2=0
cc_133 N_A_45_473#_c_170_n N_Y_c_221_n 0.0133845f $X=1.085 $Y=2.09 $X2=0 $Y2=0
cc_134 N_A_45_473#_c_170_n Y 0.0150111f $X=1.085 $Y=2.09 $X2=0 $Y2=0
cc_135 N_A_45_473#_c_172_n Y 0.016916f $X=1.21 $Y=2.51 $X2=0 $Y2=0
cc_136 N_VPWR_c_199_n Y 0.0175718f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_137 N_VPWR_c_197_n Y 0.0122421f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_138 N_Y_c_246_p N_VGND_c_253_n 0.0124106f $X=1.21 $Y=0.445 $X2=0 $Y2=0
cc_139 N_Y_M1003_d N_VGND_c_254_n 0.00354733f $X=1.07 $Y=0.235 $X2=0 $Y2=0
cc_140 N_Y_c_246_p N_VGND_c_254_n 0.0092923f $X=1.21 $Y=0.445 $X2=0 $Y2=0
cc_141 N_VGND_c_254_n A_136_47# 0.00208911f $X=1.68 $Y=0 $X2=-0.19 $Y2=-0.245
