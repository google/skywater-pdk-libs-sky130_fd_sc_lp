# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand4bb_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nand4bb_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465000 0.855000 0.835000 1.525000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 0.765000 3.720000 1.085000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.490000 1.615000 2.820000 2.150000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.615000 3.360000 2.150000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  0.679700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 2.290000 1.685000 2.330000 ;
        RECT 1.355000 2.330000 3.055000 2.520000 ;
        RECT 1.355000 2.520000 1.685000 3.065000 ;
        RECT 1.465000 0.265000 1.795000 0.675000 ;
        RECT 1.600000 0.675000 1.770000 1.940000 ;
        RECT 1.600000 1.940000 2.275000 2.110000 ;
        RECT 2.045000 2.110000 2.275000 2.330000 ;
        RECT 2.725000 2.520000 3.055000 3.065000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.265000 0.445000 0.675000 ;
      RECT 0.115000  0.675000 0.285000 1.725000 ;
      RECT 0.115000  1.725000 1.420000 1.895000 ;
      RECT 0.115000  1.895000 0.625000 3.065000 ;
      RECT 0.825000  2.075000 1.155000 3.245000 ;
      RECT 0.905000  0.085000 1.235000 0.675000 ;
      RECT 1.090000  1.225000 1.420000 1.725000 ;
      RECT 1.885000  2.700000 2.215000 3.245000 ;
      RECT 1.950000  1.090000 2.280000 1.265000 ;
      RECT 1.950000  1.265000 4.205000 1.435000 ;
      RECT 1.950000  1.435000 2.280000 1.760000 ;
      RECT 3.035000  0.085000 3.365000 0.585000 ;
      RECT 3.255000  2.330000 3.585000 3.245000 ;
      RECT 3.825000  1.435000 4.205000 3.065000 ;
      RECT 3.875000  0.295000 4.205000 0.585000 ;
      RECT 4.035000  0.585000 4.205000 1.265000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__nand4bb_lp
