* File: sky130_fd_sc_lp__or3_1.pxi.spice
* Created: Fri Aug 28 11:23:06 2020
* 
x_PM_SKY130_FD_SC_LP__OR3_1%C N_C_c_56_n N_C_M1007_g N_C_M1003_g N_C_c_59_n C C
+ C N_C_c_61_n PM_SKY130_FD_SC_LP__OR3_1%C
x_PM_SKY130_FD_SC_LP__OR3_1%B N_B_M1004_g N_B_M1006_g N_B_c_97_n N_B_c_98_n
+ N_B_c_99_n B B B N_B_c_102_n PM_SKY130_FD_SC_LP__OR3_1%B
x_PM_SKY130_FD_SC_LP__OR3_1%A N_A_M1005_g N_A_M1002_g A N_A_c_145_n N_A_c_146_n
+ PM_SKY130_FD_SC_LP__OR3_1%A
x_PM_SKY130_FD_SC_LP__OR3_1%A_47_47# N_A_47_47#_M1007_s N_A_47_47#_M1006_d
+ N_A_47_47#_M1003_s N_A_47_47#_M1001_g N_A_47_47#_M1000_g N_A_47_47#_c_188_n
+ N_A_47_47#_c_198_n N_A_47_47#_c_199_n N_A_47_47#_c_189_n N_A_47_47#_c_190_n
+ N_A_47_47#_c_191_n N_A_47_47#_c_192_n N_A_47_47#_c_193_n N_A_47_47#_c_194_n
+ N_A_47_47#_c_201_n N_A_47_47#_c_195_n PM_SKY130_FD_SC_LP__OR3_1%A_47_47#
x_PM_SKY130_FD_SC_LP__OR3_1%VPWR N_VPWR_M1005_d N_VPWR_c_271_n VPWR
+ N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_270_n N_VPWR_c_275_n
+ PM_SKY130_FD_SC_LP__OR3_1%VPWR
x_PM_SKY130_FD_SC_LP__OR3_1%X N_X_M1001_d N_X_M1000_d X X X X X X X N_X_c_296_n
+ X PM_SKY130_FD_SC_LP__OR3_1%X
x_PM_SKY130_FD_SC_LP__OR3_1%VGND N_VGND_M1007_d N_VGND_M1002_d N_VGND_c_312_n
+ N_VGND_c_313_n N_VGND_c_314_n VGND N_VGND_c_315_n N_VGND_c_316_n
+ N_VGND_c_317_n N_VGND_c_318_n PM_SKY130_FD_SC_LP__OR3_1%VGND
cc_1 VNB N_C_c_56_n 0.0221631f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.33
cc_2 VNB N_C_M1007_g 0.0266368f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.445
cc_3 VNB N_C_M1003_g 0.00839874f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.52
cc_4 VNB N_C_c_59_n 0.0192585f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.51
cc_5 VNB C 0.00908989f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_C_c_61_n 0.0188875f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.005
cc_7 VNB N_B_M1004_g 0.0096867f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.84
cc_8 VNB N_B_c_97_n 0.0188688f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.52
cc_9 VNB N_B_c_98_n 0.0265985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_99_n 0.016954f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_11 VNB B 0.00227293f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB B 0.00281079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_102_n 0.0262998f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.005
cc_14 VNB N_A_M1002_g 0.0475135f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.51
cc_15 VNB N_A_c_145_n 0.027925f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_16 VNB N_A_c_146_n 0.00179113f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_17 VNB N_A_47_47#_M1000_g 0.00774838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_47_47#_c_188_n 0.0531037f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.005
cc_19 VNB N_A_47_47#_c_189_n 0.00379815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_47_47#_c_190_n 0.0091137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_47_47#_c_191_n 0.00326668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_47_47#_c_192_n 9.40502e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_47_47#_c_193_n 0.0389185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_47_47#_c_194_n 0.0158966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_47_47#_c_195_n 0.0199601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_270_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.005
cc_27 VNB X 0.00857108f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.52
cc_28 VNB N_X_c_296_n 0.0197966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB X 0.0365685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_312_n 0.00785774f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.51
cc_31 VNB N_VGND_c_313_n 0.0154214f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_32 VNB N_VGND_c_314_n 0.00624797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_315_n 0.0195486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_316_n 0.169619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_317_n 0.019355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_318_n 0.0157008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_C_M1003_g 0.0539534f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.52
cc_38 VPB C 0.0033408f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_39 VPB N_B_M1004_g 0.0446861f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.84
cc_40 VPB B 0.00266679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_M1005_g 0.0503489f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.84
cc_42 VPB N_A_c_145_n 0.00751414f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_43 VPB N_A_c_146_n 0.00343785f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_44 VPB N_A_47_47#_M1000_g 0.0258036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_47_47#_c_188_n 0.014291f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.005
cc_46 VPB N_A_47_47#_c_198_n 0.0389246f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.84
cc_47 VPB N_A_47_47#_c_199_n 0.043299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_47_47#_c_192_n 0.00194411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_47_47#_c_201_n 0.0180061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_271_n 0.0200871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_272_n 0.0520077f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_52 VPB N_VPWR_c_273_n 0.0153759f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.005
cc_53 VPB N_VPWR_c_270_n 0.0817726f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.005
cc_54 VPB N_VPWR_c_275_n 0.0121291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB X 0.0561727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 N_C_c_59_n N_B_M1004_g 0.0635351f $X=0.605 $Y=1.51 $X2=0 $Y2=0
cc_57 C N_B_M1004_g 9.96382e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_58 N_C_M1007_g N_B_c_97_n 0.00530812f $X=0.575 $Y=0.445 $X2=0 $Y2=0
cc_59 N_C_M1007_g N_B_c_98_n 0.00247226f $X=0.575 $Y=0.445 $X2=0 $Y2=0
cc_60 C N_B_c_98_n 0.00404893f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_61 N_C_c_61_n N_B_c_98_n 0.0123588f $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_62 N_C_c_59_n N_B_c_99_n 0.0123588f $X=0.605 $Y=1.51 $X2=0 $Y2=0
cc_63 C B 0.0758793f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_64 N_C_c_61_n B 3.15738e-19 $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_65 N_C_c_56_n B 3.15738e-19 $X=0.605 $Y=1.33 $X2=0 $Y2=0
cc_66 N_C_c_59_n B 9.63227e-19 $X=0.605 $Y=1.51 $X2=0 $Y2=0
cc_67 N_C_c_56_n N_B_c_102_n 0.0123588f $X=0.605 $Y=1.33 $X2=0 $Y2=0
cc_68 N_C_M1007_g N_A_47_47#_c_188_n 0.00595625f $X=0.575 $Y=0.445 $X2=0 $Y2=0
cc_69 N_C_M1003_g N_A_47_47#_c_188_n 0.00644961f $X=0.71 $Y=2.52 $X2=0 $Y2=0
cc_70 C N_A_47_47#_c_188_n 0.0763598f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_71 N_C_c_61_n N_A_47_47#_c_188_n 0.0167061f $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_72 N_C_M1003_g N_A_47_47#_c_198_n 0.0181142f $X=0.71 $Y=2.52 $X2=0 $Y2=0
cc_73 N_C_M1003_g N_A_47_47#_c_199_n 0.0125268f $X=0.71 $Y=2.52 $X2=0 $Y2=0
cc_74 C N_A_47_47#_c_199_n 0.0147309f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_75 N_C_c_61_n N_A_47_47#_c_194_n 0.00167815f $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_76 N_C_M1003_g N_A_47_47#_c_201_n 0.00592313f $X=0.71 $Y=2.52 $X2=0 $Y2=0
cc_77 N_C_c_59_n N_A_47_47#_c_201_n 0.00327862f $X=0.605 $Y=1.51 $X2=0 $Y2=0
cc_78 C N_A_47_47#_c_201_n 0.0151399f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_79 N_C_M1003_g N_VPWR_c_272_n 0.00412289f $X=0.71 $Y=2.52 $X2=0 $Y2=0
cc_80 N_C_M1003_g N_VPWR_c_270_n 0.00476395f $X=0.71 $Y=2.52 $X2=0 $Y2=0
cc_81 N_C_M1007_g N_VGND_c_316_n 0.00779134f $X=0.575 $Y=0.445 $X2=0 $Y2=0
cc_82 C N_VGND_c_316_n 0.00617285f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_83 N_C_c_61_n N_VGND_c_316_n 2.78168e-19 $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_84 N_C_M1007_g N_VGND_c_317_n 0.00585385f $X=0.575 $Y=0.445 $X2=0 $Y2=0
cc_85 N_C_M1007_g N_VGND_c_318_n 0.00394437f $X=0.575 $Y=0.445 $X2=0 $Y2=0
cc_86 C N_VGND_c_318_n 0.0134349f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_87 N_C_c_61_n N_VGND_c_318_n 7.14317e-19 $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_88 N_B_c_97_n N_A_M1002_g 0.0186726f $X=1.212 $Y=0.765 $X2=0 $Y2=0
cc_89 B N_A_M1002_g 8.93485e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_90 N_B_c_102_n N_A_M1002_g 0.0123197f $X=1.16 $Y=0.93 $X2=0 $Y2=0
cc_91 N_B_M1004_g N_A_c_145_n 0.0595035f $X=1.15 $Y=2.52 $X2=0 $Y2=0
cc_92 N_B_c_99_n N_A_c_145_n 0.00611772f $X=1.16 $Y=1.435 $X2=0 $Y2=0
cc_93 B N_A_c_145_n 5.32097e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_94 B N_A_c_145_n 0.0010583f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_95 N_B_M1004_g N_A_c_146_n 9.12977e-19 $X=1.15 $Y=2.52 $X2=0 $Y2=0
cc_96 B N_A_c_146_n 0.0273009f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_97 N_B_M1004_g N_A_47_47#_c_198_n 0.00303308f $X=1.15 $Y=2.52 $X2=0 $Y2=0
cc_98 N_B_M1004_g N_A_47_47#_c_199_n 0.0173694f $X=1.15 $Y=2.52 $X2=0 $Y2=0
cc_99 N_B_c_99_n N_A_47_47#_c_199_n 0.00134048f $X=1.16 $Y=1.435 $X2=0 $Y2=0
cc_100 B N_A_47_47#_c_199_n 0.0250495f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_101 N_B_c_97_n N_A_47_47#_c_189_n 0.00425232f $X=1.212 $Y=0.765 $X2=0 $Y2=0
cc_102 B N_A_47_47#_c_189_n 0.024367f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_103 N_B_c_102_n N_A_47_47#_c_189_n 0.00137665f $X=1.16 $Y=0.93 $X2=0 $Y2=0
cc_104 B N_A_47_47#_c_191_n 0.0141595f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_105 N_B_c_102_n N_A_47_47#_c_191_n 0.00150393f $X=1.16 $Y=0.93 $X2=0 $Y2=0
cc_106 N_B_M1004_g N_VPWR_c_271_n 0.00262113f $X=1.15 $Y=2.52 $X2=0 $Y2=0
cc_107 N_B_M1004_g N_VPWR_c_272_n 0.00428744f $X=1.15 $Y=2.52 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_VPWR_c_270_n 0.00476395f $X=1.15 $Y=2.52 $X2=0 $Y2=0
cc_109 N_B_c_97_n N_VGND_c_313_n 0.00525069f $X=1.212 $Y=0.765 $X2=0 $Y2=0
cc_110 N_B_c_97_n N_VGND_c_316_n 0.00895133f $X=1.212 $Y=0.765 $X2=0 $Y2=0
cc_111 B N_VGND_c_316_n 0.00101398f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_112 N_B_c_97_n N_VGND_c_318_n 0.00844217f $X=1.212 $Y=0.765 $X2=0 $Y2=0
cc_113 N_B_c_98_n N_VGND_c_318_n 0.00308104f $X=1.212 $Y=0.915 $X2=0 $Y2=0
cc_114 B N_VGND_c_318_n 0.0203615f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_115 N_A_M1005_g N_A_47_47#_M1000_g 0.0101814f $X=1.61 $Y=2.52 $X2=0 $Y2=0
cc_116 N_A_c_145_n N_A_47_47#_M1000_g 0.00369338f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_117 N_A_c_146_n N_A_47_47#_M1000_g 3.71417e-19 $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A_M1005_g N_A_47_47#_c_199_n 0.0183398f $X=1.61 $Y=2.52 $X2=0 $Y2=0
cc_119 N_A_c_145_n N_A_47_47#_c_199_n 0.00121933f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_120 N_A_c_146_n N_A_47_47#_c_199_n 0.0306592f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_121 N_A_M1002_g N_A_47_47#_c_189_n 0.0132895f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_M1002_g N_A_47_47#_c_190_n 0.01283f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_123 N_A_c_145_n N_A_47_47#_c_190_n 8.67805e-19 $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_124 N_A_c_146_n N_A_47_47#_c_190_n 0.012927f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_125 N_A_M1002_g N_A_47_47#_c_191_n 0.0021362f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_c_145_n N_A_47_47#_c_191_n 0.00513529f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_127 N_A_c_146_n N_A_47_47#_c_191_n 0.0182324f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_128 N_A_M1005_g N_A_47_47#_c_192_n 0.0033415f $X=1.61 $Y=2.52 $X2=0 $Y2=0
cc_129 N_A_M1002_g N_A_47_47#_c_192_n 5.63654e-19 $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_130 N_A_c_145_n N_A_47_47#_c_192_n 0.00218533f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A_c_146_n N_A_47_47#_c_192_n 0.0209236f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A_M1002_g N_A_47_47#_c_193_n 0.00871166f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_133 N_A_c_145_n N_A_47_47#_c_193_n 0.011093f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A_c_146_n N_A_47_47#_c_193_n 3.23253e-19 $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A_M1002_g N_A_47_47#_c_195_n 0.0185394f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_136 N_A_M1005_g N_VPWR_c_271_n 0.0152266f $X=1.61 $Y=2.52 $X2=0 $Y2=0
cc_137 N_A_M1005_g N_VPWR_c_272_n 0.00356352f $X=1.61 $Y=2.52 $X2=0 $Y2=0
cc_138 N_A_M1005_g N_VPWR_c_270_n 0.00400172f $X=1.61 $Y=2.52 $X2=0 $Y2=0
cc_139 N_A_M1002_g N_VGND_c_312_n 0.00469456f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A_M1002_g N_VGND_c_313_n 0.0057945f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A_M1002_g N_VGND_c_316_n 0.0107913f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_M1002_g N_VGND_c_318_n 5.25694e-19 $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A_47_47#_c_199_n N_VPWR_M1005_d 0.00421882f $X=2.115 $Y=2.03 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A_47_47#_c_192_n N_VPWR_M1005_d 0.0014253f $X=2.27 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_47_47#_M1000_g N_VPWR_c_271_n 0.0182665f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_47_47#_c_199_n N_VPWR_c_271_n 0.0515907f $X=2.115 $Y=2.03 $X2=0 $Y2=0
cc_147 N_A_47_47#_c_198_n N_VPWR_c_272_n 0.0136179f $X=0.495 $Y=2.52 $X2=0 $Y2=0
cc_148 N_A_47_47#_M1000_g N_VPWR_c_273_n 0.00486043f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_47_47#_M1000_g N_VPWR_c_270_n 0.00917987f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_47_47#_c_198_n N_VPWR_c_270_n 0.01834f $X=0.495 $Y=2.52 $X2=0 $Y2=0
cc_151 N_A_47_47#_c_193_n X 0.00199106f $X=2.27 $Y=1.35 $X2=0 $Y2=0
cc_152 N_A_47_47#_c_195_n X 0.0032648f $X=2.292 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A_47_47#_c_195_n N_X_c_296_n 0.00500623f $X=2.292 $Y=1.185 $X2=0 $Y2=0
cc_154 N_A_47_47#_c_190_n X 0.0139703f $X=2.115 $Y=1.17 $X2=0 $Y2=0
cc_155 N_A_47_47#_c_192_n X 0.046892f $X=2.27 $Y=1.35 $X2=0 $Y2=0
cc_156 N_A_47_47#_c_193_n X 0.0189904f $X=2.27 $Y=1.35 $X2=0 $Y2=0
cc_157 N_A_47_47#_c_195_n X 0.0067549f $X=2.292 $Y=1.185 $X2=0 $Y2=0
cc_158 N_A_47_47#_c_189_n N_VGND_c_312_n 0.0335849f $X=1.57 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_47_47#_c_190_n N_VGND_c_312_n 0.0271923f $X=2.115 $Y=1.17 $X2=0 $Y2=0
cc_160 N_A_47_47#_c_193_n N_VGND_c_312_n 6.26875e-19 $X=2.27 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A_47_47#_c_195_n N_VGND_c_312_n 0.00496795f $X=2.292 $Y=1.185 $X2=0
+ $Y2=0
cc_162 N_A_47_47#_c_189_n N_VGND_c_313_n 0.0126721f $X=1.57 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_47_47#_c_195_n N_VGND_c_315_n 0.0054895f $X=2.292 $Y=1.185 $X2=0
+ $Y2=0
cc_164 N_A_47_47#_M1007_s N_VGND_c_316_n 0.0022721f $X=0.235 $Y=0.235 $X2=0
+ $Y2=0
cc_165 N_A_47_47#_M1006_d N_VGND_c_316_n 0.00351258f $X=1.43 $Y=0.235 $X2=0
+ $Y2=0
cc_166 N_A_47_47#_c_189_n N_VGND_c_316_n 0.00949526f $X=1.57 $Y=0.445 $X2=0
+ $Y2=0
cc_167 N_A_47_47#_c_194_n N_VGND_c_316_n 0.0150532f $X=0.36 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_47_47#_c_195_n N_VGND_c_316_n 0.011168f $X=2.292 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A_47_47#_c_194_n N_VGND_c_317_n 0.0219443f $X=0.36 $Y=0.445 $X2=0 $Y2=0
cc_170 N_VPWR_c_270_n N_X_M1000_d 0.00371702f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_171 N_VPWR_c_273_n X 0.0178111f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_270_n X 0.0100304f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_173 N_X_c_296_n N_VGND_c_315_n 0.0264034f $X=2.545 $Y=0.42 $X2=0 $Y2=0
cc_174 N_X_M1001_d N_VGND_c_316_n 0.00215158f $X=2.405 $Y=0.235 $X2=0 $Y2=0
cc_175 N_X_c_296_n N_VGND_c_316_n 0.0154782f $X=2.545 $Y=0.42 $X2=0 $Y2=0
