* File: sky130_fd_sc_lp__or4bb_4.pxi.spice
* Created: Fri Aug 28 11:26:44 2020
* 
x_PM_SKY130_FD_SC_LP__OR4BB_4%C_N N_C_N_c_104_n N_C_N_M1011_g N_C_N_M1014_g
+ N_C_N_c_106_n N_C_N_c_107_n C_N C_N PM_SKY130_FD_SC_LP__OR4BB_4%C_N
x_PM_SKY130_FD_SC_LP__OR4BB_4%A N_A_M1001_g N_A_M1004_g A A N_A_c_134_n
+ N_A_c_135_n PM_SKY130_FD_SC_LP__OR4BB_4%A
x_PM_SKY130_FD_SC_LP__OR4BB_4%B N_B_M1009_g N_B_M1015_g B N_B_c_170_n
+ N_B_c_171_n PM_SKY130_FD_SC_LP__OR4BB_4%B
x_PM_SKY130_FD_SC_LP__OR4BB_4%A_79_137# N_A_79_137#_M1011_s N_A_79_137#_M1014_s
+ N_A_79_137#_M1013_g N_A_79_137#_M1007_g N_A_79_137#_c_208_n
+ N_A_79_137#_c_222_n N_A_79_137#_c_214_n N_A_79_137#_c_209_n
+ N_A_79_137#_c_210_n N_A_79_137#_c_211_n PM_SKY130_FD_SC_LP__OR4BB_4%A_79_137#
x_PM_SKY130_FD_SC_LP__OR4BB_4%A_528_27# N_A_528_27#_M1012_d N_A_528_27#_M1008_d
+ N_A_528_27#_c_282_n N_A_528_27#_M1018_g N_A_528_27#_M1002_g
+ N_A_528_27#_c_284_n N_A_528_27#_c_285_n N_A_528_27#_c_286_n
+ N_A_528_27#_c_310_p N_A_528_27#_c_287_n N_A_528_27#_c_288_n
+ N_A_528_27#_c_291_n PM_SKY130_FD_SC_LP__OR4BB_4%A_528_27#
x_PM_SKY130_FD_SC_LP__OR4BB_4%A_270_53# N_A_270_53#_M1001_d N_A_270_53#_M1007_d
+ N_A_270_53#_M1002_d N_A_270_53#_M1003_g N_A_270_53#_M1000_g
+ N_A_270_53#_M1006_g N_A_270_53#_M1005_g N_A_270_53#_M1016_g
+ N_A_270_53#_M1010_g N_A_270_53#_M1017_g N_A_270_53#_M1019_g
+ N_A_270_53#_c_375_n N_A_270_53#_c_376_n N_A_270_53#_c_377_n
+ N_A_270_53#_c_378_n N_A_270_53#_c_379_n N_A_270_53#_c_389_n
+ N_A_270_53#_c_390_n N_A_270_53#_c_391_n N_A_270_53#_c_380_n
+ N_A_270_53#_c_381_n N_A_270_53#_c_457_p N_A_270_53#_c_382_n
+ N_A_270_53#_c_383_n PM_SKY130_FD_SC_LP__OR4BB_4%A_270_53#
x_PM_SKY130_FD_SC_LP__OR4BB_4%D_N N_D_N_M1012_g N_D_N_M1008_g D_N D_N
+ N_D_N_c_525_n N_D_N_c_526_n PM_SKY130_FD_SC_LP__OR4BB_4%D_N
x_PM_SKY130_FD_SC_LP__OR4BB_4%VPWR N_VPWR_M1014_d N_VPWR_M1000_d N_VPWR_M1005_d
+ N_VPWR_M1019_d N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n
+ N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n
+ VPWR N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_548_n N_VPWR_c_561_n
+ N_VPWR_c_562_n PM_SKY130_FD_SC_LP__OR4BB_4%VPWR
x_PM_SKY130_FD_SC_LP__OR4BB_4%X N_X_M1003_s N_X_M1016_s N_X_M1000_s N_X_M1010_s
+ N_X_c_624_n N_X_c_666_n N_X_c_626_n N_X_c_627_n N_X_c_670_n X X N_X_c_629_n X
+ PM_SKY130_FD_SC_LP__OR4BB_4%X
x_PM_SKY130_FD_SC_LP__OR4BB_4%VGND N_VGND_M1011_d N_VGND_M1015_d N_VGND_M1018_d
+ N_VGND_M1006_d N_VGND_M1017_d N_VGND_c_676_n N_VGND_c_677_n N_VGND_c_678_n
+ N_VGND_c_679_n N_VGND_c_680_n N_VGND_c_681_n N_VGND_c_682_n VGND
+ N_VGND_c_683_n N_VGND_c_684_n N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n
+ N_VGND_c_688_n N_VGND_c_689_n PM_SKY130_FD_SC_LP__OR4BB_4%VGND
cc_1 VNB N_C_N_c_104_n 0.0231062f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.215
cc_2 VNB N_C_N_M1014_g 0.00732341f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.045
cc_3 VNB N_C_N_c_106_n 0.0596018f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.38
cc_4 VNB N_C_N_c_107_n 0.0108499f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.38
cc_5 VNB C_N 0.0277344f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A_M1004_g 0.00473112f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.045
cc_7 VNB A 0.00626354f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.38
cc_8 VNB N_A_c_134_n 0.0313532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_135_n 0.019873f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_10 VNB N_B_M1015_g 0.0251017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_170_n 0.0242728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_c_171_n 0.00391033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_79_137#_M1007_g 0.0243414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_79_137#_c_208_n 0.00466358f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_15 VNB N_A_79_137#_c_209_n 0.00104374f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=1.665
cc_16 VNB N_A_79_137#_c_210_n 0.0259419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_79_137#_c_211_n 0.0129777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_528_27#_c_282_n 0.0180263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_528_27#_M1002_g 0.00593818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_528_27#_c_284_n 0.00429268f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_21 VNB N_A_528_27#_c_285_n 0.0474517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_528_27#_c_286_n 0.00377889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_528_27#_c_287_n 0.0188732f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=1.665
cc_24 VNB N_A_528_27#_c_288_n 0.0082772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_270_53#_M1003_g 0.0238339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_270_53#_M1006_g 0.023145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_270_53#_M1016_g 0.023118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_270_53#_M1017_g 0.0234027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_270_53#_c_375_n 0.00246282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_270_53#_c_376_n 0.00827321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_270_53#_c_377_n 0.00182398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_270_53#_c_378_n 0.00207996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_270_53#_c_379_n 0.00356289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_270_53#_c_380_n 0.00231453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_270_53#_c_381_n 8.18702e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_270_53#_c_382_n 0.00481694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_270_53#_c_383_n 0.0828377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_D_N_M1012_g 0.0334733f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.895
cc_39 VNB N_D_N_M1008_g 0.00193385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_D_N_c_525_n 0.121489f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_41 VNB N_D_N_c_526_n 0.0370865f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_42 VNB N_VPWR_c_548_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_624_n 0.00839522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB X 0.00476453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_676_n 0.0194268f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=1.295
cc_46 VNB N_VGND_c_677_n 0.00592932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_678_n 0.0187635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_679_n 0.0287009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_680_n 0.00615512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_681_n 0.0179887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_682_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_683_n 0.0184418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_684_n 0.0198281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_685_n 0.0275436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_686_n 0.360095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_687_n 0.0118081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_688_n 0.0117943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_689_n 0.0118439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_C_N_M1014_g 0.0315032f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.045
cc_60 VPB C_N 0.015078f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_61 VPB N_A_M1004_g 0.0219616f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.045
cc_62 VPB A 0.00308148f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.38
cc_63 VPB N_B_M1009_g 0.0189143f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=0.895
cc_64 VPB N_B_c_170_n 0.00635136f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_B_c_171_n 0.00312351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_79_137#_M1013_g 0.0197401f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.38
cc_67 VPB N_A_79_137#_c_208_n 0.00379278f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.38
cc_68 VPB N_A_79_137#_c_214_n 0.0137371f $X=-0.19 $Y=1.655 $X2=0.225 $Y2=1.295
cc_69 VPB N_A_79_137#_c_209_n 0.00104046f $X=-0.19 $Y=1.655 $X2=0.225 $Y2=1.665
cc_70 VPB N_A_79_137#_c_210_n 0.00836918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_528_27#_M1002_g 0.0247384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_528_27#_c_288_n 0.00384458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_528_27#_c_291_n 0.013184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_270_53#_M1000_g 0.0221988f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.38
cc_75 VPB N_A_270_53#_M1005_g 0.0187757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_270_53#_M1010_g 0.018749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_270_53#_M1019_g 0.0209949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_270_53#_c_379_n 9.47763e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_270_53#_c_389_n 0.0118115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_270_53#_c_390_n 0.0146711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_270_53#_c_391_n 0.00370501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_270_53#_c_381_n 0.0019314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A_270_53#_c_383_n 0.0141278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_D_N_M1008_g 0.031286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_D_N_c_526_n 0.0154136f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.38
cc_86 VPB N_VPWR_c_549_n 0.0318068f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.38
cc_87 VPB N_VPWR_c_550_n 0.0122412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_551_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_552_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_553_n 0.031426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_554_n 0.0613376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_555_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_556_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_557_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_558_n 0.030624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_559_n 0.0307831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_548_n 0.119204f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_561_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_562_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_X_c_626_n 0.00304538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_X_c_627_n 0.00220118f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB X 0.00122404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_X_c_629_n 0.00367691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 N_C_N_M1014_g N_A_M1004_g 0.0216928f $X=0.735 $Y=2.045 $X2=0 $Y2=0
cc_105 N_C_N_M1014_g A 0.00173431f $X=0.735 $Y=2.045 $X2=0 $Y2=0
cc_106 N_C_N_c_107_n A 0.00141897f $X=0.735 $Y=1.38 $X2=0 $Y2=0
cc_107 N_C_N_c_107_n N_A_c_134_n 0.0217256f $X=0.735 $Y=1.38 $X2=0 $Y2=0
cc_108 N_C_N_c_104_n N_A_c_135_n 0.0110383f $X=0.735 $Y=1.215 $X2=0 $Y2=0
cc_109 N_C_N_c_104_n N_A_79_137#_c_208_n 0.00572176f $X=0.735 $Y=1.215 $X2=0
+ $Y2=0
cc_110 N_C_N_M1014_g N_A_79_137#_c_208_n 0.0115643f $X=0.735 $Y=2.045 $X2=0
+ $Y2=0
cc_111 N_C_N_c_106_n N_A_79_137#_c_208_n 0.013446f $X=0.66 $Y=1.38 $X2=0 $Y2=0
cc_112 N_C_N_c_107_n N_A_79_137#_c_208_n 0.00481778f $X=0.735 $Y=1.38 $X2=0
+ $Y2=0
cc_113 C_N N_A_79_137#_c_208_n 0.0396922f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_114 N_C_N_M1014_g N_A_79_137#_c_222_n 0.0129262f $X=0.735 $Y=2.045 $X2=0
+ $Y2=0
cc_115 N_C_N_M1014_g N_A_79_137#_c_214_n 0.00509257f $X=0.735 $Y=2.045 $X2=0
+ $Y2=0
cc_116 N_C_N_c_106_n N_A_79_137#_c_214_n 0.00553104f $X=0.66 $Y=1.38 $X2=0 $Y2=0
cc_117 C_N N_A_79_137#_c_214_n 7.78181e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_118 N_C_N_c_104_n N_A_79_137#_c_211_n 0.00461409f $X=0.735 $Y=1.215 $X2=0
+ $Y2=0
cc_119 N_C_N_c_106_n N_A_79_137#_c_211_n 0.00752154f $X=0.66 $Y=1.38 $X2=0 $Y2=0
cc_120 C_N N_A_79_137#_c_211_n 7.78155e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_121 N_C_N_M1014_g N_VPWR_c_549_n 0.00329105f $X=0.735 $Y=2.045 $X2=0 $Y2=0
cc_122 N_C_N_c_104_n N_VGND_c_676_n 0.00565738f $X=0.735 $Y=1.215 $X2=0 $Y2=0
cc_123 N_C_N_c_104_n N_VGND_c_679_n 0.0036064f $X=0.735 $Y=1.215 $X2=0 $Y2=0
cc_124 N_C_N_c_104_n N_VGND_c_686_n 0.00453162f $X=0.735 $Y=1.215 $X2=0 $Y2=0
cc_125 N_A_M1004_g N_B_M1009_g 0.0679032f $X=1.275 $Y=2.465 $X2=0 $Y2=0
cc_126 A N_B_M1009_g 2.13565e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_127 A N_B_M1015_g 0.00268593f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_128 N_A_c_135_n N_B_M1015_g 0.0173582f $X=1.185 $Y=1.215 $X2=0 $Y2=0
cc_129 A N_B_c_170_n 0.00100169f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A_c_134_n N_B_c_170_n 0.0213463f $X=1.185 $Y=1.38 $X2=0 $Y2=0
cc_131 A N_B_c_171_n 0.0344293f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A_c_134_n N_B_c_171_n 0.00138391f $X=1.185 $Y=1.38 $X2=0 $Y2=0
cc_133 N_A_M1004_g N_A_79_137#_c_208_n 9.8122e-19 $X=1.275 $Y=2.465 $X2=0 $Y2=0
cc_134 A N_A_79_137#_c_208_n 0.0246512f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_135 N_A_c_134_n N_A_79_137#_c_208_n 9.85976e-19 $X=1.185 $Y=1.38 $X2=0 $Y2=0
cc_136 N_A_c_135_n N_A_79_137#_c_208_n 8.25264e-19 $X=1.185 $Y=1.215 $X2=0 $Y2=0
cc_137 N_A_M1004_g N_A_79_137#_c_222_n 0.0149226f $X=1.275 $Y=2.465 $X2=0 $Y2=0
cc_138 A N_A_79_137#_c_222_n 0.0239252f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A_c_134_n N_A_79_137#_c_222_n 6.89559e-19 $X=1.185 $Y=1.38 $X2=0 $Y2=0
cc_140 N_A_M1004_g N_A_79_137#_c_214_n 5.33613e-19 $X=1.275 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_c_135_n N_A_270_53#_c_375_n 8.16416e-19 $X=1.185 $Y=1.215 $X2=0 $Y2=0
cc_142 N_A_c_135_n N_A_270_53#_c_377_n 0.00324385f $X=1.185 $Y=1.215 $X2=0 $Y2=0
cc_143 N_A_M1004_g N_VPWR_c_549_n 0.0249555f $X=1.275 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_M1004_g N_VPWR_c_554_n 0.00486043f $X=1.275 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1004_g N_VPWR_c_548_n 0.00843372f $X=1.275 $Y=2.465 $X2=0 $Y2=0
cc_146 A N_VGND_c_676_n 0.0133392f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A_c_134_n N_VGND_c_676_n 0.00119676f $X=1.185 $Y=1.38 $X2=0 $Y2=0
cc_148 N_A_c_135_n N_VGND_c_676_n 0.00624086f $X=1.185 $Y=1.215 $X2=0 $Y2=0
cc_149 N_A_c_135_n N_VGND_c_681_n 0.00555245f $X=1.185 $Y=1.215 $X2=0 $Y2=0
cc_150 N_A_c_135_n N_VGND_c_686_n 0.0116312f $X=1.185 $Y=1.215 $X2=0 $Y2=0
cc_151 N_B_M1009_g N_A_79_137#_M1013_g 0.0707682f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_152 N_B_c_171_n N_A_79_137#_M1013_g 4.94547e-19 $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_153 N_B_M1015_g N_A_79_137#_M1007_g 0.0182471f $X=1.765 $Y=0.685 $X2=0 $Y2=0
cc_154 N_B_M1009_g N_A_79_137#_c_222_n 0.0152054f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_155 N_B_c_170_n N_A_79_137#_c_222_n 8.05279e-19 $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_156 N_B_c_171_n N_A_79_137#_c_222_n 0.0237784f $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_157 N_B_M1009_g N_A_79_137#_c_209_n 0.0011385f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B_c_170_n N_A_79_137#_c_209_n 0.00115083f $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_159 N_B_c_171_n N_A_79_137#_c_209_n 0.0259542f $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_160 N_B_c_170_n N_A_79_137#_c_210_n 0.0201104f $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_161 N_B_c_171_n N_A_79_137#_c_210_n 0.00114883f $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_162 N_B_M1015_g N_A_270_53#_c_375_n 0.0100751f $X=1.765 $Y=0.685 $X2=0 $Y2=0
cc_163 N_B_M1015_g N_A_270_53#_c_376_n 0.0131066f $X=1.765 $Y=0.685 $X2=0 $Y2=0
cc_164 N_B_c_170_n N_A_270_53#_c_376_n 3.41152e-19 $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_165 N_B_c_171_n N_A_270_53#_c_376_n 0.0136861f $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_166 N_B_M1015_g N_A_270_53#_c_377_n 6.81087e-19 $X=1.765 $Y=0.685 $X2=0 $Y2=0
cc_167 N_B_c_170_n N_A_270_53#_c_377_n 0.00101761f $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_168 N_B_c_171_n N_A_270_53#_c_377_n 0.0140434f $X=1.725 $Y=1.51 $X2=0 $Y2=0
cc_169 N_B_M1009_g N_VPWR_c_549_n 0.00501578f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_170 N_B_M1009_g N_VPWR_c_554_n 0.00585385f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_171 N_B_M1009_g N_VPWR_c_548_n 0.0111381f $X=1.725 $Y=2.465 $X2=0 $Y2=0
cc_172 N_B_M1015_g N_VGND_c_677_n 0.00177056f $X=1.765 $Y=0.685 $X2=0 $Y2=0
cc_173 N_B_M1015_g N_VGND_c_681_n 0.00549455f $X=1.765 $Y=0.685 $X2=0 $Y2=0
cc_174 N_B_M1015_g N_VGND_c_686_n 0.0105936f $X=1.765 $Y=0.685 $X2=0 $Y2=0
cc_175 N_A_79_137#_M1007_g N_A_528_27#_c_282_n 0.0223418f $X=2.285 $Y=0.685
+ $X2=0 $Y2=0
cc_176 N_A_79_137#_M1013_g N_A_528_27#_M1002_g 0.0486902f $X=2.175 $Y=2.465
+ $X2=0 $Y2=0
cc_177 N_A_79_137#_c_222_n N_A_528_27#_M1002_g 0.00152664f $X=2.1 $Y=2.01 $X2=0
+ $Y2=0
cc_178 N_A_79_137#_c_209_n N_A_528_27#_M1002_g 7.06281e-19 $X=2.265 $Y=1.51
+ $X2=0 $Y2=0
cc_179 N_A_79_137#_c_209_n N_A_528_27#_c_285_n 2.96168e-19 $X=2.265 $Y=1.51
+ $X2=0 $Y2=0
cc_180 N_A_79_137#_c_210_n N_A_528_27#_c_285_n 0.0204065f $X=2.265 $Y=1.51 $X2=0
+ $Y2=0
cc_181 N_A_79_137#_M1007_g N_A_270_53#_c_375_n 4.10624e-19 $X=2.285 $Y=0.685
+ $X2=0 $Y2=0
cc_182 N_A_79_137#_M1007_g N_A_270_53#_c_376_n 0.0144791f $X=2.285 $Y=0.685
+ $X2=0 $Y2=0
cc_183 N_A_79_137#_c_209_n N_A_270_53#_c_376_n 0.0184514f $X=2.265 $Y=1.51 $X2=0
+ $Y2=0
cc_184 N_A_79_137#_c_210_n N_A_270_53#_c_376_n 9.17626e-19 $X=2.265 $Y=1.51
+ $X2=0 $Y2=0
cc_185 N_A_79_137#_M1007_g N_A_270_53#_c_378_n 7.80435e-19 $X=2.285 $Y=0.685
+ $X2=0 $Y2=0
cc_186 N_A_79_137#_M1013_g N_A_270_53#_c_379_n 2.1886e-19 $X=2.175 $Y=2.465
+ $X2=0 $Y2=0
cc_187 N_A_79_137#_M1007_g N_A_270_53#_c_379_n 0.0037016f $X=2.285 $Y=0.685
+ $X2=0 $Y2=0
cc_188 N_A_79_137#_c_209_n N_A_270_53#_c_379_n 0.0292202f $X=2.265 $Y=1.51 $X2=0
+ $Y2=0
cc_189 N_A_79_137#_c_210_n N_A_270_53#_c_379_n 0.00204951f $X=2.265 $Y=1.51
+ $X2=0 $Y2=0
cc_190 N_A_79_137#_M1013_g N_A_270_53#_c_389_n 0.00470233f $X=2.175 $Y=2.465
+ $X2=0 $Y2=0
cc_191 N_A_79_137#_c_222_n N_A_270_53#_c_389_n 0.00705146f $X=2.1 $Y=2.01 $X2=0
+ $Y2=0
cc_192 N_A_79_137#_M1013_g N_A_270_53#_c_391_n 5.84103e-19 $X=2.175 $Y=2.465
+ $X2=0 $Y2=0
cc_193 N_A_79_137#_c_209_n N_A_270_53#_c_391_n 0.0137017f $X=2.265 $Y=1.51 $X2=0
+ $Y2=0
cc_194 N_A_79_137#_c_210_n N_A_270_53#_c_382_n 0.00285766f $X=2.265 $Y=1.51
+ $X2=0 $Y2=0
cc_195 N_A_79_137#_c_222_n N_VPWR_M1014_d 0.0109923f $X=2.1 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_79_137#_c_222_n N_VPWR_c_549_n 0.0219507f $X=2.1 $Y=2.01 $X2=0 $Y2=0
cc_197 N_A_79_137#_M1013_g N_VPWR_c_554_n 0.00585385f $X=2.175 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A_79_137#_M1013_g N_VPWR_c_548_n 0.0113476f $X=2.175 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A_79_137#_c_222_n A_270_367# 0.0122827f $X=2.1 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A_79_137#_c_222_n A_360_367# 0.0132482f $X=2.1 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_201 N_A_79_137#_c_222_n A_450_367# 0.00416623f $X=2.1 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A_79_137#_c_209_n A_450_367# 8.04744e-19 $X=2.265 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_203 N_A_79_137#_c_211_n N_VGND_c_676_n 0.0240761f $X=0.62 $Y=0.885 $X2=0
+ $Y2=0
cc_204 N_A_79_137#_M1007_g N_VGND_c_677_n 0.00309326f $X=2.285 $Y=0.685 $X2=0
+ $Y2=0
cc_205 N_A_79_137#_c_211_n N_VGND_c_679_n 0.00478516f $X=0.62 $Y=0.885 $X2=0
+ $Y2=0
cc_206 N_A_79_137#_M1007_g N_VGND_c_683_n 0.00555245f $X=2.285 $Y=0.685 $X2=0
+ $Y2=0
cc_207 N_A_79_137#_M1007_g N_VGND_c_686_n 0.010634f $X=2.285 $Y=0.685 $X2=0
+ $Y2=0
cc_208 N_A_79_137#_c_211_n N_VGND_c_686_n 0.0094663f $X=0.62 $Y=0.885 $X2=0
+ $Y2=0
cc_209 N_A_528_27#_c_282_n N_A_270_53#_M1003_g 0.0166678f $X=2.715 $Y=1.215
+ $X2=0 $Y2=0
cc_210 N_A_528_27#_c_284_n N_A_270_53#_M1003_g 0.00886843f $X=2.965 $Y=1.38
+ $X2=0 $Y2=0
cc_211 N_A_528_27#_c_285_n N_A_270_53#_M1003_g 0.0169791f $X=2.965 $Y=1.38 $X2=0
+ $Y2=0
cc_212 N_A_528_27#_c_286_n N_A_270_53#_M1003_g 0.0140569f $X=5.51 $Y=0.64 $X2=0
+ $Y2=0
cc_213 N_A_528_27#_c_286_n N_A_270_53#_M1006_g 0.0120795f $X=5.51 $Y=0.64 $X2=0
+ $Y2=0
cc_214 N_A_528_27#_c_286_n N_A_270_53#_M1016_g 0.0120795f $X=5.51 $Y=0.64 $X2=0
+ $Y2=0
cc_215 N_A_528_27#_c_286_n N_A_270_53#_M1017_g 0.0124249f $X=5.51 $Y=0.64 $X2=0
+ $Y2=0
cc_216 N_A_528_27#_c_287_n N_A_270_53#_M1017_g 7.54342e-19 $X=5.607 $Y=0.725
+ $X2=0 $Y2=0
cc_217 N_A_528_27#_c_288_n N_A_270_53#_M1017_g 0.00122807f $X=5.607 $Y=1.92
+ $X2=0 $Y2=0
cc_218 N_A_528_27#_c_291_n N_A_270_53#_M1019_g 2.65393e-19 $X=5.7 $Y=2.045 $X2=0
+ $Y2=0
cc_219 N_A_528_27#_c_282_n N_A_270_53#_c_378_n 0.0135959f $X=2.715 $Y=1.215
+ $X2=0 $Y2=0
cc_220 N_A_528_27#_c_284_n N_A_270_53#_c_378_n 0.020527f $X=2.965 $Y=1.38 $X2=0
+ $Y2=0
cc_221 N_A_528_27#_c_310_p N_A_270_53#_c_378_n 0.0140532f $X=3.13 $Y=0.64 $X2=0
+ $Y2=0
cc_222 N_A_528_27#_c_282_n N_A_270_53#_c_379_n 9.24074e-19 $X=2.715 $Y=1.215
+ $X2=0 $Y2=0
cc_223 N_A_528_27#_M1002_g N_A_270_53#_c_379_n 0.0062548f $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_224 N_A_528_27#_c_284_n N_A_270_53#_c_379_n 0.0267553f $X=2.965 $Y=1.38 $X2=0
+ $Y2=0
cc_225 N_A_528_27#_c_285_n N_A_270_53#_c_379_n 0.00797219f $X=2.965 $Y=1.38
+ $X2=0 $Y2=0
cc_226 N_A_528_27#_M1002_g N_A_270_53#_c_389_n 0.0254979f $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_227 N_A_528_27#_M1002_g N_A_270_53#_c_391_n 0.0155582f $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_228 N_A_528_27#_c_284_n N_A_270_53#_c_391_n 0.017537f $X=2.965 $Y=1.38 $X2=0
+ $Y2=0
cc_229 N_A_528_27#_c_285_n N_A_270_53#_c_391_n 0.00465084f $X=2.965 $Y=1.38
+ $X2=0 $Y2=0
cc_230 N_A_528_27#_M1002_g N_A_270_53#_c_380_n 2.51568e-19 $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_231 N_A_528_27#_c_284_n N_A_270_53#_c_380_n 0.0182558f $X=2.965 $Y=1.38 $X2=0
+ $Y2=0
cc_232 N_A_528_27#_c_285_n N_A_270_53#_c_380_n 0.00144391f $X=2.965 $Y=1.38
+ $X2=0 $Y2=0
cc_233 N_A_528_27#_c_286_n N_A_270_53#_c_380_n 0.0040696f $X=5.51 $Y=0.64 $X2=0
+ $Y2=0
cc_234 N_A_528_27#_M1002_g N_A_270_53#_c_381_n 0.0021579f $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_235 N_A_528_27#_c_282_n N_A_270_53#_c_382_n 0.00287784f $X=2.715 $Y=1.215
+ $X2=0 $Y2=0
cc_236 N_A_528_27#_c_284_n N_A_270_53#_c_382_n 0.0138549f $X=2.965 $Y=1.38 $X2=0
+ $Y2=0
cc_237 N_A_528_27#_M1002_g N_A_270_53#_c_383_n 0.00163722f $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_238 N_A_528_27#_c_284_n N_A_270_53#_c_383_n 2.47891e-19 $X=2.965 $Y=1.38
+ $X2=0 $Y2=0
cc_239 N_A_528_27#_c_285_n N_A_270_53#_c_383_n 0.00381165f $X=2.965 $Y=1.38
+ $X2=0 $Y2=0
cc_240 N_A_528_27#_c_288_n N_A_270_53#_c_383_n 2.07267e-19 $X=5.607 $Y=1.92
+ $X2=0 $Y2=0
cc_241 N_A_528_27#_c_286_n N_D_N_M1012_g 0.0109147f $X=5.51 $Y=0.64 $X2=0 $Y2=0
cc_242 N_A_528_27#_c_287_n N_D_N_M1012_g 0.00719478f $X=5.607 $Y=0.725 $X2=0
+ $Y2=0
cc_243 N_A_528_27#_c_288_n N_D_N_M1012_g 0.00861422f $X=5.607 $Y=1.92 $X2=0
+ $Y2=0
cc_244 N_A_528_27#_c_288_n N_D_N_M1008_g 0.00849301f $X=5.607 $Y=1.92 $X2=0
+ $Y2=0
cc_245 N_A_528_27#_c_291_n N_D_N_M1008_g 0.00719811f $X=5.7 $Y=2.045 $X2=0 $Y2=0
cc_246 N_A_528_27#_c_287_n N_D_N_c_525_n 0.00668076f $X=5.607 $Y=0.725 $X2=0
+ $Y2=0
cc_247 N_A_528_27#_c_288_n N_D_N_c_525_n 0.0345929f $X=5.607 $Y=1.92 $X2=0 $Y2=0
cc_248 N_A_528_27#_c_291_n N_D_N_c_525_n 0.00659753f $X=5.7 $Y=2.045 $X2=0 $Y2=0
cc_249 N_A_528_27#_c_288_n N_D_N_c_526_n 0.0575874f $X=5.607 $Y=1.92 $X2=0 $Y2=0
cc_250 N_A_528_27#_M1002_g N_VPWR_c_550_n 0.00417735f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_251 N_A_528_27#_c_291_n N_VPWR_c_553_n 0.00972606f $X=5.7 $Y=2.045 $X2=0
+ $Y2=0
cc_252 N_A_528_27#_M1002_g N_VPWR_c_554_n 0.0054895f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_253 N_A_528_27#_M1002_g N_VPWR_c_548_n 0.0116084f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_254 N_A_528_27#_c_286_n N_X_M1003_s 0.00429347f $X=5.51 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_255 N_A_528_27#_c_286_n N_X_M1016_s 0.00429347f $X=5.51 $Y=0.64 $X2=0 $Y2=0
cc_256 N_A_528_27#_c_284_n N_X_c_624_n 0.0119537f $X=2.965 $Y=1.38 $X2=0 $Y2=0
cc_257 N_A_528_27#_c_286_n N_X_c_624_n 0.101088f $X=5.51 $Y=0.64 $X2=0 $Y2=0
cc_258 N_A_528_27#_c_288_n N_X_c_624_n 0.0134498f $X=5.607 $Y=1.92 $X2=0 $Y2=0
cc_259 N_A_528_27#_c_288_n X 0.0311556f $X=5.607 $Y=1.92 $X2=0 $Y2=0
cc_260 N_A_528_27#_c_288_n N_X_c_629_n 0.00916931f $X=5.607 $Y=1.92 $X2=0 $Y2=0
cc_261 N_A_528_27#_c_284_n N_VGND_M1018_d 0.0119025f $X=2.965 $Y=1.38 $X2=0
+ $Y2=0
cc_262 N_A_528_27#_c_286_n N_VGND_M1018_d 0.00800263f $X=5.51 $Y=0.64 $X2=0
+ $Y2=0
cc_263 N_A_528_27#_c_310_p N_VGND_M1018_d 0.0065744f $X=3.13 $Y=0.64 $X2=0 $Y2=0
cc_264 N_A_528_27#_c_286_n N_VGND_M1006_d 0.00608986f $X=5.51 $Y=0.64 $X2=0
+ $Y2=0
cc_265 N_A_528_27#_c_286_n N_VGND_M1017_d 0.011438f $X=5.51 $Y=0.64 $X2=0 $Y2=0
cc_266 N_A_528_27#_c_286_n N_VGND_c_678_n 0.0126366f $X=5.51 $Y=0.64 $X2=0 $Y2=0
cc_267 N_A_528_27#_c_282_n N_VGND_c_683_n 0.00469843f $X=2.715 $Y=1.215 $X2=0
+ $Y2=0
cc_268 N_A_528_27#_c_310_p N_VGND_c_683_n 2.31449e-19 $X=3.13 $Y=0.64 $X2=0
+ $Y2=0
cc_269 N_A_528_27#_c_286_n N_VGND_c_684_n 0.013478f $X=5.51 $Y=0.64 $X2=0 $Y2=0
cc_270 N_A_528_27#_c_286_n N_VGND_c_685_n 0.00336185f $X=5.51 $Y=0.64 $X2=0
+ $Y2=0
cc_271 N_A_528_27#_c_287_n N_VGND_c_685_n 0.0159086f $X=5.607 $Y=0.725 $X2=0
+ $Y2=0
cc_272 N_A_528_27#_c_282_n N_VGND_c_686_n 0.00892035f $X=2.715 $Y=1.215 $X2=0
+ $Y2=0
cc_273 N_A_528_27#_c_286_n N_VGND_c_686_n 0.0504225f $X=5.51 $Y=0.64 $X2=0 $Y2=0
cc_274 N_A_528_27#_c_310_p N_VGND_c_686_n 0.0018498f $X=3.13 $Y=0.64 $X2=0 $Y2=0
cc_275 N_A_528_27#_c_287_n N_VGND_c_686_n 0.0129267f $X=5.607 $Y=0.725 $X2=0
+ $Y2=0
cc_276 N_A_528_27#_c_282_n N_VGND_c_687_n 0.00411335f $X=2.715 $Y=1.215 $X2=0
+ $Y2=0
cc_277 N_A_528_27#_c_286_n N_VGND_c_687_n 0.00582708f $X=5.51 $Y=0.64 $X2=0
+ $Y2=0
cc_278 N_A_528_27#_c_310_p N_VGND_c_687_n 0.0203865f $X=3.13 $Y=0.64 $X2=0 $Y2=0
cc_279 N_A_528_27#_c_286_n N_VGND_c_688_n 0.0212102f $X=5.51 $Y=0.64 $X2=0 $Y2=0
cc_280 N_A_528_27#_c_286_n N_VGND_c_689_n 0.024325f $X=5.51 $Y=0.64 $X2=0 $Y2=0
cc_281 N_A_528_27#_c_287_n N_VGND_c_689_n 0.00487979f $X=5.607 $Y=0.725 $X2=0
+ $Y2=0
cc_282 N_A_270_53#_M1017_g N_D_N_M1012_g 0.0137048f $X=4.825 $Y=0.685 $X2=0
+ $Y2=0
cc_283 N_A_270_53#_M1019_g N_D_N_M1008_g 0.00915135f $X=4.96 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_A_270_53#_c_383_n N_D_N_c_525_n 0.0228561f $X=4.825 $Y=1.49 $X2=0 $Y2=0
cc_285 N_A_270_53#_c_390_n N_VPWR_M1000_d 0.00326164f $X=3.3 $Y=1.84 $X2=0 $Y2=0
cc_286 N_A_270_53#_M1000_g N_VPWR_c_550_n 0.0155684f $X=3.67 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_A_270_53#_M1005_g N_VPWR_c_550_n 7.27171e-19 $X=4.1 $Y=2.465 $X2=0
+ $Y2=0
cc_288 N_A_270_53#_c_389_n N_VPWR_c_550_n 0.0741033f $X=2.93 $Y=1.98 $X2=0 $Y2=0
cc_289 N_A_270_53#_c_390_n N_VPWR_c_550_n 0.0220423f $X=3.3 $Y=1.84 $X2=0 $Y2=0
cc_290 N_A_270_53#_c_457_p N_VPWR_c_550_n 0.00151356f $X=4.555 $Y=1.49 $X2=0
+ $Y2=0
cc_291 N_A_270_53#_c_383_n N_VPWR_c_550_n 8.24241e-19 $X=4.825 $Y=1.49 $X2=0
+ $Y2=0
cc_292 N_A_270_53#_M1000_g N_VPWR_c_551_n 7.3e-19 $X=3.67 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A_270_53#_M1005_g N_VPWR_c_551_n 0.0143802f $X=4.1 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A_270_53#_M1010_g N_VPWR_c_551_n 0.0143802f $X=4.53 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_270_53#_M1019_g N_VPWR_c_551_n 7.3e-19 $X=4.96 $Y=2.465 $X2=0 $Y2=0
cc_296 N_A_270_53#_M1010_g N_VPWR_c_552_n 0.00486043f $X=4.53 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_A_270_53#_M1019_g N_VPWR_c_552_n 0.00486043f $X=4.96 $Y=2.465 $X2=0
+ $Y2=0
cc_298 N_A_270_53#_M1010_g N_VPWR_c_553_n 7.3e-19 $X=4.53 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A_270_53#_M1019_g N_VPWR_c_553_n 0.0154849f $X=4.96 $Y=2.465 $X2=0
+ $Y2=0
cc_300 N_A_270_53#_c_389_n N_VPWR_c_554_n 0.0210467f $X=2.93 $Y=1.98 $X2=0 $Y2=0
cc_301 N_A_270_53#_M1000_g N_VPWR_c_556_n 0.00486043f $X=3.67 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_A_270_53#_M1005_g N_VPWR_c_556_n 0.00486043f $X=4.1 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_270_53#_M1002_d N_VPWR_c_548_n 0.00215158f $X=2.79 $Y=1.835 $X2=0
+ $Y2=0
cc_304 N_A_270_53#_M1000_g N_VPWR_c_548_n 0.00824727f $X=3.67 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_A_270_53#_M1005_g N_VPWR_c_548_n 0.00824727f $X=4.1 $Y=2.465 $X2=0
+ $Y2=0
cc_306 N_A_270_53#_M1010_g N_VPWR_c_548_n 0.00824727f $X=4.53 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_270_53#_M1019_g N_VPWR_c_548_n 0.00824727f $X=4.96 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A_270_53#_c_389_n N_VPWR_c_548_n 0.0125689f $X=2.93 $Y=1.98 $X2=0 $Y2=0
cc_309 N_A_270_53#_c_391_n A_450_367# 0.00284854f $X=3.095 $Y=1.84 $X2=-0.19
+ $Y2=-0.245
cc_310 N_A_270_53#_M1003_g N_X_c_624_n 0.00474137f $X=3.415 $Y=0.685 $X2=0 $Y2=0
cc_311 N_A_270_53#_M1006_g N_X_c_624_n 0.012057f $X=3.845 $Y=0.685 $X2=0 $Y2=0
cc_312 N_A_270_53#_M1016_g N_X_c_624_n 0.012057f $X=4.395 $Y=0.685 $X2=0 $Y2=0
cc_313 N_A_270_53#_M1017_g N_X_c_624_n 0.0133686f $X=4.825 $Y=0.685 $X2=0 $Y2=0
cc_314 N_A_270_53#_c_380_n N_X_c_624_n 0.00574734f $X=3.42 $Y=1.575 $X2=0 $Y2=0
cc_315 N_A_270_53#_c_457_p N_X_c_624_n 0.0845372f $X=4.555 $Y=1.49 $X2=0 $Y2=0
cc_316 N_A_270_53#_c_383_n N_X_c_624_n 0.0110232f $X=4.825 $Y=1.49 $X2=0 $Y2=0
cc_317 N_A_270_53#_M1005_g N_X_c_626_n 0.0130971f $X=4.1 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A_270_53#_M1010_g N_X_c_626_n 0.0132616f $X=4.53 $Y=2.465 $X2=0 $Y2=0
cc_319 N_A_270_53#_c_457_p N_X_c_626_n 0.053265f $X=4.555 $Y=1.49 $X2=0 $Y2=0
cc_320 N_A_270_53#_c_383_n N_X_c_626_n 0.00289453f $X=4.825 $Y=1.49 $X2=0 $Y2=0
cc_321 N_A_270_53#_M1000_g N_X_c_627_n 8.83463e-19 $X=3.67 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A_270_53#_c_390_n N_X_c_627_n 0.00563246f $X=3.3 $Y=1.84 $X2=0 $Y2=0
cc_323 N_A_270_53#_c_381_n N_X_c_627_n 6.28717e-19 $X=3.42 $Y=1.755 $X2=0 $Y2=0
cc_324 N_A_270_53#_c_457_p N_X_c_627_n 0.0157258f $X=4.555 $Y=1.49 $X2=0 $Y2=0
cc_325 N_A_270_53#_c_383_n N_X_c_627_n 0.00299787f $X=4.825 $Y=1.49 $X2=0 $Y2=0
cc_326 N_A_270_53#_M1016_g X 8.46089e-19 $X=4.395 $Y=0.685 $X2=0 $Y2=0
cc_327 N_A_270_53#_M1010_g X 5.51633e-19 $X=4.53 $Y=2.465 $X2=0 $Y2=0
cc_328 N_A_270_53#_M1017_g X 0.00575239f $X=4.825 $Y=0.685 $X2=0 $Y2=0
cc_329 N_A_270_53#_M1019_g X 0.00381912f $X=4.96 $Y=2.465 $X2=0 $Y2=0
cc_330 N_A_270_53#_c_457_p X 0.0198181f $X=4.555 $Y=1.49 $X2=0 $Y2=0
cc_331 N_A_270_53#_c_383_n X 0.0169561f $X=4.825 $Y=1.49 $X2=0 $Y2=0
cc_332 N_A_270_53#_M1019_g N_X_c_629_n 0.0116016f $X=4.96 $Y=2.465 $X2=0 $Y2=0
cc_333 N_A_270_53#_c_383_n N_X_c_629_n 0.00327074f $X=4.825 $Y=1.49 $X2=0 $Y2=0
cc_334 N_A_270_53#_c_376_n N_VGND_M1015_d 0.00284774f $X=2.365 $Y=1.08 $X2=0
+ $Y2=0
cc_335 N_A_270_53#_c_375_n N_VGND_c_676_n 7.47134e-19 $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_336 N_A_270_53#_c_375_n N_VGND_c_677_n 0.021387f $X=1.525 $Y=0.42 $X2=0 $Y2=0
cc_337 N_A_270_53#_c_376_n N_VGND_c_677_n 0.0199561f $X=2.365 $Y=1.08 $X2=0
+ $Y2=0
cc_338 N_A_270_53#_c_378_n N_VGND_c_677_n 7.49726e-19 $X=2.5 $Y=0.42 $X2=0 $Y2=0
cc_339 N_A_270_53#_M1016_g N_VGND_c_678_n 0.00389194f $X=4.395 $Y=0.685 $X2=0
+ $Y2=0
cc_340 N_A_270_53#_M1017_g N_VGND_c_678_n 0.00389194f $X=4.825 $Y=0.685 $X2=0
+ $Y2=0
cc_341 N_A_270_53#_c_375_n N_VGND_c_681_n 0.0234992f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_342 N_A_270_53#_c_378_n N_VGND_c_683_n 0.0236643f $X=2.5 $Y=0.42 $X2=0 $Y2=0
cc_343 N_A_270_53#_M1003_g N_VGND_c_684_n 0.00389194f $X=3.415 $Y=0.685 $X2=0
+ $Y2=0
cc_344 N_A_270_53#_M1006_g N_VGND_c_684_n 0.00389194f $X=3.845 $Y=0.685 $X2=0
+ $Y2=0
cc_345 N_A_270_53#_M1003_g N_VGND_c_686_n 0.00596709f $X=3.415 $Y=0.685 $X2=0
+ $Y2=0
cc_346 N_A_270_53#_M1006_g N_VGND_c_686_n 0.00556918f $X=3.845 $Y=0.685 $X2=0
+ $Y2=0
cc_347 N_A_270_53#_M1016_g N_VGND_c_686_n 0.00556918f $X=4.395 $Y=0.685 $X2=0
+ $Y2=0
cc_348 N_A_270_53#_M1017_g N_VGND_c_686_n 0.00589032f $X=4.825 $Y=0.685 $X2=0
+ $Y2=0
cc_349 N_A_270_53#_c_375_n N_VGND_c_686_n 0.0127336f $X=1.525 $Y=0.42 $X2=0
+ $Y2=0
cc_350 N_A_270_53#_c_378_n N_VGND_c_686_n 0.0126763f $X=2.5 $Y=0.42 $X2=0 $Y2=0
cc_351 N_A_270_53#_M1003_g N_VGND_c_687_n 0.00617284f $X=3.415 $Y=0.685 $X2=0
+ $Y2=0
cc_352 N_A_270_53#_c_378_n N_VGND_c_687_n 0.00968174f $X=2.5 $Y=0.42 $X2=0 $Y2=0
cc_353 N_A_270_53#_M1006_g N_VGND_c_688_n 0.0039161f $X=3.845 $Y=0.685 $X2=0
+ $Y2=0
cc_354 N_A_270_53#_M1016_g N_VGND_c_688_n 0.0039161f $X=4.395 $Y=0.685 $X2=0
+ $Y2=0
cc_355 N_A_270_53#_M1017_g N_VGND_c_689_n 0.00647286f $X=4.825 $Y=0.685 $X2=0
+ $Y2=0
cc_356 N_D_N_M1008_g N_VPWR_c_553_n 0.00592692f $X=5.485 $Y=2.045 $X2=0 $Y2=0
cc_357 N_D_N_M1012_g N_X_c_624_n 0.00298315f $X=5.485 $Y=0.475 $X2=0 $Y2=0
cc_358 N_D_N_c_525_n X 0.00639657f $X=5.97 $Y=1.12 $X2=0 $Y2=0
cc_359 N_D_N_M1008_g N_X_c_629_n 0.0015017f $X=5.485 $Y=2.045 $X2=0 $Y2=0
cc_360 N_D_N_M1012_g N_VGND_c_685_n 0.00382387f $X=5.485 $Y=0.475 $X2=0 $Y2=0
cc_361 N_D_N_M1012_g N_VGND_c_686_n 0.00676457f $X=5.485 $Y=0.475 $X2=0 $Y2=0
cc_362 N_D_N_M1012_g N_VGND_c_689_n 0.00509838f $X=5.485 $Y=0.475 $X2=0 $Y2=0
cc_363 N_VPWR_c_548_n A_270_367# 0.0128488f $X=6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_364 N_VPWR_c_548_n A_360_367# 0.0128488f $X=6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_365 N_VPWR_c_548_n A_450_367# 0.0167135f $X=6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_366 N_VPWR_c_548_n N_X_M1000_s 0.00536646f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_367 N_VPWR_c_548_n N_X_M1010_s 0.00536646f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_368 N_VPWR_c_556_n N_X_c_666_n 0.0124525f $X=4.15 $Y=3.33 $X2=0 $Y2=0
cc_369 N_VPWR_c_548_n N_X_c_666_n 0.00730901f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_370 N_VPWR_M1005_d N_X_c_626_n 0.00176461f $X=4.175 $Y=1.835 $X2=0 $Y2=0
cc_371 N_VPWR_c_551_n N_X_c_626_n 0.0170777f $X=4.315 $Y=2.17 $X2=0 $Y2=0
cc_372 N_VPWR_c_552_n N_X_c_670_n 0.0124525f $X=5.01 $Y=3.33 $X2=0 $Y2=0
cc_373 N_VPWR_c_548_n N_X_c_670_n 0.00730901f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_374 N_VPWR_M1019_d N_X_c_629_n 0.00231219f $X=5.035 $Y=1.835 $X2=0 $Y2=0
cc_375 N_VPWR_c_553_n N_X_c_629_n 0.0126068f $X=5.175 $Y=2.17 $X2=0 $Y2=0
cc_376 N_X_c_624_n N_VGND_M1006_d 0.00354682f $X=4.89 $Y=1.02 $X2=0 $Y2=0
cc_377 N_X_c_624_n N_VGND_M1017_d 0.00693031f $X=4.89 $Y=1.02 $X2=0 $Y2=0
