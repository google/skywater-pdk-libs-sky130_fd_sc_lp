* File: sky130_fd_sc_lp__einvn_4.pxi.spice
* Created: Wed Sep  2 09:51:46 2020
* 
x_PM_SKY130_FD_SC_LP__EINVN_4%A N_A_c_109_n N_A_M1002_g N_A_M1000_g N_A_c_110_n
+ N_A_M1003_g N_A_M1001_g N_A_M1004_g N_A_M1010_g N_A_c_112_n N_A_c_113_n
+ N_A_M1009_g N_A_M1013_g N_A_c_115_n A A A A PM_SKY130_FD_SC_LP__EINVN_4%A
x_PM_SKY130_FD_SC_LP__EINVN_4%A_555_201# N_A_555_201#_M1016_d
+ N_A_555_201#_M1011_d N_A_555_201#_c_201_n N_A_555_201#_c_202_n
+ N_A_555_201#_M1007_g N_A_555_201#_c_203_n N_A_555_201#_c_204_n
+ N_A_555_201#_M1008_g N_A_555_201#_c_205_n N_A_555_201#_c_206_n
+ N_A_555_201#_M1012_g N_A_555_201#_c_207_n N_A_555_201#_c_208_n
+ N_A_555_201#_M1014_g N_A_555_201#_c_209_n N_A_555_201#_c_210_n
+ N_A_555_201#_c_211_n N_A_555_201#_c_212_n N_A_555_201#_c_213_n
+ N_A_555_201#_c_214_n N_A_555_201#_c_215_n N_A_555_201#_c_216_n
+ N_A_555_201#_c_217_n PM_SKY130_FD_SC_LP__EINVN_4%A_555_201#
x_PM_SKY130_FD_SC_LP__EINVN_4%TE_B N_TE_B_c_311_n N_TE_B_M1005_g N_TE_B_c_299_n
+ N_TE_B_c_300_n N_TE_B_c_314_n N_TE_B_M1006_g N_TE_B_c_301_n N_TE_B_c_316_n
+ N_TE_B_M1015_g N_TE_B_c_302_n N_TE_B_c_318_n N_TE_B_M1017_g N_TE_B_c_303_n
+ N_TE_B_c_304_n N_TE_B_M1016_g N_TE_B_c_321_n N_TE_B_M1011_g N_TE_B_c_306_n
+ N_TE_B_c_307_n N_TE_B_c_308_n N_TE_B_c_309_n N_TE_B_c_310_n TE_B TE_B TE_B
+ N_TE_B_c_327_n N_TE_B_c_328_n PM_SKY130_FD_SC_LP__EINVN_4%TE_B
x_PM_SKY130_FD_SC_LP__EINVN_4%A_87_367# N_A_87_367#_M1000_s N_A_87_367#_M1001_s
+ N_A_87_367#_M1013_s N_A_87_367#_M1006_s N_A_87_367#_M1017_s
+ N_A_87_367#_c_389_n N_A_87_367#_c_390_n N_A_87_367#_c_397_n
+ N_A_87_367#_c_399_n N_A_87_367#_c_401_n N_A_87_367#_c_438_p
+ N_A_87_367#_c_391_n N_A_87_367#_c_392_n N_A_87_367#_c_432_p
+ N_A_87_367#_c_393_n N_A_87_367#_c_394_n N_A_87_367#_c_404_n
+ N_A_87_367#_c_395_n PM_SKY130_FD_SC_LP__EINVN_4%A_87_367#
x_PM_SKY130_FD_SC_LP__EINVN_4%Z N_Z_M1002_d N_Z_M1004_d N_Z_M1000_d N_Z_M1010_d
+ N_Z_c_459_n N_Z_c_460_n N_Z_c_455_n N_Z_c_456_n N_Z_c_469_n N_Z_c_473_n
+ N_Z_c_476_n N_Z_c_457_n N_Z_c_458_n N_Z_c_487_n Z Z N_Z_c_489_n
+ PM_SKY130_FD_SC_LP__EINVN_4%Z
x_PM_SKY130_FD_SC_LP__EINVN_4%VPWR N_VPWR_M1005_d N_VPWR_M1015_d N_VPWR_M1011_s
+ N_VPWR_c_517_n N_VPWR_c_518_n N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n
+ N_VPWR_c_522_n VPWR N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_516_n
+ N_VPWR_c_526_n N_VPWR_c_527_n PM_SKY130_FD_SC_LP__EINVN_4%VPWR
x_PM_SKY130_FD_SC_LP__EINVN_4%A_83_69# N_A_83_69#_M1002_s N_A_83_69#_M1003_s
+ N_A_83_69#_M1009_s N_A_83_69#_M1007_d N_A_83_69#_M1012_d N_A_83_69#_c_590_n
+ N_A_83_69#_c_591_n N_A_83_69#_c_592_n N_A_83_69#_c_604_n N_A_83_69#_c_593_n
+ N_A_83_69#_c_594_n N_A_83_69#_c_595_n N_A_83_69#_c_596_n N_A_83_69#_c_622_n
+ N_A_83_69#_c_665_p N_A_83_69#_c_597_n N_A_83_69#_c_634_n N_A_83_69#_c_674_p
+ N_A_83_69#_c_598_n N_A_83_69#_c_599_n N_A_83_69#_c_640_n
+ PM_SKY130_FD_SC_LP__EINVN_4%A_83_69#
x_PM_SKY130_FD_SC_LP__EINVN_4%VGND N_VGND_M1007_s N_VGND_M1008_s N_VGND_M1014_s
+ N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n N_VGND_c_689_n
+ N_VGND_c_690_n VGND N_VGND_c_691_n N_VGND_c_692_n N_VGND_c_693_n
+ N_VGND_c_694_n N_VGND_c_695_n PM_SKY130_FD_SC_LP__EINVN_4%VGND
cc_1 VNB N_A_c_109_n 0.0216848f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.295
cc_2 VNB N_A_c_110_n 0.0163934f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.295
cc_3 VNB N_A_M1004_g 0.0190481f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=0.765
cc_4 VNB N_A_c_112_n 0.0165844f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=1.51
cc_5 VNB N_A_c_113_n 0.06053f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.51
cc_6 VNB N_A_M1009_g 0.0224865f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.765
cc_7 VNB N_A_c_115_n 0.0140279f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.51
cc_8 VNB A 0.0254475f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_9 VNB N_A_555_201#_c_201_n 0.0214187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_555_201#_c_202_n 0.0178973f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.765
cc_11 VNB N_A_555_201#_c_203_n 0.0122506f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_12 VNB N_A_555_201#_c_204_n 0.0150524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_555_201#_c_205_n 0.0121781f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=0.765
cc_14 VNB N_A_555_201#_c_206_n 0.0150524f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.675
cc_15 VNB N_A_555_201#_c_207_n 0.0203578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_555_201#_c_208_n 0.0159142f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.51
cc_17 VNB N_A_555_201#_c_209_n 0.00510736f $X=-0.19 $Y=-0.245 $X2=2.225
+ $Y2=0.765
cc_18 VNB N_A_555_201#_c_210_n 0.00510736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_555_201#_c_211_n 0.00510736f $X=-0.19 $Y=-0.245 $X2=2.225
+ $Y2=1.675
cc_20 VNB N_A_555_201#_c_212_n 0.0408084f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.465
cc_21 VNB N_A_555_201#_c_213_n 0.00404653f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_555_201#_c_214_n 0.0477137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_555_201#_c_215_n 0.00618735f $X=-0.19 $Y=-0.245 $X2=1.215
+ $Y2=1.485
cc_24 VNB N_A_555_201#_c_216_n 0.0354702f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=1.51
cc_25 VNB N_A_555_201#_c_217_n 0.0100025f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.51
cc_26 VNB N_TE_B_c_299_n 0.00669782f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.675
cc_27 VNB N_TE_B_c_300_n 0.00820714f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.465
cc_28 VNB N_TE_B_c_301_n 0.00731825f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.765
cc_29 VNB N_TE_B_c_302_n 0.00724578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_TE_B_c_303_n 0.0110621f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.675
cc_31 VNB N_TE_B_c_304_n 0.0123834f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=2.465
cc_32 VNB N_TE_B_M1016_g 0.0456557f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.345
cc_33 VNB N_TE_B_c_306_n 0.00335787f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.465
cc_34 VNB N_TE_B_c_307_n 0.00399128f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.465
cc_35 VNB N_TE_B_c_308_n 0.00399128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_TE_B_c_309_n 0.00878081f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_37 VNB N_TE_B_c_310_n 0.00325913f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_38 VNB N_Z_c_455_n 0.00361153f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=2.465
cc_39 VNB N_Z_c_456_n 0.00226834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Z_c_457_n 0.0021045f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.675
cc_41 VNB N_VPWR_c_516_n 0.243291f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.51
cc_42 VNB N_A_83_69#_c_590_n 0.0324941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_83_69#_c_591_n 0.00294772f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=2.465
cc_44 VNB N_A_83_69#_c_592_n 0.00949021f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=2.465
cc_45 VNB N_A_83_69#_c_593_n 0.00857099f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=0.765
cc_46 VNB N_A_83_69#_c_594_n 0.00843383f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=2.465
cc_47 VNB N_A_83_69#_c_595_n 0.00411264f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_48 VNB N_A_83_69#_c_596_n 0.0150614f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_49 VNB N_A_83_69#_c_597_n 9.16311e-19 $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.485
cc_50 VNB N_A_83_69#_c_598_n 0.0020362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_83_69#_c_599_n 9.39062e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_685_n 0.00842966f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_53 VNB N_VGND_c_686_n 0.012299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_687_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_688_n 0.00278533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_689_n 0.0791087f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.51
cc_57 VNB N_VGND_c_690_n 0.00510637f $X=-0.19 $Y=-0.245 $X2=2.225 $Y2=1.345
cc_58 VNB N_VGND_c_691_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_59 VNB N_VGND_c_692_n 0.0156941f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.485
cc_60 VNB N_VGND_c_693_n 0.318638f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=1.485
cc_61 VNB N_VGND_c_694_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.485
cc_62 VNB N_VGND_c_695_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.51
cc_63 VPB N_A_M1000_g 0.0253431f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=2.465
cc_64 VPB N_A_M1001_g 0.0190258f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.465
cc_65 VPB N_A_M1010_g 0.019273f $X=-0.19 $Y=1.655 $X2=1.715 $Y2=2.465
cc_66 VPB N_A_c_112_n 0.005666f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=1.51
cc_67 VPB N_A_c_113_n 0.0108876f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=1.51
cc_68 VPB N_A_M1013_g 0.0192388f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=2.465
cc_69 VPB N_A_c_115_n 7.19422e-19 $X=-0.19 $Y=1.655 $X2=2.225 $Y2=1.51
cc_70 VPB A 0.0253613f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_71 VPB N_A_555_201#_c_213_n 0.057485f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_72 VPB N_TE_B_c_311_n 0.0154105f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.295
cc_73 VPB N_TE_B_c_299_n 0.00418369f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=1.675
cc_74 VPB N_TE_B_c_300_n 0.00251208f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=2.465
cc_75 VPB N_TE_B_c_314_n 0.0153032f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=2.465
cc_76 VPB N_TE_B_c_301_n 0.00418344f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=0.765
cc_77 VPB N_TE_B_c_316_n 0.0153032f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=1.675
cc_78 VPB N_TE_B_c_302_n 0.00418369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_TE_B_c_318_n 0.0185047f $X=-0.19 $Y=1.655 $X2=1.715 $Y2=0.765
cc_80 VPB N_TE_B_c_303_n 0.00975675f $X=-0.19 $Y=1.655 $X2=1.715 $Y2=1.675
cc_81 VPB N_TE_B_c_304_n 0.00919828f $X=-0.19 $Y=1.655 $X2=1.715 $Y2=2.465
cc_82 VPB N_TE_B_c_321_n 0.0224491f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=0.765
cc_83 VPB N_TE_B_c_306_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=2.465
cc_84 VPB N_TE_B_c_307_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=2.465
cc_85 VPB N_TE_B_c_308_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_TE_B_c_309_n 0.00245158f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_87 VPB N_TE_B_c_310_n 0.00285174f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_88 VPB N_TE_B_c_327_n 0.0663598f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=1.485
cc_89 VPB N_TE_B_c_328_n 0.0114275f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=1.51
cc_90 VPB N_A_87_367#_c_389_n 0.00746637f $X=-0.19 $Y=1.655 $X2=1.715 $Y2=0.765
cc_91 VPB N_A_87_367#_c_390_n 0.037567f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_87_367#_c_391_n 0.0040407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_87_367#_c_392_n 0.00524713f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=1.51
cc_94 VPB N_A_87_367#_c_393_n 0.00524587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_87_367#_c_394_n 0.0109581f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=1.51
cc_96 VPB N_A_87_367#_c_395_n 0.00124366f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_Z_c_458_n 0.00129923f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=2.465
cc_98 VPB N_VPWR_c_517_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.465
cc_99 VPB N_VPWR_c_518_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.715 $Y2=0.765
cc_100 VPB N_VPWR_c_519_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.715 $Y2=2.465
cc_101 VPB N_VPWR_c_520_n 0.0210688f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=0.765
cc_102 VPB N_VPWR_c_521_n 0.0664745f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=2.465
cc_103 VPB N_VPWR_c_522_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=2.465
cc_104 VPB N_VPWR_c_523_n 0.0269584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_524_n 0.0177367f $X=-0.19 $Y=1.655 $X2=1.6 $Y2=1.51
cc_106 VPB N_VPWR_c_516_n 0.0747678f $X=-0.19 $Y=1.655 $X2=1.6 $Y2=1.51
cc_107 VPB N_VPWR_c_526_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_527_n 0.00545601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 N_A_M1009_g N_A_555_201#_c_215_n 0.00545324f $X=2.225 $Y=0.765 $X2=0
+ $Y2=0
cc_110 N_A_M1009_g N_A_555_201#_c_216_n 0.0061701f $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_111 N_A_M1013_g N_TE_B_c_311_n 0.0123141f $X=2.225 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_c_115_n N_TE_B_c_300_n 0.0123141f $X=2.225 $Y=1.51 $X2=0 $Y2=0
cc_113 A N_A_87_367#_c_390_n 0.0223338f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A_M1000_g N_A_87_367#_c_397_n 0.0126807f $X=0.775 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_M1001_g N_A_87_367#_c_397_n 0.0130869f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_M1010_g N_A_87_367#_c_399_n 0.00916233f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_M1013_g N_A_87_367#_c_399_n 4.70665e-19 $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_M1010_g N_A_87_367#_c_401_n 0.0102775f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_M1013_g N_A_87_367#_c_401_n 0.0119467f $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A_M1013_g N_A_87_367#_c_392_n 6.55961e-19 $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_M1010_g N_A_87_367#_c_404_n 0.00198771f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_c_109_n N_Z_c_459_n 0.00555412f $X=0.775 $Y=1.295 $X2=0 $Y2=0
cc_123 N_A_M1001_g N_Z_c_460_n 0.0103172f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_M1010_g N_Z_c_460_n 4.5114e-19 $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_c_110_n N_Z_c_455_n 0.0128367f $X=1.285 $Y=1.295 $X2=0 $Y2=0
cc_126 N_A_M1004_g N_Z_c_455_n 0.0131979f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_127 N_A_c_113_n N_Z_c_455_n 0.00244902f $X=1.79 $Y=1.51 $X2=0 $Y2=0
cc_128 A N_Z_c_455_n 0.0427906f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A_c_109_n N_Z_c_456_n 0.00453083f $X=0.775 $Y=1.295 $X2=0 $Y2=0
cc_130 N_A_c_113_n N_Z_c_456_n 0.00501355f $X=1.79 $Y=1.51 $X2=0 $Y2=0
cc_131 A N_Z_c_456_n 0.0264172f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_132 N_A_M1001_g N_Z_c_469_n 0.01115f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A_M1010_g N_Z_c_469_n 0.0147907f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A_c_113_n N_Z_c_469_n 5.78305e-19 $X=1.79 $Y=1.51 $X2=0 $Y2=0
cc_135 A N_Z_c_469_n 0.0354567f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A_M1001_g N_Z_c_473_n 7.32094e-19 $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_c_113_n N_Z_c_473_n 0.00117291f $X=1.79 $Y=1.51 $X2=0 $Y2=0
cc_138 A N_Z_c_473_n 0.0257144f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A_M1013_g N_Z_c_476_n 0.00883338f $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A_M1004_g N_Z_c_457_n 0.00243916f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_141 N_A_c_112_n N_Z_c_457_n 0.0128408f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_142 N_A_M1009_g N_Z_c_457_n 0.00659282f $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_143 N_A_c_115_n N_Z_c_457_n 0.00741099f $X=2.225 $Y=1.51 $X2=0 $Y2=0
cc_144 A N_Z_c_457_n 0.00563012f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_145 N_A_M1010_g N_Z_c_458_n 0.00444672f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_c_112_n N_Z_c_458_n 0.00861005f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_147 N_A_M1013_g N_Z_c_458_n 0.00538103f $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_c_115_n N_Z_c_458_n 0.00332755f $X=2.225 $Y=1.51 $X2=0 $Y2=0
cc_149 A N_Z_c_458_n 0.0187144f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A_c_112_n N_Z_c_487_n 0.00178083f $X=2.15 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A_M1013_g N_Z_c_487_n 0.00168611f $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_M1009_g N_Z_c_489_n 0.00863146f $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_153 N_A_M1013_g N_VPWR_c_517_n 0.00109252f $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_M1000_g N_VPWR_c_521_n 0.00357877f $X=0.775 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_M1001_g N_VPWR_c_521_n 0.00357877f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A_M1010_g N_VPWR_c_521_n 0.00357828f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_M1013_g N_VPWR_c_521_n 0.00357877f $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_M1000_g N_VPWR_c_516_n 0.00667903f $X=0.775 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A_M1001_g N_VPWR_c_516_n 0.00563058f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A_M1010_g N_VPWR_c_516_n 0.00563056f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A_M1013_g N_VPWR_c_516_n 0.00558518f $X=2.225 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_c_109_n N_A_83_69#_c_590_n 0.00350947f $X=0.775 $Y=1.295 $X2=0 $Y2=0
cc_163 A N_A_83_69#_c_590_n 0.0197536f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A_c_109_n N_A_83_69#_c_591_n 0.0133384f $X=0.775 $Y=1.295 $X2=0 $Y2=0
cc_165 N_A_c_110_n N_A_83_69#_c_591_n 0.00865124f $X=1.285 $Y=1.295 $X2=0 $Y2=0
cc_166 N_A_c_109_n N_A_83_69#_c_604_n 5.37284e-19 $X=0.775 $Y=1.295 $X2=0 $Y2=0
cc_167 N_A_c_110_n N_A_83_69#_c_604_n 0.00677031f $X=1.285 $Y=1.295 $X2=0 $Y2=0
cc_168 N_A_M1004_g N_A_83_69#_c_604_n 0.00677031f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_169 N_A_M1009_g N_A_83_69#_c_604_n 5.37284e-19 $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_170 N_A_M1004_g N_A_83_69#_c_593_n 0.00865124f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_171 N_A_M1009_g N_A_83_69#_c_593_n 0.013004f $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_172 N_A_M1009_g N_A_83_69#_c_594_n 0.00916024f $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_173 N_A_M1009_g N_A_83_69#_c_595_n 0.00441984f $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_174 N_A_c_110_n N_A_83_69#_c_598_n 0.00159238f $X=1.285 $Y=1.295 $X2=0 $Y2=0
cc_175 N_A_M1004_g N_A_83_69#_c_598_n 0.00159238f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_176 N_A_M1009_g N_A_83_69#_c_599_n 0.00363151f $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_177 N_A_c_109_n N_VGND_c_689_n 0.0029147f $X=0.775 $Y=1.295 $X2=0 $Y2=0
cc_178 N_A_c_110_n N_VGND_c_689_n 0.00291444f $X=1.285 $Y=1.295 $X2=0 $Y2=0
cc_179 N_A_M1004_g N_VGND_c_689_n 0.00291444f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_180 N_A_M1009_g N_VGND_c_689_n 0.0029147f $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_181 N_A_c_109_n N_VGND_c_693_n 0.00428931f $X=0.775 $Y=1.295 $X2=0 $Y2=0
cc_182 N_A_c_110_n N_VGND_c_693_n 0.00403101f $X=1.285 $Y=1.295 $X2=0 $Y2=0
cc_183 N_A_M1004_g N_VGND_c_693_n 0.00403101f $X=1.715 $Y=0.765 $X2=0 $Y2=0
cc_184 N_A_M1009_g N_VGND_c_693_n 0.00433096f $X=2.225 $Y=0.765 $X2=0 $Y2=0
cc_185 N_A_555_201#_c_215_n N_TE_B_c_299_n 0.00313882f $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_186 N_A_555_201#_c_216_n N_TE_B_c_299_n 0.0138318f $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_187 N_A_555_201#_c_209_n N_TE_B_c_301_n 0.0138318f $X=3.555 $Y=1.26 $X2=0
+ $Y2=0
cc_188 N_A_555_201#_c_210_n N_TE_B_c_302_n 0.0138318f $X=3.985 $Y=1.26 $X2=0
+ $Y2=0
cc_189 N_A_555_201#_c_211_n N_TE_B_c_303_n 0.0138318f $X=4.415 $Y=1.26 $X2=0
+ $Y2=0
cc_190 N_A_555_201#_c_208_n N_TE_B_M1016_g 0.0262526f $X=4.845 $Y=1.185 $X2=0
+ $Y2=0
cc_191 N_A_555_201#_c_212_n N_TE_B_M1016_g 0.019415f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_192 N_A_555_201#_c_214_n N_TE_B_M1016_g 0.013437f $X=5.49 $Y=0.42 $X2=0 $Y2=0
cc_193 N_A_555_201#_c_217_n N_TE_B_M1016_g 0.00359621f $X=5.502 $Y=1.485 $X2=0
+ $Y2=0
cc_194 N_A_555_201#_c_201_n N_TE_B_c_306_n 0.0138318f $X=3.48 $Y=1.26 $X2=0
+ $Y2=0
cc_195 N_A_555_201#_c_212_n N_TE_B_c_306_n 0.0299362f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_196 N_A_555_201#_c_203_n N_TE_B_c_307_n 0.0138318f $X=3.91 $Y=1.26 $X2=0
+ $Y2=0
cc_197 N_A_555_201#_c_205_n N_TE_B_c_308_n 0.0138318f $X=4.34 $Y=1.26 $X2=0
+ $Y2=0
cc_198 N_A_555_201#_c_207_n N_TE_B_c_309_n 0.0138318f $X=4.77 $Y=1.26 $X2=0
+ $Y2=0
cc_199 N_A_555_201#_c_213_n N_TE_B_c_310_n 0.0144719f $X=5.49 $Y=1.98 $X2=0
+ $Y2=0
cc_200 N_A_555_201#_c_212_n N_TE_B_c_328_n 0.0202992f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_201 N_A_555_201#_c_213_n N_TE_B_c_328_n 0.00199757f $X=5.49 $Y=1.98 $X2=0
+ $Y2=0
cc_202 N_A_555_201#_c_212_n N_A_87_367#_c_391_n 0.00701646f $X=5.35 $Y=1.485
+ $X2=0 $Y2=0
cc_203 N_A_555_201#_c_215_n N_A_87_367#_c_391_n 0.0241394f $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_204 N_A_555_201#_c_216_n N_A_87_367#_c_391_n 3.62792e-19 $X=2.94 $Y=1.17
+ $X2=0 $Y2=0
cc_205 N_A_555_201#_c_212_n N_A_87_367#_c_393_n 0.066557f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_206 N_A_555_201#_c_212_n N_A_87_367#_c_395_n 0.0154605f $X=5.35 $Y=1.485
+ $X2=0 $Y2=0
cc_207 N_A_555_201#_c_215_n N_Z_c_457_n 0.00758183f $X=2.94 $Y=1.17 $X2=0 $Y2=0
cc_208 N_A_555_201#_c_216_n N_Z_c_457_n 3.59623e-19 $X=2.94 $Y=1.17 $X2=0 $Y2=0
cc_209 N_A_555_201#_c_215_n N_Z_c_458_n 0.00222222f $X=2.94 $Y=1.17 $X2=0 $Y2=0
cc_210 N_A_555_201#_c_212_n N_VPWR_c_520_n 0.0188163f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_211 N_A_555_201#_c_213_n N_VPWR_c_520_n 0.0463652f $X=5.49 $Y=1.98 $X2=0
+ $Y2=0
cc_212 N_A_555_201#_c_213_n N_VPWR_c_524_n 0.0194077f $X=5.49 $Y=1.98 $X2=0
+ $Y2=0
cc_213 N_A_555_201#_M1011_d N_VPWR_c_516_n 0.00215158f $X=5.35 $Y=1.835 $X2=0
+ $Y2=0
cc_214 N_A_555_201#_c_213_n N_VPWR_c_516_n 0.0117799f $X=5.49 $Y=1.98 $X2=0
+ $Y2=0
cc_215 N_A_555_201#_c_215_n N_A_83_69#_c_595_n 0.0149977f $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_216 N_A_555_201#_c_216_n N_A_83_69#_c_595_n 0.00325523f $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_217 N_A_555_201#_c_201_n N_A_83_69#_c_596_n 0.00698732f $X=3.48 $Y=1.26 $X2=0
+ $Y2=0
cc_218 N_A_555_201#_c_202_n N_A_83_69#_c_596_n 0.0114319f $X=3.555 $Y=1.185
+ $X2=0 $Y2=0
cc_219 N_A_555_201#_c_212_n N_A_83_69#_c_596_n 0.0160012f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_220 N_A_555_201#_c_215_n N_A_83_69#_c_596_n 0.0256187f $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_221 N_A_555_201#_c_216_n N_A_83_69#_c_596_n 0.0079693f $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_222 N_A_555_201#_c_202_n N_A_83_69#_c_622_n 0.00554129f $X=3.555 $Y=1.185
+ $X2=0 $Y2=0
cc_223 N_A_555_201#_c_216_n N_A_83_69#_c_622_n 2.55384e-19 $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_224 N_A_555_201#_c_203_n N_A_83_69#_c_597_n 4.79475e-19 $X=3.91 $Y=1.26 $X2=0
+ $Y2=0
cc_225 N_A_555_201#_c_204_n N_A_83_69#_c_597_n 0.0104457f $X=3.985 $Y=1.185
+ $X2=0 $Y2=0
cc_226 N_A_555_201#_c_205_n N_A_83_69#_c_597_n 0.0047604f $X=4.34 $Y=1.26 $X2=0
+ $Y2=0
cc_227 N_A_555_201#_c_206_n N_A_83_69#_c_597_n 0.0101922f $X=4.415 $Y=1.185
+ $X2=0 $Y2=0
cc_228 N_A_555_201#_c_207_n N_A_83_69#_c_597_n 0.00577238f $X=4.77 $Y=1.26 $X2=0
+ $Y2=0
cc_229 N_A_555_201#_c_208_n N_A_83_69#_c_597_n 0.00150086f $X=4.845 $Y=1.185
+ $X2=0 $Y2=0
cc_230 N_A_555_201#_c_210_n N_A_83_69#_c_597_n 0.00167259f $X=3.985 $Y=1.26
+ $X2=0 $Y2=0
cc_231 N_A_555_201#_c_211_n N_A_83_69#_c_597_n 0.00167259f $X=4.415 $Y=1.26
+ $X2=0 $Y2=0
cc_232 N_A_555_201#_c_212_n N_A_83_69#_c_597_n 0.0631764f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_233 N_A_555_201#_c_214_n N_A_83_69#_c_597_n 0.00341507f $X=5.49 $Y=0.42 $X2=0
+ $Y2=0
cc_234 N_A_555_201#_c_202_n N_A_83_69#_c_634_n 0.00358552f $X=3.555 $Y=1.185
+ $X2=0 $Y2=0
cc_235 N_A_555_201#_c_203_n N_A_83_69#_c_634_n 0.00502885f $X=3.91 $Y=1.26 $X2=0
+ $Y2=0
cc_236 N_A_555_201#_c_209_n N_A_83_69#_c_634_n 0.00133413f $X=3.555 $Y=1.26
+ $X2=0 $Y2=0
cc_237 N_A_555_201#_c_212_n N_A_83_69#_c_634_n 0.0206864f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_238 N_A_555_201#_c_215_n N_A_83_69#_c_634_n 0.00526542f $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_239 N_A_555_201#_c_216_n N_A_83_69#_c_634_n 4.63568e-19 $X=2.94 $Y=1.17 $X2=0
+ $Y2=0
cc_240 N_A_555_201#_c_202_n N_A_83_69#_c_640_n 0.00111029f $X=3.555 $Y=1.185
+ $X2=0 $Y2=0
cc_241 N_A_555_201#_c_202_n N_VGND_c_685_n 0.00841028f $X=3.555 $Y=1.185 $X2=0
+ $Y2=0
cc_242 N_A_555_201#_c_204_n N_VGND_c_685_n 5.34794e-19 $X=3.985 $Y=1.185 $X2=0
+ $Y2=0
cc_243 N_A_555_201#_c_202_n N_VGND_c_686_n 0.00364061f $X=3.555 $Y=1.185 $X2=0
+ $Y2=0
cc_244 N_A_555_201#_c_204_n N_VGND_c_686_n 0.00486043f $X=3.985 $Y=1.185 $X2=0
+ $Y2=0
cc_245 N_A_555_201#_c_202_n N_VGND_c_687_n 6.32445e-19 $X=3.555 $Y=1.185 $X2=0
+ $Y2=0
cc_246 N_A_555_201#_c_204_n N_VGND_c_687_n 0.0112649f $X=3.985 $Y=1.185 $X2=0
+ $Y2=0
cc_247 N_A_555_201#_c_205_n N_VGND_c_687_n 5.83892e-19 $X=4.34 $Y=1.26 $X2=0
+ $Y2=0
cc_248 N_A_555_201#_c_206_n N_VGND_c_687_n 0.0112765f $X=4.415 $Y=1.185 $X2=0
+ $Y2=0
cc_249 N_A_555_201#_c_208_n N_VGND_c_687_n 6.28154e-19 $X=4.845 $Y=1.185 $X2=0
+ $Y2=0
cc_250 N_A_555_201#_c_206_n N_VGND_c_688_n 7.11292e-19 $X=4.415 $Y=1.185 $X2=0
+ $Y2=0
cc_251 N_A_555_201#_c_208_n N_VGND_c_688_n 0.0155048f $X=4.845 $Y=1.185 $X2=0
+ $Y2=0
cc_252 N_A_555_201#_c_212_n N_VGND_c_688_n 0.0193099f $X=5.35 $Y=1.485 $X2=0
+ $Y2=0
cc_253 N_A_555_201#_c_214_n N_VGND_c_688_n 0.0338343f $X=5.49 $Y=0.42 $X2=0
+ $Y2=0
cc_254 N_A_555_201#_c_206_n N_VGND_c_691_n 0.00486043f $X=4.415 $Y=1.185 $X2=0
+ $Y2=0
cc_255 N_A_555_201#_c_208_n N_VGND_c_691_n 0.00486043f $X=4.845 $Y=1.185 $X2=0
+ $Y2=0
cc_256 N_A_555_201#_c_214_n N_VGND_c_692_n 0.0178111f $X=5.49 $Y=0.42 $X2=0
+ $Y2=0
cc_257 N_A_555_201#_M1016_d N_VGND_c_693_n 0.00371702f $X=5.35 $Y=0.235 $X2=0
+ $Y2=0
cc_258 N_A_555_201#_c_202_n N_VGND_c_693_n 0.00430125f $X=3.555 $Y=1.185 $X2=0
+ $Y2=0
cc_259 N_A_555_201#_c_204_n N_VGND_c_693_n 0.00824727f $X=3.985 $Y=1.185 $X2=0
+ $Y2=0
cc_260 N_A_555_201#_c_206_n N_VGND_c_693_n 0.00824727f $X=4.415 $Y=1.185 $X2=0
+ $Y2=0
cc_261 N_A_555_201#_c_208_n N_VGND_c_693_n 0.00824727f $X=4.845 $Y=1.185 $X2=0
+ $Y2=0
cc_262 N_A_555_201#_c_214_n N_VGND_c_693_n 0.0100304f $X=5.49 $Y=0.42 $X2=0
+ $Y2=0
cc_263 N_TE_B_c_311_n N_A_87_367#_c_391_n 0.0162583f $X=2.655 $Y=1.725 $X2=0
+ $Y2=0
cc_264 N_TE_B_c_299_n N_A_87_367#_c_391_n 0.00227624f $X=3.01 $Y=1.65 $X2=0
+ $Y2=0
cc_265 N_TE_B_c_314_n N_A_87_367#_c_391_n 0.0128694f $X=3.085 $Y=1.725 $X2=0
+ $Y2=0
cc_266 N_TE_B_c_316_n N_A_87_367#_c_393_n 0.0125267f $X=3.515 $Y=1.725 $X2=0
+ $Y2=0
cc_267 N_TE_B_c_302_n N_A_87_367#_c_393_n 0.0022778f $X=3.87 $Y=1.65 $X2=0 $Y2=0
cc_268 N_TE_B_c_318_n N_A_87_367#_c_393_n 0.0126566f $X=3.945 $Y=1.725 $X2=0
+ $Y2=0
cc_269 N_TE_B_c_303_n N_A_87_367#_c_393_n 0.00456055f $X=4.445 $Y=1.65 $X2=0
+ $Y2=0
cc_270 N_TE_B_c_327_n N_A_87_367#_c_393_n 0.00157151f $X=4.61 $Y=1.91 $X2=0
+ $Y2=0
cc_271 N_TE_B_c_328_n N_A_87_367#_c_393_n 0.0140879f $X=4.61 $Y=1.91 $X2=0 $Y2=0
cc_272 N_TE_B_c_327_n N_A_87_367#_c_394_n 0.00416939f $X=4.61 $Y=1.91 $X2=0
+ $Y2=0
cc_273 N_TE_B_c_328_n N_A_87_367#_c_394_n 0.07242f $X=4.61 $Y=1.91 $X2=0 $Y2=0
cc_274 N_TE_B_c_301_n N_A_87_367#_c_395_n 0.00240029f $X=3.44 $Y=1.65 $X2=0
+ $Y2=0
cc_275 N_TE_B_c_300_n N_Z_c_458_n 0.00101917f $X=2.73 $Y=1.65 $X2=0 $Y2=0
cc_276 N_TE_B_c_311_n N_VPWR_c_517_n 0.0153918f $X=2.655 $Y=1.725 $X2=0 $Y2=0
cc_277 N_TE_B_c_314_n N_VPWR_c_517_n 0.0142189f $X=3.085 $Y=1.725 $X2=0 $Y2=0
cc_278 N_TE_B_c_316_n N_VPWR_c_517_n 7.27171e-19 $X=3.515 $Y=1.725 $X2=0 $Y2=0
cc_279 N_TE_B_c_314_n N_VPWR_c_518_n 0.00486043f $X=3.085 $Y=1.725 $X2=0 $Y2=0
cc_280 N_TE_B_c_316_n N_VPWR_c_518_n 0.00486043f $X=3.515 $Y=1.725 $X2=0 $Y2=0
cc_281 N_TE_B_c_314_n N_VPWR_c_519_n 7.27171e-19 $X=3.085 $Y=1.725 $X2=0 $Y2=0
cc_282 N_TE_B_c_316_n N_VPWR_c_519_n 0.0142189f $X=3.515 $Y=1.725 $X2=0 $Y2=0
cc_283 N_TE_B_c_318_n N_VPWR_c_519_n 0.0160927f $X=3.945 $Y=1.725 $X2=0 $Y2=0
cc_284 N_TE_B_c_304_n N_VPWR_c_520_n 0.00499972f $X=5.2 $Y=1.65 $X2=0 $Y2=0
cc_285 N_TE_B_c_321_n N_VPWR_c_520_n 0.00792822f $X=5.275 $Y=1.725 $X2=0 $Y2=0
cc_286 N_TE_B_c_327_n N_VPWR_c_520_n 0.00543664f $X=4.61 $Y=1.91 $X2=0 $Y2=0
cc_287 N_TE_B_c_328_n N_VPWR_c_520_n 0.0819993f $X=4.61 $Y=1.91 $X2=0 $Y2=0
cc_288 N_TE_B_c_311_n N_VPWR_c_521_n 0.00486043f $X=2.655 $Y=1.725 $X2=0 $Y2=0
cc_289 N_TE_B_c_318_n N_VPWR_c_523_n 0.00486043f $X=3.945 $Y=1.725 $X2=0 $Y2=0
cc_290 N_TE_B_c_328_n N_VPWR_c_523_n 0.00758553f $X=4.61 $Y=1.91 $X2=0 $Y2=0
cc_291 N_TE_B_c_321_n N_VPWR_c_524_n 0.00585385f $X=5.275 $Y=1.725 $X2=0 $Y2=0
cc_292 N_TE_B_c_311_n N_VPWR_c_516_n 0.0082726f $X=2.655 $Y=1.725 $X2=0 $Y2=0
cc_293 N_TE_B_c_314_n N_VPWR_c_516_n 0.00824727f $X=3.085 $Y=1.725 $X2=0 $Y2=0
cc_294 N_TE_B_c_316_n N_VPWR_c_516_n 0.00824727f $X=3.515 $Y=1.725 $X2=0 $Y2=0
cc_295 N_TE_B_c_318_n N_VPWR_c_516_n 0.00954696f $X=3.945 $Y=1.725 $X2=0 $Y2=0
cc_296 N_TE_B_c_321_n N_VPWR_c_516_n 0.0127914f $X=5.275 $Y=1.725 $X2=0 $Y2=0
cc_297 N_TE_B_c_328_n N_VPWR_c_516_n 0.00864285f $X=4.61 $Y=1.91 $X2=0 $Y2=0
cc_298 N_TE_B_c_300_n N_A_83_69#_c_595_n 6.44124e-19 $X=2.73 $Y=1.65 $X2=0 $Y2=0
cc_299 N_TE_B_c_300_n N_A_83_69#_c_596_n 0.00243253f $X=2.73 $Y=1.65 $X2=0 $Y2=0
cc_300 N_TE_B_c_300_n N_A_83_69#_c_599_n 0.00197688f $X=2.73 $Y=1.65 $X2=0 $Y2=0
cc_301 N_TE_B_M1016_g N_VGND_c_688_n 0.0175836f $X=5.275 $Y=0.655 $X2=0 $Y2=0
cc_302 N_TE_B_M1016_g N_VGND_c_692_n 0.00486043f $X=5.275 $Y=0.655 $X2=0 $Y2=0
cc_303 N_TE_B_M1016_g N_VGND_c_693_n 0.00918921f $X=5.275 $Y=0.655 $X2=0 $Y2=0
cc_304 N_A_87_367#_c_397_n N_Z_M1000_d 0.0049251f $X=1.405 $Y=2.99 $X2=0 $Y2=0
cc_305 N_A_87_367#_c_401_n N_Z_M1010_d 0.0049251f $X=2.345 $Y=2.99 $X2=0 $Y2=0
cc_306 N_A_87_367#_c_397_n N_Z_c_460_n 0.0203966f $X=1.405 $Y=2.99 $X2=0 $Y2=0
cc_307 N_A_87_367#_M1001_s N_Z_c_469_n 0.00332836f $X=1.36 $Y=1.835 $X2=0 $Y2=0
cc_308 N_A_87_367#_c_399_n N_Z_c_469_n 0.0160534f $X=1.5 $Y=2.425 $X2=0 $Y2=0
cc_309 N_A_87_367#_c_401_n N_Z_c_476_n 0.0203966f $X=2.345 $Y=2.99 $X2=0 $Y2=0
cc_310 N_A_87_367#_c_392_n N_Z_c_458_n 0.00953297f $X=2.535 $Y=1.84 $X2=0 $Y2=0
cc_311 N_A_87_367#_c_391_n N_VPWR_M1005_d 0.00176461f $X=3.205 $Y=1.84 $X2=-0.19
+ $Y2=1.655
cc_312 N_A_87_367#_c_393_n N_VPWR_M1015_d 0.00176461f $X=4.065 $Y=1.84 $X2=0
+ $Y2=0
cc_313 N_A_87_367#_c_391_n N_VPWR_c_517_n 0.0170777f $X=3.205 $Y=1.84 $X2=0
+ $Y2=0
cc_314 N_A_87_367#_c_432_p N_VPWR_c_518_n 0.0124525f $X=3.3 $Y=1.98 $X2=0 $Y2=0
cc_315 N_A_87_367#_c_393_n N_VPWR_c_519_n 0.0170777f $X=4.065 $Y=1.84 $X2=0
+ $Y2=0
cc_316 N_A_87_367#_c_394_n N_VPWR_c_520_n 0.00722531f $X=4.16 $Y=1.98 $X2=0
+ $Y2=0
cc_317 N_A_87_367#_c_389_n N_VPWR_c_521_n 0.0182731f $X=0.53 $Y=2.905 $X2=0
+ $Y2=0
cc_318 N_A_87_367#_c_397_n N_VPWR_c_521_n 0.0408615f $X=1.405 $Y=2.99 $X2=0
+ $Y2=0
cc_319 N_A_87_367#_c_401_n N_VPWR_c_521_n 0.037448f $X=2.345 $Y=2.99 $X2=0 $Y2=0
cc_320 N_A_87_367#_c_438_p N_VPWR_c_521_n 0.0125234f $X=2.44 $Y=2.905 $X2=0
+ $Y2=0
cc_321 N_A_87_367#_c_404_n N_VPWR_c_521_n 0.0165061f $X=1.54 $Y=2.99 $X2=0 $Y2=0
cc_322 N_A_87_367#_c_394_n N_VPWR_c_523_n 0.0160189f $X=4.16 $Y=1.98 $X2=0 $Y2=0
cc_323 N_A_87_367#_M1000_s N_VPWR_c_516_n 0.0021516f $X=0.435 $Y=1.835 $X2=0
+ $Y2=0
cc_324 N_A_87_367#_M1001_s N_VPWR_c_516_n 0.0022517f $X=1.36 $Y=1.835 $X2=0
+ $Y2=0
cc_325 N_A_87_367#_M1013_s N_VPWR_c_516_n 0.00376627f $X=2.3 $Y=1.835 $X2=0
+ $Y2=0
cc_326 N_A_87_367#_M1006_s N_VPWR_c_516_n 0.00536646f $X=3.16 $Y=1.835 $X2=0
+ $Y2=0
cc_327 N_A_87_367#_M1017_s N_VPWR_c_516_n 0.00371702f $X=4.02 $Y=1.835 $X2=0
+ $Y2=0
cc_328 N_A_87_367#_c_389_n N_VPWR_c_516_n 0.010497f $X=0.53 $Y=2.905 $X2=0 $Y2=0
cc_329 N_A_87_367#_c_397_n N_VPWR_c_516_n 0.0263785f $X=1.405 $Y=2.99 $X2=0
+ $Y2=0
cc_330 N_A_87_367#_c_401_n N_VPWR_c_516_n 0.0239065f $X=2.345 $Y=2.99 $X2=0
+ $Y2=0
cc_331 N_A_87_367#_c_438_p N_VPWR_c_516_n 0.00738676f $X=2.44 $Y=2.905 $X2=0
+ $Y2=0
cc_332 N_A_87_367#_c_432_p N_VPWR_c_516_n 0.00730901f $X=3.3 $Y=1.98 $X2=0 $Y2=0
cc_333 N_A_87_367#_c_394_n N_VPWR_c_516_n 0.0090585f $X=4.16 $Y=1.98 $X2=0 $Y2=0
cc_334 N_A_87_367#_c_404_n N_VPWR_c_516_n 0.0103368f $X=1.54 $Y=2.99 $X2=0 $Y2=0
cc_335 N_A_87_367#_c_391_n N_A_83_69#_c_595_n 0.00268372f $X=3.205 $Y=1.84 $X2=0
+ $Y2=0
cc_336 N_A_87_367#_c_392_n N_A_83_69#_c_595_n 0.00533237f $X=2.535 $Y=1.84 $X2=0
+ $Y2=0
cc_337 N_Z_M1000_d N_VPWR_c_516_n 0.00289524f $X=0.85 $Y=1.835 $X2=0 $Y2=0
cc_338 N_Z_M1010_d N_VPWR_c_516_n 0.00289524f $X=1.79 $Y=1.835 $X2=0 $Y2=0
cc_339 N_Z_c_455_n N_A_83_69#_M1003_s 0.00180746f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_340 N_Z_c_456_n N_A_83_69#_c_590_n 0.00596878f $X=1.155 $Y=1.16 $X2=0 $Y2=0
cc_341 N_Z_M1002_d N_A_83_69#_c_591_n 0.00261503f $X=0.85 $Y=0.345 $X2=0 $Y2=0
cc_342 N_Z_c_459_n N_A_83_69#_c_591_n 0.0203258f $X=0.99 $Y=0.68 $X2=0 $Y2=0
cc_343 N_Z_c_455_n N_A_83_69#_c_591_n 0.00275981f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_344 N_Z_c_455_n N_A_83_69#_c_604_n 0.0162706f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_345 N_Z_M1004_d N_A_83_69#_c_593_n 0.00261503f $X=1.79 $Y=0.345 $X2=0 $Y2=0
cc_346 N_Z_c_455_n N_A_83_69#_c_593_n 0.00275981f $X=1.845 $Y=1.16 $X2=0 $Y2=0
cc_347 N_Z_c_489_n N_A_83_69#_c_593_n 0.0253584f $X=2.01 $Y=0.68 $X2=0 $Y2=0
cc_348 N_Z_c_489_n N_A_83_69#_c_594_n 0.0100159f $X=2.01 $Y=0.68 $X2=0 $Y2=0
cc_349 N_Z_c_457_n N_A_83_69#_c_595_n 0.0150591f $X=2.06 $Y=1.5 $X2=0 $Y2=0
cc_350 N_Z_c_489_n N_A_83_69#_c_595_n 0.0135268f $X=2.01 $Y=0.68 $X2=0 $Y2=0
cc_351 N_Z_c_489_n N_A_83_69#_c_599_n 0.01423f $X=2.01 $Y=0.68 $X2=0 $Y2=0
cc_352 N_A_83_69#_c_596_n N_VGND_M1007_s 0.00579523f $X=3.605 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_353 N_A_83_69#_c_597_n N_VGND_M1008_s 0.00176461f $X=4.535 $Y=1.14 $X2=0
+ $Y2=0
cc_354 N_A_83_69#_c_593_n N_VGND_c_685_n 0.00710986f $X=2.415 $Y=0.34 $X2=0
+ $Y2=0
cc_355 N_A_83_69#_c_594_n N_VGND_c_685_n 0.005022f $X=2.51 $Y=0.49 $X2=0 $Y2=0
cc_356 N_A_83_69#_c_596_n N_VGND_c_685_n 0.0211535f $X=3.605 $Y=0.81 $X2=0 $Y2=0
cc_357 N_A_83_69#_c_596_n N_VGND_c_686_n 0.00132283f $X=3.605 $Y=0.81 $X2=0
+ $Y2=0
cc_358 N_A_83_69#_c_665_p N_VGND_c_686_n 0.0124525f $X=3.77 $Y=0.42 $X2=0 $Y2=0
cc_359 N_A_83_69#_c_640_n N_VGND_c_686_n 7.09976e-19 $X=3.735 $Y=0.81 $X2=0
+ $Y2=0
cc_360 N_A_83_69#_c_597_n N_VGND_c_687_n 0.0170776f $X=4.535 $Y=1.14 $X2=0 $Y2=0
cc_361 N_A_83_69#_c_597_n N_VGND_c_688_n 0.0040802f $X=4.535 $Y=1.14 $X2=0 $Y2=0
cc_362 N_A_83_69#_c_591_n N_VGND_c_689_n 0.0435927f $X=1.335 $Y=0.34 $X2=0 $Y2=0
cc_363 N_A_83_69#_c_592_n N_VGND_c_689_n 0.0193554f $X=0.645 $Y=0.34 $X2=0 $Y2=0
cc_364 N_A_83_69#_c_593_n N_VGND_c_689_n 0.0660734f $X=2.415 $Y=0.34 $X2=0 $Y2=0
cc_365 N_A_83_69#_c_596_n N_VGND_c_689_n 0.00758733f $X=3.605 $Y=0.81 $X2=0
+ $Y2=0
cc_366 N_A_83_69#_c_598_n N_VGND_c_689_n 0.0233745f $X=1.5 $Y=0.34 $X2=0 $Y2=0
cc_367 N_A_83_69#_c_674_p N_VGND_c_691_n 0.0124525f $X=4.63 $Y=0.42 $X2=0 $Y2=0
cc_368 N_A_83_69#_M1007_d N_VGND_c_693_n 0.00400839f $X=3.63 $Y=0.235 $X2=0
+ $Y2=0
cc_369 N_A_83_69#_M1012_d N_VGND_c_693_n 0.00536646f $X=4.49 $Y=0.235 $X2=0
+ $Y2=0
cc_370 N_A_83_69#_c_591_n N_VGND_c_693_n 0.0246836f $X=1.335 $Y=0.34 $X2=0 $Y2=0
cc_371 N_A_83_69#_c_592_n N_VGND_c_693_n 0.010497f $X=0.645 $Y=0.34 $X2=0 $Y2=0
cc_372 N_A_83_69#_c_593_n N_VGND_c_693_n 0.0370433f $X=2.415 $Y=0.34 $X2=0 $Y2=0
cc_373 N_A_83_69#_c_596_n N_VGND_c_693_n 0.016796f $X=3.605 $Y=0.81 $X2=0 $Y2=0
cc_374 N_A_83_69#_c_665_p N_VGND_c_693_n 0.00730901f $X=3.77 $Y=0.42 $X2=0 $Y2=0
cc_375 N_A_83_69#_c_674_p N_VGND_c_693_n 0.00730901f $X=4.63 $Y=0.42 $X2=0 $Y2=0
cc_376 N_A_83_69#_c_598_n N_VGND_c_693_n 0.0125806f $X=1.5 $Y=0.34 $X2=0 $Y2=0
cc_377 N_A_83_69#_c_640_n N_VGND_c_693_n 0.00178457f $X=3.735 $Y=0.81 $X2=0
+ $Y2=0
