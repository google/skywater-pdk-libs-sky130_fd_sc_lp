* File: sky130_fd_sc_lp__buflp_m.pxi.spice
* Created: Wed Sep  2 09:36:53 2020
* 
x_PM_SKY130_FD_SC_LP__BUFLP_M%A_90_94# N_A_90_94#_M1005_d N_A_90_94#_M1006_d
+ N_A_90_94#_M1004_g N_A_90_94#_M1003_g N_A_90_94#_M1001_g N_A_90_94#_M1007_g
+ N_A_90_94#_c_37_n N_A_90_94#_c_38_n N_A_90_94#_c_39_n N_A_90_94#_c_40_n
+ N_A_90_94#_c_41_n N_A_90_94#_c_42_n PM_SKY130_FD_SC_LP__BUFLP_M%A_90_94#
x_PM_SKY130_FD_SC_LP__BUFLP_M%A N_A_M1000_g N_A_M1002_g N_A_M1005_g N_A_M1006_g
+ A A A A N_A_c_98_n PM_SKY130_FD_SC_LP__BUFLP_M%A
x_PM_SKY130_FD_SC_LP__BUFLP_M%X N_X_M1004_s N_X_M1003_s X X X X X X X
+ PM_SKY130_FD_SC_LP__BUFLP_M%X
x_PM_SKY130_FD_SC_LP__BUFLP_M%VPWR N_VPWR_M1007_d N_VPWR_c_152_n VPWR
+ N_VPWR_c_153_n N_VPWR_c_154_n N_VPWR_c_151_n N_VPWR_c_156_n
+ PM_SKY130_FD_SC_LP__BUFLP_M%VPWR
x_PM_SKY130_FD_SC_LP__BUFLP_M%VGND N_VGND_M1001_d N_VGND_c_177_n VGND
+ N_VGND_c_178_n N_VGND_c_179_n N_VGND_c_180_n N_VGND_c_181_n
+ PM_SKY130_FD_SC_LP__BUFLP_M%VGND
cc_1 VNB N_A_90_94#_M1004_g 0.0232705f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.81
cc_2 VNB N_A_90_94#_M1001_g 0.0193684f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.81
cc_3 VNB N_A_90_94#_c_37_n 0.0230061f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=1.295
cc_4 VNB N_A_90_94#_c_38_n 0.0340344f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.81
cc_5 VNB N_A_90_94#_c_39_n 0.0146326f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=2.66
cc_6 VNB N_A_90_94#_c_40_n 0.00149134f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.375
cc_7 VNB N_A_90_94#_c_41_n 0.047098f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.375
cc_8 VNB N_A_90_94#_c_42_n 0.0121667f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=1.295
cc_9 VNB N_A_M1000_g 0.0348888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_M1005_g 0.0444673f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.88
cc_11 VNB A 6.94636e-19 $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.81
cc_12 VNB N_A_c_98_n 0.0171708f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.295
cc_13 VNB X 0.0543409f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.375
cc_14 VNB N_VPWR_c_151_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_177_n 0.0251758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_178_n 0.0296187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_179_n 0.0359871f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.81
cc_18 VNB N_VGND_c_180_n 0.188215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_181_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.66
cc_20 VPB N_A_90_94#_M1003_g 0.0482446f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.66
cc_21 VPB N_A_90_94#_M1007_g 0.0411664f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.66
cc_22 VPB N_A_90_94#_c_39_n 0.0592253f $X=-0.19 $Y=1.655 $X2=2.05 $Y2=2.66
cc_23 VPB N_A_90_94#_c_40_n 0.00243924f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=1.375
cc_24 VPB N_A_90_94#_c_41_n 0.0261033f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=1.375
cc_25 VPB N_A_M1002_g 0.0224776f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.375
cc_26 VPB N_A_M1006_g 0.0248784f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=1.21
cc_27 VPB A 0.00239195f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.81
cc_28 VPB N_A_c_98_n 0.0687135f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=1.295
cc_29 VPB X 0.0545352f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.375
cc_30 VPB N_VPWR_c_152_n 0.0263604f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_153_n 0.0305734f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_154_n 0.0335359f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.81
cc_33 VPB N_VPWR_c_151_n 0.0805702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_156_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.66
cc_35 N_A_90_94#_M1001_g N_A_M1000_g 0.0167142f $X=0.885 $Y=0.81 $X2=0 $Y2=0
cc_36 N_A_90_94#_c_37_n N_A_M1000_g 0.0179108f $X=1.755 $Y=1.295 $X2=0 $Y2=0
cc_37 N_A_90_94#_c_38_n N_A_M1000_g 0.00213451f $X=1.92 $Y=0.81 $X2=0 $Y2=0
cc_38 N_A_90_94#_c_40_n N_A_M1000_g 0.00180027f $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_39 N_A_90_94#_c_41_n N_A_M1000_g 0.0268715f $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_40 N_A_90_94#_M1007_g N_A_M1002_g 0.0172568f $X=0.915 $Y=2.66 $X2=0 $Y2=0
cc_41 N_A_90_94#_c_37_n N_A_M1005_g 0.0108847f $X=1.755 $Y=1.295 $X2=0 $Y2=0
cc_42 N_A_90_94#_c_38_n N_A_M1005_g 0.0163406f $X=1.92 $Y=0.81 $X2=0 $Y2=0
cc_43 N_A_90_94#_c_39_n N_A_M1005_g 0.00596098f $X=2.05 $Y=2.66 $X2=0 $Y2=0
cc_44 N_A_90_94#_c_42_n N_A_M1005_g 0.00448237f $X=1.985 $Y=1.295 $X2=0 $Y2=0
cc_45 N_A_90_94#_c_37_n A 0.0225957f $X=1.755 $Y=1.295 $X2=0 $Y2=0
cc_46 N_A_90_94#_c_39_n A 0.0868643f $X=2.05 $Y=2.66 $X2=0 $Y2=0
cc_47 N_A_90_94#_c_40_n A 0.0107407f $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_48 N_A_90_94#_c_41_n A 0.0038441f $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_49 N_A_90_94#_c_42_n A 0.00336444f $X=1.985 $Y=1.295 $X2=0 $Y2=0
cc_50 N_A_90_94#_c_37_n N_A_c_98_n 4.1732e-19 $X=1.755 $Y=1.295 $X2=0 $Y2=0
cc_51 N_A_90_94#_c_39_n N_A_c_98_n 0.0255155f $X=2.05 $Y=2.66 $X2=0 $Y2=0
cc_52 N_A_90_94#_c_40_n N_A_c_98_n 8.53431e-19 $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_53 N_A_90_94#_c_41_n N_A_c_98_n 0.0172568f $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_54 N_A_90_94#_c_42_n N_A_c_98_n 0.0057222f $X=1.985 $Y=1.295 $X2=0 $Y2=0
cc_55 N_A_90_94#_M1004_g X 0.0195448f $X=0.525 $Y=0.81 $X2=0 $Y2=0
cc_56 N_A_90_94#_M1003_g X 0.0304314f $X=0.525 $Y=2.66 $X2=0 $Y2=0
cc_57 N_A_90_94#_M1001_g X 0.00239759f $X=0.885 $Y=0.81 $X2=0 $Y2=0
cc_58 N_A_90_94#_M1007_g X 0.00402045f $X=0.915 $Y=2.66 $X2=0 $Y2=0
cc_59 N_A_90_94#_c_40_n X 0.0479173f $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_60 N_A_90_94#_c_41_n X 0.025121f $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_61 N_A_90_94#_M1003_g N_VPWR_c_152_n 0.0018473f $X=0.525 $Y=2.66 $X2=0 $Y2=0
cc_62 N_A_90_94#_M1007_g N_VPWR_c_152_n 0.013015f $X=0.915 $Y=2.66 $X2=0 $Y2=0
cc_63 N_A_90_94#_c_40_n N_VPWR_c_152_n 7.37071e-19 $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_64 N_A_90_94#_M1003_g N_VPWR_c_153_n 0.00491683f $X=0.525 $Y=2.66 $X2=0 $Y2=0
cc_65 N_A_90_94#_M1007_g N_VPWR_c_153_n 0.00426961f $X=0.915 $Y=2.66 $X2=0 $Y2=0
cc_66 N_A_90_94#_c_39_n N_VPWR_c_154_n 0.00810947f $X=2.05 $Y=2.66 $X2=0 $Y2=0
cc_67 N_A_90_94#_M1003_g N_VPWR_c_151_n 0.00517496f $X=0.525 $Y=2.66 $X2=0 $Y2=0
cc_68 N_A_90_94#_M1007_g N_VPWR_c_151_n 0.00434697f $X=0.915 $Y=2.66 $X2=0 $Y2=0
cc_69 N_A_90_94#_c_39_n N_VPWR_c_151_n 0.00864691f $X=2.05 $Y=2.66 $X2=0 $Y2=0
cc_70 N_A_90_94#_M1004_g N_VGND_c_177_n 0.00155144f $X=0.525 $Y=0.81 $X2=0 $Y2=0
cc_71 N_A_90_94#_M1001_g N_VGND_c_177_n 0.0120889f $X=0.885 $Y=0.81 $X2=0 $Y2=0
cc_72 N_A_90_94#_c_37_n N_VGND_c_177_n 0.0229055f $X=1.755 $Y=1.295 $X2=0 $Y2=0
cc_73 N_A_90_94#_c_38_n N_VGND_c_177_n 0.0149529f $X=1.92 $Y=0.81 $X2=0 $Y2=0
cc_74 N_A_90_94#_c_40_n N_VGND_c_177_n 0.0047012f $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_75 N_A_90_94#_c_41_n N_VGND_c_177_n 2.34608e-19 $X=0.825 $Y=1.375 $X2=0 $Y2=0
cc_76 N_A_90_94#_M1004_g N_VGND_c_178_n 0.00371425f $X=0.525 $Y=0.81 $X2=0 $Y2=0
cc_77 N_A_90_94#_M1001_g N_VGND_c_178_n 0.00356352f $X=0.885 $Y=0.81 $X2=0 $Y2=0
cc_78 N_A_90_94#_c_38_n N_VGND_c_179_n 0.0103857f $X=1.92 $Y=0.81 $X2=0 $Y2=0
cc_79 N_A_90_94#_M1004_g N_VGND_c_180_n 0.00400172f $X=0.525 $Y=0.81 $X2=0 $Y2=0
cc_80 N_A_90_94#_M1001_g N_VGND_c_180_n 0.00400172f $X=0.885 $Y=0.81 $X2=0 $Y2=0
cc_81 N_A_90_94#_c_38_n N_VGND_c_180_n 0.014442f $X=1.92 $Y=0.81 $X2=0 $Y2=0
cc_82 N_A_M1002_g N_VPWR_c_152_n 0.00688938f $X=1.445 $Y=2.66 $X2=0 $Y2=0
cc_83 A N_VPWR_c_152_n 0.0357675f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A_M1002_g N_VPWR_c_154_n 0.00464052f $X=1.445 $Y=2.66 $X2=0 $Y2=0
cc_85 N_A_M1006_g N_VPWR_c_154_n 0.00482473f $X=1.835 $Y=2.66 $X2=0 $Y2=0
cc_86 A N_VPWR_c_154_n 0.0104923f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_VPWR_c_151_n 0.00517496f $X=1.445 $Y=2.66 $X2=0 $Y2=0
cc_88 N_A_M1006_g N_VPWR_c_151_n 0.00517496f $X=1.835 $Y=2.66 $X2=0 $Y2=0
cc_89 A N_VPWR_c_151_n 0.0113503f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_90 N_A_M1000_g N_VGND_c_177_n 0.0125894f $X=1.315 $Y=0.81 $X2=0 $Y2=0
cc_91 N_A_M1005_g N_VGND_c_177_n 0.0018473f $X=1.705 $Y=0.81 $X2=0 $Y2=0
cc_92 N_A_M1000_g N_VGND_c_179_n 0.00356352f $X=1.315 $Y=0.81 $X2=0 $Y2=0
cc_93 N_A_M1005_g N_VGND_c_179_n 0.00412501f $X=1.705 $Y=0.81 $X2=0 $Y2=0
cc_94 N_A_M1000_g N_VGND_c_180_n 0.00400172f $X=1.315 $Y=0.81 $X2=0 $Y2=0
cc_95 N_A_M1005_g N_VGND_c_180_n 0.00476395f $X=1.705 $Y=0.81 $X2=0 $Y2=0
cc_96 X N_VPWR_c_152_n 0.014639f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_97 X N_VPWR_c_153_n 0.0113158f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_98 X N_VPWR_c_151_n 0.0121101f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_99 X N_VGND_c_177_n 0.0204182f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_100 X N_VGND_c_178_n 0.0113794f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_101 X N_VGND_c_180_n 0.0121336f $X=0.155 $Y=0.47 $X2=0 $Y2=0
