* File: sky130_fd_sc_lp__fa_4.pex.spice
* Created: Fri Aug 28 10:35:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__FA_4%A 2 5 9 13 17 21 25 29 33 35 38 39 41 42 44 45
+ 46 47 48 49 51 53 54 59 60 63 64 69 70 71
c203 64 0 1.50014e-19 $X=3.99 $Y=1.65
c204 41 0 5.06513e-20 $X=1.5 $Y=2.015
c205 29 0 1.3646e-19 $X=5.535 $Y=0.865
c206 21 0 1.31942e-19 $X=3.915 $Y=0.865
c207 9 0 8.06897e-20 $X=0.525 $Y=0.865
c208 2 0 1.98052e-19 $X=0.43 $Y=1.87
r209 70 71 10.8324 $w=5.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.65
+ $X2=3.6 $Y2=1.65
r210 69 70 10.8324 $w=5.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.65
+ $X2=3.12 $Y2=1.65
r211 63 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.77
+ $X2=3.825 $Y2=1.935
r212 63 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.77
+ $X2=3.825 $Y2=1.605
r213 62 64 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.825 $Y=1.65
+ $X2=3.99 $Y2=1.65
r214 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.77 $X2=3.825 $Y2=1.77
r215 60 71 2.82094 $w=5.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.725 $Y=1.65
+ $X2=3.6 $Y2=1.65
r216 60 62 2.25675 $w=5.28e-07 $l=1e-07 $layer=LI1_cond $X=3.725 $Y=1.65
+ $X2=3.825 $Y2=1.65
r217 59 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=1.43
+ $X2=2.445 $Y2=1.595
r218 59 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=1.43
+ $X2=2.445 $Y2=1.265
r219 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.445
+ $Y=1.43 $X2=2.445 $Y2=1.43
r220 56 69 2.48243 $w=5.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.53 $Y=1.65
+ $X2=2.64 $Y2=1.65
r221 56 58 3.15432 $w=5.3e-07 $l=1.44928e-07 $layer=LI1_cond $X=2.53 $Y=1.65
+ $X2=2.412 $Y2=1.59
r222 54 85 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.625 $Y=1.51
+ $X2=5.625 $Y2=1.675
r223 54 84 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.625 $Y=1.51
+ $X2=5.625 $Y2=1.345
r224 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.625
+ $Y=1.51 $X2=5.625 $Y2=1.51
r225 51 67 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.91 $Y=1.51
+ $X2=4.91 $Y2=1.83
r226 51 53 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=4.995 $Y=1.51
+ $X2=5.625 $Y2=1.51
r227 49 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.825 $Y=1.83
+ $X2=4.91 $Y2=1.83
r228 49 64 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.825 $Y=1.83
+ $X2=3.99 $Y2=1.83
r229 47 58 6.32636 $w=1.7e-07 $l=3.40624e-07 $layer=LI1_cond $X=2.38 $Y=1.915
+ $X2=2.412 $Y2=1.59
r230 47 48 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=2.38 $Y=1.915
+ $X2=2.38 $Y2=2.895
r231 45 48 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.295 $Y=2.985
+ $X2=2.38 $Y2=2.895
r232 45 46 38.5101 $w=1.78e-07 $l=6.25e-07 $layer=LI1_cond $X=2.295 $Y=2.985
+ $X2=1.67 $Y2=2.985
r233 44 46 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.585 $Y=2.895
+ $X2=1.67 $Y2=2.985
r234 43 44 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.585 $Y=2.1
+ $X2=1.585 $Y2=2.895
r235 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.5 $Y=2.015
+ $X2=1.585 $Y2=2.1
r236 41 42 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.5 $Y=2.015
+ $X2=0.695 $Y2=2.015
r237 39 76 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.535
+ $X2=0.43 $Y2=1.37
r238 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.425
+ $Y=1.535 $X2=0.425 $Y2=1.535
r239 36 42 32.7657 $w=8e-08 $l=2.5701e-07 $layer=LI1_cond $X=0.477 $Y=1.93
+ $X2=0.695 $Y2=2.015
r240 36 38 10.4647 $w=4.33e-07 $l=3.95e-07 $layer=LI1_cond $X=0.477 $Y=1.93
+ $X2=0.477 $Y2=1.535
r241 33 85 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.535 $Y=2.415
+ $X2=5.535 $Y2=1.675
r242 29 84 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.535 $Y=0.865
+ $X2=5.535 $Y2=1.345
r243 25 82 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.915 $Y=2.415
+ $X2=3.915 $Y2=1.935
r244 21 81 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.915 $Y=0.865
+ $X2=3.915 $Y2=1.605
r245 17 79 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.51 $Y=2.415
+ $X2=2.51 $Y2=1.595
r246 13 78 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.355 $Y=0.865
+ $X2=2.355 $Y2=1.265
r247 9 76 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.525 $Y=0.865
+ $X2=0.525 $Y2=1.37
r248 5 35 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.475 $Y=2.52
+ $X2=0.475 $Y2=2.04
r249 2 35 40.8437 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=0.43 $Y=1.87
+ $X2=0.43 $Y2=2.04
r250 1 39 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=0.43 $Y=1.54 $X2=0.43
+ $Y2=1.535
r251 1 2 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=0.43 $Y=1.54 $X2=0.43
+ $Y2=1.87
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%A_328_131# 1 2 9 13 15 17 20 22 24 27 29 31 34
+ 36 38 41 45 47 49 53 56 58 59 60 61 62 65 69 71 86 87
c204 87 0 1.57905e-19 $X=9.12 $Y=1.35
c205 69 0 3.24677e-20 $X=4.56 $Y=1.295
c206 62 0 2.49488e-19 $X=4.705 $Y=1.295
c207 56 0 1.94228e-19 $X=4.365 $Y=1.48
c208 45 0 1.98692e-19 $X=1.78 $Y=0.93
r209 85 87 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=8.93 $Y=1.35
+ $X2=9.12 $Y2=1.35
r210 85 86 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.93
+ $Y=1.35 $X2=8.93 $Y2=1.35
r211 83 85 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=8.69 $Y=1.35
+ $X2=8.93 $Y2=1.35
r212 82 83 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=8.26 $Y=1.35
+ $X2=8.69 $Y2=1.35
r213 81 86 35.0893 $w=3.33e-07 $l=1.02e-06 $layer=LI1_cond $X=7.91 $Y=1.347
+ $X2=8.93 $Y2=1.347
r214 80 82 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=7.91 $Y=1.35
+ $X2=8.26 $Y2=1.35
r215 80 81 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.91
+ $Y=1.35 $X2=7.91 $Y2=1.35
r216 77 80 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=7.83 $Y=1.35 $X2=7.91
+ $Y2=1.35
r217 71 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.295
+ $X2=7.92 $Y2=1.295
r218 69 98 11.399 $w=1.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.565 $Y=1.295
+ $X2=4.565 $Y2=1.48
r219 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=1.295
+ $X2=4.56 $Y2=1.295
r220 65 95 7.80118 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=1.295
+ $X2=1.855 $Y2=1.38
r221 65 94 3.23862 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=1.295
+ $X2=1.855 $Y2=1.21
r222 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=1.295
+ $X2=1.68 $Y2=1.295
r223 62 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=1.295
+ $X2=4.56 $Y2=1.295
r224 61 71 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=1.295
+ $X2=7.92 $Y2=1.295
r225 61 62 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=7.775 $Y=1.295
+ $X2=4.705 $Y2=1.295
r226 60 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.825 $Y=1.295
+ $X2=1.68 $Y2=1.295
r227 59 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.415 $Y=1.295
+ $X2=4.56 $Y2=1.295
r228 59 60 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=4.415 $Y=1.295
+ $X2=1.825 $Y2=1.295
r229 58 95 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.03 $Y=2.055
+ $X2=2.03 $Y2=1.38
r230 56 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.365 $Y=1.48
+ $X2=4.365 $Y2=1.645
r231 56 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.365 $Y=1.48
+ $X2=4.365 $Y2=1.315
r232 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.365
+ $Y=1.48 $X2=4.365 $Y2=1.48
r233 53 98 0.384081 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=4.475 $Y=1.48
+ $X2=4.565 $Y2=1.48
r234 53 55 6.42105 $w=1.88e-07 $l=1.1e-07 $layer=LI1_cond $X=4.475 $Y=1.48
+ $X2=4.365 $Y2=1.48
r235 47 58 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=1.977 $Y=2.192
+ $X2=1.977 $Y2=2.055
r236 47 49 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=1.977 $Y=2.192
+ $X2=1.977 $Y2=2.22
r237 45 94 9.21954 $w=3.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.77 $Y=0.93
+ $X2=1.77 $Y2=1.21
r238 39 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.12 $Y=1.515
+ $X2=9.12 $Y2=1.35
r239 39 41 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.12 $Y=1.515
+ $X2=9.12 $Y2=2.465
r240 36 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.12 $Y=1.185
+ $X2=9.12 $Y2=1.35
r241 36 38 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.12 $Y=1.185
+ $X2=9.12 $Y2=0.655
r242 32 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.69 $Y=1.515
+ $X2=8.69 $Y2=1.35
r243 32 34 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.69 $Y=1.515
+ $X2=8.69 $Y2=2.465
r244 29 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.69 $Y=1.185
+ $X2=8.69 $Y2=1.35
r245 29 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.69 $Y=1.185
+ $X2=8.69 $Y2=0.655
r246 25 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.26 $Y=1.515
+ $X2=8.26 $Y2=1.35
r247 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.26 $Y=1.515
+ $X2=8.26 $Y2=2.465
r248 22 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.26 $Y=1.185
+ $X2=8.26 $Y2=1.35
r249 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.26 $Y=1.185
+ $X2=8.26 $Y2=0.655
r250 18 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.83 $Y=1.515
+ $X2=7.83 $Y2=1.35
r251 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.83 $Y=1.515
+ $X2=7.83 $Y2=2.465
r252 15 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.83 $Y=1.185
+ $X2=7.83 $Y2=1.35
r253 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.83 $Y=1.185
+ $X2=7.83 $Y2=0.655
r254 13 76 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=4.345 $Y=2.415
+ $X2=4.345 $Y2=1.645
r255 9 75 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=4.345 $Y=0.865
+ $X2=4.345 $Y2=1.315
r256 2 49 300 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=2 $X=1.64
+ $Y=2.095 $X2=1.935 $Y2=2.22
r257 1 45 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.655 $X2=1.78 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%CIN 3 5 7 11 13 15 19 21 23 24 25 26 30
c92 26 0 8.06897e-20 $X=2.16 $Y=0.555
c93 19 0 6.40318e-20 $X=4.815 $Y=0.865
c94 3 0 1.39168e-19 $X=1.565 $Y=0.865
r95 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=0.35
+ $X2=1.515 $Y2=0.515
r96 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.515
+ $Y=0.35 $X2=1.515 $Y2=0.35
r97 30 33 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.515 $Y=0.21
+ $X2=1.515 $Y2=0.35
r98 25 26 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.452
+ $X2=2.16 $Y2=0.452
r99 25 34 5.07075 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=0.452
+ $X2=1.515 $Y2=0.452
r100 24 34 9.68052 $w=3.73e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=0.452
+ $X2=1.515 $Y2=0.452
r101 19 21 794.787 $w=1.5e-07 $l=1.55e-06 $layer=POLY_cond $X=4.815 $Y=0.865
+ $X2=4.815 $Y2=2.415
r102 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.815 $Y=0.285
+ $X2=4.815 $Y2=0.865
r103 16 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.02 $Y=0.21
+ $X2=2.945 $Y2=0.21
r104 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.74 $Y=0.21
+ $X2=4.815 $Y2=0.285
r105 15 16 881.957 $w=1.5e-07 $l=1.72e-06 $layer=POLY_cond $X=4.74 $Y=0.21
+ $X2=3.02 $Y2=0.21
r106 11 13 794.787 $w=1.5e-07 $l=1.55e-06 $layer=POLY_cond $X=2.945 $Y=0.865
+ $X2=2.945 $Y2=2.415
r107 9 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.945 $Y=0.285
+ $X2=2.945 $Y2=0.21
r108 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.945 $Y=0.285
+ $X2=2.945 $Y2=0.865
r109 8 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=0.21
+ $X2=1.515 $Y2=0.21
r110 7 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.87 $Y=0.21
+ $X2=2.945 $Y2=0.21
r111 7 8 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=2.87 $Y=0.21
+ $X2=1.68 $Y2=0.21
r112 3 5 794.787 $w=1.5e-07 $l=1.55e-06 $layer=POLY_cond $X=1.565 $Y=0.865
+ $X2=1.565 $Y2=2.415
r113 3 35 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.565 $Y=0.865
+ $X2=1.565 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%B 4 7 9 10 13 18 19 23 26 27 31 34 37 39 40 41
+ 42 46
c133 42 0 1.98052e-19 $X=1.68 $Y=1.665
c134 18 0 5.06513e-20 $X=2.15 $Y=2.415
c135 7 0 1.98692e-19 $X=1.035 $Y=0.865
r136 46 49 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.017 $Y=1.665
+ $X2=1.017 $Y2=1.83
r137 46 48 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.017 $Y=1.665
+ $X2=1.017 $Y2=1.5
r138 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.04
+ $Y=1.665 $X2=1.04 $Y2=1.665
r139 41 42 25.969 $w=2.03e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.652
+ $X2=1.68 $Y2=1.652
r140 41 47 8.65632 $w=2.03e-07 $l=1.6e-07 $layer=LI1_cond $X=1.2 $Y=1.652
+ $X2=1.04 $Y2=1.652
r141 35 37 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.995 $Y=1.91
+ $X2=2.15 $Y2=1.91
r142 31 34 794.787 $w=1.5e-07 $l=1.55e-06 $layer=POLY_cond $X=5.175 $Y=0.865
+ $X2=5.175 $Y2=2.415
r143 29 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.175 $Y=3.075
+ $X2=5.175 $Y2=2.415
r144 28 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.45 $Y=3.15
+ $X2=3.375 $Y2=3.15
r145 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.1 $Y=3.15
+ $X2=5.175 $Y2=3.075
r146 27 28 846.064 $w=1.5e-07 $l=1.65e-06 $layer=POLY_cond $X=5.1 $Y=3.15
+ $X2=3.45 $Y2=3.15
r147 23 26 794.787 $w=1.5e-07 $l=1.55e-06 $layer=POLY_cond $X=3.375 $Y=0.865
+ $X2=3.375 $Y2=2.415
r148 21 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.375 $Y=3.075
+ $X2=3.375 $Y2=3.15
r149 21 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.375 $Y=3.075
+ $X2=3.375 $Y2=2.415
r150 20 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.225 $Y=3.15
+ $X2=2.15 $Y2=3.15
r151 19 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.3 $Y=3.15
+ $X2=3.375 $Y2=3.15
r152 19 20 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=3.3 $Y=3.15
+ $X2=2.225 $Y2=3.15
r153 16 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.15 $Y=3.075
+ $X2=2.15 $Y2=3.15
r154 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=3.075
+ $X2=2.15 $Y2=2.415
r155 15 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.15 $Y=1.985
+ $X2=2.15 $Y2=1.91
r156 15 18 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.15 $Y=1.985
+ $X2=2.15 $Y2=2.415
r157 11 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.995 $Y=1.835
+ $X2=1.995 $Y2=1.91
r158 11 13 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=1.995 $Y=1.835
+ $X2=1.995 $Y2=0.865
r159 9 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.075 $Y=3.15
+ $X2=2.15 $Y2=3.15
r160 9 10 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=2.075 $Y=3.15
+ $X2=0.98 $Y2=3.15
r161 7 48 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.035 $Y=0.865
+ $X2=1.035 $Y2=1.5
r162 4 49 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.905 $Y=2.52
+ $X2=0.905 $Y2=1.83
r163 2 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=3.075
+ $X2=0.98 $Y2=3.15
r164 2 4 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.905 $Y=3.075
+ $X2=0.905 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%A_884_131# 1 2 9 13 17 21 25 29 33 37 41 45 48
+ 50 56 60 61 68
c134 60 0 6.40318e-20 $X=4.58 $Y=2.26
c135 41 0 1.94228e-19 $X=5.89 $Y=0.865
r136 67 68 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.97 $Y=1.48
+ $X2=7.4 $Y2=1.48
r137 57 67 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.88 $Y=1.48 $X2=6.97
+ $Y2=1.48
r138 57 65 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.88 $Y=1.48
+ $X2=6.54 $Y2=1.48
r139 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=1.48 $X2=6.88 $Y2=1.48
r140 54 65 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.2 $Y=1.48
+ $X2=6.54 $Y2=1.48
r141 54 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.2 $Y=1.48 $X2=6.11
+ $Y2=1.48
r142 53 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.2 $Y=1.48
+ $X2=6.88 $Y2=1.48
r143 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.2
+ $Y=1.48 $X2=6.2 $Y2=1.48
r144 51 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.06 $Y=1.48
+ $X2=5.975 $Y2=1.48
r145 51 53 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.06 $Y=1.48
+ $X2=6.2 $Y2=1.48
r146 49 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.975 $Y=1.565
+ $X2=5.975 $Y2=1.48
r147 49 50 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.975 $Y=1.565
+ $X2=5.975 $Y2=2.095
r148 48 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.975 $Y=1.395
+ $X2=5.975 $Y2=1.48
r149 47 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.975 $Y=1.03
+ $X2=5.975 $Y2=1.395
r150 46 60 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=4.745 $Y=2.18
+ $X2=4.587 $Y2=2.18
r151 45 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.89 $Y=2.18
+ $X2=5.975 $Y2=2.095
r152 45 46 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=5.89 $Y=2.18
+ $X2=4.745 $Y2=2.18
r153 41 47 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.89 $Y=0.865
+ $X2=5.975 $Y2=1.03
r154 41 43 45.05 $w=3.28e-07 $l=1.29e-06 $layer=LI1_cond $X=5.89 $Y=0.865
+ $X2=4.6 $Y2=0.865
r155 35 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.4 $Y=1.645
+ $X2=7.4 $Y2=1.48
r156 35 37 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.4 $Y=1.645
+ $X2=7.4 $Y2=2.465
r157 31 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.4 $Y=1.315
+ $X2=7.4 $Y2=1.48
r158 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.4 $Y=1.315
+ $X2=7.4 $Y2=0.655
r159 27 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=1.645
+ $X2=6.97 $Y2=1.48
r160 27 29 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.97 $Y=1.645
+ $X2=6.97 $Y2=2.465
r161 23 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.97 $Y=1.315
+ $X2=6.97 $Y2=1.48
r162 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.97 $Y=1.315
+ $X2=6.97 $Y2=0.655
r163 19 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.54 $Y=1.645
+ $X2=6.54 $Y2=1.48
r164 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.54 $Y=1.645
+ $X2=6.54 $Y2=2.465
r165 15 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.54 $Y=1.315
+ $X2=6.54 $Y2=1.48
r166 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.54 $Y=1.315
+ $X2=6.54 $Y2=0.655
r167 11 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.11 $Y=1.645
+ $X2=6.11 $Y2=1.48
r168 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.11 $Y=1.645
+ $X2=6.11 $Y2=2.465
r169 7 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.11 $Y=1.315
+ $X2=6.11 $Y2=1.48
r170 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.11 $Y=1.315
+ $X2=6.11 $Y2=0.655
r171 2 60 300 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=2.095 $X2=4.58 $Y2=2.26
r172 1 43 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.655 $X2=4.6 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%A_27_440# 1 2 7 9 11 15
r24 15 18 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.215 $Y=2.365
+ $X2=1.215 $Y2=2.445
r25 12 14 4.01803 $w=1.7e-07 $l=1.52971e-07 $layer=LI1_cond $X=0.355 $Y=2.365
+ $X2=0.225 $Y2=2.315
r26 11 15 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.11 $Y=2.365
+ $X2=1.215 $Y2=2.365
r27 11 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.11 $Y=2.365
+ $X2=0.355 $Y2=2.365
r28 7 14 3.12513 $w=2.5e-07 $l=1.37477e-07 $layer=LI1_cond $X=0.22 $Y=2.45
+ $X2=0.225 $Y2=2.315
r29 7 9 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=0.22 $Y=2.45 $X2=0.22
+ $Y2=2.685
r30 2 18 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.2 $X2=1.215 $Y2=2.445
r31 1 14 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.2 $X2=0.26 $Y2=2.345
r32 1 9 600 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.2 $X2=0.26 $Y2=2.685
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 45 51 57 61 63
+ 68 69 71 72 74 75 76 78 83 88 106 110 116 119 122 125 129
c141 129 0 6.50762e-20 $X=9.36 $Y=3.33
r142 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r143 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r144 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r145 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r146 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 114 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r148 114 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r149 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r150 111 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.64 $Y=3.33
+ $X2=8.475 $Y2=3.33
r151 111 113 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.64 $Y=3.33
+ $X2=8.88 $Y2=3.33
r152 110 128 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=9.17 $Y=3.33
+ $X2=9.385 $Y2=3.33
r153 110 113 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.17 $Y=3.33
+ $X2=8.88 $Y2=3.33
r154 109 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r156 106 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.31 $Y=3.33
+ $X2=8.475 $Y2=3.33
r157 106 108 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.31 $Y=3.33
+ $X2=7.92 $Y2=3.33
r158 105 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r159 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r160 102 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r161 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r162 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r163 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r164 96 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r165 95 98 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.52 $Y2=3.33
r166 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r167 93 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=3.33
+ $X2=3.645 $Y2=3.33
r168 93 95 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.81 $Y=3.33
+ $X2=4.08 $Y2=3.33
r169 92 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r170 92 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r171 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r172 89 119 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.745 $Y2=3.33
r173 89 91 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.12 $Y2=3.33
r174 88 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.48 $Y=3.33
+ $X2=3.645 $Y2=3.33
r175 88 91 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.48 $Y=3.33
+ $X2=3.12 $Y2=3.33
r176 87 120 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r177 87 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r178 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r179 84 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r180 84 86 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r181 83 119 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.745 $Y2=3.33
r182 83 86 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=1.2 $Y2=3.33
r183 81 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r184 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r185 78 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r186 78 80 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r187 76 99 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.52 $Y2=3.33
r188 76 96 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.08 $Y2=3.33
r189 74 104 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=7.45 $Y=3.33
+ $X2=7.44 $Y2=3.33
r190 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=3.33
+ $X2=7.615 $Y2=3.33
r191 73 108 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=7.78 $Y=3.33
+ $X2=7.92 $Y2=3.33
r192 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.78 $Y=3.33
+ $X2=7.615 $Y2=3.33
r193 71 101 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.59 $Y=3.33
+ $X2=6.48 $Y2=3.33
r194 71 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.59 $Y=3.33
+ $X2=6.755 $Y2=3.33
r195 70 104 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r196 70 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.92 $Y=3.33
+ $X2=6.755 $Y2=3.33
r197 68 98 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r198 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.895 $Y2=3.33
r199 67 101 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=6.48 $Y2=3.33
r200 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.06 $Y=3.33
+ $X2=5.895 $Y2=3.33
r201 63 66 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=9.335 $Y=2.19
+ $X2=9.335 $Y2=2.95
r202 61 128 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=9.335 $Y=3.245
+ $X2=9.385 $Y2=3.33
r203 61 66 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.335 $Y=3.245
+ $X2=9.335 $Y2=2.95
r204 57 60 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=8.475 $Y=2.19
+ $X2=8.475 $Y2=2.95
r205 55 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.475 $Y=3.245
+ $X2=8.475 $Y2=3.33
r206 55 60 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.475 $Y=3.245
+ $X2=8.475 $Y2=2.95
r207 51 54 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=7.615 $Y=2.19
+ $X2=7.615 $Y2=2.95
r208 49 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.615 $Y=3.245
+ $X2=7.615 $Y2=3.33
r209 49 54 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.615 $Y=3.245
+ $X2=7.615 $Y2=2.95
r210 45 48 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=6.755 $Y=2.19
+ $X2=6.755 $Y2=2.95
r211 43 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=3.245
+ $X2=6.755 $Y2=3.33
r212 43 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.755 $Y=3.245
+ $X2=6.755 $Y2=2.95
r213 39 42 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=5.895 $Y=2.535
+ $X2=5.895 $Y2=2.95
r214 37 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.895 $Y=3.245
+ $X2=5.895 $Y2=3.33
r215 37 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.895 $Y=3.245
+ $X2=5.895 $Y2=2.95
r216 33 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=3.245
+ $X2=3.645 $Y2=3.33
r217 33 35 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=3.645 $Y=3.245
+ $X2=3.645 $Y2=2.56
r218 29 119 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=3.245
+ $X2=2.745 $Y2=3.33
r219 29 31 51.0742 $w=2.18e-07 $l=9.75e-07 $layer=LI1_cond $X=2.745 $Y=3.245
+ $X2=2.745 $Y2=2.27
r220 25 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r221 25 27 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.715
r222 8 66 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.195
+ $Y=1.835 $X2=9.335 $Y2=2.95
r223 8 63 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=9.195
+ $Y=1.835 $X2=9.335 $Y2=2.19
r224 7 60 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=1.835 $X2=8.475 $Y2=2.95
r225 7 57 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=1.835 $X2=8.475 $Y2=2.19
r226 6 54 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.475
+ $Y=1.835 $X2=7.615 $Y2=2.95
r227 6 51 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=7.475
+ $Y=1.835 $X2=7.615 $Y2=2.19
r228 5 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.615
+ $Y=1.835 $X2=6.755 $Y2=2.95
r229 5 45 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=6.615
+ $Y=1.835 $X2=6.755 $Y2=2.19
r230 4 42 600 $w=1.7e-07 $l=9.87269e-07 $layer=licon1_PDIFF $count=1 $X=5.61
+ $Y=2.095 $X2=5.895 $Y2=2.95
r231 4 39 600 $w=1.7e-07 $l=5.64801e-07 $layer=licon1_PDIFF $count=1 $X=5.61
+ $Y=2.095 $X2=5.895 $Y2=2.535
r232 3 35 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=2.095 $X2=3.645 $Y2=2.56
r233 2 31 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=2.585
+ $Y=2.095 $X2=2.73 $Y2=2.27
r234 1 27 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.2 $X2=0.69 $Y2=2.715
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%A_604_419# 1 2 9 14 16
r25 10 14 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.275 $Y=2.18
+ $X2=3.15 $Y2=2.18
r26 9 16 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.98 $Y=2.18 $X2=4.12
+ $Y2=2.18
r27 9 10 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.98 $Y=2.18
+ $X2=3.275 $Y2=2.18
r28 2 16 300 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.095 $X2=4.13 $Y2=2.26
r29 1 14 300 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=2 $X=3.02
+ $Y=2.095 $X2=3.16 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%SUM 1 2 3 4 15 19 23 24 25 26 29 33 38 39 45
c64 38 0 1.57905e-19 $X=7.332 $Y=1.135
r65 42 45 2.24086 $w=3.58e-07 $l=7e-08 $layer=LI1_cond $X=7.395 $Y=1.735
+ $X2=7.395 $Y2=1.665
r66 39 42 3.75991 $w=2.75e-07 $l=1.22515e-07 $layer=LI1_cond $X=7.332 $Y=1.83
+ $X2=7.395 $Y2=1.735
r67 39 45 0.256098 $w=3.58e-07 $l=8e-09 $layer=LI1_cond $X=7.395 $Y=1.657
+ $X2=7.395 $Y2=1.665
r68 37 39 13.8293 $w=3.58e-07 $l=4.32e-07 $layer=LI1_cond $X=7.395 $Y=1.225
+ $X2=7.395 $Y2=1.657
r69 37 38 3.58391 $w=2.75e-07 $l=1.17346e-07 $layer=LI1_cond $X=7.395 $Y=1.225
+ $X2=7.332 $Y2=1.135
r70 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=7.185 $Y=1.98
+ $X2=7.185 $Y2=2.91
r71 31 39 3.75991 $w=2.75e-07 $l=1.88611e-07 $layer=LI1_cond $X=7.185 $Y=1.925
+ $X2=7.332 $Y2=1.83
r72 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=7.185 $Y=1.925
+ $X2=7.185 $Y2=1.98
r73 27 38 3.58391 $w=2.75e-07 $l=1.86652e-07 $layer=LI1_cond $X=7.185 $Y=1.045
+ $X2=7.332 $Y2=1.135
r74 27 29 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=7.185 $Y=1.045
+ $X2=7.185 $Y2=0.42
r75 25 39 2.70212 $w=1.9e-07 $l=2.42e-07 $layer=LI1_cond $X=7.09 $Y=1.83
+ $X2=7.332 $Y2=1.83
r76 25 26 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=7.09 $Y=1.83 $X2=6.42
+ $Y2=1.83
r77 23 38 2.90466 $w=1.8e-07 $l=2.42e-07 $layer=LI1_cond $X=7.09 $Y=1.135
+ $X2=7.332 $Y2=1.135
r78 23 24 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.09 $Y=1.135
+ $X2=6.42 $Y2=1.135
r79 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.325 $Y=1.98
+ $X2=6.325 $Y2=2.91
r80 17 26 6.81649 $w=1.9e-07 $l=1.3435e-07 $layer=LI1_cond $X=6.325 $Y=1.925
+ $X2=6.42 $Y2=1.83
r81 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.325 $Y=1.925
+ $X2=6.325 $Y2=1.98
r82 13 24 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=6.325 $Y=1.045
+ $X2=6.42 $Y2=1.135
r83 13 15 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=6.325 $Y=1.045
+ $X2=6.325 $Y2=0.42
r84 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=1.835 $X2=7.185 $Y2=2.91
r85 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=1.835 $X2=7.185 $Y2=1.98
r86 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.185
+ $Y=1.835 $X2=6.325 $Y2=2.91
r87 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.185
+ $Y=1.835 $X2=6.325 $Y2=1.98
r88 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.045
+ $Y=0.235 $X2=7.185 $Y2=0.42
r89 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.185
+ $Y=0.235 $X2=6.325 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%COUT 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41
+ 42 44 45 46
r59 45 46 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=9.387 $Y=1.295
+ $X2=9.387 $Y2=1.665
r60 44 45 9.83236 $w=4.13e-07 $l=2.85e-07 $layer=LI1_cond $X=9.387 $Y=1.01
+ $X2=9.387 $Y2=1.295
r61 43 46 4.23346 $w=2.43e-07 $l=9e-08 $layer=LI1_cond $X=9.387 $Y=1.755
+ $X2=9.387 $Y2=1.665
r62 40 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9 $Y=1.84 $X2=8.905
+ $Y2=1.84
r63 39 43 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=9.265 $Y=1.84
+ $X2=9.387 $Y2=1.755
r64 39 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.265 $Y=1.84 $X2=9
+ $Y2=1.84
r65 38 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9 $Y=0.925 $X2=8.905
+ $Y2=0.925
r66 37 44 4.1905 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=9.265 $Y=0.925
+ $X2=9.387 $Y2=0.925
r67 37 38 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.265 $Y=0.925
+ $X2=9 $Y2=0.925
r68 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=8.905 $Y=1.98
+ $X2=8.905 $Y2=2.91
r69 31 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=1.925
+ $X2=8.905 $Y2=1.84
r70 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=8.905 $Y=1.925
+ $X2=8.905 $Y2=1.98
r71 27 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=0.84
+ $X2=8.905 $Y2=0.925
r72 27 29 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=8.905 $Y=0.84
+ $X2=8.905 $Y2=0.42
r73 25 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.81 $Y=1.84
+ $X2=8.905 $Y2=1.84
r74 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.81 $Y=1.84
+ $X2=8.14 $Y2=1.84
r75 23 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.81 $Y=0.925
+ $X2=8.905 $Y2=0.925
r76 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.81 $Y=0.925
+ $X2=8.14 $Y2=0.925
r77 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=8.045 $Y=1.98
+ $X2=8.045 $Y2=2.91
r78 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.045 $Y=1.925
+ $X2=8.14 $Y2=1.84
r79 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=8.045 $Y=1.925
+ $X2=8.045 $Y2=1.98
r80 13 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.045 $Y=0.84
+ $X2=8.14 $Y2=0.925
r81 13 15 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=8.045 $Y=0.84
+ $X2=8.045 $Y2=0.42
r82 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.765
+ $Y=1.835 $X2=8.905 $Y2=2.91
r83 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.765
+ $Y=1.835 $X2=8.905 $Y2=1.98
r84 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.905
+ $Y=1.835 $X2=8.045 $Y2=2.91
r85 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.905
+ $Y=1.835 $X2=8.045 $Y2=1.98
r86 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.765
+ $Y=0.235 $X2=8.905 $Y2=0.42
r87 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.905
+ $Y=0.235 $X2=8.045 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%A_37_131# 1 2 9 11 12 14
r25 14 16 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.25 $Y=0.93
+ $X2=1.25 $Y2=1.15
r26 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=1.15
+ $X2=1.25 $Y2=1.15
r27 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.085 $Y=1.15
+ $X2=0.405 $Y2=1.15
r28 7 12 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.305 $Y=1.065
+ $X2=0.405 $Y2=1.15
r29 7 9 10.8136 $w=1.98e-07 $l=1.95e-07 $layer=LI1_cond $X=0.305 $Y=1.065
+ $X2=0.305 $Y2=0.87
r30 2 14 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.11
+ $Y=0.655 $X2=1.25 $Y2=0.93
r31 1 9 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.655 $X2=0.31 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51 53 55
+ 58 59 61 62 64 65 66 68 73 81 99 103 109 112 115 118 122
c138 39 0 1.3646e-19 $X=5.875 $Y=0.415
c139 27 0 7.40916e-20 $X=0.74 $Y=0.78
r140 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r141 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r142 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r143 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r144 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r145 107 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r146 107 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=8.4 $Y2=0
r147 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r148 104 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.64 $Y=0
+ $X2=8.475 $Y2=0
r149 104 106 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=8.64 $Y=0
+ $X2=8.88 $Y2=0
r150 103 121 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=9.17 $Y=0
+ $X2=9.385 $Y2=0
r151 103 106 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.17 $Y=0
+ $X2=8.88 $Y2=0
r152 102 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r153 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r154 99 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.31 $Y=0
+ $X2=8.475 $Y2=0
r155 99 101 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.31 $Y=0 $X2=7.92
+ $Y2=0
r156 98 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r157 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r158 95 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r159 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r160 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r161 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r162 89 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r163 88 91 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r164 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r165 86 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.775 $Y=0
+ $X2=3.61 $Y2=0
r166 86 88 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.775 $Y=0
+ $X2=4.08 $Y2=0
r167 85 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r168 85 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=2.64 $Y2=0
r169 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r170 82 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0
+ $X2=2.59 $Y2=0
r171 82 84 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=0
+ $X2=3.12 $Y2=0
r172 81 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=0
+ $X2=3.61 $Y2=0
r173 81 84 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.445 $Y=0
+ $X2=3.12 $Y2=0
r174 80 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r175 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r176 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r177 77 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r178 76 79 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r179 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r180 74 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.74 $Y2=0
r181 74 76 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.2
+ $Y2=0
r182 73 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=0
+ $X2=2.59 $Y2=0
r183 73 79 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.425 $Y=0
+ $X2=2.16 $Y2=0
r184 71 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r185 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r186 68 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0
+ $X2=0.74 $Y2=0
r187 68 70 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0
+ $X2=0.24 $Y2=0
r188 66 92 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.52
+ $Y2=0
r189 66 89 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.08
+ $Y2=0
r190 64 97 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=7.45 $Y=0 $X2=7.44
+ $Y2=0
r191 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=0 $X2=7.615
+ $Y2=0
r192 63 101 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=7.78 $Y=0 $X2=7.92
+ $Y2=0
r193 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.78 $Y=0 $X2=7.615
+ $Y2=0
r194 61 94 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.59 $Y=0 $X2=6.48
+ $Y2=0
r195 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.59 $Y=0 $X2=6.755
+ $Y2=0
r196 60 97 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.92 $Y=0 $X2=7.44
+ $Y2=0
r197 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.92 $Y=0 $X2=6.755
+ $Y2=0
r198 58 91 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.71 $Y=0 $X2=5.52
+ $Y2=0
r199 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.71 $Y=0 $X2=5.875
+ $Y2=0
r200 57 94 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.04 $Y=0 $X2=6.48
+ $Y2=0
r201 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.04 $Y=0 $X2=5.875
+ $Y2=0
r202 53 121 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=9.335 $Y=0.085
+ $X2=9.385 $Y2=0
r203 53 55 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=9.335 $Y=0.085
+ $X2=9.335 $Y2=0.53
r204 49 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.475 $Y=0.085
+ $X2=8.475 $Y2=0
r205 49 51 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.475 $Y=0.085
+ $X2=8.475 $Y2=0.53
r206 45 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.615 $Y=0.085
+ $X2=7.615 $Y2=0
r207 45 47 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.615 $Y=0.085
+ $X2=7.615 $Y2=0.36
r208 41 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=0.085
+ $X2=6.755 $Y2=0
r209 41 43 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0.085
+ $X2=6.755 $Y2=0.36
r210 37 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=0.085
+ $X2=5.875 $Y2=0
r211 37 39 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.875 $Y=0.085
+ $X2=5.875 $Y2=0.415
r212 33 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.61 $Y=0.085
+ $X2=3.61 $Y2=0
r213 33 35 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.61 $Y=0.085
+ $X2=3.61 $Y2=0.78
r214 29 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0
r215 29 31 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0.875
r216 25 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r217 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.78
r218 8 55 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=9.195
+ $Y=0.235 $X2=9.335 $Y2=0.53
r219 7 51 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=8.335
+ $Y=0.235 $X2=8.475 $Y2=0.53
r220 6 47 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.475
+ $Y=0.235 $X2=7.615 $Y2=0.36
r221 5 43 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.615
+ $Y=0.235 $X2=6.755 $Y2=0.36
r222 4 39 182 $w=1.7e-07 $l=3.65821e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.655 $X2=5.875 $Y2=0.415
r223 3 35 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.655 $X2=3.61 $Y2=0.78
r224 2 31 182 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.655 $X2=2.59 $Y2=0.875
r225 1 27 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.655 $X2=0.74 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__FA_4%A_604_131# 1 2 9 11 12 15
r22 13 15 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=4.13 $Y=1.045
+ $X2=4.13 $Y2=0.93
r23 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.025 $Y=1.13
+ $X2=4.13 $Y2=1.045
r24 11 12 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.025 $Y=1.13
+ $X2=3.265 $Y2=1.13
r25 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.16 $Y=1.045
+ $X2=3.265 $Y2=1.13
r26 7 9 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=3.16 $Y=1.045
+ $X2=3.16 $Y2=0.93
r27 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.655 $X2=4.13 $Y2=0.93
r28 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.655 $X2=3.16 $Y2=0.93
.ends

