* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o211a_0 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 VGND A2 a_257_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_257_47# B1 a_520_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR A1 a_340_485# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_520_47# C1 a_80_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_257_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_340_485# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
