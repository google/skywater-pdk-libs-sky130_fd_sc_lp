* File: sky130_fd_sc_lp__o211a_2.pex.spice
* Created: Wed Sep  2 10:13:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211A_2%C1 3 5 7 8 13
c26 13 0 1.36063e-19 $X=0.475 $Y=1.485
c27 3 0 2.2534e-19 $X=0.475 $Y=0.655
r28 11 13 25.4665 $w=3.88e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.485
+ $X2=0.475 $Y2=1.485
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.41 $X2=0.27 $Y2=1.41
r30 8 12 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.41
r31 5 13 21.1186 $w=3.88e-07 $l=3.13688e-07 $layer=POLY_cond $X=0.645 $Y=1.725
+ $X2=0.475 $Y2=1.485
r32 5 7 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.645 $Y=1.725
+ $X2=0.645 $Y2=2.465
r33 1 13 25.1189 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.475 $Y=1.245
+ $X2=0.475 $Y2=1.485
r34 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.475 $Y=1.245
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_2%B1 1 3 6 8 12
c36 8 0 2.94736e-19 $X=1.2 $Y=1.295
r37 12 14 3.59701 $w=2.68e-07 $l=2e-08 $layer=POLY_cond $X=1.095 $Y=1.35
+ $X2=1.115 $Y2=1.35
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.35 $X2=1.095 $Y2=1.35
r39 8 13 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.34 $X2=1.095
+ $Y2=1.34
r40 4 14 16.3317 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.515
+ $X2=1.115 $Y2=1.35
r41 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.115 $Y=1.515
+ $X2=1.115 $Y2=2.465
r42 1 12 46.7612 $w=2.68e-07 $l=3.32415e-07 $layer=POLY_cond $X=0.835 $Y=1.185
+ $X2=1.095 $Y2=1.35
r43 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.835 $Y=1.185
+ $X2=0.835 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_2%A2 1 3 4 6 8 9 10
c43 8 0 1.911e-20 $X=1.68 $Y=1.295
c44 1 0 6.50375e-20 $X=1.785 $Y=1.23
r45 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.395 $X2=1.68 $Y2=1.395
r46 9 10 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=2.035
r47 9 16 14.1436 $w=2.18e-07 $l=2.7e-07 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=1.395
r48 8 16 5.23838 $w=2.18e-07 $l=1e-07 $layer=LI1_cond $X=1.705 $Y=1.295
+ $X2=1.705 $Y2=1.395
r49 4 15 49.2895 $w=3.89e-07 $l=2.9904e-07 $layer=POLY_cond $X=1.785 $Y=1.64
+ $X2=1.665 $Y2=1.395
r50 4 6 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=1.785 $Y=1.64
+ $X2=1.785 $Y2=2.465
r51 1 15 39.3769 $w=3.89e-07 $l=2.16852e-07 $layer=POLY_cond $X=1.785 $Y=1.23
+ $X2=1.665 $Y2=1.395
r52 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.785 $Y=1.23
+ $X2=1.785 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_2%A1 3 7 8 9 10 15 17
c38 17 0 1.911e-20 $X=2.235 $Y=1.23
c39 15 0 3.23284e-20 $X=2.235 $Y=1.395
c40 3 0 1.95222e-19 $X=2.145 $Y=2.465
r41 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.395
+ $X2=2.235 $Y2=1.56
r42 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.395
+ $X2=2.235 $Y2=1.23
r43 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.395 $X2=2.235 $Y2=1.395
r44 9 10 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.172 $Y=1.665
+ $X2=2.172 $Y2=2.035
r45 9 16 10.5478 $w=2.93e-07 $l=2.7e-07 $layer=LI1_cond $X=2.172 $Y=1.665
+ $X2=2.172 $Y2=1.395
r46 8 16 3.90659 $w=2.93e-07 $l=1e-07 $layer=LI1_cond $X=2.172 $Y=1.295
+ $X2=2.172 $Y2=1.395
r47 7 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.215 $Y=0.7
+ $X2=2.215 $Y2=1.23
r48 3 18 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=2.145 $Y=2.465
+ $X2=2.145 $Y2=1.56
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_2%A_27_47# 1 2 3 12 16 20 24 28 32 37 38 43 46
+ 49 52 54 56 60 66
c109 60 0 1.95222e-19 $X=2.775 $Y=1.46
r110 65 66 29.0361 $w=3.32e-07 $l=2e-07 $layer=POLY_cond $X=2.915 $Y=1.462
+ $X2=3.115 $Y2=1.462
r111 61 65 20.3253 $w=3.32e-07 $l=1.4e-07 $layer=POLY_cond $X=2.775 $Y=1.462
+ $X2=2.915 $Y2=1.462
r112 61 63 13.0663 $w=3.32e-07 $l=9e-08 $layer=POLY_cond $X=2.775 $Y=1.462
+ $X2=2.685 $Y2=1.462
r113 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.775
+ $Y=1.46 $X2=2.775 $Y2=1.46
r114 57 60 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.575 $Y=1.46
+ $X2=2.775 $Y2=1.46
r115 48 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=1.625
+ $X2=2.575 $Y2=1.46
r116 48 49 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.575 $Y=1.625
+ $X2=2.575 $Y2=2.29
r117 47 56 3.51065 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.615 $Y=2.375
+ $X2=1.415 $Y2=2.375
r118 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.49 $Y=2.375
+ $X2=2.575 $Y2=2.29
r119 46 47 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.49 $Y=2.375
+ $X2=1.615 $Y2=2.375
r120 41 56 3.10218 $w=3.05e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.32 $Y=2.29
+ $X2=1.415 $Y2=2.375
r121 41 43 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=1.32 $Y=2.29
+ $X2=1.32 $Y2=1.98
r122 40 43 3.4329 $w=2.08e-07 $l=6.5e-08 $layer=LI1_cond $X=1.32 $Y=1.915
+ $X2=1.32 $Y2=1.98
r123 39 54 0.70772 $w=2.75e-07 $l=4.55719e-07 $layer=LI1_cond $X=0.705 $Y=1.777
+ $X2=0.265 $Y2=1.745
r124 38 40 6.97695 $w=2.75e-07 $l=1.83123e-07 $layer=LI1_cond $X=1.215 $Y=1.777
+ $X2=1.32 $Y2=1.915
r125 38 39 21.3726 $w=2.73e-07 $l=5.1e-07 $layer=LI1_cond $X=1.215 $Y=1.777
+ $X2=0.705 $Y2=1.777
r126 37 54 5.97828 $w=2.3e-07 $l=3.99061e-07 $layer=LI1_cond $X=0.615 $Y=1.64
+ $X2=0.265 $Y2=1.745
r127 36 52 0.716491 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=0.615 $Y=1.04
+ $X2=0.615 $Y2=0.95
r128 36 37 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=0.615 $Y=1.04
+ $X2=0.615 $Y2=1.64
r129 32 34 38.2776 $w=2.78e-07 $l=9.3e-07 $layer=LI1_cond $X=0.405 $Y=1.98
+ $X2=0.405 $Y2=2.91
r130 30 54 5.97828 $w=2.3e-07 $l=2.29565e-07 $layer=LI1_cond $X=0.405 $Y=1.915
+ $X2=0.265 $Y2=1.745
r131 30 32 2.67531 $w=2.78e-07 $l=6.5e-08 $layer=LI1_cond $X=0.405 $Y=1.915
+ $X2=0.405 $Y2=1.98
r132 26 52 21.8737 $w=1.78e-07 $l=3.55e-07 $layer=LI1_cond $X=0.26 $Y=0.95
+ $X2=0.615 $Y2=0.95
r133 26 28 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.26 $Y=0.86
+ $X2=0.26 $Y2=0.38
r134 22 66 33.3916 $w=3.32e-07 $l=2.3e-07 $layer=POLY_cond $X=3.345 $Y=1.462
+ $X2=3.115 $Y2=1.462
r135 22 24 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.345 $Y=1.625
+ $X2=3.345 $Y2=2.465
r136 18 66 21.3668 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=3.115 $Y=1.295
+ $X2=3.115 $Y2=1.462
r137 18 20 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=3.115 $Y=1.295
+ $X2=3.115 $Y2=0.7
r138 14 65 21.3668 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=2.915 $Y=1.63
+ $X2=2.915 $Y2=1.462
r139 14 16 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=2.915 $Y=1.63
+ $X2=2.915 $Y2=2.465
r140 10 63 21.3668 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=2.685 $Y=1.295
+ $X2=2.685 $Y2=1.462
r141 10 12 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=2.685 $Y=1.295
+ $X2=2.685 $Y2=0.7
r142 3 56 300 $w=1.7e-07 $l=7.1325e-07 $layer=licon1_PDIFF $count=2 $X=1.19
+ $Y=1.835 $X2=1.45 $Y2=2.43
r143 3 43 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.19
+ $Y=1.835 $X2=1.33 $Y2=1.98
r144 2 34 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.835 $X2=0.43 $Y2=2.91
r145 2 32 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.835 $X2=0.43 $Y2=1.98
r146 1 28 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_2%VPWR 1 2 3 14 18 20 22 24 32 38 41 49
r50 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r51 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 41 44 10.2649 $w=6.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.53 $Y=2.755
+ $X2=2.53 $Y2=3.33
r53 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 36 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r55 36 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 33 44 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=2.53 $Y2=3.33
r58 33 35 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 32 48 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.617 $Y2=3.33
r60 32 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r65 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 25 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=0.88 $Y2=3.33
r67 25 27 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 24 44 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.53 $Y2=3.33
r69 24 30 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 22 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 22 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r72 18 48 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.617 $Y2=3.33
r73 18 20 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=2.395
r74 14 17 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.88 $Y=2.17
+ $X2=0.88 $Y2=2.95
r75 12 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=3.33
r76 12 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.88 $Y=3.245
+ $X2=0.88 $Y2=2.95
r77 3 20 300 $w=1.7e-07 $l=6.26099e-07 $layer=licon1_PDIFF $count=2 $X=3.42
+ $Y=1.835 $X2=3.56 $Y2=2.395
r78 2 41 300 $w=1.7e-07 $l=1.1349e-06 $layer=licon1_PDIFF $count=2 $X=2.22
+ $Y=1.835 $X2=2.7 $Y2=2.755
r79 1 17 400 $w=1.7e-07 $l=1.19232e-06 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.835 $X2=0.88 $Y2=2.95
r80 1 14 400 $w=1.7e-07 $l=4.07216e-07 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.835 $X2=0.88 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_2%X 1 2 9 13 19 20 21
c27 19 0 3.23284e-20 $X=3.12 $Y=1.295
r28 21 27 3.07563 $w=4.53e-07 $l=1.17e-07 $layer=LI1_cond $X=3.257 $Y=2.01
+ $X2=3.257 $Y2=1.893
r29 20 27 5.99354 $w=4.53e-07 $l=2.28e-07 $layer=LI1_cond $X=3.257 $Y=1.665
+ $X2=3.257 $Y2=1.893
r30 20 26 4.94204 $w=4.53e-07 $l=1.88e-07 $layer=LI1_cond $X=3.257 $Y=1.665
+ $X2=3.257 $Y2=1.477
r31 19 26 6.12234 $w=2.73e-07 $l=3.22301e-07 $layer=LI1_cond $X=3.12 $Y=1.216
+ $X2=3.257 $Y2=1.477
r32 17 18 1.70629 $w=1.93e-07 $l=3e-08 $layer=LI1_cond $X=3.127 $Y=2.43
+ $X2=3.127 $Y2=2.46
r33 15 21 8.9683 $w=3.63e-07 $l=2.43e-07 $layer=LI1_cond $X=3.127 $Y=2.363
+ $X2=3.127 $Y2=2.12
r34 15 17 3.81072 $w=1.93e-07 $l=6.7e-08 $layer=LI1_cond $X=3.127 $Y=2.363
+ $X2=3.127 $Y2=2.43
r35 13 18 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=3.13 $Y=2.91
+ $X2=3.13 $Y2=2.46
r36 7 19 9.8315 $w=2.73e-07 $l=3.54318e-07 $layer=LI1_cond $X=2.9 $Y=0.955
+ $X2=3.12 $Y2=1.216
r37 7 9 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=2.9 $Y=0.955 $X2=2.9
+ $Y2=0.42
r38 2 21 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.835 $X2=3.13 $Y2=2.01
r39 2 17 600 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.835 $X2=3.13 $Y2=2.43
r40 2 13 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.835 $X2=3.13 $Y2=2.91
r41 1 9 91 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=2 $X=2.76 $Y=0.28
+ $X2=2.9 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_2%A_182_47# 1 2 9 11 12 13 15
c33 12 0 1.31705e-19 $X=1.215 $Y=0.955
r34 13 18 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=0.87
+ $X2=2.035 $Y2=0.955
r35 13 15 19.2813 $w=2.58e-07 $l=4.35e-07 $layer=LI1_cond $X=2.035 $Y=0.87
+ $X2=2.035 $Y2=0.435
r36 11 18 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.905 $Y=0.955
+ $X2=2.035 $Y2=0.955
r37 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.905 $Y=0.955
+ $X2=1.215 $Y2=0.955
r38 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.05 $Y=0.87
+ $X2=1.215 $Y2=0.955
r39 7 9 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.05 $Y=0.87 $X2=1.05
+ $Y2=0.435
r40 2 18 182 $w=1.7e-07 $l=7.41704e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.28 $X2=2 $Y2=0.955
r41 2 15 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.28 $X2=2 $Y2=0.435
r42 1 9 91 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.235 $X2=1.05 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_2%VGND 1 2 3 12 16 18 21 23 24 26 27 29 41 47
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r52 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r53 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r54 41 46 5.00713 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.537
+ $Y2=0
r55 41 43 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.12
+ $Y2=0
r56 40 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r57 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r58 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 33 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r60 32 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r61 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r62 29 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r63 29 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r64 26 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.16
+ $Y2=0
r65 26 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.45
+ $Y2=0
r66 25 43 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=3.12
+ $Y2=0
r67 25 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.45
+ $Y2=0
r68 23 36 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.2
+ $Y2=0
r69 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.57
+ $Y2=0
r70 22 39 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=2.16
+ $Y2=0
r71 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.57
+ $Y2=0
r72 18 46 3.23308 $w=3.85e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.427 $Y=0.085
+ $X2=3.537 $Y2=0
r73 18 21 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=3.427 $Y=0.085
+ $X2=3.427 $Y2=0.425
r74 14 27 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0
r75 14 16 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0.425
r76 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0
r77 10 12 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0.575
r78 3 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.19
+ $Y=0.28 $X2=3.33 $Y2=0.425
r79 2 16 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.28 $X2=2.45 $Y2=0.425
r80 1 12 182 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.28 $X2=1.57 $Y2=0.575
.ends

