* File: sky130_fd_sc_lp__a31oi_1.spice
* Created: Fri Aug 28 09:59:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a31oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a31oi_1  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1003 A_151_47# N_A3_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.2268 PD=1.05 PS=2.22 NRD=7.14 NRS=0.708 M=1 R=5.6 SA=75000.2 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1006 A_223_47# N_A2_M1006_g A_151_47# VNB NSHORT L=0.15 W=0.84 AD=0.168
+ AS=0.0882 PD=1.24 PS=1.05 NRD=20.712 NRS=7.14 M=1 R=5.6 SA=75000.6 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1007 N_Y_M1007_d N_A1_M1007_g A_223_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.168 PD=1.23 PS=1.24 NRD=5.712 NRS=20.712 M=1 R=5.6 SA=75001.1 SB=75000.7
+ A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_151_367#_M1000_d N_A3_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_151_367#_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2772 AS=0.1764 PD=1.7 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1001 N_A_151_367#_M1001_d N_A1_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2772 PD=1.54 PS=1.7 NRD=0 NRS=12.4898 M=1 R=8.4
+ SA=75001.2 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_151_367#_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4347 AS=0.1764 PD=3.21 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75000.3 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__a31oi_1.pxi.spice"
*
.ends
*
*
