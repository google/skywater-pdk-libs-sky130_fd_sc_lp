* File: sky130_fd_sc_lp__nand2_0.pex.spice
* Created: Wed Sep  2 10:02:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2_0%B 2 5 9 11 12 13 14 15 21
r33 21 23 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.005
+ $X2=0.402 $Y2=0.84
r34 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.35
+ $Y=1.005 $X2=0.35 $Y2=1.005
r35 14 15 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.035
r36 13 14 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r37 13 22 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.005
r38 12 22 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=0.925 $X2=0.26
+ $Y2=1.005
r39 9 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.545 $Y=0.445
+ $X2=0.545 $Y2=0.84
r40 5 11 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=0.505 $Y=2.63
+ $X2=0.505 $Y2=1.51
r41 2 11 47.7177 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=0.402 $Y=1.293
+ $X2=0.402 $Y2=1.51
r42 1 21 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=0.402 $Y=1.057
+ $X2=0.402 $Y2=1.005
r43 1 2 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=0.402 $Y=1.057
+ $X2=0.402 $Y2=1.293
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_0%A 3 6 9 11 12 13 14 15 21
r27 21 23 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.047 $Y=1.005
+ $X2=1.047 $Y2=0.84
r28 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.07
+ $Y=1.005 $X2=1.07 $Y2=1.005
r29 14 15 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=2.035
r30 13 14 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.17 $Y=1.295
+ $X2=1.17 $Y2=1.665
r31 13 22 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.17 $Y=1.295
+ $X2=1.17 $Y2=1.005
r32 12 22 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=1.17 $Y=0.925 $X2=1.17
+ $Y2=1.005
r33 9 11 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=0.935 $Y=2.63
+ $X2=0.935 $Y2=1.51
r34 6 11 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=1.047 $Y=1.323
+ $X2=1.047 $Y2=1.51
r35 5 21 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=1.047 $Y=1.027
+ $X2=1.047 $Y2=1.005
r36 5 6 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=1.047 $Y=1.027
+ $X2=1.047 $Y2=1.323
r37 3 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.935 $Y=0.445
+ $X2=0.935 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_0%VPWR 1 2 7 9 11 13 15 17 27
r21 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r22 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 18 23 4.5263 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r24 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 17 26 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.212 $Y2=3.33
r26 17 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r28 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 11 26 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.212 $Y2=3.33
r31 11 13 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=2.455
r32 7 23 3.0729 $w=3.1e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.217 $Y2=3.33
r33 7 9 29.3687 $w=3.08e-07 $l=7.9e-07 $layer=LI1_cond $X=0.28 $Y=3.245 $X2=0.28
+ $Y2=2.455
r34 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.31 $X2=1.15 $Y2=2.455
r35 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.31 $X2=0.29 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_0%Y 1 2 9 11 12 13 14 15 16 17 26
r25 16 17 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=2.405
+ $X2=0.71 $Y2=2.775
r26 15 16 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=2.035
+ $X2=0.71 $Y2=2.405
r27 14 15 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=1.665
+ $X2=0.71 $Y2=2.035
r28 13 14 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=1.295
+ $X2=0.71 $Y2=1.665
r29 12 13 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=0.925
+ $X2=0.71 $Y2=1.295
r30 11 26 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=0.445
+ $X2=0.71 $Y2=0.61
r31 11 12 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=0.71 $Y=0.625 $X2=0.71
+ $Y2=0.925
r32 11 26 0.792208 $w=2.08e-07 $l=1.5e-08 $layer=LI1_cond $X=0.71 $Y=0.625
+ $X2=0.71 $Y2=0.61
r33 7 11 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=0.815 $Y=0.445
+ $X2=0.71 $Y2=0.445
r34 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0.445
+ $X2=1.15 $Y2=0.445
r35 2 16 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.31 $X2=0.72 $Y2=2.465
r36 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.235 $X2=1.15 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_0%VGND 1 4 6 8 12 13
r20 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r21 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r22 10 16 4.11415 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r23 10 12 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=1.2
+ $Y2=0
r24 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r25 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r26 4 16 3.17054 $w=2.7e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.217 $Y2=0
r27 4 6 15.3659 $w=2.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.3 $Y=0.085 $X2=0.3
+ $Y2=0.445
r28 1 6 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.235 $X2=0.33 $Y2=0.445
.ends

