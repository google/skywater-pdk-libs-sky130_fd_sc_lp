* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4bb_lp A B C_N D_N VGND VNB VPB VPWR X
X0 a_274_47# C_N a_318_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1284_47# D_N a_654_355# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_823_125# a_654_355# a_86_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR C_N a_318_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_505_400# B a_1076_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VGND A a_476_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_116_47# a_86_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_505_400# a_318_409# a_612_400# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_1076_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VPWR D_N a_654_355# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 X a_86_21# a_116_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND C_N a_274_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_654_355# a_823_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND D_N a_1284_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_476_125# A a_86_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_86_21# B a_981_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_665_125# a_318_409# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 X a_86_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X18 a_86_21# a_318_409# a_665_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_612_400# a_654_355# a_86_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 a_981_125# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
