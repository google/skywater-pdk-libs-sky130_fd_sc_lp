* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
X0 Q a_796_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_383_479# a_251_475# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_574_47# a_383_479# a_646_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_646_47# a_251_475# a_754_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_796_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_646_47# a_383_479# a_785_479# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_754_47# a_796_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR GATE a_251_475# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_40_54# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_796_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_383_479# a_251_475# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 Q a_796_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND a_40_54# a_574_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_40_54# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_796_21# a_646_47# a_1043_73# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_1043_73# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VGND GATE a_251_475# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_796_21# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_785_479# a_796_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VPWR a_40_54# a_611_479# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_611_479# a_251_475# a_646_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VPWR a_646_47# a_796_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
