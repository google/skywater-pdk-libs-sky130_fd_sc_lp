* File: sky130_fd_sc_lp__sdfrtp_1.pex.spice
* Created: Fri Aug 28 11:28:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%A_35_74# 1 2 7 9 12 16 19 22 23 25 27 32 34
+ 35
c73 34 0 8.22072e-20 $X=2.51 $Y=1.98
c74 23 0 1.42315e-19 $X=1.345 $Y=0.945
r75 35 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.98
+ $X2=2.51 $Y2=2.145
r76 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.98 $X2=2.51 $Y2=1.98
r77 31 32 11.9313 $w=9.88e-07 $l=9.5e-08 $layer=LI1_cond $X=1.055 $Y=2.47
+ $X2=1.15 $Y2=2.47
r78 28 31 10.1667 $w=9.88e-07 $l=8.25e-07 $layer=LI1_cond $X=0.23 $Y=2.47
+ $X2=1.055 $Y2=2.47
r79 25 34 2.99516 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=2.425 $Y=2.06
+ $X2=2.55 $Y2=1.98
r80 25 32 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=2.425 $Y=2.06
+ $X2=1.15 $Y2=2.06
r81 23 39 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=1.345 $Y=0.945
+ $X2=1.465 $Y2=0.945
r82 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.345
+ $Y=0.945 $X2=1.345 $Y2=0.945
r83 20 27 3.57226 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.43 $Y=0.945
+ $X2=0.26 $Y2=0.945
r84 20 22 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=0.43 $Y=0.945
+ $X2=1.345 $Y2=0.945
r85 19 28 8.32829 $w=2.8e-07 $l=4.95e-07 $layer=LI1_cond $X=0.23 $Y=1.975
+ $X2=0.23 $Y2=2.47
r86 18 27 3.05675 $w=3.1e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.23 $Y=1.03
+ $X2=0.26 $Y2=0.945
r87 18 19 38.895 $w=2.78e-07 $l=9.45e-07 $layer=LI1_cond $X=0.23 $Y=1.03
+ $X2=0.23 $Y2=1.975
r88 14 27 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.86 $X2=0.26
+ $Y2=0.945
r89 14 16 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=0.26 $Y=0.86
+ $X2=0.26 $Y2=0.58
r90 12 42 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.49 $Y=2.635
+ $X2=2.49 $Y2=2.145
r91 7 39 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=0.78
+ $X2=1.465 $Y2=0.945
r92 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.465 $Y=0.78
+ $X2=1.465 $Y2=0.46
r93 2 31 150 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=4 $X=0.59
+ $Y=2.315 $X2=1.055 $Y2=2.46
r94 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.37 $X2=0.3 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%SCE 3 6 7 8 11 13 17 21 23 24 25 26 27 28
+ 35 39
c71 39 0 1.6277e-19 $X=2.395 $Y=1.295
c72 13 0 1.24551e-19 $X=1.625 $Y=2.105
r73 39 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.295
+ $X2=2.395 $Y2=1.13
r74 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.395
+ $Y=1.295 $X2=2.395 $Y2=1.295
r75 35 37 47.6426 $w=4.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.677 $Y=1.295
+ $X2=0.677 $Y2=1.13
r76 28 40 13.9347 $w=1.93e-07 $l=2.45e-07 $layer=LI1_cond $X=2.64 $Y=1.297
+ $X2=2.395 $Y2=1.297
r77 27 40 13.366 $w=1.93e-07 $l=2.35e-07 $layer=LI1_cond $X=2.16 $Y=1.297
+ $X2=2.395 $Y2=1.297
r78 26 27 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.297
+ $X2=2.16 $Y2=1.297
r79 25 26 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.297
+ $X2=1.68 $Y2=1.297
r80 24 25 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.297
+ $X2=1.2 $Y2=1.297
r81 24 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.295 $X2=0.75 $Y2=1.295
r82 21 41 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.485 $Y=0.615
+ $X2=2.485 $Y2=1.13
r83 15 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.7 $Y=2.18 $X2=1.7
+ $Y2=2.635
r84 14 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.345 $Y=2.105
+ $X2=1.27 $Y2=2.105
r85 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.625 $Y=2.105
+ $X2=1.7 $Y2=2.18
r86 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.625 $Y=2.105
+ $X2=1.345 $Y2=2.105
r87 9 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.27 $Y=2.18 $X2=1.27
+ $Y2=2.105
r88 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.27 $Y=2.18
+ $X2=1.27 $Y2=2.635
r89 7 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.195 $Y=2.105
+ $X2=1.27 $Y2=2.105
r90 7 8 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.195 $Y=2.105
+ $X2=0.915 $Y2=2.105
r91 6 8 37.7275 $w=1.5e-07 $l=2.72936e-07 $layer=POLY_cond $X=0.677 $Y=2.03
+ $X2=0.915 $Y2=2.105
r92 5 35 8.43012 $w=4.75e-07 $l=7.2e-08 $layer=POLY_cond $X=0.677 $Y=1.367
+ $X2=0.677 $Y2=1.295
r93 5 6 77.6274 $w=4.75e-07 $l=6.63e-07 $layer=POLY_cond $X=0.677 $Y=1.367
+ $X2=0.677 $Y2=2.03
r94 3 37 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.515 $Y=0.58
+ $X2=0.515 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%D 3 7 9 10 11 12 18
c35 12 0 1.24551e-19 $X=2.16 $Y=1.665
c36 7 0 8.22072e-20 $X=2.06 $Y=2.635
r37 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.655 $X2=1.825 $Y2=1.655
r38 12 19 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=2.16 $Y=1.685
+ $X2=1.825 $Y2=1.685
r39 11 19 6.96268 $w=2.38e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=1.685
+ $X2=1.825 $Y2=1.685
r40 10 11 23.0489 $w=2.38e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.685
+ $X2=1.68 $Y2=1.685
r41 9 10 23.0489 $w=2.38e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.685 $X2=1.2
+ $Y2=1.685
r42 5 18 38.3966 $w=2.95e-07 $l=3.1229e-07 $layer=POLY_cond $X=2.06 $Y=1.82
+ $X2=1.825 $Y2=1.64
r43 5 7 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.06 $Y=1.82 $X2=2.06
+ $Y2=2.635
r44 1 18 18.5736 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.825 $Y=1.46
+ $X2=1.825 $Y2=1.64
r45 1 3 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=1.825 $Y=1.46 $X2=1.825
+ $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%SCD 3 7 11 13 14 15 16 21
c46 7 0 9.78661e-20 $X=2.96 $Y=2.635
c47 3 0 3.56444e-20 $X=2.845 $Y=0.615
r48 15 16 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.137 $Y=1.665
+ $X2=3.137 $Y2=2.035
r49 14 15 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.137 $Y=1.295
+ $X2=3.137 $Y2=1.665
r50 14 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.05
+ $Y=1.34 $X2=3.05 $Y2=1.34
r51 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.05 $Y=1.68
+ $X2=3.05 $Y2=1.34
r52 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.68
+ $X2=3.05 $Y2=1.845
r53 11 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.05 $Y=1.325
+ $X2=3.05 $Y2=1.34
r54 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.992 $Y=1.175
+ $X2=2.992 $Y2=1.325
r55 7 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.96 $Y=2.635
+ $X2=2.96 $Y2=1.845
r56 3 10 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.845 $Y=0.615
+ $X2=2.845 $Y2=1.175
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%A_757_317# 1 2 9 13 14 16 19 22 23 27 28 32
+ 35 36 37 38 39 40 43 52 53 56 61 62 63
c206 40 0 1.85618e-19 $X=7.585 $Y=1.295
c207 28 0 3.68148e-20 $X=7.955 $Y=2.22
c208 27 0 2.82467e-20 $X=7.955 $Y=2.22
c209 23 0 1.53911e-19 $X=7.77 $Y=1.26
r210 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.44
+ $Y=1.26 $X2=7.44 $Y2=1.26
r211 61 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.9 $Y=1.29
+ $X2=4.9 $Y2=1.125
r212 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=1.29 $X2=4.9 $Y2=1.29
r213 56 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.75
+ $X2=3.95 $Y2=1.915
r214 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.75 $X2=3.95 $Y2=1.75
r215 53 84 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=10.38 $Y=1.295
+ $X2=10.38 $Y2=2.035
r216 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=1.295
+ $X2=10.32 $Y2=1.295
r217 49 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.295
+ $X2=7.44 $Y2=1.295
r218 46 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.295
r219 43 57 14.5656 $w=3.58e-07 $l=4.55e-07 $layer=LI1_cond $X=4.035 $Y=1.295
+ $X2=4.035 $Y2=1.75
r220 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.295
r221 40 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.295
+ $X2=7.44 $Y2=1.295
r222 39 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=10.32 $Y2=1.295
r223 39 40 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=7.585 $Y2=1.295
r224 38 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.295
+ $X2=5.04 $Y2=1.295
r225 37 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.295 $Y=1.295
+ $X2=7.44 $Y2=1.295
r226 37 38 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=7.295 $Y=1.295
+ $X2=5.185 $Y2=1.295
r227 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.295
+ $X2=4.08 $Y2=1.295
r228 35 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=5.04 $Y2=1.295
r229 35 36 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=4.225 $Y2=1.295
r230 34 53 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=10.38 $Y=1.165
+ $X2=10.38 $Y2=1.295
r231 32 34 2.82206 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=10.395 $Y=1.08
+ $X2=10.395 $Y2=1.165
r232 28 69 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=7.955 $Y=2.22
+ $X2=7.815 $Y2=2.22
r233 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.955
+ $Y=2.22 $X2=7.955 $Y2=2.22
r234 24 27 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=7.855 $Y=2.18
+ $X2=7.955 $Y2=2.18
r235 23 68 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=7.77 $Y=1.26
+ $X2=7.44 $Y2=1.26
r236 22 24 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.855 $Y=2.055
+ $X2=7.855 $Y2=2.18
r237 21 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.855 $Y=1.425
+ $X2=7.77 $Y2=1.26
r238 21 22 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=7.855 $Y=1.425
+ $X2=7.855 $Y2=2.055
r239 17 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.815 $Y=2.385
+ $X2=7.815 $Y2=2.22
r240 17 19 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=7.815 $Y=2.385
+ $X2=7.815 $Y2=2.875
r241 14 67 53.3511 $w=2.62e-07 $l=3.63249e-07 $layer=POLY_cond $X=7.15 $Y=1.095
+ $X2=7.44 $Y2=1.26
r242 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.15 $Y=1.095
+ $X2=7.15 $Y2=0.665
r243 13 63 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.88 $Y=0.805
+ $X2=4.88 $Y2=1.125
r244 9 59 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.97 $Y=2.525
+ $X2=3.97 $Y2=1.915
r245 2 84 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=10.325
+ $Y=1.835 $X2=10.45 $Y2=2.035
r246 1 32 182 $w=1.7e-07 $l=7.84156e-07 $layer=licon1_NDIFF $count=1 $X=10.265
+ $Y=0.365 $X2=10.41 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%A_937_333# 1 2 9 11 15 18 20 21 26 28 29 31
+ 33 42 44 48
c98 44 0 2.9296e-19 $X=6.74 $Y=1.685
c99 33 0 1.16283e-19 $X=4.87 $Y=1.685
c100 31 0 5.31087e-20 $X=6.98 $Y=2.055
c101 28 0 1.85378e-20 $X=6.745 $Y=1.96
r102 39 42 10.2148 $w=2.18e-07 $l=1.95e-07 $layer=LI1_cond $X=6.74 $Y=0.465
+ $X2=6.935 $Y2=0.465
r103 37 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.83
+ $X2=5.015 $Y2=1.83
r104 37 45 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.85 $Y=1.83 $X2=4.76
+ $Y2=1.83
r105 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.83 $X2=4.85 $Y2=1.83
r106 33 36 5.76222 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=4.87 $Y=1.685
+ $X2=4.87 $Y2=1.83
r107 29 31 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=6.835 $Y=2.055
+ $X2=6.98 $Y2=2.055
r108 28 29 6.82297 $w=1.9e-07 $l=1.32571e-07 $layer=LI1_cond $X=6.745 $Y=1.96
+ $X2=6.835 $Y2=2.055
r109 27 44 4.81226 $w=1.85e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.745 $Y=1.77
+ $X2=6.74 $Y2=1.685
r110 27 28 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=6.745 $Y=1.77
+ $X2=6.745 $Y2=1.96
r111 24 44 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=6.74 $Y=1.6
+ $X2=6.74 $Y2=1.685
r112 24 26 43.1962 $w=1.88e-07 $l=7.4e-07 $layer=LI1_cond $X=6.74 $Y=1.6
+ $X2=6.74 $Y2=0.86
r113 23 39 1.59589 $w=1.9e-07 $l=1.1e-07 $layer=LI1_cond $X=6.74 $Y=0.575
+ $X2=6.74 $Y2=0.465
r114 23 26 16.6364 $w=1.88e-07 $l=2.85e-07 $layer=LI1_cond $X=6.74 $Y=0.575
+ $X2=6.74 $Y2=0.86
r115 22 33 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.015 $Y=1.685
+ $X2=4.87 $Y2=1.685
r116 21 44 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.645 $Y=1.685
+ $X2=6.74 $Y2=1.685
r117 21 22 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=6.645 $Y=1.685
+ $X2=5.015 $Y2=1.685
r118 19 20 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.365 $Y=1.275
+ $X2=5.365 $Y2=1.425
r119 18 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.38 $Y=1.695
+ $X2=5.38 $Y2=1.425
r120 15 19 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.35 $Y=0.805 $X2=5.35
+ $Y2=1.275
r121 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.305 $Y=1.77
+ $X2=5.38 $Y2=1.695
r122 11 48 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.305 $Y=1.77
+ $X2=5.015 $Y2=1.77
r123 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.76 $Y=1.995
+ $X2=4.76 $Y2=1.83
r124 7 9 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.76 $Y=1.995
+ $X2=4.76 $Y2=2.525
r125 2 31 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.895 $X2=6.98 $Y2=2.055
r126 1 42 182 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=1 $X=6.6
+ $Y=0.345 $X2=6.935 $Y2=0.47
r127 1 26 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=6.6
+ $Y=0.345 $X2=6.74 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%RESET_B 3 7 8 9 12 13 15 16 18 20 21 22 28
+ 31 35 37 38 39 41 42 45 46 47 49 50 51 53 56 57 62 64 70
c211 70 0 6.31513e-20 $X=9.24 $Y=2.34
c212 38 0 1.11215e-19 $X=3.472 $Y=2.205
c213 31 0 2.92081e-20 $X=9.015 $Y=0.805
c214 16 0 1.14005e-19 $X=5.785 $Y=0.18
c215 15 0 5.71712e-20 $X=3.845 $Y=1.195
c216 12 0 9.02003e-20 $X=3.77 $Y=1.27
r217 62 64 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=5.942 $Y=2.04
+ $X2=5.942 $Y2=1.875
r218 56 57 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=5.965 $Y=2.035
+ $X2=5.965 $Y2=2.32
r219 56 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.965
+ $Y=2.04 $X2=5.965 $Y2=2.04
r220 54 70 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=9.105 $Y=2.34
+ $X2=9.24 $Y2=2.34
r221 54 67 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.105 $Y=2.34
+ $X2=9.015 $Y2=2.34
r222 53 55 8.41379 $w=3.19e-07 $l=2.2e-07 $layer=LI1_cond $X=9.105 $Y=2.34
+ $X2=9.105 $Y2=2.56
r223 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.105
+ $Y=2.34 $X2=9.105 $Y2=2.34
r224 50 55 4.42298 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.94 $Y=2.56
+ $X2=9.105 $Y2=2.56
r225 50 51 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.94 $Y=2.56
+ $X2=8.285 $Y2=2.56
r226 48 51 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.16 $Y=2.645
+ $X2=8.285 $Y2=2.56
r227 48 49 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=8.16 $Y=2.645
+ $X2=8.16 $Y2=2.905
r228 46 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.035 $Y=2.99
+ $X2=8.16 $Y2=2.905
r229 46 47 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=8.035 $Y=2.99
+ $X2=6.95 $Y2=2.99
r230 45 47 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.86 $Y=2.905
+ $X2=6.95 $Y2=2.99
r231 44 45 25.5707 $w=1.78e-07 $l=4.15e-07 $layer=LI1_cond $X=6.86 $Y=2.49
+ $X2=6.86 $Y2=2.905
r232 43 57 4.90495 $w=1.7e-07 $l=1.77989e-07 $layer=LI1_cond $X=6.13 $Y=2.405
+ $X2=5.965 $Y2=2.432
r233 42 44 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.77 $Y=2.405
+ $X2=6.86 $Y2=2.49
r234 42 43 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.77 $Y=2.405
+ $X2=6.13 $Y2=2.405
r235 41 64 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=5.83 $Y=1.245
+ $X2=5.83 $Y2=1.875
r236 40 41 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.845 $Y=1.095
+ $X2=5.845 $Y2=1.245
r237 37 38 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=3.472 $Y=2.055
+ $X2=3.472 $Y2=2.205
r238 33 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.24 $Y=2.505
+ $X2=9.24 $Y2=2.34
r239 33 35 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.24 $Y=2.505
+ $X2=9.24 $Y2=2.875
r240 29 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.015 $Y=2.175
+ $X2=9.015 $Y2=2.34
r241 29 31 702.489 $w=1.5e-07 $l=1.37e-06 $layer=POLY_cond $X=9.015 $Y=2.175
+ $X2=9.015 $Y2=0.805
r242 28 40 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.86 $Y=0.775
+ $X2=5.86 $Y2=1.095
r243 25 28 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.86 $Y=0.255
+ $X2=5.86 $Y2=0.775
r244 21 62 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=5.942 $Y=2.13
+ $X2=5.942 $Y2=2.04
r245 21 22 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=5.755 $Y=2.13
+ $X2=5.375 $Y2=2.13
r246 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.3 $Y=2.205
+ $X2=5.375 $Y2=2.13
r247 18 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.3 $Y=2.205
+ $X2=5.3 $Y2=2.525
r248 17 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.92 $Y=0.18
+ $X2=3.845 $Y2=0.18
r249 16 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.785 $Y=0.18
+ $X2=5.86 $Y2=0.255
r250 16 17 956.309 $w=1.5e-07 $l=1.865e-06 $layer=POLY_cond $X=5.785 $Y=0.18
+ $X2=3.92 $Y2=0.18
r251 14 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.845 $Y=0.255
+ $X2=3.845 $Y2=0.18
r252 14 15 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.845 $Y=0.255
+ $X2=3.845 $Y2=1.195
r253 12 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.77 $Y=1.27
+ $X2=3.845 $Y2=1.195
r254 12 13 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.77 $Y=1.27
+ $X2=3.575 $Y2=1.27
r255 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.5 $Y=1.345
+ $X2=3.575 $Y2=1.27
r256 10 37 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.5 $Y=1.345
+ $X2=3.5 $Y2=2.055
r257 8 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=0.18
+ $X2=3.845 $Y2=0.18
r258 8 9 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=3.77 $Y=0.18
+ $X2=3.395 $Y2=0.18
r259 7 38 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.445 $Y=2.635
+ $X2=3.445 $Y2=2.205
r260 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.32 $Y=0.255
+ $X2=3.395 $Y2=0.18
r261 1 3 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.32 $Y=0.255
+ $X2=3.32 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%A_809_463# 1 2 3 12 16 19 20 21 24 28 32 35
+ 39
c115 35 0 1.11215e-19 $X=4.287 $Y=2.25
c116 21 0 5.71712e-20 $X=4.555 $Y=0.89
c117 20 0 1.16283e-19 $X=6.145 $Y=0.89
c118 16 0 5.31087e-20 $X=6.765 $Y=2.315
r119 35 37 7.71264 $w=4.35e-07 $l=2.75e-07 $layer=LI1_cond $X=4.287 $Y=2.25
+ $X2=4.287 $Y2=2.525
r120 33 39 29.1096 $w=3.56e-07 $l=2.15e-07 $layer=POLY_cond $X=6.31 $Y=1.402
+ $X2=6.525 $Y2=1.402
r121 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.31
+ $Y=1.335 $X2=6.31 $Y2=1.335
r122 30 32 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.31 $Y=0.995
+ $X2=6.31 $Y2=1.335
r123 26 28 8.2628 $w=2.63e-07 $l=1.9e-07 $layer=LI1_cond $X=5.497 $Y=2.335
+ $X2=5.497 $Y2=2.525
r124 25 35 6.29128 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=4.555 $Y=2.25
+ $X2=4.287 $Y2=2.25
r125 24 26 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=5.365 $Y=2.25
+ $X2=5.497 $Y2=2.335
r126 24 25 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.365 $Y=2.25
+ $X2=4.555 $Y2=2.25
r127 21 23 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=4.555 $Y=0.89
+ $X2=4.665 $Y2=0.89
r128 20 30 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=6.145 $Y=0.89
+ $X2=6.31 $Y2=0.995
r129 20 23 78.1645 $w=2.08e-07 $l=1.48e-06 $layer=LI1_cond $X=6.145 $Y=0.89
+ $X2=4.665 $Y2=0.89
r130 19 35 9.32629 $w=4.35e-07 $l=2.52357e-07 $layer=LI1_cond $X=4.47 $Y=2.085
+ $X2=4.287 $Y2=2.25
r131 18 21 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.47 $Y=0.995
+ $X2=4.555 $Y2=0.89
r132 18 19 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=2.085
r133 14 39 32.4944 $w=3.56e-07 $l=3.36927e-07 $layer=POLY_cond $X=6.765 $Y=1.635
+ $X2=6.525 $Y2=1.402
r134 14 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.765 $Y=1.635
+ $X2=6.765 $Y2=2.315
r135 10 39 23.0368 $w=1.5e-07 $l=2.32e-07 $layer=POLY_cond $X=6.525 $Y=1.17
+ $X2=6.525 $Y2=1.402
r136 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.525 $Y=1.17
+ $X2=6.525 $Y2=0.665
r137 3 28 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.375
+ $Y=2.315 $X2=5.515 $Y2=2.525
r138 2 37 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=2.315 $X2=4.185 $Y2=2.525
r139 1 23 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.595 $X2=4.665 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%A_865_255# 1 2 10 13 15 16 20 21 22 25 29
+ 33 36 38 39 42 43 44 46 51 53 55 56 57 58 64
c201 56 0 6.7118e-20 $X=10.8 $Y=1.51
c202 55 0 1.23014e-19 $X=10.8 $Y=1.51
c203 53 0 2.24062e-19 $X=8.37 $Y=1.65
c204 38 0 1.80416e-19 $X=7.815 $Y=1.635
c205 22 0 1.54882e-19 $X=7.27 $Y=1.71
c206 21 0 2.82467e-20 $X=7.815 $Y=1.71
r207 68 70 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=10.625 $Y=1.51
+ $X2=10.665 $Y2=1.51
r208 61 64 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=11.29 $Y=1.085
+ $X2=11.465 $Y2=1.085
r209 58 60 8.95413 $w=4.36e-07 $l=3.2e-07 $layer=LI1_cond $X=11.21 $Y=2.455
+ $X2=11.21 $Y2=2.775
r210 56 70 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=10.8 $Y=1.51
+ $X2=10.665 $Y2=1.51
r211 55 57 10.1645 $w=6.63e-07 $l=1.65e-07 $layer=LI1_cond $X=11.047 $Y=1.51
+ $X2=11.047 $Y2=1.345
r212 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.8
+ $Y=1.51 $X2=10.8 $Y2=1.51
r213 50 53 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=1.65
+ $X2=8.37 $Y2=1.65
r214 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.205
+ $Y=1.65 $X2=8.205 $Y2=1.65
r215 47 61 1.35108 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=11.29 $Y=1.185
+ $X2=11.29 $Y2=1.085
r216 47 57 9.85859 $w=1.78e-07 $l=1.6e-07 $layer=LI1_cond $X=11.29 $Y=1.185
+ $X2=11.29 $Y2=1.345
r217 46 58 3.0058 $w=6.65e-07 $l=2.01057e-07 $layer=LI1_cond $X=11.047 $Y=2.37
+ $X2=11.21 $Y2=2.455
r218 45 55 3.00369 $w=6.63e-07 $l=1.67e-07 $layer=LI1_cond $X=11.047 $Y=1.677
+ $X2=11.047 $Y2=1.51
r219 45 46 12.4644 $w=6.63e-07 $l=6.93e-07 $layer=LI1_cond $X=11.047 $Y=1.677
+ $X2=11.047 $Y2=2.37
r220 43 58 6.30541 $w=1.7e-07 $l=4.95e-07 $layer=LI1_cond $X=10.715 $Y=2.455
+ $X2=11.21 $Y2=2.455
r221 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.715 $Y=2.455
+ $X2=10.045 $Y2=2.455
r222 42 44 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=9.922 $Y=2.37
+ $X2=10.045 $Y2=2.455
r223 41 42 30.3398 $w=2.43e-07 $l=6.45e-07 $layer=LI1_cond $X=9.922 $Y=1.725
+ $X2=9.922 $Y2=2.37
r224 39 41 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=9.8 $Y=1.64
+ $X2=9.922 $Y2=1.725
r225 39 53 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=9.8 $Y=1.64
+ $X2=8.37 $Y2=1.64
r226 37 51 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.995 $Y=1.65
+ $X2=8.205 $Y2=1.65
r227 37 38 13.5877 $w=2.4e-07 $l=1.8735e-07 $layer=POLY_cond $X=7.995 $Y=1.65
+ $X2=7.815 $Y2=1.635
r228 35 36 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.425 $Y=1.275
+ $X2=4.425 $Y2=1.425
r229 31 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.665 $Y=1.675
+ $X2=10.665 $Y2=1.51
r230 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.665 $Y=1.675
+ $X2=10.665 $Y2=2.465
r231 27 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.625 $Y=1.345
+ $X2=10.625 $Y2=1.51
r232 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.625 $Y=1.345
+ $X2=10.625 $Y2=0.785
r233 23 38 12.1617 $w=1.5e-07 $l=1.95576e-07 $layer=POLY_cond $X=7.92 $Y=1.485
+ $X2=7.815 $Y2=1.635
r234 23 25 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.92 $Y=1.485
+ $X2=7.92 $Y2=0.775
r235 21 38 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=7.815 $Y=1.71
+ $X2=7.815 $Y2=1.635
r236 21 22 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.815 $Y=1.71
+ $X2=7.27 $Y2=1.71
r237 18 20 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.195 $Y=3.075
+ $X2=7.195 $Y2=2.315
r238 17 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.195 $Y=1.785
+ $X2=7.27 $Y2=1.71
r239 17 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.195 $Y=1.785
+ $X2=7.195 $Y2=2.315
r240 15 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.12 $Y=3.15
+ $X2=7.195 $Y2=3.075
r241 15 16 1356.27 $w=1.5e-07 $l=2.645e-06 $layer=POLY_cond $X=7.12 $Y=3.15
+ $X2=4.475 $Y2=3.15
r242 13 35 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.45 $Y=0.805 $X2=4.45
+ $Y2=1.275
r243 10 36 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=4.4 $Y=2.525
+ $X2=4.4 $Y2=1.425
r244 8 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.4 $Y=3.075
+ $X2=4.475 $Y2=3.15
r245 8 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.4 $Y=3.075 $X2=4.4
+ $Y2=2.525
r246 2 60 600 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=11.325
+ $Y=1.835 $X2=11.465 $Y2=2.775
r247 1 64 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=11.325
+ $Y=0.365 $X2=11.465 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%A_1445_69# 1 2 7 9 12 16 20 24 26 28 31 33
+ 35 37 38 42 44 46 47 48 50 62 63 64 69 70
c204 69 0 3.17486e-19 $X=12.29 $Y=1.08
c205 44 0 1.85618e-19 $X=8.32 $Y=1.22
c206 35 0 9.19974e-20 $X=7.41 $Y=2.04
c207 33 0 8.84191e-20 $X=7.445 $Y=1.79
r208 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.29
+ $Y=1.08 $X2=12.29 $Y2=1.08
r209 66 69 24.3384 $w=1.78e-07 $l=3.95e-07 $layer=LI1_cond $X=11.895 $Y=1.075
+ $X2=12.29 $Y2=1.075
r210 62 75 4.53008 $w=2.66e-07 $l=2.5e-08 $layer=POLY_cond $X=9.645 $Y=1.29
+ $X2=9.67 $Y2=1.29
r211 61 64 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=9.645 $Y=1.26
+ $X2=9.96 $Y2=1.26
r212 61 63 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=9.645 $Y=1.26
+ $X2=9.48 $Y2=1.26
r213 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.645
+ $Y=1.29 $X2=9.645 $Y2=1.29
r214 50 66 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=11.895 $Y=0.985
+ $X2=11.895 $Y2=1.075
r215 49 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.895 $Y=0.815
+ $X2=11.895 $Y2=0.985
r216 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.81 $Y=0.73
+ $X2=11.895 $Y2=0.815
r217 47 48 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=11.81 $Y=0.73
+ $X2=10.045 $Y2=0.73
r218 46 64 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.96 $Y=1.135
+ $X2=9.96 $Y2=1.26
r219 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.96 $Y=0.815
+ $X2=10.045 $Y2=0.73
r220 45 46 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.96 $Y=0.815
+ $X2=9.96 $Y2=1.135
r221 44 63 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=8.32 $Y=1.22
+ $X2=9.48 $Y2=1.22
r222 42 44 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.215 $Y=1.135
+ $X2=8.32 $Y2=1.22
r223 41 42 11.619 $w=2.08e-07 $l=2.2e-07 $layer=LI1_cond $X=8.215 $Y=0.915
+ $X2=8.215 $Y2=1.135
r224 38 40 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.53 $Y=0.83
+ $X2=7.705 $Y2=0.83
r225 37 41 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.11 $Y=0.83
+ $X2=8.215 $Y2=0.915
r226 37 40 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.11 $Y=0.83
+ $X2=7.705 $Y2=0.83
r227 33 56 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.445 $Y=1.705
+ $X2=7.09 $Y2=1.705
r228 33 35 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=7.445 $Y=1.79
+ $X2=7.445 $Y2=2.04
r229 29 38 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.4 $Y=0.83
+ $X2=7.53 $Y2=0.83
r230 29 53 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.4 $Y=0.83
+ $X2=7.09 $Y2=0.83
r231 29 31 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=7.4 $Y=0.745
+ $X2=7.4 $Y2=0.49
r232 28 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=1.62
+ $X2=7.09 $Y2=1.705
r233 27 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=0.915
+ $X2=7.09 $Y2=0.83
r234 27 28 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.09 $Y=0.915
+ $X2=7.09 $Y2=1.62
r235 25 70 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=12.29 $Y=1.42
+ $X2=12.29 $Y2=1.08
r236 25 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.29 $Y=1.42
+ $X2=12.29 $Y2=1.585
r237 24 70 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=12.29 $Y=1.065
+ $X2=12.29 $Y2=1.08
r238 23 24 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=12.327 $Y=0.915
+ $X2=12.327 $Y2=1.065
r239 20 23 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=12.455 $Y=0.445
+ $X2=12.455 $Y2=0.915
r240 16 26 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=12.38 $Y=2.155
+ $X2=12.38 $Y2=1.585
r241 10 75 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.67 $Y=1.455
+ $X2=9.67 $Y2=1.29
r242 10 12 728.128 $w=1.5e-07 $l=1.42e-06 $layer=POLY_cond $X=9.67 $Y=1.455
+ $X2=9.67 $Y2=2.875
r243 7 62 48.9248 $w=2.66e-07 $l=3.4271e-07 $layer=POLY_cond $X=9.375 $Y=1.125
+ $X2=9.645 $Y2=1.29
r244 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.375 $Y=1.125
+ $X2=9.375 $Y2=0.805
r245 2 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.27
+ $Y=1.895 $X2=7.41 $Y2=2.04
r246 1 40 182 $w=1.7e-07 $l=6.84124e-07 $layer=licon1_NDIFF $count=1 $X=7.225
+ $Y=0.345 $X2=7.705 $Y2=0.83
r247 1 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.225
+ $Y=0.345 $X2=7.365 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%A_1641_21# 1 2 10 13 15 16 17 18 20 21 25
+ 29 31 34 39 40 45 47
c113 34 0 6.31513e-20 $X=8.565 $Y=1.99
c114 29 0 2.92081e-20 $X=9.705 $Y=0.365
c115 18 0 3.41158e-19 $X=8.355 $Y=1.17
r116 39 40 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.49 $Y=2.91
+ $X2=9.49 $Y2=2.745
r117 37 45 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.565 $Y=2.22
+ $X2=8.655 $Y2=2.22
r118 37 42 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=8.565 $Y=2.22
+ $X2=8.405 $Y2=2.22
r119 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.565
+ $Y=2.22 $X2=8.565 $Y2=2.22
r120 34 36 10.3926 $w=2.7e-07 $l=2.3e-07 $layer=LI1_cond $X=8.565 $Y=1.99
+ $X2=8.565 $Y2=2.22
r121 32 47 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=9.99 $Y=0.35
+ $X2=9.99 $Y2=0.18
r122 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.99
+ $Y=0.35 $X2=9.99 $Y2=0.35
r123 29 31 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=9.705 $Y=0.365
+ $X2=9.99 $Y2=0.365
r124 27 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.535 $Y=2.075
+ $X2=9.535 $Y2=2.745
r125 23 29 6.94494 $w=2.2e-07 $l=1.87083e-07 $layer=LI1_cond $X=9.565 $Y=0.475
+ $X2=9.705 $Y2=0.365
r126 23 25 13.3766 $w=2.78e-07 $l=3.25e-07 $layer=LI1_cond $X=9.565 $Y=0.475
+ $X2=9.565 $Y2=0.8
r127 22 34 3.44395 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.73 $Y=1.99
+ $X2=8.565 $Y2=1.99
r128 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.45 $Y=1.99
+ $X2=9.535 $Y2=2.075
r129 21 22 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=9.45 $Y=1.99
+ $X2=8.73 $Y2=1.99
r130 20 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.655 $Y=2.055
+ $X2=8.655 $Y2=2.22
r131 19 20 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=8.655 $Y=1.245
+ $X2=8.655 $Y2=2.055
r132 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.58 $Y=1.17
+ $X2=8.655 $Y2=1.245
r133 17 18 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=8.58 $Y=1.17
+ $X2=8.355 $Y2=1.17
r134 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.825 $Y=0.18
+ $X2=9.99 $Y2=0.18
r135 15 16 753.766 $w=1.5e-07 $l=1.47e-06 $layer=POLY_cond $X=9.825 $Y=0.18
+ $X2=8.355 $Y2=0.18
r136 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.405 $Y=2.385
+ $X2=8.405 $Y2=2.22
r137 11 13 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=8.405 $Y=2.385
+ $X2=8.405 $Y2=2.875
r138 8 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.28 $Y=1.095
+ $X2=8.355 $Y2=1.17
r139 8 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.28 $Y=1.095
+ $X2=8.28 $Y2=0.775
r140 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.28 $Y=0.255
+ $X2=8.355 $Y2=0.18
r141 7 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=8.28 $Y=0.255
+ $X2=8.28 $Y2=0.775
r142 2 39 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=9.315
+ $Y=2.665 $X2=9.455 $Y2=2.91
r143 1 25 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=9.45
+ $Y=0.595 $X2=9.59 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%CLK 3 7 9 11 12 13 14 18 22
c44 22 0 2.35026e-19 $X=11.715 $Y=1.51
r45 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.715
+ $Y=1.51 $X2=11.715 $Y2=1.51
r46 18 21 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.715 $Y=1.42
+ $X2=11.715 $Y2=1.51
r47 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.715 $Y=2.035
+ $X2=11.715 $Y2=2.405
r48 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.715 $Y=1.665
+ $X2=11.715 $Y2=2.035
r49 12 22 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=11.715 $Y=1.665
+ $X2=11.715 $Y2=1.51
r50 10 11 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.325 $Y=1.42
+ $X2=11.25 $Y2=1.42
r51 9 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.55 $Y=1.42
+ $X2=11.715 $Y2=1.42
r52 9 10 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=11.55 $Y=1.42
+ $X2=11.325 $Y2=1.42
r53 5 11 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.25 $Y=1.495
+ $X2=11.25 $Y2=1.42
r54 5 7 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=11.25 $Y=1.495
+ $X2=11.25 $Y2=2.465
r55 1 11 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.25 $Y=1.345
+ $X2=11.25 $Y2=1.42
r56 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.25 $Y=1.345
+ $X2=11.25 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%A_2408_367# 1 2 9 13 17 21 23 24 25 26 30
+ 31
c57 30 0 1.96847e-19 $X=12.83 $Y=1.47
c58 23 0 2.77631e-20 $X=12.665 $Y=1.76
c59 9 0 2.89723e-19 $X=12.965 $Y=0.655
r60 31 34 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=12.852 $Y=1.47
+ $X2=12.852 $Y2=1.635
r61 31 33 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=12.852 $Y=1.47
+ $X2=12.852 $Y2=1.305
r62 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.83
+ $Y=1.47 $X2=12.83 $Y2=1.47
r63 28 30 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=12.79 $Y=1.675
+ $X2=12.79 $Y2=1.47
r64 27 30 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=12.79 $Y=0.815
+ $X2=12.79 $Y2=1.47
r65 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.665 $Y=0.73
+ $X2=12.79 $Y2=0.815
r66 25 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.665 $Y=0.73
+ $X2=12.405 $Y2=0.73
r67 23 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.665 $Y=1.76
+ $X2=12.79 $Y2=1.675
r68 23 24 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=12.665 $Y=1.76
+ $X2=12.26 $Y2=1.76
r69 19 26 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=12.277 $Y=0.645
+ $X2=12.405 $Y2=0.73
r70 19 21 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=12.277 $Y=0.645
+ $X2=12.277 $Y2=0.44
r71 15 24 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=12.155 $Y=1.845
+ $X2=12.26 $Y2=1.76
r72 15 17 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=12.155 $Y=1.845
+ $X2=12.155 $Y2=1.98
r73 13 34 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=12.965 $Y=2.465
+ $X2=12.965 $Y2=1.635
r74 9 33 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=12.965 $Y=0.655
+ $X2=12.965 $Y2=1.305
r75 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.04
+ $Y=1.835 $X2=12.165 $Y2=1.98
r76 1 21 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=12.115
+ $Y=0.235 $X2=12.24 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 41 45 49
+ 53 58 59 60 69 73 81 94 99 109 110 113 116 119 124 127 129 132 135
c150 53 0 1.67908e-19 $X=12.595 $Y=2.1
r151 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r152 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r153 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r154 126 127 9.89636 $w=5.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=3.135
+ $X2=9.19 $Y2=3.135
r155 123 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r156 122 126 3.09699 $w=5.58e-07 $l=1.45e-07 $layer=LI1_cond $X=8.88 $Y=3.135
+ $X2=9.025 $Y2=3.135
r157 122 124 15.4496 $w=5.58e-07 $l=4.25e-07 $layer=LI1_cond $X=8.88 $Y=3.135
+ $X2=8.455 $Y2=3.135
r158 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r159 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r160 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r161 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r162 110 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r163 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r164 107 135 11.0851 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=12.915 $Y=3.33
+ $X2=12.672 $Y2=3.33
r165 107 109 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.915 $Y=3.33
+ $X2=13.2 $Y2=3.33
r166 106 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r167 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r168 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r169 103 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r170 102 105 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r171 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r172 100 132 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=10.877 $Y2=3.33
r173 100 102 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=11.04 $Y=3.33
+ $X2=11.28 $Y2=3.33
r174 99 135 11.0851 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=12.43 $Y=3.33
+ $X2=12.672 $Y2=3.33
r175 99 105 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=12.43 $Y=3.33
+ $X2=12.24 $Y2=3.33
r176 98 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r177 98 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r178 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r179 95 129 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.05 $Y=3.33
+ $X2=9.92 $Y2=3.33
r180 95 97 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=10.05 $Y=3.33
+ $X2=10.32 $Y2=3.33
r181 94 132 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=10.715 $Y=3.33
+ $X2=10.877 $Y2=3.33
r182 94 97 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.715 $Y=3.33
+ $X2=10.32 $Y2=3.33
r183 93 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r184 92 124 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=8.455 $Y2=3.33
r185 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r186 90 93 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r187 89 92 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r188 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r189 87 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.435 $Y2=3.33
r190 87 89 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r191 85 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r192 85 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r193 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r194 82 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.195 $Y=3.33
+ $X2=5.03 $Y2=3.33
r195 82 84 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=5.195 $Y=3.33
+ $X2=6 $Y2=3.33
r196 81 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.27 $Y=3.33
+ $X2=6.435 $Y2=3.33
r197 81 84 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.27 $Y=3.33 $X2=6
+ $Y2=3.33
r198 80 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r199 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r200 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r201 77 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r202 76 79 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r203 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r204 74 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.205 $Y2=3.33
r205 74 76 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.6 $Y2=3.33
r206 73 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=5.03 $Y2=3.33
r207 73 79 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=4.56 $Y2=3.33
r208 72 114 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r209 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r210 69 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=3.33
+ $X2=3.205 $Y2=3.33
r211 69 71 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r212 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r213 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r214 64 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r215 63 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r216 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r217 60 90 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r218 60 120 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r219 58 67 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.2 $Y2=3.33
r220 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.485 $Y2=3.33
r221 57 71 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.65 $Y=3.33 $X2=1.68
+ $Y2=3.33
r222 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=1.485 $Y2=3.33
r223 53 56 9.98787 $w=4.83e-07 $l=4.05e-07 $layer=LI1_cond $X=12.672 $Y=2.1
+ $X2=12.672 $Y2=2.505
r224 51 135 1.99554 $w=4.85e-07 $l=8.5e-08 $layer=LI1_cond $X=12.672 $Y=3.245
+ $X2=12.672 $Y2=3.33
r225 51 56 18.2494 $w=4.83e-07 $l=7.4e-07 $layer=LI1_cond $X=12.672 $Y=3.245
+ $X2=12.672 $Y2=2.505
r226 47 132 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=10.877 $Y=3.245
+ $X2=10.877 $Y2=3.33
r227 47 49 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=10.877 $Y=3.245
+ $X2=10.877 $Y2=2.875
r228 43 129 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.92 $Y=3.245
+ $X2=9.92 $Y2=3.33
r229 43 45 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=9.92 $Y=3.245
+ $X2=9.92 $Y2=2.875
r230 41 129 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.79 $Y=3.33
+ $X2=9.92 $Y2=3.33
r231 41 127 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=9.79 $Y=3.33
+ $X2=9.19 $Y2=3.33
r232 37 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=3.245
+ $X2=6.435 $Y2=3.33
r233 37 39 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.435 $Y=3.245
+ $X2=6.435 $Y2=2.755
r234 33 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=3.245
+ $X2=5.03 $Y2=3.33
r235 33 35 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.03 $Y=3.245
+ $X2=5.03 $Y2=2.61
r236 29 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=3.245
+ $X2=3.205 $Y2=3.33
r237 29 31 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=3.205 $Y=3.245
+ $X2=3.205 $Y2=2.77
r238 25 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=3.245
+ $X2=1.485 $Y2=3.33
r239 25 27 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=1.485 $Y=3.245
+ $X2=1.485 $Y2=2.46
r240 8 56 300 $w=1.7e-07 $l=8.04083e-07 $layer=licon1_PDIFF $count=2 $X=12.455
+ $Y=1.835 $X2=12.75 $Y2=2.505
r241 8 53 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=12.455
+ $Y=1.835 $X2=12.595 $Y2=2.1
r242 7 49 600 $w=1.7e-07 $l=1.12641e-06 $layer=licon1_PDIFF $count=1 $X=10.74
+ $Y=1.835 $X2=10.92 $Y2=2.875
r243 6 45 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=9.745
+ $Y=2.665 $X2=9.885 $Y2=2.875
r244 5 126 300 $w=1.7e-07 $l=6.76609e-07 $layer=licon1_PDIFF $count=2 $X=8.48
+ $Y=2.665 $X2=9.025 $Y2=2.96
r245 4 39 600 $w=1.7e-07 $l=9.29677e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.895 $X2=6.435 $Y2=2.755
r246 3 35 600 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_PDIFF $count=1 $X=4.835
+ $Y=2.315 $X2=5.03 $Y2=2.61
r247 2 31 600 $w=1.7e-07 $l=5.33268e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=2.315 $X2=3.205 $Y2=2.77
r248 1 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.345
+ $Y=2.315 $X2=1.485 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%A_380_50# 1 2 3 4 15 17 20 23 26 31 32 34
+ 36
c96 34 0 9.78661e-20 $X=3.72 $Y=2.46
c97 32 0 8.87678e-20 $X=3.582 $Y=0.9
c98 23 0 2.10427e-19 $X=4.015 $Y=0.9
r99 36 38 4.43636 $w=1.98e-07 $l=8e-08 $layer=LI1_cond $X=4.115 $Y=0.82
+ $X2=4.115 $Y2=0.9
r100 26 28 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.155 $Y=0.7 $X2=2.155
+ $Y2=0.9
r101 24 32 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=3.685 $Y=0.9
+ $X2=3.582 $Y2=0.9
r102 23 38 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.015 $Y=0.9 $X2=4.115
+ $Y2=0.9
r103 23 24 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.015 $Y=0.9
+ $X2=3.685 $Y2=0.9
r104 20 34 3.77418 $w=2.45e-07 $l=1.252e-07 $layer=LI1_cond $X=3.582 $Y=2.295
+ $X2=3.652 $Y2=2.39
r105 19 32 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.582 $Y=0.985
+ $X2=3.582 $Y2=0.9
r106 19 20 70.8736 $w=2.03e-07 $l=1.31e-06 $layer=LI1_cond $X=3.582 $Y=0.985
+ $X2=3.582 $Y2=2.295
r107 18 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.44 $Y=2.4
+ $X2=2.275 $Y2=2.4
r108 17 34 2.68609 $w=1.7e-07 $l=1.76929e-07 $layer=LI1_cond $X=3.48 $Y=2.4
+ $X2=3.652 $Y2=2.39
r109 17 18 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.48 $Y=2.4
+ $X2=2.44 $Y2=2.4
r110 16 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=0.9
+ $X2=2.155 $Y2=0.9
r111 15 32 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=3.48 $Y=0.9
+ $X2=3.582 $Y2=0.9
r112 15 16 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=3.48 $Y=0.9
+ $X2=2.32 $Y2=0.9
r113 4 34 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=3.52
+ $Y=2.315 $X2=3.72 $Y2=2.46
r114 3 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.135
+ $Y=2.315 $X2=2.275 $Y2=2.46
r115 2 36 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.595 $X2=4.13 $Y2=0.82
r116 1 26 182 $w=1.7e-07 $l=5.6325e-07 $layer=licon1_NDIFF $count=1 $X=1.9
+ $Y=0.25 $X2=2.155 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%Q 1 2 7 8 9 10 11 12 20
r11 12 36 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=13.22 $Y=2.775
+ $X2=13.22 $Y2=2.91
r12 11 12 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.22 $Y=2.405
+ $X2=13.22 $Y2=2.775
r13 10 11 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=13.22 $Y=1.98
+ $X2=13.22 $Y2=2.405
r14 9 10 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=13.22 $Y=1.665
+ $X2=13.22 $Y2=1.98
r15 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.22 $Y=1.295
+ $X2=13.22 $Y2=1.665
r16 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.22 $Y=0.925
+ $X2=13.22 $Y2=1.295
r17 7 20 21.555 $w=2.68e-07 $l=5.05e-07 $layer=LI1_cond $X=13.22 $Y=0.925
+ $X2=13.22 $Y2=0.42
r18 2 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=13.04
+ $Y=1.835 $X2=13.18 $Y2=2.91
r19 2 10 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.04
+ $Y=1.835 $X2=13.18 $Y2=1.98
r20 1 20 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=13.04
+ $Y=0.235 $X2=13.18 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 49 51 56 77 81 91 92 95 98 101 104
c139 92 0 5.91316e-20 $X=13.2 $Y=0
c140 56 0 1.18827e-19 $X=3.405 $Y=0
c141 25 0 9.02003e-20 $X=3.57 $Y=0.55
c142 2 0 9.64219e-20 $X=3.395 $Y=0.405
r143 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r144 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r145 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r146 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r147 92 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r148 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r149 89 104 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.915 $Y=0
+ $X2=12.745 $Y2=0
r150 89 91 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.915 $Y=0
+ $X2=13.2 $Y2=0
r151 88 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r152 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r153 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.24 $Y2=0
r154 85 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r155 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=0 $X2=12.24
+ $Y2=0
r156 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r157 82 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=10.92 $Y2=0
r158 82 84 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=11.28 $Y2=0
r159 81 104 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.575 $Y=0
+ $X2=12.745 $Y2=0
r160 81 87 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=12.575 $Y=0
+ $X2=12.24 $Y2=0
r161 80 102 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=10.8 $Y2=0
r162 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r163 77 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=10.92 $Y2=0
r164 77 79 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=8.88 $Y2=0
r165 76 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r166 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r167 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r168 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r169 70 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r170 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r171 67 70 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r172 67 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r173 66 69 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r174 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r175 64 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.57
+ $Y2=0
r176 64 66 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=4.08
+ $Y2=0
r177 63 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r178 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r179 60 63 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r180 60 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r181 59 62 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r182 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r183 57 95 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.747 $Y2=0
r184 57 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.2
+ $Y2=0
r185 56 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.57
+ $Y2=0
r186 56 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=0
+ $X2=3.12 $Y2=0
r187 54 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r188 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r189 51 95 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.747
+ $Y2=0
r190 51 53 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.24
+ $Y2=0
r191 49 76 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=8.4
+ $Y2=0
r192 49 73 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.48 $Y2=0
r193 47 75 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.49 $Y=0 $X2=8.4
+ $Y2=0
r194 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.49 $Y=0 $X2=8.655
+ $Y2=0
r195 46 79 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=8.82 $Y=0 $X2=8.88
+ $Y2=0
r196 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.82 $Y=0 $X2=8.655
+ $Y2=0
r197 44 69 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.145 $Y=0 $X2=6
+ $Y2=0
r198 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=0 $X2=6.31
+ $Y2=0
r199 43 72 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.475 $Y=0 $X2=6.48
+ $Y2=0
r200 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.475 $Y=0 $X2=6.31
+ $Y2=0
r201 39 104 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=12.745 $Y=0.085
+ $X2=12.745 $Y2=0
r202 39 41 9.66018 $w=3.38e-07 $l=2.85e-07 $layer=LI1_cond $X=12.745 $Y=0.085
+ $X2=12.745 $Y2=0.37
r203 35 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0
r204 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0.38
r205 31 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.655 $Y=0.085
+ $X2=8.655 $Y2=0
r206 31 33 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=8.655 $Y=0.085
+ $X2=8.655 $Y2=0.8
r207 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.31 $Y=0.085
+ $X2=6.31 $Y2=0
r208 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.31 $Y=0.085
+ $X2=6.31 $Y2=0.515
r209 23 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0
r210 23 25 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0.55
r211 19 95 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.747 $Y=0.085
+ $X2=0.747 $Y2=0
r212 19 21 17.189 $w=2.93e-07 $l=4.4e-07 $layer=LI1_cond $X=0.747 $Y=0.085
+ $X2=0.747 $Y2=0.525
r213 6 41 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=12.53
+ $Y=0.235 $X2=12.75 $Y2=0.37
r214 5 37 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=10.7
+ $Y=0.365 $X2=10.92 $Y2=0.38
r215 4 33 182 $w=1.7e-07 $l=4.00625e-07 $layer=licon1_NDIFF $count=1 $X=8.355
+ $Y=0.565 $X2=8.655 $Y2=0.8
r216 3 29 182 $w=1.7e-07 $l=3.99218e-07 $layer=licon1_NDIFF $count=1 $X=5.935
+ $Y=0.565 $X2=6.31 $Y2=0.515
r217 2 25 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=3.395
+ $Y=0.405 $X2=3.57 $Y2=0.55
r218 1 21 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.37 $X2=0.73 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_1%noxref_24 1 2 7 9 14
c28 7 0 1.6277e-19 $X=2.895 $Y=0.35
r29 14 17 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.06 $Y=0.35
+ $X2=3.06 $Y2=0.53
r30 9 12 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.25 $Y=0.35 $X2=1.25
+ $Y2=0.43
r31 8 9 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.355 $Y=0.35 $X2=1.25
+ $Y2=0.35
r32 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=0.35
+ $X2=3.06 $Y2=0.35
r33 7 8 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=2.895 $Y=0.35
+ $X2=1.355 $Y2=0.35
r34 2 17 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.92
+ $Y=0.405 $X2=3.06 $Y2=0.53
r35 1 12 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.25 $X2=1.25 $Y2=0.43
.ends

