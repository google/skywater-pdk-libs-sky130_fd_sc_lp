* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__buflp_0 A VGND VNB VPB VPWR X
X0 VPWR a_36_120# a_315_446# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_36_120# A a_128_490# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_128_490# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_36_120# A a_123_120# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_315_446# a_36_120# X VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VGND a_36_120# a_287_120# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_123_120# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_287_120# a_36_120# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
