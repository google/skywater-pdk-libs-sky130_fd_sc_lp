* File: sky130_fd_sc_lp__maj3_0.pxi.spice
* Created: Wed Sep  2 09:59:17 2020
* 
x_PM_SKY130_FD_SC_LP__MAJ3_0%A N_A_c_75_n N_A_M1012_g N_A_M1010_g N_A_c_70_n
+ N_A_M1001_g N_A_M1008_g N_A_c_78_n A A N_A_c_73_n N_A_c_74_n
+ PM_SKY130_FD_SC_LP__MAJ3_0%A
x_PM_SKY130_FD_SC_LP__MAJ3_0%B N_B_M1002_g N_B_M1006_g N_B_M1007_g N_B_M1004_g B
+ B N_B_c_123_n PM_SKY130_FD_SC_LP__MAJ3_0%B
x_PM_SKY130_FD_SC_LP__MAJ3_0%C N_C_M1013_g N_C_c_168_n N_C_c_169_n N_C_M1000_g
+ N_C_M1011_g N_C_M1005_g N_C_c_166_n C N_C_c_173_n PM_SKY130_FD_SC_LP__MAJ3_0%C
x_PM_SKY130_FD_SC_LP__MAJ3_0%A_28_431# N_A_28_431#_M1000_s N_A_28_431#_M1002_d
+ N_A_28_431#_M1013_s N_A_28_431#_M1006_d N_A_28_431#_c_223_n
+ N_A_28_431#_M1003_g N_A_28_431#_M1009_g N_A_28_431#_c_225_n
+ N_A_28_431#_c_226_n N_A_28_431#_c_235_n N_A_28_431#_c_236_n
+ N_A_28_431#_c_227_n N_A_28_431#_c_238_n N_A_28_431#_c_239_n
+ N_A_28_431#_c_240_n N_A_28_431#_c_228_n N_A_28_431#_c_229_n
+ N_A_28_431#_c_230_n N_A_28_431#_c_241_n N_A_28_431#_c_231_n
+ PM_SKY130_FD_SC_LP__MAJ3_0%A_28_431#
x_PM_SKY130_FD_SC_LP__MAJ3_0%VPWR N_VPWR_M1012_d N_VPWR_M1005_d N_VPWR_c_325_n
+ N_VPWR_c_326_n N_VPWR_c_327_n VPWR N_VPWR_c_328_n N_VPWR_c_329_n
+ N_VPWR_c_330_n N_VPWR_c_324_n N_VPWR_c_332_n N_VPWR_c_333_n
+ PM_SKY130_FD_SC_LP__MAJ3_0%VPWR
x_PM_SKY130_FD_SC_LP__MAJ3_0%X N_X_M1003_d N_X_M1009_d N_X_c_374_n X X X
+ PM_SKY130_FD_SC_LP__MAJ3_0%X
x_PM_SKY130_FD_SC_LP__MAJ3_0%VGND N_VGND_M1010_d N_VGND_M1011_d N_VGND_c_391_n
+ N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n VGND N_VGND_c_395_n
+ N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n PM_SKY130_FD_SC_LP__MAJ3_0%VGND
cc_1 VNB N_A_M1010_g 0.0205246f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=0.495
cc_2 VNB N_A_c_70_n 0.00412086f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.895
cc_3 VNB N_A_M1001_g 0.0204979f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=0.495
cc_4 VNB N_A_M1008_g 0.00401174f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=2.365
cc_5 VNB N_A_c_73_n 0.0689791f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.07
cc_6 VNB N_A_c_74_n 0.0114923f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.07
cc_7 VNB N_B_M1002_g 0.0194687f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.365
cc_8 VNB N_B_M1006_g 0.00344334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B_M1007_g 0.0203812f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=0.495
cc_10 VNB N_B_M1004_g 0.00392238f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=2.365
cc_11 VNB B 0.0162752f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.97
cc_12 VNB N_B_c_123_n 0.0607769f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_C_M1000_g 0.0562473f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.895
cc_14 VNB N_C_M1011_g 0.0493377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C_c_166_n 0.0201131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_28_431#_c_223_n 0.025238f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.575
cc_17 VNB N_A_28_431#_M1003_g 0.0373418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_28_431#_c_225_n 0.00385357f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_19 VNB N_A_28_431#_c_226_n 0.0460128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_28_431#_c_227_n 0.00671706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_28_431#_c_228_n 0.00387159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_28_431#_c_229_n 0.0184926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_28_431#_c_230_n 0.0371924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_28_431#_c_231_n 0.008423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_324_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_374_n 0.0351671f $X=-0.19 $Y=-0.245 $X2=1.49 $Y2=0.905
cc_27 VNB X 0.050293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_391_n 0.00412757f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.895
cc_29 VNB N_VGND_c_392_n 0.012099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_393_n 0.0340274f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=2.365
cc_31 VNB N_VGND_c_394_n 0.00397464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_395_n 0.0321407f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.97
cc_33 VNB N_VGND_c_396_n 0.0246225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_397_n 0.246063f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.24
cc_35 VNB N_VGND_c_398_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_A_c_75_n 0.0164394f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.045
cc_37 VPB N_A_c_70_n 0.0125095f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.895
cc_38 VPB N_A_M1008_g 0.0345763f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=2.365
cc_39 VPB N_A_c_78_n 0.0236325f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.97
cc_40 VPB N_B_M1006_g 0.0306294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_B_M1004_g 0.0312149f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=2.365
cc_42 VPB N_C_M1013_g 0.0619253f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=0.905
cc_43 VPB N_C_c_168_n 0.155374f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=0.495
cc_44 VPB N_C_c_169_n 0.0155689f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=0.495
cc_45 VPB N_C_M1011_g 0.0336922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_C_c_166_n 0.00422773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB C 0.0172677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_C_c_173_n 0.0440662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_28_431#_M1009_g 0.0232445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_28_431#_c_225_n 0.0145398f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_51 VPB N_A_28_431#_c_226_n 0.00478473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_28_431#_c_235_n 0.0308959f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.07
cc_53 VPB N_A_28_431#_c_236_n 0.0251471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_28_431#_c_227_n 0.0012338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_28_431#_c_238_n 0.00346978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_28_431#_c_239_n 0.0222616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_28_431#_c_240_n 0.00940387f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_28_431#_c_241_n 0.0132078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_325_n 0.0240932f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.895
cc_60 VPB N_VPWR_c_326_n 0.0230304f $X=-0.19 $Y=1.655 $X2=1.49 $Y2=0.495
cc_61 VPB N_VPWR_c_327_n 6.80727e-19 $X=-0.19 $Y=1.655 $X2=1.52 $Y2=2.365
cc_62 VPB N_VPWR_c_328_n 0.0333738f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.97
cc_63 VPB N_VPWR_c_329_n 0.0505532f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_330_n 0.0192183f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.24
cc_65 VPB N_VPWR_c_324_n 0.0627428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_332_n 0.00595541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_333_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB X 0.0426394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 N_A_M1001_g N_B_M1002_g 0.0332194f $X=1.49 $Y=0.495 $X2=0 $Y2=0
cc_70 N_A_M1008_g N_B_M1006_g 0.0387231f $X=1.52 $Y=2.365 $X2=0 $Y2=0
cc_71 N_A_c_73_n N_B_c_123_n 0.0719425f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_72 N_A_c_74_n N_B_c_123_n 6.20639e-19 $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_73 N_A_c_70_n N_C_M1013_g 0.00690307f $X=1.06 $Y=1.895 $X2=0 $Y2=0
cc_74 N_A_c_78_n N_C_M1013_g 0.0486796f $X=1.06 $Y=1.97 $X2=0 $Y2=0
cc_75 N_A_c_75_n N_C_c_168_n 0.00929759f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_76 N_A_M1008_g N_C_c_168_n 0.00929759f $X=1.52 $Y=2.365 $X2=0 $Y2=0
cc_77 N_A_M1010_g N_C_M1000_g 0.0401911f $X=1.06 $Y=0.495 $X2=0 $Y2=0
cc_78 N_A_c_74_n N_C_M1000_g 0.0259622f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_79 N_A_c_73_n N_C_c_166_n 0.0401911f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_80 N_A_c_74_n N_C_c_166_n 0.00360631f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_81 N_A_c_74_n N_A_28_431#_c_226_n 0.0335394f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_82 N_A_c_78_n N_A_28_431#_c_235_n 0.00242745f $X=1.06 $Y=1.97 $X2=0 $Y2=0
cc_83 N_A_c_70_n N_A_28_431#_c_236_n 0.00800457f $X=1.06 $Y=1.895 $X2=0 $Y2=0
cc_84 N_A_M1008_g N_A_28_431#_c_236_n 0.0171048f $X=1.52 $Y=2.365 $X2=0 $Y2=0
cc_85 N_A_c_78_n N_A_28_431#_c_236_n 0.0161388f $X=1.06 $Y=1.97 $X2=0 $Y2=0
cc_86 N_A_c_73_n N_A_28_431#_c_236_n 0.00336371f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_87 N_A_c_74_n N_A_28_431#_c_236_n 0.0695078f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_88 N_A_M1001_g N_A_28_431#_c_227_n 0.00736278f $X=1.49 $Y=0.495 $X2=0 $Y2=0
cc_89 N_A_c_73_n N_A_28_431#_c_227_n 0.00492368f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_90 N_A_c_74_n N_A_28_431#_c_227_n 0.0511081f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_91 N_A_M1008_g N_A_28_431#_c_238_n 0.00238439f $X=1.52 $Y=2.365 $X2=0 $Y2=0
cc_92 N_A_M1010_g N_A_28_431#_c_230_n 0.0012945f $X=1.06 $Y=0.495 $X2=0 $Y2=0
cc_93 N_A_c_74_n N_A_28_431#_c_230_n 0.00116472f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_94 N_A_M1001_g N_A_28_431#_c_231_n 0.00351584f $X=1.49 $Y=0.495 $X2=0 $Y2=0
cc_95 N_A_c_75_n N_VPWR_c_325_n 0.0100714f $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_96 N_A_M1008_g N_VPWR_c_325_n 0.0100714f $X=1.52 $Y=2.365 $X2=0 $Y2=0
cc_97 N_A_c_78_n N_VPWR_c_325_n 0.00335117f $X=1.06 $Y=1.97 $X2=0 $Y2=0
cc_98 N_A_c_75_n N_VPWR_c_324_n 8.12218e-19 $X=0.86 $Y=2.045 $X2=0 $Y2=0
cc_99 N_A_M1008_g N_VPWR_c_324_n 8.12218e-19 $X=1.52 $Y=2.365 $X2=0 $Y2=0
cc_100 N_A_M1010_g N_VGND_c_391_n 0.0128622f $X=1.06 $Y=0.495 $X2=0 $Y2=0
cc_101 N_A_M1001_g N_VGND_c_391_n 0.0107512f $X=1.49 $Y=0.495 $X2=0 $Y2=0
cc_102 N_A_c_73_n N_VGND_c_391_n 0.00266929f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_103 N_A_c_74_n N_VGND_c_391_n 0.027631f $X=1.35 $Y=1.07 $X2=0 $Y2=0
cc_104 N_A_M1001_g N_VGND_c_393_n 0.00445056f $X=1.49 $Y=0.495 $X2=0 $Y2=0
cc_105 N_A_M1010_g N_VGND_c_395_n 0.00445056f $X=1.06 $Y=0.495 $X2=0 $Y2=0
cc_106 N_A_M1010_g N_VGND_c_397_n 0.00804604f $X=1.06 $Y=0.495 $X2=0 $Y2=0
cc_107 N_A_M1001_g N_VGND_c_397_n 0.00804604f $X=1.49 $Y=0.495 $X2=0 $Y2=0
cc_108 N_B_M1006_g N_C_c_168_n 0.00917428f $X=1.88 $Y=2.365 $X2=0 $Y2=0
cc_109 N_B_M1004_g N_C_c_168_n 0.00917428f $X=2.31 $Y=2.365 $X2=0 $Y2=0
cc_110 N_B_M1007_g N_C_M1011_g 0.157788f $X=2.31 $Y=0.495 $X2=0 $Y2=0
cc_111 B N_C_M1011_g 0.0258531f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B_M1004_g C 0.00110422f $X=2.31 $Y=2.365 $X2=0 $Y2=0
cc_113 B N_A_28_431#_M1003_g 0.00485878f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B_M1002_g N_A_28_431#_c_227_n 0.00487611f $X=1.88 $Y=0.495 $X2=0 $Y2=0
cc_115 N_B_M1006_g N_A_28_431#_c_227_n 0.00455805f $X=1.88 $Y=2.365 $X2=0 $Y2=0
cc_116 N_B_M1007_g N_A_28_431#_c_227_n 9.41713e-19 $X=2.31 $Y=0.495 $X2=0 $Y2=0
cc_117 N_B_M1004_g N_A_28_431#_c_227_n 9.41713e-19 $X=2.31 $Y=2.365 $X2=0 $Y2=0
cc_118 B N_A_28_431#_c_227_n 0.0487691f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_119 N_B_c_123_n N_A_28_431#_c_227_n 0.0165892f $X=2.21 $Y=1.07 $X2=0 $Y2=0
cc_120 N_B_M1006_g N_A_28_431#_c_238_n 0.0156315f $X=1.88 $Y=2.365 $X2=0 $Y2=0
cc_121 N_B_M1004_g N_A_28_431#_c_238_n 0.0156117f $X=2.31 $Y=2.365 $X2=0 $Y2=0
cc_122 N_B_M1004_g N_A_28_431#_c_239_n 0.010699f $X=2.31 $Y=2.365 $X2=0 $Y2=0
cc_123 N_B_M1006_g N_A_28_431#_c_240_n 0.0157438f $X=1.88 $Y=2.365 $X2=0 $Y2=0
cc_124 N_B_M1004_g N_A_28_431#_c_240_n 0.00283017f $X=2.31 $Y=2.365 $X2=0 $Y2=0
cc_125 B N_A_28_431#_c_240_n 0.0538656f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B_c_123_n N_A_28_431#_c_240_n 0.00257849f $X=2.21 $Y=1.07 $X2=0 $Y2=0
cc_127 B N_A_28_431#_c_228_n 0.0351049f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_128 B N_A_28_431#_c_229_n 0.00293095f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B_M1002_g N_A_28_431#_c_231_n 0.0156057f $X=1.88 $Y=0.495 $X2=0 $Y2=0
cc_130 N_B_M1007_g N_A_28_431#_c_231_n 0.00867914f $X=2.31 $Y=0.495 $X2=0 $Y2=0
cc_131 B N_A_28_431#_c_231_n 0.017517f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B_c_123_n N_A_28_431#_c_231_n 0.00263677f $X=2.21 $Y=1.07 $X2=0 $Y2=0
cc_133 N_B_M1006_g N_VPWR_c_324_n 8.12218e-19 $X=1.88 $Y=2.365 $X2=0 $Y2=0
cc_134 N_B_M1004_g N_VPWR_c_324_n 8.12218e-19 $X=2.31 $Y=2.365 $X2=0 $Y2=0
cc_135 N_B_M1002_g N_VGND_c_391_n 0.0012465f $X=1.88 $Y=0.495 $X2=0 $Y2=0
cc_136 N_B_M1007_g N_VGND_c_392_n 0.00210322f $X=2.31 $Y=0.495 $X2=0 $Y2=0
cc_137 B N_VGND_c_392_n 0.00282302f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_138 N_B_M1002_g N_VGND_c_393_n 0.00327726f $X=1.88 $Y=0.495 $X2=0 $Y2=0
cc_139 N_B_M1007_g N_VGND_c_393_n 0.00501304f $X=2.31 $Y=0.495 $X2=0 $Y2=0
cc_140 N_B_M1002_g N_VGND_c_397_n 0.00481846f $X=1.88 $Y=0.495 $X2=0 $Y2=0
cc_141 N_B_M1007_g N_VGND_c_397_n 0.00939373f $X=2.31 $Y=0.495 $X2=0 $Y2=0
cc_142 N_C_M1011_g N_A_28_431#_M1003_g 0.025307f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_143 N_C_M1011_g N_A_28_431#_M1009_g 0.0202985f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_144 N_C_M1000_g N_A_28_431#_c_226_n 0.0158852f $X=0.67 $Y=0.495 $X2=0 $Y2=0
cc_145 N_C_c_166_n N_A_28_431#_c_226_n 0.00839044f $X=0.67 $Y=1.58 $X2=0 $Y2=0
cc_146 N_C_M1013_g N_A_28_431#_c_235_n 0.0180376f $X=0.5 $Y=2.365 $X2=0 $Y2=0
cc_147 N_C_M1013_g N_A_28_431#_c_236_n 0.0147704f $X=0.5 $Y=2.365 $X2=0 $Y2=0
cc_148 N_C_c_166_n N_A_28_431#_c_236_n 0.00521054f $X=0.67 $Y=1.58 $X2=0 $Y2=0
cc_149 N_C_c_168_n N_A_28_431#_c_238_n 0.00600475f $X=2.595 $Y=3.02 $X2=0 $Y2=0
cc_150 N_C_M1011_g N_A_28_431#_c_238_n 0.00257113f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_151 N_C_M1011_g N_A_28_431#_c_239_n 0.0150768f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_152 N_C_M1011_g N_A_28_431#_c_228_n 0.00178277f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_153 N_C_M1011_g N_A_28_431#_c_229_n 0.0422703f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_154 N_C_M1000_g N_A_28_431#_c_230_n 0.0100528f $X=0.67 $Y=0.495 $X2=0 $Y2=0
cc_155 N_C_M1013_g N_A_28_431#_c_241_n 0.0049947f $X=0.5 $Y=2.365 $X2=0 $Y2=0
cc_156 N_C_M1011_g N_A_28_431#_c_231_n 0.00124336f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_157 N_C_M1013_g N_VPWR_c_325_n 0.0074879f $X=0.5 $Y=2.365 $X2=0 $Y2=0
cc_158 N_C_c_168_n N_VPWR_c_325_n 0.0327904f $X=2.595 $Y=3.02 $X2=0 $Y2=0
cc_159 N_C_M1011_g N_VPWR_c_326_n 0.00201006f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_160 C N_VPWR_c_326_n 0.0299087f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_161 N_C_c_173_n N_VPWR_c_326_n 0.00893458f $X=2.76 $Y=2.9 $X2=0 $Y2=0
cc_162 N_C_M1011_g N_VPWR_c_327_n 0.00537229f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_163 C N_VPWR_c_327_n 0.00660146f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_164 N_C_c_173_n N_VPWR_c_327_n 5.13949e-19 $X=2.76 $Y=2.9 $X2=0 $Y2=0
cc_165 N_C_c_169_n N_VPWR_c_328_n 0.0173226f $X=0.575 $Y=3.02 $X2=0 $Y2=0
cc_166 N_C_c_168_n N_VPWR_c_329_n 0.037424f $X=2.595 $Y=3.02 $X2=0 $Y2=0
cc_167 C N_VPWR_c_329_n 0.0245092f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_168 N_C_c_168_n N_VPWR_c_324_n 0.0688504f $X=2.595 $Y=3.02 $X2=0 $Y2=0
cc_169 N_C_c_169_n N_VPWR_c_324_n 0.00844206f $X=0.575 $Y=3.02 $X2=0 $Y2=0
cc_170 C N_VPWR_c_324_n 0.0133281f $X=2.555 $Y=2.69 $X2=0 $Y2=0
cc_171 N_C_c_173_n N_VPWR_c_324_n 0.00767005f $X=2.76 $Y=2.9 $X2=0 $Y2=0
cc_172 N_C_M1000_g N_VGND_c_391_n 0.00213595f $X=0.67 $Y=0.495 $X2=0 $Y2=0
cc_173 N_C_M1011_g N_VGND_c_392_n 0.0120232f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_174 N_C_M1011_g N_VGND_c_393_n 0.00445056f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_175 N_C_M1000_g N_VGND_c_395_n 0.00501304f $X=0.67 $Y=0.495 $X2=0 $Y2=0
cc_176 N_C_M1000_g N_VGND_c_397_n 0.0101917f $X=0.67 $Y=0.495 $X2=0 $Y2=0
cc_177 N_C_M1011_g N_VGND_c_397_n 0.0079903f $X=2.67 $Y=0.495 $X2=0 $Y2=0
cc_178 N_A_28_431#_c_235_n N_VPWR_c_325_n 0.0137622f $X=0.285 $Y=2.365 $X2=0
+ $Y2=0
cc_179 N_A_28_431#_c_236_n N_VPWR_c_325_n 0.0234462f $X=1.695 $Y=1.84 $X2=0
+ $Y2=0
cc_180 N_A_28_431#_c_238_n N_VPWR_c_325_n 0.0137622f $X=2.095 $Y=2.365 $X2=0
+ $Y2=0
cc_181 N_A_28_431#_M1009_g N_VPWR_c_326_n 0.0124083f $X=3.22 $Y=2.255 $X2=0
+ $Y2=0
cc_182 N_A_28_431#_M1009_g N_VPWR_c_327_n 0.00901099f $X=3.22 $Y=2.255 $X2=0
+ $Y2=0
cc_183 N_A_28_431#_c_225_n N_VPWR_c_327_n 8.61336e-19 $X=3.125 $Y=1.775 $X2=0
+ $Y2=0
cc_184 N_A_28_431#_c_238_n N_VPWR_c_327_n 0.0113777f $X=2.095 $Y=2.365 $X2=0
+ $Y2=0
cc_185 N_A_28_431#_c_239_n N_VPWR_c_327_n 0.0323691f $X=2.955 $Y=1.84 $X2=0
+ $Y2=0
cc_186 N_A_28_431#_c_235_n N_VPWR_c_328_n 0.00541334f $X=0.285 $Y=2.365 $X2=0
+ $Y2=0
cc_187 N_A_28_431#_c_238_n N_VPWR_c_329_n 0.00533533f $X=2.095 $Y=2.365 $X2=0
+ $Y2=0
cc_188 N_A_28_431#_M1009_g N_VPWR_c_330_n 4.63495e-19 $X=3.22 $Y=2.255 $X2=0
+ $Y2=0
cc_189 N_A_28_431#_M1009_g N_VPWR_c_324_n 6.08924e-19 $X=3.22 $Y=2.255 $X2=0
+ $Y2=0
cc_190 N_A_28_431#_c_235_n N_VPWR_c_324_n 0.00911923f $X=0.285 $Y=2.365 $X2=0
+ $Y2=0
cc_191 N_A_28_431#_c_238_n N_VPWR_c_324_n 0.00790535f $X=2.095 $Y=2.365 $X2=0
+ $Y2=0
cc_192 N_A_28_431#_M1003_g N_X_c_374_n 0.00706665f $X=3.1 $Y=0.495 $X2=0 $Y2=0
cc_193 N_A_28_431#_c_228_n N_X_c_374_n 0.00620631f $X=3.12 $Y=1.27 $X2=0 $Y2=0
cc_194 N_A_28_431#_c_229_n N_X_c_374_n 0.00112824f $X=3.12 $Y=1.27 $X2=0 $Y2=0
cc_195 N_A_28_431#_M1003_g X 0.0119667f $X=3.1 $Y=0.495 $X2=0 $Y2=0
cc_196 N_A_28_431#_c_239_n X 0.0133392f $X=2.955 $Y=1.84 $X2=0 $Y2=0
cc_197 N_A_28_431#_c_228_n X 0.0481012f $X=3.12 $Y=1.27 $X2=0 $Y2=0
cc_198 N_A_28_431#_c_229_n X 0.0342531f $X=3.12 $Y=1.27 $X2=0 $Y2=0
cc_199 N_A_28_431#_c_230_n N_VGND_c_391_n 0.0150171f $X=0.455 $Y=0.495 $X2=0
+ $Y2=0
cc_200 N_A_28_431#_c_231_n N_VGND_c_391_n 0.0273445f $X=2.095 $Y=0.495 $X2=0
+ $Y2=0
cc_201 N_A_28_431#_M1003_g N_VGND_c_392_n 0.00286943f $X=3.1 $Y=0.495 $X2=0
+ $Y2=0
cc_202 N_A_28_431#_c_228_n N_VGND_c_392_n 6.34075e-19 $X=3.12 $Y=1.27 $X2=0
+ $Y2=0
cc_203 N_A_28_431#_c_231_n N_VGND_c_392_n 0.0156946f $X=2.095 $Y=0.495 $X2=0
+ $Y2=0
cc_204 N_A_28_431#_c_231_n N_VGND_c_393_n 0.0361968f $X=2.095 $Y=0.495 $X2=0
+ $Y2=0
cc_205 N_A_28_431#_c_230_n N_VGND_c_395_n 0.0324583f $X=0.455 $Y=0.495 $X2=0
+ $Y2=0
cc_206 N_A_28_431#_M1003_g N_VGND_c_396_n 0.00501304f $X=3.1 $Y=0.495 $X2=0
+ $Y2=0
cc_207 N_A_28_431#_M1003_g N_VGND_c_397_n 0.010164f $X=3.1 $Y=0.495 $X2=0 $Y2=0
cc_208 N_A_28_431#_c_230_n N_VGND_c_397_n 0.0190199f $X=0.455 $Y=0.495 $X2=0
+ $Y2=0
cc_209 N_A_28_431#_c_231_n N_VGND_c_397_n 0.0208169f $X=2.095 $Y=0.495 $X2=0
+ $Y2=0
cc_210 N_A_28_431#_c_231_n A_313_57# 0.00422865f $X=2.095 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_211 N_VPWR_c_326_n X 0.00766846f $X=3.19 $Y=3.245 $X2=0 $Y2=0
cc_212 N_VPWR_c_327_n X 0.0266866f $X=3.19 $Y=2.292 $X2=0 $Y2=0
cc_213 N_VPWR_c_330_n X 0.00413386f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_c_324_n X 0.00698862f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_215 N_X_c_374_n N_VGND_c_392_n 0.019296f $X=3.59 $Y=0.495 $X2=0 $Y2=0
cc_216 N_X_c_374_n N_VGND_c_396_n 0.0366886f $X=3.59 $Y=0.495 $X2=0 $Y2=0
cc_217 N_X_c_374_n N_VGND_c_397_n 0.0215075f $X=3.59 $Y=0.495 $X2=0 $Y2=0
