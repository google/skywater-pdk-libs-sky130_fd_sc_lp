* File: sky130_fd_sc_lp__a22oi_2.spice
* Created: Wed Sep  2 09:23:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22oi_2.pex.spice"
.subckt sky130_fd_sc_lp__a22oi_2  VNB VPB A1 A2 B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A1_M1002_g N_A_179_47#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.7 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_179_47#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1848 AS=0.1176 PD=1.28 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1007_d N_A2_M1009_g N_A_179_47#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1848 AS=0.1176 PD=1.28 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75002.6 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A1_M1003_g N_A_179_47#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2016 AS=0.1176 PD=1.32 PS=1.12 NRD=12.852 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1008 N_A_595_47#_M1008_d N_B1_M1008_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.2016 PD=1.23 PS=1.32 NRD=4.284 NRS=15.708 M=1 R=5.6 SA=75002.3
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1006 N_A_595_47#_M1008_d N_B2_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1176 PD=1.23 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1012 N_A_595_47#_M1012_d N_B2_M1012_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1011 N_A_595_47#_M1012_d N_B1_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_49_367#_M1004_d N_A1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.31185 PD=3.05 PS=1.755 NRD=0 NRS=17.9664 M=1 R=8.4 SA=75000.2
+ SB=75003.9 A=0.189 P=2.82 MULT=1
MM1001 N_A_49_367#_M1001_d N_A2_M1001_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.31185 PD=1.54 PS=1.755 NRD=0 NRS=15.6221 M=1 R=8.4 SA=75000.8
+ SB=75003.3 A=0.189 P=2.82 MULT=1
MM1013 N_A_49_367#_M1001_d N_A2_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.473675 PD=1.54 PS=2.085 NRD=0 NRS=29.3136 M=1 R=8.4 SA=75001.3
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1014 N_A_49_367#_M1014_d N_A1_M1014_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.473675 PD=1.54 PS=2.085 NRD=0 NRS=41.8231 M=1 R=8.4 SA=75002.1
+ SB=75002 A=0.189 P=2.82 MULT=1
MM1000 N_A_49_367#_M1014_d N_B1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=6.2449 M=1 R=8.4 SA=75002.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1000_s N_B2_M1005_g N_A_49_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003 SB=75001.1
+ A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1010_d N_B2_M1010_g N_A_49_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1015 N_A_49_367#_M1015_d N_B1_M1015_g N_Y_M1010_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__a22oi_2.pxi.spice"
*
.ends
*
*
