* File: sky130_fd_sc_lp__mux2i_m.pxi.spice
* Created: Wed Sep  2 10:01:37 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2I_M%S N_S_M1004_g N_S_M1005_g N_S_c_76_n N_S_M1000_g
+ N_S_c_83_n N_S_M1003_g N_S_c_77_n N_S_c_78_n N_S_c_85_n N_S_c_86_n N_S_c_87_n
+ N_S_c_88_n N_S_c_98_p N_S_c_89_n N_S_c_90_n N_S_c_141_p N_S_c_91_n N_S_c_92_n
+ S S S N_S_c_80_n PM_SKY130_FD_SC_LP__MUX2I_M%S
x_PM_SKY130_FD_SC_LP__MUX2I_M%A_55_125# N_A_55_125#_M1004_s N_A_55_125#_M1005_s
+ N_A_55_125#_M1008_g N_A_55_125#_M1006_g N_A_55_125#_c_193_n
+ N_A_55_125#_c_194_n N_A_55_125#_c_187_n N_A_55_125#_c_195_n
+ N_A_55_125#_c_188_n N_A_55_125#_c_189_n N_A_55_125#_c_198_n
+ N_A_55_125#_c_199_n N_A_55_125#_c_190_n N_A_55_125#_c_191_n
+ PM_SKY130_FD_SC_LP__MUX2I_M%A_55_125#
x_PM_SKY130_FD_SC_LP__MUX2I_M%A1 N_A1_M1001_g N_A1_M1009_g N_A1_c_250_n
+ N_A1_c_251_n N_A1_c_252_n A1 A1 A1 N_A1_c_259_n N_A1_c_255_n N_A1_c_256_n
+ PM_SKY130_FD_SC_LP__MUX2I_M%A1
x_PM_SKY130_FD_SC_LP__MUX2I_M%A0 N_A0_M1007_g N_A0_c_320_n N_A0_c_321_n
+ N_A0_c_322_n N_A0_M1002_g A0 PM_SKY130_FD_SC_LP__MUX2I_M%A0
x_PM_SKY130_FD_SC_LP__MUX2I_M%VPWR N_VPWR_M1005_d N_VPWR_M1003_d N_VPWR_c_371_n
+ N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_375_n VPWR
+ N_VPWR_c_376_n N_VPWR_c_370_n PM_SKY130_FD_SC_LP__MUX2I_M%VPWR
x_PM_SKY130_FD_SC_LP__MUX2I_M%Y N_Y_M1007_d N_Y_M1001_d N_Y_c_411_n N_Y_c_412_n
+ N_Y_c_413_n N_Y_c_408_n N_Y_c_409_n N_Y_c_434_n Y
+ PM_SKY130_FD_SC_LP__MUX2I_M%Y
x_PM_SKY130_FD_SC_LP__MUX2I_M%VGND N_VGND_M1004_d N_VGND_M1000_d N_VGND_c_475_n
+ N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n VGND N_VGND_c_479_n
+ N_VGND_c_480_n N_VGND_c_481_n N_VGND_c_482_n PM_SKY130_FD_SC_LP__MUX2I_M%VGND
cc_1 VNB N_S_M1004_g 0.0518629f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.835
cc_2 VNB N_S_c_76_n 0.0203027f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=1.155
cc_3 VNB N_S_c_77_n 0.0309262f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.23
cc_4 VNB N_S_c_78_n 0.0129426f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.23
cc_5 VNB S 0.0301596f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.21
cc_6 VNB N_S_c_80_n 0.0291475f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=1.32
cc_7 VNB N_A_55_125#_M1008_g 0.0326581f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=1.155
cc_8 VNB N_A_55_125#_c_187_n 0.0209742f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=1.66
cc_9 VNB N_A_55_125#_c_188_n 0.0068201f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.16
cc_10 VNB N_A_55_125#_c_189_n 0.0210702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_55_125#_c_190_n 0.0108174f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=2.41
cc_12 VNB N_A_55_125#_c_191_n 0.0108135f $X=-0.19 $Y=-0.245 $X2=3.047 $Y2=2.325
cc_13 VNB N_A1_c_250_n 0.00350568f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=0.835
cc_14 VNB N_A1_c_251_n 0.0099885f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.975
cc_15 VNB N_A1_c_252_n 0.0466524f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.695
cc_16 VNB A1 0.0139825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A1 0.00222741f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.23
cc_18 VNB N_A1_c_255_n 0.0161728f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.385
cc_19 VNB N_A1_c_256_n 0.00369457f $X=-0.19 $Y=-0.245 $X2=3.047 $Y2=2.325
cc_20 VNB N_A0_M1007_g 0.0262554f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.835
cc_21 VNB N_A0_c_320_n 0.0260199f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.325
cc_22 VNB N_A0_c_321_n 0.0104248f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.695
cc_23 VNB N_A0_c_322_n 0.0233601f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.695
cc_24 VNB N_VPWR_c_370_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.38 $Y2=2.495
cc_25 VNB N_Y_c_408_n 0.0180375f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=0.835
cc_26 VNB N_Y_c_409_n 0.00942702f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.695
cc_27 VNB Y 0.00233508f $X=-0.19 $Y=-0.245 $X2=2.975 $Y2=1.66
cc_28 VNB N_VGND_c_475_n 0.0254251f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=1.155
cc_29 VNB N_VGND_c_476_n 0.0352133f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.695
cc_30 VNB N_VGND_c_477_n 0.0258507f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.23
cc_31 VNB N_VGND_c_478_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.23
cc_32 VNB N_VGND_c_479_n 0.0407669f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.16
cc_33 VNB N_VGND_c_480_n 0.0158267f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=2.895
cc_34 VNB N_VGND_c_481_n 0.237989f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=2.98
cc_35 VNB N_VGND_c_482_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.38 $Y2=2.895
cc_36 VPB N_S_M1004_g 0.0202468f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.835
cc_37 VPB N_S_M1005_g 0.0246896f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.695
cc_38 VPB N_S_c_83_n 0.0420398f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=1.975
cc_39 VPB N_S_M1003_g 0.0402656f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.695
cc_40 VPB N_S_c_85_n 4.13128e-19 $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.16
cc_41 VPB N_S_c_86_n 0.0362168f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.16
cc_42 VPB N_S_c_87_n 0.0132434f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.385
cc_43 VPB N_S_c_88_n 0.00228669f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.385
cc_44 VPB N_S_c_89_n 0.00909982f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=2.98
cc_45 VPB N_S_c_90_n 0.00232339f $X=-0.19 $Y=1.655 $X2=1.505 $Y2=2.98
cc_46 VPB N_S_c_91_n 0.0137071f $X=-0.19 $Y=1.655 $X2=2.89 $Y2=2.41
cc_47 VPB N_S_c_92_n 0.00298641f $X=-0.19 $Y=1.655 $X2=2.465 $Y2=2.41
cc_48 VPB S 0.0299356f $X=-0.19 $Y=1.655 $X2=3.035 $Y2=1.21
cc_49 VPB N_A_55_125#_M1006_g 0.0266762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_55_125#_c_193_n 0.0134965f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=1.23
cc_51 VPB N_A_55_125#_c_194_n 0.010897f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=1.975
cc_52 VPB N_A_55_125#_c_195_n 0.0433817f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.3
cc_53 VPB N_A_55_125#_c_188_n 0.00787718f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.16
cc_54 VPB N_A_55_125#_c_189_n 0.0125329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_55_125#_c_198_n 0.0112073f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.385
cc_56 VPB N_A_55_125#_c_199_n 7.44524e-19 $X=-0.19 $Y=1.655 $X2=1.42 $Y2=2.895
cc_57 VPB N_A_55_125#_c_191_n 0.00470152f $X=-0.19 $Y=1.655 $X2=3.047 $Y2=2.325
cc_58 VPB N_A1_M1001_g 0.0305687f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.835
cc_59 VPB A1 0.0101506f $X=-0.19 $Y=1.655 $X2=2.81 $Y2=1.23
cc_60 VPB N_A1_c_259_n 0.0303388f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.3
cc_61 VPB N_A0_c_322_n 0.021733f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.695
cc_62 VPB N_A0_M1002_g 0.0427869f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=1.155
cc_63 VPB N_VPWR_c_371_n 0.0100304f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=1.155
cc_64 VPB N_VPWR_c_372_n 0.0161782f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=0.835
cc_65 VPB N_VPWR_c_373_n 0.0262448f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.695
cc_66 VPB N_VPWR_c_374_n 0.025469f $X=-0.19 $Y=1.655 $X2=2.81 $Y2=1.23
cc_67 VPB N_VPWR_c_375_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=1.23
cc_68 VPB N_VPWR_c_376_n 0.0415546f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.16
cc_69 VPB N_VPWR_c_370_n 0.0742372f $X=-0.19 $Y=1.655 $X2=2.38 $Y2=2.495
cc_70 VPB N_Y_c_411_n 0.00330766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_Y_c_412_n 0.00924924f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=1.155
cc_72 VPB N_Y_c_413_n 0.00283826f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=0.835
cc_73 VPB N_Y_c_409_n 0.00398867f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.695
cc_74 N_S_M1004_g N_A_55_125#_M1008_g 0.0218964f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_75 N_S_c_85_n N_A_55_125#_M1006_g 7.90629e-19 $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_76 N_S_c_86_n N_A_55_125#_M1006_g 0.0227743f $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_77 N_S_c_87_n N_A_55_125#_M1006_g 0.0153286f $X=1.335 $Y=2.385 $X2=0 $Y2=0
cc_78 N_S_c_98_p N_A_55_125#_M1006_g 0.00163774f $X=1.42 $Y=2.895 $X2=0 $Y2=0
cc_79 N_S_c_90_n N_A_55_125#_M1006_g 9.8105e-19 $X=1.505 $Y=2.98 $X2=0 $Y2=0
cc_80 N_S_M1004_g N_A_55_125#_c_193_n 0.00796992f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_81 N_S_c_85_n N_A_55_125#_c_194_n 5.7537e-19 $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_82 N_S_c_86_n N_A_55_125#_c_194_n 0.00561827f $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_83 N_S_c_87_n N_A_55_125#_c_194_n 9.23898e-19 $X=1.335 $Y=2.385 $X2=0 $Y2=0
cc_84 N_S_M1004_g N_A_55_125#_c_187_n 0.0129694f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_85 N_S_M1004_g N_A_55_125#_c_195_n 0.007754f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_86 N_S_M1005_g N_A_55_125#_c_195_n 0.00490306f $X=0.695 $Y=2.695 $X2=0 $Y2=0
cc_87 N_S_c_85_n N_A_55_125#_c_195_n 0.0208633f $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_88 N_S_c_86_n N_A_55_125#_c_195_n 0.00808144f $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_89 N_S_c_88_n N_A_55_125#_c_195_n 0.0136718f $X=0.69 $Y=2.385 $X2=0 $Y2=0
cc_90 N_S_M1004_g N_A_55_125#_c_188_n 0.0243263f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_91 N_S_c_85_n N_A_55_125#_c_188_n 0.0100463f $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_92 N_S_c_86_n N_A_55_125#_c_188_n 0.00502734f $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_93 N_S_c_87_n N_A_55_125#_c_188_n 0.0153744f $X=1.335 $Y=2.385 $X2=0 $Y2=0
cc_94 N_S_M1004_g N_A_55_125#_c_189_n 0.0213329f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_95 N_S_c_87_n N_A_55_125#_c_189_n 0.00303138f $X=1.335 $Y=2.385 $X2=0 $Y2=0
cc_96 N_S_M1005_g N_A_55_125#_c_199_n 0.00283645f $X=0.695 $Y=2.695 $X2=0 $Y2=0
cc_97 N_S_c_86_n N_A_55_125#_c_199_n 0.00300031f $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_98 N_S_c_88_n N_A_55_125#_c_199_n 0.0072764f $X=0.69 $Y=2.385 $X2=0 $Y2=0
cc_99 N_S_M1004_g N_A_55_125#_c_190_n 0.00316375f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_100 N_S_c_87_n N_A1_M1001_g 0.00446609f $X=1.335 $Y=2.385 $X2=0 $Y2=0
cc_101 N_S_c_98_p N_A1_M1001_g 0.00871927f $X=1.42 $Y=2.895 $X2=0 $Y2=0
cc_102 N_S_c_89_n N_A1_M1001_g 0.0119783f $X=2.295 $Y=2.98 $X2=0 $Y2=0
cc_103 N_S_c_90_n N_A1_M1001_g 0.00122434f $X=1.505 $Y=2.98 $X2=0 $Y2=0
cc_104 N_S_c_76_n N_A1_c_252_n 8.26e-19 $X=2.55 $Y=1.155 $X2=0 $Y2=0
cc_105 N_S_c_85_n A1 0.00338609f $X=0.605 $Y=2.16 $X2=0 $Y2=0
cc_106 N_S_c_87_n A1 0.0132659f $X=1.335 $Y=2.385 $X2=0 $Y2=0
cc_107 N_S_c_76_n N_A1_c_255_n 0.0182877f $X=2.55 $Y=1.155 $X2=0 $Y2=0
cc_108 N_S_c_83_n N_A0_c_322_n 0.00313324f $X=2.645 $Y=1.975 $X2=0 $Y2=0
cc_109 N_S_c_80_n N_A0_c_322_n 0.0054627f $X=2.975 $Y=1.32 $X2=0 $Y2=0
cc_110 N_S_c_83_n N_A0_M1002_g 0.0400342f $X=2.645 $Y=1.975 $X2=0 $Y2=0
cc_111 N_S_c_98_p N_A0_M1002_g 9.65411e-19 $X=1.42 $Y=2.895 $X2=0 $Y2=0
cc_112 N_S_c_89_n N_A0_M1002_g 0.0142058f $X=2.295 $Y=2.98 $X2=0 $Y2=0
cc_113 N_S_c_92_n N_A0_M1002_g 0.0014918f $X=2.465 $Y=2.41 $X2=0 $Y2=0
cc_114 N_S_c_91_n N_VPWR_M1003_d 0.00355458f $X=2.89 $Y=2.41 $X2=0 $Y2=0
cc_115 N_S_M1005_g N_VPWR_c_371_n 0.00494176f $X=0.695 $Y=2.695 $X2=0 $Y2=0
cc_116 N_S_c_87_n N_VPWR_c_371_n 0.0221854f $X=1.335 $Y=2.385 $X2=0 $Y2=0
cc_117 N_S_c_90_n N_VPWR_c_371_n 0.0133632f $X=1.505 $Y=2.98 $X2=0 $Y2=0
cc_118 N_S_c_83_n N_VPWR_c_373_n 3.37915e-19 $X=2.645 $Y=1.975 $X2=0 $Y2=0
cc_119 N_S_M1003_g N_VPWR_c_373_n 0.00879194f $X=2.645 $Y=2.695 $X2=0 $Y2=0
cc_120 N_S_c_89_n N_VPWR_c_373_n 0.00952362f $X=2.295 $Y=2.98 $X2=0 $Y2=0
cc_121 N_S_c_141_p N_VPWR_c_373_n 0.0104107f $X=2.38 $Y=2.895 $X2=0 $Y2=0
cc_122 N_S_c_91_n N_VPWR_c_373_n 0.0268203f $X=2.89 $Y=2.41 $X2=0 $Y2=0
cc_123 N_S_M1005_g N_VPWR_c_374_n 0.00514239f $X=0.695 $Y=2.695 $X2=0 $Y2=0
cc_124 N_S_M1003_g N_VPWR_c_376_n 0.00537957f $X=2.645 $Y=2.695 $X2=0 $Y2=0
cc_125 N_S_c_89_n N_VPWR_c_376_n 0.0593089f $X=2.295 $Y=2.98 $X2=0 $Y2=0
cc_126 N_S_c_90_n N_VPWR_c_376_n 0.0114622f $X=1.505 $Y=2.98 $X2=0 $Y2=0
cc_127 N_S_M1005_g N_VPWR_c_370_n 0.00528353f $X=0.695 $Y=2.695 $X2=0 $Y2=0
cc_128 N_S_M1003_g N_VPWR_c_370_n 0.00528353f $X=2.645 $Y=2.695 $X2=0 $Y2=0
cc_129 N_S_c_87_n N_VPWR_c_370_n 0.011097f $X=1.335 $Y=2.385 $X2=0 $Y2=0
cc_130 N_S_c_88_n N_VPWR_c_370_n 0.00172654f $X=0.69 $Y=2.385 $X2=0 $Y2=0
cc_131 N_S_c_89_n N_VPWR_c_370_n 0.0360943f $X=2.295 $Y=2.98 $X2=0 $Y2=0
cc_132 N_S_c_90_n N_VPWR_c_370_n 0.00657784f $X=1.505 $Y=2.98 $X2=0 $Y2=0
cc_133 N_S_c_91_n N_VPWR_c_370_n 0.0153667f $X=2.89 $Y=2.41 $X2=0 $Y2=0
cc_134 N_S_c_89_n N_Y_M1001_d 0.00429432f $X=2.295 $Y=2.98 $X2=0 $Y2=0
cc_135 N_S_M1003_g N_Y_c_411_n 9.71648e-19 $X=2.645 $Y=2.695 $X2=0 $Y2=0
cc_136 N_S_c_87_n N_Y_c_411_n 0.00662267f $X=1.335 $Y=2.385 $X2=0 $Y2=0
cc_137 N_S_c_98_p N_Y_c_411_n 0.00185951f $X=1.42 $Y=2.895 $X2=0 $Y2=0
cc_138 N_S_c_92_n N_Y_c_411_n 0.0126451f $X=2.465 $Y=2.41 $X2=0 $Y2=0
cc_139 N_S_M1003_g N_Y_c_412_n 0.00735882f $X=2.645 $Y=2.695 $X2=0 $Y2=0
cc_140 N_S_c_78_n N_Y_c_412_n 0.00160128f $X=2.625 $Y=1.23 $X2=0 $Y2=0
cc_141 N_S_c_91_n N_Y_c_412_n 0.0179246f $X=2.89 $Y=2.41 $X2=0 $Y2=0
cc_142 N_S_c_92_n N_Y_c_412_n 0.0137878f $X=2.465 $Y=2.41 $X2=0 $Y2=0
cc_143 S N_Y_c_412_n 0.0135722f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_144 N_S_c_76_n N_Y_c_408_n 0.0101527f $X=2.55 $Y=1.155 $X2=0 $Y2=0
cc_145 N_S_c_77_n N_Y_c_408_n 0.00293164f $X=2.81 $Y=1.23 $X2=0 $Y2=0
cc_146 N_S_c_78_n N_Y_c_408_n 0.00453783f $X=2.625 $Y=1.23 $X2=0 $Y2=0
cc_147 S N_Y_c_408_n 0.00516207f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_148 N_S_c_83_n N_Y_c_409_n 0.00716793f $X=2.645 $Y=1.975 $X2=0 $Y2=0
cc_149 N_S_c_77_n N_Y_c_409_n 0.00326106f $X=2.81 $Y=1.23 $X2=0 $Y2=0
cc_150 N_S_c_78_n N_Y_c_409_n 0.00531691f $X=2.625 $Y=1.23 $X2=0 $Y2=0
cc_151 S N_Y_c_409_n 0.0527964f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_152 N_S_c_80_n N_Y_c_409_n 0.00381671f $X=2.975 $Y=1.32 $X2=0 $Y2=0
cc_153 N_S_c_98_p N_Y_c_434_n 0.0123021f $X=1.42 $Y=2.895 $X2=0 $Y2=0
cc_154 N_S_c_89_n N_Y_c_434_n 0.0228671f $X=2.295 $Y=2.98 $X2=0 $Y2=0
cc_155 N_S_c_76_n Y 0.00535962f $X=2.55 $Y=1.155 $X2=0 $Y2=0
cc_156 N_S_c_141_p A_452_497# 0.00564067f $X=2.38 $Y=2.895 $X2=-0.19 $Y2=-0.245
cc_157 N_S_c_91_n A_452_497# 9.40906e-19 $X=2.89 $Y=2.41 $X2=-0.19 $Y2=-0.245
cc_158 N_S_M1004_g N_VGND_c_475_n 0.00523461f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_159 N_S_c_76_n N_VGND_c_476_n 0.0101236f $X=2.55 $Y=1.155 $X2=0 $Y2=0
cc_160 N_S_c_77_n N_VGND_c_476_n 0.00778126f $X=2.81 $Y=1.23 $X2=0 $Y2=0
cc_161 S N_VGND_c_476_n 0.00232903f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_162 N_S_M1004_g N_VGND_c_477_n 0.00415323f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_163 N_S_c_76_n N_VGND_c_479_n 0.00345209f $X=2.55 $Y=1.155 $X2=0 $Y2=0
cc_164 N_S_M1004_g N_VGND_c_481_n 0.00469432f $X=0.635 $Y=0.835 $X2=0 $Y2=0
cc_165 N_S_c_76_n N_VGND_c_481_n 0.00394323f $X=2.55 $Y=1.155 $X2=0 $Y2=0
cc_166 N_A_55_125#_M1006_g N_A1_M1001_g 0.0313464f $X=1.205 $Y=2.695 $X2=0 $Y2=0
cc_167 N_A_55_125#_c_189_n A1 0.00920247f $X=1.085 $Y=1.59 $X2=0 $Y2=0
cc_168 N_A_55_125#_c_193_n A1 0.00920247f $X=1.19 $Y=1.995 $X2=0 $Y2=0
cc_169 N_A_55_125#_c_194_n A1 0.00169877f $X=1.19 $Y=2.145 $X2=0 $Y2=0
cc_170 N_A_55_125#_c_188_n A1 0.0262435f $X=1.085 $Y=1.59 $X2=0 $Y2=0
cc_171 N_A_55_125#_c_193_n N_A1_c_259_n 0.0108499f $X=1.19 $Y=1.995 $X2=0 $Y2=0
cc_172 N_A_55_125#_c_194_n N_A1_c_259_n 0.0313464f $X=1.19 $Y=2.145 $X2=0 $Y2=0
cc_173 N_A_55_125#_M1008_g N_A1_c_256_n 0.00920247f $X=1.175 $Y=0.835 $X2=0
+ $Y2=0
cc_174 N_A_55_125#_M1008_g N_A0_M1007_g 0.0299408f $X=1.175 $Y=0.835 $X2=0 $Y2=0
cc_175 N_A_55_125#_c_189_n N_A0_c_321_n 0.0325611f $X=1.085 $Y=1.59 $X2=0 $Y2=0
cc_176 N_A_55_125#_M1006_g N_VPWR_c_371_n 0.00631778f $X=1.205 $Y=2.695 $X2=0
+ $Y2=0
cc_177 N_A_55_125#_c_198_n N_VPWR_c_374_n 0.005097f $X=0.34 $Y=2.755 $X2=0 $Y2=0
cc_178 N_A_55_125#_c_199_n N_VPWR_c_374_n 0.00745538f $X=0.48 $Y=2.755 $X2=0
+ $Y2=0
cc_179 N_A_55_125#_M1006_g N_VPWR_c_376_n 0.00447026f $X=1.205 $Y=2.695 $X2=0
+ $Y2=0
cc_180 N_A_55_125#_M1006_g N_VPWR_c_370_n 0.00443817f $X=1.205 $Y=2.695 $X2=0
+ $Y2=0
cc_181 N_A_55_125#_c_198_n N_VPWR_c_370_n 0.00580745f $X=0.34 $Y=2.755 $X2=0
+ $Y2=0
cc_182 N_A_55_125#_c_199_n N_VPWR_c_370_n 0.00992023f $X=0.48 $Y=2.755 $X2=0
+ $Y2=0
cc_183 N_A_55_125#_M1008_g N_VGND_c_475_n 0.00146868f $X=1.175 $Y=0.835 $X2=0
+ $Y2=0
cc_184 N_A_55_125#_c_188_n N_VGND_c_475_n 0.0105778f $X=1.085 $Y=1.59 $X2=0
+ $Y2=0
cc_185 N_A_55_125#_c_189_n N_VGND_c_475_n 0.00264012f $X=1.085 $Y=1.59 $X2=0
+ $Y2=0
cc_186 N_A_55_125#_M1008_g N_VGND_c_479_n 0.00415323f $X=1.175 $Y=0.835 $X2=0
+ $Y2=0
cc_187 N_A_55_125#_M1008_g N_VGND_c_481_n 0.00469432f $X=1.175 $Y=0.835 $X2=0
+ $Y2=0
cc_188 N_A_55_125#_c_190_n N_VGND_c_481_n 0.0144247f $X=0.4 $Y=0.9 $X2=0 $Y2=0
cc_189 N_A1_c_251_n N_A0_M1007_g 0.00395799f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_190 N_A1_c_252_n N_A0_M1007_g 0.00128806f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_191 A1 N_A0_M1007_g 0.00994403f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A1_c_255_n N_A0_M1007_g 0.0105588f $X=1.985 $Y=0.515 $X2=0 $Y2=0
cc_193 N_A1_c_256_n N_A0_M1007_g 0.016746f $X=1.56 $Y=1.21 $X2=0 $Y2=0
cc_194 A1 N_A0_c_320_n 0.00227303f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_195 A1 N_A0_c_320_n 0.00961882f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A1_c_255_n N_A0_c_320_n 0.00911688f $X=1.985 $Y=0.515 $X2=0 $Y2=0
cc_197 A1 N_A0_c_321_n 0.00243408f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_198 A1 N_A0_c_321_n 0.00519819f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_199 N_A1_c_259_n N_A0_c_321_n 0.0217071f $X=1.655 $Y=1.94 $X2=0 $Y2=0
cc_200 A1 N_A0_c_322_n 0.00534063f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_201 N_A1_c_259_n N_A0_c_322_n 0.00668953f $X=1.655 $Y=1.94 $X2=0 $Y2=0
cc_202 N_A1_M1001_g N_A0_M1002_g 0.0188993f $X=1.565 $Y=2.695 $X2=0 $Y2=0
cc_203 A1 N_A0_M1002_g 7.11441e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_204 N_A1_c_259_n N_A0_M1002_g 0.00990077f $X=1.655 $Y=1.94 $X2=0 $Y2=0
cc_205 A1 A0 0.0123593f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_206 N_A1_M1001_g N_VPWR_c_371_n 3.00552e-19 $X=1.565 $Y=2.695 $X2=0 $Y2=0
cc_207 N_A1_M1001_g N_VPWR_c_376_n 8.9499e-19 $X=1.565 $Y=2.695 $X2=0 $Y2=0
cc_208 N_A1_M1001_g N_Y_c_411_n 0.0047523f $X=1.565 $Y=2.695 $X2=0 $Y2=0
cc_209 N_A1_M1001_g N_Y_c_413_n 6.76209e-19 $X=1.565 $Y=2.695 $X2=0 $Y2=0
cc_210 A1 N_Y_c_413_n 0.0119527f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_211 N_A1_c_259_n N_Y_c_413_n 0.00104448f $X=1.655 $Y=1.94 $X2=0 $Y2=0
cc_212 N_A1_M1001_g N_Y_c_434_n 0.00192484f $X=1.565 $Y=2.695 $X2=0 $Y2=0
cc_213 A1 N_Y_c_434_n 0.00243387f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_214 N_A1_c_259_n N_Y_c_434_n 0.00194409f $X=1.655 $Y=1.94 $X2=0 $Y2=0
cc_215 N_A1_c_251_n Y 0.0183264f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_216 N_A1_c_252_n Y 0.00383445f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_217 A1 Y 0.00571834f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_218 N_A1_c_255_n Y 0.0186557f $X=1.985 $Y=0.515 $X2=0 $Y2=0
cc_219 N_A1_c_256_n Y 0.0283728f $X=1.56 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A1_c_250_n N_VGND_c_475_n 0.0106161f $X=1.525 $Y=0.35 $X2=0 $Y2=0
cc_221 N_A1_c_256_n N_VGND_c_475_n 0.0168669f $X=1.56 $Y=1.21 $X2=0 $Y2=0
cc_222 N_A1_c_251_n N_VGND_c_476_n 0.00677895f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_223 N_A1_c_252_n N_VGND_c_476_n 0.00469138f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_224 N_A1_c_255_n N_VGND_c_476_n 0.00100666f $X=1.985 $Y=0.515 $X2=0 $Y2=0
cc_225 N_A1_c_250_n N_VGND_c_479_n 0.0114622f $X=1.525 $Y=0.35 $X2=0 $Y2=0
cc_226 N_A1_c_251_n N_VGND_c_479_n 0.0369241f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_227 N_A1_c_252_n N_VGND_c_479_n 0.00651318f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_228 N_A1_c_250_n N_VGND_c_481_n 0.00657784f $X=1.525 $Y=0.35 $X2=0 $Y2=0
cc_229 N_A1_c_251_n N_VGND_c_481_n 0.0218433f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_230 N_A1_c_252_n N_VGND_c_481_n 0.0100587f $X=1.985 $Y=0.35 $X2=0 $Y2=0
cc_231 N_A1_c_256_n A_250_125# 0.00440902f $X=1.56 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_232 N_A0_M1002_g N_VPWR_c_376_n 8.76173e-19 $X=2.185 $Y=2.695 $X2=0 $Y2=0
cc_233 N_A0_M1002_g N_Y_c_411_n 0.00900562f $X=2.185 $Y=2.695 $X2=0 $Y2=0
cc_234 N_A0_c_322_n N_Y_c_412_n 0.00246373f $X=2.185 $Y=1.875 $X2=0 $Y2=0
cc_235 N_A0_M1002_g N_Y_c_412_n 0.0128022f $X=2.185 $Y=2.695 $X2=0 $Y2=0
cc_236 A0 N_Y_c_412_n 0.0165118f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_237 N_A0_c_320_n N_Y_c_413_n 0.00260364f $X=2.03 $Y=1.49 $X2=0 $Y2=0
cc_238 N_A0_c_322_n N_Y_c_413_n 0.00218375f $X=2.185 $Y=1.875 $X2=0 $Y2=0
cc_239 N_A0_M1002_g N_Y_c_413_n 0.00157994f $X=2.185 $Y=2.695 $X2=0 $Y2=0
cc_240 A0 N_Y_c_413_n 0.00648476f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_241 N_A0_c_322_n N_Y_c_408_n 0.0024123f $X=2.185 $Y=1.875 $X2=0 $Y2=0
cc_242 A0 N_Y_c_408_n 0.0048087f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_243 N_A0_c_322_n N_Y_c_409_n 0.00827594f $X=2.185 $Y=1.875 $X2=0 $Y2=0
cc_244 N_A0_M1002_g N_Y_c_409_n 0.00181979f $X=2.185 $Y=2.695 $X2=0 $Y2=0
cc_245 A0 N_Y_c_409_n 0.0154775f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A0_M1002_g N_Y_c_434_n 0.00469903f $X=2.185 $Y=2.695 $X2=0 $Y2=0
cc_247 N_A0_M1007_g Y 0.0010211f $X=1.535 $Y=0.835 $X2=0 $Y2=0
cc_248 N_A0_c_320_n Y 0.00488662f $X=2.03 $Y=1.49 $X2=0 $Y2=0
cc_249 N_A0_c_322_n Y 0.00444733f $X=2.185 $Y=1.875 $X2=0 $Y2=0
cc_250 A0 Y 0.00903112f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_251 N_A0_M1007_g N_VGND_c_479_n 3.33984e-19 $X=1.535 $Y=0.835 $X2=0 $Y2=0
cc_252 N_Y_c_408_n N_VGND_c_476_n 0.00693121f $X=2.54 $Y=1.14 $X2=0 $Y2=0
cc_253 Y N_VGND_c_476_n 0.00733374f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_254 Y N_VGND_c_479_n 0.00155229f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_255 Y N_VGND_c_481_n 0.00292789f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_256 Y A_416_125# 0.00605058f $X=2.075 $Y=0.84 $X2=-0.19 $Y2=-0.245
