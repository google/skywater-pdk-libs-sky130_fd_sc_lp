* File: sky130_fd_sc_lp__o211a_lp.spice
* Created: Wed Sep  2 10:14:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o211a_lp.pex.spice"
.subckt sky130_fd_sc_lp__o211a_lp  VNB VPB A1 A2 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A1_M1010_g N_A_27_144#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.1197 PD=0.86 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_27_144#_M1002_d N_A2_M1002_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0924 PD=0.7 PS=0.86 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_318_144# N_B1_M1008_g N_A_27_144#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_232_419#_M1006_d N_C1_M1006_g A_318_144# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_606_47# N_A_232_419#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_232_419#_M1001_g A_606_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_134_419# N_A1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1003 N_A_232_419#_M1003_d N_A2_M1003_g A_134_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_A_232_419#_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.195 AS=0.14 PD=1.39 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1005 N_A_232_419#_M1005_d N_C1_M1005_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.195 PD=2.57 PS=1.39 NRD=0 NRS=21.67 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1004 N_X_M1004_d N_A_232_419#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX11_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o211a_lp.pxi.spice"
*
.ends
*
*
