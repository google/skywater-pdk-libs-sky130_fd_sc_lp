* File: sky130_fd_sc_lp__o31a_m.pxi.spice
* Created: Fri Aug 28 11:16:00 2020
* 
x_PM_SKY130_FD_SC_LP__O31A_M%A1 N_A1_M1000_g N_A1_M1008_g N_A1_c_71_n
+ N_A1_c_75_n A1 A1 N_A1_c_73_n PM_SKY130_FD_SC_LP__O31A_M%A1
x_PM_SKY130_FD_SC_LP__O31A_M%A_95_153# N_A_95_153#_M1005_d N_A_95_153#_M1009_d
+ N_A_95_153#_c_108_n N_A_95_153#_M1003_g N_A_95_153#_c_110_n
+ N_A_95_153#_M1006_g N_A_95_153#_c_115_n N_A_95_153#_c_116_n
+ N_A_95_153#_c_111_n N_A_95_153#_c_112_n N_A_95_153#_c_117_n
+ N_A_95_153#_c_118_n N_A_95_153#_c_119_n N_A_95_153#_c_120_n
+ N_A_95_153#_c_113_n N_A_95_153#_c_122_n N_A_95_153#_c_123_n
+ PM_SKY130_FD_SC_LP__O31A_M%A_95_153#
x_PM_SKY130_FD_SC_LP__O31A_M%A2 N_A2_M1004_g N_A2_M1001_g N_A2_c_184_n
+ N_A2_c_188_n A2 A2 A2 A2 N_A2_c_186_n PM_SKY130_FD_SC_LP__O31A_M%A2
x_PM_SKY130_FD_SC_LP__O31A_M%A3 N_A3_M1009_g N_A3_M1007_g N_A3_c_228_n
+ N_A3_c_229_n A3 N_A3_c_231_n PM_SKY130_FD_SC_LP__O31A_M%A3
x_PM_SKY130_FD_SC_LP__O31A_M%B1 N_B1_M1005_g N_B1_M1002_g N_B1_c_267_n
+ N_B1_c_268_n N_B1_c_269_n B1 B1 B1 N_B1_c_271_n PM_SKY130_FD_SC_LP__O31A_M%B1
x_PM_SKY130_FD_SC_LP__O31A_M%X N_X_M1006_s N_X_M1003_s N_X_c_303_n X X
+ PM_SKY130_FD_SC_LP__O31A_M%X
x_PM_SKY130_FD_SC_LP__O31A_M%VPWR N_VPWR_M1003_d N_VPWR_M1002_d N_VPWR_c_326_n
+ N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n VPWR N_VPWR_c_330_n
+ N_VPWR_c_331_n N_VPWR_c_325_n N_VPWR_c_333_n PM_SKY130_FD_SC_LP__O31A_M%VPWR
x_PM_SKY130_FD_SC_LP__O31A_M%VGND N_VGND_M1006_d N_VGND_M1001_d N_VGND_c_358_n
+ N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n VGND
+ N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n PM_SKY130_FD_SC_LP__O31A_M%VGND
x_PM_SKY130_FD_SC_LP__O31A_M%A_239_47# N_A_239_47#_M1000_d N_A_239_47#_M1007_d
+ N_A_239_47#_c_412_n N_A_239_47#_c_407_n N_A_239_47#_c_408_n
+ N_A_239_47#_c_411_n PM_SKY130_FD_SC_LP__O31A_M%A_239_47#
cc_1 VNB N_A1_M1000_g 0.0386706f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.445
cc_2 VNB N_A1_c_71_n 0.0206545f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.66
cc_3 VNB A1 0.00770822f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_4 VNB N_A1_c_73_n 0.0158945f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.32
cc_5 VNB N_A_95_153#_c_108_n 0.0104998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_95_153#_M1003_g 0.0303582f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.825
cc_7 VNB N_A_95_153#_c_110_n 0.019492f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_8 VNB N_A_95_153#_c_111_n 0.0221915f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.295
cc_9 VNB N_A_95_153#_c_112_n 0.00724238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_95_153#_c_113_n 0.0488037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_M1001_g 0.0373102f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.195
cc_12 VNB N_A2_c_184_n 0.0206235f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.66
cc_13 VNB A2 0.00530206f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_14 VNB N_A2_c_186_n 0.0153576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_M1009_g 0.00270614f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.445
cc_16 VNB N_A3_M1007_g 0.0261518f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.195
cc_17 VNB N_A3_c_228_n 0.0189297f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.66
cc_18 VNB N_A3_c_229_n 0.0159579f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.825
cc_19 VNB A3 0.00783899f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_20 VNB N_A3_c_231_n 0.0154759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_M1002_g 0.0126482f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.195
cc_22 VNB N_B1_c_267_n 0.0207147f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.32
cc_23 VNB N_B1_c_268_n 0.0252921f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.155
cc_24 VNB N_B1_c_269_n 0.0176217f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.66
cc_25 VNB B1 0.00230619f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.825
cc_26 VNB N_B1_c_271_n 0.018997f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.32
cc_27 VNB N_X_c_303_n 8.39306e-19 $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.32
cc_28 VNB X 0.0130763f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.66
cc_29 VNB X 0.0337823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_325_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_358_n 0.00435083f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.32
cc_32 VNB N_VGND_c_359_n 0.0158981f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.66
cc_33 VNB N_VGND_c_360_n 0.00286637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_361_n 0.0250674f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.32
cc_35 VNB N_VGND_c_362_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.32
cc_36 VNB N_VGND_c_363_n 0.0419555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_364_n 0.198733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_365_n 0.00522083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_239_47#_c_407_n 0.018487f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.66
cc_40 VNB N_A_239_47#_c_408_n 0.00784206f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.825
cc_41 VPB N_A1_M1008_g 0.0186082f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.195
cc_42 VPB N_A1_c_75_n 0.0152753f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.825
cc_43 VPB A1 0.00802994f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_44 VPB N_A_95_153#_M1003_g 0.0524629f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.825
cc_45 VPB N_A_95_153#_c_115_n 0.0371078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_95_153#_c_116_n 0.0150294f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.32
cc_47 VPB N_A_95_153#_c_117_n 0.0267425f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.32
cc_48 VPB N_A_95_153#_c_118_n 0.0103818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_95_153#_c_119_n 0.033368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_95_153#_c_120_n 0.00612432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_95_153#_c_113_n 0.00780757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_95_153#_c_122_n 0.0101849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_95_153#_c_123_n 0.0501092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A2_M1004_g 0.017802f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=0.445
cc_55 VPB N_A2_c_188_n 0.0153258f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.825
cc_56 VPB A2 0.00563486f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_57 VPB N_A3_M1009_g 0.0309155f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=0.445
cc_58 VPB N_B1_M1002_g 0.0354637f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.195
cc_59 VPB X 0.0285561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_326_n 0.0238704f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.32
cc_61 VPB N_VPWR_c_327_n 0.059817f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_62 VPB N_VPWR_c_328_n 0.026328f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_329_n 0.00401341f $X=-0.19 $Y=1.655 $X2=1.03 $Y2=1.32
cc_64 VPB N_VPWR_c_330_n 0.0442063f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.665
cc_65 VPB N_VPWR_c_331_n 0.0155085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_325_n 0.0979274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_333_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 N_A1_M1000_g N_A_95_153#_c_108_n 0.00777798f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_69 N_A1_M1008_g N_A_95_153#_M1003_g 0.0144032f $X=1.12 $Y=2.195 $X2=0 $Y2=0
cc_70 A1 N_A_95_153#_M1003_g 0.00189429f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A1_c_73_n N_A_95_153#_M1003_g 0.039541f $X=1.03 $Y=1.32 $X2=0 $Y2=0
cc_72 N_A1_M1000_g N_A_95_153#_c_110_n 0.0213828f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_73 N_A1_M1008_g N_A_95_153#_c_115_n 0.00928116f $X=1.12 $Y=2.195 $X2=0 $Y2=0
cc_74 N_A1_M1008_g N_A_95_153#_c_122_n 0.00113739f $X=1.12 $Y=2.195 $X2=0 $Y2=0
cc_75 N_A1_M1008_g N_A2_M1004_g 0.0208031f $X=1.12 $Y=2.195 $X2=0 $Y2=0
cc_76 N_A1_M1000_g N_A2_M1001_g 0.0332774f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A1_c_71_n N_A2_c_184_n 0.0208031f $X=1.03 $Y=1.66 $X2=0 $Y2=0
cc_78 N_A1_c_75_n N_A2_c_188_n 0.0208031f $X=1.03 $Y=1.825 $X2=0 $Y2=0
cc_79 N_A1_M1008_g A2 0.00271493f $X=1.12 $Y=2.195 $X2=0 $Y2=0
cc_80 A1 A2 0.0464404f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A1_c_73_n A2 6.2776e-19 $X=1.03 $Y=1.32 $X2=0 $Y2=0
cc_82 A1 N_A2_c_186_n 0.00448675f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A1_c_73_n N_A2_c_186_n 0.0208031f $X=1.03 $Y=1.32 $X2=0 $Y2=0
cc_84 N_A1_M1000_g X 0.00173874f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A1_M1008_g X 0.00131362f $X=1.12 $Y=2.195 $X2=0 $Y2=0
cc_86 A1 X 0.0277547f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A1_c_73_n X 0.00218263f $X=1.03 $Y=1.32 $X2=0 $Y2=0
cc_88 N_A1_M1008_g N_VPWR_c_326_n 0.00448819f $X=1.12 $Y=2.195 $X2=0 $Y2=0
cc_89 N_A1_c_75_n N_VPWR_c_326_n 0.00366294f $X=1.03 $Y=1.825 $X2=0 $Y2=0
cc_90 A1 N_VPWR_c_326_n 0.00140381f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A1_M1000_g N_VGND_c_358_n 0.00151442f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_92 A1 N_VGND_c_358_n 0.00163238f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A1_c_73_n N_VGND_c_358_n 0.00272142f $X=1.03 $Y=1.32 $X2=0 $Y2=0
cc_94 N_A1_M1000_g N_VGND_c_359_n 0.00585385f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A1_M1000_g N_VGND_c_360_n 7.33522e-19 $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A1_M1000_g N_VGND_c_364_n 0.0107511f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A1_M1000_g N_A_239_47#_c_408_n 0.00287294f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_98 A1 N_A_239_47#_c_408_n 0.0031716f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A_95_153#_c_117_n N_A2_M1004_g 0.00216092f $X=2.13 $Y=2.755 $X2=0 $Y2=0
cc_100 N_A_95_153#_c_122_n N_A2_M1004_g 0.00191288f $X=1.315 $Y=2.755 $X2=0
+ $Y2=0
cc_101 N_A_95_153#_c_123_n N_A2_M1004_g 0.00417602f $X=1.315 $Y=2.85 $X2=0 $Y2=0
cc_102 N_A_95_153#_c_117_n A2 0.0215268f $X=2.13 $Y=2.755 $X2=0 $Y2=0
cc_103 N_A_95_153#_c_118_n A2 0.013731f $X=2.235 $Y=2.26 $X2=0 $Y2=0
cc_104 N_A_95_153#_c_120_n A2 0.0087114f $X=2.34 $Y=1.89 $X2=0 $Y2=0
cc_105 N_A_95_153#_c_117_n N_A3_M1009_g 0.0064666f $X=2.13 $Y=2.755 $X2=0 $Y2=0
cc_106 N_A_95_153#_c_118_n N_A3_M1009_g 0.00278082f $X=2.235 $Y=2.26 $X2=0 $Y2=0
cc_107 N_A_95_153#_c_120_n N_A3_M1009_g 0.00233939f $X=2.34 $Y=1.89 $X2=0 $Y2=0
cc_108 N_A_95_153#_c_120_n N_A3_c_229_n 0.00400544f $X=2.34 $Y=1.89 $X2=0 $Y2=0
cc_109 N_A_95_153#_c_120_n A3 0.00868331f $X=2.34 $Y=1.89 $X2=0 $Y2=0
cc_110 N_A_95_153#_c_113_n A3 0.00243559f $X=3 $Y=0.51 $X2=0 $Y2=0
cc_111 N_A_95_153#_c_118_n N_B1_M1002_g 0.0073705f $X=2.235 $Y=2.26 $X2=0 $Y2=0
cc_112 N_A_95_153#_c_119_n N_B1_M1002_g 0.0188309f $X=2.915 $Y=1.89 $X2=0 $Y2=0
cc_113 N_A_95_153#_c_113_n N_B1_M1002_g 0.0104852f $X=3 $Y=0.51 $X2=0 $Y2=0
cc_114 N_A_95_153#_c_113_n N_B1_c_267_n 0.00414168f $X=3 $Y=0.51 $X2=0 $Y2=0
cc_115 N_A_95_153#_c_119_n N_B1_c_269_n 0.00327698f $X=2.915 $Y=1.89 $X2=0 $Y2=0
cc_116 N_A_95_153#_M1005_d B1 0.00263467f $X=2.635 $Y=0.235 $X2=0 $Y2=0
cc_117 N_A_95_153#_c_119_n B1 0.00762042f $X=2.915 $Y=1.89 $X2=0 $Y2=0
cc_118 N_A_95_153#_c_113_n B1 0.0675409f $X=3 $Y=0.51 $X2=0 $Y2=0
cc_119 N_A_95_153#_c_113_n N_B1_c_271_n 0.0164112f $X=3 $Y=0.51 $X2=0 $Y2=0
cc_120 N_A_95_153#_c_110_n N_X_c_303_n 0.00329851f $X=0.69 $Y=0.765 $X2=0 $Y2=0
cc_121 N_A_95_153#_c_111_n X 0.00817335f $X=0.69 $Y=0.84 $X2=0 $Y2=0
cc_122 N_A_95_153#_c_108_n X 0.00701822f $X=0.565 $Y=1.065 $X2=0 $Y2=0
cc_123 N_A_95_153#_M1003_g X 0.0412851f $X=0.58 $Y=2.195 $X2=0 $Y2=0
cc_124 N_A_95_153#_c_111_n X 0.0012965f $X=0.69 $Y=0.84 $X2=0 $Y2=0
cc_125 N_A_95_153#_c_112_n X 0.00500952f $X=0.565 $Y=1.155 $X2=0 $Y2=0
cc_126 N_A_95_153#_M1003_g N_VPWR_c_326_n 0.0175001f $X=0.58 $Y=2.195 $X2=0
+ $Y2=0
cc_127 N_A_95_153#_c_115_n N_VPWR_c_326_n 0.0207528f $X=1.15 $Y=2.85 $X2=0 $Y2=0
cc_128 N_A_95_153#_c_122_n N_VPWR_c_326_n 0.0258293f $X=1.315 $Y=2.755 $X2=0
+ $Y2=0
cc_129 N_A_95_153#_c_123_n N_VPWR_c_326_n 0.00508672f $X=1.315 $Y=2.85 $X2=0
+ $Y2=0
cc_130 N_A_95_153#_c_117_n N_VPWR_c_327_n 0.0108854f $X=2.13 $Y=2.755 $X2=0
+ $Y2=0
cc_131 N_A_95_153#_c_118_n N_VPWR_c_327_n 0.0280279f $X=2.235 $Y=2.26 $X2=0
+ $Y2=0
cc_132 N_A_95_153#_c_119_n N_VPWR_c_327_n 0.0235655f $X=2.915 $Y=1.89 $X2=0
+ $Y2=0
cc_133 N_A_95_153#_c_116_n N_VPWR_c_328_n 0.0072474f $X=0.655 $Y=2.85 $X2=0
+ $Y2=0
cc_134 N_A_95_153#_c_115_n N_VPWR_c_330_n 0.00445258f $X=1.15 $Y=2.85 $X2=0
+ $Y2=0
cc_135 N_A_95_153#_c_117_n N_VPWR_c_330_n 0.0226623f $X=2.13 $Y=2.755 $X2=0
+ $Y2=0
cc_136 N_A_95_153#_c_122_n N_VPWR_c_330_n 0.0160528f $X=1.315 $Y=2.755 $X2=0
+ $Y2=0
cc_137 N_A_95_153#_c_123_n N_VPWR_c_330_n 0.0059602f $X=1.315 $Y=2.85 $X2=0
+ $Y2=0
cc_138 N_A_95_153#_c_116_n N_VPWR_c_325_n 0.012474f $X=0.655 $Y=2.85 $X2=0 $Y2=0
cc_139 N_A_95_153#_c_117_n N_VPWR_c_325_n 0.02783f $X=2.13 $Y=2.755 $X2=0 $Y2=0
cc_140 N_A_95_153#_c_122_n N_VPWR_c_325_n 0.010655f $X=1.315 $Y=2.755 $X2=0
+ $Y2=0
cc_141 N_A_95_153#_c_123_n N_VPWR_c_325_n 0.00813556f $X=1.315 $Y=2.85 $X2=0
+ $Y2=0
cc_142 N_A_95_153#_c_110_n N_VGND_c_358_n 0.00288714f $X=0.69 $Y=0.765 $X2=0
+ $Y2=0
cc_143 N_A_95_153#_c_110_n N_VGND_c_361_n 0.00585385f $X=0.69 $Y=0.765 $X2=0
+ $Y2=0
cc_144 N_A_95_153#_c_111_n N_VGND_c_361_n 9.62948e-19 $X=0.69 $Y=0.84 $X2=0
+ $Y2=0
cc_145 N_A_95_153#_c_113_n N_VGND_c_363_n 0.00833313f $X=3 $Y=0.51 $X2=0 $Y2=0
cc_146 N_A_95_153#_M1005_d N_VGND_c_364_n 0.0094357f $X=2.635 $Y=0.235 $X2=0
+ $Y2=0
cc_147 N_A_95_153#_c_110_n N_VGND_c_364_n 0.0118894f $X=0.69 $Y=0.765 $X2=0
+ $Y2=0
cc_148 N_A_95_153#_c_111_n N_VGND_c_364_n 9.62037e-19 $X=0.69 $Y=0.84 $X2=0
+ $Y2=0
cc_149 N_A_95_153#_c_113_n N_VGND_c_364_n 0.00696426f $X=3 $Y=0.51 $X2=0 $Y2=0
cc_150 N_A_95_153#_c_113_n N_A_239_47#_c_411_n 0.00389536f $X=3 $Y=0.51 $X2=0
+ $Y2=0
cc_151 N_A2_M1004_g N_A3_M1009_g 0.0184434f $X=1.48 $Y=2.195 $X2=0 $Y2=0
cc_152 N_A2_c_188_n N_A3_M1009_g 0.0139728f $X=1.57 $Y=1.825 $X2=0 $Y2=0
cc_153 N_A2_M1001_g N_A3_M1007_g 0.020285f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_154 A2 N_A3_c_228_n 0.00119496f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_155 N_A2_c_186_n N_A3_c_228_n 0.0139728f $X=1.57 $Y=1.32 $X2=0 $Y2=0
cc_156 N_A2_c_184_n N_A3_c_229_n 0.0139728f $X=1.57 $Y=1.66 $X2=0 $Y2=0
cc_157 A2 N_A3_c_229_n 0.0123909f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A2_M1001_g A3 8.40661e-19 $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_159 A2 A3 0.027705f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A2_c_186_n A3 4.35554e-19 $X=1.57 $Y=1.32 $X2=0 $Y2=0
cc_161 N_A2_M1001_g N_A3_c_231_n 0.00873831f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_162 A2 N_VPWR_c_326_n 0.0124385f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_163 A2 A_311_397# 0.00556047f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_164 N_A2_M1001_g N_VGND_c_359_n 0.00414412f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A2_M1001_g N_VGND_c_360_n 0.00643429f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A2_M1001_g N_VGND_c_364_n 0.00486498f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A2_M1001_g N_A_239_47#_c_412_n 2.1266e-19 $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A2_M1001_g N_A_239_47#_c_407_n 0.0129476f $X=1.55 $Y=0.445 $X2=0 $Y2=0
cc_169 A2 N_A_239_47#_c_407_n 0.013408f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A2_c_186_n N_A_239_47#_c_407_n 0.00189471f $X=1.57 $Y=1.32 $X2=0 $Y2=0
cc_171 N_A2_c_186_n N_A_239_47#_c_408_n 0.00138418f $X=1.57 $Y=1.32 $X2=0 $Y2=0
cc_172 N_A3_M1009_g N_B1_M1002_g 0.0202538f $X=2.02 $Y=2.195 $X2=0 $Y2=0
cc_173 N_A3_c_229_n N_B1_M1002_g 0.0141865f $X=2.11 $Y=1.605 $X2=0 $Y2=0
cc_174 N_A3_M1007_g N_B1_c_267_n 0.018168f $X=2.075 $Y=0.445 $X2=0 $Y2=0
cc_175 A3 N_B1_c_268_n 0.0018924f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_176 N_A3_c_231_n N_B1_c_268_n 0.0141865f $X=2.11 $Y=1.1 $X2=0 $Y2=0
cc_177 N_A3_c_228_n N_B1_c_269_n 0.0141865f $X=2.11 $Y=1.44 $X2=0 $Y2=0
cc_178 N_A3_M1007_g B1 7.29443e-19 $X=2.075 $Y=0.445 $X2=0 $Y2=0
cc_179 A3 B1 0.0201847f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A3_c_231_n B1 9.73789e-19 $X=2.11 $Y=1.1 $X2=0 $Y2=0
cc_181 N_A3_M1007_g N_VGND_c_360_n 0.00443559f $X=2.075 $Y=0.445 $X2=0 $Y2=0
cc_182 N_A3_M1007_g N_VGND_c_363_n 0.00429465f $X=2.075 $Y=0.445 $X2=0 $Y2=0
cc_183 N_A3_M1007_g N_VGND_c_364_n 0.00638334f $X=2.075 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A3_M1007_g N_A_239_47#_c_407_n 0.0122335f $X=2.075 $Y=0.445 $X2=0 $Y2=0
cc_185 A3 N_A_239_47#_c_407_n 0.024567f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A3_c_231_n N_A_239_47#_c_407_n 0.00518598f $X=2.11 $Y=1.1 $X2=0 $Y2=0
cc_187 N_A3_M1007_g N_A_239_47#_c_411_n 2.16198e-19 $X=2.075 $Y=0.445 $X2=0
+ $Y2=0
cc_188 N_B1_M1002_g N_VPWR_c_327_n 0.00836635f $X=2.56 $Y=2.195 $X2=0 $Y2=0
cc_189 N_B1_M1002_g N_VPWR_c_325_n 0.00330899f $X=2.56 $Y=2.195 $X2=0 $Y2=0
cc_190 N_B1_c_267_n N_VGND_c_363_n 0.0048701f $X=2.65 $Y=0.765 $X2=0 $Y2=0
cc_191 B1 N_VGND_c_363_n 0.00426263f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_192 N_B1_c_271_n N_VGND_c_363_n 0.00185549f $X=2.65 $Y=0.93 $X2=0 $Y2=0
cc_193 N_B1_c_267_n N_VGND_c_364_n 0.00974176f $X=2.65 $Y=0.765 $X2=0 $Y2=0
cc_194 B1 N_VGND_c_364_n 0.00568396f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_195 N_B1_c_271_n N_VGND_c_364_n 0.00213938f $X=2.65 $Y=0.93 $X2=0 $Y2=0
cc_196 N_B1_c_267_n N_A_239_47#_c_407_n 0.00142304f $X=2.65 $Y=0.765 $X2=0 $Y2=0
cc_197 B1 N_A_239_47#_c_407_n 0.0131547f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_198 N_B1_c_267_n N_A_239_47#_c_411_n 0.00142799f $X=2.65 $Y=0.765 $X2=0 $Y2=0
cc_199 B1 N_A_239_47#_c_411_n 0.013246f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_200 X N_VPWR_c_326_n 0.010245f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_201 N_X_c_303_n N_VGND_c_361_n 0.00877924f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_202 X N_VGND_c_361_n 0.00399781f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_203 N_X_M1006_s N_VGND_c_364_n 0.00272007f $X=0.35 $Y=0.235 $X2=0 $Y2=0
cc_204 N_X_c_303_n N_VGND_c_364_n 0.00770513f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_205 X N_VGND_c_364_n 0.00630506f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_206 N_X_c_303_n N_A_239_47#_c_412_n 2.54064e-19 $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_207 N_X_c_303_n N_A_239_47#_c_408_n 0.00556613f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_208 N_VGND_c_364_n N_A_239_47#_M1000_d 0.00369956f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_209 N_VGND_c_364_n N_A_239_47#_M1007_d 0.00674488f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_359_n N_A_239_47#_c_412_n 0.0081737f $X=1.62 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_364_n N_A_239_47#_c_412_n 0.00762225f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_212 N_VGND_c_359_n N_A_239_47#_c_407_n 0.002793f $X=1.62 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_c_360_n N_A_239_47#_c_407_n 0.02169f $X=1.785 $Y=0.38 $X2=0 $Y2=0
cc_214 N_VGND_c_363_n N_A_239_47#_c_407_n 0.00372557f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_c_364_n N_A_239_47#_c_407_n 0.0115499f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_363_n N_A_239_47#_c_411_n 0.0077266f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_364_n N_A_239_47#_c_411_n 0.00688934f $X=3.12 $Y=0 $X2=0 $Y2=0
