* File: sky130_fd_sc_lp__and4_lp.pex.spice
* Created: Wed Sep  2 09:33:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4_LP%D 3 5 6 9 13 20 22 23 24 35
c42 22 0 8.05769e-20 $X=0.72 $Y=1.295
c43 20 0 1.80104e-19 $X=0.855 $Y=1.835
r44 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.405 $X2=0.585 $Y2=1.405
r45 23 24 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=2.035
r46 23 36 4.38001 $w=7.08e-07 $l=2.6e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=1.405
r47 22 36 1.85308 $w=7.08e-07 $l=1.1e-07 $layer=LI1_cond $X=0.48 $Y=1.295
+ $X2=0.48 $Y2=1.405
r48 19 35 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.585 $Y=1.76
+ $X2=0.585 $Y2=1.405
r49 19 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.585 $Y=1.835
+ $X2=0.855 $Y2=1.835
r50 16 19 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.495 $Y=1.835
+ $X2=0.585 $Y2=1.835
r51 15 35 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.585 $Y=1.39
+ $X2=0.585 $Y2=1.405
r52 11 13 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.075 $Y=1.24
+ $X2=1.075 $Y2=0.485
r53 7 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.855 $Y=1.91
+ $X2=0.855 $Y2=1.835
r54 7 9 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=0.855 $Y=1.91
+ $X2=0.855 $Y2=2.635
r55 6 15 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.75 $Y=1.315
+ $X2=0.585 $Y2=1.39
r56 5 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1 $Y=1.315
+ $X2=1.075 $Y2=1.24
r57 5 6 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1 $Y=1.315 $X2=0.75
+ $Y2=1.315
r58 1 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.91
+ $X2=0.495 $Y2=1.835
r59 1 3 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=0.495 $Y=1.91
+ $X2=0.495 $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP%C 3 7 11 16 17 21 22 23 24 38
c54 38 0 8.05769e-20 $X=1.555 $Y=1.275
c55 21 0 1.80104e-19 $X=1.68 $Y=0.555
c56 17 0 1.87633e-19 $X=1.645 $Y=1.705
r57 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.555
+ $Y=1.275 $X2=1.555 $Y2=1.275
r58 23 24 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.44 $Y=1.295
+ $X2=1.44 $Y2=1.665
r59 23 39 0.336923 $w=7.08e-07 $l=2e-08 $layer=LI1_cond $X=1.44 $Y=1.295
+ $X2=1.44 $Y2=1.275
r60 22 39 5.89616 $w=7.08e-07 $l=3.5e-07 $layer=LI1_cond $X=1.44 $Y=0.925
+ $X2=1.44 $Y2=1.275
r61 21 22 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.44 $Y=0.555
+ $X2=1.44 $Y2=0.925
r62 20 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.555 $Y=1.11
+ $X2=1.555 $Y2=1.275
r63 16 38 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.555 $Y=1.63
+ $X2=1.555 $Y2=1.275
r64 16 17 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.555 $Y=1.705
+ $X2=1.645 $Y2=1.705
r65 13 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.285 $Y=1.705
+ $X2=1.555 $Y2=1.705
r66 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.645 $Y=1.78
+ $X2=1.645 $Y2=1.705
r67 9 11 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.645 $Y=1.78
+ $X2=1.645 $Y2=2.635
r68 7 20 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.465 $Y=0.485
+ $X2=1.465 $Y2=1.11
r69 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.285 $Y=1.78
+ $X2=1.285 $Y2=1.705
r70 1 3 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.285 $Y=1.78
+ $X2=1.285 $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP%B 3 6 9 13 18 20 21 22 23 29
r55 29 31 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.127 $Y=1.36
+ $X2=2.127 $Y2=1.195
r56 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.13 $Y=1.295
+ $X2=2.13 $Y2=1.665
r57 22 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.13
+ $Y=1.36 $X2=2.13 $Y2=1.36
r58 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.13 $Y=0.925
+ $X2=2.13 $Y2=1.295
r59 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.13 $Y=0.555
+ $X2=2.13 $Y2=0.925
r60 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.435 $Y=1.865
+ $X2=2.435 $Y2=1.79
r61 11 13 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.435 $Y=1.865
+ $X2=2.435 $Y2=2.635
r62 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.075 $Y=1.865
+ $X2=2.075 $Y2=1.79
r63 7 9 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.075 $Y=1.865
+ $X2=2.075 $Y2=2.635
r64 6 18 157.932 $w=1.5e-07 $l=3.08e-07 $layer=POLY_cond $X=2.127 $Y=1.79
+ $X2=2.435 $Y2=1.79
r65 6 15 26.6638 $w=1.5e-07 $l=5.2e-08 $layer=POLY_cond $X=2.127 $Y=1.79
+ $X2=2.075 $Y2=1.79
r66 5 29 0.344503 $w=3.35e-07 $l=2e-09 $layer=POLY_cond $X=2.127 $Y=1.362
+ $X2=2.127 $Y2=1.36
r67 5 6 60.8048 $w=3.35e-07 $l=3.53e-07 $layer=POLY_cond $X=2.127 $Y=1.362
+ $X2=2.127 $Y2=1.715
r68 3 31 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.035 $Y=0.485
+ $X2=2.035 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP%A 1 3 4 5 9 10 12 13 15 17 19 20 21 22 23 24
+ 28
r72 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.955
+ $Y=1.39 $X2=2.955 $Y2=1.39
r73 24 29 2.94557 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=1.56
+ $X2=2.955 $Y2=1.56
r74 23 29 5.62335 $w=6.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.64 $Y=1.56
+ $X2=2.955 $Y2=1.56
r75 20 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.955 $Y=1.73
+ $X2=2.955 $Y2=1.39
r76 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.73
+ $X2=2.955 $Y2=1.895
r77 19 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.225
+ $X2=2.955 $Y2=1.39
r78 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.225 $Y=2.315
+ $X2=3.225 $Y2=2.635
r79 14 22 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.94 $Y=2.24
+ $X2=2.865 $Y2=2.24
r80 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.15 $Y=2.24
+ $X2=3.225 $Y2=2.315
r81 13 14 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.15 $Y=2.24
+ $X2=2.94 $Y2=2.24
r82 10 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=2.315
+ $X2=2.865 $Y2=2.24
r83 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.865 $Y=2.315
+ $X2=2.865 $Y2=2.635
r84 9 22 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=2.165
+ $X2=2.865 $Y2=2.24
r85 9 21 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.865 $Y=2.165
+ $X2=2.865 $Y2=1.895
r86 6 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.865 $Y=0.955
+ $X2=2.865 $Y2=1.225
r87 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.79 $Y=0.88
+ $X2=2.865 $Y2=0.955
r88 4 5 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.79 $Y=0.88 $X2=2.5
+ $Y2=0.88
r89 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.425 $Y=0.805
+ $X2=2.5 $Y2=0.88
r90 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.425 $Y=0.805
+ $X2=2.425 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP%A_186_485# 1 2 3 12 16 20 24 28 29 32 36 38
+ 39 40 42 43 45 47 48 50 53 54
c121 28 0 1.87633e-19 $X=2.485 $Y=2.15
r122 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.615
+ $Y=1.05 $X2=3.615 $Y2=1.05
r123 47 48 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.07 $Y=2.635
+ $X2=1.07 $Y2=2.405
r124 45 54 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.49 $Y=2.065
+ $X2=3.49 $Y2=1.555
r125 43 54 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=3.592 $Y=1.368
+ $X2=3.592 $Y2=1.555
r126 42 52 2.54787 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=3.592 $Y=1.055
+ $X2=3.592 $Y2=0.97
r127 42 43 9.61906 $w=3.73e-07 $l=3.13e-07 $layer=LI1_cond $X=3.592 $Y=1.055
+ $X2=3.592 $Y2=1.368
r128 41 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=2.15
+ $X2=2.65 $Y2=2.15
r129 40 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.405 $Y=2.15
+ $X2=3.49 $Y2=2.065
r130 40 41 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.405 $Y=2.15
+ $X2=2.815 $Y2=2.15
r131 38 52 5.60532 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=3.405 $Y=0.97
+ $X2=3.592 $Y2=0.97
r132 38 39 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.405 $Y=0.97
+ $X2=2.805 $Y2=0.97
r133 34 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=2.235
+ $X2=2.65 $Y2=2.15
r134 34 36 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.65 $Y=2.235 $X2=2.65
+ $Y2=2.635
r135 30 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.64 $Y=0.885
+ $X2=2.805 $Y2=0.97
r136 30 32 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.64 $Y=0.885 $X2=2.64
+ $Y2=0.485
r137 28 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.485 $Y=2.15
+ $X2=2.65 $Y2=2.15
r138 28 29 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.485 $Y=2.15
+ $X2=1.235 $Y2=2.15
r139 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.235
+ $X2=1.235 $Y2=2.15
r140 26 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.15 $Y=2.235
+ $X2=1.15 $Y2=2.405
r141 22 53 76.1577 $w=3.35e-07 $l=6.2155e-07 $layer=POLY_cond $X=4.045 $Y=1.555
+ $X2=3.785 $Y2=1.05
r142 22 24 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=4.045 $Y=1.555
+ $X2=4.045 $Y2=2.635
r143 18 53 27.2383 $w=3.35e-07 $l=2.20624e-07 $layer=POLY_cond $X=3.915 $Y=0.885
+ $X2=3.785 $Y2=1.05
r144 18 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.915 $Y=0.885
+ $X2=3.915 $Y2=0.485
r145 14 53 76.1577 $w=3.35e-07 $l=5.66282e-07 $layer=POLY_cond $X=3.655 $Y=1.555
+ $X2=3.785 $Y2=1.05
r146 14 16 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=3.655 $Y=1.555
+ $X2=3.655 $Y2=2.635
r147 10 53 27.2383 $w=3.35e-07 $l=2.6e-07 $layer=POLY_cond $X=3.525 $Y=1.05
+ $X2=3.785 $Y2=1.05
r148 10 12 205.106 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.525 $Y=1.05
+ $X2=3.525 $Y2=0.485
r149 3 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.51
+ $Y=2.425 $X2=2.65 $Y2=2.635
r150 2 47 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=2.425 $X2=1.07 $Y2=2.635
r151 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.275 $X2=2.64 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP%VPWR 1 2 3 10 12 16 20 23 24 25 34 43 44 50
r55 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 44 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 41 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.44 $Y2=3.33
r60 41 43 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r62 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r64 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 34 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.44 $Y2=3.33
r66 34 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 33 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r68 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 30 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r72 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 27 47 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r74 27 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 25 40 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r76 25 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 23 32 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.68 $Y2=3.33
r78 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.86 $Y2=3.33
r79 22 36 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.16 $Y2=3.33
r80 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.86 $Y2=3.33
r81 18 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=3.33
r82 18 20 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=2.635
r83 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=3.245
+ $X2=1.86 $Y2=3.33
r84 14 16 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=1.86 $Y=3.245
+ $X2=1.86 $Y2=2.635
r85 10 47 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r86 10 12 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.635
r87 3 20 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=2.425 $X2=3.44 $Y2=2.635
r88 2 16 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.72
+ $Y=2.425 $X2=1.86 $Y2=2.635
r89 1 12 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.425 $X2=0.28 $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP%X 1 2 7 8 9 10 11 12 13 35
r20 13 52 2.35846 $w=7.08e-07 $l=1.4e-07 $layer=LI1_cond $X=4.32 $Y=2.775
+ $X2=4.32 $Y2=2.635
r21 12 52 3.87462 $w=7.08e-07 $l=2.3e-07 $layer=LI1_cond $X=4.32 $Y=2.405
+ $X2=4.32 $Y2=2.635
r22 11 12 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=4.32 $Y=2.035
+ $X2=4.32 $Y2=2.405
r23 10 11 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=4.32 $Y=1.665
+ $X2=4.32 $Y2=2.035
r24 9 10 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=4.32 $Y=1.295
+ $X2=4.32 $Y2=1.665
r25 8 9 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=4.32 $Y=0.925 $X2=4.32
+ $Y2=1.295
r26 8 35 2.19 $w=7.08e-07 $l=1.3e-07 $layer=LI1_cond $X=4.32 $Y=0.925 $X2=4.32
+ $Y2=0.795
r27 7 35 5.77805 $w=7.1e-07 $l=3.1e-07 $layer=LI1_cond $X=4.32 $Y=0.485 $X2=4.32
+ $Y2=0.795
r28 2 52 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=2.425 $X2=4.26 $Y2=2.635
r29 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.275 $X2=4.13 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP%VGND 1 2 9 13 16 17 18 20 36 37 40
r41 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r43 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r44 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r45 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r46 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r47 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r49 27 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r50 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 25 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r52 25 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.2
+ $Y2=0
r53 23 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 20 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r56 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r57 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r58 18 28 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r59 16 30 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.12
+ $Y2=0
r60 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.31
+ $Y2=0
r61 15 33 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.6
+ $Y2=0
r62 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.31
+ $Y2=0
r63 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=0.085
+ $X2=3.31 $Y2=0
r64 11 13 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.31 $Y=0.085 $X2=3.31
+ $Y2=0.485
r65 7 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0
r66 7 9 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0.485
r67 2 13 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.165
+ $Y=0.275 $X2=3.31 $Y2=0.485
r68 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.275 $X2=0.75 $Y2=0.485
.ends

