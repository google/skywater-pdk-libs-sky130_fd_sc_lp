* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or3_2 A B C VGND VNB VPB VPWR X
X0 a_132_367# B a_207_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_207_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND B a_35_60# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_35_60# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 X a_35_60# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_35_60# C a_132_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_35_60# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_35_60# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR a_35_60# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_35_60# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
