* File: sky130_fd_sc_lp__a2111o_lp.pxi.spice
* Created: Wed Sep  2 09:16:31 2020
* 
x_PM_SKY130_FD_SC_LP__A2111O_LP%D1 N_D1_M1001_g N_D1_M1000_g N_D1_c_106_n
+ N_D1_M1014_g N_D1_c_108_n N_D1_c_109_n D1 D1 N_D1_c_110_n N_D1_c_111_n
+ PM_SKY130_FD_SC_LP__A2111O_LP%D1
x_PM_SKY130_FD_SC_LP__A2111O_LP%C1 N_C1_M1006_g N_C1_c_151_n N_C1_M1007_g
+ N_C1_c_152_n N_C1_c_153_n N_C1_M1002_g N_C1_c_154_n C1 C1 N_C1_c_156_n
+ N_C1_c_157_n PM_SKY130_FD_SC_LP__A2111O_LP%C1
x_PM_SKY130_FD_SC_LP__A2111O_LP%A_27_409# N_A_27_409#_M1014_d
+ N_A_27_409#_M1009_s N_A_27_409#_M1005_d N_A_27_409#_M1000_s
+ N_A_27_409#_M1013_g N_A_27_409#_M1015_g N_A_27_409#_M1008_g
+ N_A_27_409#_c_222_n N_A_27_409#_c_223_n N_A_27_409#_c_224_n
+ N_A_27_409#_c_209_n N_A_27_409#_c_210_n N_A_27_409#_c_211_n
+ N_A_27_409#_c_212_n N_A_27_409#_c_213_n N_A_27_409#_c_214_n
+ N_A_27_409#_c_215_n N_A_27_409#_c_216_n N_A_27_409#_c_217_n
+ N_A_27_409#_c_218_n N_A_27_409#_c_219_n N_A_27_409#_c_220_n
+ PM_SKY130_FD_SC_LP__A2111O_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__A2111O_LP%B1 N_B1_c_343_n N_B1_M1009_g N_B1_M1011_g
+ N_B1_c_344_n N_B1_c_345_n N_B1_M1010_g N_B1_c_346_n N_B1_c_347_n N_B1_c_353_n
+ N_B1_c_348_n B1 B1 N_B1_c_350_n PM_SKY130_FD_SC_LP__A2111O_LP%B1
x_PM_SKY130_FD_SC_LP__A2111O_LP%A2 N_A2_c_403_n N_A2_M1003_g N_A2_M1004_g
+ N_A2_c_405_n A2 A2 N_A2_c_407_n PM_SKY130_FD_SC_LP__A2111O_LP%A2
x_PM_SKY130_FD_SC_LP__A2111O_LP%A1 N_A1_M1005_g N_A1_M1012_g N_A1_c_447_n
+ N_A1_c_452_n A1 A1 N_A1_c_449_n PM_SKY130_FD_SC_LP__A2111O_LP%A1
x_PM_SKY130_FD_SC_LP__A2111O_LP%A_232_409# N_A_232_409#_M1006_d
+ N_A_232_409#_M1011_s N_A_232_409#_c_480_n N_A_232_409#_c_481_n
+ N_A_232_409#_c_482_n N_A_232_409#_c_483_n N_A_232_409#_c_484_n
+ N_A_232_409#_c_487_n N_A_232_409#_c_503_n
+ PM_SKY130_FD_SC_LP__A2111O_LP%A_232_409#
x_PM_SKY130_FD_SC_LP__A2111O_LP%VPWR N_VPWR_M1015_s N_VPWR_M1003_d
+ N_VPWR_c_521_n N_VPWR_c_522_n N_VPWR_c_523_n N_VPWR_c_524_n VPWR
+ N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_520_n N_VPWR_c_528_n
+ PM_SKY130_FD_SC_LP__A2111O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A2111O_LP%X N_X_M1008_d N_X_M1015_d N_X_c_564_n
+ N_X_c_565_n N_X_c_579_n X PM_SKY130_FD_SC_LP__A2111O_LP%X
x_PM_SKY130_FD_SC_LP__A2111O_LP%A_739_409# N_A_739_409#_M1011_d
+ N_A_739_409#_M1012_d N_A_739_409#_c_593_n N_A_739_409#_c_594_n
+ N_A_739_409#_c_595_n N_A_739_409#_c_596_n N_A_739_409#_c_597_n
+ PM_SKY130_FD_SC_LP__A2111O_LP%A_739_409#
x_PM_SKY130_FD_SC_LP__A2111O_LP%VGND N_VGND_M1001_s N_VGND_M1002_d
+ N_VGND_M1010_d N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_630_n N_VGND_c_631_n
+ N_VGND_c_632_n N_VGND_c_633_n VGND N_VGND_c_634_n N_VGND_c_635_n
+ N_VGND_c_636_n N_VGND_c_637_n PM_SKY130_FD_SC_LP__A2111O_LP%VGND
cc_1 VNB N_D1_M1001_g 0.0219544f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_2 VNB N_D1_M1000_g 0.00938167f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_3 VNB N_D1_c_106_n 0.0206992f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.86
cc_4 VNB N_D1_M1014_g 0.0157113f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_5 VNB N_D1_c_108_n 0.0176301f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.86
cc_6 VNB N_D1_c_109_n 0.0230745f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.525
cc_7 VNB N_D1_c_110_n 0.0411494f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.02
cc_8 VNB N_D1_c_111_n 0.0312454f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.02
cc_9 VNB N_C1_c_151_n 0.0135266f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.525
cc_10 VNB N_C1_c_152_n 0.0190111f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.86
cc_11 VNB N_C1_c_153_n 0.013722f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_12 VNB N_C1_c_154_n 0.00437176f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.935
cc_13 VNB C1 0.00171029f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.86
cc_14 VNB N_C1_c_156_n 0.0528942f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_C1_c_157_n 0.0195346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_409#_M1013_g 0.0335128f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.935
cc_17 VNB N_A_27_409#_M1008_g 0.0222349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_409#_c_209_n 0.0013378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_409#_c_210_n 0.012121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_409#_c_211_n 0.0140079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_409#_c_212_n 0.00148114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_409#_c_213_n 0.00914236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_409#_c_214_n 0.00901275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_409#_c_215_n 0.0317179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_409#_c_216_n 0.0240181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_409#_c_217_n 0.00444224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_409#_c_218_n 0.0125242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_409#_c_219_n 0.0120361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_409#_c_220_n 0.146118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B1_c_343_n 0.0175029f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.785
cc_31 VNB N_B1_c_344_n 0.0167543f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.86
cc_32 VNB N_B1_c_345_n 0.0138901f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_33 VNB N_B1_c_346_n 0.0166377f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.86
cc_34 VNB N_B1_c_347_n 0.0267148f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_35 VNB N_B1_c_348_n 0.0057254f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.525
cc_36 VNB B1 0.00463468f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_37 VNB N_B1_c_350_n 0.0145555f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.02
cc_38 VNB N_A2_c_403_n 0.0207968f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_39 VNB N_A2_M1004_g 0.0358192f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.86
cc_40 VNB N_A2_c_405_n 9.4531e-19 $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.785
cc_41 VNB A2 0.00243157f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_42 VNB N_A2_c_407_n 0.0231439f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_43 VNB N_A1_M1005_g 0.0448828f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_44 VNB N_A1_c_447_n 0.023616f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.785
cc_45 VNB A1 0.0310519f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.935
cc_46 VNB N_A1_c_449_n 0.0170897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VPWR_c_520_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_X_c_564_n 0.00876658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_X_c_565_n 0.00378311f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_50 VNB N_VGND_c_628_n 0.0110036f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.86
cc_51 VNB N_VGND_c_629_n 0.0218419f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.445
cc_52 VNB N_VGND_c_630_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.86
cc_53 VNB N_VGND_c_631_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_54 VNB N_VGND_c_632_n 0.0334731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_633_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.02
cc_56 VNB N_VGND_c_634_n 0.0477599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_635_n 0.0322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_636_n 0.288583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_637_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VPB N_D1_M1000_g 0.0516533f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_61 VPB N_D1_c_111_n 0.00824848f $X=-0.19 $Y=1.655 $X2=0.365 $Y2=1.02
cc_62 VPB N_C1_M1006_g 0.0362158f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_63 VPB C1 0.00218802f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.86
cc_64 VPB N_C1_c_156_n 0.0254696f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_65 VPB N_A_27_409#_M1015_g 0.0366955f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.525
cc_66 VPB N_A_27_409#_c_222_n 0.0101883f $X=-0.19 $Y=1.655 $X2=0.365 $Y2=1.02
cc_67 VPB N_A_27_409#_c_223_n 0.0353271f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.02
cc_68 VPB N_A_27_409#_c_224_n 0.00148891f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.295
cc_69 VPB N_A_27_409#_c_210_n 0.00705308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_27_409#_c_212_n 0.00523215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_27_409#_c_220_n 0.028695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_B1_M1011_g 0.0351794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_B1_c_347_n 0.00234379f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.375
cc_74 VPB N_B1_c_353_n 0.0183683f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.375
cc_75 VPB B1 0.0022214f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_76 VPB N_A2_M1003_g 0.0290319f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.525
cc_77 VPB N_A2_c_405_n 0.0191764f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.785
cc_78 VPB A2 7.45984e-19 $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.445
cc_79 VPB N_A1_M1012_g 0.037865f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_80 VPB N_A1_c_447_n 0.00180504f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.785
cc_81 VPB N_A1_c_452_n 0.0144588f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.445
cc_82 VPB A1 0.0136064f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.935
cc_83 VPB N_A_232_409#_c_480_n 0.0101911f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.86
cc_84 VPB N_A_232_409#_c_481_n 0.00928687f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.445
cc_85 VPB N_A_232_409#_c_482_n 0.0437198f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.935
cc_86 VPB N_A_232_409#_c_483_n 0.0186711f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=1.525
cc_87 VPB N_A_232_409#_c_484_n 0.0226067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_521_n 0.0099948f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.86
cc_89 VPB N_VPWR_c_522_n 0.00417436f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.445
cc_90 VPB N_VPWR_c_523_n 0.0578323f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.86
cc_91 VPB N_VPWR_c_524_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.375
cc_92 VPB N_VPWR_c_525_n 0.0544846f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_93 VPB N_VPWR_c_526_n 0.0229838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_520_n 0.0883157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_528_n 0.00620906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_X_c_564_n 0.00906934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB X 0.00898414f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.935
cc_98 VPB N_A_739_409#_c_593_n 0.00946742f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_99 VPB N_A_739_409#_c_594_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.86
cc_100 VPB N_A_739_409#_c_595_n 0.00584497f $X=-0.19 $Y=1.655 $X2=0.885
+ $Y2=0.785
cc_101 VPB N_A_739_409#_c_596_n 0.00978367f $X=-0.19 $Y=1.655 $X2=0.885
+ $Y2=0.445
cc_102 VPB N_A_739_409#_c_597_n 0.0353271f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.935
cc_103 N_D1_M1000_g N_C1_M1006_g 0.0472883f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_104 N_D1_M1014_g N_C1_c_151_n 0.0105817f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_105 N_D1_c_106_n N_C1_c_154_n 0.0105817f $X=0.81 $Y=0.86 $X2=0 $Y2=0
cc_106 N_D1_c_106_n N_C1_c_156_n 0.00280779f $X=0.81 $Y=0.86 $X2=0 $Y2=0
cc_107 N_D1_c_109_n N_C1_c_156_n 0.0472883f $X=0.435 $Y=1.525 $X2=0 $Y2=0
cc_108 N_D1_c_110_n N_C1_c_156_n 0.00619905f $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_109 N_D1_c_110_n N_C1_c_157_n 0.00250361f $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_110 N_D1_M1000_g N_A_27_409#_c_222_n 0.0012099f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_111 N_D1_c_109_n N_A_27_409#_c_222_n 0.00100339f $X=0.435 $Y=1.525 $X2=0
+ $Y2=0
cc_112 N_D1_c_111_n N_A_27_409#_c_222_n 0.0228694f $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_113 N_D1_M1000_g N_A_27_409#_c_223_n 0.0176529f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_114 N_D1_M1000_g N_A_27_409#_c_224_n 0.0222274f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_115 N_D1_c_111_n N_A_27_409#_c_224_n 0.00474601f $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_116 N_D1_M1001_g N_A_27_409#_c_209_n 0.00606143f $X=0.495 $Y=0.445 $X2=0
+ $Y2=0
cc_117 N_D1_c_106_n N_A_27_409#_c_209_n 0.00344443f $X=0.81 $Y=0.86 $X2=0 $Y2=0
cc_118 N_D1_M1014_g N_A_27_409#_c_209_n 0.0129052f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_119 N_D1_c_109_n N_A_27_409#_c_210_n 0.00896031f $X=0.435 $Y=1.525 $X2=0
+ $Y2=0
cc_120 N_D1_c_110_n N_A_27_409#_c_210_n 0.00357569f $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_121 N_D1_c_111_n N_A_27_409#_c_210_n 0.0572896f $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_122 N_D1_c_106_n N_A_27_409#_c_217_n 0.0114482f $X=0.81 $Y=0.86 $X2=0 $Y2=0
cc_123 N_D1_c_110_n N_A_27_409#_c_217_n 7.358e-19 $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_124 N_D1_c_111_n N_A_27_409#_c_217_n 0.011068f $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_125 N_D1_M1000_g N_A_232_409#_c_480_n 8.27996e-19 $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_126 N_D1_M1000_g N_A_232_409#_c_481_n 0.00231035f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_127 N_D1_M1000_g N_A_232_409#_c_487_n 7.28154e-19 $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_128 N_D1_M1000_g N_VPWR_c_525_n 0.0086001f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_129 N_D1_M1000_g N_VPWR_c_520_n 0.0163652f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_130 N_D1_M1001_g N_VGND_c_629_n 0.0127913f $X=0.495 $Y=0.445 $X2=0 $Y2=0
cc_131 N_D1_M1014_g N_VGND_c_629_n 0.00161202f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_132 N_D1_c_108_n N_VGND_c_629_n 0.0064747f $X=0.385 $Y=0.86 $X2=0 $Y2=0
cc_133 N_D1_c_111_n N_VGND_c_629_n 0.0266616f $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_134 N_D1_M1001_g N_VGND_c_632_n 0.00486043f $X=0.495 $Y=0.445 $X2=0 $Y2=0
cc_135 N_D1_M1014_g N_VGND_c_632_n 0.00359757f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_136 N_D1_M1001_g N_VGND_c_636_n 0.00573768f $X=0.495 $Y=0.445 $X2=0 $Y2=0
cc_137 N_D1_c_106_n N_VGND_c_636_n 0.00107318f $X=0.81 $Y=0.86 $X2=0 $Y2=0
cc_138 N_D1_M1014_g N_VGND_c_636_n 0.00533371f $X=0.885 $Y=0.445 $X2=0 $Y2=0
cc_139 N_D1_c_111_n N_VGND_c_636_n 0.00372933f $X=0.365 $Y=1.02 $X2=0 $Y2=0
cc_140 N_C1_c_153_n N_A_27_409#_M1013_g 0.0179726f $X=1.675 $Y=0.73 $X2=0 $Y2=0
cc_141 N_C1_c_157_n N_A_27_409#_M1013_g 0.00279816f $X=1.15 $Y=1.175 $X2=0 $Y2=0
cc_142 N_C1_M1006_g N_A_27_409#_c_223_n 0.00375854f $X=1.035 $Y=2.545 $X2=0
+ $Y2=0
cc_143 N_C1_M1006_g N_A_27_409#_c_224_n 8.51849e-19 $X=1.035 $Y=2.545 $X2=0
+ $Y2=0
cc_144 N_C1_c_151_n N_A_27_409#_c_209_n 0.00877411f $X=1.315 $Y=0.73 $X2=0 $Y2=0
cc_145 N_C1_c_153_n N_A_27_409#_c_209_n 0.00144802f $X=1.675 $Y=0.73 $X2=0 $Y2=0
cc_146 N_C1_c_154_n N_A_27_409#_c_209_n 0.00580246f $X=1.315 $Y=0.805 $X2=0
+ $Y2=0
cc_147 C1 N_A_27_409#_c_210_n 0.0482234f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_148 N_C1_c_156_n N_A_27_409#_c_210_n 0.0102014f $X=1.225 $Y=1.34 $X2=0 $Y2=0
cc_149 N_C1_c_157_n N_A_27_409#_c_210_n 0.00342318f $X=1.15 $Y=1.175 $X2=0 $Y2=0
cc_150 N_C1_c_152_n N_A_27_409#_c_211_n 0.0163715f $X=1.6 $Y=0.805 $X2=0 $Y2=0
cc_151 N_C1_c_154_n N_A_27_409#_c_211_n 0.00357648f $X=1.315 $Y=0.805 $X2=0
+ $Y2=0
cc_152 C1 N_A_27_409#_c_211_n 0.00897633f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_153 N_C1_c_157_n N_A_27_409#_c_211_n 0.00529657f $X=1.15 $Y=1.175 $X2=0 $Y2=0
cc_154 C1 N_A_27_409#_c_212_n 0.0268001f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_155 N_C1_c_157_n N_A_27_409#_c_212_n 0.00575281f $X=1.15 $Y=1.175 $X2=0 $Y2=0
cc_156 N_C1_c_154_n N_A_27_409#_c_217_n 7.83618e-19 $X=1.315 $Y=0.805 $X2=0
+ $Y2=0
cc_157 C1 N_A_27_409#_c_217_n 0.0172817f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_158 N_C1_c_156_n N_A_27_409#_c_217_n 0.00762581f $X=1.225 $Y=1.34 $X2=0 $Y2=0
cc_159 N_C1_c_157_n N_A_27_409#_c_217_n 0.00242554f $X=1.15 $Y=1.175 $X2=0 $Y2=0
cc_160 N_C1_c_152_n N_A_27_409#_c_220_n 0.00139458f $X=1.6 $Y=0.805 $X2=0 $Y2=0
cc_161 C1 N_A_27_409#_c_220_n 0.00290253f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_162 N_C1_c_157_n N_A_27_409#_c_220_n 0.0253441f $X=1.15 $Y=1.175 $X2=0 $Y2=0
cc_163 N_C1_M1006_g N_A_232_409#_c_480_n 0.0063703f $X=1.035 $Y=2.545 $X2=0
+ $Y2=0
cc_164 C1 N_A_232_409#_c_480_n 0.0214646f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_165 N_C1_c_156_n N_A_232_409#_c_480_n 0.00177874f $X=1.225 $Y=1.34 $X2=0
+ $Y2=0
cc_166 N_C1_M1006_g N_A_232_409#_c_481_n 0.0110688f $X=1.035 $Y=2.545 $X2=0
+ $Y2=0
cc_167 N_C1_M1006_g N_A_232_409#_c_487_n 0.00361451f $X=1.035 $Y=2.545 $X2=0
+ $Y2=0
cc_168 N_C1_M1006_g N_VPWR_c_521_n 0.00233601f $X=1.035 $Y=2.545 $X2=0 $Y2=0
cc_169 N_C1_M1006_g N_VPWR_c_525_n 0.0086001f $X=1.035 $Y=2.545 $X2=0 $Y2=0
cc_170 N_C1_M1006_g N_VPWR_c_520_n 0.0166232f $X=1.035 $Y=2.545 $X2=0 $Y2=0
cc_171 N_C1_c_151_n N_VGND_c_630_n 0.00231629f $X=1.315 $Y=0.73 $X2=0 $Y2=0
cc_172 N_C1_c_153_n N_VGND_c_630_n 0.0119143f $X=1.675 $Y=0.73 $X2=0 $Y2=0
cc_173 N_C1_c_151_n N_VGND_c_632_n 0.00549284f $X=1.315 $Y=0.73 $X2=0 $Y2=0
cc_174 N_C1_c_152_n N_VGND_c_632_n 4.87571e-19 $X=1.6 $Y=0.805 $X2=0 $Y2=0
cc_175 N_C1_c_153_n N_VGND_c_632_n 0.00486043f $X=1.675 $Y=0.73 $X2=0 $Y2=0
cc_176 N_C1_c_151_n N_VGND_c_636_n 0.00612472f $X=1.315 $Y=0.73 $X2=0 $Y2=0
cc_177 N_C1_c_152_n N_VGND_c_636_n 6.51792e-19 $X=1.6 $Y=0.805 $X2=0 $Y2=0
cc_178 N_C1_c_153_n N_VGND_c_636_n 0.00436085f $X=1.675 $Y=0.73 $X2=0 $Y2=0
cc_179 N_A_27_409#_c_214_n N_B1_c_343_n 0.0110491f $X=3.26 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A_27_409#_c_215_n N_B1_c_344_n 0.0167004f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_181 N_A_27_409#_c_214_n N_B1_c_345_n 0.00170639f $X=3.26 $Y=0.495 $X2=0 $Y2=0
cc_182 N_A_27_409#_c_215_n N_B1_c_346_n 0.00373203f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_183 N_A_27_409#_c_218_n N_B1_c_346_n 9.68574e-19 $X=2.75 $Y=0.99 $X2=0 $Y2=0
cc_184 N_A_27_409#_c_219_n N_B1_c_346_n 0.0016279f $X=3.26 $Y=0.91 $X2=0 $Y2=0
cc_185 N_A_27_409#_c_214_n N_B1_c_348_n 0.00296195f $X=3.26 $Y=0.495 $X2=0 $Y2=0
cc_186 N_A_27_409#_c_215_n N_B1_c_348_n 0.00407103f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_187 N_A_27_409#_c_219_n N_B1_c_348_n 0.00209642f $X=3.26 $Y=0.91 $X2=0 $Y2=0
cc_188 N_A_27_409#_c_220_n N_B1_c_348_n 0.00862297f $X=2.465 $Y=1.307 $X2=0
+ $Y2=0
cc_189 N_A_27_409#_c_215_n B1 0.0216694f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_190 N_A_27_409#_c_218_n B1 0.0109442f $X=2.75 $Y=0.99 $X2=0 $Y2=0
cc_191 N_A_27_409#_c_219_n B1 0.00491731f $X=3.26 $Y=0.91 $X2=0 $Y2=0
cc_192 N_A_27_409#_c_220_n B1 0.00159028f $X=2.465 $Y=1.307 $X2=0 $Y2=0
cc_193 N_A_27_409#_c_215_n N_B1_c_350_n 4.43313e-19 $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_194 N_A_27_409#_c_218_n N_B1_c_350_n 0.00135979f $X=2.75 $Y=0.99 $X2=0 $Y2=0
cc_195 N_A_27_409#_c_219_n N_B1_c_350_n 2.64278e-19 $X=3.26 $Y=0.91 $X2=0 $Y2=0
cc_196 N_A_27_409#_c_220_n N_B1_c_350_n 0.00817366f $X=2.465 $Y=1.307 $X2=0
+ $Y2=0
cc_197 N_A_27_409#_c_215_n N_A2_M1004_g 0.0142104f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_198 N_A_27_409#_c_216_n N_A2_M1004_g 0.0019649f $X=4.87 $Y=0.495 $X2=0 $Y2=0
cc_199 N_A_27_409#_c_215_n A2 0.0247881f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_200 N_A_27_409#_c_215_n N_A2_c_407_n 0.00174562f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_201 N_A_27_409#_c_215_n N_A1_M1005_g 0.0124846f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_202 N_A_27_409#_c_216_n N_A1_M1005_g 0.0130843f $X=4.87 $Y=0.495 $X2=0 $Y2=0
cc_203 N_A_27_409#_c_215_n A1 0.0483714f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_204 N_A_27_409#_c_215_n N_A1_c_449_n 0.0048437f $X=4.705 $Y=0.91 $X2=0 $Y2=0
cc_205 N_A_27_409#_c_224_n A_134_409# 0.00570883f $X=0.71 $Y=2.11 $X2=-0.19
+ $Y2=-0.245
cc_206 N_A_27_409#_M1015_g N_A_232_409#_c_480_n 0.00779127f $X=2.265 $Y=2.45
+ $X2=0 $Y2=0
cc_207 N_A_27_409#_c_224_n N_A_232_409#_c_480_n 0.00529447f $X=0.71 $Y=2.11
+ $X2=0 $Y2=0
cc_208 N_A_27_409#_M1015_g N_A_232_409#_c_481_n 0.00395264f $X=2.265 $Y=2.45
+ $X2=0 $Y2=0
cc_209 N_A_27_409#_M1015_g N_A_232_409#_c_482_n 0.0238696f $X=2.265 $Y=2.45
+ $X2=0 $Y2=0
cc_210 N_A_27_409#_c_212_n N_A_232_409#_c_482_n 0.0101213f $X=1.89 $Y=1.285
+ $X2=0 $Y2=0
cc_211 N_A_27_409#_c_220_n N_A_232_409#_c_482_n 0.00338882f $X=2.465 $Y=1.307
+ $X2=0 $Y2=0
cc_212 N_A_27_409#_M1015_g N_VPWR_c_521_n 0.0199425f $X=2.265 $Y=2.45 $X2=0
+ $Y2=0
cc_213 N_A_27_409#_M1015_g N_VPWR_c_523_n 0.0085504f $X=2.265 $Y=2.45 $X2=0
+ $Y2=0
cc_214 N_A_27_409#_c_223_n N_VPWR_c_525_n 0.0220321f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_215 N_A_27_409#_M1015_g N_VPWR_c_520_n 0.00817624f $X=2.265 $Y=2.45 $X2=0
+ $Y2=0
cc_216 N_A_27_409#_c_223_n N_VPWR_c_520_n 0.0125808f $X=0.28 $Y=2.9 $X2=0 $Y2=0
cc_217 N_A_27_409#_M1013_g N_X_c_564_n 0.00572464f $X=2.105 $Y=0.445 $X2=0 $Y2=0
cc_218 N_A_27_409#_M1015_g N_X_c_564_n 0.00848914f $X=2.265 $Y=2.45 $X2=0 $Y2=0
cc_219 N_A_27_409#_M1008_g N_X_c_564_n 0.00819445f $X=2.465 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A_27_409#_c_211_n N_X_c_564_n 0.0130055f $X=1.725 $Y=0.91 $X2=0 $Y2=0
cc_221 N_A_27_409#_c_212_n N_X_c_564_n 0.0546282f $X=1.89 $Y=1.285 $X2=0 $Y2=0
cc_222 N_A_27_409#_c_218_n N_X_c_564_n 0.046437f $X=2.75 $Y=0.99 $X2=0 $Y2=0
cc_223 N_A_27_409#_c_220_n N_X_c_564_n 0.0363387f $X=2.465 $Y=1.307 $X2=0 $Y2=0
cc_224 N_A_27_409#_M1008_g N_X_c_565_n 0.0154349f $X=2.465 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A_27_409#_c_214_n N_X_c_565_n 0.0253054f $X=3.26 $Y=0.495 $X2=0 $Y2=0
cc_226 N_A_27_409#_c_218_n N_X_c_565_n 0.0196036f $X=2.75 $Y=0.99 $X2=0 $Y2=0
cc_227 N_A_27_409#_c_220_n N_X_c_565_n 0.00194564f $X=2.465 $Y=1.307 $X2=0 $Y2=0
cc_228 N_A_27_409#_M1015_g N_X_c_579_n 0.0177462f $X=2.265 $Y=2.45 $X2=0 $Y2=0
cc_229 N_A_27_409#_c_218_n X 0.00698534f $X=2.75 $Y=0.99 $X2=0 $Y2=0
cc_230 N_A_27_409#_c_220_n X 0.00697141f $X=2.465 $Y=1.307 $X2=0 $Y2=0
cc_231 N_A_27_409#_c_209_n N_VGND_c_629_n 0.0236358f $X=1.1 $Y=0.47 $X2=0 $Y2=0
cc_232 N_A_27_409#_M1013_g N_VGND_c_630_n 0.00976183f $X=2.105 $Y=0.445 $X2=0
+ $Y2=0
cc_233 N_A_27_409#_M1008_g N_VGND_c_630_n 0.00158408f $X=2.465 $Y=0.445 $X2=0
+ $Y2=0
cc_234 N_A_27_409#_c_209_n N_VGND_c_630_n 0.0132397f $X=1.1 $Y=0.47 $X2=0 $Y2=0
cc_235 N_A_27_409#_c_211_n N_VGND_c_630_n 0.0227656f $X=1.725 $Y=0.91 $X2=0
+ $Y2=0
cc_236 N_A_27_409#_c_220_n N_VGND_c_630_n 9.7121e-19 $X=2.465 $Y=1.307 $X2=0
+ $Y2=0
cc_237 N_A_27_409#_c_214_n N_VGND_c_631_n 0.0127138f $X=3.26 $Y=0.495 $X2=0
+ $Y2=0
cc_238 N_A_27_409#_c_215_n N_VGND_c_631_n 0.0200008f $X=4.705 $Y=0.91 $X2=0
+ $Y2=0
cc_239 N_A_27_409#_c_216_n N_VGND_c_631_n 0.0120387f $X=4.87 $Y=0.495 $X2=0
+ $Y2=0
cc_240 N_A_27_409#_c_209_n N_VGND_c_632_n 0.0305995f $X=1.1 $Y=0.47 $X2=0 $Y2=0
cc_241 N_A_27_409#_M1013_g N_VGND_c_634_n 0.00486043f $X=2.105 $Y=0.445 $X2=0
+ $Y2=0
cc_242 N_A_27_409#_M1008_g N_VGND_c_634_n 0.00359964f $X=2.465 $Y=0.445 $X2=0
+ $Y2=0
cc_243 N_A_27_409#_c_214_n N_VGND_c_634_n 0.0220321f $X=3.26 $Y=0.495 $X2=0
+ $Y2=0
cc_244 N_A_27_409#_c_216_n N_VGND_c_635_n 0.0220321f $X=4.87 $Y=0.495 $X2=0
+ $Y2=0
cc_245 N_A_27_409#_M1014_d N_VGND_c_636_n 0.0022543f $X=0.96 $Y=0.235 $X2=0
+ $Y2=0
cc_246 N_A_27_409#_M1013_g N_VGND_c_636_n 0.00814425f $X=2.105 $Y=0.445 $X2=0
+ $Y2=0
cc_247 N_A_27_409#_M1008_g N_VGND_c_636_n 0.00661248f $X=2.465 $Y=0.445 $X2=0
+ $Y2=0
cc_248 N_A_27_409#_c_209_n N_VGND_c_636_n 0.0205958f $X=1.1 $Y=0.47 $X2=0 $Y2=0
cc_249 N_A_27_409#_c_211_n N_VGND_c_636_n 0.0147838f $X=1.725 $Y=0.91 $X2=0
+ $Y2=0
cc_250 N_A_27_409#_c_213_n N_VGND_c_636_n 0.00627113f $X=3.095 $Y=0.91 $X2=0
+ $Y2=0
cc_251 N_A_27_409#_c_214_n N_VGND_c_636_n 0.0125808f $X=3.26 $Y=0.495 $X2=0
+ $Y2=0
cc_252 N_A_27_409#_c_215_n N_VGND_c_636_n 0.0300466f $X=4.705 $Y=0.91 $X2=0
+ $Y2=0
cc_253 N_A_27_409#_c_216_n N_VGND_c_636_n 0.0125808f $X=4.87 $Y=0.495 $X2=0
+ $Y2=0
cc_254 N_A_27_409#_c_218_n N_VGND_c_636_n 0.00293632f $X=2.75 $Y=0.99 $X2=0
+ $Y2=0
cc_255 N_A_27_409#_c_209_n A_114_47# 0.00442806f $X=1.1 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_256 N_B1_c_347_n N_A2_c_403_n 0.0120198f $X=3.53 $Y=1.68 $X2=0 $Y2=0
cc_257 N_B1_M1011_g N_A2_M1003_g 0.0172401f $X=3.57 $Y=2.545 $X2=0 $Y2=0
cc_258 N_B1_c_345_n N_A2_M1004_g 0.0197172f $X=3.835 $Y=0.78 $X2=0 $Y2=0
cc_259 N_B1_c_346_n N_A2_M1004_g 0.00501416f $X=3.53 $Y=1.175 $X2=0 $Y2=0
cc_260 N_B1_c_353_n N_A2_c_405_n 0.0120198f $X=3.53 $Y=1.845 $X2=0 $Y2=0
cc_261 B1 A2 0.0438819f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_262 N_B1_c_350_n A2 8.23261e-19 $X=3.53 $Y=1.34 $X2=0 $Y2=0
cc_263 B1 N_A2_c_407_n 0.0042029f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_264 N_B1_c_350_n N_A2_c_407_n 0.0120198f $X=3.53 $Y=1.34 $X2=0 $Y2=0
cc_265 N_B1_M1011_g N_A_232_409#_c_483_n 0.00632946f $X=3.57 $Y=2.545 $X2=0
+ $Y2=0
cc_266 N_B1_c_353_n N_A_232_409#_c_483_n 6.13682e-19 $X=3.53 $Y=1.845 $X2=0
+ $Y2=0
cc_267 B1 N_A_232_409#_c_483_n 0.00867382f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_268 N_B1_M1011_g N_A_232_409#_c_484_n 0.00951569f $X=3.57 $Y=2.545 $X2=0
+ $Y2=0
cc_269 N_B1_M1011_g N_A_232_409#_c_503_n 0.00293538f $X=3.57 $Y=2.545 $X2=0
+ $Y2=0
cc_270 N_B1_M1011_g N_VPWR_c_522_n 8.49223e-19 $X=3.57 $Y=2.545 $X2=0 $Y2=0
cc_271 N_B1_M1011_g N_VPWR_c_523_n 0.00826654f $X=3.57 $Y=2.545 $X2=0 $Y2=0
cc_272 N_B1_M1011_g N_VPWR_c_520_n 0.0158042f $X=3.57 $Y=2.545 $X2=0 $Y2=0
cc_273 N_B1_c_343_n N_X_c_565_n 8.6009e-19 $X=3.475 $Y=0.78 $X2=0 $Y2=0
cc_274 N_B1_M1011_g X 0.00292976f $X=3.57 $Y=2.545 $X2=0 $Y2=0
cc_275 N_B1_M1011_g N_A_739_409#_c_593_n 0.00366581f $X=3.57 $Y=2.545 $X2=0
+ $Y2=0
cc_276 B1 N_A_739_409#_c_593_n 0.00372527f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_277 N_B1_M1011_g N_A_739_409#_c_594_n 0.0156174f $X=3.57 $Y=2.545 $X2=0 $Y2=0
cc_278 N_B1_c_343_n N_VGND_c_631_n 0.00189426f $X=3.475 $Y=0.78 $X2=0 $Y2=0
cc_279 N_B1_c_345_n N_VGND_c_631_n 0.0106455f $X=3.835 $Y=0.78 $X2=0 $Y2=0
cc_280 N_B1_c_343_n N_VGND_c_634_n 0.00502664f $X=3.475 $Y=0.78 $X2=0 $Y2=0
cc_281 N_B1_c_344_n N_VGND_c_634_n 4.57848e-19 $X=3.76 $Y=0.855 $X2=0 $Y2=0
cc_282 N_B1_c_345_n N_VGND_c_634_n 0.00445056f $X=3.835 $Y=0.78 $X2=0 $Y2=0
cc_283 N_B1_c_343_n N_VGND_c_636_n 0.00651958f $X=3.475 $Y=0.78 $X2=0 $Y2=0
cc_284 N_B1_c_344_n N_VGND_c_636_n 6.33118e-19 $X=3.76 $Y=0.855 $X2=0 $Y2=0
cc_285 N_B1_c_345_n N_VGND_c_636_n 0.0041956f $X=3.835 $Y=0.78 $X2=0 $Y2=0
cc_286 N_A2_M1004_g N_A1_M1005_g 0.0224031f $X=4.265 $Y=0.495 $X2=0 $Y2=0
cc_287 N_A2_M1003_g N_A1_M1012_g 0.0326465f $X=4.1 $Y=2.545 $X2=0 $Y2=0
cc_288 N_A2_c_403_n N_A1_c_447_n 0.0224031f $X=4.137 $Y=1.643 $X2=0 $Y2=0
cc_289 N_A2_c_405_n N_A1_c_452_n 0.0224031f $X=4.137 $Y=1.845 $X2=0 $Y2=0
cc_290 A2 A1 0.0540775f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_291 N_A2_c_407_n A1 0.00521108f $X=4.1 $Y=1.34 $X2=0 $Y2=0
cc_292 A2 N_A1_c_449_n 5.88676e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_293 N_A2_c_407_n N_A1_c_449_n 0.0224031f $X=4.1 $Y=1.34 $X2=0 $Y2=0
cc_294 N_A2_M1003_g N_VPWR_c_522_n 0.0163992f $X=4.1 $Y=2.545 $X2=0 $Y2=0
cc_295 N_A2_M1003_g N_VPWR_c_523_n 0.00769046f $X=4.1 $Y=2.545 $X2=0 $Y2=0
cc_296 N_A2_M1003_g N_VPWR_c_520_n 0.0134474f $X=4.1 $Y=2.545 $X2=0 $Y2=0
cc_297 N_A2_M1003_g N_A_739_409#_c_593_n 9.81754e-19 $X=4.1 $Y=2.545 $X2=0 $Y2=0
cc_298 N_A2_c_405_n N_A_739_409#_c_593_n 3.03142e-19 $X=4.137 $Y=1.845 $X2=0
+ $Y2=0
cc_299 A2 N_A_739_409#_c_593_n 0.00534367f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_300 N_A2_M1003_g N_A_739_409#_c_594_n 0.0159281f $X=4.1 $Y=2.545 $X2=0 $Y2=0
cc_301 N_A2_M1003_g N_A_739_409#_c_595_n 0.0182584f $X=4.1 $Y=2.545 $X2=0 $Y2=0
cc_302 N_A2_c_405_n N_A_739_409#_c_595_n 0.00338858f $X=4.137 $Y=1.845 $X2=0
+ $Y2=0
cc_303 A2 N_A_739_409#_c_595_n 0.0192947f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_304 N_A2_M1003_g N_A_739_409#_c_597_n 8.97659e-19 $X=4.1 $Y=2.545 $X2=0 $Y2=0
cc_305 N_A2_M1004_g N_VGND_c_631_n 0.0109044f $X=4.265 $Y=0.495 $X2=0 $Y2=0
cc_306 N_A2_M1004_g N_VGND_c_635_n 0.00445056f $X=4.265 $Y=0.495 $X2=0 $Y2=0
cc_307 N_A2_M1004_g N_VGND_c_636_n 0.0042789f $X=4.265 $Y=0.495 $X2=0 $Y2=0
cc_308 N_A1_M1012_g N_VPWR_c_522_n 0.00680165f $X=4.705 $Y=2.545 $X2=0 $Y2=0
cc_309 N_A1_M1012_g N_VPWR_c_526_n 0.0086001f $X=4.705 $Y=2.545 $X2=0 $Y2=0
cc_310 N_A1_M1012_g N_VPWR_c_520_n 0.0164378f $X=4.705 $Y=2.545 $X2=0 $Y2=0
cc_311 N_A1_M1012_g N_A_739_409#_c_594_n 9.07015e-19 $X=4.705 $Y=2.545 $X2=0
+ $Y2=0
cc_312 N_A1_M1012_g N_A_739_409#_c_595_n 0.0189917f $X=4.705 $Y=2.545 $X2=0
+ $Y2=0
cc_313 A1 N_A_739_409#_c_595_n 0.0271277f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_314 N_A1_M1012_g N_A_739_409#_c_596_n 0.00114325f $X=4.705 $Y=2.545 $X2=0
+ $Y2=0
cc_315 N_A1_c_452_n N_A_739_409#_c_596_n 0.00213543f $X=4.745 $Y=1.845 $X2=0
+ $Y2=0
cc_316 A1 N_A_739_409#_c_596_n 0.028933f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_317 N_A1_M1012_g N_A_739_409#_c_597_n 0.0147872f $X=4.705 $Y=2.545 $X2=0
+ $Y2=0
cc_318 N_A1_M1005_g N_VGND_c_631_n 0.0019059f $X=4.655 $Y=0.495 $X2=0 $Y2=0
cc_319 N_A1_M1005_g N_VGND_c_635_n 0.00502664f $X=4.655 $Y=0.495 $X2=0 $Y2=0
cc_320 N_A1_M1005_g N_VGND_c_636_n 0.00642785f $X=4.655 $Y=0.495 $X2=0 $Y2=0
cc_321 N_A_232_409#_c_482_n N_VPWR_M1015_s 0.00719074f $X=3.14 $Y=2.445
+ $X2=-0.19 $Y2=1.655
cc_322 N_A_232_409#_c_481_n N_VPWR_c_521_n 0.0172695f $X=1.3 $Y=2.9 $X2=0 $Y2=0
cc_323 N_A_232_409#_c_482_n N_VPWR_c_521_n 0.0204535f $X=3.14 $Y=2.445 $X2=0
+ $Y2=0
cc_324 N_A_232_409#_c_484_n N_VPWR_c_523_n 0.0220321f $X=3.305 $Y=2.9 $X2=0
+ $Y2=0
cc_325 N_A_232_409#_c_481_n N_VPWR_c_525_n 0.0220321f $X=1.3 $Y=2.9 $X2=0 $Y2=0
cc_326 N_A_232_409#_c_481_n N_VPWR_c_520_n 0.0125808f $X=1.3 $Y=2.9 $X2=0 $Y2=0
cc_327 N_A_232_409#_c_482_n N_VPWR_c_520_n 0.0485484f $X=3.14 $Y=2.445 $X2=0
+ $Y2=0
cc_328 N_A_232_409#_c_484_n N_VPWR_c_520_n 0.0125808f $X=3.305 $Y=2.9 $X2=0
+ $Y2=0
cc_329 N_A_232_409#_c_482_n N_X_M1015_d 0.00789112f $X=3.14 $Y=2.445 $X2=0 $Y2=0
cc_330 N_A_232_409#_c_482_n N_X_c_579_n 0.0111946f $X=3.14 $Y=2.445 $X2=0 $Y2=0
cc_331 N_A_232_409#_c_482_n X 0.0223717f $X=3.14 $Y=2.445 $X2=0 $Y2=0
cc_332 N_A_232_409#_c_483_n X 0.00756497f $X=3.305 $Y=2.19 $X2=0 $Y2=0
cc_333 N_A_232_409#_c_483_n N_A_739_409#_c_593_n 0.0119061f $X=3.305 $Y=2.19
+ $X2=0 $Y2=0
cc_334 N_A_232_409#_c_483_n N_A_739_409#_c_594_n 0.0108061f $X=3.305 $Y=2.19
+ $X2=0 $Y2=0
cc_335 N_A_232_409#_c_484_n N_A_739_409#_c_594_n 0.0352186f $X=3.305 $Y=2.9
+ $X2=0 $Y2=0
cc_336 N_A_232_409#_c_503_n N_A_739_409#_c_594_n 0.0119061f $X=3.305 $Y=2.445
+ $X2=0 $Y2=0
cc_337 N_VPWR_c_522_n N_A_739_409#_c_594_n 0.0454646f $X=4.365 $Y=2.54 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_523_n N_A_739_409#_c_594_n 0.021949f $X=4.2 $Y=3.33 $X2=0 $Y2=0
cc_339 N_VPWR_c_520_n N_A_739_409#_c_594_n 0.0124703f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_340 N_VPWR_M1003_d N_A_739_409#_c_595_n 0.00262408f $X=4.225 $Y=2.045 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_522_n N_A_739_409#_c_595_n 0.0204924f $X=4.365 $Y=2.54 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_522_n N_A_739_409#_c_597_n 0.0181941f $X=4.365 $Y=2.54 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_526_n N_A_739_409#_c_597_n 0.0220321f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_520_n N_A_739_409#_c_597_n 0.0125808f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_345 N_X_c_565_n N_VGND_c_634_n 0.0346699f $X=2.68 $Y=0.455 $X2=0 $Y2=0
cc_346 N_X_M1008_d N_VGND_c_636_n 0.00233022f $X=2.54 $Y=0.235 $X2=0 $Y2=0
cc_347 N_X_c_565_n N_VGND_c_636_n 0.0225227f $X=2.68 $Y=0.455 $X2=0 $Y2=0
cc_348 N_X_c_564_n A_436_47# 2.77635e-19 $X=2.32 $Y=1.92 $X2=-0.19 $Y2=-0.245
cc_349 N_X_c_565_n A_436_47# 0.00122016f $X=2.68 $Y=0.455 $X2=-0.19 $Y2=-0.245
cc_350 N_VGND_c_636_n A_114_47# 0.00566796f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
cc_351 N_VGND_c_636_n A_278_47# 0.00303453f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
cc_352 N_VGND_c_636_n A_436_47# 0.00359567f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
