* File: sky130_fd_sc_lp__and4bb_1.spice
* Created: Wed Sep  2 09:34:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4bb_1.pex.spice"
.subckt sky130_fd_sc_lp__and4bb_1  VNB VPB A_N B_N C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_N_M1009_g N_A_27_51#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_196_51#_M1000_d N_B_N_M1000_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1013 A_427_131# N_A_27_51#_M1013_g N_A_344_131#_M1013_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1007 A_499_131# N_A_196_51#_M1007_g A_427_131# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1002 A_607_131# N_C_M1002_g A_499_131# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=39.996 M=1 R=2.8 SA=75001.1 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_D_M1010_g A_607_131# VNB NSHORT L=0.15 W=0.42 AD=0.0896
+ AS=0.0441 PD=0.81 PS=0.63 NRD=9.996 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1012 N_X_M1012_d N_A_344_131#_M1012_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=4.284 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_27_51#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_196_51#_M1005_d N_B_N_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_344_131#_M1006_d N_A_27_51#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_196_51#_M1004_g N_A_344_131#_M1006_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=7.0329 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_344_131#_M1001_d N_C_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=11.7215 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_D_M1008_g N_A_344_131#_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0588 PD=0.8175 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1011 N_X_M1011_d N_A_344_131#_M1011_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=4.9447 M=1 R=8.4 SA=75000.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__and4bb_1.pxi.spice"
*
.ends
*
*
