# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__a21bo_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a21bo_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 1.250000 1.925000 1.550000 ;
        RECT 1.595000 1.550000 2.825000 1.720000 ;
        RECT 2.495000 1.720000 2.825000 1.935000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.280000 1.355000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.035000 3.335000 1.780000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.265000 0.445000 0.715000 ;
        RECT 0.090000 0.715000 0.260000 2.025000 ;
        RECT 0.090000 2.025000 0.495000 3.065000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.840000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 4.030000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.440000  0.895000 2.055000 1.065000 ;
      RECT 0.440000  1.065000 0.845000 1.565000 ;
      RECT 0.675000  1.565000 0.845000 1.960000 ;
      RECT 0.675000  1.960000 2.095000 2.130000 ;
      RECT 0.695000  2.310000 1.025000 3.245000 ;
      RECT 0.905000  0.085000 1.235000 0.715000 ;
      RECT 1.235000  2.310000 1.565000 2.895000 ;
      RECT 1.235000  2.895000 2.655000 3.065000 ;
      RECT 1.725000  0.265000 2.055000 0.895000 ;
      RECT 1.765000  2.130000 2.095000 2.715000 ;
      RECT 2.250000  0.685000 3.715000 0.855000 ;
      RECT 2.250000  0.855000 2.580000 1.135000 ;
      RECT 2.325000  2.115000 2.655000 2.895000 ;
      RECT 2.515000  0.085000 2.845000 0.505000 ;
      RECT 2.855000  2.115000 3.185000 3.245000 ;
      RECT 3.305000  0.265000 3.635000 0.685000 ;
      RECT 3.385000  2.075000 3.715000 3.065000 ;
      RECT 3.545000  0.855000 3.715000 2.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__a21bo_lp
END LIBRARY
