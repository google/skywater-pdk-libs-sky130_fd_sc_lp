* File: sky130_fd_sc_lp__iso0n_lp2.pex.spice
* Created: Fri Aug 28 10:40:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__ISO0N_LP2%A 1 2 3 5 9 17 18 22 23
c41 2 0 2.72973e-20 $X=0.455 $Y=1.03
r42 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=1.12 $X2=0.29 $Y2=1.12
r43 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r44 17 23 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.12
r45 13 22 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.29 $Y=1.475
+ $X2=0.29 $Y2=1.12
r46 11 22 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.29 $Y=1.105
+ $X2=0.29 $Y2=1.12
r47 7 9 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.685 $Y=0.955
+ $X2=0.685 $Y2=0.535
r48 3 13 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.635 $Y=1.55
+ $X2=0.29 $Y2=1.55
r49 3 5 228.577 $w=2.5e-07 $l=9.2e-07 $layer=POLY_cond $X=0.635 $Y=1.625
+ $X2=0.635 $Y2=2.545
r50 2 11 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.455 $Y=1.03
+ $X2=0.29 $Y2=1.105
r51 1 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.61 $Y=1.03
+ $X2=0.685 $Y2=0.955
r52 1 2 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.61 $Y=1.03
+ $X2=0.455 $Y2=1.03
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0N_LP2%SLEEP_B 3 7 9 10 14
r43 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.165 $Y=1.68
+ $X2=1.165 $Y2=1.515
r44 9 10 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=1.165 $Y=1.68
+ $X2=1.68 $Y2=1.68
r45 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.68 $X2=1.165 $Y2=1.68
r46 5 14 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.165 $Y=1.845
+ $X2=1.165 $Y2=1.68
r47 5 7 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.165 $Y=1.845 $X2=1.165
+ $Y2=2.545
r48 3 16 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.075 $Y=0.535
+ $X2=1.075 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0N_LP2%A_65_65# 1 2 9 13 17 20 25 29 33 35 37 38
+ 41
r77 37 38 8.71334 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.857 $Y=2.19
+ $X2=0.857 $Y2=2.025
r78 30 41 21.0218 $w=3.21e-07 $l=1.4e-07 $layer=POLY_cond $X=1.555 $Y=1.202
+ $X2=1.695 $Y2=1.202
r79 30 39 7.50779 $w=3.21e-07 $l=5e-08 $layer=POLY_cond $X=1.555 $Y=1.202
+ $X2=1.505 $Y2=1.202
r80 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.555
+ $Y=1.11 $X2=1.555 $Y2=1.11
r81 27 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=1.11
+ $X2=0.735 $Y2=1.11
r82 27 29 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=0.82 $Y=1.11
+ $X2=1.555 $Y2=1.11
r83 23 37 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=0.857 $Y=2.232
+ $X2=0.857 $Y2=2.19
r84 23 25 18.5502 $w=4.13e-07 $l=6.68e-07 $layer=LI1_cond $X=0.857 $Y=2.232
+ $X2=0.857 $Y2=2.9
r85 21 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=1.275
+ $X2=0.735 $Y2=1.11
r86 21 38 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.735 $Y=1.275
+ $X2=0.735 $Y2=2.025
r87 20 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=0.945
+ $X2=0.735 $Y2=1.11
r88 19 33 9.10704 $w=3.55e-07 $l=3.62181e-07 $layer=LI1_cond $X=0.735 $Y=0.765
+ $X2=0.47 $Y2=0.535
r89 19 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.735 $Y=0.765
+ $X2=0.735 $Y2=0.945
r90 15 41 30.0312 $w=3.21e-07 $l=3.42708e-07 $layer=POLY_cond $X=1.895 $Y=0.945
+ $X2=1.695 $Y2=1.202
r91 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.895 $Y=0.945
+ $X2=1.895 $Y2=0.535
r92 11 41 8.70639 $w=2.5e-07 $l=2.58e-07 $layer=POLY_cond $X=1.695 $Y=1.46
+ $X2=1.695 $Y2=1.202
r93 11 13 269.572 $w=2.5e-07 $l=1.085e-06 $layer=POLY_cond $X=1.695 $Y=1.46
+ $X2=1.695 $Y2=2.545
r94 7 39 20.5661 $w=1.5e-07 $l=2.57e-07 $layer=POLY_cond $X=1.505 $Y=0.945
+ $X2=1.505 $Y2=1.202
r95 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.505 $Y=0.945
+ $X2=1.505 $Y2=0.535
r96 2 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.76
+ $Y=2.045 $X2=0.9 $Y2=2.19
r97 2 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.76
+ $Y=2.045 $X2=0.9 $Y2=2.9
r98 1 33 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.325
+ $Y=0.325 $X2=0.47 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0N_LP2%VPWR 1 2 7 9 15 20 21 22 29 30
r29 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 24 33 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=3.33
+ $X2=0.235 $Y2=3.33
r32 24 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=0.47 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 22 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 22 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 22 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 20 26 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.2 $Y2=3.33
r37 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.43 $Y2=3.33
r38 19 29 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.43 $Y2=3.33
r40 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.43 $Y=2.19 $X2=1.43
+ $Y2=2.9
r41 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.43 $Y=3.245
+ $X2=1.43 $Y2=3.33
r42 13 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.43 $Y=3.245
+ $X2=1.43 $Y2=2.9
r43 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.305 $Y=2.19
+ $X2=0.305 $Y2=2.9
r44 7 33 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.235 $Y2=3.33
r45 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.305 $Y2=2.9
r46 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.29
+ $Y=2.045 $X2=1.43 $Y2=2.9
r47 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.29
+ $Y=2.045 $X2=1.43 $Y2=2.19
r48 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.045 $X2=0.305 $Y2=2.9
r49 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.045 $X2=0.305 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0N_LP2%X 1 2 9 12 13 14 15 16 17 42
r21 42 43 3.50689 $w=4.78e-07 $l=1e-08 $layer=LI1_cond $X=2.035 $Y=2.035
+ $X2=2.035 $Y2=2.025
r22 33 46 1.86887 $w=4.78e-07 $l=7.5e-08 $layer=LI1_cond $X=2.035 $Y=2.265
+ $X2=2.035 $Y2=2.19
r23 17 39 3.11479 $w=4.78e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=2.775
+ $X2=2.035 $Y2=2.9
r24 16 17 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.035 $Y=2.405
+ $X2=2.035 $Y2=2.775
r25 16 33 3.48856 $w=4.78e-07 $l=1.4e-07 $layer=LI1_cond $X=2.035 $Y=2.405
+ $X2=2.035 $Y2=2.265
r26 15 46 2.94036 $w=4.78e-07 $l=1.18e-07 $layer=LI1_cond $X=2.035 $Y=2.072
+ $X2=2.035 $Y2=2.19
r27 15 42 0.921977 $w=4.78e-07 $l=3.7e-08 $layer=LI1_cond $X=2.035 $Y=2.072
+ $X2=2.035 $Y2=2.035
r28 15 43 1.90404 $w=2.28e-07 $l=3.8e-08 $layer=LI1_cond $X=2.16 $Y=1.987
+ $X2=2.16 $Y2=2.025
r29 14 15 16.1342 $w=2.28e-07 $l=3.22e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.987
r30 13 14 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.665
r31 12 13 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=1.295
r32 11 12 8.01699 $w=2.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=0.765
+ $X2=2.16 $Y2=0.925
r33 9 11 9.10257 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.11 $Y=0.535
+ $X2=2.11 $Y2=0.765
r34 2 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=2.045 $X2=1.96 $Y2=2.19
r35 2 39 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.82
+ $Y=2.045 $X2=1.96 $Y2=2.9
r36 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.97
+ $Y=0.325 $X2=2.11 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0N_LP2%KAGND 1 4 7
c25 4 0 2.72973e-20 $X=1.2 $Y=0.558
r26 4 7 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0.555 $X2=1.2
+ $Y2=0.555
r27 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.15
+ $Y=0.325 $X2=1.29 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__ISO0N_LP2%VGND 1 5 8 15
r18 5 8 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r19 4 8 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r20 4 5 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r21 1 15 5.20833e-05 $w=2.4e-06 $l=1e-09 $layer=MET1_cond $X=1.2 $Y=0.122
+ $X2=1.2 $Y2=0.123
r22 1 5 0.00635417 $w=2.4e-06 $l=1.22e-07 $layer=MET1_cond $X=1.2 $Y=0.122
+ $X2=1.2 $Y2=0
.ends

