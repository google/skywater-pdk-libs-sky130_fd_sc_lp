* NGSPICE file created from sky130_fd_sc_lp__o22ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_341_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=6.678e+11p pd=6.1e+06u as=2.646e+11p ps=2.94e+06u
M1001 VGND A2 a_27_69# VNB nshort w=840000u l=150000u
+  ad=5.208e+11p pd=2.92e+06u as=7.35e+11p ps=6.79e+06u
M1002 a_341_367# A2 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=8.127e+11p ps=3.81e+06u
M1003 Y B1 a_27_69# VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1004 Y B2 a_110_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1005 a_27_69# B2 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_69# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_110_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

