* File: sky130_fd_sc_lp__a221oi_0.pex.spice
* Created: Fri Aug 28 09:53:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221OI_0%C1 3 6 9 11 12 13 14 19
c41 19 0 1.91845e-19 $X=0.615 $Y=1.375
c42 3 0 2.64969e-20 $X=0.5 $Y=0.445
r43 19 21 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.602 $Y=1.375
+ $X2=0.602 $Y2=1.21
r44 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.615
+ $Y=1.375 $X2=0.615 $Y2=1.375
r45 14 22 5.46897 $w=2.9e-07 $l=1.3e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.675 $Y2=1.905
r46 13 22 9.53746 $w=2.88e-07 $l=2.4e-07 $layer=LI1_cond $X=0.675 $Y=1.665
+ $X2=0.675 $Y2=1.905
r47 13 20 11.5244 $w=2.88e-07 $l=2.9e-07 $layer=LI1_cond $X=0.675 $Y=1.665
+ $X2=0.675 $Y2=1.375
r48 12 20 3.17915 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=0.675 $Y=1.295
+ $X2=0.675 $Y2=1.375
r49 9 11 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=0.705 $Y=2.755
+ $X2=0.705 $Y2=1.88
r50 6 11 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.602 $Y=1.703
+ $X2=0.602 $Y2=1.88
r51 5 19 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.602 $Y=1.387
+ $X2=0.602 $Y2=1.375
r52 5 6 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.602 $Y=1.387
+ $X2=0.602 $Y2=1.703
r53 3 21 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.5 $Y=0.445 $X2=0.5
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_0%B2 3 7 11 12 13 14 19 21 29
c56 21 0 3.57768e-19 $X=1.182 $Y=1.377
c57 19 0 1.62018e-19 $X=1.155 $Y=1.5
c58 7 0 1.93782e-19 $X=1.135 $Y=2.755
r59 21 29 2.59844 $w=3.85e-07 $l=8.2e-08 $layer=LI1_cond $X=1.182 $Y=1.377
+ $X2=1.182 $Y2=1.295
r60 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.155
+ $Y=1.5 $X2=1.155 $Y2=1.5
r61 14 20 4.93904 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.182 $Y=1.665
+ $X2=1.182 $Y2=1.5
r62 13 29 0.0637076 $w=3.83e-07 $l=2e-09 $layer=LI1_cond $X=1.182 $Y=1.293
+ $X2=1.182 $Y2=1.295
r63 13 20 3.6519 $w=3.83e-07 $l=1.22e-07 $layer=LI1_cond $X=1.182 $Y=1.378
+ $X2=1.182 $Y2=1.5
r64 13 21 0.0299336 $w=3.83e-07 $l=1e-09 $layer=LI1_cond $X=1.182 $Y=1.378
+ $X2=1.182 $Y2=1.377
r65 11 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.155 $Y=1.84
+ $X2=1.155 $Y2=1.5
r66 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.84
+ $X2=1.155 $Y2=2.005
r67 10 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.335
+ $X2=1.155 $Y2=1.5
r68 7 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.135 $Y=2.755
+ $X2=1.135 $Y2=2.005
r69 3 10 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.065 $Y=0.445
+ $X2=1.065 $Y2=1.335
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_0%B1 3 4 6 8 11 14 15 17 18 20 21 22 23 31 33
+ 35
r58 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=0.93
+ $X2=1.515 $Y2=0.765
r59 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.515
+ $Y=0.93 $X2=1.515 $Y2=0.93
r60 23 35 5.10519 $w=2.35e-07 $l=2.27e-07 $layer=LI1_cond $X=2.977 $Y=0.897
+ $X2=2.75 $Y2=0.897
r61 22 35 5.39441 $w=2.33e-07 $l=1.1e-07 $layer=LI1_cond $X=2.64 $Y=0.897
+ $X2=2.75 $Y2=0.897
r62 21 22 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0.897
+ $X2=2.64 $Y2=0.897
r63 20 21 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.897
+ $X2=2.16 $Y2=0.897
r64 20 32 8.09162 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=0.897
+ $X2=1.515 $Y2=0.897
r65 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.975
+ $Y=1.53 $X2=2.975 $Y2=1.53
r66 15 23 2.6538 $w=4.55e-07 $l=1.18e-07 $layer=LI1_cond $X=2.977 $Y=1.015
+ $X2=2.977 $Y2=0.897
r67 15 17 13.538 $w=4.53e-07 $l=5.15e-07 $layer=LI1_cond $X=2.977 $Y=1.015
+ $X2=2.977 $Y2=1.53
r68 13 18 54.4068 $w=3.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.965 $Y=1.86
+ $X2=2.965 $Y2=1.53
r69 13 14 48.0802 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.965 $Y=1.86
+ $X2=2.965 $Y2=2.035
r70 9 11 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.695 $Y=2.275
+ $X2=2.865 $Y2=2.275
r71 8 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=2.2
+ $X2=2.865 $Y2=2.275
r72 8 14 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=2.2
+ $X2=2.865 $Y2=2.035
r73 4 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.695 $Y=2.35
+ $X2=2.695 $Y2=2.275
r74 4 6 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.695 $Y=2.35
+ $X2=2.695 $Y2=2.755
r75 3 33 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.455 $Y=0.445
+ $X2=1.455 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_0%A1 3 7 11 13 14 15 19
c50 14 0 1.06357e-19 $X=1.68 $Y=1.295
c51 11 0 1.39426e-19 $X=1.802 $Y=1.485
r52 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73 $Y=1.5
+ $X2=1.73 $Y2=1.5
r53 15 20 5.43295 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.72 $Y2=1.5
r54 14 20 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.72 $Y=1.295
+ $X2=1.72 $Y2=1.5
r55 12 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.73 $Y=1.84
+ $X2=1.73 $Y2=1.5
r56 12 13 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.84
+ $X2=1.73 $Y2=2.005
r57 11 19 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.73 $Y=1.485
+ $X2=1.73 $Y2=1.5
r58 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.802 $Y=1.335
+ $X2=1.802 $Y2=1.485
r59 7 10 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.965 $Y=0.445
+ $X2=1.965 $Y2=1.335
r60 3 13 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.695 $Y=2.755
+ $X2=1.695 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_0%A2 3 5 9 11 12 19 21
c43 9 0 1.06357e-19 $X=2.355 $Y=0.445
c44 3 0 1.86641e-19 $X=2.195 $Y=2.755
r45 19 22 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.825
+ $X2=2.35 $Y2=1.99
r46 19 21 20.2458 $w=4.6e-07 $l=1.3e-07 $layer=POLY_cond $X=2.35 $Y=1.825
+ $X2=2.35 $Y2=1.695
r47 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.825 $X2=2.415 $Y2=1.825
r48 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.485 $X2=2.415 $Y2=1.485
r49 12 20 3.71597 $w=5.13e-07 $l=1.6e-07 $layer=LI1_cond $X=2.322 $Y=1.665
+ $X2=2.322 $Y2=1.825
r50 12 17 4.18047 $w=5.13e-07 $l=1.8e-07 $layer=LI1_cond $X=2.322 $Y=1.665
+ $X2=2.322 $Y2=1.485
r51 11 17 4.41272 $w=5.13e-07 $l=1.9e-07 $layer=LI1_cond $X=2.322 $Y=1.295
+ $X2=2.322 $Y2=1.485
r52 7 16 38.5818 $w=3.27e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.355 $Y=1.32
+ $X2=2.415 $Y2=1.485
r53 7 9 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=2.355 $Y=1.32
+ $X2=2.355 $Y2=0.445
r54 5 16 2.19091 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.415 $Y=1.5
+ $X2=2.415 $Y2=1.485
r55 5 21 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.415 $Y=1.5
+ $X2=2.415 $Y2=1.695
r56 3 22 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.195 $Y=2.755
+ $X2=2.195 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_0%Y 1 2 3 12 15 16 18 20 21 22 23 24 25 26 27
+ 48
c50 25 0 1.93782e-19 $X=0.155 $Y=2.32
c51 20 0 1.62018e-19 $X=1 $Y=0.895
r52 48 55 0.54102 $w=2.03e-07 $l=1e-08 $layer=LI1_cond $X=0.257 $Y=2.405
+ $X2=0.257 $Y2=2.415
r53 27 49 16.5351 $w=2.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.72 $Y=0.895
+ $X2=0.39 $Y2=0.895
r54 26 57 4.66471 $w=4.98e-07 $l=1.95e-07 $layer=LI1_cond $X=0.405 $Y=2.775
+ $X2=0.405 $Y2=2.58
r55 25 57 3.06196 $w=4.98e-07 $l=1.28e-07 $layer=LI1_cond $X=0.405 $Y=2.452
+ $X2=0.405 $Y2=2.58
r56 25 55 5.16693 $w=4.98e-07 $l=3.7e-08 $layer=LI1_cond $X=0.405 $Y=2.452
+ $X2=0.405 $Y2=2.415
r57 25 48 2.05588 $w=2.03e-07 $l=3.8e-08 $layer=LI1_cond $X=0.257 $Y=2.367
+ $X2=0.257 $Y2=2.405
r58 24 25 17.9619 $w=2.03e-07 $l=3.32e-07 $layer=LI1_cond $X=0.257 $Y=2.035
+ $X2=0.257 $Y2=2.367
r59 23 24 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=2.035
r60 22 23 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.295
+ $X2=0.257 $Y2=1.665
r61 21 49 1.18299 $w=2.3e-07 $l=1.18e-07 $layer=LI1_cond $X=0.272 $Y=0.895
+ $X2=0.39 $Y2=0.895
r62 21 22 11.11 $w=3.73e-07 $l=2.85e-07 $layer=LI1_cond $X=0.257 $Y=1.01
+ $X2=0.257 $Y2=1.295
r63 20 27 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=0.895 $X2=0.72
+ $Y2=0.895
r64 16 18 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=1.17 $Y=0.445
+ $X2=1.715 $Y2=0.445
r65 15 20 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.085 $Y=0.78
+ $X2=1 $Y2=0.895
r66 14 16 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.085 $Y=0.61
+ $X2=1.17 $Y2=0.445
r67 14 15 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.085 $Y=0.61
+ $X2=1.085 $Y2=0.78
r68 10 21 5.35987 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=0.272 $Y=0.78
+ $X2=0.272 $Y2=0.895
r69 10 12 16.4284 $w=2.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.272 $Y=0.78
+ $X2=0.272 $Y2=0.445
r70 3 57 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.365
+ $Y=2.435 $X2=0.49 $Y2=2.58
r71 2 18 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.235 $X2=1.715 $Y2=0.445
r72 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_0%A_156_487# 1 2 7 9 11 15
c36 15 0 1.86641e-19 $X=2.98 $Y=2.58
r37 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.98 $Y=2.305
+ $X2=2.98 $Y2=2.58
r38 12 17 2.80567 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.145 $Y=2.22
+ $X2=0.985 $Y2=2.22
r39 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.815 $Y=2.22
+ $X2=2.98 $Y2=2.305
r40 11 12 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=2.815 $Y=2.22
+ $X2=1.145 $Y2=2.22
r41 7 17 10.0942 $w=3.2e-07 $l=2.45e-07 $layer=LI1_cond $X=0.985 $Y=2.465
+ $X2=0.985 $Y2=2.22
r42 7 9 3.42132 $w=3.18e-07 $l=9.5e-08 $layer=LI1_cond $X=0.985 $Y=2.465
+ $X2=0.985 $Y2=2.56
r43 2 15 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=2.77
+ $Y=2.435 $X2=2.98 $Y2=2.58
r44 1 9 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=0.78
+ $Y=2.435 $X2=0.92 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_0%A_242_487# 1 2 9 14 16
r21 10 14 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=2.565
+ $X2=1.48 $Y2=2.565
r22 9 16 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=2.565
+ $X2=2.48 $Y2=2.565
r23 9 10 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.315 $Y=2.565
+ $X2=1.645 $Y2=2.565
r24 2 16 300 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.435 $X2=2.48 $Y2=2.59
r25 1 14 300 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_PDIFF $count=2 $X=1.21
+ $Y=2.435 $X2=1.48 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_0%VPWR 1 6 9 10 11 24 25
r34 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 22 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 21 24 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r37 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 14 18 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 11 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 11 15 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 11 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 9 18 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.98 $Y2=3.33
r45 8 21 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=1.98 $Y2=3.33
r47 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=3.245 $X2=1.98
+ $Y2=3.33
r48 4 6 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.98 $Y=3.245 $X2=1.98
+ $Y2=2.925
r49 1 6 600 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=2.435 $X2=1.98 $Y2=2.925
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_0%VGND 1 2 9 13 15 17 22 32 33 36 39
r39 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r42 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.57
+ $Y2=0
r44 30 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=3.12
+ $Y2=0
r45 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r46 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r47 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r49 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 23 36 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.72
+ $Y2=0
r51 23 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.2
+ $Y2=0
r52 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.57
+ $Y2=0
r53 22 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.16
+ $Y2=0
r54 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r55 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r56 17 36 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.72
+ $Y2=0
r57 17 19 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.24
+ $Y2=0
r58 15 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r59 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r60 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=0.085
+ $X2=2.57 $Y2=0
r61 11 13 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.57 $Y=0.085
+ $X2=2.57 $Y2=0.445
r62 7 36 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r63 7 9 18.8582 $w=2.18e-07 $l=3.6e-07 $layer=LI1_cond $X=0.72 $Y=0.085 $X2=0.72
+ $Y2=0.445
r64 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.235 $X2=2.57 $Y2=0.445
r65 1 9 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.745 $Y2=0.445
.ends

