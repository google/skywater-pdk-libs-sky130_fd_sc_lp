* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfxbp_2 CLK D VGND VNB VPB VPWR Q Q_N
X0 VGND a_1513_137# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_537_119# a_110_70# a_669_499# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND CLK a_110_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_236_463# a_110_70# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 Q a_1169_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_670_93# a_236_463# a_982_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1157_453# a_1169_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND a_1169_93# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_429_119# a_236_463# a_537_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 Q_N a_1513_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND a_537_119# a_670_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_537_119# a_236_463# a_628_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_1169_93# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VPWR a_537_119# a_670_93# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 a_982_369# a_236_463# a_1157_453# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_429_119# a_110_70# a_537_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_982_369# a_110_70# a_1125_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_982_369# a_1169_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_1513_137# a_1169_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_236_463# a_110_70# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_982_369# a_1169_93# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 Q a_1169_93# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_1513_137# a_1169_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_670_93# a_110_70# a_982_369# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X24 a_628_119# a_670_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VPWR CLK a_110_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 VGND D a_429_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 Q_N a_1513_137# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_669_499# a_670_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VPWR a_1513_137# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 VPWR D a_429_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_1125_119# a_1169_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
