* File: sky130_fd_sc_lp__and2b_lp.pxi.spice
* Created: Wed Sep  2 09:31:14 2020
* 
x_PM_SKY130_FD_SC_LP__AND2B_LP%A_108_127# N_A_108_127#_M1004_d
+ N_A_108_127#_M1000_d N_A_108_127#_c_53_n N_A_108_127#_M1006_g
+ N_A_108_127#_M1008_g N_A_108_127#_c_55_n N_A_108_127#_M1003_g
+ N_A_108_127#_c_56_n N_A_108_127#_c_57_n N_A_108_127#_c_58_n
+ N_A_108_127#_c_65_p N_A_108_127#_c_99_p N_A_108_127#_c_59_n
+ N_A_108_127#_c_66_p N_A_108_127#_c_60_n
+ PM_SKY130_FD_SC_LP__AND2B_LP%A_108_127#
x_PM_SKY130_FD_SC_LP__AND2B_LP%B N_B_M1000_g N_B_M1001_g B N_B_c_123_n
+ N_B_c_124_n PM_SKY130_FD_SC_LP__AND2B_LP%B
x_PM_SKY130_FD_SC_LP__AND2B_LP%A_378_159# N_A_378_159#_M1007_d
+ N_A_378_159#_M1002_d N_A_378_159#_M1004_g N_A_378_159#_M1009_g
+ N_A_378_159#_c_162_n N_A_378_159#_c_163_n N_A_378_159#_c_170_n
+ N_A_378_159#_c_164_n N_A_378_159#_c_165_n N_A_378_159#_c_166_n
+ PM_SKY130_FD_SC_LP__AND2B_LP%A_378_159#
x_PM_SKY130_FD_SC_LP__AND2B_LP%A_N N_A_N_M1005_g N_A_N_M1002_g N_A_N_M1007_g A_N
+ N_A_N_c_216_n N_A_N_c_217_n PM_SKY130_FD_SC_LP__AND2B_LP%A_N
x_PM_SKY130_FD_SC_LP__AND2B_LP%X N_X_M1006_s N_X_M1008_s X X X X X X X
+ PM_SKY130_FD_SC_LP__AND2B_LP%X
x_PM_SKY130_FD_SC_LP__AND2B_LP%VPWR N_VPWR_M1008_d N_VPWR_M1009_d N_VPWR_c_264_n
+ N_VPWR_c_265_n N_VPWR_c_266_n N_VPWR_c_267_n VPWR N_VPWR_c_268_n
+ N_VPWR_c_269_n N_VPWR_c_263_n N_VPWR_c_271_n PM_SKY130_FD_SC_LP__AND2B_LP%VPWR
x_PM_SKY130_FD_SC_LP__AND2B_LP%VGND N_VGND_M1003_d N_VGND_M1005_s N_VGND_c_307_n
+ N_VGND_c_308_n N_VGND_c_309_n VGND N_VGND_c_310_n N_VGND_c_311_n
+ N_VGND_c_312_n N_VGND_c_313_n N_VGND_c_314_n PM_SKY130_FD_SC_LP__AND2B_LP%VGND
cc_1 VNB N_A_108_127#_c_53_n 0.0193148f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_2 VNB N_A_108_127#_M1008_g 0.00196579f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.595
cc_3 VNB N_A_108_127#_c_55_n 0.0164459f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.295
cc_4 VNB N_A_108_127#_c_56_n 2.1104e-19 $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.46
cc_5 VNB N_A_108_127#_c_57_n 0.024045f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=1.34
cc_6 VNB N_A_108_127#_c_58_n 0.00757196f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.34
cc_7 VNB N_A_108_127#_c_59_n 0.00769864f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=1.135
cc_8 VNB N_A_108_127#_c_60_n 0.0461199f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.46
cc_9 VNB N_B_M1001_g 0.0375725f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_10 VNB N_B_c_123_n 0.0106801f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.595
cc_11 VNB N_B_c_124_n 0.00355824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_378_159#_M1004_g 0.0291412f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.975
cc_13 VNB N_A_378_159#_c_162_n 0.00393603f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.975
cc_14 VNB N_A_378_159#_c_163_n 0.0125076f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.33
cc_15 VNB N_A_378_159#_c_164_n 0.0448385f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=2.415
cc_16 VNB N_A_378_159#_c_165_n 0.00945573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_378_159#_c_166_n 0.0197773f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=1.255
cc_18 VNB N_A_N_M1005_g 0.0356142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_N_M1002_g 0.0232257f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_20 VNB N_A_N_M1007_g 0.0347471f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.595
cc_21 VNB N_A_N_c_216_n 0.00381974f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.46
cc_22 VNB N_A_N_c_217_n 0.0442528f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.46
cc_23 VNB X 0.0634061f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.295
cc_24 VNB N_VPWR_c_263_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_307_n 0.0358815f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.975
cc_26 VNB N_VGND_c_308_n 0.02253f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.595
cc_27 VNB N_VGND_c_309_n 0.0233443f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.975
cc_28 VNB N_VGND_c_310_n 0.0328155f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.46
cc_29 VNB N_VGND_c_311_n 0.0279964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_312_n 0.230946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_313_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.18 $Y2=1.135
cc_32 VNB N_VGND_c_314_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=2.495
cc_33 VPB N_A_108_127#_M1008_g 0.0487024f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.595
cc_34 VPB N_A_108_127#_c_56_n 0.00337807f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.46
cc_35 VPB N_B_M1000_g 0.0258601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_B_c_123_n 0.0201218f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.595
cc_37 VPB N_B_c_124_n 0.00444913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_378_159#_M1009_g 0.0269253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_378_159#_c_162_n 0.00507851f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.975
cc_40 VPB N_A_378_159#_c_163_n 0.0223715f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.33
cc_41 VPB N_A_378_159#_c_170_n 0.0436279f $X=-0.19 $Y=1.655 $X2=2.015 $Y2=1.34
cc_42 VPB N_A_378_159#_c_165_n 0.0201054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_N_M1002_g 0.0499988f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.295
cc_44 VPB X 0.0724483f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.295
cc_45 VPB N_VPWR_c_264_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.975
cc_46 VPB N_VPWR_c_265_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_266_n 0.0240582f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.975
cc_48 VPB N_VPWR_c_267_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.425
cc_49 VPB N_VPWR_c_268_n 0.0256171f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.415
cc_50 VPB N_VPWR_c_269_n 0.0282344f $X=-0.19 $Y=1.655 $X2=2.18 $Y2=1.135
cc_51 VPB N_VPWR_c_263_n 0.0541667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_271_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.46
cc_53 N_A_108_127#_M1008_g N_B_M1000_g 0.0242383f $X=0.75 $Y=2.595 $X2=0 $Y2=0
cc_54 N_A_108_127#_c_56_n N_B_M1000_g 0.00493206f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_55 N_A_108_127#_c_65_p N_B_M1000_g 0.0149613f $X=1.585 $Y=2.415 $X2=0 $Y2=0
cc_56 N_A_108_127#_c_66_p N_B_M1000_g 0.0163585f $X=1.75 $Y=2.495 $X2=0 $Y2=0
cc_57 N_A_108_127#_c_55_n N_B_M1001_g 0.0240618f $X=1.005 $Y=1.295 $X2=0 $Y2=0
cc_58 N_A_108_127#_c_56_n N_B_M1001_g 0.00107644f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_59 N_A_108_127#_c_57_n N_B_M1001_g 0.0153453f $X=2.015 $Y=1.34 $X2=0 $Y2=0
cc_60 N_A_108_127#_c_59_n N_B_M1001_g 0.00138391f $X=2.18 $Y=1.135 $X2=0 $Y2=0
cc_61 N_A_108_127#_M1008_g N_B_c_123_n 0.00693037f $X=0.75 $Y=2.595 $X2=0 $Y2=0
cc_62 N_A_108_127#_c_56_n N_B_c_123_n 0.00264599f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_63 N_A_108_127#_c_57_n N_B_c_123_n 0.00123714f $X=2.015 $Y=1.34 $X2=0 $Y2=0
cc_64 N_A_108_127#_c_60_n N_B_c_123_n 0.00107535f $X=1.005 $Y=1.46 $X2=0 $Y2=0
cc_65 N_A_108_127#_M1000_d N_B_c_124_n 0.00206558f $X=1.61 $Y=2.095 $X2=0 $Y2=0
cc_66 N_A_108_127#_M1008_g N_B_c_124_n 8.01838e-19 $X=0.75 $Y=2.595 $X2=0 $Y2=0
cc_67 N_A_108_127#_c_56_n N_B_c_124_n 0.0330933f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_68 N_A_108_127#_c_57_n N_B_c_124_n 0.0356373f $X=2.015 $Y=1.34 $X2=0 $Y2=0
cc_69 N_A_108_127#_c_65_p N_B_c_124_n 0.0160348f $X=1.585 $Y=2.415 $X2=0 $Y2=0
cc_70 N_A_108_127#_c_66_p N_B_c_124_n 0.0127378f $X=1.75 $Y=2.495 $X2=0 $Y2=0
cc_71 N_A_108_127#_c_57_n N_A_378_159#_M1004_g 0.0156801f $X=2.015 $Y=1.34 $X2=0
+ $Y2=0
cc_72 N_A_108_127#_c_59_n N_A_378_159#_M1004_g 0.00812896f $X=2.18 $Y=1.135
+ $X2=0 $Y2=0
cc_73 N_A_108_127#_c_66_p N_A_378_159#_M1009_g 0.0142146f $X=1.75 $Y=2.495 $X2=0
+ $Y2=0
cc_74 N_A_108_127#_c_57_n N_A_378_159#_c_162_n 0.0288298f $X=2.015 $Y=1.34 $X2=0
+ $Y2=0
cc_75 N_A_108_127#_c_57_n N_A_378_159#_c_163_n 0.00647338f $X=2.015 $Y=1.34
+ $X2=0 $Y2=0
cc_76 N_A_108_127#_c_59_n N_A_N_M1005_g 0.00593991f $X=2.18 $Y=1.135 $X2=0 $Y2=0
cc_77 N_A_108_127#_c_57_n N_A_N_M1002_g 6.38942e-19 $X=2.015 $Y=1.34 $X2=0 $Y2=0
cc_78 N_A_108_127#_c_57_n N_A_N_c_216_n 0.012706f $X=2.015 $Y=1.34 $X2=0 $Y2=0
cc_79 N_A_108_127#_c_59_n N_A_N_c_216_n 0.0166362f $X=2.18 $Y=1.135 $X2=0 $Y2=0
cc_80 N_A_108_127#_c_57_n N_A_N_c_217_n 0.00121981f $X=2.015 $Y=1.34 $X2=0 $Y2=0
cc_81 N_A_108_127#_c_53_n X 0.0175525f $X=0.615 $Y=1.295 $X2=0 $Y2=0
cc_82 N_A_108_127#_M1008_g X 0.0176179f $X=0.75 $Y=2.595 $X2=0 $Y2=0
cc_83 N_A_108_127#_c_55_n X 0.00218011f $X=1.005 $Y=1.295 $X2=0 $Y2=0
cc_84 N_A_108_127#_c_56_n X 0.0594398f $X=0.915 $Y=1.46 $X2=0 $Y2=0
cc_85 N_A_108_127#_c_58_n X 0.013389f $X=1.08 $Y=1.34 $X2=0 $Y2=0
cc_86 N_A_108_127#_c_60_n X 0.0136219f $X=1.005 $Y=1.46 $X2=0 $Y2=0
cc_87 N_A_108_127#_c_56_n N_VPWR_M1008_d 0.00332407f $X=0.915 $Y=1.46 $X2=-0.19
+ $Y2=-0.245
cc_88 N_A_108_127#_c_65_p N_VPWR_M1008_d 0.0129141f $X=1.585 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_89 N_A_108_127#_c_99_p N_VPWR_M1008_d 0.00187712f $X=1.08 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_90 N_A_108_127#_M1008_g N_VPWR_c_264_n 0.0132094f $X=0.75 $Y=2.595 $X2=0
+ $Y2=0
cc_91 N_A_108_127#_c_65_p N_VPWR_c_264_n 0.00747743f $X=1.585 $Y=2.415 $X2=0
+ $Y2=0
cc_92 N_A_108_127#_c_99_p N_VPWR_c_264_n 0.0142457f $X=1.08 $Y=2.415 $X2=0 $Y2=0
cc_93 N_A_108_127#_c_66_p N_VPWR_c_264_n 0.0153132f $X=1.75 $Y=2.495 $X2=0 $Y2=0
cc_94 N_A_108_127#_c_66_p N_VPWR_c_265_n 0.0491014f $X=1.75 $Y=2.495 $X2=0 $Y2=0
cc_95 N_A_108_127#_M1008_g N_VPWR_c_266_n 0.008763f $X=0.75 $Y=2.595 $X2=0 $Y2=0
cc_96 N_A_108_127#_c_66_p N_VPWR_c_268_n 0.0177952f $X=1.75 $Y=2.495 $X2=0 $Y2=0
cc_97 N_A_108_127#_M1000_d N_VPWR_c_263_n 0.00223819f $X=1.61 $Y=2.095 $X2=0
+ $Y2=0
cc_98 N_A_108_127#_M1008_g N_VPWR_c_263_n 0.0124997f $X=0.75 $Y=2.595 $X2=0
+ $Y2=0
cc_99 N_A_108_127#_c_65_p N_VPWR_c_263_n 0.0128532f $X=1.585 $Y=2.415 $X2=0
+ $Y2=0
cc_100 N_A_108_127#_c_99_p N_VPWR_c_263_n 0.00408f $X=1.08 $Y=2.415 $X2=0 $Y2=0
cc_101 N_A_108_127#_c_66_p N_VPWR_c_263_n 0.0123247f $X=1.75 $Y=2.495 $X2=0
+ $Y2=0
cc_102 N_A_108_127#_c_53_n N_VGND_c_307_n 0.00124234f $X=0.615 $Y=1.295 $X2=0
+ $Y2=0
cc_103 N_A_108_127#_c_55_n N_VGND_c_307_n 0.00972358f $X=1.005 $Y=1.295 $X2=0
+ $Y2=0
cc_104 N_A_108_127#_c_57_n N_VGND_c_307_n 0.0205044f $X=2.015 $Y=1.34 $X2=0
+ $Y2=0
cc_105 N_A_108_127#_c_58_n N_VGND_c_307_n 0.00189912f $X=1.08 $Y=1.34 $X2=0
+ $Y2=0
cc_106 N_A_108_127#_c_59_n N_VGND_c_309_n 0.0183994f $X=2.18 $Y=1.135 $X2=0
+ $Y2=0
cc_107 N_A_108_127#_c_53_n N_VGND_c_310_n 0.00290919f $X=0.615 $Y=1.295 $X2=0
+ $Y2=0
cc_108 N_A_108_127#_c_55_n N_VGND_c_310_n 0.00289826f $X=1.005 $Y=1.295 $X2=0
+ $Y2=0
cc_109 N_A_108_127#_c_53_n N_VGND_c_312_n 0.0034881f $X=0.615 $Y=1.295 $X2=0
+ $Y2=0
cc_110 N_A_108_127#_c_55_n N_VGND_c_312_n 0.00363223f $X=1.005 $Y=1.295 $X2=0
+ $Y2=0
cc_111 N_A_108_127#_c_57_n A_313_153# 0.00736402f $X=2.015 $Y=1.34 $X2=-0.19
+ $Y2=-0.245
cc_112 N_B_M1001_g N_A_378_159#_M1004_g 0.0315204f $X=1.49 $Y=0.975 $X2=0 $Y2=0
cc_113 N_B_M1000_g N_A_378_159#_M1009_g 0.0237813f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_114 N_B_c_123_n N_A_378_159#_c_162_n 2.79725e-19 $X=1.485 $Y=1.77 $X2=0 $Y2=0
cc_115 N_B_c_124_n N_A_378_159#_c_162_n 0.027098f $X=1.485 $Y=1.77 $X2=0 $Y2=0
cc_116 N_B_c_123_n N_A_378_159#_c_163_n 0.0174906f $X=1.485 $Y=1.77 $X2=0 $Y2=0
cc_117 N_B_c_124_n N_A_378_159#_c_163_n 0.00798638f $X=1.485 $Y=1.77 $X2=0 $Y2=0
cc_118 N_B_M1000_g N_VPWR_c_264_n 0.00754036f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_119 N_B_M1000_g N_VPWR_c_265_n 0.00186723f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_120 N_B_c_124_n N_VPWR_c_265_n 0.00172177f $X=1.485 $Y=1.77 $X2=0 $Y2=0
cc_121 N_B_M1000_g N_VPWR_c_268_n 0.00939541f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_122 N_B_M1000_g N_VPWR_c_263_n 0.0099576f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_123 N_B_M1001_g N_VGND_c_307_n 0.00370971f $X=1.49 $Y=0.975 $X2=0 $Y2=0
cc_124 N_B_M1001_g N_VGND_c_308_n 0.00348629f $X=1.49 $Y=0.975 $X2=0 $Y2=0
cc_125 N_B_M1001_g N_VGND_c_309_n 0.00101844f $X=1.49 $Y=0.975 $X2=0 $Y2=0
cc_126 N_B_M1001_g N_VGND_c_312_n 0.00432409f $X=1.49 $Y=0.975 $X2=0 $Y2=0
cc_127 N_A_378_159#_M1004_g N_A_N_M1005_g 0.0119659f $X=1.965 $Y=1.135 $X2=0
+ $Y2=0
cc_128 N_A_378_159#_c_166_n N_A_N_M1005_g 0.0010756f $X=3.08 $Y=0.445 $X2=0
+ $Y2=0
cc_129 N_A_378_159#_M1004_g N_A_N_M1002_g 0.00664675f $X=1.965 $Y=1.135 $X2=0
+ $Y2=0
cc_130 N_A_378_159#_M1009_g N_A_N_M1002_g 0.0245063f $X=2.015 $Y=2.595 $X2=0
+ $Y2=0
cc_131 N_A_378_159#_c_162_n N_A_N_M1002_g 0.0243616f $X=2.77 $Y=1.77 $X2=0 $Y2=0
cc_132 N_A_378_159#_c_163_n N_A_N_M1002_g 0.018168f $X=2.14 $Y=1.77 $X2=0 $Y2=0
cc_133 N_A_378_159#_c_170_n N_A_N_M1002_g 0.0283345f $X=2.935 $Y=2.24 $X2=0
+ $Y2=0
cc_134 N_A_378_159#_c_164_n N_A_N_M1002_g 0.00494093f $X=3.16 $Y=1.605 $X2=0
+ $Y2=0
cc_135 N_A_378_159#_c_165_n N_A_N_M1002_g 0.00844008f $X=3.007 $Y=1.77 $X2=0
+ $Y2=0
cc_136 N_A_378_159#_c_164_n N_A_N_M1007_g 0.0197461f $X=3.16 $Y=1.605 $X2=0
+ $Y2=0
cc_137 N_A_378_159#_c_166_n N_A_N_M1007_g 0.00841368f $X=3.08 $Y=0.445 $X2=0
+ $Y2=0
cc_138 N_A_378_159#_c_162_n N_A_N_c_216_n 0.0167695f $X=2.77 $Y=1.77 $X2=0 $Y2=0
cc_139 N_A_378_159#_c_164_n N_A_N_c_216_n 0.0234184f $X=3.16 $Y=1.605 $X2=0
+ $Y2=0
cc_140 N_A_378_159#_c_165_n N_A_N_c_216_n 0.00661051f $X=3.007 $Y=1.77 $X2=0
+ $Y2=0
cc_141 N_A_378_159#_c_162_n N_A_N_c_217_n 0.0053064f $X=2.77 $Y=1.77 $X2=0 $Y2=0
cc_142 N_A_378_159#_c_165_n N_A_N_c_217_n 0.00426553f $X=3.007 $Y=1.77 $X2=0
+ $Y2=0
cc_143 N_A_378_159#_M1009_g N_VPWR_c_265_n 0.0262782f $X=2.015 $Y=2.595 $X2=0
+ $Y2=0
cc_144 N_A_378_159#_c_162_n N_VPWR_c_265_n 0.0239317f $X=2.77 $Y=1.77 $X2=0
+ $Y2=0
cc_145 N_A_378_159#_c_163_n N_VPWR_c_265_n 0.0036453f $X=2.14 $Y=1.77 $X2=0
+ $Y2=0
cc_146 N_A_378_159#_c_170_n N_VPWR_c_265_n 0.0448599f $X=2.935 $Y=2.24 $X2=0
+ $Y2=0
cc_147 N_A_378_159#_M1009_g N_VPWR_c_268_n 0.00840199f $X=2.015 $Y=2.595 $X2=0
+ $Y2=0
cc_148 N_A_378_159#_c_170_n N_VPWR_c_269_n 0.019758f $X=2.935 $Y=2.24 $X2=0
+ $Y2=0
cc_149 N_A_378_159#_M1002_d N_VPWR_c_263_n 0.0023218f $X=2.795 $Y=2.095 $X2=0
+ $Y2=0
cc_150 N_A_378_159#_M1009_g N_VPWR_c_263_n 0.0136033f $X=2.015 $Y=2.595 $X2=0
+ $Y2=0
cc_151 N_A_378_159#_c_170_n N_VPWR_c_263_n 0.012508f $X=2.935 $Y=2.24 $X2=0
+ $Y2=0
cc_152 N_A_378_159#_c_166_n N_VGND_c_309_n 0.0120387f $X=3.08 $Y=0.445 $X2=0
+ $Y2=0
cc_153 N_A_378_159#_c_166_n N_VGND_c_311_n 0.0165089f $X=3.08 $Y=0.445 $X2=0
+ $Y2=0
cc_154 N_A_378_159#_M1007_d N_VGND_c_312_n 0.00234843f $X=2.94 $Y=0.235 $X2=0
+ $Y2=0
cc_155 N_A_378_159#_M1004_g N_VGND_c_312_n 0.00393927f $X=1.965 $Y=1.135 $X2=0
+ $Y2=0
cc_156 N_A_378_159#_c_166_n N_VGND_c_312_n 0.0122765f $X=3.08 $Y=0.445 $X2=0
+ $Y2=0
cc_157 N_A_N_M1002_g N_VPWR_c_265_n 0.0141887f $X=2.67 $Y=2.595 $X2=0 $Y2=0
cc_158 N_A_N_M1002_g N_VPWR_c_269_n 0.00939541f $X=2.67 $Y=2.595 $X2=0 $Y2=0
cc_159 N_A_N_M1002_g N_VPWR_c_263_n 0.0175815f $X=2.67 $Y=2.595 $X2=0 $Y2=0
cc_160 N_A_N_M1005_g N_VGND_c_309_n 0.0155215f $X=2.475 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_N_M1007_g N_VGND_c_309_n 0.0024608f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_N_M1005_g N_VGND_c_311_n 0.00486043f $X=2.475 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_N_M1007_g N_VGND_c_311_n 0.00550269f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A_N_M1005_g N_VGND_c_312_n 0.00823808f $X=2.475 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_N_M1007_g N_VGND_c_312_n 0.0110006f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_166 X N_VPWR_c_266_n 0.0295251f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_167 N_X_M1008_s N_VPWR_c_263_n 0.0042346f $X=0.34 $Y=2.095 $X2=0 $Y2=0
cc_168 X N_VPWR_c_263_n 0.0171356f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_169 X N_VGND_c_307_n 0.02244f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_170 X N_VGND_c_310_n 0.0144859f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_171 X N_VGND_c_312_n 0.0154459f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_172 N_VGND_c_312_n A_510_47# 0.010279f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
