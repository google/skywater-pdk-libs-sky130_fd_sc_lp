* File: sky130_fd_sc_lp__a21bo_m.pxi.spice
* Created: Wed Sep  2 09:19:05 2020
* 
x_PM_SKY130_FD_SC_LP__A21BO_M%A_80_72# N_A_80_72#_M1000_d N_A_80_72#_M1003_s
+ N_A_80_72#_M1002_g N_A_80_72#_c_87_n N_A_80_72#_M1008_g N_A_80_72#_c_89_n
+ N_A_80_72#_c_82_n N_A_80_72#_c_83_n N_A_80_72#_c_91_n N_A_80_72#_c_92_n
+ N_A_80_72#_c_93_n N_A_80_72#_c_84_n N_A_80_72#_c_85_n N_A_80_72#_c_131_p
+ N_A_80_72#_c_86_n PM_SKY130_FD_SC_LP__A21BO_M%A_80_72#
x_PM_SKY130_FD_SC_LP__A21BO_M%B1_N N_B1_N_c_175_n N_B1_N_M1006_g N_B1_N_c_180_n
+ N_B1_N_M1001_g N_B1_N_c_181_n N_B1_N_c_176_n N_B1_N_c_182_n N_B1_N_c_177_n
+ B1_N B1_N B1_N N_B1_N_c_178_n N_B1_N_c_179_n PM_SKY130_FD_SC_LP__A21BO_M%B1_N
x_PM_SKY130_FD_SC_LP__A21BO_M%A_196_98# N_A_196_98#_M1006_d N_A_196_98#_M1001_d
+ N_A_196_98#_c_232_n N_A_196_98#_c_233_n N_A_196_98#_c_240_n
+ N_A_196_98#_c_241_n N_A_196_98#_M1000_g N_A_196_98#_c_242_n
+ N_A_196_98#_M1003_g N_A_196_98#_c_234_n N_A_196_98#_c_243_n
+ N_A_196_98#_c_244_n N_A_196_98#_c_235_n N_A_196_98#_c_236_n
+ N_A_196_98#_c_237_n N_A_196_98#_c_275_n N_A_196_98#_c_245_n
+ N_A_196_98#_c_238_n PM_SKY130_FD_SC_LP__A21BO_M%A_196_98#
x_PM_SKY130_FD_SC_LP__A21BO_M%A1 N_A1_M1004_g N_A1_M1009_g N_A1_c_309_n
+ N_A1_c_310_n N_A1_c_311_n A1 A1 N_A1_c_313_n PM_SKY130_FD_SC_LP__A21BO_M%A1
x_PM_SKY130_FD_SC_LP__A21BO_M%A2 N_A2_M1005_g N_A2_M1007_g N_A2_c_353_n
+ N_A2_c_354_n A2 A2 A2 N_A2_c_356_n PM_SKY130_FD_SC_LP__A21BO_M%A2
x_PM_SKY130_FD_SC_LP__A21BO_M%X N_X_M1002_s N_X_M1008_s X X X X X X X
+ PM_SKY130_FD_SC_LP__A21BO_M%X
x_PM_SKY130_FD_SC_LP__A21BO_M%VPWR N_VPWR_M1008_d N_VPWR_M1009_d N_VPWR_c_400_n
+ N_VPWR_c_401_n N_VPWR_c_402_n VPWR N_VPWR_c_403_n N_VPWR_c_404_n
+ N_VPWR_c_399_n N_VPWR_c_406_n N_VPWR_c_407_n PM_SKY130_FD_SC_LP__A21BO_M%VPWR
x_PM_SKY130_FD_SC_LP__A21BO_M%A_419_439# N_A_419_439#_M1003_d
+ N_A_419_439#_M1007_d N_A_419_439#_c_438_n N_A_419_439#_c_439_n
+ N_A_419_439#_c_440_n N_A_419_439#_c_441_n
+ PM_SKY130_FD_SC_LP__A21BO_M%A_419_439#
x_PM_SKY130_FD_SC_LP__A21BO_M%VGND N_VGND_M1002_d N_VGND_M1000_s N_VGND_M1005_d
+ N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n N_VGND_c_461_n
+ N_VGND_c_462_n VGND N_VGND_c_463_n N_VGND_c_464_n N_VGND_c_465_n
+ N_VGND_c_466_n PM_SKY130_FD_SC_LP__A21BO_M%VGND
cc_1 VNB N_A_80_72#_M1002_g 0.0485141f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.7
cc_2 VNB N_A_80_72#_c_82_n 0.00299759f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.64
cc_3 VNB N_A_80_72#_c_83_n 0.0207787f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.64
cc_4 VNB N_A_80_72#_c_84_n 0.0100452f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.71
cc_5 VNB N_A_80_72#_c_85_n 0.00104894f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.71
cc_6 VNB N_A_80_72#_c_86_n 0.0127772f $X=-0.19 $Y=-0.245 $X2=2.71 $Y2=1.625
cc_7 VNB N_B1_N_c_175_n 0.0200585f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=0.235
cc_8 VNB N_B1_N_c_176_n 0.0363536f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.968
cc_9 VNB N_B1_N_c_177_n 0.00916355f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.64
cc_10 VNB N_B1_N_c_178_n 0.0256706f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.71
cc_11 VNB N_B1_N_c_179_n 0.00159713f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.71
cc_12 VNB N_A_196_98#_c_232_n 0.0236272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_196_98#_c_233_n 0.011152f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.968
cc_14 VNB N_A_196_98#_c_234_n 0.0179646f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.42
cc_15 VNB N_A_196_98#_c_235_n 0.0176857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_196_98#_c_236_n 7.49658e-19 $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.34
cc_17 VNB N_A_196_98#_c_237_n 0.0207833f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.64
cc_18 VNB N_A_196_98#_c_238_n 0.0201463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1009_g 0.0152185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_309_n 0.0169629f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.7
cc_21 VNB N_A1_c_310_n 0.0216313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_c_311_n 0.0157762f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.652
cc_23 VNB A1 0.00982101f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.968
cc_24 VNB N_A1_c_313_n 0.0153068f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=2.145
cc_25 VNB N_A2_M1005_g 0.0267554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_M1007_g 0.00804854f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.475
cc_27 VNB N_A2_c_353_n 0.0308374f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.652
cc_28 VNB N_A2_c_354_n 0.0326343f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.145
cc_29 VNB A2 0.00888511f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.855
cc_30 VNB N_A2_c_356_n 0.0358078f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.64
cc_31 VNB X 0.00314671f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.475
cc_32 VNB X 0.0364486f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.7
cc_33 VNB N_VPWR_c_399_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.71
cc_34 VNB N_VGND_c_457_n 0.0176322f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.968
cc_35 VNB N_VGND_c_458_n 0.00981922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_459_n 0.0120484f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.335
cc_37 VNB N_VGND_c_460_n 0.00485511f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.64
cc_38 VNB N_VGND_c_461_n 0.0194756f $X=-0.19 $Y=-0.245 $X2=1.7 $Y2=2.42
cc_39 VNB N_VGND_c_462_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.42
cc_40 VNB N_VGND_c_463_n 0.0208909f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=0.39
cc_41 VNB N_VGND_c_464_n 0.0276253f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=2.42
cc_42 VNB N_VGND_c_465_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_466_n 0.210838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_A_80_72#_c_87_n 0.0251366f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.968
cc_45 VPB N_A_80_72#_M1008_g 0.0421388f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.855
cc_46 VPB N_A_80_72#_c_89_n 0.0199055f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=2.145
cc_47 VPB N_A_80_72#_c_82_n 0.00303017f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.64
cc_48 VPB N_A_80_72#_c_91_n 0.0225865f $X=-0.19 $Y=1.655 $X2=1.7 $Y2=2.42
cc_49 VPB N_A_80_72#_c_92_n 0.0016311f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.42
cc_50 VPB N_A_80_72#_c_93_n 0.00343959f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.335
cc_51 VPB N_A_80_72#_c_84_n 0.0103381f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=1.71
cc_52 VPB N_B1_N_c_180_n 0.0196003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_B1_N_c_181_n 0.0349133f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.7
cc_54 VPB N_B1_N_c_182_n 0.0214345f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B1_N_c_177_n 0.00867502f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.64
cc_56 VPB N_B1_N_c_179_n 0.00470253f $X=-0.19 $Y=1.655 $X2=1.91 $Y2=1.71
cc_57 VPB N_A_196_98#_c_233_n 0.0153004f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.968
cc_58 VPB N_A_196_98#_c_240_n 0.017614f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.145
cc_59 VPB N_A_196_98#_c_241_n 0.0194804f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.855
cc_60 VPB N_A_196_98#_c_242_n 0.0179893f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.335
cc_61 VPB N_A_196_98#_c_243_n 0.0164801f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=0.39
cc_62 VPB N_A_196_98#_c_244_n 0.045059f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=0.39
cc_63 VPB N_A_196_98#_c_245_n 0.0369378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A1_M1009_g 0.040098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A2_M1007_g 0.0520312f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.475
cc_66 VPB A2 0.00677664f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.855
cc_67 VPB X 0.046458f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.7
cc_68 VPB N_VPWR_c_400_n 0.00580687f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.7
cc_69 VPB N_VPWR_c_401_n 0.0499714f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.652
cc_70 VPB N_VPWR_c_402_n 0.0352866f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.855
cc_71 VPB N_VPWR_c_403_n 0.019019f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.64
cc_72 VPB N_VPWR_c_404_n 0.0209183f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.335
cc_73 VPB N_VPWR_c_399_n 0.0810832f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=1.71
cc_74 VPB N_VPWR_c_406_n 0.00401277f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=0.39
cc_75 VPB N_VPWR_c_407_n 0.00401341f $X=-0.19 $Y=1.655 $X2=2.71 $Y2=0.495
cc_76 VPB N_A_419_439#_c_438_n 8.22023e-19 $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.7
cc_77 VPB N_A_419_439#_c_439_n 0.0192003f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.652
cc_78 VPB N_A_419_439#_c_440_n 0.00319687f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.968
cc_79 VPB N_A_419_439#_c_441_n 0.00224906f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.855
cc_80 N_A_80_72#_M1002_g N_B1_N_c_175_n 0.0206039f $X=0.475 $Y=0.7 $X2=-0.19
+ $Y2=-0.245
cc_81 N_A_80_72#_M1008_g N_B1_N_c_181_n 0.00285365f $X=0.475 $Y=2.855 $X2=0
+ $Y2=0
cc_82 N_A_80_72#_c_89_n N_B1_N_c_181_n 0.00964261f $X=0.577 $Y=2.145 $X2=0 $Y2=0
cc_83 N_A_80_72#_c_82_n N_B1_N_c_181_n 0.0026952f $X=0.59 $Y=1.64 $X2=0 $Y2=0
cc_84 N_A_80_72#_c_91_n N_B1_N_c_181_n 0.00588293f $X=1.7 $Y=2.42 $X2=0 $Y2=0
cc_85 N_A_80_72#_c_93_n N_B1_N_c_181_n 2.62871e-19 $X=1.805 $Y=2.335 $X2=0 $Y2=0
cc_86 N_A_80_72#_M1008_g N_B1_N_c_182_n 0.0218163f $X=0.475 $Y=2.855 $X2=0 $Y2=0
cc_87 N_A_80_72#_c_91_n N_B1_N_c_182_n 0.0151453f $X=1.7 $Y=2.42 $X2=0 $Y2=0
cc_88 N_A_80_72#_c_87_n N_B1_N_c_177_n 0.00964261f $X=0.577 $Y=1.968 $X2=0 $Y2=0
cc_89 N_A_80_72#_c_91_n N_B1_N_c_177_n 0.00234067f $X=1.7 $Y=2.42 $X2=0 $Y2=0
cc_90 N_A_80_72#_c_85_n N_B1_N_c_177_n 2.45122e-19 $X=1.91 $Y=1.71 $X2=0 $Y2=0
cc_91 N_A_80_72#_M1002_g N_B1_N_c_178_n 0.00579551f $X=0.475 $Y=0.7 $X2=0 $Y2=0
cc_92 N_A_80_72#_c_82_n N_B1_N_c_178_n 0.00223414f $X=0.59 $Y=1.64 $X2=0 $Y2=0
cc_93 N_A_80_72#_c_83_n N_B1_N_c_178_n 0.00964261f $X=0.59 $Y=1.64 $X2=0 $Y2=0
cc_94 N_A_80_72#_M1002_g N_B1_N_c_179_n 0.00274944f $X=0.475 $Y=0.7 $X2=0 $Y2=0
cc_95 N_A_80_72#_c_82_n N_B1_N_c_179_n 0.020184f $X=0.59 $Y=1.64 $X2=0 $Y2=0
cc_96 N_A_80_72#_c_83_n N_B1_N_c_179_n 0.00232014f $X=0.59 $Y=1.64 $X2=0 $Y2=0
cc_97 N_A_80_72#_c_91_n N_B1_N_c_179_n 0.011439f $X=1.7 $Y=2.42 $X2=0 $Y2=0
cc_98 N_A_80_72#_c_93_n N_B1_N_c_179_n 0.0122209f $X=1.805 $Y=2.335 $X2=0 $Y2=0
cc_99 N_A_80_72#_c_85_n N_B1_N_c_179_n 0.00666441f $X=1.91 $Y=1.71 $X2=0 $Y2=0
cc_100 N_A_80_72#_c_93_n N_A_196_98#_c_233_n 0.00328703f $X=1.805 $Y=2.335 $X2=0
+ $Y2=0
cc_101 N_A_80_72#_c_85_n N_A_196_98#_c_233_n 0.00791002f $X=1.91 $Y=1.71 $X2=0
+ $Y2=0
cc_102 N_A_80_72#_c_93_n N_A_196_98#_c_240_n 0.00735206f $X=1.805 $Y=2.335 $X2=0
+ $Y2=0
cc_103 N_A_80_72#_c_84_n N_A_196_98#_c_240_n 0.00665737f $X=2.625 $Y=1.71 $X2=0
+ $Y2=0
cc_104 N_A_80_72#_c_93_n N_A_196_98#_c_241_n 0.00494361f $X=1.805 $Y=2.335 $X2=0
+ $Y2=0
cc_105 N_A_80_72#_c_93_n N_A_196_98#_c_242_n 9.83928e-19 $X=1.805 $Y=2.335 $X2=0
+ $Y2=0
cc_106 N_A_80_72#_c_84_n N_A_196_98#_c_234_n 0.00182341f $X=2.625 $Y=1.71 $X2=0
+ $Y2=0
cc_107 N_A_80_72#_c_85_n N_A_196_98#_c_234_n 0.00158749f $X=1.91 $Y=1.71 $X2=0
+ $Y2=0
cc_108 N_A_80_72#_c_91_n N_A_196_98#_c_243_n 0.0455245f $X=1.7 $Y=2.42 $X2=0
+ $Y2=0
cc_109 N_A_80_72#_c_93_n N_A_196_98#_c_243_n 0.00265749f $X=1.805 $Y=2.335 $X2=0
+ $Y2=0
cc_110 N_A_80_72#_c_91_n N_A_196_98#_c_244_n 8.05967e-19 $X=1.7 $Y=2.42 $X2=0
+ $Y2=0
cc_111 N_A_80_72#_c_85_n N_A_196_98#_c_236_n 0.0134493f $X=1.91 $Y=1.71 $X2=0
+ $Y2=0
cc_112 N_A_80_72#_c_91_n N_A_196_98#_c_245_n 0.0145705f $X=1.7 $Y=2.42 $X2=0
+ $Y2=0
cc_113 N_A_80_72#_c_93_n N_A_196_98#_c_245_n 0.00557714f $X=1.805 $Y=2.335 $X2=0
+ $Y2=0
cc_114 N_A_80_72#_c_93_n N_A1_M1009_g 0.00341463f $X=1.805 $Y=2.335 $X2=0 $Y2=0
cc_115 N_A_80_72#_c_84_n N_A1_M1009_g 0.0139767f $X=2.625 $Y=1.71 $X2=0 $Y2=0
cc_116 N_A_80_72#_c_131_p N_A1_c_309_n 0.0105642f $X=2.625 $Y=0.39 $X2=0 $Y2=0
cc_117 N_A_80_72#_c_86_n N_A1_c_309_n 0.00571762f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_118 N_A_80_72#_c_84_n N_A1_c_311_n 0.00122414f $X=2.625 $Y=1.71 $X2=0 $Y2=0
cc_119 N_A_80_72#_c_84_n A1 0.0272823f $X=2.625 $Y=1.71 $X2=0 $Y2=0
cc_120 N_A_80_72#_c_131_p A1 0.0172732f $X=2.625 $Y=0.39 $X2=0 $Y2=0
cc_121 N_A_80_72#_c_86_n A1 0.0485778f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_122 N_A_80_72#_c_131_p N_A1_c_313_n 8.05846e-19 $X=2.625 $Y=0.39 $X2=0 $Y2=0
cc_123 N_A_80_72#_c_86_n N_A1_c_313_n 0.00888143f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_124 N_A_80_72#_c_131_p N_A2_M1005_g 0.00552813f $X=2.625 $Y=0.39 $X2=0 $Y2=0
cc_125 N_A_80_72#_c_86_n N_A2_M1005_g 0.0151479f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_126 N_A_80_72#_c_84_n N_A2_M1007_g 0.00264499f $X=2.625 $Y=1.71 $X2=0 $Y2=0
cc_127 N_A_80_72#_c_86_n N_A2_c_353_n 0.00512044f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_128 N_A_80_72#_c_84_n A2 0.0103428f $X=2.625 $Y=1.71 $X2=0 $Y2=0
cc_129 N_A_80_72#_c_86_n A2 0.054768f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_130 N_A_80_72#_c_86_n N_A2_c_356_n 0.00560108f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_131 N_A_80_72#_M1002_g X 4.64676e-19 $X=0.475 $Y=0.7 $X2=0 $Y2=0
cc_132 N_A_80_72#_M1002_g X 0.0560871f $X=0.475 $Y=0.7 $X2=0 $Y2=0
cc_133 N_A_80_72#_c_82_n X 0.0587877f $X=0.59 $Y=1.64 $X2=0 $Y2=0
cc_134 N_A_80_72#_c_92_n X 0.0130058f $X=0.675 $Y=2.42 $X2=0 $Y2=0
cc_135 N_A_80_72#_M1008_g N_VPWR_c_400_n 0.00286392f $X=0.475 $Y=2.855 $X2=0
+ $Y2=0
cc_136 N_A_80_72#_c_89_n N_VPWR_c_400_n 4.65832e-19 $X=0.577 $Y=2.145 $X2=0
+ $Y2=0
cc_137 N_A_80_72#_c_91_n N_VPWR_c_400_n 0.00624333f $X=1.7 $Y=2.42 $X2=0 $Y2=0
cc_138 N_A_80_72#_c_92_n N_VPWR_c_400_n 0.00504797f $X=0.675 $Y=2.42 $X2=0 $Y2=0
cc_139 N_A_80_72#_M1008_g N_VPWR_c_403_n 0.00555245f $X=0.475 $Y=2.855 $X2=0
+ $Y2=0
cc_140 N_A_80_72#_M1008_g N_VPWR_c_399_n 0.00993957f $X=0.475 $Y=2.855 $X2=0
+ $Y2=0
cc_141 N_A_80_72#_c_91_n N_VPWR_c_399_n 0.00798893f $X=1.7 $Y=2.42 $X2=0 $Y2=0
cc_142 N_A_80_72#_c_92_n N_VPWR_c_399_n 0.00327625f $X=0.675 $Y=2.42 $X2=0 $Y2=0
cc_143 N_A_80_72#_c_93_n N_VPWR_c_399_n 0.00704238f $X=1.805 $Y=2.335 $X2=0
+ $Y2=0
cc_144 N_A_80_72#_c_93_n N_A_419_439#_c_438_n 0.00314476f $X=1.805 $Y=2.335
+ $X2=0 $Y2=0
cc_145 N_A_80_72#_c_84_n N_A_419_439#_c_439_n 0.0331913f $X=2.625 $Y=1.71 $X2=0
+ $Y2=0
cc_146 N_A_80_72#_c_93_n N_A_419_439#_c_440_n 0.0117033f $X=1.805 $Y=2.335 $X2=0
+ $Y2=0
cc_147 N_A_80_72#_c_84_n N_A_419_439#_c_440_n 0.0166893f $X=2.625 $Y=1.71 $X2=0
+ $Y2=0
cc_148 N_A_80_72#_M1002_g N_VGND_c_457_n 0.00296421f $X=0.475 $Y=0.7 $X2=0 $Y2=0
cc_149 N_A_80_72#_c_82_n N_VGND_c_457_n 0.00222866f $X=0.59 $Y=1.64 $X2=0 $Y2=0
cc_150 N_A_80_72#_c_83_n N_VGND_c_457_n 0.00274745f $X=0.59 $Y=1.64 $X2=0 $Y2=0
cc_151 N_A_80_72#_c_131_p N_VGND_c_460_n 0.0159098f $X=2.625 $Y=0.39 $X2=0 $Y2=0
cc_152 N_A_80_72#_c_86_n N_VGND_c_460_n 0.00335563f $X=2.71 $Y=1.625 $X2=0 $Y2=0
cc_153 N_A_80_72#_M1002_g N_VGND_c_461_n 0.0049405f $X=0.475 $Y=0.7 $X2=0 $Y2=0
cc_154 N_A_80_72#_c_131_p N_VGND_c_464_n 0.0367462f $X=2.625 $Y=0.39 $X2=0 $Y2=0
cc_155 N_A_80_72#_M1000_d N_VGND_c_466_n 0.00481524f $X=1.985 $Y=0.235 $X2=0
+ $Y2=0
cc_156 N_A_80_72#_M1002_g N_VGND_c_466_n 0.00508379f $X=0.475 $Y=0.7 $X2=0 $Y2=0
cc_157 N_A_80_72#_c_131_p N_VGND_c_466_n 0.0271572f $X=2.625 $Y=0.39 $X2=0 $Y2=0
cc_158 N_A_80_72#_c_131_p A_499_47# 0.00409729f $X=2.625 $Y=0.39 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A_80_72#_c_86_n A_499_47# 0.0018001f $X=2.71 $Y=1.625 $X2=-0.19
+ $Y2=-0.245
cc_160 N_B1_N_c_176_n N_A_196_98#_c_232_n 0.0113968f $X=1.2 $Y=1.175 $X2=0 $Y2=0
cc_161 N_B1_N_c_179_n N_A_196_98#_c_232_n 0.00277674f $X=1.2 $Y=1.19 $X2=0 $Y2=0
cc_162 N_B1_N_c_181_n N_A_196_98#_c_233_n 0.00554605f $X=1.11 $Y=2.385 $X2=0
+ $Y2=0
cc_163 N_B1_N_c_177_n N_A_196_98#_c_233_n 0.0113968f $X=1.2 $Y=1.695 $X2=0 $Y2=0
cc_164 N_B1_N_c_179_n N_A_196_98#_c_233_n 0.00185448f $X=1.2 $Y=1.19 $X2=0 $Y2=0
cc_165 N_B1_N_c_181_n N_A_196_98#_c_241_n 0.0144764f $X=1.11 $Y=2.385 $X2=0
+ $Y2=0
cc_166 N_B1_N_c_179_n N_A_196_98#_c_241_n 0.00168199f $X=1.2 $Y=1.19 $X2=0 $Y2=0
cc_167 N_B1_N_c_178_n N_A_196_98#_c_234_n 0.0113968f $X=1.2 $Y=1.19 $X2=0 $Y2=0
cc_168 N_B1_N_c_182_n N_A_196_98#_c_243_n 0.00443343f $X=1.11 $Y=2.46 $X2=0
+ $Y2=0
cc_169 N_B1_N_c_180_n N_A_196_98#_c_244_n 0.00519109f $X=0.905 $Y=2.535 $X2=0
+ $Y2=0
cc_170 N_B1_N_c_176_n N_A_196_98#_c_235_n 0.00370026f $X=1.2 $Y=1.175 $X2=0
+ $Y2=0
cc_171 N_B1_N_c_179_n N_A_196_98#_c_235_n 0.00448758f $X=1.2 $Y=1.19 $X2=0 $Y2=0
cc_172 N_B1_N_c_176_n N_A_196_98#_c_236_n 0.00152445f $X=1.2 $Y=1.175 $X2=0
+ $Y2=0
cc_173 N_B1_N_c_179_n N_A_196_98#_c_236_n 0.0133535f $X=1.2 $Y=1.19 $X2=0 $Y2=0
cc_174 N_B1_N_c_175_n N_A_196_98#_c_237_n 0.00462977f $X=0.905 $Y=1.025 $X2=0
+ $Y2=0
cc_175 N_B1_N_c_176_n N_A_196_98#_c_275_n 0.00462268f $X=1.2 $Y=1.175 $X2=0
+ $Y2=0
cc_176 N_B1_N_c_179_n N_A_196_98#_c_275_n 0.00855326f $X=1.2 $Y=1.19 $X2=0 $Y2=0
cc_177 N_B1_N_c_180_n N_A_196_98#_c_245_n 0.0053742f $X=0.905 $Y=2.535 $X2=0
+ $Y2=0
cc_178 N_B1_N_c_182_n N_A_196_98#_c_245_n 0.0144764f $X=1.11 $Y=2.46 $X2=0 $Y2=0
cc_179 N_B1_N_c_180_n N_VPWR_c_400_n 0.00286392f $X=0.905 $Y=2.535 $X2=0 $Y2=0
cc_180 N_B1_N_c_180_n N_VPWR_c_401_n 0.00555245f $X=0.905 $Y=2.535 $X2=0 $Y2=0
cc_181 N_B1_N_c_180_n N_VPWR_c_399_n 0.00696322f $X=0.905 $Y=2.535 $X2=0 $Y2=0
cc_182 N_B1_N_c_182_n N_VPWR_c_399_n 7.32236e-19 $X=1.11 $Y=2.46 $X2=0 $Y2=0
cc_183 N_B1_N_c_175_n N_VGND_c_457_n 0.00329204f $X=0.905 $Y=1.025 $X2=0 $Y2=0
cc_184 N_B1_N_c_175_n N_VGND_c_458_n 0.00311925f $X=0.905 $Y=1.025 $X2=0 $Y2=0
cc_185 N_B1_N_c_175_n N_VGND_c_463_n 0.0049405f $X=0.905 $Y=1.025 $X2=0 $Y2=0
cc_186 N_B1_N_c_175_n N_VGND_c_466_n 0.00508379f $X=0.905 $Y=1.025 $X2=0 $Y2=0
cc_187 N_A_196_98#_c_233_n N_A1_M1009_g 0.00552718f $X=1.7 $Y=1.935 $X2=0 $Y2=0
cc_188 N_A_196_98#_c_240_n N_A1_M1009_g 0.0206188f $X=1.945 $Y=2.01 $X2=0 $Y2=0
cc_189 N_A_196_98#_c_235_n N_A1_c_309_n 4.26763e-19 $X=1.705 $Y=0.76 $X2=0 $Y2=0
cc_190 N_A_196_98#_c_238_n N_A1_c_309_n 0.0159852f $X=1.805 $Y=0.765 $X2=0 $Y2=0
cc_191 N_A_196_98#_c_232_n N_A1_c_310_n 0.0138696f $X=1.805 $Y=1.255 $X2=0 $Y2=0
cc_192 N_A_196_98#_c_234_n N_A1_c_311_n 0.0138696f $X=1.805 $Y=1.435 $X2=0 $Y2=0
cc_193 N_A_196_98#_c_235_n A1 0.00596809f $X=1.705 $Y=0.76 $X2=0 $Y2=0
cc_194 N_A_196_98#_c_236_n A1 0.039745f $X=1.79 $Y=0.93 $X2=0 $Y2=0
cc_195 N_A_196_98#_c_237_n A1 0.00486431f $X=1.79 $Y=0.93 $X2=0 $Y2=0
cc_196 N_A_196_98#_c_236_n N_A1_c_313_n 5.06095e-19 $X=1.79 $Y=0.93 $X2=0 $Y2=0
cc_197 N_A_196_98#_c_237_n N_A1_c_313_n 0.0138696f $X=1.79 $Y=0.93 $X2=0 $Y2=0
cc_198 N_A_196_98#_c_242_n N_VPWR_c_401_n 0.00370896f $X=2.02 $Y=2.085 $X2=0
+ $Y2=0
cc_199 N_A_196_98#_c_243_n N_VPWR_c_401_n 0.0352571f $X=1.57 $Y=2.94 $X2=0 $Y2=0
cc_200 N_A_196_98#_c_244_n N_VPWR_c_401_n 0.00617531f $X=1.57 $Y=2.94 $X2=0
+ $Y2=0
cc_201 N_A_196_98#_c_242_n N_VPWR_c_399_n 0.00445256f $X=2.02 $Y=2.085 $X2=0
+ $Y2=0
cc_202 N_A_196_98#_c_243_n N_VPWR_c_399_n 0.0251483f $X=1.57 $Y=2.94 $X2=0 $Y2=0
cc_203 N_A_196_98#_c_244_n N_VPWR_c_399_n 0.00817244f $X=1.57 $Y=2.94 $X2=0
+ $Y2=0
cc_204 N_A_196_98#_c_242_n N_A_419_439#_c_438_n 4.03889e-19 $X=2.02 $Y=2.085
+ $X2=0 $Y2=0
cc_205 N_A_196_98#_c_240_n N_A_419_439#_c_440_n 0.00179855f $X=1.945 $Y=2.01
+ $X2=0 $Y2=0
cc_206 N_A_196_98#_c_235_n N_VGND_c_458_n 0.0220416f $X=1.705 $Y=0.76 $X2=0
+ $Y2=0
cc_207 N_A_196_98#_c_237_n N_VGND_c_458_n 0.00114803f $X=1.79 $Y=0.93 $X2=0
+ $Y2=0
cc_208 N_A_196_98#_c_238_n N_VGND_c_458_n 0.00928197f $X=1.805 $Y=0.765 $X2=0
+ $Y2=0
cc_209 N_A_196_98#_c_235_n N_VGND_c_463_n 0.00509422f $X=1.705 $Y=0.76 $X2=0
+ $Y2=0
cc_210 N_A_196_98#_c_275_n N_VGND_c_463_n 0.00484261f $X=1.12 $Y=0.68 $X2=0
+ $Y2=0
cc_211 N_A_196_98#_c_235_n N_VGND_c_464_n 2.3697e-19 $X=1.705 $Y=0.76 $X2=0
+ $Y2=0
cc_212 N_A_196_98#_c_238_n N_VGND_c_464_n 0.00471611f $X=1.805 $Y=0.765 $X2=0
+ $Y2=0
cc_213 N_A_196_98#_c_235_n N_VGND_c_466_n 0.0104085f $X=1.705 $Y=0.76 $X2=0
+ $Y2=0
cc_214 N_A_196_98#_c_275_n N_VGND_c_466_n 0.00668611f $X=1.12 $Y=0.68 $X2=0
+ $Y2=0
cc_215 N_A_196_98#_c_238_n N_VGND_c_466_n 0.00805858f $X=1.805 $Y=0.765 $X2=0
+ $Y2=0
cc_216 N_A1_c_309_n N_A2_M1005_g 0.0352862f $X=2.36 $Y=0.765 $X2=0 $Y2=0
cc_217 A1 N_A2_M1005_g 2.00237e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_218 N_A1_c_313_n N_A2_M1005_g 0.00693958f $X=2.36 $Y=0.93 $X2=0 $Y2=0
cc_219 N_A1_M1009_g N_A2_M1007_g 0.0196794f $X=2.45 $Y=2.405 $X2=0 $Y2=0
cc_220 N_A1_c_310_n N_A2_c_353_n 0.00693958f $X=2.36 $Y=1.27 $X2=0 $Y2=0
cc_221 N_A1_c_311_n N_A2_c_354_n 0.0196794f $X=2.36 $Y=1.435 $X2=0 $Y2=0
cc_222 N_A1_c_310_n N_A2_c_356_n 0.0196794f $X=2.36 $Y=1.27 $X2=0 $Y2=0
cc_223 N_A1_M1009_g N_VPWR_c_401_n 0.00370896f $X=2.45 $Y=2.405 $X2=0 $Y2=0
cc_224 N_A1_M1009_g N_VPWR_c_402_n 0.00329204f $X=2.45 $Y=2.405 $X2=0 $Y2=0
cc_225 N_A1_M1009_g N_VPWR_c_399_n 0.00445256f $X=2.45 $Y=2.405 $X2=0 $Y2=0
cc_226 N_A1_M1009_g N_A_419_439#_c_438_n 6.71115e-19 $X=2.45 $Y=2.405 $X2=0
+ $Y2=0
cc_227 N_A1_M1009_g N_A_419_439#_c_439_n 0.0144058f $X=2.45 $Y=2.405 $X2=0 $Y2=0
cc_228 N_A1_c_309_n N_VGND_c_458_n 0.00105055f $X=2.36 $Y=0.765 $X2=0 $Y2=0
cc_229 N_A1_c_309_n N_VGND_c_464_n 0.00364081f $X=2.36 $Y=0.765 $X2=0 $Y2=0
cc_230 N_A1_c_309_n N_VGND_c_466_n 0.00548428f $X=2.36 $Y=0.765 $X2=0 $Y2=0
cc_231 N_A2_M1007_g N_VPWR_c_402_n 0.00329204f $X=2.88 $Y=2.405 $X2=0 $Y2=0
cc_232 N_A2_M1007_g N_VPWR_c_404_n 0.00370896f $X=2.88 $Y=2.405 $X2=0 $Y2=0
cc_233 N_A2_M1007_g N_VPWR_c_399_n 0.00445256f $X=2.88 $Y=2.405 $X2=0 $Y2=0
cc_234 N_A2_M1007_g N_A_419_439#_c_439_n 0.0205654f $X=2.88 $Y=2.405 $X2=0 $Y2=0
cc_235 N_A2_c_354_n N_A_419_439#_c_439_n 0.00163535f $X=3.015 $Y=1.51 $X2=0
+ $Y2=0
cc_236 A2 N_A_419_439#_c_439_n 0.0167857f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_237 N_A2_M1007_g N_A_419_439#_c_441_n 0.00143084f $X=2.88 $Y=2.405 $X2=0
+ $Y2=0
cc_238 N_A2_M1005_g N_VGND_c_460_n 0.00574314f $X=2.81 $Y=0.445 $X2=0 $Y2=0
cc_239 N_A2_c_353_n N_VGND_c_460_n 0.00135706f $X=2.98 $Y=0.99 $X2=0 $Y2=0
cc_240 A2 N_VGND_c_460_n 0.00977736f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_241 N_A2_M1005_g N_VGND_c_464_n 0.00496782f $X=2.81 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A2_M1005_g N_VGND_c_466_n 0.00954337f $X=2.81 $Y=0.445 $X2=0 $Y2=0
cc_243 N_A2_c_353_n N_VGND_c_466_n 0.00284108f $X=2.98 $Y=0.99 $X2=0 $Y2=0
cc_244 A2 N_VGND_c_466_n 0.00222711f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_245 X N_VPWR_c_403_n 0.00997412f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_246 X N_VPWR_c_399_n 0.00780853f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_247 X N_VGND_c_457_n 0.00123197f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_248 X N_VGND_c_461_n 0.00617805f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_249 X N_VGND_c_466_n 0.00706876f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_250 N_VPWR_c_399_n N_A_419_439#_c_438_n 0.00810724f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_402_n N_A_419_439#_c_439_n 0.0146902f $X=2.665 $Y=2.49 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_399_n N_A_419_439#_c_441_n 0.00810724f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_253 N_VGND_c_466_n A_499_47# 0.00194154f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
