* File: sky130_fd_sc_lp__clkbuflp_4.pex.spice
* Created: Fri Aug 28 10:15:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_4%A 3 7 11 15 17 18 28
c46 3 0 2.20622e-20 $X=0.475 $Y=0.555
r47 27 28 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.835 $Y=1.4
+ $X2=1.055 $Y2=1.4
r48 25 27 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.565 $Y=1.4
+ $X2=0.835 $Y2=1.4
r49 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.565
+ $Y=1.4 $X2=0.565 $Y2=1.4
r50 23 25 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.525 $Y=1.4 $X2=0.565
+ $Y2=1.4
r51 21 23 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.475 $Y=1.4 $X2=0.525
+ $Y2=1.4
r52 18 26 6.625 $w=4.88e-07 $l=3.43402e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.42 $Y2=1.4
r53 17 26 2.625 $w=4.88e-07 $l=1.05e-07 $layer=LI1_cond $X=0.42 $Y=1.295
+ $X2=0.42 $Y2=1.4
r54 13 28 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.565
+ $X2=1.055 $Y2=1.4
r55 13 15 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.055 $Y=1.565
+ $X2=1.055 $Y2=2.585
r56 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=1.4
r57 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=0.555
r58 5 23 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.565
+ $X2=0.525 $Y2=1.4
r59 5 7 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=0.525 $Y=1.565
+ $X2=0.525 $Y2=2.585
r60 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=1.4
r61 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_4%A_130_417# 1 2 9 13 17 21 25 29 33 37 41
+ 45 51 55 56 57 67
c115 57 0 2.20622e-20 $X=1.057 $Y=1.37
r116 66 67 40.7324 $w=3.4e-07 $l=2.4e-07 $layer=POLY_cond $X=2.935 $Y=1.375
+ $X2=3.175 $Y2=1.375
r117 65 66 49.2183 $w=3.4e-07 $l=2.9e-07 $layer=POLY_cond $X=2.645 $Y=1.375
+ $X2=2.935 $Y2=1.375
r118 64 65 11.8803 $w=3.4e-07 $l=7e-08 $layer=POLY_cond $X=2.575 $Y=1.375
+ $X2=2.645 $Y2=1.375
r119 63 64 72.9789 $w=3.4e-07 $l=4.3e-07 $layer=POLY_cond $X=2.145 $Y=1.375
+ $X2=2.575 $Y2=1.375
r120 62 63 5.09155 $w=3.4e-07 $l=3e-08 $layer=POLY_cond $X=2.115 $Y=1.375
+ $X2=2.145 $Y2=1.375
r121 58 60 33.9437 $w=3.4e-07 $l=2e-07 $layer=POLY_cond $X=1.585 $Y=1.375
+ $X2=1.785 $Y2=1.375
r122 55 56 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.84 $Y=2.23
+ $X2=0.84 $Y2=2.065
r123 52 62 25.4577 $w=3.4e-07 $l=1.5e-07 $layer=POLY_cond $X=1.965 $Y=1.375
+ $X2=2.115 $Y2=1.375
r124 52 60 30.5493 $w=3.4e-07 $l=1.8e-07 $layer=POLY_cond $X=1.965 $Y=1.375
+ $X2=1.785 $Y2=1.375
r125 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.965
+ $Y=1.37 $X2=1.965 $Y2=1.37
r126 49 57 0.466467 $w=3.3e-07 $l=1.73e-07 $layer=LI1_cond $X=1.23 $Y=1.37
+ $X2=1.057 $Y2=1.37
r127 49 51 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=1.23 $Y=1.37
+ $X2=1.965 $Y2=1.37
r128 47 57 6.31733 $w=2.57e-07 $l=2.03912e-07 $layer=LI1_cond $X=0.97 $Y=1.535
+ $X2=1.057 $Y2=1.37
r129 47 56 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.97 $Y=1.535
+ $X2=0.97 $Y2=2.065
r130 43 57 6.31733 $w=2.57e-07 $l=1.65e-07 $layer=LI1_cond $X=1.057 $Y=1.205
+ $X2=1.057 $Y2=1.37
r131 43 45 27.2244 $w=3.43e-07 $l=8.15e-07 $layer=LI1_cond $X=1.057 $Y=1.205
+ $X2=1.057 $Y2=0.39
r132 39 55 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=0.84 $Y=2.28 $X2=0.84
+ $Y2=2.23
r133 39 41 16.8846 $w=4.28e-07 $l=6.3e-07 $layer=LI1_cond $X=0.84 $Y=2.28
+ $X2=0.84 $Y2=2.91
r134 35 67 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.175 $Y=1.545
+ $X2=3.175 $Y2=1.375
r135 35 37 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=3.175 $Y=1.545
+ $X2=3.175 $Y2=2.585
r136 31 66 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.935 $Y=1.205
+ $X2=2.935 $Y2=1.375
r137 31 33 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.935 $Y=1.205
+ $X2=2.935 $Y2=0.51
r138 27 65 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.645 $Y=1.545
+ $X2=2.645 $Y2=1.375
r139 27 29 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.645 $Y=1.545
+ $X2=2.645 $Y2=2.585
r140 23 64 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.575 $Y=1.205
+ $X2=2.575 $Y2=1.375
r141 23 25 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.575 $Y=1.205
+ $X2=2.575 $Y2=0.51
r142 19 63 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.145 $Y=1.205
+ $X2=2.145 $Y2=1.375
r143 19 21 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.145 $Y=1.205
+ $X2=2.145 $Y2=0.51
r144 15 62 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.115 $Y=1.545
+ $X2=2.115 $Y2=1.375
r145 15 17 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.115 $Y=1.545
+ $X2=2.115 $Y2=2.585
r146 11 60 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.785 $Y=1.205
+ $X2=1.785 $Y2=1.375
r147 11 13 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.785 $Y=1.205
+ $X2=1.785 $Y2=0.51
r148 7 58 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.585 $Y=1.545
+ $X2=1.585 $Y2=1.375
r149 7 9 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.585 $Y=1.545
+ $X2=1.585 $Y2=2.585
r150 2 55 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.085 $X2=0.79 $Y2=2.23
r151 2 41 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.085 $X2=0.79 $Y2=2.91
r152 1 45 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.235 $X2=1.05 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_4%VPWR 1 2 3 4 13 15 21 27 31 33 38 39 41
+ 42 43 52 61
r56 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 55 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r60 52 60 4.52492 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.557 $Y2=3.33
r61 52 54 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r64 48 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r65 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 45 57 4.43563 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r67 45 47 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 43 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 43 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 41 50 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.38 $Y2=3.33
r72 40 54 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.38 $Y2=3.33
r74 38 47 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.2 $Y2=3.33
r75 38 39 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.355 $Y2=3.33
r76 37 50 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r77 37 39 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.355 $Y2=3.33
r78 33 36 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.44 $Y=2.23
+ $X2=3.44 $Y2=2.91
r79 31 60 3.24126 $w=3.3e-07 $l=1.53734e-07 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.557 $Y2=3.33
r80 31 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=2.91
r81 27 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.38 $Y=2.23
+ $X2=2.38 $Y2=2.91
r82 25 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=3.33
r83 25 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=2.91
r84 21 24 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.355 $Y=2.23
+ $X2=1.355 $Y2=2.91
r85 19 39 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=3.33
r86 19 24 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=2.91
r87 15 18 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=0.275 $Y=2.23
+ $X2=0.275 $Y2=2.91
r88 13 57 3.08204 $w=3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.212 $Y2=3.33
r89 13 18 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.91
r90 4 36 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=2.085 $X2=3.44 $Y2=2.91
r91 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=2.085 $X2=3.44 $Y2=2.23
r92 3 30 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=2.085 $X2=2.38 $Y2=2.91
r93 3 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=2.085 $X2=2.38 $Y2=2.23
r94 2 24 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=2.085 $X2=1.32 $Y2=2.91
r95 2 21 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=2.085 $X2=1.32 $Y2=2.23
r96 1 18 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.085 $X2=0.26 $Y2=2.91
r97 1 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.085 $X2=0.26 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_4%X 1 2 3 12 17 20 24 25 26 28 30 48 56 62
+ 68
r64 48 68 0.868121 $w=6.18e-07 $l=4.5e-08 $layer=LI1_cond $X=3.12 $Y=1.48
+ $X2=3.075 $Y2=1.48
r65 43 62 11.6006 $w=7.03e-07 $l=2.1e-07 $layer=LI1_cond $X=2.565 $Y=1.522
+ $X2=2.355 $Y2=1.522
r66 28 68 0.543556 $w=7.03e-07 $l=2e-08 $layer=LI1_cond $X=3.055 $Y=1.522
+ $X2=3.075 $Y2=1.522
r67 28 66 2.46002 $w=7.03e-07 $l=1.45e-07 $layer=LI1_cond $X=3.055 $Y=1.522
+ $X2=2.91 $Y2=1.522
r68 28 30 8.87413 $w=6.18e-07 $l=4.6e-07 $layer=LI1_cond $X=3.14 $Y=1.48 $X2=3.6
+ $Y2=1.48
r69 28 48 0.385832 $w=6.18e-07 $l=2e-08 $layer=LI1_cond $X=3.14 $Y=1.48 $X2=3.12
+ $Y2=1.48
r70 26 66 4.58073 $w=7.03e-07 $l=2.7e-07 $layer=LI1_cond $X=2.64 $Y=1.522
+ $X2=2.91 $Y2=1.522
r71 26 43 1.27242 $w=7.03e-07 $l=7.5e-08 $layer=LI1_cond $X=2.64 $Y=1.522
+ $X2=2.565 $Y2=1.522
r72 25 43 6.72258 $w=4.18e-07 $l=2.45e-07 $layer=LI1_cond $X=2.565 $Y=0.925
+ $X2=2.565 $Y2=1.17
r73 25 60 7.40856 $w=4.18e-07 $l=2.7e-07 $layer=LI1_cond $X=2.565 $Y=0.925
+ $X2=2.565 $Y2=0.655
r74 24 60 2.9929 $w=5.78e-07 $l=1e-07 $layer=LI1_cond $X=2.485 $Y=0.555
+ $X2=2.485 $Y2=0.655
r75 24 56 1.34043 $w=5.78e-07 $l=6.5e-08 $layer=LI1_cond $X=2.485 $Y=0.555
+ $X2=2.485 $Y2=0.49
r76 20 22 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.91 $Y=2.23
+ $X2=2.91 $Y2=2.91
r77 18 66 5.19532 $w=3.3e-07 $l=3.53e-07 $layer=LI1_cond $X=2.91 $Y=1.875
+ $X2=2.91 $Y2=1.522
r78 18 20 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.91 $Y=1.875
+ $X2=2.91 $Y2=2.23
r79 17 62 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.015 $Y=1.79
+ $X2=2.355 $Y2=1.79
r80 12 14 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.85 $Y=2.23
+ $X2=1.85 $Y2=2.91
r81 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.85 $Y=1.875
+ $X2=2.015 $Y2=1.79
r82 10 12 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.85 $Y=1.875
+ $X2=1.85 $Y2=2.23
r83 3 22 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=2.085 $X2=2.91 $Y2=2.91
r84 3 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=2.085 $X2=2.91 $Y2=2.23
r85 2 14 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.085 $X2=1.85 $Y2=2.91
r86 2 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.085 $X2=1.85 $Y2=2.23
r87 1 56 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.22
+ $Y=0.235 $X2=2.36 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_4%VGND 1 2 3 10 12 16 20 22 24 29 36 37 43
+ 46
r47 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r49 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 37 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r51 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r52 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.15
+ $Y2=0
r53 34 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.6
+ $Y2=0
r54 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r55 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r56 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.57
+ $Y2=0
r57 30 32 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=2.64
+ $Y2=0
r58 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=3.15
+ $Y2=0
r59 29 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=2.64
+ $Y2=0
r60 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r61 28 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r62 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r63 25 40 4.43563 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r64 25 27 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=1.2
+ $Y2=0
r65 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.57
+ $Y2=0
r66 24 27 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.2
+ $Y2=0
r67 22 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r68 22 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r69 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=0.085
+ $X2=3.15 $Y2=0
r70 18 20 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.15 $Y=0.085
+ $X2=3.15 $Y2=0.49
r71 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0
r72 14 16 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0.49
r73 10 40 3.08204 $w=3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.212 $Y2=0
r74 10 12 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.39
r75 3 20 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.235 $X2=3.15 $Y2=0.49
r76 2 16 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=1.57 $Y2=0.49
r77 1 12 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

