* File: sky130_fd_sc_lp__sdfbbn_2.pex.spice
* Created: Fri Aug 28 11:27:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%SCD 2 5 8 11 13 16 18 21 22
r37 21 23 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=1.38 $X2=0.42
+ $Y2=1.215
r38 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.38 $X2=0.385 $Y2=1.38
r39 18 22 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.55
+ $X2=0.385 $Y2=1.55
r40 14 16 48.7128 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=0.545 $Y=2.2
+ $X2=0.64 $Y2=2.2
r41 9 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.64 $Y=2.275
+ $X2=0.64 $Y2=2.2
r42 9 11 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=0.64 $Y=2.275
+ $X2=0.64 $Y2=2.725
r43 8 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.545 $Y=2.125
+ $X2=0.545 $Y2=2.2
r44 8 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.545 $Y=2.125
+ $X2=0.545 $Y2=1.885
r45 5 23 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.545 $Y=0.805
+ $X2=0.545 $Y2=1.215
r46 2 13 50.5417 $w=4e-07 $l=2e-07 $layer=POLY_cond $X=0.42 $Y=1.685 $X2=0.42
+ $Y2=1.885
r47 1 21 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=0.42 $Y=1.415 $X2=0.42
+ $Y2=1.38
r48 1 2 37.5404 $w=4e-07 $l=2.7e-07 $layer=POLY_cond $X=0.42 $Y=1.415 $X2=0.42
+ $Y2=1.685
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%D 3 6 9 10 11 12 13 14 19
r47 13 14 14.4055 $w=2.98e-07 $l=3.75e-07 $layer=LI1_cond $X=1.645 $Y=1.29
+ $X2=1.645 $Y2=1.665
r48 13 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.29 $X2=1.63 $Y2=1.29
r49 12 13 14.0214 $w=2.98e-07 $l=3.65e-07 $layer=LI1_cond $X=1.645 $Y=0.925
+ $X2=1.645 $Y2=1.29
r50 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.63 $Y=1.63
+ $X2=1.63 $Y2=1.29
r51 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.63
+ $X2=1.63 $Y2=1.795
r52 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.125
+ $X2=1.63 $Y2=1.29
r53 6 11 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=1.54 $Y=2.725
+ $X2=1.54 $Y2=1.795
r54 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.54 $Y=0.805 $X2=1.54
+ $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_407_93# 1 2 9 11 13 18 25 26 28 29 30 32
c69 13 0 8.92047e-20 $X=2.11 $Y=2.725
r70 30 35 2.89128 $w=5e-07 $l=1.7e-07 $layer=LI1_cond $X=3.195 $Y=1.515
+ $X2=3.195 $Y2=1.685
r71 30 32 16.9843 $w=4.98e-07 $l=7.1e-07 $layer=LI1_cond $X=3.195 $Y=1.515
+ $X2=3.195 $Y2=0.805
r72 28 35 4.25188 $w=3.4e-07 $l=2.5e-07 $layer=LI1_cond $X=2.945 $Y=1.685
+ $X2=3.195 $Y2=1.685
r73 28 29 12.3718 $w=3.38e-07 $l=3.65e-07 $layer=LI1_cond $X=2.945 $Y=1.685
+ $X2=2.58 $Y2=1.685
r74 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.415
+ $Y=1.35 $X2=2.415 $Y2=1.35
r75 23 29 6.999 $w=3.4e-07 $l=2.25078e-07 $layer=LI1_cond $X=2.452 $Y=1.515
+ $X2=2.58 $Y2=1.685
r76 23 25 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.452 $Y=1.515
+ $X2=2.452 $Y2=1.35
r77 22 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.415 $Y=1.69
+ $X2=2.415 $Y2=1.35
r78 18 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.415 $Y=1.335
+ $X2=2.415 $Y2=1.35
r79 15 18 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=2.11 $Y=1.26
+ $X2=2.415 $Y2=1.26
r80 11 22 73.505 $w=2e-07 $l=3.75786e-07 $layer=POLY_cond $X=2.11 $Y=2.005
+ $X2=2.415 $Y2=1.847
r81 11 13 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.11 $Y=2.005
+ $X2=2.11 $Y2=2.725
r82 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.11 $Y=1.185
+ $X2=2.11 $Y2=1.26
r83 7 9 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.11 $Y=1.185 $X2=2.11
+ $Y2=0.805
r84 2 35 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.535 $X2=3.28 $Y2=1.685
r85 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.97
+ $Y=0.595 $X2=3.11 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%SCE 4 6 7 8 11 16 19 21 24 26 29
r74 29 31 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.042 $Y=1.38
+ $X2=1.042 $Y2=1.215
r75 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.06
+ $Y=1.38 $X2=1.06 $Y2=1.38
r76 26 30 2.49927 $w=6.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.55 $X2=1.06
+ $Y2=1.55
r77 22 24 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2.895 $Y=1.165
+ $X2=3.065 $Y2=1.165
r78 17 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.065 $Y=1.24
+ $X2=3.065 $Y2=1.165
r79 17 19 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.065 $Y=1.24
+ $X2=3.065 $Y2=1.855
r80 14 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.895 $Y=1.09
+ $X2=2.895 $Y2=1.165
r81 14 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.895 $Y=1.09
+ $X2=2.895 $Y2=0.805
r82 13 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.895 $Y=0.255
+ $X2=2.895 $Y2=0.805
r83 11 21 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.15 $Y=2.725
+ $X2=1.15 $Y2=1.885
r84 7 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.82 $Y=0.18
+ $X2=2.895 $Y2=0.255
r85 7 8 928.106 $w=1.5e-07 $l=1.81e-06 $layer=POLY_cond $X=2.82 $Y=0.18 $X2=1.01
+ $Y2=0.18
r86 6 21 49.3547 $w=3.65e-07 $l=1.82e-07 $layer=POLY_cond $X=1.042 $Y=1.703
+ $X2=1.042 $Y2=1.885
r87 5 29 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=1.042 $Y=1.397
+ $X2=1.042 $Y2=1.38
r88 5 6 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=1.042 $Y=1.397
+ $X2=1.042 $Y2=1.703
r89 4 31 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.935 $Y=0.805
+ $X2=0.935 $Y2=1.215
r90 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.935 $Y=0.255
+ $X2=1.01 $Y2=0.18
r91 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.935 $Y=0.255
+ $X2=0.935 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%CLK_N 3 7 11 12 13 14 18
r34 13 14 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=4.035 $Y=1.275
+ $X2=4.035 $Y2=1.665
r35 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.035
+ $Y=1.275 $X2=4.035 $Y2=1.275
r36 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.035 $Y=1.615
+ $X2=4.035 $Y2=1.275
r37 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.035 $Y=1.615
+ $X2=4.035 $Y2=1.78
r38 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.035 $Y=1.11
+ $X2=4.035 $Y2=1.275
r39 7 12 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=4.125 $Y=2.375
+ $X2=4.125 $Y2=1.78
r40 3 10 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.125 $Y=0.685
+ $X2=4.125 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_840_95# 1 2 10 14 15 16 17 18 21 26 29 30
+ 32 33 34 38 40 42 46 47 49 50 52 53 54 56 57 58 60 61 62 65 66 73 77 88
c219 77 0 1.2181e-19 $X=10.955 $Y=1.51
c220 66 0 3.07529e-20 $X=11.855 $Y=1.865
c221 65 0 1.22987e-19 $X=11.855 $Y=1.865
c222 47 0 1.09444e-19 $X=6.855 $Y=1.38
c223 33 0 1.28128e-19 $X=5.235 $Y=1.34
r224 77 88 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.955 $Y=1.51
+ $X2=10.955 $Y2=1.345
r225 76 78 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=10.9 $Y=1.51
+ $X2=10.9 $Y2=1.675
r226 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.955
+ $Y=1.51 $X2=10.955 $Y2=1.51
r227 73 76 8.64332 $w=4.38e-07 $l=3.3e-07 $layer=LI1_cond $X=10.9 $Y=1.18
+ $X2=10.9 $Y2=1.51
r228 71 72 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.605
+ $Y=1.17 $X2=4.605 $Y2=1.17
r229 69 71 15.9919 $w=3.7e-07 $l=4.85e-07 $layer=LI1_cond $X=4.472 $Y=0.685
+ $X2=4.472 $Y2=1.17
r230 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.855
+ $Y=1.865 $X2=11.855 $Y2=1.865
r231 63 65 35.9702 $w=3.28e-07 $l=1.03e-06 $layer=LI1_cond $X=11.855 $Y=2.895
+ $X2=11.855 $Y2=1.865
r232 61 63 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.69 $Y=2.98
+ $X2=11.855 $Y2=2.895
r233 61 62 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=11.69 $Y=2.98
+ $X2=10.85 $Y2=2.98
r234 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.765 $Y=2.895
+ $X2=10.85 $Y2=2.98
r235 60 78 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=10.765 $Y=2.895
+ $X2=10.765 $Y2=1.675
r236 57 73 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=10.68 $Y=1.18
+ $X2=10.9 $Y2=1.18
r237 57 58 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=10.68 $Y=1.18
+ $X2=10.025 $Y2=1.18
r238 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.94 $Y=1.095
+ $X2=10.025 $Y2=1.18
r239 55 56 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=9.94 $Y=0.435
+ $X2=9.94 $Y2=1.095
r240 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.855 $Y=0.35
+ $X2=9.94 $Y2=0.435
r241 53 54 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=9.855 $Y=0.35
+ $X2=8.145 $Y2=0.35
r242 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.06 $Y=0.435
+ $X2=8.145 $Y2=0.35
r243 51 52 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.06 $Y=0.435
+ $X2=8.06 $Y2=0.83
r244 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.975 $Y=0.915
+ $X2=8.06 $Y2=0.83
r245 49 50 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=7.975 $Y=0.915
+ $X2=6.945 $Y2=0.915
r246 47 83 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.855 $Y=1.38
+ $X2=6.72 $Y2=1.38
r247 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.855
+ $Y=1.38 $X2=6.855 $Y2=1.38
r248 44 50 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=6.857 $Y=1
+ $X2=6.945 $Y2=0.915
r249 44 46 24.0831 $w=1.73e-07 $l=3.8e-07 $layer=LI1_cond $X=6.857 $Y=1
+ $X2=6.857 $Y2=1.38
r250 40 71 0.304073 $w=3.7e-07 $l=1.28452e-07 $layer=LI1_cond $X=4.597 $Y=1.177
+ $X2=4.472 $Y2=1.17
r251 40 42 34.1724 $w=3.43e-07 $l=1.023e-06 $layer=LI1_cond $X=4.597 $Y=1.177
+ $X2=4.597 $Y2=2.2
r252 38 66 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=11.855 $Y=2.305
+ $X2=11.855 $Y2=1.865
r253 35 38 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=11.49 $Y=2.38
+ $X2=11.855 $Y2=2.38
r254 33 72 50.3087 $w=6.7e-07 $l=6.3e-07 $layer=POLY_cond $X=5.235 $Y=1.34
+ $X2=4.605 $Y2=1.34
r255 33 34 11.9686 $w=6.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.235 $Y=1.34
+ $X2=5.31 $Y2=1.34
r256 30 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.49 $Y=2.455
+ $X2=11.49 $Y2=2.38
r257 30 32 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.49 $Y=2.455
+ $X2=11.49 $Y2=2.74
r258 29 88 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.015 $Y=0.915
+ $X2=11.015 $Y2=1.345
r259 24 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.72 $Y=1.215
+ $X2=6.72 $Y2=1.38
r260 24 26 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.72 $Y=1.215
+ $X2=6.72 $Y2=0.895
r261 23 26 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.72 $Y=0.26
+ $X2=6.72 $Y2=0.895
r262 19 21 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=6.29 $Y=3.06
+ $X2=6.29 $Y2=2.525
r263 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.215 $Y=3.135
+ $X2=6.29 $Y2=3.06
r264 17 18 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=6.215 $Y=3.135
+ $X2=5.385 $Y2=3.135
r265 15 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.645 $Y=0.185
+ $X2=6.72 $Y2=0.26
r266 15 16 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=6.645 $Y=0.185
+ $X2=5.385 $Y2=0.185
r267 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.31 $Y=3.06
+ $X2=5.385 $Y2=3.135
r268 12 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.31 $Y=3.06
+ $X2=5.31 $Y2=2.665
r269 11 34 56.3093 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.31 $Y=1.675
+ $X2=5.31 $Y2=1.34
r270 11 14 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=5.31 $Y=1.675
+ $X2=5.31 $Y2=2.665
r271 8 34 56.3093 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.31 $Y=1.005
+ $X2=5.31 $Y2=1.34
r272 8 10 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=5.31 $Y=1.005
+ $X2=5.31 $Y2=0.545
r273 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.31 $Y=0.26
+ $X2=5.385 $Y2=0.185
r274 7 10 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.31 $Y=0.26
+ $X2=5.31 $Y2=0.545
r275 2 42 300 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_PDIFF $count=2 $X=4.2
+ $Y=2.055 $X2=4.51 $Y2=2.2
r276 1 69 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.475 $X2=4.34 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_1423_401# 1 2 9 13 17 21 25 30 32 36 43
+ 44 46 48 49 50 53
c124 50 0 1.26967e-19 $X=10.17 $Y=1.575
c125 36 0 8.25457e-20 $X=7.565 $Y=1.99
r126 49 57 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=10.375 $Y=1.57
+ $X2=10.375 $Y2=1.735
r127 49 56 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=10.375 $Y=1.57
+ $X2=10.375 $Y2=1.405
r128 48 50 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.335 $Y=1.575
+ $X2=10.17 $Y2=1.575
r129 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.335
+ $Y=1.57 $X2=10.335 $Y2=1.57
r130 42 44 9.76211 $w=6.78e-07 $l=5.55e-07 $layer=LI1_cond $X=8.69 $Y=2.415
+ $X2=9.245 $Y2=2.415
r131 42 43 10.6764 $w=6.78e-07 $l=1.65e-07 $layer=LI1_cond $X=8.69 $Y=2.415
+ $X2=8.525 $Y2=2.415
r132 37 53 38.6272 $w=2.87e-07 $l=2.3e-07 $layer=POLY_cond $X=7.565 $Y=1.99
+ $X2=7.335 $Y2=1.99
r133 36 39 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=7.565 $Y=1.99
+ $X2=7.565 $Y2=2.16
r134 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.565
+ $Y=1.99 $X2=7.565 $Y2=1.99
r135 34 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.33 $Y=1.53
+ $X2=9.245 $Y2=1.53
r136 34 50 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=9.33 $Y=1.53
+ $X2=10.17 $Y2=1.53
r137 32 44 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=9.245 $Y=2.075
+ $X2=9.245 $Y2=2.415
r138 31 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.245 $Y=1.615
+ $X2=9.245 $Y2=1.53
r139 31 32 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=9.245 $Y=1.615
+ $X2=9.245 $Y2=2.075
r140 30 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.245 $Y=1.445
+ $X2=9.245 $Y2=1.53
r141 29 30 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.245 $Y=1.225
+ $X2=9.245 $Y2=1.445
r142 25 29 7.10164 $w=2.18e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.16 $Y=1.095
+ $X2=9.245 $Y2=1.225
r143 25 27 7.09196 $w=2.58e-07 $l=1.6e-07 $layer=LI1_cond $X=9.16 $Y=1.095 $X2=9
+ $Y2=1.095
r144 24 39 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=7.655 $Y=2.16
+ $X2=7.565 $Y2=2.16
r145 24 43 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=7.655 $Y=2.16
+ $X2=8.525 $Y2=2.16
r146 21 57 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.505 $Y=2.315
+ $X2=10.505 $Y2=1.735
r147 17 56 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=10.505 $Y=0.915
+ $X2=10.505 $Y2=1.405
r148 11 53 17.9292 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.335 $Y=1.825
+ $X2=7.335 $Y2=1.99
r149 11 13 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=7.335 $Y=1.825
+ $X2=7.335 $Y2=0.895
r150 7 53 24.3519 $w=2.87e-07 $l=2.26164e-07 $layer=POLY_cond $X=7.19 $Y=2.155
+ $X2=7.335 $Y2=1.99
r151 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.19 $Y=2.155
+ $X2=7.19 $Y2=2.525
r152 2 42 300 $w=1.7e-07 $l=4.64354e-07 $layer=licon1_PDIFF $count=2 $X=8.41
+ $Y=1.895 $X2=8.69 $Y2=2.24
r153 1 27 182 $w=1.7e-07 $l=7.58436e-07 $layer=licon1_NDIFF $count=1 $X=8.8
+ $Y=0.465 $X2=9 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%SET_B 1 3 6 10 12 13 15 18 20 22 23 29 30
+ 33 34 37 39
c132 33 0 1.38231e-19 $X=8.275 $Y=1.38
c133 23 0 1.4512e-19 $X=8.545 $Y=1.295
c134 22 0 1.78884e-19 $X=12.575 $Y=1.295
c135 18 0 3.77964e-20 $X=13.065 $Y=2.105
c136 13 0 6.75576e-20 $X=13.065 $Y=2.18
r137 37 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.785 $Y=1.51
+ $X2=12.785 $Y2=1.675
r138 37 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.785 $Y=1.51
+ $X2=12.785 $Y2=1.345
r139 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.785
+ $Y=1.51 $X2=12.785 $Y2=1.51
r140 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.275 $Y=1.38
+ $X2=8.275 $Y2=1.545
r141 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.275
+ $Y=1.38 $X2=8.275 $Y2=1.38
r142 30 38 7.18189 $w=3.43e-07 $l=2.15e-07 $layer=LI1_cond $X=12.777 $Y=1.295
+ $X2=12.777 $Y2=1.51
r143 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=1.295
+ $X2=12.72 $Y2=1.295
r144 25 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.295
+ $X2=8.4 $Y2=1.295
r145 23 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=1.295
+ $X2=8.4 $Y2=1.295
r146 22 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.575 $Y=1.295
+ $X2=12.72 $Y2=1.295
r147 22 23 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=12.575 $Y=1.295
+ $X2=8.545 $Y2=1.295
r148 20 38 5.17764 $w=3.43e-07 $l=1.55e-07 $layer=LI1_cond $X=12.777 $Y=1.665
+ $X2=12.777 $Y2=1.51
r149 16 18 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=12.875 $Y=2.105
+ $X2=13.065 $Y2=2.105
r150 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.065 $Y=2.18
+ $X2=13.065 $Y2=2.105
r151 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=13.065 $Y=2.18
+ $X2=13.065 $Y2=2.675
r152 12 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.875 $Y=2.03
+ $X2=12.875 $Y2=2.105
r153 12 40 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=12.875 $Y=2.03
+ $X2=12.875 $Y2=1.675
r154 10 39 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.795 $Y=0.915
+ $X2=12.795 $Y2=1.345
r155 6 35 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=8.335 $Y=2.315
+ $X2=8.335 $Y2=1.545
r156 1 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.275 $Y=1.215
+ $X2=8.275 $Y2=1.38
r157 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.275 $Y=1.215
+ $X2=8.275 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_1273_137# 1 2 9 13 17 21 23 26 27 28 29
+ 33 34 36 37
c111 36 0 1.09444e-19 $X=6.585 $Y=2.16
c112 34 0 2.20873e-19 $X=8.815 $Y=1.57
c113 33 0 2.83351e-19 $X=8.815 $Y=1.57
c114 29 0 1.92809e-19 $X=8.705 $Y=1.81
c115 26 0 1.18451e-19 $X=7.21 $Y=2.075
r116 37 39 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.92 $Y=1.56
+ $X2=7.92 $Y2=1.81
r117 34 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.815 $Y=1.57
+ $X2=8.815 $Y2=1.735
r118 34 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.815 $Y=1.57
+ $X2=8.815 $Y2=1.405
r119 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.815
+ $Y=1.57 $X2=8.815 $Y2=1.57
r120 31 33 6.49559 $w=2.73e-07 $l=1.55e-07 $layer=LI1_cond $X=8.842 $Y=1.725
+ $X2=8.842 $Y2=1.57
r121 30 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.005 $Y=1.81
+ $X2=7.92 $Y2=1.81
r122 29 31 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=8.705 $Y=1.81
+ $X2=8.842 $Y2=1.725
r123 29 30 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.705 $Y=1.81
+ $X2=8.005 $Y2=1.81
r124 27 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.835 $Y=1.56
+ $X2=7.92 $Y2=1.56
r125 27 28 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=7.835 $Y=1.56
+ $X2=7.295 $Y2=1.56
r126 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.21 $Y=1.645
+ $X2=7.295 $Y2=1.56
r127 25 26 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.21 $Y=1.645
+ $X2=7.21 $Y2=2.075
r128 24 36 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.75 $Y=2.16
+ $X2=6.585 $Y2=2.16
r129 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.125 $Y=2.16
+ $X2=7.21 $Y2=2.075
r130 23 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.125 $Y=2.16
+ $X2=6.75 $Y2=2.16
r131 19 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.585 $Y=2.245
+ $X2=6.585 $Y2=2.16
r132 19 21 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.585 $Y=2.245
+ $X2=6.585 $Y2=2.525
r133 15 36 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.505 $Y=2.075
+ $X2=6.585 $Y2=2.16
r134 15 17 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=6.505 $Y=2.075
+ $X2=6.505 $Y2=0.895
r135 13 43 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.905 $Y=2.315
+ $X2=8.905 $Y2=1.735
r136 9 42 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.725 $Y=0.785
+ $X2=8.725 $Y2=1.405
r137 2 21 600 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_PDIFF $count=1 $X=6.365
+ $Y=2.315 $X2=6.585 $Y2=2.525
r138 1 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.365
+ $Y=0.685 $X2=6.505 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_978_67# 1 2 7 8 11 13 18 19 20 24 25 26
+ 28 29 30 31 33 35 37 38 42 43 46
c132 35 0 1.06469e-20 $X=6.29 $Y=1.87
c133 24 0 1.22987e-19 $X=10.98 $Y=2.56
c134 18 0 2.24221e-19 $X=6.8 $Y=2.525
r135 46 48 8.73685 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.035 $Y=0.545
+ $X2=5.035 $Y2=0.775
r136 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.78
+ $Y=1.48 $X2=5.78 $Y2=1.48
r137 40 42 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=5.752 $Y=1.815
+ $X2=5.752 $Y2=1.48
r138 39 50 3.9577 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=5.2 $Y=1.9
+ $X2=5.075 $Y2=1.98
r139 38 40 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=5.615 $Y=1.9
+ $X2=5.752 $Y2=1.815
r140 38 39 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.615 $Y=1.9
+ $X2=5.2 $Y2=1.9
r141 37 50 3.18546 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.075 $Y=1.815
+ $X2=5.075 $Y2=1.98
r142 37 48 47.9416 $w=2.48e-07 $l=1.04e-06 $layer=LI1_cond $X=5.075 $Y=1.815
+ $X2=5.075 $Y2=0.775
r143 34 43 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=5.78 $Y=1.795
+ $X2=5.78 $Y2=1.48
r144 31 33 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.76 $Y=1.31
+ $X2=11.76 $Y2=1.025
r145 29 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.685 $Y=1.385
+ $X2=11.76 $Y2=1.31
r146 29 30 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=11.685 $Y=1.385
+ $X2=11.48 $Y2=1.385
r147 27 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.405 $Y=1.46
+ $X2=11.48 $Y2=1.385
r148 27 28 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=11.405 $Y=1.46
+ $X2=11.405 $Y2=1.915
r149 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.33 $Y=1.99
+ $X2=11.405 $Y2=1.915
r150 25 26 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=11.33 $Y=1.99
+ $X2=11.055 $Y2=1.99
r151 22 24 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=10.98 $Y=3.075
+ $X2=10.98 $Y2=2.56
r152 21 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.98 $Y=2.065
+ $X2=11.055 $Y2=1.99
r153 21 24 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.98 $Y=2.065
+ $X2=10.98 $Y2=2.56
r154 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.905 $Y=3.15
+ $X2=10.98 $Y2=3.075
r155 19 20 2066.45 $w=1.5e-07 $l=4.03e-06 $layer=POLY_cond $X=10.905 $Y=3.15
+ $X2=6.875 $Y2=3.15
r156 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.8 $Y=3.075
+ $X2=6.875 $Y2=3.15
r157 16 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.8 $Y=3.075
+ $X2=6.8 $Y2=2.525
r158 15 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.8 $Y=1.945
+ $X2=6.8 $Y2=2.525
r159 14 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.365 $Y=1.87
+ $X2=6.29 $Y2=1.87
r160 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.725 $Y=1.87
+ $X2=6.8 $Y2=1.945
r161 13 14 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.725 $Y=1.87
+ $X2=6.365 $Y2=1.87
r162 9 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.29 $Y=1.795
+ $X2=6.29 $Y2=1.87
r163 9 11 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=6.29 $Y=1.795 $X2=6.29
+ $Y2=0.895
r164 8 34 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.945 $Y=1.87
+ $X2=5.78 $Y2=1.795
r165 7 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.215 $Y=1.87
+ $X2=6.29 $Y2=1.87
r166 7 8 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.215 $Y=1.87
+ $X2=5.945 $Y2=1.87
r167 2 50 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=1.835 $X2=5.035 $Y2=1.98
r168 1 46 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.335 $X2=5.035 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_2415_137# 1 2 7 9 14 18 22 24 28 32 34 37
+ 39 40 41 42 43 46 48 50 53 55 56 57 61 65 68 69 72 74 75 79 83 85 86 90 94 96
c206 75 0 1.88236e-20 $X=12.395 $Y=2.125
c207 74 0 1.05354e-19 $X=12.395 $Y=2.125
c208 57 0 8.16742e-20 $X=13.115 $Y=2.205
c209 18 0 1.49913e-19 $X=15.355 $Y=2.465
r210 96 97 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=15.33 $Y=1.38
+ $X2=15.33 $Y2=1.305
r211 91 99 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.33 $Y=1.47
+ $X2=15.33 $Y2=1.635
r212 91 96 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=15.33 $Y=1.47
+ $X2=15.33 $Y2=1.38
r213 90 91 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.33
+ $Y=1.47 $X2=15.33 $Y2=1.47
r214 87 90 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=15.22 $Y=1.47
+ $X2=15.33 $Y2=1.47
r215 84 85 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=13.657 $Y=0.995
+ $X2=13.657 $Y2=1.165
r216 82 83 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=13.28 $Y=2.4
+ $X2=13.28 $Y2=2.475
r217 79 82 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=13.28 $Y=2.205
+ $X2=13.28 $Y2=2.4
r218 75 95 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.395 $Y=2.125
+ $X2=12.395 $Y2=2.29
r219 75 94 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.395 $Y=2.125
+ $X2=12.395 $Y2=1.96
r220 74 77 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=12.395 $Y=2.125
+ $X2=12.395 $Y2=2.205
r221 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.395
+ $Y=2.125 $X2=12.395 $Y2=2.125
r222 71 87 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.22 $Y=1.635
+ $X2=15.22 $Y2=1.47
r223 71 72 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=15.22 $Y=1.635
+ $X2=15.22 $Y2=2.39
r224 70 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.835 $Y=2.475
+ $X2=13.75 $Y2=2.475
r225 69 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.135 $Y=2.475
+ $X2=15.22 $Y2=2.39
r226 69 70 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=15.135 $Y=2.475
+ $X2=13.835 $Y2=2.475
r227 68 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.75 $Y=2.39
+ $X2=13.75 $Y2=2.475
r228 68 85 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=13.75 $Y=2.39
+ $X2=13.75 $Y2=1.165
r229 65 84 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=13.645 $Y=0.815
+ $X2=13.645 $Y2=0.995
r230 62 83 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.445 $Y=2.475
+ $X2=13.28 $Y2=2.475
r231 61 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.665 $Y=2.475
+ $X2=13.75 $Y2=2.475
r232 61 62 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=13.665 $Y=2.475
+ $X2=13.445 $Y2=2.475
r233 58 77 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.56 $Y=2.205
+ $X2=12.395 $Y2=2.205
r234 57 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.115 $Y=2.205
+ $X2=13.28 $Y2=2.205
r235 57 58 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=13.115 $Y=2.205
+ $X2=12.56 $Y2=2.205
r236 51 53 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=12.15 $Y=1.385
+ $X2=12.305 $Y2=1.385
r237 48 50 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=16.805 $Y=1.905
+ $X2=16.805 $Y2=2.3
r238 44 46 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=16.805 $Y=0.795
+ $X2=16.805 $Y2=0.445
r239 42 48 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.73 $Y=1.83
+ $X2=16.805 $Y2=1.905
r240 42 43 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=16.73 $Y=1.83
+ $X2=16.4 $Y2=1.83
r241 40 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.73 $Y=0.87
+ $X2=16.805 $Y2=0.795
r242 40 41 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=16.73 $Y=0.87
+ $X2=16.4 $Y2=0.87
r243 39 43 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.325 $Y=1.755
+ $X2=16.4 $Y2=1.83
r244 38 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.325 $Y=1.455
+ $X2=16.325 $Y2=1.38
r245 38 39 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=16.325 $Y=1.455
+ $X2=16.325 $Y2=1.755
r246 37 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.325 $Y=1.305
+ $X2=16.325 $Y2=1.38
r247 36 41 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.325 $Y=0.945
+ $X2=16.4 $Y2=0.87
r248 36 37 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=16.325 $Y=0.945
+ $X2=16.325 $Y2=1.305
r249 35 55 12.05 $w=1.5e-07 $l=7.8e-08 $layer=POLY_cond $X=15.865 $Y=1.38
+ $X2=15.787 $Y2=1.38
r250 34 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.25 $Y=1.38
+ $X2=16.325 $Y2=1.38
r251 34 35 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=16.25 $Y=1.38
+ $X2=15.865 $Y2=1.38
r252 30 55 12.05 $w=1.5e-07 $l=7.64853e-08 $layer=POLY_cond $X=15.79 $Y=1.305
+ $X2=15.787 $Y2=1.38
r253 30 32 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=15.79 $Y=1.305
+ $X2=15.79 $Y2=0.685
r254 26 55 12.05 $w=1.5e-07 $l=7.59934e-08 $layer=POLY_cond $X=15.785 $Y=1.455
+ $X2=15.787 $Y2=1.38
r255 26 28 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=15.785 $Y=1.455
+ $X2=15.785 $Y2=2.465
r256 25 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.495 $Y=1.38
+ $X2=15.33 $Y2=1.38
r257 24 55 12.05 $w=1.5e-07 $l=7.7e-08 $layer=POLY_cond $X=15.71 $Y=1.38
+ $X2=15.787 $Y2=1.38
r258 24 25 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=15.71 $Y=1.38
+ $X2=15.495 $Y2=1.38
r259 22 97 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=15.36 $Y=0.685
+ $X2=15.36 $Y2=1.305
r260 18 99 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=15.355 $Y=2.465
+ $X2=15.355 $Y2=1.635
r261 14 95 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=12.335 $Y=2.74
+ $X2=12.335 $Y2=2.29
r262 10 53 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.305 $Y=1.46
+ $X2=12.305 $Y2=1.385
r263 10 94 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=12.305 $Y=1.46
+ $X2=12.305 $Y2=1.96
r264 7 51 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.15 $Y=1.31
+ $X2=12.15 $Y2=1.385
r265 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.15 $Y=1.31
+ $X2=12.15 $Y2=1.025
r266 2 82 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=13.14
+ $Y=2.255 $X2=13.28 $Y2=2.4
r267 1 65 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=13.46
+ $Y=0.595 $X2=13.645 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_2211_428# 1 2 9 13 17 20 22 23 26 33 34
c90 22 0 2.25888e-20 $X=11.195 $Y=2.415
c91 13 0 8.16742e-20 $X=13.495 $Y=2.675
r92 34 38 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=13.365 $Y=1.625
+ $X2=13.365 $Y2=1.79
r93 34 37 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=13.365 $Y=1.625
+ $X2=13.365 $Y2=1.46
r94 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.325
+ $Y=1.625 $X2=13.325 $Y2=1.625
r95 30 33 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=13.215 $Y=1.625
+ $X2=13.325 $Y2=1.625
r96 28 29 14.5736 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=11.465 $Y=0.915
+ $X2=11.465 $Y2=1.255
r97 26 28 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=11.465 $Y=0.74
+ $X2=11.465 $Y2=0.915
r98 23 29 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=11.385 $Y=2.12
+ $X2=11.385 $Y2=1.255
r99 22 23 12.2403 $w=4.38e-07 $l=2.95e-07 $layer=LI1_cond $X=11.25 $Y=2.415
+ $X2=11.25 $Y2=2.12
r100 20 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.215 $Y=1.46
+ $X2=13.215 $Y2=1.625
r101 19 20 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=13.215 $Y=1
+ $X2=13.215 $Y2=1.46
r102 18 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.63 $Y=0.915
+ $X2=11.465 $Y2=0.915
r103 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.13 $Y=0.915
+ $X2=13.215 $Y2=1
r104 17 18 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=13.13 $Y=0.915
+ $X2=11.63 $Y2=0.915
r105 13 38 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=13.495 $Y=2.675
+ $X2=13.495 $Y2=1.79
r106 9 37 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=13.385 $Y=0.915
+ $X2=13.385 $Y2=1.46
r107 2 22 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=11.055
+ $Y=2.14 $X2=11.195 $Y2=2.415
r108 1 26 91 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_NDIFF $count=2 $X=11.09
+ $Y=0.595 $X2=11.465 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_1840_21# 1 2 10 13 15 16 20 25 28 30 31
+ 34 35 36 38 44
c110 13 0 1.92809e-19 $X=9.295 $Y=2.315
r111 36 38 13.3683 $w=2.48e-07 $l=2.9e-07 $layer=LI1_cond $X=14.34 $Y=2.085
+ $X2=14.63 $Y2=2.085
r112 35 45 81.7318 $w=5.3e-07 $l=5.05e-07 $layer=POLY_cond $X=14.075 $Y=1.54
+ $X2=14.075 $Y2=2.045
r113 35 44 47.4091 $w=5.3e-07 $l=1.65e-07 $layer=POLY_cond $X=14.075 $Y=1.54
+ $X2=14.075 $Y2=1.375
r114 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.175
+ $Y=1.54 $X2=14.175 $Y2=1.54
r115 32 36 6.96842 $w=2.5e-07 $l=2.16666e-07 $layer=LI1_cond $X=14.177 $Y=1.96
+ $X2=14.34 $Y2=2.085
r116 32 34 14.8931 $w=3.23e-07 $l=4.2e-07 $layer=LI1_cond $X=14.177 $Y=1.96
+ $X2=14.177 $Y2=1.54
r117 31 42 18.1416 $w=3.08e-07 $l=6.02656e-07 $layer=LI1_cond $X=14.177 $Y=1.165
+ $X2=14.635 $Y2=0.83
r118 31 34 13.2974 $w=3.23e-07 $l=3.75e-07 $layer=LI1_cond $X=14.177 $Y=1.165
+ $X2=14.177 $Y2=1.54
r119 30 44 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=13.885 $Y=1.22
+ $X2=13.885 $Y2=1.375
r120 29 30 59.9724 $w=1.75e-07 $l=1.5e-07 $layer=POLY_cond $X=13.872 $Y=1.07
+ $X2=13.872 $Y2=1.22
r121 27 28 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=9.285 $Y=1.18
+ $X2=9.285 $Y2=1.33
r122 25 45 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=13.885 $Y=2.675
+ $X2=13.885 $Y2=2.045
r123 20 29 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=13.86 $Y=0.675
+ $X2=13.86 $Y2=1.07
r124 17 20 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=13.86 $Y=0.255
+ $X2=13.86 $Y2=0.675
r125 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.785 $Y=0.18
+ $X2=13.86 $Y2=0.255
r126 15 16 2274.12 $w=1.5e-07 $l=4.435e-06 $layer=POLY_cond $X=13.785 $Y=0.18
+ $X2=9.35 $Y2=0.18
r127 13 28 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=9.295 $Y=2.315
+ $X2=9.295 $Y2=1.33
r128 10 27 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.275 $Y=0.785
+ $X2=9.275 $Y2=1.18
r129 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.275 $Y=0.255
+ $X2=9.35 $Y2=0.18
r130 7 10 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.275 $Y=0.255
+ $X2=9.275 $Y2=0.785
r131 2 38 600 $w=1.7e-07 $l=3.48999e-07 $layer=licon1_PDIFF $count=1 $X=14.5
+ $Y=1.835 $X2=14.63 $Y2=2.125
r132 1 42 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=14.49
+ $Y=0.685 $X2=14.635 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%RESET_B 1 3 7 9 13
c38 13 0 1.76153e-19 $X=14.755 $Y=1.51
c39 7 0 2.68377e-20 $X=14.85 $Y=0.895
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.755
+ $Y=1.51 $X2=14.755 $Y2=1.51
r41 9 13 4.52224 $w=3.93e-07 $l=1.55e-07 $layer=LI1_cond $X=14.722 $Y=1.665
+ $X2=14.722 $Y2=1.51
r42 5 12 38.6139 $w=3.32e-07 $l=2.06325e-07 $layer=POLY_cond $X=14.85 $Y=1.345
+ $X2=14.757 $Y2=1.51
r43 5 7 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=14.85 $Y=1.345
+ $X2=14.85 $Y2=0.895
r44 1 12 38.6139 $w=3.32e-07 $l=2.04316e-07 $layer=POLY_cond $X=14.845 $Y=1.675
+ $X2=14.757 $Y2=1.51
r45 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=14.845 $Y=1.675
+ $X2=14.845 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_3289_47# 1 2 7 9 12 14 16 18 21 23 26 30
+ 34 37 41
r66 40 41 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=17.315 $Y=1.35
+ $X2=17.39 $Y2=1.35
r67 35 40 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=17.1 $Y=1.35
+ $X2=17.315 $Y2=1.35
r68 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.1
+ $Y=1.35 $X2=17.1 $Y2=1.35
r69 32 37 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=16.755 $Y=1.35
+ $X2=16.59 $Y2=1.35
r70 32 34 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=16.755 $Y=1.35
+ $X2=17.1 $Y2=1.35
r71 28 37 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=16.59 $Y=1.515
+ $X2=16.59 $Y2=1.35
r72 28 30 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=16.59 $Y=1.515
+ $X2=16.59 $Y2=2.125
r73 24 37 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=16.59 $Y=1.185
+ $X2=16.59 $Y2=1.35
r74 24 26 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=16.59 $Y=1.185
+ $X2=16.59 $Y2=0.445
r75 19 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.745 $Y=1.335
+ $X2=17.745 $Y2=1.26
r76 19 21 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=17.745 $Y=1.335
+ $X2=17.745 $Y2=2.465
r77 16 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.745 $Y=1.185
+ $X2=17.745 $Y2=1.26
r78 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=17.745 $Y=1.185
+ $X2=17.745 $Y2=0.655
r79 14 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.67 $Y=1.26
+ $X2=17.745 $Y2=1.26
r80 14 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=17.67 $Y=1.26
+ $X2=17.39 $Y2=1.26
r81 10 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=17.315 $Y=1.515
+ $X2=17.315 $Y2=1.35
r82 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=17.315 $Y=1.515
+ $X2=17.315 $Y2=2.465
r83 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=17.315 $Y=1.185
+ $X2=17.315 $Y2=1.35
r84 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=17.315 $Y=1.185
+ $X2=17.315 $Y2=0.655
r85 2 30 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=16.46
+ $Y=1.98 $X2=16.59 $Y2=2.125
r86 1 26 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=16.445
+ $Y=0.235 $X2=16.59 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_56_481# 1 2 9 11 12 14 15 16 19
c50 11 0 8.92047e-20 $X=1.3 $Y=2.15
r51 17 19 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.325 $Y=2.895
+ $X2=2.325 $Y2=2.55
r52 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.16 $Y=2.98
+ $X2=2.325 $Y2=2.895
r53 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.16 $Y=2.98 $X2=1.47
+ $Y2=2.98
r54 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.385 $Y=2.895
+ $X2=1.47 $Y2=2.98
r55 13 14 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.385 $Y=2.235
+ $X2=1.385 $Y2=2.895
r56 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.3 $Y=2.15
+ $X2=1.385 $Y2=2.235
r57 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.3 $Y=2.15 $X2=0.59
+ $Y2=2.15
r58 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.425 $Y=2.235
+ $X2=0.59 $Y2=2.15
r59 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.425 $Y=2.235
+ $X2=0.425 $Y2=2.55
r60 2 19 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.185
+ $Y=2.405 $X2=2.325 $Y2=2.55
r61 1 9 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=2.405 $X2=0.425 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 39 43 47 51
+ 55 59 63 67 71 75 81 87 89 94 95 97 98 100 101 103 104 106 107 108 123 143 147
+ 152 157 162 167 173 176 179 182 185 188 192
r192 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=3.33 $X2=18
+ $Y2=3.33
r193 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r194 185 186 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r195 182 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r196 179 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r197 176 177 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=12.72
+ $Y=3.33 $X2=12.72 $Y2=3.33
r198 173 174 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r199 171 192 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=3.33
+ $X2=18 $Y2=3.33
r200 171 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=3.33
+ $X2=17.04 $Y2=3.33
r201 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=3.33
+ $X2=17.52 $Y2=3.33
r202 168 188 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.185 $Y=3.33
+ $X2=17.06 $Y2=3.33
r203 168 170 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=17.185 $Y=3.33
+ $X2=17.52 $Y2=3.33
r204 167 191 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=17.875 $Y=3.33
+ $X2=18.057 $Y2=3.33
r205 167 170 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=17.875 $Y=3.33
+ $X2=17.52 $Y2=3.33
r206 166 189 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=17.04 $Y2=3.33
r207 166 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=16.08 $Y2=3.33
r208 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r209 163 185 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.195 $Y=3.33
+ $X2=16.07 $Y2=3.33
r210 163 165 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=16.195 $Y=3.33
+ $X2=16.56 $Y2=3.33
r211 162 188 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.935 $Y=3.33
+ $X2=17.06 $Y2=3.33
r212 162 165 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=16.935 $Y=3.33
+ $X2=16.56 $Y2=3.33
r213 161 186 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.08 $Y2=3.33
r214 161 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=15.12 $Y2=3.33
r215 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r216 158 182 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.305 $Y=3.33
+ $X2=15.14 $Y2=3.33
r217 158 160 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.305 $Y=3.33
+ $X2=15.6 $Y2=3.33
r218 157 185 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.945 $Y=3.33
+ $X2=16.07 $Y2=3.33
r219 157 160 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=15.945 $Y=3.33
+ $X2=15.6 $Y2=3.33
r220 156 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r221 156 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r222 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r223 153 179 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.265 $Y=3.33
+ $X2=14.1 $Y2=3.33
r224 153 155 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=14.265 $Y=3.33
+ $X2=14.64 $Y2=3.33
r225 152 182 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.975 $Y=3.33
+ $X2=15.14 $Y2=3.33
r226 152 155 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.975 $Y=3.33
+ $X2=14.64 $Y2=3.33
r227 151 180 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r228 151 177 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=12.72 $Y2=3.33
r229 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r230 148 176 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.935 $Y=3.33
+ $X2=12.81 $Y2=3.33
r231 148 150 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=12.935 $Y=3.33
+ $X2=13.68 $Y2=3.33
r232 147 179 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.935 $Y=3.33
+ $X2=14.1 $Y2=3.33
r233 147 150 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=13.935 $Y=3.33
+ $X2=13.68 $Y2=3.33
r234 146 177 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=12.72 $Y2=3.33
r235 145 146 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r236 143 176 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.685 $Y=3.33
+ $X2=12.81 $Y2=3.33
r237 143 145 185.61 $w=1.68e-07 $l=2.845e-06 $layer=LI1_cond $X=12.685 $Y=3.33
+ $X2=9.84 $Y2=3.33
r238 142 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r239 141 142 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r240 138 141 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r241 138 139 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r242 136 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r243 135 136 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r244 133 136 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r245 133 174 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r246 132 135 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r247 132 133 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r248 130 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.69 $Y=3.33
+ $X2=5.525 $Y2=3.33
r249 130 132 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.69 $Y=3.33
+ $X2=6 $Y2=3.33
r250 129 174 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r251 128 129 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r252 126 129 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r253 125 128 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r254 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r255 123 173 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.36 $Y=3.33
+ $X2=5.525 $Y2=3.33
r256 123 128 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.36 $Y=3.33
+ $X2=5.04 $Y2=3.33
r257 122 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r258 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r259 119 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r260 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r261 116 119 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r262 115 118 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r263 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r264 112 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r265 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r266 108 142 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=9.36 $Y2=3.33
r267 108 139 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=8.4 $Y2=3.33
r268 107 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.675 $Y=3.33
+ $X2=9.84 $Y2=3.33
r269 106 141 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=9.51 $Y=3.33
+ $X2=9.36 $Y2=3.33
r270 106 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.51 $Y=3.33
+ $X2=9.675 $Y2=3.33
r271 103 135 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.955 $Y=3.33
+ $X2=7.92 $Y2=3.33
r272 103 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.955 $Y=3.33
+ $X2=8.12 $Y2=3.33
r273 102 138 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.285 $Y=3.33
+ $X2=8.4 $Y2=3.33
r274 102 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.285 $Y=3.33
+ $X2=8.12 $Y2=3.33
r275 100 121 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.6 $Y2=3.33
r276 100 101 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.77 $Y2=3.33
r277 99 125 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.895 $Y=3.33
+ $X2=4.08 $Y2=3.33
r278 99 101 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.895 $Y=3.33
+ $X2=3.77 $Y2=3.33
r279 97 118 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r280 97 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.72 $Y=3.33
+ $X2=2.885 $Y2=3.33
r281 96 121 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=3.6 $Y2=3.33
r282 96 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=2.885 $Y2=3.33
r283 94 111 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.77 $Y=3.33
+ $X2=0.72 $Y2=3.33
r284 94 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=3.33
+ $X2=0.935 $Y2=3.33
r285 93 115 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=1.2
+ $Y2=3.33
r286 93 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=0.935 $Y2=3.33
r287 89 92 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=18 $Y=1.98 $X2=18
+ $Y2=2.95
r288 87 191 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=18 $Y=3.245
+ $X2=18.057 $Y2=3.33
r289 87 92 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=18 $Y=3.245 $X2=18
+ $Y2=2.95
r290 84 86 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=17.06 $Y=2.465
+ $X2=17.06 $Y2=2.95
r291 81 84 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=17.06 $Y=1.98
+ $X2=17.06 $Y2=2.465
r292 79 188 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=17.06 $Y=3.245
+ $X2=17.06 $Y2=3.33
r293 79 86 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=17.06 $Y=3.245
+ $X2=17.06 $Y2=2.95
r294 75 78 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=16.07 $Y=1.98
+ $X2=16.07 $Y2=2.95
r295 73 185 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.07 $Y=3.245
+ $X2=16.07 $Y2=3.33
r296 73 78 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=16.07 $Y=3.245
+ $X2=16.07 $Y2=2.95
r297 69 182 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.14 $Y=3.245
+ $X2=15.14 $Y2=3.33
r298 69 71 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=15.14 $Y=3.245
+ $X2=15.14 $Y2=2.925
r299 65 179 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.1 $Y=3.245
+ $X2=14.1 $Y2=3.33
r300 65 67 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=14.1 $Y=3.245
+ $X2=14.1 $Y2=2.925
r301 61 176 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.81 $Y=3.245
+ $X2=12.81 $Y2=3.33
r302 61 63 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=12.81 $Y=3.245
+ $X2=12.81 $Y2=2.79
r303 57 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.675 $Y=3.245
+ $X2=9.675 $Y2=3.33
r304 57 59 42.0816 $w=3.28e-07 $l=1.205e-06 $layer=LI1_cond $X=9.675 $Y=3.245
+ $X2=9.675 $Y2=2.04
r305 53 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.12 $Y=3.245
+ $X2=8.12 $Y2=3.33
r306 53 55 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=8.12 $Y=3.245
+ $X2=8.12 $Y2=2.59
r307 49 173 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.525 $Y=3.245
+ $X2=5.525 $Y2=3.33
r308 49 51 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=5.525 $Y=3.245
+ $X2=5.525 $Y2=2.84
r309 45 101 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=3.245
+ $X2=3.77 $Y2=3.33
r310 45 47 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=3.77 $Y=3.245
+ $X2=3.77 $Y2=2.55
r311 41 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=3.245
+ $X2=2.885 $Y2=3.33
r312 41 43 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=2.885 $Y=3.245
+ $X2=2.885 $Y2=2.59
r313 37 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=3.245
+ $X2=0.935 $Y2=3.33
r314 37 39 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=0.935 $Y=3.245
+ $X2=0.935 $Y2=2.74
r315 12 92 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=17.82
+ $Y=1.835 $X2=17.96 $Y2=2.95
r316 12 89 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=17.82
+ $Y=1.835 $X2=17.96 $Y2=1.98
r317 11 86 600 $w=1.7e-07 $l=1.07438e-06 $layer=licon1_PDIFF $count=1 $X=16.88
+ $Y=1.98 $X2=17.1 $Y2=2.95
r318 11 84 600 $w=1.7e-07 $l=5.84744e-07 $layer=licon1_PDIFF $count=1 $X=16.88
+ $Y=1.98 $X2=17.1 $Y2=2.465
r319 11 81 600 $w=1.7e-07 $l=2.2e-07 $layer=licon1_PDIFF $count=1 $X=16.88
+ $Y=1.98 $X2=17.1 $Y2=1.98
r320 10 78 400 $w=1.7e-07 $l=1.19699e-06 $layer=licon1_PDIFF $count=1 $X=15.86
+ $Y=1.835 $X2=16.03 $Y2=2.95
r321 10 75 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=15.86
+ $Y=1.835 $X2=16.03 $Y2=1.98
r322 9 71 600 $w=1.7e-07 $l=1.19495e-06 $layer=licon1_PDIFF $count=1 $X=14.92
+ $Y=1.835 $X2=15.14 $Y2=2.925
r323 8 67 600 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=1 $X=13.96
+ $Y=2.255 $X2=14.1 $Y2=2.925
r324 7 63 600 $w=1.7e-07 $l=5.54977e-07 $layer=licon1_PDIFF $count=1 $X=12.41
+ $Y=2.53 $X2=12.85 $Y2=2.79
r325 6 59 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=9.37
+ $Y=1.895 $X2=9.675 $Y2=2.04
r326 5 55 600 $w=1.7e-07 $l=9.82929e-07 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=2.315 $X2=8.12 $Y2=2.59
r327 4 51 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=2.345 $X2=5.525 $Y2=2.84
r328 3 47 600 $w=1.7e-07 $l=5.56215e-07 $layer=licon1_PDIFF $count=1 $X=3.68
+ $Y=2.055 $X2=3.81 $Y2=2.55
r329 2 43 600 $w=1.7e-07 $l=1.12517e-06 $layer=licon1_PDIFF $count=1 $X=2.74
+ $Y=1.535 $X2=2.885 $Y2=2.59
r330 1 39 600 $w=1.7e-07 $l=4.3119e-07 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=2.405 $X2=0.935 $Y2=2.74
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_202_119# 1 2 3 4 15 17 18 21 24 25 28 29
+ 30 32 34 36 37 39 44 45
c138 45 0 1.52322e-19 $X=6.155 $Y=2.525
c139 44 0 1.28128e-19 $X=5.91 $Y=2.525
c140 34 0 1.58976e-19 $X=5.18 $Y=2.41
r141 43 45 2.08014 $w=4.58e-07 $l=8e-08 $layer=LI1_cond $X=6.075 $Y=2.525
+ $X2=6.155 $Y2=2.525
r142 43 44 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.075 $Y=2.525
+ $X2=5.91 $Y2=2.525
r143 39 41 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6.075 $Y=0.895
+ $X2=6.075 $Y2=1.125
r144 36 45 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=6.155 $Y=2.295
+ $X2=6.155 $Y2=2.525
r145 36 41 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=6.155 $Y=2.295
+ $X2=6.155 $Y2=1.125
r146 34 44 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.18 $Y=2.41
+ $X2=5.91 $Y2=2.41
r147 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.095 $Y=2.495
+ $X2=5.18 $Y2=2.41
r148 31 32 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.095 $Y=2.495
+ $X2=5.095 $Y2=2.895
r149 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.01 $Y=2.98
+ $X2=5.095 $Y2=2.895
r150 29 30 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.01 $Y=2.98
+ $X2=4.245 $Y2=2.98
r151 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.16 $Y=2.895
+ $X2=4.245 $Y2=2.98
r152 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.16 $Y=2.205
+ $X2=4.16 $Y2=2.895
r153 26 37 2.76166 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=2.145 $Y=2.12
+ $X2=1.897 $Y2=2.12
r154 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.075 $Y=2.12
+ $X2=4.16 $Y2=2.205
r155 25 26 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=4.075 $Y=2.12
+ $X2=2.145 $Y2=2.12
r156 24 37 3.70735 $w=2.5e-07 $l=2.01057e-07 $layer=LI1_cond $X=2.06 $Y=2.035
+ $X2=1.897 $Y2=2.12
r157 23 24 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.06 $Y=0.63
+ $X2=2.06 $Y2=2.035
r158 19 37 3.70735 $w=2.5e-07 $l=1.19143e-07 $layer=LI1_cond $X=1.815 $Y=2.205
+ $X2=1.897 $Y2=2.12
r159 19 21 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.815 $Y=2.205
+ $X2=1.815 $Y2=2.59
r160 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.975 $Y=0.545
+ $X2=2.06 $Y2=0.63
r161 17 18 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.975 $Y=0.545
+ $X2=1.315 $Y2=0.545
r162 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.15 $Y=0.63
+ $X2=1.315 $Y2=0.545
r163 13 15 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.15 $Y=0.63
+ $X2=1.15 $Y2=0.805
r164 4 43 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=5.945
+ $Y=2.315 $X2=6.075 $Y2=2.525
r165 3 21 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=1.615
+ $Y=2.405 $X2=1.815 $Y2=2.59
r166 2 39 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=5.945
+ $Y=0.685 $X2=6.075 $Y2=0.895
r167 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.595 $X2=1.15 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%Q_N 1 2 9 13 14 15 16 24 34
c39 34 0 5.30782e-20 $X=15.625 $Y=1.815
r40 21 24 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=15.625 $Y=1.955
+ $X2=15.625 $Y2=1.98
r41 16 31 5.14483 $w=2.78e-07 $l=1.25e-07 $layer=LI1_cond $X=15.625 $Y=2.775
+ $X2=15.625 $Y2=2.9
r42 15 16 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=15.625 $Y=2.405
+ $X2=15.625 $Y2=2.775
r43 14 21 0.123476 $w=2.78e-07 $l=3e-09 $layer=LI1_cond $X=15.625 $Y=1.952
+ $X2=15.625 $Y2=1.955
r44 14 34 7.40445 $w=2.78e-07 $l=1.37e-07 $layer=LI1_cond $X=15.625 $Y=1.952
+ $X2=15.625 $Y2=1.815
r45 14 15 15.1464 $w=2.78e-07 $l=3.68e-07 $layer=LI1_cond $X=15.625 $Y=2.037
+ $X2=15.625 $Y2=2.405
r46 14 24 2.34604 $w=2.78e-07 $l=5.7e-08 $layer=LI1_cond $X=15.625 $Y=2.037
+ $X2=15.625 $Y2=1.98
r47 13 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=15.68 $Y=1.125
+ $X2=15.68 $Y2=1.815
r48 7 13 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=15.587 $Y=0.948
+ $X2=15.587 $Y2=1.125
r49 7 9 16.8159 $w=3.53e-07 $l=5.18e-07 $layer=LI1_cond $X=15.587 $Y=0.948
+ $X2=15.587 $Y2=0.43
r50 2 31 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=15.43
+ $Y=1.835 $X2=15.57 $Y2=2.9
r51 2 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.43
+ $Y=1.835 $X2=15.57 $Y2=1.98
r52 1 9 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=15.435
+ $Y=0.265 $X2=15.575 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%Q 1 2 7 8 9 10 11 12 13 22
r20 13 40 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=17.53 $Y=2.775
+ $X2=17.53 $Y2=2.9
r21 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.53 $Y=2.405
+ $X2=17.53 $Y2=2.775
r22 11 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=17.53 $Y=1.98
+ $X2=17.53 $Y2=2.405
r23 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=17.53 $Y=1.665
+ $X2=17.53 $Y2=1.98
r24 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.53 $Y=1.295
+ $X2=17.53 $Y2=1.665
r25 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.53 $Y=0.925
+ $X2=17.53 $Y2=1.295
r26 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=17.53 $Y=0.555
+ $X2=17.53 $Y2=0.925
r27 7 22 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=17.53 $Y=0.555
+ $X2=17.53 $Y2=0.43
r28 2 40 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=17.39
+ $Y=1.835 $X2=17.53 $Y2=2.9
r29 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=17.39
+ $Y=1.835 $X2=17.53 $Y2=1.98
r30 1 22 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=17.39
+ $Y=0.235 $X2=17.53 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%VGND 1 2 3 4 5 6 7 8 9 10 11 34 36 40 44 48
+ 52 56 60 64 70 74 78 80 83 84 86 87 89 90 91 93 105 119 133 140 145 150 159
+ 162 165 168 171 174 178
r185 177 178 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=0 $X2=18
+ $Y2=0
r186 174 175 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=0
+ $X2=17.04 $Y2=0
r187 171 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r188 168 169 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r189 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r190 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r191 159 160 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r192 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r193 154 178 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=0
+ $X2=18 $Y2=0
r194 154 175 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.52 $Y=0
+ $X2=17.04 $Y2=0
r195 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r196 151 174 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.185 $Y=0
+ $X2=17.06 $Y2=0
r197 151 153 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=17.185 $Y=0
+ $X2=17.52 $Y2=0
r198 150 177 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=17.875 $Y=0
+ $X2=18.057 $Y2=0
r199 150 153 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=17.875 $Y=0
+ $X2=17.52 $Y2=0
r200 149 175 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=17.04 $Y2=0
r201 149 172 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=16.08 $Y2=0
r202 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r203 146 171 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.195 $Y=0
+ $X2=16.07 $Y2=0
r204 146 148 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=16.195 $Y=0
+ $X2=16.56 $Y2=0
r205 145 174 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.935 $Y=0
+ $X2=17.06 $Y2=0
r206 145 148 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=16.935 $Y=0
+ $X2=16.56 $Y2=0
r207 144 172 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.08 $Y2=0
r208 144 169 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=15.12 $Y2=0
r209 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r210 141 168 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.23 $Y=0
+ $X2=15.105 $Y2=0
r211 141 143 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=15.23 $Y=0
+ $X2=15.6 $Y2=0
r212 140 171 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.945 $Y=0
+ $X2=16.07 $Y2=0
r213 140 143 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=15.945 $Y=0
+ $X2=15.6 $Y2=0
r214 139 169 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r215 138 139 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r216 136 139 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=14.64 $Y2=0
r217 135 138 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=12.72 $Y=0
+ $X2=14.64 $Y2=0
r218 135 136 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r219 133 168 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.98 $Y=0
+ $X2=15.105 $Y2=0
r220 133 138 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=14.98 $Y=0
+ $X2=14.64 $Y2=0
r221 132 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r222 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r223 129 132 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=12.24 $Y2=0
r224 129 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r225 128 131 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=10.8 $Y=0
+ $X2=12.24 $Y2=0
r226 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r227 126 165 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.455 $Y=0
+ $X2=10.33 $Y2=0
r228 126 128 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.455 $Y=0
+ $X2=10.8 $Y2=0
r229 125 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r230 124 125 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r231 121 124 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r232 121 122 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r233 119 165 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.205 $Y=0
+ $X2=10.33 $Y2=0
r234 119 124 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=10.205 $Y=0
+ $X2=9.84 $Y2=0
r235 118 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r236 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r237 115 118 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=0 $X2=7.44
+ $Y2=0
r238 115 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r239 114 117 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=0 $X2=7.44
+ $Y2=0
r240 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r241 112 162 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.71 $Y=0
+ $X2=5.545 $Y2=0
r242 112 114 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.71 $Y=0 $X2=6
+ $Y2=0
r243 111 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r244 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r245 108 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r246 107 110 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r247 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r248 105 162 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.38 $Y=0
+ $X2=5.545 $Y2=0
r249 105 110 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.38 $Y=0
+ $X2=5.04 $Y2=0
r250 104 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.08 $Y2=0
r251 104 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=2.64 $Y2=0
r252 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r253 101 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=0
+ $X2=2.49 $Y2=0
r254 101 103 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=2.655 $Y=0
+ $X2=3.6 $Y2=0
r255 100 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r256 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r257 97 100 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=2.16 $Y2=0
r258 97 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r259 96 99 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r260 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r261 94 156 4.62984 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=0.495 $Y=0
+ $X2=0.247 $Y2=0
r262 94 96 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.495 $Y=0
+ $X2=0.72 $Y2=0
r263 93 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0
+ $X2=2.49 $Y2=0
r264 93 99 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0
+ $X2=2.16 $Y2=0
r265 91 125 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=9.84 $Y2=0
r266 91 122 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=7.92 $Y2=0
r267 89 131 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=12.335 $Y=0
+ $X2=12.24 $Y2=0
r268 89 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.335 $Y=0
+ $X2=12.5 $Y2=0
r269 88 135 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=12.665 $Y=0
+ $X2=12.72 $Y2=0
r270 88 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.665 $Y=0
+ $X2=12.5 $Y2=0
r271 86 117 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.465 $Y=0
+ $X2=7.44 $Y2=0
r272 86 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.465 $Y=0 $X2=7.63
+ $Y2=0
r273 85 121 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.795 $Y=0
+ $X2=7.92 $Y2=0
r274 85 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=0 $X2=7.63
+ $Y2=0
r275 83 103 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.6
+ $Y2=0
r276 83 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.83
+ $Y2=0
r277 82 107 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=0
+ $X2=4.08 $Y2=0
r278 82 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.83
+ $Y2=0
r279 78 177 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=18 $Y=0.085
+ $X2=18.057 $Y2=0
r280 78 80 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=18 $Y=0.085 $X2=18
+ $Y2=0.38
r281 74 76 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=17.06 $Y=0.38
+ $X2=17.06 $Y2=0.84
r282 72 174 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=17.06 $Y=0.085
+ $X2=17.06 $Y2=0
r283 72 74 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=17.06 $Y=0.085
+ $X2=17.06 $Y2=0.38
r284 68 171 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.07 $Y=0.085
+ $X2=16.07 $Y2=0
r285 68 70 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=16.07 $Y=0.085
+ $X2=16.07 $Y2=0.41
r286 64 66 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=15.105 $Y=0.41
+ $X2=15.105 $Y2=0.96
r287 62 168 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.105 $Y=0.085
+ $X2=15.105 $Y2=0
r288 62 64 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=15.105 $Y=0.085
+ $X2=15.105 $Y2=0.41
r289 58 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.5 $Y=0.085
+ $X2=12.5 $Y2=0
r290 58 60 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=12.5 $Y=0.085 $X2=12.5
+ $Y2=0.485
r291 54 165 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.33 $Y=0.085
+ $X2=10.33 $Y2=0
r292 54 56 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=10.33 $Y=0.085
+ $X2=10.33 $Y2=0.745
r293 50 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.63 $Y=0.085
+ $X2=7.63 $Y2=0
r294 50 52 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=7.63 $Y=0.085 $X2=7.63
+ $Y2=0.485
r295 46 162 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.545 $Y=0.085
+ $X2=5.545 $Y2=0
r296 46 48 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=5.545 $Y=0.085
+ $X2=5.545 $Y2=0.545
r297 42 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0
r298 42 44 20.9535 $w=3.28e-07 $l=6e-07 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0.685
r299 38 159 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0
r300 38 40 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0.79
r301 34 156 3.13634 $w=3.3e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.247 $Y2=0
r302 34 36 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.33 $Y2=0.805
r303 11 80 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=17.82
+ $Y=0.235 $X2=17.96 $Y2=0.38
r304 10 76 182 $w=1.7e-07 $l=7.06488e-07 $layer=licon1_NDIFF $count=1 $X=16.88
+ $Y=0.235 $X2=17.1 $Y2=0.84
r305 10 74 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=16.88
+ $Y=0.235 $X2=17.1 $Y2=0.38
r306 9 70 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=15.865
+ $Y=0.265 $X2=16.03 $Y2=0.41
r307 8 66 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=14.925
+ $Y=0.685 $X2=15.145 $Y2=0.96
r308 8 64 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=14.925
+ $Y=0.685 $X2=15.145 $Y2=0.41
r309 7 60 182 $w=1.7e-07 $l=4.46822e-07 $layer=licon1_NDIFF $count=1 $X=12.225
+ $Y=0.815 $X2=12.5 $Y2=0.485
r310 6 56 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=10.145
+ $Y=0.595 $X2=10.29 $Y2=0.745
r311 5 52 182 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_NDIFF $count=1 $X=7.41
+ $Y=0.685 $X2=7.63 $Y2=0.485
r312 4 48 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=5.385
+ $Y=0.335 $X2=5.545 $Y2=0.545
r313 3 44 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.685
+ $Y=0.475 $X2=3.83 $Y2=0.685
r314 2 40 182 $w=1.7e-07 $l=3.90512e-07 $layer=licon1_NDIFF $count=1 $X=2.185
+ $Y=0.595 $X2=2.49 $Y2=0.79
r315 1 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.595 $X2=0.33 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_1670_93# 1 2 7 9 14
c22 7 0 3.17754e-19 $X=9.345 $Y=0.7
r23 14 17 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=9.51 $Y=0.7 $X2=9.51
+ $Y2=0.785
r24 9 12 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=8.49 $Y=0.7 $X2=8.49
+ $Y2=0.805
r25 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.655 $Y=0.7 $X2=8.49
+ $Y2=0.7
r26 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.345 $Y=0.7 $X2=9.51
+ $Y2=0.7
r27 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.345 $Y=0.7 $X2=8.655
+ $Y2=0.7
r28 2 17 182 $w=1.7e-07 $l=3.91918e-07 $layer=licon1_NDIFF $count=1 $X=9.35
+ $Y=0.465 $X2=9.51 $Y2=0.785
r29 1 12 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=8.35
+ $Y=0.465 $X2=8.49 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBN_2%A_2574_119# 1 2 7 11 13
r26 13 16 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=13.09 $Y=0.35
+ $X2=13.09 $Y2=0.485
r27 9 11 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=14.115 $Y=0.435
+ $X2=14.115 $Y2=0.575
r28 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.255 $Y=0.35
+ $X2=13.09 $Y2=0.35
r29 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.99 $Y=0.35
+ $X2=14.115 $Y2=0.435
r30 7 8 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=13.99 $Y=0.35
+ $X2=13.255 $Y2=0.35
r31 2 11 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=13.935
+ $Y=0.355 $X2=14.075 $Y2=0.575
r32 1 16 182 $w=1.7e-07 $l=2.69444e-07 $layer=licon1_NDIFF $count=1 $X=12.87
+ $Y=0.595 $X2=13.09 $Y2=0.485
.ends

