* File: sky130_fd_sc_lp__nand2_2.pxi.spice
* Created: Wed Sep  2 10:02:43 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2_2%B N_B_M1001_g N_B_M1003_g N_B_M1005_g N_B_M1006_g
+ B B N_B_c_46_n PM_SKY130_FD_SC_LP__NAND2_2%B
x_PM_SKY130_FD_SC_LP__NAND2_2%A N_A_M1002_g N_A_M1000_g N_A_M1007_g N_A_M1004_g
+ A A N_A_c_86_n PM_SKY130_FD_SC_LP__NAND2_2%A
x_PM_SKY130_FD_SC_LP__NAND2_2%VPWR N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_M1004_s
+ N_VPWR_c_131_n N_VPWR_c_132_n N_VPWR_c_133_n N_VPWR_c_134_n N_VPWR_c_135_n
+ VPWR N_VPWR_c_136_n N_VPWR_c_137_n N_VPWR_c_138_n N_VPWR_c_130_n
+ PM_SKY130_FD_SC_LP__NAND2_2%VPWR
x_PM_SKY130_FD_SC_LP__NAND2_2%Y N_Y_M1002_d N_Y_M1003_s N_Y_M1000_d N_Y_c_173_n
+ N_Y_c_195_n N_Y_c_175_n N_Y_c_179_n N_Y_c_199_n N_Y_c_171_n N_Y_c_168_n
+ N_Y_c_169_n N_Y_c_189_n Y PM_SKY130_FD_SC_LP__NAND2_2%Y
x_PM_SKY130_FD_SC_LP__NAND2_2%A_27_65# N_A_27_65#_M1001_d N_A_27_65#_M1005_d
+ N_A_27_65#_M1007_s N_A_27_65#_c_211_n N_A_27_65#_c_212_n N_A_27_65#_c_213_n
+ N_A_27_65#_c_214_n N_A_27_65#_c_215_n N_A_27_65#_c_216_n
+ PM_SKY130_FD_SC_LP__NAND2_2%A_27_65#
x_PM_SKY130_FD_SC_LP__NAND2_2%VGND N_VGND_M1001_s N_VGND_c_245_n VGND
+ N_VGND_c_246_n N_VGND_c_247_n N_VGND_c_248_n N_VGND_c_249_n
+ PM_SKY130_FD_SC_LP__NAND2_2%VGND
cc_1 VNB N_B_M1001_g 0.0262168f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.745
cc_2 VNB N_B_M1005_g 0.0194982f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.745
cc_3 VNB B 0.0141308f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_B_c_46_n 0.0381828f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.51
cc_5 VNB N_A_M1002_g 0.0198596f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.745
cc_6 VNB N_A_M1007_g 0.023346f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.745
cc_7 VNB A 0.00446349f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_A_c_86_n 0.033906f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.51
cc_9 VNB N_VPWR_c_130_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_Y_c_168_n 0.014502f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.51
cc_11 VNB N_Y_c_169_n 0.00228591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB Y 0.0227708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_65#_c_211_n 0.0312591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_65#_c_212_n 0.00626417f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_15 VNB N_A_27_65#_c_213_n 0.00985882f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_16 VNB N_A_27_65#_c_214_n 0.0127794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_65#_c_215_n 0.00171451f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_18 VNB N_A_27_65#_c_216_n 0.0181406f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.51
cc_19 VNB N_VGND_c_245_n 0.00280617f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_20 VNB N_VGND_c_246_n 0.0161944f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.745
cc_21 VNB N_VGND_c_247_n 0.0398879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_248_n 0.163532f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_23 VNB N_VGND_c_249_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.51
cc_24 VPB N_B_M1003_g 0.0235869f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_25 VPB N_B_M1006_g 0.0185012f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_26 VPB B 0.0114172f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_27 VPB N_B_c_46_n 0.00505318f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.51
cc_28 VPB N_A_M1000_g 0.0180979f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_29 VPB N_A_M1004_g 0.0209722f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_30 VPB A 0.00465098f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_31 VPB N_A_c_86_n 0.00486532f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.51
cc_32 VPB N_VPWR_c_131_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.745
cc_33 VPB N_VPWR_c_132_n 0.0481737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_133_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_35 VPB N_VPWR_c_134_n 0.0154435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_135_n 0.0352012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_136_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.51
cc_38 VPB N_VPWR_c_137_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.582
cc_39 VPB N_VPWR_c_138_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_130_n 0.0499569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_Y_c_171_n 0.0152982f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.51
cc_42 VPB Y 0.0138034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 N_B_M1005_g N_A_M1002_g 0.0242562f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_44 N_B_M1006_g N_A_M1000_g 0.0242562f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_45 B A 0.0296441f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_46 N_B_c_46_n A 0.00268875f $X=0.905 $Y=1.51 $X2=0 $Y2=0
cc_47 B N_A_c_86_n 2.94915e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_48 N_B_c_46_n N_A_c_86_n 0.0242562f $X=0.905 $Y=1.51 $X2=0 $Y2=0
cc_49 N_B_M1003_g N_VPWR_c_132_n 0.0186161f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_50 N_B_M1006_g N_VPWR_c_132_n 7.28867e-19 $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_51 B N_VPWR_c_132_n 0.0252291f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_52 N_B_M1003_g N_VPWR_c_133_n 6.77662e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_53 N_B_M1006_g N_VPWR_c_133_n 0.0143066f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_54 N_B_M1003_g N_VPWR_c_136_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_55 N_B_M1006_g N_VPWR_c_136_n 0.00486043f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_56 N_B_M1003_g N_VPWR_c_130_n 0.00824727f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_57 N_B_M1006_g N_VPWR_c_130_n 0.00824727f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_58 B N_Y_c_173_n 0.0154121f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_59 N_B_c_46_n N_Y_c_173_n 6.52992e-19 $X=0.905 $Y=1.51 $X2=0 $Y2=0
cc_60 N_B_M1006_g N_Y_c_175_n 0.0129876f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_61 B N_Y_c_175_n 0.00899385f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_62 N_B_M1001_g N_A_27_65#_c_211_n 0.00354556f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_63 N_B_M1001_g N_A_27_65#_c_212_n 0.0138099f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_64 N_B_M1005_g N_A_27_65#_c_212_n 0.0137533f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_65 B N_A_27_65#_c_212_n 0.0424795f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_66 N_B_c_46_n N_A_27_65#_c_212_n 0.00243542f $X=0.905 $Y=1.51 $X2=0 $Y2=0
cc_67 B N_A_27_65#_c_213_n 0.0230248f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_68 N_B_M1005_g N_A_27_65#_c_215_n 4.93056e-19 $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_69 N_B_M1001_g N_VGND_c_245_n 0.0124264f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_70 N_B_M1005_g N_VGND_c_245_n 0.0103937f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_71 N_B_M1001_g N_VGND_c_246_n 0.00414769f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_72 N_B_M1005_g N_VGND_c_247_n 0.00414769f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_73 N_B_M1001_g N_VGND_c_248_n 0.00823375f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_74 N_B_M1005_g N_VGND_c_248_n 0.0078848f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_VPWR_c_133_n 0.0143066f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_76 N_A_M1004_g N_VPWR_c_133_n 6.77662e-19 $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A_M1000_g N_VPWR_c_135_n 6.80491e-19 $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_VPWR_c_135_n 0.0168603f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A_M1000_g N_VPWR_c_137_n 0.00486043f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A_M1004_g N_VPWR_c_137_n 0.00486043f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_81 N_A_M1000_g N_VPWR_c_130_n 0.00824727f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A_M1004_g N_VPWR_c_130_n 0.00824727f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A_M1000_g N_Y_c_175_n 0.0122227f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_84 A N_Y_c_175_n 0.0229862f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_85 N_A_M1002_g N_Y_c_179_n 0.00517467f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_86 N_A_M1007_g N_Y_c_179_n 0.0112499f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_87 N_A_M1004_g N_Y_c_171_n 0.0141385f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_88 A N_Y_c_171_n 0.0118538f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_M1007_g N_Y_c_168_n 0.0110435f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_90 A N_Y_c_168_n 0.0081885f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_Y_c_169_n 0.0030426f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_92 N_A_M1007_g N_Y_c_169_n 0.0016823f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_93 A N_Y_c_169_n 0.0274989f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_94 N_A_c_86_n N_Y_c_169_n 0.00252688f $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_95 A N_Y_c_189_n 0.0154121f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_96 N_A_c_86_n N_Y_c_189_n 6.52992e-19 $X=1.765 $Y=1.51 $X2=0 $Y2=0
cc_97 N_A_M1007_g Y 0.0212269f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_98 A Y 0.0277703f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_99 N_A_M1002_g N_A_27_65#_c_212_n 6.57126e-19 $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_100 A N_A_27_65#_c_212_n 0.00929846f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A_M1002_g N_A_27_65#_c_214_n 0.0117775f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_102 N_A_M1007_g N_A_27_65#_c_214_n 0.0127933f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_103 N_A_M1002_g N_VGND_c_245_n 5.62244e-19 $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_104 N_A_M1002_g N_VGND_c_247_n 0.0030414f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_105 N_A_M1007_g N_VGND_c_247_n 0.0030414f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_106 N_A_M1002_g N_VGND_c_248_n 0.00435814f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_107 N_A_M1007_g N_VGND_c_248_n 0.00475332f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_108 N_VPWR_c_130_n N_Y_M1003_s 0.00536646f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_109 N_VPWR_c_130_n N_Y_M1000_d 0.00536646f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_110 N_VPWR_c_136_n N_Y_c_195_n 0.0124525f $X=0.955 $Y=3.33 $X2=0 $Y2=0
cc_111 N_VPWR_c_130_n N_Y_c_195_n 0.00730901f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_112 N_VPWR_M1006_d N_Y_c_175_n 0.00423879f $X=0.98 $Y=1.835 $X2=0 $Y2=0
cc_113 N_VPWR_c_133_n N_Y_c_175_n 0.0163515f $X=1.12 $Y=2.4 $X2=0 $Y2=0
cc_114 N_VPWR_c_137_n N_Y_c_199_n 0.0124525f $X=1.815 $Y=3.33 $X2=0 $Y2=0
cc_115 N_VPWR_c_130_n N_Y_c_199_n 0.00730901f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_116 N_VPWR_M1004_s N_Y_c_171_n 0.00508822f $X=1.84 $Y=1.835 $X2=0 $Y2=0
cc_117 N_VPWR_c_135_n N_Y_c_171_n 0.0232056f $X=1.98 $Y=2.4 $X2=0 $Y2=0
cc_118 N_VPWR_M1004_s Y 0.00143604f $X=1.84 $Y=1.835 $X2=0 $Y2=0
cc_119 N_Y_c_168_n N_A_27_65#_M1007_s 0.00403f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_120 N_Y_c_175_n N_A_27_65#_c_212_n 0.00380868f $X=1.455 $Y=2.005 $X2=0 $Y2=0
cc_121 N_Y_c_169_n N_A_27_65#_c_212_n 0.0104195f $X=1.715 $Y=1.16 $X2=0 $Y2=0
cc_122 N_Y_M1002_d N_A_27_65#_c_214_n 0.00176461f $X=1.41 $Y=0.325 $X2=0 $Y2=0
cc_123 N_Y_c_179_n N_A_27_65#_c_214_n 0.0159398f $X=1.55 $Y=0.69 $X2=0 $Y2=0
cc_124 N_Y_c_168_n N_A_27_65#_c_214_n 0.00280043f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_125 N_Y_c_168_n N_A_27_65#_c_216_n 0.0273201f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_27_65#_c_212_n N_VGND_M1001_s 0.00176461f $X=1.035 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_27_65#_c_211_n N_VGND_c_245_n 0.0232759f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A_27_65#_c_212_n N_VGND_c_245_n 0.0170777f $X=1.035 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_27_65#_c_215_n N_VGND_c_245_n 0.00876136f $X=1.205 $Y=0.35 $X2=0
+ $Y2=0
cc_130 N_A_27_65#_c_211_n N_VGND_c_246_n 0.0140356f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_131 N_A_27_65#_c_214_n N_VGND_c_247_n 0.063047f $X=1.895 $Y=0.35 $X2=0 $Y2=0
cc_132 N_A_27_65#_c_215_n N_VGND_c_247_n 0.0114622f $X=1.205 $Y=0.35 $X2=0 $Y2=0
cc_133 N_A_27_65#_c_211_n N_VGND_c_248_n 0.00977851f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_134 N_A_27_65#_c_214_n N_VGND_c_248_n 0.0371481f $X=1.895 $Y=0.35 $X2=0 $Y2=0
cc_135 N_A_27_65#_c_215_n N_VGND_c_248_n 0.00657784f $X=1.205 $Y=0.35 $X2=0
+ $Y2=0
