* File: sky130_fd_sc_lp__sdlclkp_lp.pex.spice
* Created: Fri Aug 28 11:31:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%GATE 1 3 6 8 10 11 15 17
c34 17 0 8.43713e-20 $X=0.875 $Y=1.37
c35 15 0 7.30689e-20 $X=0.39 $Y=1.2
r36 17 18 0.728097 $w=6.62e-07 $l=1e-08 $layer=POLY_cond $X=0.875 $Y=1.37
+ $X2=0.885 $Y2=1.37
r37 16 17 27.6677 $w=6.62e-07 $l=3.8e-07 $layer=POLY_cond $X=0.495 $Y=1.37
+ $X2=0.875 $Y2=1.37
r38 14 16 7.64502 $w=6.62e-07 $l=1.05e-07 $layer=POLY_cond $X=0.39 $Y=1.37
+ $X2=0.495 $Y2=1.37
r39 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.39 $Y=1.2
+ $X2=0.39 $Y2=1.2
r40 11 15 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=1.37
+ $X2=0.39 $Y2=1.37
r41 8 18 38.6408 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.885 $Y=1.035
+ $X2=0.885 $Y2=1.37
r42 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.885 $Y=1.035
+ $X2=0.885 $Y2=0.715
r43 4 17 25.6903 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.875 $Y=1.705
+ $X2=0.875 $Y2=1.37
r44 4 6 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.875 $Y=1.705
+ $X2=0.875 $Y2=2.38
r45 1 16 38.6408 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.495 $Y=1.035
+ $X2=0.495 $Y2=1.37
r46 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.495 $Y=1.035
+ $X2=0.495 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%SCE 1 3 8 10 12 14 15 16 17 21 22 23
c56 15 0 7.30689e-20 $X=1.315 $Y=1.075
c57 10 0 1.92286e-19 $X=1.6 $Y=1.075
r58 21 24 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.555
+ $X2=1.405 $Y2=1.72
r59 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.555
+ $X2=1.405 $Y2=1.39
r60 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.405
+ $Y=1.555 $X2=1.405 $Y2=1.555
r61 16 17 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.327 $Y=1.665
+ $X2=1.327 $Y2=2.035
r62 16 22 2.71276 $w=4.83e-07 $l=1.1e-07 $layer=LI1_cond $X=1.327 $Y=1.665
+ $X2=1.327 $Y2=1.555
r63 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.675 $Y=1 $X2=1.675
+ $Y2=0.715
r64 11 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.39 $Y=1.075
+ $X2=1.315 $Y2=1.075
r65 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.6 $Y=1.075
+ $X2=1.675 $Y2=1
r66 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.6 $Y=1.075
+ $X2=1.39 $Y2=1.075
r67 8 24 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.365 $Y=2.38
+ $X2=1.365 $Y2=1.72
r68 4 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.315 $Y=1.15
+ $X2=1.315 $Y2=1.075
r69 4 23 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.315 $Y=1.15
+ $X2=1.315 $Y2=1.39
r70 1 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.315 $Y=1 $X2=1.315
+ $Y2=1.075
r71 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.315 $Y=1 $X2=1.315
+ $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_356_278# 1 2 9 11 13 15 16 18 20 21 23
+ 25 27 30 32 33 34 40 43 44 45 47 48 53 60 63 64 67 68 73
c180 68 0 4.27658e-20 $X=6 $Y=2.06
c181 60 0 1.14082e-19 $X=3.895 $Y=1.66
c182 34 0 6.80345e-20 $X=3.055 $Y=0.82
c183 30 0 1.70279e-19 $X=3.895 $Y=2.525
c184 25 0 3.33038e-20 $X=3.555 $Y=0.745
c185 23 0 1.58242e-19 $X=3.48 $Y=0.82
r186 72 73 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=2.105 $Y=1.555
+ $X2=2.11 $Y2=1.555
r187 67 68 7.28026 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=2.225 $X2=6
+ $Y2=2.06
r188 62 64 1.5601 $w=4.58e-07 $l=6e-08 $layer=LI1_cond $X=5.88 $Y=1.17 $X2=5.94
+ $Y2=1.17
r189 62 63 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.88 $Y=1.17
+ $X2=5.715 $Y2=1.17
r190 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.895
+ $Y=1.66 $X2=3.895 $Y2=1.66
r191 53 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.49 $Y=2.35
+ $X2=2.49 $Y2=2.52
r192 51 64 5.34566 $w=2.1e-07 $l=2.3e-07 $layer=LI1_cond $X=5.94 $Y=1.4 $X2=5.94
+ $Y2=1.17
r193 51 68 34.8571 $w=2.08e-07 $l=6.6e-07 $layer=LI1_cond $X=5.94 $Y=1.4
+ $X2=5.94 $Y2=2.06
r194 50 59 13.8 $w=3.05e-07 $l=4.36789e-07 $layer=LI1_cond $X=4.145 $Y=1.315
+ $X2=3.937 $Y2=1.66
r195 50 63 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=4.145 $Y=1.315
+ $X2=5.715 $Y2=1.315
r196 47 59 8.97136 $w=3.05e-07 $l=2.17991e-07 $layer=LI1_cond $X=4.06 $Y=1.825
+ $X2=3.937 $Y2=1.66
r197 47 48 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.06 $Y=1.825
+ $X2=4.06 $Y2=2.435
r198 46 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=2.52
+ $X2=2.49 $Y2=2.52
r199 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.975 $Y=2.52
+ $X2=4.06 $Y2=2.435
r200 45 46 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.975 $Y=2.52
+ $X2=2.575 $Y2=2.52
r201 43 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=2.35
+ $X2=2.49 $Y2=2.35
r202 43 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.405 $Y=2.35
+ $X2=2.11 $Y2=2.35
r203 41 72 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.945 $Y=1.555
+ $X2=2.105 $Y2=1.555
r204 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.945
+ $Y=1.555 $X2=1.945 $Y2=1.555
r205 38 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=2.265
+ $X2=2.11 $Y2=2.35
r206 38 40 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.945 $Y=2.265
+ $X2=1.945 $Y2=1.555
r207 34 36 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=3.055 $Y=0.82
+ $X2=3.055 $Y2=1.075
r208 28 60 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.895 $Y=1.825
+ $X2=3.895 $Y2=1.66
r209 28 30 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.895 $Y=1.825
+ $X2=3.895 $Y2=2.525
r210 25 27 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.555 $Y=0.745 $X2=3.555
+ $Y2=0.445
r211 24 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=0.82
+ $X2=3.055 $Y2=0.82
r212 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.48 $Y=0.82
+ $X2=3.555 $Y2=0.745
r213 23 24 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.48 $Y=0.82
+ $X2=3.13 $Y2=0.82
r214 22 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.54 $Y=1.075
+ $X2=2.465 $Y2=1.075
r215 21 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.075
+ $X2=3.055 $Y2=1.075
r216 21 22 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.98 $Y=1.075
+ $X2=2.54 $Y2=1.075
r217 18 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.465 $Y=1
+ $X2=2.465 $Y2=1.075
r218 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.465 $Y=1 $X2=2.465
+ $Y2=0.715
r219 17 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.18 $Y=1.075
+ $X2=2.105 $Y2=1.075
r220 16 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.39 $Y=1.075
+ $X2=2.465 $Y2=1.075
r221 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.39 $Y=1.075
+ $X2=2.18 $Y2=1.075
r222 15 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.105 $Y=1.39
+ $X2=2.105 $Y2=1.555
r223 14 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.105 $Y=1.15
+ $X2=2.105 $Y2=1.075
r224 14 15 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.105 $Y=1.15
+ $X2=2.105 $Y2=1.39
r225 11 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.105 $Y=1
+ $X2=2.105 $Y2=1.075
r226 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.105 $Y=1 $X2=2.105
+ $Y2=0.715
r227 7 73 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.72
+ $X2=2.11 $Y2=1.555
r228 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.11 $Y=1.72 $X2=2.11
+ $Y2=2.38
r229 2 67 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.855
+ $Y=2.08 $X2=6 $Y2=2.225
r230 1 62 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.735
+ $Y=0.96 $X2=5.88 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_447_376# 1 2 7 9 11 15 19 22 25 30 36
c76 15 0 1.35974e-19 $X=3.985 $Y=0.445
r77 34 36 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.76 $Y=0.78
+ $X2=2.885 $Y2=0.78
r78 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.035
+ $Y=1.555 $X2=3.035 $Y2=1.555
r79 28 30 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.885 $Y=1.555
+ $X2=3.035 $Y2=1.555
r80 26 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.455 $Y=1.555
+ $X2=2.885 $Y2=1.555
r81 25 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=1.39
+ $X2=2.885 $Y2=1.555
r82 24 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=0.945
+ $X2=2.885 $Y2=0.78
r83 24 25 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.885 $Y=0.945
+ $X2=2.885 $Y2=1.39
r84 20 26 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=1.72
+ $X2=2.455 $Y2=1.555
r85 20 22 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.455 $Y=1.72 $X2=2.455
+ $Y2=1.92
r86 19 31 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.24 $Y=1.555
+ $X2=3.035 $Y2=1.555
r87 17 19 89.0394 $w=2.03e-07 $l=3.75e-07 $layer=POLY_cond $X=3.365 $Y=1.18
+ $X2=3.365 $Y2=1.555
r88 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.985 $Y=1.105
+ $X2=3.985 $Y2=0.445
r89 12 17 9.92004 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=3.49 $Y=1.18
+ $X2=3.365 $Y2=1.18
r90 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.91 $Y=1.18
+ $X2=3.985 $Y2=1.105
r91 11 12 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.91 $Y=1.18
+ $X2=3.49 $Y2=1.18
r92 7 19 33.6572 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.72
+ $X2=3.365 $Y2=1.555
r93 7 9 200.005 $w=2.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.365 $Y=1.72
+ $X2=3.365 $Y2=2.525
r94 2 22 600 $w=1.7e-07 $l=2.39165e-07 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.88 $X2=2.455 $Y2=1.92
r95 1 34 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=2.54
+ $Y=0.505 $X2=2.76 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_860_21# 1 2 9 13 15 17 20 24 27 28 30
+ 31 34 36 39 41 42 45 46 50 52 58 60 62 63 70
c167 63 0 6.92102e-20 $X=7.92 $Y=1.48
c168 41 0 1.79113e-19 $X=6.43 $Y=2.49
c169 36 0 6.75081e-20 $X=6.225 $Y=0.59
c170 31 0 1.70279e-19 $X=4.655 $Y=2.415
c171 20 0 4.59691e-20 $X=7.325 $Y=2.58
r172 63 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.92 $Y=1.48
+ $X2=7.755 $Y2=1.48
r173 62 65 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.92 $Y=1.48
+ $X2=7.92 $Y2=1.645
r174 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.92
+ $Y=1.48 $X2=7.92 $Y2=1.48
r175 56 58 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.31 $Y=1.665
+ $X2=6.43 $Y2=1.665
r176 52 54 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.61 $Y=0.47
+ $X2=5.61 $Y2=0.59
r177 49 50 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.255 $Y=2.495
+ $X2=5.255 $Y2=2.575
r178 46 49 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.255 $Y=2.415
+ $X2=5.255 $Y2=2.495
r179 45 65 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=7.84 $Y=2.49
+ $X2=7.84 $Y2=1.645
r180 43 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.515 $Y=2.575
+ $X2=6.43 $Y2=2.575
r181 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.755 $Y=2.575
+ $X2=7.84 $Y2=2.49
r182 42 43 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.755 $Y=2.575
+ $X2=6.515 $Y2=2.575
r183 41 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=2.49
+ $X2=6.43 $Y2=2.575
r184 40 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=1.75
+ $X2=6.43 $Y2=1.665
r185 40 41 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.43 $Y=1.75
+ $X2=6.43 $Y2=2.49
r186 39 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.31 $Y=1.58
+ $X2=6.31 $Y2=1.665
r187 38 39 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=6.31 $Y=0.675
+ $X2=6.31 $Y2=1.58
r188 37 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=0.59
+ $X2=5.61 $Y2=0.59
r189 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.225 $Y=0.59
+ $X2=6.31 $Y2=0.675
r190 36 37 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.225 $Y=0.59
+ $X2=5.775 $Y2=0.59
r191 35 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.42 $Y=2.575
+ $X2=5.255 $Y2=2.575
r192 34 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.345 $Y=2.575
+ $X2=6.43 $Y2=2.575
r193 34 35 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.345 $Y=2.575
+ $X2=5.42 $Y2=2.575
r194 30 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.09 $Y=2.415
+ $X2=5.255 $Y2=2.415
r195 30 31 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.09 $Y=2.415
+ $X2=4.655 $Y2=2.415
r196 28 68 31.9397 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=4.477 $Y=1.7
+ $X2=4.477 $Y2=1.865
r197 28 67 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=4.477 $Y=1.7
+ $X2=4.477 $Y2=1.535
r198 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.49
+ $Y=1.7 $X2=4.49 $Y2=1.7
r199 25 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.49 $Y=2.33
+ $X2=4.655 $Y2=2.415
r200 25 27 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=4.49 $Y=2.33
+ $X2=4.49 $Y2=1.7
r201 23 24 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=7.45 $Y=1.53
+ $X2=7.325 $Y2=1.53
r202 23 70 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=7.45 $Y=1.53
+ $X2=7.755 $Y2=1.53
r203 18 24 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=7.325 $Y=1.605
+ $X2=7.325 $Y2=1.53
r204 18 20 242.242 $w=2.5e-07 $l=9.75e-07 $layer=POLY_cond $X=7.325 $Y=1.605
+ $X2=7.325 $Y2=2.58
r205 15 24 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=7.275 $Y=1.455
+ $X2=7.325 $Y2=1.53
r206 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.275 $Y=1.455
+ $X2=7.275 $Y2=1.17
r207 13 68 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.425 $Y=2.525
+ $X2=4.425 $Y2=1.865
r208 9 67 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=4.375 $Y=0.445
+ $X2=4.375 $Y2=1.535
r209 2 49 300 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_PDIFF $count=2 $X=5.115
+ $Y=2.025 $X2=5.255 $Y2=2.495
r210 1 52 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=5.47
+ $Y=0.235 $X2=5.61 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_698_405# 1 2 9 11 13 14 16 18 21 24 31
+ 34 35 36
c82 36 0 5.23495e-20 $X=4.935 $Y=0.907
c83 24 0 6.17323e-20 $X=3.935 $Y=0.965
c84 18 0 1.36704e-19 $X=3.465 $Y=2.005
c85 14 0 6.75081e-20 $X=5.395 $Y=0.735
r86 38 39 2.40199 $w=3.01e-07 $l=1.5e-08 $layer=POLY_cond $X=4.99 $Y=0.977
+ $X2=5.005 $Y2=0.977
r87 35 39 15.2126 $w=3.01e-07 $l=9.5e-08 $layer=POLY_cond $X=5.1 $Y=0.977
+ $X2=5.005 $Y2=0.977
r88 34 36 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=5.1 $Y=0.907
+ $X2=4.935 $Y2=0.907
r89 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.1
+ $Y=0.93 $X2=5.1 $Y2=0.93
r90 28 31 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=2.13
+ $X2=3.63 $Y2=2.13
r91 24 36 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.935 $Y=0.965
+ $X2=4.935 $Y2=0.965
r92 19 24 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.81 $Y=0.965
+ $X2=3.935 $Y2=0.965
r93 19 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.81 $Y=0.965
+ $X2=3.465 $Y2=0.965
r94 19 21 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.81 $Y=0.88
+ $X2=3.81 $Y2=0.47
r95 18 28 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.465 $Y=2.005
+ $X2=3.465 $Y2=2.13
r96 17 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=1.05
+ $X2=3.465 $Y2=0.965
r97 17 18 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.465 $Y=1.05
+ $X2=3.465 $Y2=2.005
r98 14 35 47.2392 $w=3.01e-07 $l=3.98014e-07 $layer=POLY_cond $X=5.395 $Y=0.735
+ $X2=5.1 $Y2=0.977
r99 14 16 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.395 $Y=0.735
+ $X2=5.395 $Y2=0.445
r100 11 39 19.0468 $w=1.5e-07 $l=2.42e-07 $layer=POLY_cond $X=5.005 $Y=0.735
+ $X2=5.005 $Y2=0.977
r101 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.005 $Y=0.735
+ $X2=5.005 $Y2=0.445
r102 7 38 7.2153 $w=2.5e-07 $l=2.43e-07 $layer=POLY_cond $X=4.99 $Y=1.22
+ $X2=4.99 $Y2=0.977
r103 7 9 324.232 $w=2.5e-07 $l=1.305e-06 $layer=POLY_cond $X=4.99 $Y=1.22
+ $X2=4.99 $Y2=2.525
r104 2 31 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=2.025 $X2=3.63 $Y2=2.17
r105 1 21 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.235 $X2=3.77 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%CLK 1 3 5 8 10 12 13 15 17 19 25 26 29
c72 13 0 1.79113e-19 $X=6.795 $Y=1.605
c73 10 0 4.27658e-20 $X=6.455 $Y=1.455
r74 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.49
+ $Y=1.7 $X2=5.49 $Y2=1.7
r75 29 32 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.49 $Y=1.61 $X2=5.49
+ $Y2=1.7
r76 26 33 0.629515 $w=5.68e-07 $l=3e-08 $layer=LI1_cond $X=5.52 $Y=1.865
+ $X2=5.49 $Y2=1.865
r77 25 33 9.44272 $w=5.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.04 $Y=1.865
+ $X2=5.49 $Y2=1.865
r78 17 24 7.26674 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=6.885 $Y=1.455
+ $X2=6.885 $Y2=1.57
r79 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.885 $Y=1.455
+ $X2=6.885 $Y2=1.17
r80 13 24 23.9669 $w=1.81e-07 $l=9e-08 $layer=POLY_cond $X=6.795 $Y=1.57
+ $X2=6.885 $Y2=1.57
r81 13 22 90.5414 $w=1.81e-07 $l=3.4e-07 $layer=POLY_cond $X=6.795 $Y=1.57
+ $X2=6.455 $Y2=1.57
r82 13 15 242.242 $w=2.5e-07 $l=9.75e-07 $layer=POLY_cond $X=6.795 $Y=1.605
+ $X2=6.795 $Y2=2.58
r83 10 22 7.26674 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=6.455 $Y=1.455
+ $X2=6.455 $Y2=1.57
r84 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.455 $Y=1.455
+ $X2=6.455 $Y2=1.17
r85 6 22 50.5967 $w=1.81e-07 $l=1.9e-07 $layer=POLY_cond $X=6.265 $Y=1.57
+ $X2=6.455 $Y2=1.57
r86 6 20 45.2707 $w=1.81e-07 $l=1.7e-07 $layer=POLY_cond $X=6.265 $Y=1.57
+ $X2=6.095 $Y2=1.57
r87 6 8 222.366 $w=2.5e-07 $l=8.95e-07 $layer=POLY_cond $X=6.265 $Y=1.685
+ $X2=6.265 $Y2=2.58
r88 3 20 7.26674 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=6.095 $Y=1.455
+ $X2=6.095 $Y2=1.57
r89 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.095 $Y=1.455
+ $X2=6.095 $Y2=1.17
r90 2 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.655 $Y=1.61
+ $X2=5.49 $Y2=1.61
r91 1 20 21.5288 $w=1.81e-07 $l=9.28709e-08 $layer=POLY_cond $X=6.02 $Y=1.61
+ $X2=6.095 $Y2=1.57
r92 1 2 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=6.02 $Y=1.61 $X2=5.655
+ $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_1384_416# 1 2 7 9 10 12 13 15 16 17 19
+ 23 24 25 27 30 37
c77 24 0 6.92102e-20 $X=7.775 $Y=1.02
r78 37 38 55.787 $w=3.24e-07 $l=3.75e-07 $layer=POLY_cond $X=8.025 $Y=0.92
+ $X2=8.4 $Y2=0.92
r79 31 37 12.6451 $w=3.24e-07 $l=8.5e-08 $layer=POLY_cond $X=7.94 $Y=0.92
+ $X2=8.025 $Y2=0.92
r80 30 33 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.94 $Y=0.94 $X2=7.94
+ $Y2=1.02
r81 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.94
+ $Y=0.94 $X2=7.94 $Y2=0.94
r82 24 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.775 $Y=1.02
+ $X2=7.94 $Y2=1.02
r83 24 25 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.775 $Y=1.02
+ $X2=7.575 $Y2=1.02
r84 21 27 22.875 $w=2.08e-07 $l=3.9e-07 $layer=LI1_cond $X=7.45 $Y=2.185
+ $X2=7.06 $Y2=2.185
r85 21 23 41.027 $w=2.48e-07 $l=8.9e-07 $layer=LI1_cond $X=7.45 $Y=2.06 $X2=7.45
+ $Y2=1.17
r86 20 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.45 $Y=1.105
+ $X2=7.575 $Y2=1.02
r87 20 23 2.99635 $w=2.48e-07 $l=6.5e-08 $layer=LI1_cond $X=7.45 $Y=1.105
+ $X2=7.45 $Y2=1.17
r88 18 38 20.7868 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=8.4 $Y=1.105
+ $X2=8.4 $Y2=0.92
r89 18 19 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=8.4 $Y=1.105 $X2=8.4
+ $Y2=1.855
r90 16 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.325 $Y=1.93
+ $X2=8.4 $Y2=1.855
r91 16 17 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=8.325 $Y=1.93
+ $X2=8.14 $Y2=1.93
r92 13 37 20.7868 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=8.025 $Y=0.735
+ $X2=8.025 $Y2=0.92
r93 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.025 $Y=0.735
+ $X2=8.025 $Y2=0.45
r94 10 17 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=8.015 $Y=2.005
+ $X2=8.14 $Y2=1.93
r95 10 12 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.015 $Y=2.005
+ $X2=8.015 $Y2=2.58
r96 7 31 40.9105 $w=3.24e-07 $l=3.55668e-07 $layer=POLY_cond $X=7.665 $Y=0.735
+ $X2=7.94 $Y2=0.92
r97 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.665 $Y=0.735
+ $X2=7.665 $Y2=0.45
r98 2 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.92
+ $Y=2.08 $X2=7.06 $Y2=2.225
r99 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.35
+ $Y=0.96 $X2=7.49 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_93_376# 1 2 3 4 14 17 21 23 27 30 31 32
+ 34 35 38 39 43
c109 43 0 1.35974e-19 $X=3.34 $Y=0.35
c110 31 0 3.33038e-20 $X=3.175 $Y=0.35
c111 30 0 2.6032e-19 $X=2.32 $Y=1.04
c112 17 0 8.43713e-20 $X=1.1 $Y=0.715
r113 43 46 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.34 $Y=0.35
+ $X2=3.34 $Y2=0.47
r114 34 35 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.675 $Y=2.05
+ $X2=0.675 $Y2=1.885
r115 31 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=0.35
+ $X2=3.34 $Y2=0.35
r116 31 32 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.175 $Y=0.35
+ $X2=2.405 $Y2=0.35
r117 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.32 $Y=0.435
+ $X2=2.405 $Y2=0.35
r118 29 30 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.32 $Y=0.435
+ $X2=2.32 $Y2=1.04
r119 25 39 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.14 $Y=2.915
+ $X2=2.14 $Y2=2.7
r120 25 27 38.7841 $w=2.58e-07 $l=8.75e-07 $layer=LI1_cond $X=2.225 $Y=2.915
+ $X2=3.1 $Y2=2.915
r121 24 38 4.03347 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.265 $Y=1.125
+ $X2=1 $Y2=1.125
r122 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.235 $Y=1.125
+ $X2=2.32 $Y2=1.04
r123 23 24 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=2.235 $Y=1.125
+ $X2=1.265 $Y2=1.125
r124 22 37 5.94789 $w=1.7e-07 $l=2.56924e-07 $layer=LI1_cond $X=0.905 $Y=2.7
+ $X2=0.675 $Y2=2.757
r125 21 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.7
+ $X2=2.14 $Y2=2.7
r126 21 22 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=2.055 $Y=2.7
+ $X2=0.905 $Y2=2.7
r127 19 38 2.73602 $w=3.5e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.82 $Y=1.21
+ $X2=1 $Y2=1.125
r128 19 35 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.82 $Y=1.21
+ $X2=0.82 $Y2=1.885
r129 15 38 2.73602 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1 $Y=1.04 $X2=1
+ $Y2=1.125
r130 15 17 7.33444 $w=5.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1 $Y=1.04 $X2=1
+ $Y2=0.715
r131 14 37 2.94286 $w=4.6e-07 $l=1.42e-07 $layer=LI1_cond $X=0.675 $Y=2.615
+ $X2=0.675 $Y2=2.757
r132 13 34 1.69011 $w=4.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.675 $Y=2.115
+ $X2=0.675 $Y2=2.05
r133 13 14 13.0009 $w=4.58e-07 $l=5e-07 $layer=LI1_cond $X=0.675 $Y=2.115
+ $X2=0.675 $Y2=2.615
r134 4 27 600 $w=1.7e-07 $l=9.19647e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=2.025 $X2=3.1 $Y2=2.875
r135 3 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.465
+ $Y=1.88 $X2=0.61 $Y2=2.735
r136 3 34 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=0.465
+ $Y=1.88 $X2=0.61 $Y2=2.05
r137 2 46 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=3.195
+ $Y=0.235 $X2=3.34 $Y2=0.47
r138 1 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.505 $X2=1.1 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%VPWR 1 2 3 4 15 19 23 26 27 28 30 38 43
+ 56 57 60 67 70
r91 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r92 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r94 60 63 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.71 $Y=3.05 $X2=1.71
+ $Y2=3.33
r95 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r96 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r97 54 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r98 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r99 51 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.53 $Y2=3.33
r100 51 53 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=7.44 $Y2=3.33
r101 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r102 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r103 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r104 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r105 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r106 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r107 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.69 $Y2=3.33
r108 44 46 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 43 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.365 $Y=3.33
+ $X2=6.53 $Y2=3.33
r110 43 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.365 $Y=3.33
+ $X2=6 $Y2=3.33
r111 42 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r113 39 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.71 $Y2=3.33
r114 39 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 38 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.69 $Y2=3.33
r116 38 41 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 37 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r118 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 33 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 32 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r121 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r122 30 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.71 $Y2=3.33
r123 30 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 28 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 28 42 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 26 53 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.505 $Y=3.33
+ $X2=7.44 $Y2=3.33
r127 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.505 $Y=3.33
+ $X2=7.67 $Y2=3.33
r128 25 56 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=8.4 $Y2=3.33
r129 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.67 $Y2=3.33
r130 21 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=3.245
+ $X2=7.67 $Y2=3.33
r131 21 23 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=7.67 $Y=3.245
+ $X2=7.67 $Y2=3.005
r132 17 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=3.245
+ $X2=6.53 $Y2=3.33
r133 17 19 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=6.53 $Y=3.245
+ $X2=6.53 $Y2=2.93
r134 13 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=3.245
+ $X2=4.69 $Y2=3.33
r135 13 15 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=4.69 $Y=3.245
+ $X2=4.69 $Y2=2.86
r136 4 23 600 $w=1.7e-07 $l=1.02914e-06 $layer=licon1_PDIFF $count=1 $X=7.45
+ $Y=2.08 $X2=7.67 $Y2=3.005
r137 3 19 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=6.39
+ $Y=2.08 $X2=6.53 $Y2=2.93
r138 2 15 600 $w=1.7e-07 $l=9.02289e-07 $layer=licon1_PDIFF $count=1 $X=4.55
+ $Y=2.025 $X2=4.69 $Y2=2.86
r139 1 60 600 $w=1.7e-07 $l=1.27526e-06 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.88 $X2=1.71 $Y2=3.05
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%GCLK 1 2 7 8 9 10 11 12 32
c26 11 0 4.59691e-20 $X=8.315 $Y=1.95
r27 33 45 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=8.315 $Y=2.26
+ $X2=8.315 $Y2=2.225
r28 32 43 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=8.4 $Y=2.035 $X2=8.4
+ $Y2=2.06
r29 12 33 4.4225 $w=4e-07 $l=1.45e-07 $layer=LI1_cond $X=8.315 $Y=2.405
+ $X2=8.315 $Y2=2.26
r30 11 45 3.8895 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=8.315 $Y=2.09
+ $X2=8.315 $Y2=2.225
r31 11 43 2.92847 $w=3.98e-07 $l=3e-08 $layer=LI1_cond $X=8.315 $Y=2.09
+ $X2=8.315 $Y2=2.06
r32 11 32 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=8.4 $Y=2.005 $X2=8.4
+ $Y2=2.035
r33 10 11 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.4 $Y=1.665 $X2=8.4
+ $Y2=2.005
r34 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.4 $Y=1.295 $X2=8.4
+ $Y2=1.665
r35 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.4 $Y=0.925 $X2=8.4
+ $Y2=1.295
r36 7 21 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.4 $Y=0.43 $X2=8.4
+ $Y2=0.595
r37 7 37 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=8.4 $Y=0.43 $X2=8.24
+ $Y2=0.43
r38 7 8 15.4327 $w=2.28e-07 $l=3.08e-07 $layer=LI1_cond $X=8.4 $Y=0.617 $X2=8.4
+ $Y2=0.925
r39 7 21 1.10234 $w=2.28e-07 $l=2.2e-08 $layer=LI1_cond $X=8.4 $Y=0.617 $X2=8.4
+ $Y2=0.595
r40 2 45 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.14
+ $Y=2.08 $X2=8.28 $Y2=2.225
r41 1 37 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=8.1 $Y=0.24
+ $X2=8.24 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_LP%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40
+ 41 42 51 65 71 72 78 81
c106 72 0 2.15376e-20 $X=8.4 $Y=0
r107 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r108 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r109 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r110 72 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r111 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r112 69 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=0 $X2=7.43
+ $Y2=0
r113 69 71 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=7.595 $Y=0 $X2=8.4
+ $Y2=0
r114 68 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r115 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r116 65 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.265 $Y=0 $X2=7.43
+ $Y2=0
r117 65 67 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.265 $Y=0
+ $X2=6.96 $Y2=0
r118 64 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r119 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r120 61 64 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r121 61 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r122 60 63 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r123 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r124 58 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.59
+ $Y2=0
r125 58 60 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=5.04 $Y2=0
r126 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r127 54 57 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r128 53 56 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r129 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r130 51 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.59
+ $Y2=0
r131 51 56 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.08
+ $Y2=0
r132 50 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r133 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r134 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r135 47 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r136 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r137 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r138 44 75 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r139 44 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r140 42 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r141 42 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r142 40 63 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=6.585 $Y=0
+ $X2=6.48 $Y2=0
r143 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.585 $Y=0 $X2=6.71
+ $Y2=0
r144 39 67 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.835 $Y=0
+ $X2=6.96 $Y2=0
r145 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.835 $Y=0 $X2=6.71
+ $Y2=0
r146 37 49 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.725 $Y=0 $X2=1.68
+ $Y2=0
r147 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=0 $X2=1.89
+ $Y2=0
r148 36 53 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=2.16 $Y2=0
r149 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=1.89
+ $Y2=0
r150 32 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=0.085
+ $X2=7.43 $Y2=0
r151 32 34 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.43 $Y=0.085
+ $X2=7.43 $Y2=0.45
r152 28 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.71 $Y=0.085
+ $X2=6.71 $Y2=0
r153 28 30 50.016 $w=2.48e-07 $l=1.085e-06 $layer=LI1_cond $X=6.71 $Y=0.085
+ $X2=6.71 $Y2=1.17
r154 24 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0
r155 24 26 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.59 $Y=0.085
+ $X2=4.59 $Y2=0.445
r156 20 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.89 $Y=0.085
+ $X2=1.89 $Y2=0
r157 20 22 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=1.89 $Y=0.085
+ $X2=1.89 $Y2=0.67
r158 16 75 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r159 16 18 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.67
r160 5 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.285
+ $Y=0.24 $X2=7.43 $Y2=0.45
r161 4 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.53
+ $Y=0.96 $X2=6.67 $Y2=1.17
r162 3 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.45
+ $Y=0.235 $X2=4.59 $Y2=0.445
r163 2 22 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.505 $X2=1.89 $Y2=0.67
r164 1 18 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.505 $X2=0.28 $Y2=0.67
.ends

