* File: sky130_fd_sc_lp__a211oi_4.pex.spice
* Created: Fri Aug 28 09:48:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211OI_4%A2 3 5 7 10 12 14 17 19 21 24 28 30 32 33
+ 35 36 38 39 40 54
c111 36 0 8.73804e-20 $X=3.595 $Y=1.44
c112 24 0 1.47759e-19 $X=3.505 $Y=0.655
r113 54 55 7.97636 $w=4.23e-07 $l=7e-08 $layer=POLY_cond $X=1.355 $Y=1.51
+ $X2=1.425 $Y2=1.51
r114 52 54 5.6974 $w=4.23e-07 $l=5e-08 $layer=POLY_cond $X=1.305 $Y=1.51
+ $X2=1.355 $Y2=1.51
r115 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.305
+ $Y=1.46 $X2=1.305 $Y2=1.46
r116 50 52 35.3239 $w=4.23e-07 $l=3.1e-07 $layer=POLY_cond $X=0.995 $Y=1.51
+ $X2=1.305 $Y2=1.51
r117 49 50 7.97636 $w=4.23e-07 $l=7e-08 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.995 $Y2=1.51
r118 48 49 41.0213 $w=4.23e-07 $l=3.6e-07 $layer=POLY_cond $X=0.565 $Y=1.51
+ $X2=0.925 $Y2=1.51
r119 47 48 7.97636 $w=4.23e-07 $l=7e-08 $layer=POLY_cond $X=0.495 $Y=1.51
+ $X2=0.565 $Y2=1.51
r120 45 47 23.9291 $w=4.23e-07 $l=2.1e-07 $layer=POLY_cond $X=0.285 $Y=1.51
+ $X2=0.495 $Y2=1.51
r121 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.285
+ $Y=1.46 $X2=0.285 $Y2=1.46
r122 40 53 2.75015 $w=4.38e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.305 $Y2=1.565
r123 39 40 12.5721 $w=4.38e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r124 39 46 11.3935 $w=4.38e-07 $l=4.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.285 $Y2=1.565
r125 38 46 1.17863 $w=4.38e-07 $l=4.5e-08 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.285 $Y2=1.565
r126 36 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.44
+ $X2=3.595 $Y2=1.605
r127 36 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.44
+ $X2=3.595 $Y2=1.275
r128 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.595
+ $Y=1.44 $X2=3.595 $Y2=1.44
r129 32 53 3.14303 $w=4.38e-07 $l=1.2e-07 $layer=LI1_cond $X=1.425 $Y=1.565
+ $X2=1.305 $Y2=1.565
r130 32 33 10.2759 $w=4.38e-07 $l=2.2e-07 $layer=LI1_cond $X=1.425 $Y=1.565
+ $X2=1.645 $Y2=1.565
r131 30 35 11.5345 $w=2.75e-07 $l=3.40911e-07 $layer=LI1_cond $X=3.385 $Y=1.7
+ $X2=3.572 $Y2=1.44
r132 30 33 113.519 $w=1.68e-07 $l=1.74e-06 $layer=LI1_cond $X=3.385 $Y=1.7
+ $X2=1.645 $Y2=1.7
r133 28 58 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.625 $Y=2.465
+ $X2=3.625 $Y2=1.605
r134 24 57 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.505 $Y=0.655
+ $X2=3.505 $Y2=1.275
r135 19 55 27.2344 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.425 $Y=1.725
+ $X2=1.425 $Y2=1.51
r136 19 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.425 $Y=1.725
+ $X2=1.425 $Y2=2.465
r137 15 54 27.2344 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.355 $Y=1.295
+ $X2=1.355 $Y2=1.51
r138 15 17 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.355 $Y=1.295
+ $X2=1.355 $Y2=0.655
r139 12 50 27.2344 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.995 $Y=1.725
+ $X2=0.995 $Y2=1.51
r140 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.995 $Y=1.725
+ $X2=0.995 $Y2=2.465
r141 8 49 27.2344 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.925 $Y=1.295
+ $X2=0.925 $Y2=1.51
r142 8 10 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.925 $Y=1.295
+ $X2=0.925 $Y2=0.655
r143 5 48 27.2344 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.565 $Y=1.725
+ $X2=0.565 $Y2=1.51
r144 5 7 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.565 $Y=1.725
+ $X2=0.565 $Y2=2.465
r145 1 47 27.2344 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.51
r146 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 50
c76 31 0 8.73804e-20 $X=3.12 $Y=1.295
r77 50 51 10.6435 $w=3.17e-07 $l=7e-08 $layer=POLY_cond $X=3.075 $Y=1.35
+ $X2=3.145 $Y2=1.35
r78 48 50 8.36278 $w=3.17e-07 $l=5.5e-08 $layer=POLY_cond $X=3.02 $Y=1.35
+ $X2=3.075 $Y2=1.35
r79 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.02
+ $Y=1.35 $X2=3.02 $Y2=1.35
r80 46 48 46.3754 $w=3.17e-07 $l=3.05e-07 $layer=POLY_cond $X=2.715 $Y=1.35
+ $X2=3.02 $Y2=1.35
r81 45 46 10.6435 $w=3.17e-07 $l=7e-08 $layer=POLY_cond $X=2.645 $Y=1.35
+ $X2=2.715 $Y2=1.35
r82 43 45 46.3754 $w=3.17e-07 $l=3.05e-07 $layer=POLY_cond $X=2.34 $Y=1.35
+ $X2=2.645 $Y2=1.35
r83 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.34
+ $Y=1.35 $X2=2.34 $Y2=1.35
r84 41 43 8.36278 $w=3.17e-07 $l=5.5e-08 $layer=POLY_cond $X=2.285 $Y=1.35
+ $X2=2.34 $Y2=1.35
r85 40 41 10.6435 $w=3.17e-07 $l=7e-08 $layer=POLY_cond $X=2.215 $Y=1.35
+ $X2=2.285 $Y2=1.35
r86 38 40 32.6909 $w=3.17e-07 $l=2.15e-07 $layer=POLY_cond $X=2 $Y=1.35
+ $X2=2.215 $Y2=1.35
r87 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2 $Y=1.35
+ $X2=2 $Y2=1.35
r88 36 38 22.0473 $w=3.17e-07 $l=1.45e-07 $layer=POLY_cond $X=1.855 $Y=1.35
+ $X2=2 $Y2=1.35
r89 35 36 10.6435 $w=3.17e-07 $l=7e-08 $layer=POLY_cond $X=1.785 $Y=1.35
+ $X2=1.855 $Y2=1.35
r90 31 49 4.34884 $w=2.63e-07 $l=1e-07 $layer=LI1_cond $X=3.12 $Y=1.312 $X2=3.02
+ $Y2=1.312
r91 30 49 16.5256 $w=2.63e-07 $l=3.8e-07 $layer=LI1_cond $X=2.64 $Y=1.312
+ $X2=3.02 $Y2=1.312
r92 30 44 13.0465 $w=2.63e-07 $l=3e-07 $layer=LI1_cond $X=2.64 $Y=1.312 $X2=2.34
+ $Y2=1.312
r93 29 44 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=2.16 $Y=1.312
+ $X2=2.34 $Y2=1.312
r94 29 39 6.95815 $w=2.63e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=1.312 $X2=2
+ $Y2=1.312
r95 25 51 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.515
+ $X2=3.145 $Y2=1.35
r96 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.145 $Y=1.515
+ $X2=3.145 $Y2=2.465
r97 22 50 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.185
+ $X2=3.075 $Y2=1.35
r98 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.075 $Y=1.185
+ $X2=3.075 $Y2=0.655
r99 18 46 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.515
+ $X2=2.715 $Y2=1.35
r100 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.715 $Y=1.515
+ $X2=2.715 $Y2=2.465
r101 15 45 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.185
+ $X2=2.645 $Y2=1.35
r102 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.645 $Y=1.185
+ $X2=2.645 $Y2=0.655
r103 11 41 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.515
+ $X2=2.285 $Y2=1.35
r104 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.285 $Y=1.515
+ $X2=2.285 $Y2=2.465
r105 8 40 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.185
+ $X2=2.215 $Y2=1.35
r106 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.215 $Y=1.185
+ $X2=2.215 $Y2=0.655
r107 4 36 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.855 $Y2=1.35
r108 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.855 $Y2=2.465
r109 1 35 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.185
+ $X2=1.785 $Y2=1.35
r110 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.785 $Y=1.185
+ $X2=1.785 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_4%B1 1 3 6 8 10 13 15 17 20 24 27 29 31 35 37
+ 38 39 53 56 66 68
r117 53 54 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=4.905 $Y=1.35
+ $X2=4.915 $Y2=1.35
r118 52 66 2.64495 $w=3.03e-07 $l=7e-08 $layer=LI1_cond $X=4.825 $Y=1.362
+ $X2=4.895 $Y2=1.362
r119 51 53 11.7561 $w=3.28e-07 $l=8e-08 $layer=POLY_cond $X=4.825 $Y=1.35
+ $X2=4.905 $Y2=1.35
r120 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.825
+ $Y=1.35 $X2=4.825 $Y2=1.35
r121 49 51 49.9634 $w=3.28e-07 $l=3.4e-07 $layer=POLY_cond $X=4.485 $Y=1.35
+ $X2=4.825 $Y2=1.35
r122 48 49 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=4.475 $Y=1.35
+ $X2=4.485 $Y2=1.35
r123 46 48 48.4939 $w=3.28e-07 $l=3.3e-07 $layer=POLY_cond $X=4.145 $Y=1.35
+ $X2=4.475 $Y2=1.35
r124 44 46 13.2256 $w=3.28e-07 $l=9e-08 $layer=POLY_cond $X=4.055 $Y=1.35
+ $X2=4.145 $Y2=1.35
r125 43 44 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=4.045 $Y=1.35
+ $X2=4.055 $Y2=1.35
r126 39 68 8.11487 $w=4.28e-07 $l=1.4e-07 $layer=LI1_cond $X=5.04 $Y=1.3
+ $X2=5.18 $Y2=1.3
r127 39 66 4.87572 $w=4.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.04 $Y=1.3
+ $X2=4.895 $Y2=1.3
r128 38 52 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=4.56 $Y=1.362
+ $X2=4.825 $Y2=1.362
r129 37 38 18.1368 $w=3.03e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.362
+ $X2=4.56 $Y2=1.362
r130 37 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.145
+ $Y=1.35 $X2=4.145 $Y2=1.35
r131 35 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.145 $Y=1.35
+ $X2=7.145 $Y2=1.515
r132 35 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.145 $Y=1.35
+ $X2=7.145 $Y2=1.185
r133 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.145
+ $Y=1.35 $X2=7.145 $Y2=1.35
r134 31 34 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=7.11 $Y=1.17
+ $X2=7.11 $Y2=1.35
r135 29 31 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.98 $Y=1.17
+ $X2=7.11 $Y2=1.17
r136 29 68 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=6.98 $Y=1.17
+ $X2=5.18 $Y2=1.17
r137 27 57 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.065 $Y=2.465
+ $X2=7.065 $Y2=1.515
r138 24 56 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.055 $Y=0.655
+ $X2=7.055 $Y2=1.185
r139 18 54 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.915 $Y=1.515
+ $X2=4.915 $Y2=1.35
r140 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.915 $Y=1.515
+ $X2=4.915 $Y2=2.465
r141 15 53 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=1.185
+ $X2=4.905 $Y2=1.35
r142 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.905 $Y=1.185
+ $X2=4.905 $Y2=0.655
r143 11 49 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.485 $Y=1.515
+ $X2=4.485 $Y2=1.35
r144 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.485 $Y=1.515
+ $X2=4.485 $Y2=2.465
r145 8 48 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.475 $Y=1.185
+ $X2=4.475 $Y2=1.35
r146 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.475 $Y=1.185
+ $X2=4.475 $Y2=0.655
r147 4 44 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.055 $Y=1.515
+ $X2=4.055 $Y2=1.35
r148 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.055 $Y=1.515
+ $X2=4.055 $Y2=2.465
r149 1 43 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.045 $Y=1.185
+ $X2=4.045 $Y2=1.35
r150 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.045 $Y=1.185
+ $X2=4.045 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_4%C1 3 7 11 15 19 23 27 31 38 41 42 58 60 67
+ 69
c94 11 0 5.86634e-20 $X=5.765 $Y=0.655
r95 60 67 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=5.975 $Y=1.595
+ $X2=6 $Y2=1.595
r96 57 58 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.625 $Y=1.51
+ $X2=6.635 $Y2=1.51
r97 52 53 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.765 $Y=1.51
+ $X2=5.775 $Y2=1.51
r98 50 52 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.515 $Y=1.51
+ $X2=5.765 $Y2=1.51
r99 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.515
+ $Y=1.51 $X2=5.515 $Y2=1.51
r100 48 50 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=5.345 $Y=1.51
+ $X2=5.515 $Y2=1.51
r101 46 48 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.335 $Y=1.51
+ $X2=5.345 $Y2=1.51
r102 42 69 5.33071 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=6.03 $Y=1.595
+ $X2=6.145 $Y2=1.595
r103 42 67 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=6.03 $Y=1.595 $X2=6
+ $Y2=1.595
r104 42 60 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=5.945 $Y=1.595
+ $X2=5.975 $Y2=1.595
r105 41 42 14.4055 $w=3.38e-07 $l=4.25e-07 $layer=LI1_cond $X=5.52 $Y=1.595
+ $X2=5.945 $Y2=1.595
r106 41 51 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=5.52 $Y=1.595
+ $X2=5.515 $Y2=1.595
r107 39 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.535 $Y=1.51
+ $X2=6.625 $Y2=1.51
r108 39 55 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=6.535 $Y=1.51
+ $X2=6.205 $Y2=1.51
r109 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.535
+ $Y=1.51 $X2=6.535 $Y2=1.51
r110 36 55 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.195 $Y=1.51
+ $X2=6.205 $Y2=1.51
r111 36 53 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=6.195 $Y=1.51
+ $X2=5.775 $Y2=1.51
r112 35 38 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=6.195 $Y=1.535
+ $X2=6.535 $Y2=1.535
r113 35 69 2.61919 $w=2.18e-07 $l=5e-08 $layer=LI1_cond $X=6.195 $Y=1.535
+ $X2=6.145 $Y2=1.535
r114 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.195
+ $Y=1.51 $X2=6.195 $Y2=1.51
r115 29 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.635 $Y=1.675
+ $X2=6.635 $Y2=1.51
r116 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.635 $Y=1.675
+ $X2=6.635 $Y2=2.465
r117 25 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.625 $Y=1.345
+ $X2=6.625 $Y2=1.51
r118 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.625 $Y=1.345
+ $X2=6.625 $Y2=0.655
r119 21 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.675
+ $X2=6.205 $Y2=1.51
r120 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.205 $Y=1.675
+ $X2=6.205 $Y2=2.465
r121 17 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.345
+ $X2=6.195 $Y2=1.51
r122 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.195 $Y=1.345
+ $X2=6.195 $Y2=0.655
r123 13 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.775 $Y=1.675
+ $X2=5.775 $Y2=1.51
r124 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.775 $Y=1.675
+ $X2=5.775 $Y2=2.465
r125 9 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.765 $Y=1.345
+ $X2=5.765 $Y2=1.51
r126 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.765 $Y=1.345
+ $X2=5.765 $Y2=0.655
r127 5 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.345 $Y=1.675
+ $X2=5.345 $Y2=1.51
r128 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.345 $Y=1.675
+ $X2=5.345 $Y2=2.465
r129 1 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.335 $Y=1.345
+ $X2=5.335 $Y2=1.51
r130 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.335 $Y=1.345
+ $X2=5.335 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_4%A_45_367# 1 2 3 4 5 6 7 22 24 26 30 32 36
+ 38 42 44 46 48 50 56 57 58 60 65 67 69
r93 72 73 3.23894 $w=2.26e-07 $l=6e-08 $layer=LI1_cond $X=3.82 $Y=1.98 $X2=3.82
+ $Y2=2.04
r94 70 72 10.2566 $w=2.26e-07 $l=1.9e-07 $layer=LI1_cond $X=3.82 $Y=1.79
+ $X2=3.82 $Y2=1.98
r95 58 75 3.18275 $w=3.3e-07 $l=2.05e-07 $layer=LI1_cond $X=7.3 $Y=2.575 $X2=7.3
+ $Y2=2.37
r96 58 60 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=7.3 $Y=2.575
+ $X2=7.3 $Y2=2.95
r97 56 75 3.80378 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=7.135 $Y=2.45
+ $X2=7.3 $Y2=2.37
r98 56 57 107.408 $w=2.48e-07 $l=2.33e-06 $layer=LI1_cond $X=7.135 $Y=2.45
+ $X2=4.805 $Y2=2.45
r99 53 57 6.88375 $w=2.5e-07 $l=1.69558e-07 $layer=LI1_cond $X=4.7 $Y=2.325
+ $X2=4.805 $Y2=2.45
r100 53 55 18.2208 $w=2.08e-07 $l=3.45e-07 $layer=LI1_cond $X=4.7 $Y=2.325
+ $X2=4.7 $Y2=1.98
r101 52 55 5.54545 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=4.7 $Y=1.875
+ $X2=4.7 $Y2=1.98
r102 51 70 2.4068 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.945 $Y=1.79
+ $X2=3.82 $Y2=1.79
r103 50 52 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.595 $Y=1.79
+ $X2=4.7 $Y2=1.875
r104 50 51 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.595 $Y=1.79
+ $X2=3.945 $Y2=1.79
r105 46 73 4.28604 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=2.125
+ $X2=3.82 $Y2=2.04
r106 46 48 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=3.82 $Y=2.125
+ $X2=3.82 $Y2=2.45
r107 45 69 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.025 $Y=2.04
+ $X2=2.93 $Y2=2.04
r108 44 73 2.4068 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.695 $Y=2.04
+ $X2=3.82 $Y2=2.04
r109 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.695 $Y=2.04
+ $X2=3.025 $Y2=2.04
r110 40 69 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=2.125
+ $X2=2.93 $Y2=2.04
r111 40 42 45.2392 $w=1.88e-07 $l=7.75e-07 $layer=LI1_cond $X=2.93 $Y=2.125
+ $X2=2.93 $Y2=2.9
r112 39 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.165 $Y=2.04
+ $X2=2.07 $Y2=2.04
r113 38 69 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.835 $Y=2.04
+ $X2=2.93 $Y2=2.04
r114 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.835 $Y=2.04
+ $X2=2.165 $Y2=2.04
r115 34 67 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.125
+ $X2=2.07 $Y2=2.04
r116 34 36 45.823 $w=1.88e-07 $l=7.85e-07 $layer=LI1_cond $X=2.07 $Y=2.125
+ $X2=2.07 $Y2=2.91
r117 33 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.305 $Y=2.04
+ $X2=1.21 $Y2=2.04
r118 32 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.975 $Y=2.04
+ $X2=2.07 $Y2=2.04
r119 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=2.04
+ $X2=1.305 $Y2=2.04
r120 28 65 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=2.125
+ $X2=1.21 $Y2=2.04
r121 28 30 45.823 $w=1.88e-07 $l=7.85e-07 $layer=LI1_cond $X=1.21 $Y=2.125
+ $X2=1.21 $Y2=2.91
r122 27 63 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.445 $Y=2.04
+ $X2=0.315 $Y2=2.04
r123 26 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.115 $Y=2.04
+ $X2=1.21 $Y2=2.04
r124 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.04
+ $X2=0.445 $Y2=2.04
r125 22 63 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.315 $Y=2.125
+ $X2=0.315 $Y2=2.04
r126 22 24 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=0.315 $Y=2.125
+ $X2=0.315 $Y2=2.91
r127 7 75 400 $w=1.7e-07 $l=4.88493e-07 $layer=licon1_PDIFF $count=1 $X=7.14
+ $Y=1.835 $X2=7.3 $Y2=2.25
r128 7 60 400 $w=1.7e-07 $l=1.19232e-06 $layer=licon1_PDIFF $count=1 $X=7.14
+ $Y=1.835 $X2=7.3 $Y2=2.95
r129 6 55 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.56
+ $Y=1.835 $X2=4.7 $Y2=1.98
r130 5 72 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=1.835 $X2=3.84 $Y2=1.98
r131 5 48 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=3.7
+ $Y=1.835 $X2=3.84 $Y2=2.45
r132 4 69 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.835 $X2=2.93 $Y2=2.12
r133 4 42 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.835 $X2=2.93 $Y2=2.9
r134 3 67 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.835 $X2=2.07 $Y2=2.12
r135 3 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.835 $X2=2.07 $Y2=2.91
r136 2 65 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.835 $X2=1.21 $Y2=2.12
r137 2 30 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.835 $X2=1.21 $Y2=2.91
r138 1 63 400 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.835 $X2=0.35 $Y2=2.12
r139 1 24 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.835 $X2=0.35 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_4%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 35 37
+ 42 58 59 62 65
r100 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r103 55 58 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r104 55 56 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 53 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r106 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r107 50 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r108 50 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 47 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.64 $Y2=3.33
r111 47 49 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=2.16 $Y2=3.33
r112 46 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r113 46 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r114 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r115 43 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r116 43 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r117 42 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=3.33
+ $X2=1.64 $Y2=3.33
r118 42 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 40 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r121 37 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r122 37 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r123 35 59 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=7.44 $Y2=3.33
r124 35 56 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r125 33 52 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.12 $Y2=3.33
r126 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.36 $Y2=3.33
r127 32 55 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=3.6 $Y2=3.33
r128 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=3.36 $Y2=3.33
r129 30 49 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.5 $Y2=3.33
r131 29 52 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=3.12 $Y2=3.33
r132 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=2.5 $Y2=3.33
r133 25 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=3.245
+ $X2=3.36 $Y2=3.33
r134 25 27 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=3.36 $Y=3.245
+ $X2=3.36 $Y2=2.41
r135 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=3.245 $X2=2.5
+ $Y2=3.33
r136 21 23 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=2.5 $Y=3.245
+ $X2=2.5 $Y2=2.41
r137 17 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=3.245
+ $X2=1.64 $Y2=3.33
r138 17 19 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=1.64 $Y=3.245
+ $X2=1.64 $Y2=2.4
r139 13 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r140 13 15 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.4
r141 4 27 300 $w=1.7e-07 $l=6.4119e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=1.835 $X2=3.36 $Y2=2.41
r142 3 23 300 $w=1.7e-07 $l=6.4119e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=1.835 $X2=2.5 $Y2=2.41
r143 2 19 300 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=2.4
r144 1 15 300 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=2 $X=0.64
+ $Y=1.835 $X2=0.78 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_4%A_826_367# 1 2 3 4 13 15 23
r26 21 23 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.99 $Y=2.91
+ $X2=6.85 $Y2=2.91
r27 19 21 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.13 $Y=2.91
+ $X2=5.99 $Y2=2.91
r28 17 26 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=4.375 $Y=2.91
+ $X2=4.27 $Y2=2.91
r29 17 19 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=4.375 $Y=2.91
+ $X2=5.13 $Y2=2.91
r30 13 26 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=2.745
+ $X2=4.27 $Y2=2.91
r31 13 15 28.2554 $w=2.08e-07 $l=5.35e-07 $layer=LI1_cond $X=4.27 $Y=2.745
+ $X2=4.27 $Y2=2.21
r32 4 23 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.71
+ $Y=1.835 $X2=6.85 $Y2=2.91
r33 3 21 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.85
+ $Y=1.835 $X2=5.99 $Y2=2.91
r34 2 19 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.99
+ $Y=1.835 $X2=5.13 $Y2=2.91
r35 1 26 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.13
+ $Y=1.835 $X2=4.27 $Y2=2.91
r36 1 15 300 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=2 $X=4.13
+ $Y=1.835 $X2=4.27 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_4%Y 1 2 3 4 5 6 7 8 27 29 33 35 37 43 45 47
+ 51 53 56 57 58 59 65 66 67 72 79 83 88
c142 66 0 1.47759e-19 $X=4.08 $Y=0.925
c143 57 0 5.86634e-20 $X=5.12 $Y=0.82
r144 79 83 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=4.583 $Y=0.867
+ $X2=4.56 $Y2=0.867
r145 74 77 38.8667 $w=2.53e-07 $l=8.6e-07 $layer=LI1_cond $X=2 $Y=0.882 $X2=2.86
+ $Y2=0.882
r146 67 88 5.77195 $w=2.83e-07 $l=1.11e-07 $layer=LI1_cond $X=4.614 $Y=0.867
+ $X2=4.725 $Y2=0.867
r147 67 79 1.25353 $w=2.83e-07 $l=3.1e-08 $layer=LI1_cond $X=4.614 $Y=0.867
+ $X2=4.583 $Y2=0.867
r148 67 83 1.25353 $w=2.83e-07 $l=3.1e-08 $layer=LI1_cond $X=4.529 $Y=0.867
+ $X2=4.56 $Y2=0.867
r149 67 80 7.03597 $w=2.83e-07 $l=1.74e-07 $layer=LI1_cond $X=4.529 $Y=0.867
+ $X2=4.355 $Y2=0.867
r150 66 72 5.63431 $w=2.7e-07 $l=1.57321e-07 $layer=LI1_cond $X=4.205 $Y=0.867
+ $X2=4.055 $Y2=0.882
r151 66 80 5.63431 $w=2.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.205 $Y=0.867
+ $X2=4.355 $Y2=0.867
r152 66 72 1.35582 $w=2.53e-07 $l=3e-08 $layer=LI1_cond $X=4.025 $Y=0.882
+ $X2=4.055 $Y2=0.882
r153 66 77 52.6508 $w=2.53e-07 $l=1.165e-06 $layer=LI1_cond $X=4.025 $Y=0.882
+ $X2=2.86 $Y2=0.882
r154 62 63 2.30489 $w=2.98e-07 $l=6e-08 $layer=LI1_cond $X=6.465 $Y=1.98
+ $X2=6.465 $Y2=2.04
r155 59 62 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=6.465 $Y=1.9
+ $X2=6.465 $Y2=1.98
r156 55 56 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=7.495 $Y=0.915
+ $X2=7.495 $Y2=1.815
r157 54 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=0.83
+ $X2=6.84 $Y2=0.83
r158 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.41 $Y=0.83
+ $X2=7.495 $Y2=0.915
r159 53 54 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.41 $Y=0.83
+ $X2=7.005 $Y2=0.83
r160 49 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.745
+ $X2=6.84 $Y2=0.83
r161 49 51 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=6.84 $Y=0.745
+ $X2=6.84 $Y2=0.37
r162 48 59 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.615 $Y=1.9 $X2=6.465
+ $Y2=1.9
r163 47 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.41 $Y=1.9
+ $X2=7.495 $Y2=1.815
r164 47 48 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=7.41 $Y=1.9
+ $X2=6.615 $Y2=1.9
r165 46 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=0.83
+ $X2=5.98 $Y2=0.83
r166 45 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=0.83
+ $X2=6.84 $Y2=0.83
r167 45 46 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.675 $Y=0.83
+ $X2=6.145 $Y2=0.83
r168 41 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=0.745
+ $X2=5.98 $Y2=0.83
r169 41 43 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.98 $Y=0.745
+ $X2=5.98 $Y2=0.37
r170 37 63 2.82627 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=6.315 $Y=2.04
+ $X2=6.465 $Y2=2.04
r171 37 39 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=6.315 $Y=2.04
+ $X2=5.56 $Y2=2.04
r172 36 57 8.26956 $w=1.8e-07 $l=1.69926e-07 $layer=LI1_cond $X=5.285 $Y=0.83
+ $X2=5.12 $Y2=0.82
r173 35 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=0.83
+ $X2=5.98 $Y2=0.83
r174 35 36 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.815 $Y=0.83
+ $X2=5.285 $Y2=0.83
r175 31 57 0.718145 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=5.12 $Y=0.725
+ $X2=5.12 $Y2=0.82
r176 31 33 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.12 $Y=0.725
+ $X2=5.12 $Y2=0.37
r177 29 57 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.955 $Y=0.82
+ $X2=5.12 $Y2=0.82
r178 29 88 13.4258 $w=1.88e-07 $l=2.3e-07 $layer=LI1_cond $X=4.955 $Y=0.82
+ $X2=4.725 $Y2=0.82
r179 25 66 0.966048 $w=3e-07 $l=1.42e-07 $layer=LI1_cond $X=4.205 $Y=0.725
+ $X2=4.205 $Y2=0.867
r180 25 27 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=4.205 $Y=0.725
+ $X2=4.205 $Y2=0.42
r181 8 62 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.28
+ $Y=1.835 $X2=6.42 $Y2=1.98
r182 7 39 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=1.835 $X2=5.56 $Y2=2.04
r183 6 51 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=6.7
+ $Y=0.235 $X2=6.84 $Y2=0.37
r184 5 43 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=5.84
+ $Y=0.235 $X2=5.98 $Y2=0.37
r185 4 33 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=4.98
+ $Y=0.235 $X2=5.12 $Y2=0.37
r186 3 66 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=4.12
+ $Y=0.235 $X2=4.26 $Y2=0.845
r187 3 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.12
+ $Y=0.235 $X2=4.26 $Y2=0.42
r188 2 77 182 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_NDIFF $count=1 $X=2.72
+ $Y=0.235 $X2=2.86 $Y2=0.885
r189 1 74 182 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.235 $X2=2 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_4%VGND 1 2 3 4 5 6 7 22 24 28 32 34 38 40 44
+ 48 50 52 55 56 57 59 64 73 81 84 87 90 94
r126 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r127 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r128 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r129 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r130 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r131 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r132 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r133 76 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r134 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r135 73 93 3.95965 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=7.175 $Y=0
+ $X2=7.427 $Y2=0
r136 73 75 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.175 $Y=0
+ $X2=6.96 $Y2=0
r137 72 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r138 72 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r139 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r140 69 90 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.645 $Y=0 $X2=5.55
+ $Y2=0
r141 69 71 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.645 $Y=0 $X2=6
+ $Y2=0
r142 68 85 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r143 68 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r144 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r145 65 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r146 65 67 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=1.68 $Y2=0
r147 64 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.72
+ $Y2=0
r148 64 67 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=1.68 $Y2=0
r149 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r150 63 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r151 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r152 60 78 4.45492 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=0
+ $X2=0.207 $Y2=0
r153 60 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.415 $Y=0
+ $X2=0.72 $Y2=0
r154 59 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r155 59 62 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r156 57 88 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=4.56
+ $Y2=0
r157 57 85 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r158 55 71 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.315 $Y=0 $X2=6
+ $Y2=0
r159 55 56 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.315 $Y=0 $X2=6.41
+ $Y2=0
r160 54 75 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=6.96 $Y2=0
r161 54 56 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.505 $Y=0 $X2=6.41
+ $Y2=0
r162 50 93 3.25257 $w=2.6e-07 $l=1.58915e-07 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.427 $Y2=0
r163 50 52 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=7.305 $Y=0.085
+ $X2=7.305 $Y2=0.41
r164 46 56 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0
r165 46 48 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0.39
r166 42 90 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0
r167 42 44 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0.41
r168 41 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.785 $Y=0 $X2=4.655
+ $Y2=0
r169 40 90 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.455 $Y=0 $X2=5.55
+ $Y2=0
r170 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.455 $Y=0
+ $X2=4.785 $Y2=0
r171 36 87 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.655 $Y=0.085
+ $X2=4.655 $Y2=0
r172 36 38 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=4.655 $Y=0.085
+ $X2=4.655 $Y2=0.39
r173 35 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.72
+ $Y2=0
r174 34 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.525 $Y=0 $X2=4.655
+ $Y2=0
r175 34 35 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.525 $Y=0 $X2=3.885
+ $Y2=0
r176 30 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0
r177 30 32 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0.45
r178 26 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r179 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.38
r180 22 78 3.06275 $w=3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.207 $Y2=0
r181 22 24 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.38
r182 7 52 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=7.13
+ $Y=0.235 $X2=7.27 $Y2=0.41
r183 6 48 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=6.27
+ $Y=0.235 $X2=6.41 $Y2=0.39
r184 5 44 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=5.41
+ $Y=0.235 $X2=5.55 $Y2=0.41
r185 4 38 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.55
+ $Y=0.235 $X2=4.69 $Y2=0.39
r186 3 32 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=3.58
+ $Y=0.235 $X2=3.72 $Y2=0.45
r187 2 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1
+ $Y=0.235 $X2=1.14 $Y2=0.38
r188 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.235 $X2=0.28 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_4%A_114_47# 1 2 3 4 15 17 18 19 27
r33 25 27 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.43 $Y=0.42
+ $X2=3.29 $Y2=0.42
r34 23 30 2.73294 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=1.665 $Y=0.42
+ $X2=1.57 $Y2=0.42
r35 23 25 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.665 $Y=0.42
+ $X2=2.43 $Y2=0.42
r36 20 22 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.57 $Y=1.005
+ $X2=1.57 $Y2=0.95
r37 19 30 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=0.585
+ $X2=1.57 $Y2=0.42
r38 19 22 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=1.57 $Y=0.585
+ $X2=1.57 $Y2=0.95
r39 17 20 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.475 $Y=1.09
+ $X2=1.57 $Y2=1.005
r40 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.475 $Y=1.09
+ $X2=0.805 $Y2=1.09
r41 13 18 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.695 $Y=1.005
+ $X2=0.805 $Y2=1.09
r42 13 15 30.6445 $w=2.18e-07 $l=5.85e-07 $layer=LI1_cond $X=0.695 $Y=1.005
+ $X2=0.695 $Y2=0.42
r43 4 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.235 $X2=3.29 $Y2=0.42
r44 3 25 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.29
+ $Y=0.235 $X2=2.43 $Y2=0.42
r45 2 30 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.42
r46 2 22 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.95
r47 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.42
.ends

