* File: sky130_fd_sc_lp__isobufsrc_1.pxi.spice
* Created: Wed Sep  2 09:58:29 2020
* 
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_1%A N_A_M1002_g N_A_c_43_n N_A_M1003_g A A
+ PM_SKY130_FD_SC_LP__ISOBUFSRC_1%A
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_1%SLEEP N_SLEEP_M1004_g N_SLEEP_M1005_g SLEEP
+ N_SLEEP_c_68_n N_SLEEP_c_69_n PM_SKY130_FD_SC_LP__ISOBUFSRC_1%SLEEP
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_1%A_79_47# N_A_79_47#_M1002_s N_A_79_47#_M1003_s
+ N_A_79_47#_M1000_g N_A_79_47#_M1001_g N_A_79_47#_c_102_n N_A_79_47#_c_110_n
+ N_A_79_47#_c_103_n N_A_79_47#_c_104_n N_A_79_47#_c_105_n N_A_79_47#_c_106_n
+ N_A_79_47#_c_107_n N_A_79_47#_c_108_n PM_SKY130_FD_SC_LP__ISOBUFSRC_1%A_79_47#
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_1%VPWR N_VPWR_M1003_d N_VPWR_c_163_n VPWR
+ N_VPWR_c_164_n N_VPWR_c_165_n N_VPWR_c_162_n N_VPWR_c_167_n
+ PM_SKY130_FD_SC_LP__ISOBUFSRC_1%VPWR
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_1%X N_X_M1004_d N_X_M1000_d N_X_c_189_n
+ N_X_c_190_n N_X_c_193_n X X X X X X N_X_c_184_n X X
+ PM_SKY130_FD_SC_LP__ISOBUFSRC_1%X
x_PM_SKY130_FD_SC_LP__ISOBUFSRC_1%VGND N_VGND_M1002_d N_VGND_M1001_d
+ N_VGND_c_221_n N_VGND_c_222_n N_VGND_c_223_n N_VGND_c_224_n N_VGND_c_225_n
+ VGND N_VGND_c_226_n N_VGND_c_227_n PM_SKY130_FD_SC_LP__ISOBUFSRC_1%VGND
cc_1 VNB N_A_M1002_g 0.0577821f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.445
cc_2 VNB N_A_c_43_n 0.033798f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.675
cc_3 VNB A 0.0233953f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_SLEEP_M1004_g 0.0252435f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.445
cc_5 VNB N_SLEEP_c_68_n 0.0243624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_SLEEP_c_69_n 0.00185986f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.51
cc_7 VNB N_A_79_47#_M1000_g 0.00696454f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_A_79_47#_c_102_n 0.0362414f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.587
cc_9 VNB N_A_79_47#_c_103_n 0.0160786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_79_47#_c_104_n 0.00968934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_79_47#_c_105_n 8.3509e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_79_47#_c_106_n 0.00914334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_79_47#_c_107_n 0.0335936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_79_47#_c_108_n 0.0187964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_162_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_X_c_184_n 0.0110339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB X 0.0370578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_221_n 0.00424491f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_VGND_c_222_n 0.0146919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_223_n 0.0160508f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.51
cc_21 VNB N_VGND_c_224_n 0.0240173f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.587
cc_22 VNB N_VGND_c_225_n 0.00701746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_226_n 0.0148157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_227_n 0.160429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VPB N_A_c_43_n 0.00889775f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.675
cc_26 VPB N_A_M1003_g 0.0317374f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=2.045
cc_27 VPB A 0.0198536f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_28 VPB N_SLEEP_M1005_g 0.0204408f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=2.045
cc_29 VPB N_SLEEP_c_68_n 0.00638147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_SLEEP_c_69_n 0.00269256f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.51
cc_31 VPB N_A_79_47#_M1000_g 0.0219297f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_32 VPB N_A_79_47#_c_110_n 0.0109886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_A_79_47#_c_105_n 0.00137696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_163_n 0.0312943f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=2.045
cc_35 VPB N_VPWR_c_164_n 0.0326924f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_36 VPB N_VPWR_c_165_n 0.0327687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_162_n 0.079895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_167_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB X 0.0125749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB X 0.00849495f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB X 0.0427581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 N_A_M1002_g N_SLEEP_M1004_g 0.0210846f $X=0.735 $Y=0.445 $X2=0 $Y2=0
cc_43 N_A_M1003_g N_SLEEP_M1005_g 0.0202207f $X=0.8 $Y=2.045 $X2=0 $Y2=0
cc_44 N_A_c_43_n N_SLEEP_c_68_n 0.0188044f $X=0.8 $Y=1.675 $X2=0 $Y2=0
cc_45 A N_SLEEP_c_68_n 5.15864e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_46 N_A_c_43_n N_SLEEP_c_69_n 0.0017587f $X=0.8 $Y=1.675 $X2=0 $Y2=0
cc_47 A N_SLEEP_c_69_n 0.0278008f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_48 N_A_M1002_g N_A_79_47#_c_102_n 0.0132293f $X=0.735 $Y=0.445 $X2=0 $Y2=0
cc_49 N_A_c_43_n N_A_79_47#_c_110_n 0.00135528f $X=0.8 $Y=1.675 $X2=0 $Y2=0
cc_50 N_A_M1003_g N_A_79_47#_c_110_n 0.0145687f $X=0.8 $Y=2.045 $X2=0 $Y2=0
cc_51 A N_A_79_47#_c_110_n 0.032229f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_52 N_A_M1002_g N_A_79_47#_c_103_n 0.016819f $X=0.735 $Y=0.445 $X2=0 $Y2=0
cc_53 N_A_c_43_n N_A_79_47#_c_103_n 0.0014324f $X=0.8 $Y=1.675 $X2=0 $Y2=0
cc_54 A N_A_79_47#_c_103_n 0.0176433f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_55 N_A_c_43_n N_A_79_47#_c_104_n 0.00385139f $X=0.8 $Y=1.675 $X2=0 $Y2=0
cc_56 A N_A_79_47#_c_104_n 0.0232392f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_57 N_A_M1003_g N_VPWR_c_163_n 0.0020569f $X=0.8 $Y=2.045 $X2=0 $Y2=0
cc_58 N_A_M1002_g N_VGND_c_221_n 0.0186229f $X=0.735 $Y=0.445 $X2=0 $Y2=0
cc_59 N_A_M1002_g N_VGND_c_224_n 0.00525069f $X=0.735 $Y=0.445 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_VGND_c_227_n 0.0101608f $X=0.735 $Y=0.445 $X2=0 $Y2=0
cc_61 N_SLEEP_c_68_n N_A_79_47#_M1000_g 0.0622505f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_62 N_SLEEP_M1005_g N_A_79_47#_c_110_n 0.0163944f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_63 N_SLEEP_c_68_n N_A_79_47#_c_110_n 9.45883e-19 $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_64 N_SLEEP_c_69_n N_A_79_47#_c_110_n 0.0269704f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_65 N_SLEEP_M1004_g N_A_79_47#_c_103_n 0.0142735f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_66 N_SLEEP_c_68_n N_A_79_47#_c_103_n 0.00443399f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_67 N_SLEEP_c_69_n N_A_79_47#_c_103_n 0.0281593f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_68 N_SLEEP_c_68_n N_A_79_47#_c_105_n 0.00372476f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_69 N_SLEEP_M1004_g N_A_79_47#_c_106_n 0.00387666f $X=1.34 $Y=0.655 $X2=0
+ $Y2=0
cc_70 N_SLEEP_c_69_n N_A_79_47#_c_106_n 0.0249209f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_71 N_SLEEP_M1004_g N_A_79_47#_c_107_n 0.0622505f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_72 N_SLEEP_c_69_n N_A_79_47#_c_107_n 3.76098e-19 $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_73 N_SLEEP_M1004_g N_A_79_47#_c_108_n 0.0146764f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_74 N_SLEEP_M1005_g N_VPWR_c_163_n 0.0236468f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_75 N_SLEEP_M1005_g N_VPWR_c_165_n 0.00486043f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_76 N_SLEEP_M1005_g N_VPWR_c_162_n 0.00818711f $X=1.34 $Y=2.465 $X2=0 $Y2=0
cc_77 N_SLEEP_M1004_g N_X_c_189_n 0.00210081f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_78 N_SLEEP_M1004_g N_X_c_190_n 0.00544733f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_79 N_SLEEP_M1004_g N_VGND_c_221_n 0.00386418f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_80 N_SLEEP_M1004_g N_VGND_c_223_n 4.78045e-19 $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_81 N_SLEEP_M1004_g N_VGND_c_226_n 0.0054895f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_82 N_SLEEP_M1004_g N_VGND_c_227_n 0.0103177f $X=1.34 $Y=0.655 $X2=0 $Y2=0
cc_83 N_A_79_47#_c_110_n N_VPWR_M1003_d 0.00781403f $X=1.585 $Y=2.03 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_79_47#_M1000_g N_VPWR_c_163_n 0.00351016f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_79_47#_c_110_n N_VPWR_c_163_n 0.0223387f $X=1.585 $Y=2.03 $X2=0 $Y2=0
cc_86 N_A_79_47#_M1000_g N_VPWR_c_165_n 0.00585385f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_79_47#_M1000_g N_VPWR_c_162_n 0.0119837f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_88 N_A_79_47#_c_110_n A_283_367# 0.00569383f $X=1.585 $Y=2.03 $X2=-0.19
+ $Y2=-0.245
cc_89 N_A_79_47#_c_103_n N_X_c_189_n 0.0133344f $X=1.585 $Y=1.17 $X2=0 $Y2=0
cc_90 N_A_79_47#_c_106_n N_X_c_189_n 0.00533216f $X=1.735 $Y=1.17 $X2=0 $Y2=0
cc_91 N_A_79_47#_c_106_n N_X_c_193_n 0.0149345f $X=1.735 $Y=1.17 $X2=0 $Y2=0
cc_92 N_A_79_47#_c_107_n N_X_c_193_n 0.00211584f $X=1.79 $Y=1.35 $X2=0 $Y2=0
cc_93 N_A_79_47#_c_108_n N_X_c_193_n 0.0116558f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_94 N_A_79_47#_M1000_g X 0.0328587f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A_79_47#_c_110_n X 0.0183112f $X=1.585 $Y=2.03 $X2=0 $Y2=0
cc_96 N_A_79_47#_c_105_n X 0.00787294f $X=1.67 $Y=1.92 $X2=0 $Y2=0
cc_97 N_A_79_47#_c_107_n X 0.00112164f $X=1.79 $Y=1.35 $X2=0 $Y2=0
cc_98 N_A_79_47#_M1000_g X 0.00547213f $X=1.7 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_79_47#_c_105_n X 0.0145256f $X=1.67 $Y=1.92 $X2=0 $Y2=0
cc_100 N_A_79_47#_c_106_n X 0.0335658f $X=1.735 $Y=1.17 $X2=0 $Y2=0
cc_101 N_A_79_47#_c_107_n X 0.00812269f $X=1.79 $Y=1.35 $X2=0 $Y2=0
cc_102 N_A_79_47#_c_108_n X 0.00650334f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_103 N_A_79_47#_c_102_n N_VGND_c_221_n 0.0350253f $X=0.52 $Y=0.45 $X2=0 $Y2=0
cc_104 N_A_79_47#_c_103_n N_VGND_c_221_n 0.0346938f $X=1.585 $Y=1.17 $X2=0 $Y2=0
cc_105 N_A_79_47#_c_108_n N_VGND_c_223_n 0.00919683f $X=1.79 $Y=1.185 $X2=0
+ $Y2=0
cc_106 N_A_79_47#_c_102_n N_VGND_c_224_n 0.0152359f $X=0.52 $Y=0.45 $X2=0 $Y2=0
cc_107 N_A_79_47#_c_108_n N_VGND_c_226_n 0.00366311f $X=1.79 $Y=1.185 $X2=0
+ $Y2=0
cc_108 N_A_79_47#_M1002_s N_VGND_c_227_n 0.00342267f $X=0.395 $Y=0.235 $X2=0
+ $Y2=0
cc_109 N_A_79_47#_c_102_n N_VGND_c_227_n 0.0102663f $X=0.52 $Y=0.45 $X2=0 $Y2=0
cc_110 N_A_79_47#_c_108_n N_VGND_c_227_n 0.00436859f $X=1.79 $Y=1.185 $X2=0
+ $Y2=0
cc_111 N_VPWR_c_162_n A_283_367# 0.00899413f $X=2.16 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_112 N_VPWR_c_162_n N_X_M1000_d 0.00929756f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_113 N_VPWR_c_163_n X 0.0211817f $X=1.125 $Y=2.42 $X2=0 $Y2=0
cc_114 N_VPWR_c_165_n X 0.0273486f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_115 N_VPWR_c_162_n X 0.0150845f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_116 N_X_c_193_n N_VGND_M1001_d 0.00629056f $X=2.055 $Y=0.83 $X2=0 $Y2=0
cc_117 N_X_c_184_n N_VGND_M1001_d 0.00111246f $X=2.185 $Y=0.915 $X2=0 $Y2=0
cc_118 X N_VGND_M1001_d 0.00244175f $X=2.16 $Y=0.925 $X2=0 $Y2=0
cc_119 N_X_c_184_n N_VGND_c_222_n 0.00270734f $X=2.185 $Y=0.915 $X2=0 $Y2=0
cc_120 N_X_c_193_n N_VGND_c_223_n 0.0137194f $X=2.055 $Y=0.83 $X2=0 $Y2=0
cc_121 N_X_c_184_n N_VGND_c_223_n 0.00829742f $X=2.185 $Y=0.915 $X2=0 $Y2=0
cc_122 N_X_c_190_n N_VGND_c_226_n 0.0156591f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_123 N_X_c_193_n N_VGND_c_226_n 0.00191958f $X=2.055 $Y=0.83 $X2=0 $Y2=0
cc_124 N_X_M1004_d N_VGND_c_227_n 0.00245675f $X=1.415 $Y=0.235 $X2=0 $Y2=0
cc_125 N_X_c_190_n N_VGND_c_227_n 0.00983963f $X=1.555 $Y=0.42 $X2=0 $Y2=0
cc_126 N_X_c_193_n N_VGND_c_227_n 0.00467209f $X=2.055 $Y=0.83 $X2=0 $Y2=0
cc_127 N_X_c_184_n N_VGND_c_227_n 0.00505278f $X=2.185 $Y=0.915 $X2=0 $Y2=0
