* File: sky130_fd_sc_lp__a31o_1.pex.spice
* Created: Fri Aug 28 09:59:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31O_1%A_80_21# 1 2 9 12 16 17 19 20 23 25 29 33 35
+ 36 39
r74 35 37 1.41596 $w=4.33e-07 $l=5e-09 $layer=LI1_cond $X=3.047 $Y=1.98
+ $X2=3.047 $Y2=1.985
r75 35 36 8.80985 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=3.047 $Y=1.98
+ $X2=3.047 $Y2=1.815
r76 31 36 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.18 $Y=1.04
+ $X2=3.18 $Y2=1.815
r77 29 37 36.759 $w=2.88e-07 $l=9.25e-07 $layer=LI1_cond $X=2.975 $Y=2.91
+ $X2=2.975 $Y2=1.985
r78 26 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.62 $Y=0.955
+ $X2=2.455 $Y2=0.955
r79 25 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.095 $Y=0.955
+ $X2=3.18 $Y2=1.04
r80 25 26 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.095 $Y=0.955
+ $X2=2.62 $Y2=0.955
r81 21 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.455 $Y=0.87
+ $X2=2.455 $Y2=0.955
r82 21 23 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.455 $Y=0.87
+ $X2=2.455 $Y2=0.42
r83 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=0.955
+ $X2=2.455 $Y2=0.955
r84 19 20 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=2.29 $Y=0.955
+ $X2=0.765 $Y2=0.955
r85 17 40 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.582 $Y=1.35
+ $X2=0.582 $Y2=1.515
r86 17 39 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.582 $Y=1.35
+ $X2=0.582 $Y2=1.185
r87 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.35 $X2=0.6 $Y2=1.35
r88 14 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.64 $Y=1.04
+ $X2=0.765 $Y2=0.955
r89 14 16 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.64 $Y=1.04
+ $X2=0.64 $Y2=1.35
r90 12 40 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.515 $Y=2.465
+ $X2=0.515 $Y2=1.515
r91 9 39 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.655
+ $X2=0.475 $Y2=1.185
r92 2 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=1.835 $X2=2.955 $Y2=1.98
r93 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.815
+ $Y=1.835 $X2=2.955 $Y2=2.91
r94 1 23 91 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=2 $X=2.275
+ $Y=0.235 $X2=2.455 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_1%A3 3 7 9 10 11 12 13 21 25 27
c43 27 0 1.17581e-19 $X=1.2 $Y=1.665
r44 25 27 1.16746 $w=1.88e-07 $l=2e-08 $layer=LI1_cond $X=1.19 $Y=1.645 $X2=1.19
+ $Y2=1.665
r45 21 24 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.375
+ $X2=1.16 $Y2=1.54
r46 21 23 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.375
+ $X2=1.16 $Y2=1.21
r47 12 13 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=2.405
+ $X2=1.19 $Y2=2.775
r48 11 12 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=2.035
+ $X2=1.19 $Y2=2.405
r49 10 25 3.75361 $w=3.55e-07 $l=4.55961e-08 $layer=LI1_cond $X=1.16 $Y=1.612
+ $X2=1.19 $Y2=1.645
r50 10 11 19.7301 $w=1.88e-07 $l=3.38e-07 $layer=LI1_cond $X=1.19 $Y=1.697
+ $X2=1.19 $Y2=2.035
r51 10 27 1.86794 $w=1.88e-07 $l=3.2e-08 $layer=LI1_cond $X=1.19 $Y=1.697
+ $X2=1.19 $Y2=1.665
r52 9 10 10.8941 $w=3.55e-07 $l=3.17e-07 $layer=LI1_cond $X=1.16 $Y=1.295
+ $X2=1.16 $Y2=1.612
r53 9 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.375 $X2=1.18 $Y2=1.375
r54 7 24 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.27 $Y=2.465
+ $X2=1.27 $Y2=1.54
r55 3 23 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.27 $Y=0.655
+ $X2=1.27 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_1%A2 3 6 8 11 13
r38 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.72 $Y=1.35
+ $X2=1.72 $Y2=1.515
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.72 $Y=1.35
+ $X2=1.72 $Y2=1.185
r40 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.35 $X2=1.72 $Y2=1.35
r41 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.755 $Y=2.465
+ $X2=1.755 $Y2=1.515
r42 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.66 $Y=0.655
+ $X2=1.66 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_1%A1 3 7 9 12 13
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.375
+ $X2=2.29 $Y2=1.54
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.375
+ $X2=2.29 $Y2=1.21
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.375 $X2=2.29 $Y2=1.375
r37 9 13 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.16 $Y=1.375
+ $X2=2.29 $Y2=1.375
r38 7 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.31 $Y=2.465
+ $X2=2.31 $Y2=1.54
r39 3 14 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.2 $Y=0.655 $X2=2.2
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_1%B1 3 7 9 12 13
r29 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.375
+ $X2=2.83 $Y2=1.54
r30 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.375
+ $X2=2.83 $Y2=1.21
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.83
+ $Y=1.375 $X2=2.83 $Y2=1.375
r32 9 13 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.64 $Y=1.375
+ $X2=2.83 $Y2=1.375
r33 7 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.74 $Y=2.465
+ $X2=2.74 $Y2=1.54
r34 3 14 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.74 $Y=0.655
+ $X2=2.74 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_1%X 1 2 7 8 9 10 11 12 13 24 34
r16 34 47 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=0.215 $Y=1.665
+ $X2=0.215 $Y2=1.695
r17 13 44 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=0.245 $Y=2.775
+ $X2=0.245 $Y2=2.91
r18 12 13 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.245 $Y=2.405
+ $X2=0.245 $Y2=2.775
r19 11 12 15.3059 $w=3.18e-07 $l=4.25e-07 $layer=LI1_cond $X=0.245 $Y=1.98
+ $X2=0.245 $Y2=2.405
r20 11 35 4.50173 $w=3.18e-07 $l=1.25e-07 $layer=LI1_cond $X=0.245 $Y=1.98
+ $X2=0.245 $Y2=1.855
r21 10 35 4.78984 $w=3.18e-07 $l=1.33e-07 $layer=LI1_cond $X=0.245 $Y=1.722
+ $X2=0.245 $Y2=1.855
r22 10 47 1.41141 $w=3.18e-07 $l=2.7e-08 $layer=LI1_cond $X=0.245 $Y=1.722
+ $X2=0.245 $Y2=1.695
r23 10 34 1.24109 $w=2.58e-07 $l=2.8e-08 $layer=LI1_cond $X=0.215 $Y=1.637
+ $X2=0.215 $Y2=1.665
r24 9 10 15.1591 $w=2.58e-07 $l=3.42e-07 $layer=LI1_cond $X=0.215 $Y=1.295
+ $X2=0.215 $Y2=1.637
r25 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=0.925
+ $X2=0.215 $Y2=1.295
r26 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=0.555
+ $X2=0.215 $Y2=0.925
r27 7 24 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.215 $Y=0.555
+ $X2=0.215 $Y2=0.42
r28 2 44 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.835 $X2=0.3 $Y2=2.91
r29 2 11 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.835 $X2=0.3 $Y2=1.98
r30 1 24 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_1%VPWR 1 2 9 15 19 21 26 33 34 37 40
r45 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 34 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 31 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.03 $Y2=3.33
r50 31 33 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 27 37 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.775 $Y2=3.33
r52 27 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=2.03 $Y2=3.33
r54 26 29 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 24 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 21 37 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.775 $Y2=3.33
r58 21 23 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 19 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 19 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 19 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 15 18 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=2.03 $Y=2.135
+ $X2=2.03 $Y2=2.95
r63 13 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=3.33
r64 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=2.95
r65 9 12 37.2623 $w=2.98e-07 $l=9.7e-07 $layer=LI1_cond $X=0.775 $Y=1.98
+ $X2=0.775 $Y2=2.95
r66 7 37 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=3.245
+ $X2=0.775 $Y2=3.33
r67 7 12 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.775 $Y=3.245
+ $X2=0.775 $Y2=2.95
r68 2 18 400 $w=1.7e-07 $l=1.21088e-06 $layer=licon1_PDIFF $count=1 $X=1.83
+ $Y=1.835 $X2=2.03 $Y2=2.95
r69 2 15 400 $w=1.7e-07 $l=3.87298e-07 $layer=licon1_PDIFF $count=1 $X=1.83
+ $Y=1.835 $X2=2.03 $Y2=2.135
r70 1 12 400 $w=1.7e-07 $l=1.22005e-06 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.835 $X2=0.81 $Y2=2.95
r71 1 9 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.835 $X2=0.81 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_1%A_269_367# 1 2 9 13 14 17
r35 17 19 36.3313 $w=2.93e-07 $l=9.3e-07 $layer=LI1_cond $X=2.512 $Y=1.98
+ $X2=2.512 $Y2=2.91
r36 15 17 3.90659 $w=2.93e-07 $l=1e-07 $layer=LI1_cond $X=2.512 $Y=1.88
+ $X2=2.512 $Y2=1.98
r37 13 15 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=2.365 $Y=1.795
+ $X2=2.512 $Y2=1.88
r38 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.365 $Y=1.795
+ $X2=1.695 $Y2=1.795
r39 9 11 44.6572 $w=2.38e-07 $l=9.3e-07 $layer=LI1_cond $X=1.575 $Y=1.98
+ $X2=1.575 $Y2=2.91
r40 7 14 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.575 $Y=1.88
+ $X2=1.695 $Y2=1.795
r41 7 9 4.80185 $w=2.38e-07 $l=1e-07 $layer=LI1_cond $X=1.575 $Y=1.88 $X2=1.575
+ $Y2=1.98
r42 2 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.835 $X2=2.525 $Y2=2.91
r43 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.835 $X2=2.525 $Y2=1.98
r44 1 11 400 $w=1.7e-07 $l=1.16844e-06 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=1.835 $X2=1.54 $Y2=2.91
r45 1 9 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=1.345
+ $Y=1.835 $X2=1.54 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_1%VGND 1 2 7 9 11 13 18 34
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r36 26 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r37 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r38 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 19 21 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=1.22 $Y=0 $X2=2.64
+ $Y2=0
r40 18 33 4.51706 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=3.075
+ $Y2=0
r41 18 21 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.64
+ $Y2=0
r42 16 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r43 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 13 30 9.89561 $w=6.93e-07 $l=5.75e-07 $layer=LI1_cond $X=0.872 $Y=0
+ $X2=0.872 $Y2=0.575
r45 13 19 9.27432 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=0.872 $Y=0 $X2=1.22
+ $Y2=0
r46 13 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 13 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 13 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r49 11 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 11 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r51 7 33 3.24911 $w=3.3e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=3.075 $Y2=0
r52 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0.575
r53 2 9 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.235 $X2=2.955 $Y2=0.575
r54 1 30 91 $w=1.7e-07 $l=6.53242e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=1.055 $Y2=0.575
.ends

