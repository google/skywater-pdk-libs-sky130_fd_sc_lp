* File: sky130_fd_sc_lp__o2bb2a_2.pex.spice
* Created: Wed Sep  2 10:21:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%B1 3 7 11 12 13 16
r29 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.16 $X2=0.585 $Y2=1.16
r30 13 17 2.41001 $w=6.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.33
+ $X2=0.585 $Y2=1.33
r31 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.585 $Y=1.5
+ $X2=0.585 $Y2=1.16
r32 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.5
+ $X2=0.585 $Y2=1.665
r33 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=0.995
+ $X2=0.585 $Y2=1.16
r34 7 12 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.675 $Y=2.155
+ $X2=0.675 $Y2=1.665
r35 3 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.675 $Y=0.445
+ $X2=0.675 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%B2 3 7 11 12 13 16
c38 13 0 1.02291e-19 $X=1.2 $Y=1.295
r39 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.125
+ $Y=1.16 $X2=1.125 $Y2=1.16
r40 13 17 1.33889 $w=6.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.2 $Y=1.33
+ $X2=1.125 $Y2=1.33
r41 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.125 $Y=1.5
+ $X2=1.125 $Y2=1.16
r42 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.125 $Y=1.5
+ $X2=1.125 $Y2=1.665
r43 10 16 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.125 $Y=0.995
+ $X2=1.125 $Y2=1.16
r44 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.145 $Y=0.445
+ $X2=1.145 $Y2=0.995
r45 3 12 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.035 $Y=2.155
+ $X2=1.035 $Y2=1.665
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%A_300_21# 1 2 9 13 16 17 20 24 28 30
c69 20 0 1.40662e-19 $X=1.98 $Y=1.5
c70 9 0 1.55732e-19 $X=1.575 $Y=0.445
r71 26 30 4.59179 $w=2.87e-07 $l=1.66958e-07 $layer=LI1_cond $X=2.76 $Y=1.585
+ $X2=2.662 $Y2=1.46
r72 26 28 23.0574 $w=1.88e-07 $l=3.95e-07 $layer=LI1_cond $X=2.76 $Y=1.585
+ $X2=2.76 $Y2=1.98
r73 22 30 4.59179 $w=2.87e-07 $l=1.25e-07 $layer=LI1_cond $X=2.662 $Y=1.335
+ $X2=2.662 $Y2=1.46
r74 22 24 26.6409 $w=3.83e-07 $l=8.9e-07 $layer=LI1_cond $X=2.662 $Y=1.335
+ $X2=2.662 $Y2=0.445
r75 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.98
+ $Y=1.5 $X2=1.98 $Y2=1.5
r76 17 30 1.85035 $w=2.5e-07 $l=1.92e-07 $layer=LI1_cond $X=2.47 $Y=1.46
+ $X2=2.662 $Y2=1.46
r77 17 19 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=2.47 $Y=1.46
+ $X2=1.98 $Y2=1.46
r78 15 20 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.65 $Y=1.5 $X2=1.98
+ $Y2=1.5
r79 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.65 $Y=1.5
+ $X2=1.575 $Y2=1.5
r80 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.575 $Y=1.665
+ $X2=1.575 $Y2=1.5
r81 11 13 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.575 $Y=1.665
+ $X2=1.575 $Y2=2.155
r82 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.575 $Y=1.335
+ $X2=1.575 $Y2=1.5
r83 7 9 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.575 $Y=1.335
+ $X2=1.575 $Y2=0.445
r84 2 28 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.63
+ $Y=1.835 $X2=2.77 $Y2=1.98
r85 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.51
+ $Y=0.235 $X2=2.635 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%A2_N 3 5 7 8 9 11 12
c44 11 0 1.55732e-19 $X=2.16 $Y=0.555
r45 12 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.205
+ $Y=0.93 $X2=2.205 $Y2=0.93
r46 11 12 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.182 $Y=0.555
+ $X2=2.182 $Y2=0.925
r47 9 10 67.7095 $w=2.1e-07 $l=2.95e-07 $layer=POLY_cond $X=2.555 $Y=0.915
+ $X2=2.85 $Y2=0.915
r48 8 16 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=2.48 $Y=0.93
+ $X2=2.205 $Y2=0.93
r49 8 9 17.3036 $w=3.3e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.48 $Y=0.93
+ $X2=2.555 $Y2=0.915
r50 5 10 10.701 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.85 $Y=0.765 $X2=2.85
+ $Y2=0.915
r51 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.85 $Y=0.765 $X2=2.85
+ $Y2=0.445
r52 1 9 10.701 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.555 $Y=1.095
+ $X2=2.555 $Y2=0.915
r53 1 3 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=2.555 $Y=1.095
+ $X2=2.555 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%A1_N 3 7 9 10 11 20
r43 18 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.12 $Y=1.35 $X2=3.21
+ $Y2=1.35
r44 15 18 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.985 $Y=1.35
+ $X2=3.12 $Y2=1.35
r45 11 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.35 $X2=3.12 $Y2=1.35
r46 10 11 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=0.925
+ $X2=3.13 $Y2=1.295
r47 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=0.555
+ $X2=3.13 $Y2=0.925
r48 5 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.185
+ $X2=3.21 $Y2=1.35
r49 5 7 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.21 $Y=1.185 $X2=3.21
+ $Y2=0.445
r50 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.985 $Y=1.515
+ $X2=2.985 $Y2=1.35
r51 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.985 $Y=1.515
+ $X2=2.985 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%A_222_367# 1 2 7 9 12 14 16 19 23 26 27 29
+ 31 34 35 36 38 39 40 43 46 54
c127 46 0 1.40662e-19 $X=1.14 $Y=1.835
r128 53 54 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.795 $Y=1.35
+ $X2=4.225 $Y2=1.35
r129 44 53 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.66 $Y=1.35
+ $X2=3.795 $Y2=1.35
r130 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=1.35 $X2=3.66 $Y2=1.35
r131 41 43 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.62 $Y=1.685
+ $X2=3.62 $Y2=1.35
r132 39 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.495 $Y=1.77
+ $X2=3.62 $Y2=1.685
r133 39 40 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.495 $Y=1.77
+ $X2=3.205 $Y2=1.77
r134 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.12 $Y=1.855
+ $X2=3.205 $Y2=1.77
r135 37 38 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.12 $Y=1.855
+ $X2=3.12 $Y2=2.665
r136 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.035 $Y=2.75
+ $X2=3.12 $Y2=2.665
r137 35 36 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.035 $Y=2.75
+ $X2=2.495 $Y2=2.75
r138 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.41 $Y=2.665
+ $X2=2.495 $Y2=2.75
r139 33 34 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.41 $Y=1.925
+ $X2=2.41 $Y2=2.665
r140 29 47 14.4834 $w=1.68e-07 $l=2.22e-07 $layer=LI1_cond $X=1.777 $Y=1.08
+ $X2=1.555 $Y2=1.08
r141 29 31 26.9721 $w=2.33e-07 $l=5.5e-07 $layer=LI1_cond $X=1.777 $Y=0.995
+ $X2=1.777 $Y2=0.445
r142 28 46 4.00616 $w=1.7e-07 $l=5.17494e-07 $layer=LI1_cond $X=1.655 $Y=1.84
+ $X2=1.14 $Y2=1.835
r143 27 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.325 $Y=1.84
+ $X2=2.41 $Y2=1.925
r144 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.325 $Y=1.84
+ $X2=1.655 $Y2=1.84
r145 26 46 2.75409 $w=3.47e-07 $l=4.53238e-07 $layer=LI1_cond $X=1.555 $Y=1.755
+ $X2=1.14 $Y2=1.835
r146 25 47 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=1.165
+ $X2=1.555 $Y2=1.08
r147 25 26 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=1.555 $Y=1.165
+ $X2=1.555 $Y2=1.755
r148 21 46 2.75409 $w=3.47e-07 $l=2.98629e-07 $layer=LI1_cond $X=1.397 $Y=1.925
+ $X2=1.14 $Y2=1.835
r149 21 23 1.27737 $w=5.13e-07 $l=5.5e-08 $layer=LI1_cond $X=1.397 $Y=1.925
+ $X2=1.397 $Y2=1.98
r150 17 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.225 $Y=1.515
+ $X2=4.225 $Y2=1.35
r151 17 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.225 $Y=1.515
+ $X2=4.225 $Y2=2.465
r152 14 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.225 $Y=1.185
+ $X2=4.225 $Y2=1.35
r153 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.225 $Y=1.185
+ $X2=4.225 $Y2=0.655
r154 10 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.515
+ $X2=3.795 $Y2=1.35
r155 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.795 $Y=1.515
+ $X2=3.795 $Y2=2.465
r156 7 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.185
+ $X2=3.795 $Y2=1.35
r157 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.795 $Y=1.185
+ $X2=3.795 $Y2=0.655
r158 2 23 300 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.835 $X2=1.305 $Y2=1.98
r159 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=0.235 $X2=1.79 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%VPWR 1 2 3 4 15 19 23 27 29 34 35 37 38 39
+ 50 57 63 67
r58 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 61 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 61 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r62 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 58 63 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.56 $Y2=3.33
r64 58 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 57 66 3.9252 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.577 $Y2=3.33
r66 57 60 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 56 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r68 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r69 52 55 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r70 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 50 63 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.56 $Y2=3.33
r72 50 55 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 49 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r77 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r80 39 56 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r81 39 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 37 48 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.99 $Y2=3.33
r84 36 52 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=2.16 $Y2=3.33
r85 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=1.99 $Y2=3.33
r86 34 42 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=0.295 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.295 $Y=3.33
+ $X2=0.46 $Y2=3.33
r88 33 45 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.72 $Y2=3.33
r89 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.46 $Y2=3.33
r90 29 32 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=4.48 $Y=1.98
+ $X2=4.48 $Y2=2.95
r91 27 66 3.21796 $w=2.5e-07 $l=1.32868e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.577 $Y2=3.33
r92 27 32 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=2.95
r93 23 26 13.2375 $w=3.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.56 $Y=2.11
+ $X2=3.56 $Y2=2.535
r94 21 63 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=3.33
r95 21 26 22.1144 $w=3.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=2.535
r96 17 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=3.33
r97 17 19 35.7956 $w=3.28e-07 $l=1.025e-06 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=2.22
r98 13 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.46 $Y=3.245
+ $X2=0.46 $Y2=3.33
r99 13 15 44.177 $w=3.28e-07 $l=1.265e-06 $layer=LI1_cond $X=0.46 $Y=3.245
+ $X2=0.46 $Y2=1.98
r100 4 32 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.3
+ $Y=1.835 $X2=4.44 $Y2=2.95
r101 4 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.3
+ $Y=1.835 $X2=4.44 $Y2=1.98
r102 3 26 300 $w=1.7e-07 $l=9.24121e-07 $layer=licon1_PDIFF $count=2 $X=3.06
+ $Y=1.835 $X2=3.58 $Y2=2.535
r103 3 23 600 $w=1.7e-07 $l=6.01997e-07 $layer=licon1_PDIFF $count=1 $X=3.06
+ $Y=1.835 $X2=3.54 $Y2=2.11
r104 2 19 600 $w=1.7e-07 $l=5.28323e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.835 $X2=1.99 $Y2=2.22
r105 1 15 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.335
+ $Y=1.835 $X2=0.46 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%X 1 2 7 8 9 10 11 12 13 22
r17 13 40 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.05 $Y=2.775
+ $X2=4.05 $Y2=2.91
r18 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.05 $Y=2.405
+ $X2=4.05 $Y2=2.775
r19 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.05 $Y=1.98
+ $X2=4.05 $Y2=2.405
r20 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.05 $Y=1.665
+ $X2=4.05 $Y2=1.98
r21 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.05 $Y=1.295
+ $X2=4.05 $Y2=1.665
r22 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.05 $Y=0.925 $X2=4.05
+ $Y2=1.295
r23 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.05 $Y=0.555 $X2=4.05
+ $Y2=0.925
r24 7 22 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.05 $Y=0.555
+ $X2=4.05 $Y2=0.42
r25 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.835 $X2=4.01 $Y2=2.91
r26 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.835 $X2=4.01 $Y2=1.98
r27 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.87
+ $Y=0.235 $X2=4.01 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%A_67_47# 1 2 9 11 12 15
r24 13 15 9.87808 $w=2.43e-07 $l=2.1e-07 $layer=LI1_cond $X=1.367 $Y=0.655
+ $X2=1.367 $Y2=0.445
r25 11 13 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=1.245 $Y=0.74
+ $X2=1.367 $Y2=0.655
r26 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.245 $Y=0.74
+ $X2=0.575 $Y2=0.74
r27 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.435 $Y=0.655
+ $X2=0.575 $Y2=0.74
r28 7 9 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=0.435 $Y=0.655
+ $X2=0.435 $Y2=0.445
r29 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.22
+ $Y=0.235 $X2=1.36 $Y2=0.445
r30 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.335
+ $Y=0.235 $X2=0.46 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_2%VGND 1 2 3 12 16 20 22 25 26 27 33 40 46 50
r63 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r64 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r65 44 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r66 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r67 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r68 41 46 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=3.575
+ $Y2=0
r69 41 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.745 $Y=0 $X2=4.08
+ $Y2=0
r70 40 49 3.9252 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.577
+ $Y2=0
r71 40 43 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.08
+ $Y2=0
r72 39 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r73 38 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r74 35 38 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r75 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r76 33 46 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.575
+ $Y2=0
r77 33 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.12
+ $Y2=0
r78 31 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r79 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r80 27 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r81 27 36 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r82 25 30 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=0 $X2=0.72
+ $Y2=0
r83 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.745 $Y=0 $X2=0.91
+ $Y2=0
r84 24 35 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=1.2
+ $Y2=0
r85 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=0.91
+ $Y2=0
r86 20 49 3.21796 $w=2.5e-07 $l=1.32868e-07 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.577 $Y2=0
r87 20 22 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.48 $Y=0.085
+ $X2=4.48 $Y2=0.38
r88 16 18 15.9308 $w=3.38e-07 $l=4.7e-07 $layer=LI1_cond $X=3.575 $Y=0.38
+ $X2=3.575 $Y2=0.85
r89 14 46 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0
r90 14 16 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0.38
r91 10 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.91 $Y=0.085
+ $X2=0.91 $Y2=0
r92 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.91 $Y=0.085
+ $X2=0.91 $Y2=0.38
r93 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.3
+ $Y=0.235 $X2=4.44 $Y2=0.38
r94 2 18 182 $w=1.7e-07 $l=7.48098e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.58 $Y2=0.85
r95 2 16 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.51 $Y2=0.38
r96 1 12 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.75
+ $Y=0.235 $X2=0.91 $Y2=0.38
.ends

