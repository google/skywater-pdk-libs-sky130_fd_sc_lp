* File: sky130_fd_sc_lp__a21o_lp.pxi.spice
* Created: Wed Sep  2 09:20:14 2020
* 
x_PM_SKY130_FD_SC_LP__A21O_LP%A2 N_A2_M1003_g N_A2_M1006_g A2 A2 N_A2_c_61_n
+ N_A2_c_62_n PM_SKY130_FD_SC_LP__A21O_LP%A2
x_PM_SKY130_FD_SC_LP__A21O_LP%A1 N_A1_M1005_g N_A1_c_89_n N_A1_M1008_g
+ N_A1_c_90_n A1 A1 N_A1_c_91_n N_A1_c_92_n PM_SKY130_FD_SC_LP__A21O_LP%A1
x_PM_SKY130_FD_SC_LP__A21O_LP%B1 N_B1_M1001_g N_B1_M1007_g N_B1_M1009_g
+ N_B1_c_129_n N_B1_c_130_n B1 B1 N_B1_c_132_n PM_SKY130_FD_SC_LP__A21O_LP%B1
x_PM_SKY130_FD_SC_LP__A21O_LP%A_218_57# N_A_218_57#_M1005_d N_A_218_57#_M1007_d
+ N_A_218_57#_c_178_n N_A_218_57#_M1002_g N_A_218_57#_c_179_n
+ N_A_218_57#_M1004_g N_A_218_57#_c_180_n N_A_218_57#_M1000_g
+ N_A_218_57#_c_182_n N_A_218_57#_c_183_n N_A_218_57#_c_184_n
+ N_A_218_57#_c_188_n N_A_218_57#_c_189_n N_A_218_57#_c_185_n
+ N_A_218_57#_c_186_n PM_SKY130_FD_SC_LP__A21O_LP%A_218_57#
x_PM_SKY130_FD_SC_LP__A21O_LP%A_33_409# N_A_33_409#_M1003_s N_A_33_409#_M1008_d
+ N_A_33_409#_c_250_n N_A_33_409#_c_251_n N_A_33_409#_c_252_n
+ N_A_33_409#_c_253_n PM_SKY130_FD_SC_LP__A21O_LP%A_33_409#
x_PM_SKY130_FD_SC_LP__A21O_LP%VPWR N_VPWR_M1003_d N_VPWR_M1000_s N_VPWR_c_281_n
+ N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n VPWR N_VPWR_c_285_n
+ N_VPWR_c_280_n N_VPWR_c_287_n PM_SKY130_FD_SC_LP__A21O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A21O_LP%X N_X_M1004_d N_X_M1000_d N_X_c_319_n X X X X
+ N_X_c_318_n PM_SKY130_FD_SC_LP__A21O_LP%X
x_PM_SKY130_FD_SC_LP__A21O_LP%VGND N_VGND_M1006_s N_VGND_M1009_d N_VGND_c_335_n
+ N_VGND_c_336_n N_VGND_c_337_n VGND N_VGND_c_338_n N_VGND_c_339_n
+ N_VGND_c_340_n N_VGND_c_341_n PM_SKY130_FD_SC_LP__A21O_LP%VGND
cc_1 VNB N_A2_M1006_g 0.0446542f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.495
cc_2 VNB N_A2_c_61_n 0.0625546f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_3 VNB N_A2_c_62_n 0.0297987f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_4 VNB N_A1_M1005_g 0.0355564f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.545
cc_5 VNB N_A1_c_89_n 0.00161387f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.11
cc_6 VNB N_A1_c_90_n 0.0218195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A1_c_91_n 0.0157887f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.78
cc_8 VNB N_A1_c_92_n 0.00912353f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.275
cc_9 VNB N_B1_M1001_g 0.0317853f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.545
cc_10 VNB N_B1_M1009_g 0.0291846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_c_129_n 0.0245519f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.78
cc_12 VNB N_B1_c_130_n 0.00192862f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_13 VNB B1 2.87194e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_132_n 0.0274124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_218_57#_c_178_n 0.0155418f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.495
cc_16 VNB N_A_218_57#_c_179_n 0.0198961f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_A_218_57#_c_180_n 0.0874408f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.275
cc_18 VNB N_A_218_57#_M1000_g 0.0143172f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_19 VNB N_A_218_57#_c_182_n 0.00353811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_218_57#_c_183_n 0.00639569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_218_57#_c_184_n 0.0114616f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_22 VNB N_A_218_57#_c_185_n 0.00364134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_218_57#_c_186_n 0.0235183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_280_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB X 0.00387738f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.11
cc_26 VNB N_X_c_318_n 0.0598407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_335_n 0.0155295f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.495
cc_28 VNB N_VGND_c_336_n 0.0249264f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_29 VNB N_VGND_c_337_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.275
cc_30 VNB N_VGND_c_338_n 0.0406624f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.78
cc_31 VNB N_VGND_c_339_n 0.0304129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_340_n 0.221236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_341_n 0.00497896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_A2_M1003_g 0.0413391f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.545
cc_35 VPB N_A2_c_61_n 0.0187581f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_36 VPB N_A2_c_62_n 0.0085757f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_37 VPB N_A1_c_89_n 0.0112934f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.11
cc_38 VPB N_A1_M1008_g 0.0307811f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.495
cc_39 VPB N_A1_c_92_n 0.00207587f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.275
cc_40 VPB N_B1_M1007_g 0.0353222f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.495
cc_41 VPB N_B1_c_130_n 0.0130549f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.295
cc_42 VPB B1 8.2657e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_218_57#_M1000_g 0.0485539f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_44 VPB N_A_218_57#_c_188_n 0.0137625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_218_57#_c_189_n 0.0109364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_218_57#_c_185_n 0.00968523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_33_409#_c_250_n 0.0372257f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_48 VPB N_A_33_409#_c_251_n 0.017172f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.275
cc_49 VPB N_A_33_409#_c_252_n 0.00954711f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_50 VPB N_A_33_409#_c_253_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.78
cc_51 VPB N_VPWR_c_281_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_282_n 0.0184261f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_53 VPB N_VPWR_c_283_n 0.0359279f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.295
cc_54 VPB N_VPWR_c_284_n 0.00598038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_285_n 0.0197141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_280_n 0.0647956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_287_n 0.0248585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_X_c_319_n 0.0496579f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_59 VPB X 0.00538525f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.11
cc_60 N_A2_M1006_g N_A1_M1005_g 0.0295506f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_61 N_A2_c_62_n N_A1_M1005_g 0.00198195f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_62 N_A2_M1003_g N_A1_M1008_g 0.0312016f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_63 N_A2_M1003_g N_A1_c_90_n 0.0295506f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_64 N_A2_c_61_n N_A1_c_91_n 0.0295506f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_65 N_A2_c_61_n N_A1_c_92_n 0.00290961f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_66 N_A2_c_62_n N_A1_c_92_n 0.0258963f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_67 N_A2_M1003_g N_A_33_409#_c_250_n 0.0165939f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_68 N_A2_M1003_g N_A_33_409#_c_251_n 0.0224516f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_69 N_A2_c_62_n N_A_33_409#_c_251_n 0.00501052f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_70 N_A2_M1003_g N_A_33_409#_c_252_n 0.00217317f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_71 N_A2_c_61_n N_A_33_409#_c_252_n 0.00177069f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_72 N_A2_c_62_n N_A_33_409#_c_252_n 0.0267187f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_73 N_A2_M1003_g N_A_33_409#_c_253_n 9.13404e-19 $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_74 N_A2_M1003_g N_VPWR_c_281_n 0.0184761f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_75 N_A2_M1003_g N_VPWR_c_280_n 0.0141028f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_76 N_A2_M1003_g N_VPWR_c_287_n 0.00769046f $X=0.575 $Y=2.545 $X2=0 $Y2=0
cc_77 N_A2_M1006_g N_VGND_c_336_n 0.0162616f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_78 N_A2_c_61_n N_VGND_c_336_n 0.00213498f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_79 N_A2_c_62_n N_VGND_c_336_n 0.0146189f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_80 N_A2_M1006_g N_VGND_c_338_n 0.00445056f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_81 N_A2_M1006_g N_VGND_c_340_n 0.00804604f $X=0.625 $Y=0.495 $X2=0 $Y2=0
cc_82 N_A1_M1005_g N_B1_M1001_g 0.0201384f $X=1.015 $Y=0.495 $X2=0 $Y2=0
cc_83 N_A1_M1008_g N_B1_M1007_g 0.0195028f $X=1.105 $Y=2.545 $X2=0 $Y2=0
cc_84 N_A1_c_91_n N_B1_c_129_n 0.0118705f $X=1.105 $Y=1.29 $X2=0 $Y2=0
cc_85 N_A1_c_92_n N_B1_c_129_n 0.00416906f $X=1.105 $Y=1.29 $X2=0 $Y2=0
cc_86 N_A1_c_89_n N_B1_c_130_n 0.0118705f $X=1.105 $Y=1.795 $X2=0 $Y2=0
cc_87 N_A1_c_91_n B1 7.81732e-19 $X=1.105 $Y=1.29 $X2=0 $Y2=0
cc_88 N_A1_c_92_n B1 0.04827f $X=1.105 $Y=1.29 $X2=0 $Y2=0
cc_89 N_A1_c_90_n N_B1_c_132_n 0.0118705f $X=1.105 $Y=1.63 $X2=0 $Y2=0
cc_90 N_A1_M1005_g N_A_218_57#_c_182_n 0.00777625f $X=1.015 $Y=0.495 $X2=0 $Y2=0
cc_91 N_A1_M1005_g N_A_218_57#_c_184_n 0.00526606f $X=1.015 $Y=0.495 $X2=0 $Y2=0
cc_92 N_A1_c_91_n N_A_218_57#_c_184_n 5.0243e-19 $X=1.105 $Y=1.29 $X2=0 $Y2=0
cc_93 N_A1_c_92_n N_A_218_57#_c_184_n 0.00949618f $X=1.105 $Y=1.29 $X2=0 $Y2=0
cc_94 N_A1_M1008_g N_A_218_57#_c_189_n 2.76446e-19 $X=1.105 $Y=2.545 $X2=0 $Y2=0
cc_95 N_A1_M1008_g N_A_33_409#_c_250_n 9.13404e-19 $X=1.105 $Y=2.545 $X2=0 $Y2=0
cc_96 N_A1_c_89_n N_A_33_409#_c_251_n 5.78893e-19 $X=1.105 $Y=1.795 $X2=0 $Y2=0
cc_97 N_A1_M1008_g N_A_33_409#_c_251_n 0.0194258f $X=1.105 $Y=2.545 $X2=0 $Y2=0
cc_98 N_A1_c_92_n N_A_33_409#_c_251_n 0.0286772f $X=1.105 $Y=1.29 $X2=0 $Y2=0
cc_99 N_A1_M1008_g N_A_33_409#_c_253_n 0.0164338f $X=1.105 $Y=2.545 $X2=0 $Y2=0
cc_100 N_A1_M1008_g N_VPWR_c_281_n 0.0174292f $X=1.105 $Y=2.545 $X2=0 $Y2=0
cc_101 N_A1_M1008_g N_VPWR_c_283_n 0.00769046f $X=1.105 $Y=2.545 $X2=0 $Y2=0
cc_102 N_A1_M1008_g N_VPWR_c_280_n 0.0134474f $X=1.105 $Y=2.545 $X2=0 $Y2=0
cc_103 N_A1_M1005_g N_VGND_c_336_n 0.00221874f $X=1.015 $Y=0.495 $X2=0 $Y2=0
cc_104 N_A1_M1005_g N_VGND_c_338_n 0.0053602f $X=1.015 $Y=0.495 $X2=0 $Y2=0
cc_105 N_A1_M1005_g N_VGND_c_340_n 0.0106011f $X=1.015 $Y=0.495 $X2=0 $Y2=0
cc_106 N_B1_M1009_g N_A_218_57#_c_178_n 0.0174634f $X=1.945 $Y=0.495 $X2=0 $Y2=0
cc_107 N_B1_c_129_n N_A_218_57#_c_180_n 0.0174634f $X=1.945 $Y=1.2 $X2=0 $Y2=0
cc_108 B1 N_A_218_57#_c_180_n 2.73877e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B1_c_132_n N_A_218_57#_c_180_n 0.00439647f $X=1.675 $Y=1.29 $X2=0 $Y2=0
cc_110 N_B1_M1001_g N_A_218_57#_c_182_n 0.0101326f $X=1.585 $Y=0.495 $X2=0 $Y2=0
cc_111 N_B1_M1009_g N_A_218_57#_c_182_n 0.00179788f $X=1.945 $Y=0.495 $X2=0
+ $Y2=0
cc_112 N_B1_M1001_g N_A_218_57#_c_183_n 0.00795118f $X=1.585 $Y=0.495 $X2=0
+ $Y2=0
cc_113 N_B1_M1009_g N_A_218_57#_c_183_n 0.0130223f $X=1.945 $Y=0.495 $X2=0 $Y2=0
cc_114 N_B1_c_129_n N_A_218_57#_c_183_n 2.06304e-19 $X=1.945 $Y=1.2 $X2=0 $Y2=0
cc_115 B1 N_A_218_57#_c_183_n 0.0227314f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_116 N_B1_M1001_g N_A_218_57#_c_184_n 0.00300966f $X=1.585 $Y=0.495 $X2=0
+ $Y2=0
cc_117 B1 N_A_218_57#_c_184_n 0.00193735f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B1_M1007_g N_A_218_57#_c_188_n 0.0143689f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_119 N_B1_M1007_g N_A_218_57#_c_189_n 0.00466771f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_120 N_B1_c_130_n N_A_218_57#_c_189_n 5.96441e-19 $X=1.675 $Y=1.795 $X2=0
+ $Y2=0
cc_121 B1 N_A_218_57#_c_189_n 0.00719112f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B1_M1007_g N_A_218_57#_c_185_n 0.00701028f $X=1.635 $Y=2.545 $X2=0
+ $Y2=0
cc_123 N_B1_c_130_n N_A_218_57#_c_185_n 0.00439059f $X=1.675 $Y=1.795 $X2=0
+ $Y2=0
cc_124 N_B1_M1009_g N_A_218_57#_c_186_n 0.00964151f $X=1.945 $Y=0.495 $X2=0
+ $Y2=0
cc_125 B1 N_A_218_57#_c_186_n 0.0508983f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B1_c_132_n N_A_218_57#_c_186_n 0.00439059f $X=1.675 $Y=1.29 $X2=0 $Y2=0
cc_127 N_B1_M1007_g N_A_33_409#_c_251_n 0.0043772f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_128 B1 N_A_33_409#_c_251_n 0.00193735f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B1_M1007_g N_A_33_409#_c_253_n 0.0164995f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_130 N_B1_M1007_g N_VPWR_c_281_n 8.61967e-19 $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_131 N_B1_M1007_g N_VPWR_c_282_n 0.00307416f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_132 N_B1_M1007_g N_VPWR_c_283_n 0.00826654f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_133 N_B1_M1007_g N_VPWR_c_280_n 0.0158042f $X=1.635 $Y=2.545 $X2=0 $Y2=0
cc_134 N_B1_M1001_g N_VGND_c_337_n 0.00175817f $X=1.585 $Y=0.495 $X2=0 $Y2=0
cc_135 N_B1_M1009_g N_VGND_c_337_n 0.00984956f $X=1.945 $Y=0.495 $X2=0 $Y2=0
cc_136 N_B1_M1001_g N_VGND_c_338_n 0.00502664f $X=1.585 $Y=0.495 $X2=0 $Y2=0
cc_137 N_B1_M1009_g N_VGND_c_338_n 0.00445056f $X=1.945 $Y=0.495 $X2=0 $Y2=0
cc_138 N_B1_M1001_g N_VGND_c_340_n 0.00574098f $X=1.585 $Y=0.495 $X2=0 $Y2=0
cc_139 N_B1_M1009_g N_VGND_c_340_n 0.00409056f $X=1.945 $Y=0.495 $X2=0 $Y2=0
cc_140 N_A_218_57#_c_189_n N_A_33_409#_c_251_n 0.00860423f $X=1.9 $Y=2.19 $X2=0
+ $Y2=0
cc_141 N_A_218_57#_c_185_n N_A_33_409#_c_251_n 0.00178561f $X=1.962 $Y=2.025
+ $X2=0 $Y2=0
cc_142 N_A_218_57#_c_189_n N_A_33_409#_c_253_n 0.0620783f $X=1.9 $Y=2.19 $X2=0
+ $Y2=0
cc_143 N_A_218_57#_c_180_n N_VPWR_c_282_n 0.00377837f $X=2.815 $Y=1.485 $X2=0
+ $Y2=0
cc_144 N_A_218_57#_M1000_g N_VPWR_c_282_n 0.0272973f $X=2.815 $Y=2.48 $X2=0
+ $Y2=0
cc_145 N_A_218_57#_c_185_n N_VPWR_c_282_n 0.0852029f $X=1.962 $Y=2.025 $X2=0
+ $Y2=0
cc_146 N_A_218_57#_c_186_n N_VPWR_c_282_n 0.0100249f $X=2.325 $Y=0.86 $X2=0
+ $Y2=0
cc_147 N_A_218_57#_c_188_n N_VPWR_c_283_n 0.0304602f $X=1.9 $Y=2.9 $X2=0 $Y2=0
cc_148 N_A_218_57#_M1000_g N_VPWR_c_285_n 0.00687065f $X=2.815 $Y=2.48 $X2=0
+ $Y2=0
cc_149 N_A_218_57#_M1000_g N_VPWR_c_280_n 0.013111f $X=2.815 $Y=2.48 $X2=0 $Y2=0
cc_150 N_A_218_57#_c_188_n N_VPWR_c_280_n 0.0174175f $X=1.9 $Y=2.9 $X2=0 $Y2=0
cc_151 N_A_218_57#_M1000_g N_X_c_319_n 0.0308063f $X=2.815 $Y=2.48 $X2=0 $Y2=0
cc_152 N_A_218_57#_M1000_g X 0.0161393f $X=2.815 $Y=2.48 $X2=0 $Y2=0
cc_153 N_A_218_57#_c_178_n N_X_c_318_n 0.00185142f $X=2.375 $Y=0.815 $X2=0 $Y2=0
cc_154 N_A_218_57#_c_179_n N_X_c_318_n 0.0127775f $X=2.765 $Y=0.815 $X2=0 $Y2=0
cc_155 N_A_218_57#_c_180_n N_X_c_318_n 0.031339f $X=2.815 $Y=1.485 $X2=0 $Y2=0
cc_156 N_A_218_57#_M1000_g N_X_c_318_n 0.00399057f $X=2.815 $Y=2.48 $X2=0 $Y2=0
cc_157 N_A_218_57#_c_185_n N_X_c_318_n 0.00834543f $X=1.962 $Y=2.025 $X2=0 $Y2=0
cc_158 N_A_218_57#_c_186_n N_X_c_318_n 0.0534137f $X=2.325 $Y=0.86 $X2=0 $Y2=0
cc_159 N_A_218_57#_c_182_n N_VGND_c_336_n 0.0127119f $X=1.37 $Y=0.495 $X2=0
+ $Y2=0
cc_160 N_A_218_57#_c_178_n N_VGND_c_337_n 0.0100745f $X=2.375 $Y=0.815 $X2=0
+ $Y2=0
cc_161 N_A_218_57#_c_179_n N_VGND_c_337_n 0.00176437f $X=2.765 $Y=0.815 $X2=0
+ $Y2=0
cc_162 N_A_218_57#_c_182_n N_VGND_c_337_n 0.0110409f $X=1.37 $Y=0.495 $X2=0
+ $Y2=0
cc_163 N_A_218_57#_c_183_n N_VGND_c_337_n 0.00164881f $X=2.02 $Y=0.86 $X2=0
+ $Y2=0
cc_164 N_A_218_57#_c_186_n N_VGND_c_337_n 0.0206789f $X=2.325 $Y=0.86 $X2=0
+ $Y2=0
cc_165 N_A_218_57#_c_182_n N_VGND_c_338_n 0.0220321f $X=1.37 $Y=0.495 $X2=0
+ $Y2=0
cc_166 N_A_218_57#_c_178_n N_VGND_c_339_n 0.00445056f $X=2.375 $Y=0.815 $X2=0
+ $Y2=0
cc_167 N_A_218_57#_c_179_n N_VGND_c_339_n 0.00502664f $X=2.765 $Y=0.815 $X2=0
+ $Y2=0
cc_168 N_A_218_57#_c_178_n N_VGND_c_340_n 0.00414878f $X=2.375 $Y=0.815 $X2=0
+ $Y2=0
cc_169 N_A_218_57#_c_179_n N_VGND_c_340_n 0.0101752f $X=2.765 $Y=0.815 $X2=0
+ $Y2=0
cc_170 N_A_218_57#_c_182_n N_VGND_c_340_n 0.0125808f $X=1.37 $Y=0.495 $X2=0
+ $Y2=0
cc_171 N_A_218_57#_c_183_n N_VGND_c_340_n 0.0151124f $X=2.02 $Y=0.86 $X2=0 $Y2=0
cc_172 N_A_218_57#_c_186_n N_VGND_c_340_n 0.0130537f $X=2.325 $Y=0.86 $X2=0
+ $Y2=0
cc_173 N_A_33_409#_c_251_n N_VPWR_M1003_d 0.00180746f $X=1.205 $Y=2.06 $X2=-0.19
+ $Y2=1.655
cc_174 N_A_33_409#_c_250_n N_VPWR_c_281_n 0.0487591f $X=0.31 $Y=2.19 $X2=0 $Y2=0
cc_175 N_A_33_409#_c_251_n N_VPWR_c_281_n 0.0163515f $X=1.205 $Y=2.06 $X2=0
+ $Y2=0
cc_176 N_A_33_409#_c_253_n N_VPWR_c_281_n 0.0487591f $X=1.37 $Y=2.19 $X2=0 $Y2=0
cc_177 N_A_33_409#_c_253_n N_VPWR_c_283_n 0.021949f $X=1.37 $Y=2.19 $X2=0 $Y2=0
cc_178 N_A_33_409#_c_250_n N_VPWR_c_280_n 0.0125808f $X=0.31 $Y=2.19 $X2=0 $Y2=0
cc_179 N_A_33_409#_c_253_n N_VPWR_c_280_n 0.0124703f $X=1.37 $Y=2.19 $X2=0 $Y2=0
cc_180 N_A_33_409#_c_250_n N_VPWR_c_287_n 0.0220321f $X=0.31 $Y=2.19 $X2=0 $Y2=0
cc_181 N_VPWR_c_282_n N_X_c_319_n 0.0685263f $X=2.55 $Y=2.125 $X2=0 $Y2=0
cc_182 N_VPWR_c_285_n N_X_c_319_n 0.0158357f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_280_n N_X_c_319_n 0.0121432f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_184 N_X_c_318_n N_VGND_c_337_n 0.0106706f $X=2.98 $Y=0.495 $X2=0 $Y2=0
cc_185 N_X_c_318_n N_VGND_c_339_n 0.0287746f $X=2.98 $Y=0.495 $X2=0 $Y2=0
cc_186 N_X_c_318_n N_VGND_c_340_n 0.0164501f $X=2.98 $Y=0.495 $X2=0 $Y2=0
