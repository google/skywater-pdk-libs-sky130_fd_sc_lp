# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand3b_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nand3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.345000 0.830000 1.750000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 1.345000 1.720000 1.735000 ;
        RECT 1.530000 1.735000 3.330000 1.905000 ;
        RECT 2.520000 1.345000 3.330000 1.735000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 1.345000 1.360000 1.750000 ;
        RECT 1.190000 1.750000 1.360000 2.075000 ;
        RECT 1.190000 2.075000 3.790000 2.245000 ;
        RECT 3.540000 1.345000 3.790000 2.075000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.453200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.225000 2.415000 4.235000 2.585000 ;
        RECT 1.225000 2.585000 1.555000 3.075000 ;
        RECT 2.240000 0.935000 2.570000 1.005000 ;
        RECT 2.240000 1.005000 4.235000 1.175000 ;
        RECT 2.245000 2.585000 2.575000 3.075000 ;
        RECT 3.235000 2.585000 3.565000 3.075000 ;
        RECT 3.960000 1.175000 4.235000 2.415000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
        RECT 0.775000  0.085000 1.105000 0.835000 ;
        RECT 3.665000  0.085000 3.995000 0.835000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.320000 3.415000 ;
        RECT 0.735000 1.920000 1.020000 3.245000 ;
        RECT 1.735000 2.755000 2.065000 3.245000 ;
        RECT 2.745000 2.755000 3.065000 3.245000 ;
        RECT 3.735000 2.755000 3.995000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.825000 0.565000 1.005000 ;
      RECT 0.090000 1.005000 2.060000 1.175000 ;
      RECT 0.090000 1.175000 0.260000 1.920000 ;
      RECT 0.090000 1.920000 0.565000 2.200000 ;
      RECT 1.275000 0.255000 3.495000 0.425000 ;
      RECT 1.275000 0.425000 1.535000 0.835000 ;
      RECT 1.705000 0.595000 3.095000 0.765000 ;
      RECT 1.705000 0.765000 2.035000 0.835000 ;
      RECT 1.890000 1.175000 2.060000 1.345000 ;
      RECT 1.890000 1.345000 2.350000 1.565000 ;
      RECT 2.765000 0.765000 3.095000 0.835000 ;
      RECT 3.265000 0.425000 3.495000 0.835000 ;
  END
END sky130_fd_sc_lp__nand3b_2
