* File: sky130_fd_sc_lp__mux2i_m.spice
* Created: Fri Aug 28 10:45:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2i_m.pex.spice"
.subckt sky130_fd_sc_lp__mux2i_m  VNB VPB S A1 A0 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_S_M1004_g N_A_55_125#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=17.136 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1008 A_250_125# N_A_55_125#_M1008_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_A0_M1007_g A_250_125# VNB NSHORT L=0.15 W=0.42 AD=0.0672
+ AS=0.0441 PD=0.74 PS=0.63 NRD=11.424 NRS=14.28 M=1 R=2.8 SA=75001.1 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1009 A_416_125# N_A1_M1009_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.42 AD=0.08295
+ AS=0.0672 PD=0.815 PS=0.74 NRD=40.704 NRS=0 M=1 R=2.8 SA=75001.6 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_S_M1000_g A_416_125# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.08295 PD=1.37 PS=0.815 NRD=0 NRS=40.704 M=1 R=2.8 SA=75002.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_S_M1005_g N_A_55_125#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0756 AS=0.1113 PD=0.78 PS=1.37 NRD=37.5088 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1006 A_256_497# N_A_55_125#_M1006_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0756 PD=0.63 PS=0.78 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A1_M1001_g A_256_497# VPB PHIGHVT L=0.15 W=0.42 AD=0.0987
+ AS=0.0441 PD=0.89 PS=0.63 NRD=44.5417 NRS=23.443 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 A_452_497# N_A0_M1002_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0651
+ AS=0.0987 PD=0.73 PS=0.89 NRD=46.886 NRS=44.5417 M=1 R=2.8 SA=75001.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_S_M1003_g A_452_497# VPB PHIGHVT L=0.15 W=0.42 AD=0.1512
+ AS=0.0651 PD=1.56 PS=0.73 NRD=44.5417 NRS=46.886 M=1 R=2.8 SA=75002.1
+ SB=75000.3 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_74 VPB 0 2.58154e-19 $X=0 $Y=3.085
c_474 A_452_497# 0 1.6591e-19 $X=2.26 $Y=2.485
*
.include "sky130_fd_sc_lp__mux2i_m.pxi.spice"
*
.ends
*
*
