* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_286_492# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_80_21# B2 a_592_492# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_237_131# A2_N a_286_492# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND A1_N a_237_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_80_21# a_286_492# a_506_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_592_492# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_506_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR A1_N a_286_492# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR a_286_492# a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND B1 a_506_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
