* File: sky130_fd_sc_lp__nor4bb_2.pxi.spice
* Created: Fri Aug 28 10:59:02 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4BB_2%C_N N_C_N_M1006_g N_C_N_c_119_n N_C_N_M1014_g
+ N_C_N_c_121_n C_N C_N N_C_N_c_118_n PM_SKY130_FD_SC_LP__NOR4BB_2%C_N
x_PM_SKY130_FD_SC_LP__NOR4BB_2%D_N N_D_N_M1011_g N_D_N_M1007_g N_D_N_c_153_n
+ N_D_N_c_154_n D_N D_N D_N N_D_N_c_151_n PM_SKY130_FD_SC_LP__NOR4BB_2%D_N
x_PM_SKY130_FD_SC_LP__NOR4BB_2%A_286_512# N_A_286_512#_M1007_d
+ N_A_286_512#_M1011_d N_A_286_512#_c_187_n N_A_286_512#_c_188_n
+ N_A_286_512#_M1012_g N_A_286_512#_M1005_g N_A_286_512#_c_190_n
+ N_A_286_512#_c_191_n N_A_286_512#_M1015_g N_A_286_512#_M1016_g
+ N_A_286_512#_c_193_n N_A_286_512#_c_194_n N_A_286_512#_c_195_n
+ N_A_286_512#_c_196_n N_A_286_512#_c_202_n N_A_286_512#_c_197_n
+ N_A_286_512#_c_198_n PM_SKY130_FD_SC_LP__NOR4BB_2%A_286_512#
x_PM_SKY130_FD_SC_LP__NOR4BB_2%A_45_164# N_A_45_164#_M1006_s N_A_45_164#_M1014_s
+ N_A_45_164#_M1000_g N_A_45_164#_M1001_g N_A_45_164#_M1010_g
+ N_A_45_164#_M1017_g N_A_45_164#_c_268_n N_A_45_164#_c_269_n
+ N_A_45_164#_c_285_n N_A_45_164#_c_270_n N_A_45_164#_c_271_n
+ N_A_45_164#_c_272_n N_A_45_164#_c_273_n N_A_45_164#_c_274_n
+ N_A_45_164#_c_275_n N_A_45_164#_c_280_n N_A_45_164#_c_276_n
+ N_A_45_164#_c_277_n PM_SKY130_FD_SC_LP__NOR4BB_2%A_45_164#
x_PM_SKY130_FD_SC_LP__NOR4BB_2%B N_B_c_375_n N_B_M1002_g N_B_c_379_n N_B_M1009_g
+ N_B_c_376_n N_B_M1008_g N_B_c_380_n N_B_M1019_g B N_B_c_378_n
+ PM_SKY130_FD_SC_LP__NOR4BB_2%B
x_PM_SKY130_FD_SC_LP__NOR4BB_2%A N_A_c_427_n N_A_M1004_g N_A_M1003_g N_A_c_429_n
+ N_A_M1018_g N_A_M1013_g A N_A_c_432_n PM_SKY130_FD_SC_LP__NOR4BB_2%A
x_PM_SKY130_FD_SC_LP__NOR4BB_2%VPWR N_VPWR_M1014_d N_VPWR_M1003_s N_VPWR_c_464_n
+ VPWR N_VPWR_c_465_n N_VPWR_c_466_n N_VPWR_c_467_n N_VPWR_c_463_n
+ N_VPWR_c_469_n N_VPWR_c_470_n PM_SKY130_FD_SC_LP__NOR4BB_2%VPWR
x_PM_SKY130_FD_SC_LP__NOR4BB_2%A_463_355# N_A_463_355#_M1005_s
+ N_A_463_355#_M1016_s N_A_463_355#_M1017_s N_A_463_355#_c_526_n
+ N_A_463_355#_c_527_n N_A_463_355#_c_528_n N_A_463_355#_c_549_p
+ N_A_463_355#_c_539_n N_A_463_355#_c_529_n
+ PM_SKY130_FD_SC_LP__NOR4BB_2%A_463_355#
x_PM_SKY130_FD_SC_LP__NOR4BB_2%Y N_Y_M1012_d N_Y_M1000_d N_Y_M1002_d N_Y_M1004_s
+ N_Y_M1005_d N_Y_c_570_n N_Y_c_640_p N_Y_c_560_n N_Y_c_643_p N_Y_c_598_n
+ N_Y_c_641_p N_Y_c_561_n N_Y_c_642_p N_Y_c_566_n N_Y_c_562_n Y Y Y N_Y_c_569_n
+ Y N_Y_c_564_n N_Y_c_565_n PM_SKY130_FD_SC_LP__NOR4BB_2%Y
x_PM_SKY130_FD_SC_LP__NOR4BB_2%A_718_355# N_A_718_355#_M1001_d
+ N_A_718_355#_M1009_d N_A_718_355#_c_658_n N_A_718_355#_c_656_n
+ N_A_718_355#_c_657_n N_A_718_355#_c_664_n N_A_718_355#_c_666_n
+ PM_SKY130_FD_SC_LP__NOR4BB_2%A_718_355#
x_PM_SKY130_FD_SC_LP__NOR4BB_2%A_919_367# N_A_919_367#_M1009_s
+ N_A_919_367#_M1019_s N_A_919_367#_M1013_d N_A_919_367#_c_685_n
+ N_A_919_367#_c_686_n N_A_919_367#_c_687_n N_A_919_367#_c_706_n
+ N_A_919_367#_c_688_n N_A_919_367#_c_689_n N_A_919_367#_c_690_n
+ PM_SKY130_FD_SC_LP__NOR4BB_2%A_919_367#
x_PM_SKY130_FD_SC_LP__NOR4BB_2%VGND N_VGND_M1006_d N_VGND_M1012_s N_VGND_M1015_s
+ N_VGND_M1010_s N_VGND_M1008_s N_VGND_M1018_d N_VGND_c_724_n N_VGND_c_725_n
+ N_VGND_c_726_n N_VGND_c_727_n N_VGND_c_728_n N_VGND_c_729_n N_VGND_c_730_n
+ N_VGND_c_731_n N_VGND_c_732_n N_VGND_c_733_n VGND N_VGND_c_734_n
+ N_VGND_c_735_n N_VGND_c_736_n N_VGND_c_737_n N_VGND_c_738_n N_VGND_c_739_n
+ N_VGND_c_740_n N_VGND_c_741_n PM_SKY130_FD_SC_LP__NOR4BB_2%VGND
cc_1 VNB N_C_N_M1006_g 0.0396254f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.03
cc_2 VNB C_N 0.0022907f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_C_N_c_118_n 0.0133419f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.745
cc_4 VNB N_D_N_M1007_g 0.0363319f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.25
cc_5 VNB D_N 0.00493775f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_6 VNB N_D_N_c_151_n 0.0106925f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.665
cc_7 VNB N_A_286_512#_c_187_n 0.0165744f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.25
cc_8 VNB N_A_286_512#_c_188_n 0.0182959f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.77
cc_9 VNB N_A_286_512#_M1005_g 0.0126761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_286_512#_c_190_n 0.00865608f $X=-0.19 $Y=-0.245 $X2=0.687
+ $Y2=1.745
cc_11 VNB N_A_286_512#_c_191_n 0.0152683f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.745
cc_12 VNB N_A_286_512#_M1016_g 0.0111757f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.035
cc_13 VNB N_A_286_512#_c_193_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_286_512#_c_194_n 0.00515988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_286_512#_c_195_n 0.0119041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_286_512#_c_196_n 0.00122342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_286_512#_c_197_n 0.011277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_286_512#_c_198_n 0.061513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_45_164#_M1000_g 0.0189243f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.77
cc_20 VNB N_A_45_164#_M1001_g 4.86587e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_21 VNB N_A_45_164#_M1010_g 0.0224043f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.745
cc_22 VNB N_A_45_164#_M1017_g 5.2124e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_45_164#_c_268_n 0.0148251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_45_164#_c_269_n 0.025846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_45_164#_c_270_n 0.0232689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_45_164#_c_271_n 0.0038146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_45_164#_c_272_n 0.00140509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_45_164#_c_273_n 0.00353453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_45_164#_c_274_n 0.011434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_45_164#_c_275_n 0.00770964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_45_164#_c_276_n 0.0122378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_45_164#_c_277_n 0.044789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B_c_375_n 0.0187913f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.58
cc_34 VNB N_B_c_376_n 0.0150696f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.25
cc_35 VNB B 0.00474685f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_36 VNB N_B_c_378_n 0.0919711f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.665
cc_37 VNB N_A_c_427_n 0.0150696f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.58
cc_38 VNB N_A_M1003_g 0.0073278f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=2.053
cc_39 VNB N_A_c_429_n 0.0211802f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.77
cc_40 VNB N_A_M1013_g 0.0111859f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_41 VNB A 0.0194913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_c_432_n 0.0617508f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=1.665
cc_43 VNB N_VPWR_c_463_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_560_n 0.00216928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_561_n 0.00423232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_562_n 2.0355e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB Y 0.00389014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_Y_c_564_n 0.00314596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_Y_c_565_n 0.00354532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_724_n 0.0442689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_725_n 0.0127197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_726_n 3.08929e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_727_n 3.08929e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_728_n 0.0135555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_729_n 0.0330598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_730_n 0.0370827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_731_n 0.00510277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_732_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_733_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_734_n 0.0217138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_735_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_736_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_737_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_738_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_739_n 0.0156681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_740_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_741_n 0.363938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VPB N_C_N_c_119_n 0.0232987f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=2.053
cc_69 VPB N_C_N_M1014_g 0.0362436f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.77
cc_70 VPB N_C_N_c_121_n 0.0242504f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=2.25
cc_71 VPB C_N 0.00306065f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_72 VPB N_C_N_c_118_n 0.0103739f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.745
cc_73 VPB N_D_N_M1011_g 0.0354992f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.03
cc_74 VPB N_D_N_c_153_n 0.0253637f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=2.25
cc_75 VPB N_D_N_c_154_n 0.0187906f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_76 VPB D_N 0.0085266f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_77 VPB N_D_N_c_151_n 0.00675366f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.665
cc_78 VPB N_A_286_512#_M1005_g 0.0240353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_286_512#_M1016_g 0.0191767f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=2.035
cc_80 VPB N_A_286_512#_c_196_n 0.0250701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_286_512#_c_202_n 0.0115146f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_286_512#_c_197_n 0.0027677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A_286_512#_c_198_n 0.00211245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_45_164#_M1001_g 0.0198827f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_85 VPB N_A_45_164#_M1017_g 0.023651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_45_164#_c_280_n 0.0133196f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_45_164#_c_276_n 0.0487329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_B_c_379_n 0.0195571f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_B_c_380_n 0.0153124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_B_c_378_n 0.0142161f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.665
cc_91 VPB N_A_M1003_g 0.0184452f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=2.053
cc_92 VPB N_A_M1013_g 0.0241666f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_93 VPB N_VPWR_c_464_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.77
cc_94 VPB N_VPWR_c_465_n 0.0201014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_466_n 0.109489f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=1.665
cc_96 VPB N_VPWR_c_467_n 0.0160123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_463_n 0.0856684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_469_n 0.0182392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_470_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_463_355#_c_526_n 0.0183994f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_101 VPB N_A_463_355#_c_527_n 0.00447377f $X=-0.19 $Y=1.655 $X2=0.687
+ $Y2=1.745
cc_102 VPB N_A_463_355#_c_528_n 0.00646416f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.745
cc_103 VPB N_A_463_355#_c_529_n 0.00835169f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_Y_c_566_n 0.00236237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB Y 0.00102628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB Y 0.00511172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_Y_c_569_n 0.00100022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_718_355#_c_656_n 0.0129206f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=2.25
cc_109 VPB N_A_718_355#_c_657_n 0.00233177f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_110 VPB N_A_919_367#_c_685_n 0.00901164f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_111 VPB N_A_919_367#_c_686_n 0.00258254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_919_367#_c_687_n 0.00251156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_919_367#_c_688_n 0.0155021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_919_367#_c_689_n 0.0461643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_919_367#_c_690_n 0.00253228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 N_C_N_M1014_g N_D_N_M1011_g 0.00696352f $X=0.585 $Y=2.77 $X2=0 $Y2=0
cc_117 N_C_N_M1006_g N_D_N_M1007_g 0.0084128f $X=0.565 $Y=1.03 $X2=0 $Y2=0
cc_118 N_C_N_c_119_n N_D_N_c_153_n 0.00948435f $X=0.687 $Y=2.053 $X2=0 $Y2=0
cc_119 N_C_N_c_121_n N_D_N_c_154_n 0.00948435f $X=0.687 $Y=2.25 $X2=0 $Y2=0
cc_120 N_C_N_M1014_g D_N 0.00243758f $X=0.585 $Y=2.77 $X2=0 $Y2=0
cc_121 C_N D_N 0.0527537f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_122 N_C_N_c_118_n D_N 0.00457903f $X=0.72 $Y=1.745 $X2=0 $Y2=0
cc_123 C_N N_D_N_c_151_n 6.98618e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_124 N_C_N_c_118_n N_D_N_c_151_n 0.00948435f $X=0.72 $Y=1.745 $X2=0 $Y2=0
cc_125 N_C_N_M1006_g N_A_45_164#_c_269_n 0.02044f $X=0.565 $Y=1.03 $X2=0 $Y2=0
cc_126 C_N N_A_45_164#_c_269_n 0.0220631f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_127 N_C_N_c_118_n N_A_45_164#_c_269_n 0.00169903f $X=0.72 $Y=1.745 $X2=0
+ $Y2=0
cc_128 N_C_N_M1006_g N_A_45_164#_c_285_n 0.00246364f $X=0.565 $Y=1.03 $X2=0
+ $Y2=0
cc_129 N_C_N_M1006_g N_A_45_164#_c_271_n 3.45997e-19 $X=0.565 $Y=1.03 $X2=0
+ $Y2=0
cc_130 N_C_N_M1006_g N_A_45_164#_c_276_n 0.0248607f $X=0.565 $Y=1.03 $X2=0 $Y2=0
cc_131 N_C_N_M1014_g N_A_45_164#_c_276_n 0.0104469f $X=0.585 $Y=2.77 $X2=0 $Y2=0
cc_132 C_N N_A_45_164#_c_276_n 0.0511703f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_133 N_C_N_M1014_g N_VPWR_c_465_n 0.00398346f $X=0.585 $Y=2.77 $X2=0 $Y2=0
cc_134 N_C_N_M1014_g N_VPWR_c_463_n 0.00790879f $X=0.585 $Y=2.77 $X2=0 $Y2=0
cc_135 N_C_N_M1014_g N_VPWR_c_469_n 0.0139715f $X=0.585 $Y=2.77 $X2=0 $Y2=0
cc_136 N_C_N_c_121_n N_VPWR_c_469_n 0.00130531f $X=0.687 $Y=2.25 $X2=0 $Y2=0
cc_137 C_N N_VPWR_c_469_n 0.00933005f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_138 N_C_N_M1006_g N_VGND_c_724_n 0.0130153f $X=0.565 $Y=1.03 $X2=0 $Y2=0
cc_139 N_C_N_M1006_g N_VGND_c_734_n 0.00270981f $X=0.565 $Y=1.03 $X2=0 $Y2=0
cc_140 N_C_N_M1006_g N_VGND_c_741_n 0.00351741f $X=0.565 $Y=1.03 $X2=0 $Y2=0
cc_141 N_D_N_M1007_g N_A_286_512#_c_195_n 0.00454874f $X=1.425 $Y=1.03 $X2=0
+ $Y2=0
cc_142 N_D_N_M1011_g N_A_286_512#_c_196_n 0.00844048f $X=1.355 $Y=2.77 $X2=0
+ $Y2=0
cc_143 N_D_N_c_153_n N_A_286_512#_c_196_n 0.00940801f $X=1.335 $Y=2.085 $X2=0
+ $Y2=0
cc_144 N_D_N_M1011_g N_A_286_512#_c_202_n 4.3369e-19 $X=1.355 $Y=2.77 $X2=0
+ $Y2=0
cc_145 N_D_N_c_154_n N_A_286_512#_c_202_n 6.65526e-19 $X=1.335 $Y=2.25 $X2=0
+ $Y2=0
cc_146 N_D_N_M1007_g N_A_286_512#_c_197_n 0.0094262f $X=1.425 $Y=1.03 $X2=0
+ $Y2=0
cc_147 D_N N_A_286_512#_c_197_n 0.0378031f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_148 N_D_N_M1007_g N_A_286_512#_c_198_n 0.0150469f $X=1.425 $Y=1.03 $X2=0
+ $Y2=0
cc_149 N_D_N_M1007_g N_A_45_164#_c_269_n 0.00310555f $X=1.425 $Y=1.03 $X2=0
+ $Y2=0
cc_150 D_N N_A_45_164#_c_269_n 0.0211507f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_151 N_D_N_c_151_n N_A_45_164#_c_269_n 9.78483e-19 $X=1.335 $Y=1.745 $X2=0
+ $Y2=0
cc_152 N_D_N_M1007_g N_A_45_164#_c_270_n 0.0155411f $X=1.425 $Y=1.03 $X2=0 $Y2=0
cc_153 D_N N_A_45_164#_c_276_n 0.00825978f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_154 N_D_N_M1011_g N_VPWR_c_466_n 0.00398346f $X=1.355 $Y=2.77 $X2=0 $Y2=0
cc_155 N_D_N_M1011_g N_VPWR_c_463_n 0.00453171f $X=1.355 $Y=2.77 $X2=0 $Y2=0
cc_156 D_N N_VPWR_c_463_n 0.00459418f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_157 N_D_N_M1011_g N_VPWR_c_469_n 0.0114177f $X=1.355 $Y=2.77 $X2=0 $Y2=0
cc_158 N_D_N_c_154_n N_VPWR_c_469_n 3.85962e-19 $X=1.335 $Y=2.25 $X2=0 $Y2=0
cc_159 D_N N_VPWR_c_469_n 0.0194355f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_160 N_D_N_M1007_g N_VGND_c_724_n 7.86974e-19 $X=1.425 $Y=1.03 $X2=0 $Y2=0
cc_161 N_D_N_M1007_g N_VGND_c_730_n 5.40682e-19 $X=1.425 $Y=1.03 $X2=0 $Y2=0
cc_162 N_A_286_512#_c_191_n N_A_45_164#_M1000_g 0.0210178f $X=3.085 $Y=1.185
+ $X2=0 $Y2=0
cc_163 N_A_286_512#_M1016_g N_A_45_164#_M1001_g 0.0247311f $X=3.085 $Y=2.405
+ $X2=0 $Y2=0
cc_164 N_A_286_512#_c_195_n N_A_45_164#_c_269_n 0.00149669f $X=1.805 $Y=1.13
+ $X2=0 $Y2=0
cc_165 N_A_286_512#_c_197_n N_A_45_164#_c_269_n 0.00626643f $X=2.04 $Y=1.095
+ $X2=0 $Y2=0
cc_166 N_A_286_512#_M1007_d N_A_45_164#_c_270_n 0.00221647f $X=1.5 $Y=0.82 $X2=0
+ $Y2=0
cc_167 N_A_286_512#_c_187_n N_A_45_164#_c_270_n 0.00251691f $X=2.58 $Y=1.26
+ $X2=0 $Y2=0
cc_168 N_A_286_512#_c_195_n N_A_45_164#_c_270_n 0.0204318f $X=1.805 $Y=1.13
+ $X2=0 $Y2=0
cc_169 N_A_286_512#_c_197_n N_A_45_164#_c_270_n 0.0319359f $X=2.04 $Y=1.095
+ $X2=0 $Y2=0
cc_170 N_A_286_512#_c_198_n N_A_45_164#_c_270_n 0.00931138f $X=2.04 $Y=1.095
+ $X2=0 $Y2=0
cc_171 N_A_286_512#_c_187_n N_A_45_164#_c_272_n 0.0131537f $X=2.58 $Y=1.26 $X2=0
+ $Y2=0
cc_172 N_A_286_512#_c_188_n N_A_45_164#_c_272_n 0.00418027f $X=2.655 $Y=1.185
+ $X2=0 $Y2=0
cc_173 N_A_286_512#_c_197_n N_A_45_164#_c_272_n 0.0237754f $X=2.04 $Y=1.095
+ $X2=0 $Y2=0
cc_174 N_A_286_512#_c_198_n N_A_45_164#_c_272_n 0.00291253f $X=2.04 $Y=1.095
+ $X2=0 $Y2=0
cc_175 N_A_286_512#_c_187_n N_A_45_164#_c_273_n 0.00184943f $X=2.58 $Y=1.26
+ $X2=0 $Y2=0
cc_176 N_A_286_512#_c_197_n N_A_45_164#_c_273_n 0.0139155f $X=2.04 $Y=1.095
+ $X2=0 $Y2=0
cc_177 N_A_286_512#_c_198_n N_A_45_164#_c_273_n 0.00139869f $X=2.04 $Y=1.095
+ $X2=0 $Y2=0
cc_178 N_A_286_512#_M1005_g N_A_45_164#_c_274_n 0.0186434f $X=2.655 $Y=2.405
+ $X2=0 $Y2=0
cc_179 N_A_286_512#_c_190_n N_A_45_164#_c_274_n 0.00234667f $X=3.01 $Y=1.26
+ $X2=0 $Y2=0
cc_180 N_A_286_512#_M1016_g N_A_45_164#_c_274_n 0.00994322f $X=3.085 $Y=2.405
+ $X2=0 $Y2=0
cc_181 N_A_286_512#_c_194_n N_A_45_164#_c_277_n 0.0236429f $X=3.085 $Y=1.26
+ $X2=0 $Y2=0
cc_182 N_A_286_512#_M1005_g N_VPWR_c_466_n 0.00319878f $X=2.655 $Y=2.405 $X2=0
+ $Y2=0
cc_183 N_A_286_512#_M1016_g N_VPWR_c_466_n 0.00319878f $X=3.085 $Y=2.405 $X2=0
+ $Y2=0
cc_184 N_A_286_512#_c_202_n N_VPWR_c_466_n 0.0228997f $X=1.89 $Y=2.835 $X2=0
+ $Y2=0
cc_185 N_A_286_512#_M1005_g N_VPWR_c_463_n 0.00555719f $X=2.655 $Y=2.405 $X2=0
+ $Y2=0
cc_186 N_A_286_512#_M1016_g N_VPWR_c_463_n 0.00477297f $X=3.085 $Y=2.405 $X2=0
+ $Y2=0
cc_187 N_A_286_512#_c_202_n N_VPWR_c_463_n 0.018252f $X=1.89 $Y=2.835 $X2=0
+ $Y2=0
cc_188 N_A_286_512#_c_202_n N_VPWR_c_469_n 0.0145806f $X=1.89 $Y=2.835 $X2=0
+ $Y2=0
cc_189 N_A_286_512#_c_187_n N_A_463_355#_c_526_n 0.00340356f $X=2.58 $Y=1.26
+ $X2=0 $Y2=0
cc_190 N_A_286_512#_M1005_g N_A_463_355#_c_526_n 0.00412626f $X=2.655 $Y=2.405
+ $X2=0 $Y2=0
cc_191 N_A_286_512#_c_196_n N_A_463_355#_c_526_n 0.0480201f $X=1.89 $Y=2.67
+ $X2=0 $Y2=0
cc_192 N_A_286_512#_c_202_n N_A_463_355#_c_526_n 0.0133428f $X=1.89 $Y=2.835
+ $X2=0 $Y2=0
cc_193 N_A_286_512#_M1005_g N_A_463_355#_c_527_n 0.0120163f $X=2.655 $Y=2.405
+ $X2=0 $Y2=0
cc_194 N_A_286_512#_M1016_g N_A_463_355#_c_527_n 0.0116614f $X=3.085 $Y=2.405
+ $X2=0 $Y2=0
cc_195 N_A_286_512#_c_202_n N_A_463_355#_c_528_n 0.00578441f $X=1.89 $Y=2.835
+ $X2=0 $Y2=0
cc_196 N_A_286_512#_M1005_g N_Y_c_570_n 0.00979852f $X=2.655 $Y=2.405 $X2=0
+ $Y2=0
cc_197 N_A_286_512#_M1016_g N_Y_c_570_n 0.0106715f $X=3.085 $Y=2.405 $X2=0 $Y2=0
cc_198 N_A_286_512#_c_188_n N_Y_c_560_n 8.31293e-19 $X=2.655 $Y=1.185 $X2=0
+ $Y2=0
cc_199 N_A_286_512#_c_190_n N_Y_c_560_n 0.00240919f $X=3.01 $Y=1.26 $X2=0 $Y2=0
cc_200 N_A_286_512#_M1005_g N_Y_c_566_n 0.00628289f $X=2.655 $Y=2.405 $X2=0
+ $Y2=0
cc_201 N_A_286_512#_M1016_g N_Y_c_566_n 0.00193846f $X=3.085 $Y=2.405 $X2=0
+ $Y2=0
cc_202 N_A_286_512#_M1016_g Y 0.0111034f $X=3.085 $Y=2.405 $X2=0 $Y2=0
cc_203 N_A_286_512#_c_191_n N_Y_c_564_n 0.0130505f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_204 N_A_286_512#_c_187_n N_VGND_c_725_n 4.08248e-19 $X=2.58 $Y=1.26 $X2=0
+ $Y2=0
cc_205 N_A_286_512#_c_188_n N_VGND_c_725_n 0.00859225f $X=2.655 $Y=1.185 $X2=0
+ $Y2=0
cc_206 N_A_286_512#_c_191_n N_VGND_c_725_n 5.16405e-19 $X=3.085 $Y=1.185 $X2=0
+ $Y2=0
cc_207 N_A_286_512#_c_188_n N_VGND_c_726_n 6.11179e-19 $X=2.655 $Y=1.185 $X2=0
+ $Y2=0
cc_208 N_A_286_512#_c_191_n N_VGND_c_726_n 0.0100402f $X=3.085 $Y=1.185 $X2=0
+ $Y2=0
cc_209 N_A_286_512#_c_188_n N_VGND_c_732_n 0.00486043f $X=2.655 $Y=1.185 $X2=0
+ $Y2=0
cc_210 N_A_286_512#_c_191_n N_VGND_c_732_n 0.00486043f $X=3.085 $Y=1.185 $X2=0
+ $Y2=0
cc_211 N_A_286_512#_c_188_n N_VGND_c_741_n 0.00824727f $X=2.655 $Y=1.185 $X2=0
+ $Y2=0
cc_212 N_A_286_512#_c_191_n N_VGND_c_741_n 0.00824727f $X=3.085 $Y=1.185 $X2=0
+ $Y2=0
cc_213 N_A_45_164#_c_277_n B 6.57013e-19 $X=3.985 $Y=1.42 $X2=0 $Y2=0
cc_214 N_A_45_164#_M1010_g N_B_c_378_n 0.00171112f $X=3.945 $Y=0.655 $X2=0 $Y2=0
cc_215 N_A_45_164#_c_277_n N_B_c_378_n 0.010182f $X=3.985 $Y=1.42 $X2=0 $Y2=0
cc_216 N_A_45_164#_c_280_n N_VPWR_c_465_n 0.0100339f $X=0.37 $Y=2.77 $X2=0 $Y2=0
cc_217 N_A_45_164#_M1001_g N_VPWR_c_466_n 0.00519759f $X=3.515 $Y=2.405 $X2=0
+ $Y2=0
cc_218 N_A_45_164#_M1017_g N_VPWR_c_466_n 0.00319872f $X=3.985 $Y=2.405 $X2=0
+ $Y2=0
cc_219 N_A_45_164#_M1001_g N_VPWR_c_463_n 0.0102085f $X=3.515 $Y=2.405 $X2=0
+ $Y2=0
cc_220 N_A_45_164#_M1017_g N_VPWR_c_463_n 0.00561909f $X=3.985 $Y=2.405 $X2=0
+ $Y2=0
cc_221 N_A_45_164#_c_280_n N_VPWR_c_463_n 0.00995805f $X=0.37 $Y=2.77 $X2=0
+ $Y2=0
cc_222 N_A_45_164#_c_273_n N_A_463_355#_c_526_n 0.010641f $X=2.555 $Y=1.42 $X2=0
+ $Y2=0
cc_223 N_A_45_164#_M1001_g N_A_463_355#_c_527_n 3.39252e-19 $X=3.515 $Y=2.405
+ $X2=0 $Y2=0
cc_224 N_A_45_164#_M1001_g N_A_463_355#_c_539_n 0.0130502f $X=3.515 $Y=2.405
+ $X2=0 $Y2=0
cc_225 N_A_45_164#_M1017_g N_A_463_355#_c_539_n 0.0129345f $X=3.985 $Y=2.405
+ $X2=0 $Y2=0
cc_226 N_A_45_164#_M1001_g N_Y_c_570_n 7.61713e-19 $X=3.515 $Y=2.405 $X2=0 $Y2=0
cc_227 N_A_45_164#_c_272_n N_Y_c_560_n 0.00626198f $X=2.47 $Y=1.335 $X2=0 $Y2=0
cc_228 N_A_45_164#_c_274_n N_Y_c_560_n 0.0160413f $X=3.66 $Y=1.42 $X2=0 $Y2=0
cc_229 N_A_45_164#_c_274_n N_Y_c_566_n 0.0274572f $X=3.66 $Y=1.42 $X2=0 $Y2=0
cc_230 N_A_45_164#_M1000_g Y 4.36066e-19 $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_231 N_A_45_164#_M1001_g Y 4.58092e-19 $X=3.515 $Y=2.405 $X2=0 $Y2=0
cc_232 N_A_45_164#_M1010_g Y 0.00283117f $X=3.945 $Y=0.655 $X2=0 $Y2=0
cc_233 N_A_45_164#_M1017_g Y 0.00309119f $X=3.985 $Y=2.405 $X2=0 $Y2=0
cc_234 N_A_45_164#_c_274_n Y 0.0130894f $X=3.66 $Y=1.42 $X2=0 $Y2=0
cc_235 N_A_45_164#_c_277_n Y 0.0157363f $X=3.985 $Y=1.42 $X2=0 $Y2=0
cc_236 N_A_45_164#_M1001_g Y 0.0105698f $X=3.515 $Y=2.405 $X2=0 $Y2=0
cc_237 N_A_45_164#_M1017_g Y 0.00670073f $X=3.985 $Y=2.405 $X2=0 $Y2=0
cc_238 N_A_45_164#_c_274_n Y 0.0562338f $X=3.66 $Y=1.42 $X2=0 $Y2=0
cc_239 N_A_45_164#_c_277_n Y 0.00534784f $X=3.985 $Y=1.42 $X2=0 $Y2=0
cc_240 N_A_45_164#_M1017_g N_Y_c_569_n 0.00479471f $X=3.985 $Y=2.405 $X2=0 $Y2=0
cc_241 N_A_45_164#_M1000_g N_Y_c_564_n 0.0132616f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_242 N_A_45_164#_c_274_n N_Y_c_564_n 0.0620149f $X=3.66 $Y=1.42 $X2=0 $Y2=0
cc_243 N_A_45_164#_c_277_n N_Y_c_564_n 0.0017253f $X=3.985 $Y=1.42 $X2=0 $Y2=0
cc_244 N_A_45_164#_M1010_g N_Y_c_565_n 0.0192234f $X=3.945 $Y=0.655 $X2=0 $Y2=0
cc_245 N_A_45_164#_c_277_n N_Y_c_565_n 0.00277671f $X=3.985 $Y=1.42 $X2=0 $Y2=0
cc_246 N_A_45_164#_M1001_g N_A_718_355#_c_658_n 0.00532675f $X=3.515 $Y=2.405
+ $X2=0 $Y2=0
cc_247 N_A_45_164#_M1017_g N_A_718_355#_c_658_n 0.0111086f $X=3.985 $Y=2.405
+ $X2=0 $Y2=0
cc_248 N_A_45_164#_M1017_g N_A_718_355#_c_656_n 0.0136715f $X=3.985 $Y=2.405
+ $X2=0 $Y2=0
cc_249 N_A_45_164#_M1001_g N_A_718_355#_c_657_n 0.00199419f $X=3.515 $Y=2.405
+ $X2=0 $Y2=0
cc_250 N_A_45_164#_M1017_g N_A_718_355#_c_657_n 5.87871e-19 $X=3.985 $Y=2.405
+ $X2=0 $Y2=0
cc_251 N_A_45_164#_M1017_g N_A_919_367#_c_685_n 0.00372553f $X=3.985 $Y=2.405
+ $X2=0 $Y2=0
cc_252 N_A_45_164#_M1017_g N_A_919_367#_c_687_n 0.00108969f $X=3.985 $Y=2.405
+ $X2=0 $Y2=0
cc_253 N_A_45_164#_c_285_n N_VGND_M1006_d 0.00738123f $X=1.21 $Y=1.24 $X2=-0.19
+ $Y2=-0.245
cc_254 N_A_45_164#_c_270_n N_VGND_M1012_s 0.00495319f $X=2.385 $Y=0.745 $X2=0
+ $Y2=0
cc_255 N_A_45_164#_c_272_n N_VGND_M1012_s 0.00654923f $X=2.47 $Y=1.335 $X2=0
+ $Y2=0
cc_256 N_A_45_164#_c_269_n N_VGND_c_724_n 0.0251924f $X=1.125 $Y=1.325 $X2=0
+ $Y2=0
cc_257 N_A_45_164#_c_285_n N_VGND_c_724_n 0.0183479f $X=1.21 $Y=1.24 $X2=0 $Y2=0
cc_258 N_A_45_164#_c_271_n N_VGND_c_724_n 0.0150371f $X=1.295 $Y=0.745 $X2=0
+ $Y2=0
cc_259 N_A_45_164#_c_270_n N_VGND_c_725_n 0.0201648f $X=2.385 $Y=0.745 $X2=0
+ $Y2=0
cc_260 N_A_45_164#_M1000_g N_VGND_c_726_n 0.0100379f $X=3.515 $Y=0.655 $X2=0
+ $Y2=0
cc_261 N_A_45_164#_M1010_g N_VGND_c_726_n 6.10768e-19 $X=3.945 $Y=0.655 $X2=0
+ $Y2=0
cc_262 N_A_45_164#_c_270_n N_VGND_c_730_n 0.0169405f $X=2.385 $Y=0.745 $X2=0
+ $Y2=0
cc_263 N_A_45_164#_c_271_n N_VGND_c_730_n 0.00327186f $X=1.295 $Y=0.745 $X2=0
+ $Y2=0
cc_264 N_A_45_164#_M1000_g N_VGND_c_738_n 0.00486043f $X=3.515 $Y=0.655 $X2=0
+ $Y2=0
cc_265 N_A_45_164#_M1010_g N_VGND_c_738_n 0.00486043f $X=3.945 $Y=0.655 $X2=0
+ $Y2=0
cc_266 N_A_45_164#_M1000_g N_VGND_c_739_n 5.83998e-19 $X=3.515 $Y=0.655 $X2=0
+ $Y2=0
cc_267 N_A_45_164#_M1010_g N_VGND_c_739_n 0.0129174f $X=3.945 $Y=0.655 $X2=0
+ $Y2=0
cc_268 N_A_45_164#_M1000_g N_VGND_c_741_n 0.00824727f $X=3.515 $Y=0.655 $X2=0
+ $Y2=0
cc_269 N_A_45_164#_M1010_g N_VGND_c_741_n 0.004522f $X=3.945 $Y=0.655 $X2=0
+ $Y2=0
cc_270 N_A_45_164#_c_268_n N_VGND_c_741_n 0.00954814f $X=0.35 $Y=1.03 $X2=0
+ $Y2=0
cc_271 N_A_45_164#_c_270_n N_VGND_c_741_n 0.0287897f $X=2.385 $Y=0.745 $X2=0
+ $Y2=0
cc_272 N_A_45_164#_c_271_n N_VGND_c_741_n 0.00506459f $X=1.295 $Y=0.745 $X2=0
+ $Y2=0
cc_273 N_B_c_376_n N_A_c_427_n 0.0154827f $X=5.285 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_274 N_B_c_378_n N_A_M1003_g 0.024206f $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_275 N_B_c_378_n N_A_c_432_n 0.0262037f $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_276 N_B_c_380_n N_VPWR_c_464_n 0.00138929f $X=5.365 $Y=1.725 $X2=0 $Y2=0
cc_277 N_B_c_379_n N_VPWR_c_466_n 0.00357842f $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_278 N_B_c_380_n N_VPWR_c_466_n 0.00547432f $X=5.365 $Y=1.725 $X2=0 $Y2=0
cc_279 N_B_c_379_n N_VPWR_c_463_n 0.00675085f $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_280 N_B_c_380_n N_VPWR_c_463_n 0.00990114f $X=5.365 $Y=1.725 $X2=0 $Y2=0
cc_281 N_B_c_375_n N_Y_c_598_n 0.0120695f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_282 B N_Y_c_598_n 0.023535f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_283 N_B_c_378_n N_Y_c_598_n 0.00739756f $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_284 N_B_c_376_n N_Y_c_561_n 0.00938454f $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_285 N_B_c_378_n N_Y_c_561_n 0.00910935f $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_286 N_B_c_375_n N_Y_c_562_n 0.00734515f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_287 N_B_c_376_n N_Y_c_562_n 2.39771e-19 $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_288 B N_Y_c_562_n 0.00363741f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_289 N_B_c_378_n N_Y_c_562_n 0.0106656f $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_290 N_B_c_375_n Y 2.94875e-19 $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_291 B Y 0.0266512f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_292 N_B_c_378_n Y 0.00401225f $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_293 N_B_c_379_n N_Y_c_569_n 4.96414e-19 $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_294 N_B_c_378_n N_Y_c_569_n 3.81235e-19 $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_295 N_B_c_375_n N_Y_c_565_n 0.00245601f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_296 N_B_c_379_n N_A_718_355#_c_656_n 0.0125611f $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_297 N_B_c_379_n N_A_718_355#_c_664_n 5.89773e-19 $X=4.935 $Y=1.725 $X2=0
+ $Y2=0
cc_298 N_B_c_380_n N_A_718_355#_c_664_n 0.00193114f $X=5.365 $Y=1.725 $X2=0
+ $Y2=0
cc_299 N_B_c_379_n N_A_718_355#_c_666_n 0.0155223f $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_300 N_B_c_380_n N_A_718_355#_c_666_n 0.00951647f $X=5.365 $Y=1.725 $X2=0
+ $Y2=0
cc_301 N_B_c_379_n N_A_919_367#_c_686_n 0.0113732f $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_302 N_B_c_380_n N_A_919_367#_c_686_n 0.0104512f $X=5.365 $Y=1.725 $X2=0 $Y2=0
cc_303 N_B_c_378_n N_A_919_367#_c_686_n 0.0205981f $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_304 B N_A_919_367#_c_687_n 0.0134257f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_305 N_B_c_378_n N_A_919_367#_c_687_n 0.0101945f $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_306 N_B_c_375_n N_VGND_c_727_n 6.15012e-19 $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_307 N_B_c_376_n N_VGND_c_727_n 0.0109991f $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_308 N_B_c_378_n N_VGND_c_727_n 2.65959e-19 $X=5.285 $Y=1.455 $X2=0 $Y2=0
cc_309 N_B_c_375_n N_VGND_c_735_n 0.00486043f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_310 N_B_c_376_n N_VGND_c_735_n 0.00486043f $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_311 N_B_c_375_n N_VGND_c_739_n 0.012932f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_312 N_B_c_376_n N_VGND_c_739_n 5.83998e-19 $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_313 N_B_c_375_n N_VGND_c_741_n 0.00450478f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_314 N_B_c_376_n N_VGND_c_741_n 0.00824727f $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_315 N_A_M1003_g N_VPWR_c_464_n 0.0168412f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_316 N_A_M1013_g N_VPWR_c_464_n 0.0176671f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_317 N_A_M1003_g N_VPWR_c_466_n 0.00486043f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A_M1013_g N_VPWR_c_467_n 0.00486043f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_319 N_A_M1003_g N_VPWR_c_463_n 0.0082726f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_320 N_A_M1013_g N_VPWR_c_463_n 0.00919827f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_321 N_A_c_427_n N_Y_c_561_n 0.00990953f $X=5.715 $Y=1.185 $X2=0 $Y2=0
cc_322 N_A_c_429_n N_Y_c_561_n 0.00349191f $X=6.145 $Y=1.185 $X2=0 $Y2=0
cc_323 A N_Y_c_561_n 0.00401496f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_324 N_A_c_432_n N_Y_c_561_n 0.0136269f $X=6.225 $Y=1.35 $X2=0 $Y2=0
cc_325 N_A_M1003_g N_A_919_367#_c_688_n 0.0154654f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_326 N_A_M1013_g N_A_919_367#_c_688_n 0.016638f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_327 A N_A_919_367#_c_688_n 0.0332854f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_328 N_A_c_432_n N_A_919_367#_c_688_n 0.00849533f $X=6.225 $Y=1.35 $X2=0 $Y2=0
cc_329 N_A_c_432_n N_A_919_367#_c_690_n 8.81383e-19 $X=6.225 $Y=1.35 $X2=0 $Y2=0
cc_330 N_A_c_427_n N_VGND_c_727_n 0.0110093f $X=5.715 $Y=1.185 $X2=0 $Y2=0
cc_331 N_A_c_429_n N_VGND_c_727_n 6.28154e-19 $X=6.145 $Y=1.185 $X2=0 $Y2=0
cc_332 N_A_c_427_n N_VGND_c_729_n 6.64931e-19 $X=5.715 $Y=1.185 $X2=0 $Y2=0
cc_333 N_A_c_429_n N_VGND_c_729_n 0.0163045f $X=6.145 $Y=1.185 $X2=0 $Y2=0
cc_334 A N_VGND_c_729_n 0.0246699f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_335 N_A_c_432_n N_VGND_c_729_n 0.00619872f $X=6.225 $Y=1.35 $X2=0 $Y2=0
cc_336 N_A_c_427_n N_VGND_c_736_n 0.00486043f $X=5.715 $Y=1.185 $X2=0 $Y2=0
cc_337 N_A_c_429_n N_VGND_c_736_n 0.00486043f $X=6.145 $Y=1.185 $X2=0 $Y2=0
cc_338 N_A_c_427_n N_VGND_c_741_n 0.00824727f $X=5.715 $Y=1.185 $X2=0 $Y2=0
cc_339 N_A_c_429_n N_VGND_c_741_n 0.00824727f $X=6.145 $Y=1.185 $X2=0 $Y2=0
cc_340 N_VPWR_c_466_n N_A_463_355#_c_527_n 0.0572829f $X=5.845 $Y=3.33 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_463_n N_A_463_355#_c_527_n 0.0319816f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_466_n N_A_463_355#_c_528_n 0.0186386f $X=5.845 $Y=3.33 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_463_n N_A_463_355#_c_528_n 0.0101082f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_463_n N_A_718_355#_M1009_d 0.00223559f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_466_n N_A_718_355#_c_656_n 0.0661868f $X=5.845 $Y=3.33 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_463_n N_A_718_355#_c_656_n 0.0389906f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_466_n N_A_718_355#_c_657_n 0.0237238f $X=5.845 $Y=3.33 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_463_n N_A_718_355#_c_657_n 0.0128032f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_466_n N_A_718_355#_c_664_n 0.01906f $X=5.845 $Y=3.33 $X2=0 $Y2=0
cc_350 N_VPWR_c_463_n N_A_718_355#_c_664_n 0.0124545f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_463_n N_A_919_367#_M1009_s 0.0021598f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_352 N_VPWR_c_463_n N_A_919_367#_M1019_s 0.00536646f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_353 N_VPWR_c_463_n N_A_919_367#_M1013_d 0.00371702f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_354 N_VPWR_c_466_n N_A_919_367#_c_706_n 0.0124525f $X=5.845 $Y=3.33 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_463_n N_A_919_367#_c_706_n 0.00730901f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_356 N_VPWR_M1003_s N_A_919_367#_c_688_n 0.00176461f $X=5.87 $Y=1.835 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_464_n N_A_919_367#_c_688_n 0.0170777f $X=6.01 $Y=2.11 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_467_n N_A_919_367#_c_689_n 0.0178111f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_463_n N_A_919_367#_c_689_n 0.0100304f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_360 N_A_463_355#_c_527_n N_Y_M1005_d 0.00176461f $X=3.205 $Y=2.99 $X2=0 $Y2=0
cc_361 N_A_463_355#_c_527_n N_Y_c_570_n 0.0159805f $X=3.205 $Y=2.99 $X2=0 $Y2=0
cc_362 N_A_463_355#_c_526_n N_Y_c_566_n 0.00455684f $X=2.44 $Y=1.92 $X2=0 $Y2=0
cc_363 N_A_463_355#_M1016_s Y 0.00176461f $X=3.16 $Y=1.775 $X2=0 $Y2=0
cc_364 N_A_463_355#_c_549_p Y 0.0135055f $X=3.31 $Y=2.185 $X2=0 $Y2=0
cc_365 N_A_463_355#_c_539_n Y 0.0308231f $X=4.085 $Y=2.1 $X2=0 $Y2=0
cc_366 N_A_463_355#_M1017_s N_Y_c_569_n 0.00218937f $X=4.06 $Y=1.775 $X2=0 $Y2=0
cc_367 N_A_463_355#_c_539_n N_Y_c_569_n 0.00484117f $X=4.085 $Y=2.1 $X2=0 $Y2=0
cc_368 N_A_463_355#_c_529_n N_Y_c_569_n 0.0102316f $X=4.2 $Y=2.18 $X2=0 $Y2=0
cc_369 N_A_463_355#_c_539_n N_A_718_355#_M1001_d 0.00418803f $X=4.085 $Y=2.1
+ $X2=-0.19 $Y2=1.655
cc_370 N_A_463_355#_c_539_n N_A_718_355#_c_658_n 0.0173659f $X=4.085 $Y=2.1
+ $X2=0 $Y2=0
cc_371 N_A_463_355#_M1017_s N_A_718_355#_c_656_n 0.002818f $X=4.06 $Y=1.775
+ $X2=0 $Y2=0
cc_372 N_A_463_355#_c_529_n N_A_718_355#_c_656_n 0.0189969f $X=4.2 $Y=2.18 $X2=0
+ $Y2=0
cc_373 N_A_463_355#_c_527_n N_A_718_355#_c_657_n 0.00902112f $X=3.205 $Y=2.99
+ $X2=0 $Y2=0
cc_374 N_A_463_355#_c_529_n N_A_919_367#_c_685_n 0.0547101f $X=4.2 $Y=2.18 $X2=0
+ $Y2=0
cc_375 Y N_A_718_355#_M1001_d 0.00219516f $X=3.995 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_376 N_Y_c_598_n N_A_919_367#_c_686_n 0.00150027f $X=4.885 $Y=0.927 $X2=0
+ $Y2=0
cc_377 N_Y_c_561_n N_A_919_367#_c_686_n 0.0105313f $X=5.835 $Y=1.15 $X2=0 $Y2=0
cc_378 N_Y_c_562_n N_A_919_367#_c_686_n 0.0100284f $X=5.025 $Y=0.927 $X2=0 $Y2=0
cc_379 N_Y_c_598_n N_A_919_367#_c_687_n 0.00181628f $X=4.885 $Y=0.927 $X2=0
+ $Y2=0
cc_380 N_Y_c_569_n N_A_919_367#_c_687_n 0.00939809f $X=4.112 $Y=1.675 $X2=0
+ $Y2=0
cc_381 N_Y_c_561_n N_A_919_367#_c_688_n 0.0122066f $X=5.835 $Y=1.15 $X2=0 $Y2=0
cc_382 N_Y_c_561_n N_A_919_367#_c_690_n 0.00803354f $X=5.835 $Y=1.15 $X2=0 $Y2=0
cc_383 N_Y_c_564_n N_VGND_M1015_s 0.00176461f $X=3.635 $Y=1.002 $X2=0 $Y2=0
cc_384 N_Y_c_598_n N_VGND_M1010_s 0.0179193f $X=4.885 $Y=0.927 $X2=0 $Y2=0
cc_385 N_Y_c_565_n N_VGND_M1010_s 0.00302344f $X=4.23 $Y=1.002 $X2=0 $Y2=0
cc_386 N_Y_c_561_n N_VGND_M1008_s 0.00180746f $X=5.835 $Y=1.15 $X2=0 $Y2=0
cc_387 N_Y_c_564_n N_VGND_c_726_n 0.0170777f $X=3.635 $Y=1.002 $X2=0 $Y2=0
cc_388 N_Y_c_561_n N_VGND_c_727_n 0.0163515f $X=5.835 $Y=1.15 $X2=0 $Y2=0
cc_389 N_Y_c_640_p N_VGND_c_732_n 0.0124525f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_390 N_Y_c_641_p N_VGND_c_735_n 0.0124525f $X=5.07 $Y=0.42 $X2=0 $Y2=0
cc_391 N_Y_c_642_p N_VGND_c_736_n 0.0124525f $X=5.93 $Y=0.42 $X2=0 $Y2=0
cc_392 N_Y_c_643_p N_VGND_c_738_n 0.0123249f $X=3.73 $Y=0.42 $X2=0 $Y2=0
cc_393 N_Y_c_565_n N_VGND_c_739_n 0.0554478f $X=4.23 $Y=1.002 $X2=0 $Y2=0
cc_394 N_Y_M1012_d N_VGND_c_741_n 0.00536646f $X=2.73 $Y=0.235 $X2=0 $Y2=0
cc_395 N_Y_M1000_d N_VGND_c_741_n 0.00405668f $X=3.59 $Y=0.235 $X2=0 $Y2=0
cc_396 N_Y_M1002_d N_VGND_c_741_n 0.00408418f $X=4.93 $Y=0.235 $X2=0 $Y2=0
cc_397 N_Y_M1004_s N_VGND_c_741_n 0.00536646f $X=5.79 $Y=0.235 $X2=0 $Y2=0
cc_398 N_Y_c_640_p N_VGND_c_741_n 0.00730901f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_399 N_Y_c_643_p N_VGND_c_741_n 0.00728036f $X=3.73 $Y=0.42 $X2=0 $Y2=0
cc_400 N_Y_c_598_n N_VGND_c_741_n 0.00219744f $X=4.885 $Y=0.927 $X2=0 $Y2=0
cc_401 N_Y_c_641_p N_VGND_c_741_n 0.00730901f $X=5.07 $Y=0.42 $X2=0 $Y2=0
cc_402 N_Y_c_642_p N_VGND_c_741_n 0.00730901f $X=5.93 $Y=0.42 $X2=0 $Y2=0
cc_403 N_Y_c_562_n N_VGND_c_741_n 0.00293069f $X=5.025 $Y=0.927 $X2=0 $Y2=0
cc_404 N_Y_c_565_n N_VGND_c_741_n 0.00794901f $X=4.23 $Y=1.002 $X2=0 $Y2=0
cc_405 N_A_718_355#_c_656_n N_A_919_367#_M1009_s 0.00495471f $X=4.985 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_406 N_A_718_355#_c_656_n N_A_919_367#_c_685_n 0.0189128f $X=4.985 $Y=2.99
+ $X2=0 $Y2=0
cc_407 N_A_718_355#_M1009_d N_A_919_367#_c_686_n 0.00176461f $X=5.01 $Y=1.835
+ $X2=0 $Y2=0
cc_408 N_A_718_355#_c_666_n N_A_919_367#_c_686_n 0.0170777f $X=5.15 $Y=2.11
+ $X2=0 $Y2=0
