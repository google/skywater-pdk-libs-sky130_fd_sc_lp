* File: sky130_fd_sc_lp__o311a_lp.pxi.spice
* Created: Wed Sep  2 10:23:17 2020
* 
x_PM_SKY130_FD_SC_LP__O311A_LP%A_84_115# N_A_84_115#_M1004_d N_A_84_115#_M1010_d
+ N_A_84_115#_M1005_d N_A_84_115#_c_73_n N_A_84_115#_M1001_g N_A_84_115#_M1009_g
+ N_A_84_115#_M1011_g N_A_84_115#_c_74_n N_A_84_115#_c_80_n N_A_84_115#_c_75_n
+ N_A_84_115#_c_76_n N_A_84_115#_c_83_n N_A_84_115#_c_89_p N_A_84_115#_c_131_p
+ N_A_84_115#_c_110_p N_A_84_115#_c_77_n N_A_84_115#_c_78_n N_A_84_115#_c_85_n
+ N_A_84_115#_c_102_p N_A_84_115#_c_86_n PM_SKY130_FD_SC_LP__O311A_LP%A_84_115#
x_PM_SKY130_FD_SC_LP__O311A_LP%A1 N_A1_M1012_g N_A1_M1006_g N_A1_c_165_n
+ N_A1_c_166_n A1 N_A1_c_168_n N_A1_c_169_n PM_SKY130_FD_SC_LP__O311A_LP%A1
x_PM_SKY130_FD_SC_LP__O311A_LP%A2 N_A2_M1003_g N_A2_M1002_g A2 N_A2_c_208_n
+ PM_SKY130_FD_SC_LP__O311A_LP%A2
x_PM_SKY130_FD_SC_LP__O311A_LP%A3 N_A3_M1010_g N_A3_M1007_g A3 N_A3_c_246_n
+ PM_SKY130_FD_SC_LP__O311A_LP%A3
x_PM_SKY130_FD_SC_LP__O311A_LP%B1 N_B1_M1000_g N_B1_M1008_g B1 N_B1_c_282_n
+ N_B1_c_283_n PM_SKY130_FD_SC_LP__O311A_LP%B1
x_PM_SKY130_FD_SC_LP__O311A_LP%C1 N_C1_c_318_n N_C1_M1004_g N_C1_M1005_g
+ N_C1_c_319_n C1 N_C1_c_320_n N_C1_c_321_n N_C1_c_322_n
+ PM_SKY130_FD_SC_LP__O311A_LP%C1
x_PM_SKY130_FD_SC_LP__O311A_LP%X N_X_M1001_s N_X_M1009_s N_X_c_357_n N_X_c_354_n
+ X X X PM_SKY130_FD_SC_LP__O311A_LP%X
x_PM_SKY130_FD_SC_LP__O311A_LP%VPWR N_VPWR_M1009_d N_VPWR_M1000_d N_VPWR_c_377_n
+ N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n VPWR N_VPWR_c_381_n
+ N_VPWR_c_376_n N_VPWR_c_383_n PM_SKY130_FD_SC_LP__O311A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O311A_LP%VGND N_VGND_M1011_d N_VGND_M1002_d N_VGND_c_425_n
+ N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n VGND N_VGND_c_429_n
+ N_VGND_c_430_n N_VGND_c_431_n N_VGND_c_432_n PM_SKY130_FD_SC_LP__O311A_LP%VGND
x_PM_SKY130_FD_SC_LP__O311A_LP%A_273_141# N_A_273_141#_M1006_d
+ N_A_273_141#_M1007_d N_A_273_141#_c_464_n N_A_273_141#_c_465_n
+ N_A_273_141#_c_466_n PM_SKY130_FD_SC_LP__O311A_LP%A_273_141#
cc_1 VNB N_A_84_115#_c_73_n 0.0307487f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.2
cc_2 VNB N_A_84_115#_c_74_n 0.0237717f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.35
cc_3 VNB N_A_84_115#_c_75_n 0.00314989f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.43
cc_4 VNB N_A_84_115#_c_76_n 0.0237302f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.43
cc_5 VNB N_A_84_115#_c_77_n 0.0249458f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=0.905
cc_6 VNB N_A_84_115#_c_78_n 0.0294298f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=2.1
cc_7 VNB N_A1_c_165_n 0.0157117f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.2
cc_8 VNB N_A1_c_166_n 0.0135841f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.915
cc_9 VNB A1 0.00317003f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.915
cc_10 VNB N_A1_c_168_n 0.00954431f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.595
cc_11 VNB N_A1_c_169_n 0.0139524f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.2
cc_12 VNB N_A2_M1002_g 0.0374391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A2 0.00219679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_208_n 0.00951667f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.915
cc_15 VNB N_A3_M1007_g 0.0353254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A3 8.962e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_c_246_n 0.0113653f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.915
cc_18 VNB N_B1_M1008_g 0.0345835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_282_n 0.0109495f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.915
cc_20 VNB N_B1_c_283_n 0.00385043f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.935
cc_21 VNB N_C1_c_318_n 0.0195873f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=0.705
cc_22 VNB N_C1_c_319_n 0.0173709f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.915
cc_23 VNB N_C1_c_320_n 0.00976901f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.2
cc_24 VNB N_C1_c_321_n 0.00387077f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.915
cc_25 VNB N_C1_c_322_n 0.0145002f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.915
cc_26 VNB N_X_c_354_n 0.0266464f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.935
cc_27 VNB X 0.0246326f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.595
cc_28 VNB X 0.00666148f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.43
cc_29 VNB N_VPWR_c_376_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.1
cc_30 VNB N_VGND_c_425_n 0.0293963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_426_n 0.0385937f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.935
cc_32 VNB N_VGND_c_427_n 0.0286968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_428_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.2
cc_34 VNB N_VGND_c_429_n 0.0207228f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.935
cc_35 VNB N_VGND_c_430_n 0.0514828f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.935
cc_36 VNB N_VGND_c_431_n 0.266571f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.1
cc_37 VNB N_VGND_c_432_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_273_141#_c_464_n 0.0220371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_273_141#_c_465_n 0.00394084f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.915
cc_40 VNB N_A_273_141#_c_466_n 0.0135735f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.595
cc_41 VPB N_A_84_115#_M1009_g 0.029543f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.595
cc_42 VPB N_A_84_115#_c_80_n 0.0161899f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.935
cc_43 VPB N_A_84_115#_c_75_n 6.15811e-19 $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.43
cc_44 VPB N_A_84_115#_c_76_n 0.00717714f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.43
cc_45 VPB N_A_84_115#_c_83_n 0.00159614f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.1
cc_46 VPB N_A_84_115#_c_78_n 0.0210831f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=2.1
cc_47 VPB N_A_84_115#_c_85_n 0.00119146f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.935
cc_48 VPB N_A_84_115#_c_86_n 0.0388736f $X=-0.19 $Y=1.655 $X2=3.54 $Y2=2.265
cc_49 VPB N_A1_M1012_g 0.0271762f $X=-0.19 $Y=1.655 $X2=3.4 $Y2=2.095
cc_50 VPB A1 7.39101e-19 $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.915
cc_51 VPB N_A1_c_168_n 0.0203031f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.595
cc_52 VPB N_A2_M1003_g 0.026558f $X=-0.19 $Y=1.655 $X2=3.4 $Y2=2.095
cc_53 VPB A2 7.48576e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A2_c_208_n 0.0203221f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.915
cc_55 VPB N_A3_M1010_g 0.0296778f $X=-0.19 $Y=1.655 $X2=3.4 $Y2=2.095
cc_56 VPB A3 0.00165706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A3_c_246_n 0.0160112f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.915
cc_58 VPB N_B1_M1000_g 0.0269272f $X=-0.19 $Y=1.655 $X2=3.4 $Y2=2.095
cc_59 VPB N_B1_c_282_n 0.0184058f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.915
cc_60 VPB N_B1_c_283_n 0.00249228f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.935
cc_61 VPB N_C1_M1005_g 0.0301967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_C1_c_320_n 0.0201046f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.2
cc_63 VPB N_C1_c_321_n 0.00268919f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.915
cc_64 VPB N_X_c_357_n 0.0378297f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.915
cc_65 VPB N_X_c_354_n 0.0214884f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.935
cc_66 VPB N_VPWR_c_377_n 0.00283282f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.915
cc_67 VPB N_VPWR_c_378_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.595
cc_68 VPB N_VPWR_c_379_n 0.0545752f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.915
cc_69 VPB N_VPWR_c_380_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.915
cc_70 VPB N_VPWR_c_381_n 0.0198732f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.935
cc_71 VPB N_VPWR_c_376_n 0.045096f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.1
cc_72 VPB N_VPWR_c_383_n 0.0239046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 N_A_84_115#_M1009_g N_A1_M1012_g 0.0353532f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_74 N_A_84_115#_c_80_n N_A1_M1012_g 6.84611e-19 $X=0.6 $Y=1.935 $X2=0 $Y2=0
cc_75 N_A_84_115#_c_89_p N_A1_M1012_g 0.0226332f $X=2.295 $Y=2.185 $X2=0 $Y2=0
cc_76 N_A_84_115#_c_85_n N_A1_M1012_g 0.00366421f $X=0.63 $Y=1.935 $X2=0 $Y2=0
cc_77 N_A_84_115#_c_73_n N_A1_c_165_n 0.0104551f $X=0.495 $Y=1.2 $X2=0 $Y2=0
cc_78 N_A_84_115#_c_74_n N_A1_c_166_n 0.00882243f $X=0.675 $Y=1.35 $X2=0 $Y2=0
cc_79 N_A_84_115#_c_75_n N_A1_c_166_n 4.35602e-19 $X=0.615 $Y=1.43 $X2=0 $Y2=0
cc_80 N_A_84_115#_c_75_n A1 0.0283725f $X=0.615 $Y=1.43 $X2=0 $Y2=0
cc_81 N_A_84_115#_c_76_n A1 5.323e-19 $X=0.615 $Y=1.43 $X2=0 $Y2=0
cc_82 N_A_84_115#_c_89_p A1 0.0201562f $X=2.295 $Y=2.185 $X2=0 $Y2=0
cc_83 N_A_84_115#_c_75_n N_A1_c_168_n 0.00188269f $X=0.615 $Y=1.43 $X2=0 $Y2=0
cc_84 N_A_84_115#_c_76_n N_A1_c_168_n 0.0206381f $X=0.615 $Y=1.43 $X2=0 $Y2=0
cc_85 N_A_84_115#_c_75_n N_A1_c_169_n 0.00409763f $X=0.615 $Y=1.43 $X2=0 $Y2=0
cc_86 N_A_84_115#_c_76_n N_A1_c_169_n 0.00650037f $X=0.615 $Y=1.43 $X2=0 $Y2=0
cc_87 N_A_84_115#_c_89_p N_A2_M1003_g 0.022271f $X=2.295 $Y=2.185 $X2=0 $Y2=0
cc_88 N_A_84_115#_c_102_p N_A2_M1003_g 0.00341252f $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_89 N_A_84_115#_c_89_p A2 0.0208926f $X=2.295 $Y=2.185 $X2=0 $Y2=0
cc_90 N_A_84_115#_c_89_p N_A2_c_208_n 4.20092e-19 $X=2.295 $Y=2.185 $X2=0 $Y2=0
cc_91 N_A_84_115#_c_89_p N_A3_M1010_g 0.0189985f $X=2.295 $Y=2.185 $X2=0 $Y2=0
cc_92 N_A_84_115#_c_102_p N_A3_M1010_g 0.0202005f $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_93 N_A_84_115#_c_89_p A3 0.0139163f $X=2.295 $Y=2.185 $X2=0 $Y2=0
cc_94 N_A_84_115#_c_102_p A3 0.00281361f $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_95 N_A_84_115#_c_102_p N_A3_c_246_n 0.00230525f $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_96 N_A_84_115#_c_110_p N_B1_M1000_g 0.0186609f $X=3.455 $Y=2.185 $X2=0 $Y2=0
cc_97 N_A_84_115#_c_102_p N_B1_M1000_g 0.0170439f $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_98 N_A_84_115#_c_77_n N_B1_M1008_g 8.90029e-19 $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_99 N_A_84_115#_c_110_p N_B1_c_282_n 0.00199529f $X=3.455 $Y=2.185 $X2=0 $Y2=0
cc_100 N_A_84_115#_c_110_p N_B1_c_283_n 0.0161465f $X=3.455 $Y=2.185 $X2=0 $Y2=0
cc_101 N_A_84_115#_c_102_p N_B1_c_283_n 0.0053697f $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_102 N_A_84_115#_c_77_n N_C1_c_318_n 0.00631841f $X=3.58 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_84_115#_c_78_n N_C1_c_318_n 0.00304886f $X=3.665 $Y=2.1 $X2=-0.19
+ $Y2=-0.245
cc_104 N_A_84_115#_c_110_p N_C1_M1005_g 0.0200748f $X=3.455 $Y=2.185 $X2=0 $Y2=0
cc_105 N_A_84_115#_c_78_n N_C1_M1005_g 0.00633844f $X=3.665 $Y=2.1 $X2=0 $Y2=0
cc_106 N_A_84_115#_c_102_p N_C1_M1005_g 9.91286e-19 $X=2.46 $Y=2.265 $X2=0 $Y2=0
cc_107 N_A_84_115#_c_77_n N_C1_c_319_n 0.00362229f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_108 N_A_84_115#_c_78_n N_C1_c_319_n 0.0110014f $X=3.665 $Y=2.1 $X2=0 $Y2=0
cc_109 N_A_84_115#_c_77_n N_C1_c_320_n 0.00257889f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_110 N_A_84_115#_c_78_n N_C1_c_320_n 0.00804858f $X=3.665 $Y=2.1 $X2=0 $Y2=0
cc_111 N_A_84_115#_c_86_n N_C1_c_320_n 0.00105123f $X=3.54 $Y=2.265 $X2=0 $Y2=0
cc_112 N_A_84_115#_c_110_p N_C1_c_321_n 0.0246194f $X=3.455 $Y=2.185 $X2=0 $Y2=0
cc_113 N_A_84_115#_c_77_n N_C1_c_321_n 0.00843191f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_114 N_A_84_115#_c_78_n N_C1_c_321_n 0.0282569f $X=3.665 $Y=2.1 $X2=0 $Y2=0
cc_115 N_A_84_115#_c_78_n N_C1_c_322_n 2.06648e-19 $X=3.665 $Y=2.1 $X2=0 $Y2=0
cc_116 N_A_84_115#_M1009_g N_X_c_357_n 0.022679f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_117 N_A_84_115#_c_131_p N_X_c_357_n 0.0118901f $X=0.81 $Y=2.185 $X2=0 $Y2=0
cc_118 N_A_84_115#_c_85_n N_X_c_357_n 6.45782e-19 $X=0.63 $Y=1.935 $X2=0 $Y2=0
cc_119 N_A_84_115#_c_73_n N_X_c_354_n 0.020737f $X=0.495 $Y=1.2 $X2=0 $Y2=0
cc_120 N_A_84_115#_M1009_g N_X_c_354_n 0.00303969f $X=0.56 $Y=2.595 $X2=0 $Y2=0
cc_121 N_A_84_115#_c_75_n N_X_c_354_n 0.0484794f $X=0.615 $Y=1.43 $X2=0 $Y2=0
cc_122 N_A_84_115#_c_83_n N_X_c_354_n 0.00519041f $X=0.725 $Y=2.1 $X2=0 $Y2=0
cc_123 N_A_84_115#_c_73_n X 0.00980611f $X=0.495 $Y=1.2 $X2=0 $Y2=0
cc_124 N_A_84_115#_c_73_n X 0.00407909f $X=0.495 $Y=1.2 $X2=0 $Y2=0
cc_125 N_A_84_115#_c_89_p N_VPWR_M1009_d 0.00843554f $X=2.295 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_126 N_A_84_115#_c_131_p N_VPWR_M1009_d 7.59612e-19 $X=0.81 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_84_115#_c_110_p N_VPWR_M1000_d 0.00630649f $X=3.455 $Y=2.185 $X2=0
+ $Y2=0
cc_128 N_A_84_115#_M1009_g N_VPWR_c_377_n 0.0203558f $X=0.56 $Y=2.595 $X2=0
+ $Y2=0
cc_129 N_A_84_115#_c_80_n N_VPWR_c_377_n 2.71602e-19 $X=0.6 $Y=1.935 $X2=0 $Y2=0
cc_130 N_A_84_115#_c_89_p N_VPWR_c_377_n 0.013451f $X=2.295 $Y=2.185 $X2=0 $Y2=0
cc_131 N_A_84_115#_c_131_p N_VPWR_c_377_n 0.0077692f $X=0.81 $Y=2.185 $X2=0
+ $Y2=0
cc_132 N_A_84_115#_c_110_p N_VPWR_c_378_n 0.016484f $X=3.455 $Y=2.185 $X2=0
+ $Y2=0
cc_133 N_A_84_115#_c_102_p N_VPWR_c_378_n 0.0389751f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_134 N_A_84_115#_c_102_p N_VPWR_c_379_n 0.0178162f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_135 N_A_84_115#_c_86_n N_VPWR_c_381_n 0.0194114f $X=3.54 $Y=2.265 $X2=0 $Y2=0
cc_136 N_A_84_115#_M1010_d N_VPWR_c_376_n 0.0023187f $X=2.32 $Y=2.095 $X2=0
+ $Y2=0
cc_137 N_A_84_115#_M1005_d N_VPWR_c_376_n 0.0042346f $X=3.4 $Y=2.095 $X2=0 $Y2=0
cc_138 N_A_84_115#_M1009_g N_VPWR_c_376_n 0.0145374f $X=0.56 $Y=2.595 $X2=0
+ $Y2=0
cc_139 N_A_84_115#_c_102_p N_VPWR_c_376_n 0.0123708f $X=2.46 $Y=2.265 $X2=0
+ $Y2=0
cc_140 N_A_84_115#_c_86_n N_VPWR_c_376_n 0.0113316f $X=3.54 $Y=2.265 $X2=0 $Y2=0
cc_141 N_A_84_115#_M1009_g N_VPWR_c_383_n 0.00840199f $X=0.56 $Y=2.595 $X2=0
+ $Y2=0
cc_142 N_A_84_115#_c_89_p A_258_419# 0.0096152f $X=2.295 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_84_115#_c_89_p A_356_419# 0.0127797f $X=2.295 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A_84_115#_c_73_n N_VGND_c_425_n 0.0124358f $X=0.495 $Y=1.2 $X2=0 $Y2=0
cc_145 N_A_84_115#_c_73_n N_VGND_c_427_n 0.00636678f $X=0.495 $Y=1.2 $X2=0 $Y2=0
cc_146 N_A_84_115#_c_77_n N_VGND_c_430_n 0.00877597f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_147 N_A_84_115#_c_73_n N_VGND_c_431_n 0.0075243f $X=0.495 $Y=1.2 $X2=0 $Y2=0
cc_148 N_A_84_115#_c_77_n N_VGND_c_431_n 0.0163788f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_149 N_A_84_115#_c_77_n N_A_273_141#_c_465_n 0.0115237f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_150 N_A_84_115#_c_73_n N_A_273_141#_c_466_n 4.24401e-19 $X=0.495 $Y=1.2 $X2=0
+ $Y2=0
cc_151 N_A1_M1012_g N_A2_M1003_g 0.078246f $X=1.165 $Y=2.595 $X2=0 $Y2=0
cc_152 N_A1_c_165_n N_A2_M1002_g 0.0161269f $X=1.267 $Y=1.2 $X2=0 $Y2=0
cc_153 N_A1_c_169_n N_A2_M1002_g 0.00994519f $X=1.155 $Y=1.59 $X2=0 $Y2=0
cc_154 A1 A2 0.0235844f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A1_c_168_n A2 0.00114936f $X=1.155 $Y=1.755 $X2=0 $Y2=0
cc_156 N_A1_c_169_n A2 2.52374e-19 $X=1.155 $Y=1.59 $X2=0 $Y2=0
cc_157 A1 N_A2_c_208_n 0.00114936f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A1_c_168_n N_A2_c_208_n 0.0201104f $X=1.155 $Y=1.755 $X2=0 $Y2=0
cc_159 N_A1_M1012_g N_X_c_357_n 9.77743e-19 $X=1.165 $Y=2.595 $X2=0 $Y2=0
cc_160 N_A1_M1012_g N_VPWR_c_377_n 0.00685982f $X=1.165 $Y=2.595 $X2=0 $Y2=0
cc_161 N_A1_M1012_g N_VPWR_c_379_n 0.00975641f $X=1.165 $Y=2.595 $X2=0 $Y2=0
cc_162 N_A1_M1012_g N_VPWR_c_376_n 0.017165f $X=1.165 $Y=2.595 $X2=0 $Y2=0
cc_163 N_A1_c_165_n N_VGND_c_425_n 0.00421329f $X=1.267 $Y=1.2 $X2=0 $Y2=0
cc_164 A1 N_VGND_c_425_n 0.00693215f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A1_c_168_n N_VGND_c_425_n 0.00103275f $X=1.155 $Y=1.755 $X2=0 $Y2=0
cc_166 N_A1_c_165_n N_VGND_c_429_n 0.00362007f $X=1.267 $Y=1.2 $X2=0 $Y2=0
cc_167 N_A1_c_165_n N_VGND_c_431_n 0.00447875f $X=1.267 $Y=1.2 $X2=0 $Y2=0
cc_168 N_A1_c_165_n N_A_273_141#_c_466_n 0.0131957f $X=1.267 $Y=1.2 $X2=0 $Y2=0
cc_169 N_A1_c_169_n N_A_273_141#_c_466_n 5.49821e-19 $X=1.155 $Y=1.59 $X2=0
+ $Y2=0
cc_170 N_A2_M1003_g N_A3_M1010_g 0.0634372f $X=1.655 $Y=2.595 $X2=0 $Y2=0
cc_171 N_A2_M1002_g N_A3_M1007_g 0.0222435f $X=1.72 $Y=0.915 $X2=0 $Y2=0
cc_172 A2 A3 0.0245445f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_173 N_A2_c_208_n A3 0.00163127f $X=1.695 $Y=1.755 $X2=0 $Y2=0
cc_174 N_A2_M1002_g N_A3_c_246_n 0.00183251f $X=1.72 $Y=0.915 $X2=0 $Y2=0
cc_175 A2 N_A3_c_246_n 6.55032e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_176 N_A2_c_208_n N_A3_c_246_n 0.0207127f $X=1.695 $Y=1.755 $X2=0 $Y2=0
cc_177 A2 N_B1_c_283_n 0.00110615f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A2_M1003_g N_VPWR_c_379_n 0.00975641f $X=1.655 $Y=2.595 $X2=0 $Y2=0
cc_179 N_A2_M1003_g N_VPWR_c_376_n 0.0171404f $X=1.655 $Y=2.595 $X2=0 $Y2=0
cc_180 N_A2_M1002_g N_VGND_c_426_n 0.0053352f $X=1.72 $Y=0.915 $X2=0 $Y2=0
cc_181 N_A2_M1002_g N_VGND_c_429_n 0.00362007f $X=1.72 $Y=0.915 $X2=0 $Y2=0
cc_182 N_A2_M1002_g N_VGND_c_431_n 0.00447875f $X=1.72 $Y=0.915 $X2=0 $Y2=0
cc_183 N_A2_M1002_g N_A_273_141#_c_464_n 0.0117247f $X=1.72 $Y=0.915 $X2=0 $Y2=0
cc_184 A2 N_A_273_141#_c_464_n 0.0135548f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A2_c_208_n N_A_273_141#_c_464_n 4.00036e-19 $X=1.695 $Y=1.755 $X2=0
+ $Y2=0
cc_186 N_A2_M1002_g N_A_273_141#_c_465_n 8.77766e-19 $X=1.72 $Y=0.915 $X2=0
+ $Y2=0
cc_187 N_A2_M1002_g N_A_273_141#_c_466_n 0.010922f $X=1.72 $Y=0.915 $X2=0 $Y2=0
cc_188 A2 N_A_273_141#_c_466_n 0.0117423f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A2_c_208_n N_A_273_141#_c_466_n 7.93511e-19 $X=1.695 $Y=1.755 $X2=0
+ $Y2=0
cc_190 N_A3_M1007_g N_B1_M1008_g 0.0275045f $X=2.31 $Y=0.915 $X2=0 $Y2=0
cc_191 N_A3_c_246_n N_B1_M1008_g 0.00181869f $X=2.235 $Y=1.715 $X2=0 $Y2=0
cc_192 N_A3_M1010_g N_B1_c_282_n 0.0278932f $X=2.195 $Y=2.595 $X2=0 $Y2=0
cc_193 A3 N_B1_c_282_n 2.8802e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A3_c_246_n N_B1_c_282_n 0.0180269f $X=2.235 $Y=1.715 $X2=0 $Y2=0
cc_195 N_A3_M1010_g N_B1_c_283_n 4.37882e-19 $X=2.195 $Y=2.595 $X2=0 $Y2=0
cc_196 A3 N_B1_c_283_n 0.0261249f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A3_c_246_n N_B1_c_283_n 0.002041f $X=2.235 $Y=1.715 $X2=0 $Y2=0
cc_198 N_A3_M1010_g N_VPWR_c_378_n 0.00116955f $X=2.195 $Y=2.595 $X2=0 $Y2=0
cc_199 N_A3_M1010_g N_VPWR_c_379_n 0.00939541f $X=2.195 $Y=2.595 $X2=0 $Y2=0
cc_200 N_A3_M1010_g N_VPWR_c_376_n 0.0163116f $X=2.195 $Y=2.595 $X2=0 $Y2=0
cc_201 N_A3_M1007_g N_VGND_c_426_n 0.00533553f $X=2.31 $Y=0.915 $X2=0 $Y2=0
cc_202 N_A3_M1007_g N_VGND_c_430_n 0.00362548f $X=2.31 $Y=0.915 $X2=0 $Y2=0
cc_203 N_A3_M1007_g N_VGND_c_431_n 0.00447875f $X=2.31 $Y=0.915 $X2=0 $Y2=0
cc_204 N_A3_M1007_g N_A_273_141#_c_464_n 0.0152876f $X=2.31 $Y=0.915 $X2=0 $Y2=0
cc_205 A3 N_A_273_141#_c_464_n 0.0222762f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_206 N_A3_c_246_n N_A_273_141#_c_464_n 0.00497414f $X=2.235 $Y=1.715 $X2=0
+ $Y2=0
cc_207 N_A3_M1007_g N_A_273_141#_c_465_n 0.00912377f $X=2.31 $Y=0.915 $X2=0
+ $Y2=0
cc_208 N_A3_M1007_g N_A_273_141#_c_466_n 8.82758e-19 $X=2.31 $Y=0.915 $X2=0
+ $Y2=0
cc_209 N_B1_M1008_g N_C1_c_318_n 0.0468515f $X=2.74 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_210 N_B1_M1000_g N_C1_M1005_g 0.0415946f $X=2.735 $Y=2.595 $X2=0 $Y2=0
cc_211 N_B1_c_282_n N_C1_c_320_n 0.0204348f $X=2.775 $Y=1.755 $X2=0 $Y2=0
cc_212 N_B1_c_283_n N_C1_c_320_n 2.8686e-19 $X=2.775 $Y=1.755 $X2=0 $Y2=0
cc_213 N_B1_c_282_n N_C1_c_321_n 0.00220756f $X=2.775 $Y=1.755 $X2=0 $Y2=0
cc_214 N_B1_c_283_n N_C1_c_321_n 0.0298996f $X=2.775 $Y=1.755 $X2=0 $Y2=0
cc_215 N_B1_M1008_g N_C1_c_322_n 0.00991548f $X=2.74 $Y=0.915 $X2=0 $Y2=0
cc_216 N_B1_M1000_g N_VPWR_c_378_n 0.0196534f $X=2.735 $Y=2.595 $X2=0 $Y2=0
cc_217 N_B1_M1000_g N_VPWR_c_379_n 0.00855241f $X=2.735 $Y=2.595 $X2=0 $Y2=0
cc_218 N_B1_M1000_g N_VPWR_c_376_n 0.013998f $X=2.735 $Y=2.595 $X2=0 $Y2=0
cc_219 N_B1_M1008_g N_VGND_c_430_n 0.00362548f $X=2.74 $Y=0.915 $X2=0 $Y2=0
cc_220 N_B1_M1008_g N_VGND_c_431_n 0.00447875f $X=2.74 $Y=0.915 $X2=0 $Y2=0
cc_221 N_B1_M1008_g N_A_273_141#_c_464_n 0.00557684f $X=2.74 $Y=0.915 $X2=0
+ $Y2=0
cc_222 N_B1_c_282_n N_A_273_141#_c_464_n 3.83651e-19 $X=2.775 $Y=1.755 $X2=0
+ $Y2=0
cc_223 N_B1_c_283_n N_A_273_141#_c_464_n 0.013491f $X=2.775 $Y=1.755 $X2=0 $Y2=0
cc_224 N_B1_M1008_g N_A_273_141#_c_465_n 0.0103136f $X=2.74 $Y=0.915 $X2=0 $Y2=0
cc_225 N_C1_M1005_g N_VPWR_c_378_n 0.0185319f $X=3.275 $Y=2.595 $X2=0 $Y2=0
cc_226 N_C1_M1005_g N_VPWR_c_381_n 0.00915325f $X=3.275 $Y=2.595 $X2=0 $Y2=0
cc_227 N_C1_M1005_g N_VPWR_c_376_n 0.0160116f $X=3.275 $Y=2.595 $X2=0 $Y2=0
cc_228 N_C1_c_318_n N_VGND_c_430_n 0.00362453f $X=3.1 $Y=1.2 $X2=0 $Y2=0
cc_229 N_C1_c_318_n N_VGND_c_431_n 0.00447875f $X=3.1 $Y=1.2 $X2=0 $Y2=0
cc_230 N_C1_c_319_n N_A_273_141#_c_464_n 7.86571e-19 $X=3.225 $Y=1.275 $X2=0
+ $Y2=0
cc_231 N_C1_c_318_n N_A_273_141#_c_465_n 0.00182516f $X=3.1 $Y=1.2 $X2=0 $Y2=0
cc_232 N_X_c_357_n N_VPWR_c_377_n 0.0407944f $X=0.295 $Y=2.28 $X2=0 $Y2=0
cc_233 N_X_M1009_s N_VPWR_c_376_n 0.0023218f $X=0.15 $Y=2.095 $X2=0 $Y2=0
cc_234 N_X_c_357_n N_VPWR_c_376_n 0.0136688f $X=0.295 $Y=2.28 $X2=0 $Y2=0
cc_235 N_X_c_357_n N_VPWR_c_383_n 0.0217808f $X=0.295 $Y=2.28 $X2=0 $Y2=0
cc_236 X N_VGND_c_425_n 0.0223022f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_237 X N_VGND_c_427_n 0.0111942f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_238 X N_VGND_c_431_n 0.0119466f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_239 N_VPWR_c_376_n A_258_419# 0.010279f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_240 N_VPWR_c_376_n A_356_419# 0.0124205f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_241 N_VGND_c_426_n N_A_273_141#_c_464_n 0.0259275f $X=2.015 $Y=0.85 $X2=0
+ $Y2=0
cc_242 N_VGND_c_426_n N_A_273_141#_c_465_n 0.0127661f $X=2.015 $Y=0.85 $X2=0
+ $Y2=0
cc_243 N_VGND_c_430_n N_A_273_141#_c_465_n 0.00590248f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_244 N_VGND_c_431_n N_A_273_141#_c_465_n 0.00953571f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_245 N_VGND_c_425_n N_A_273_141#_c_466_n 0.0286387f $X=1.07 $Y=0.885 $X2=0
+ $Y2=0
cc_246 N_VGND_c_426_n N_A_273_141#_c_466_n 0.0128339f $X=2.015 $Y=0.85 $X2=0
+ $Y2=0
cc_247 N_VGND_c_429_n N_A_273_141#_c_466_n 0.00584742f $X=1.85 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_c_431_n N_A_273_141#_c_466_n 0.00950558f $X=3.6 $Y=0 $X2=0 $Y2=0
