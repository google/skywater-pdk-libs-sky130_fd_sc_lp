* File: sky130_fd_sc_lp__nand3b_2.pex.spice
* Created: Wed Sep  2 10:04:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3B_2%A_N 3 7 9 12
r31 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.51
+ $X2=0.525 $Y2=1.675
r32 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.51
+ $X2=0.525 $Y2=1.345
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.51 $X2=0.525 $Y2=1.51
r34 9 13 5.5488 $w=4.03e-07 $l=1.95e-07 $layer=LI1_cond $X=0.72 $Y=1.547
+ $X2=0.525 $Y2=1.547
r35 7 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.615 $Y=2.045
+ $X2=0.615 $Y2=1.675
r36 3 14 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=0.615 $Y=0.985
+ $X2=0.615 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_2%C 3 7 11 15 17 18 21 22 24 25 29 42
c97 17 0 1.97015e-19 $X=3.54 $Y=2.16
c98 7 0 1.78576e-19 $X=1.175 $Y=2.465
r99 29 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.51
+ $X2=1.085 $Y2=1.675
r100 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.51
+ $X2=1.085 $Y2=1.345
r101 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.51 $X2=1.085 $Y2=1.51
r102 25 42 2.13415 $w=4.03e-07 $l=7.5e-08 $layer=LI1_cond $X=1.2 $Y=1.547
+ $X2=1.275 $Y2=1.547
r103 25 42 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=1.275 $Y=1.75
+ $X2=1.275 $Y2=1.547
r104 25 30 3.27237 $w=4.03e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.547
+ $X2=1.085 $Y2=1.547
r105 24 25 15.3752 $w=2.63e-07 $l=3.25e-07 $layer=LI1_cond $X=1.275 $Y=2.075
+ $X2=1.275 $Y2=1.75
r106 22 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.51
+ $X2=3.705 $Y2=1.675
r107 22 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.51
+ $X2=3.705 $Y2=1.345
r108 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.51 $X2=3.705 $Y2=1.51
r109 19 21 26.0452 $w=2.48e-07 $l=5.65e-07 $layer=LI1_cond $X=3.665 $Y=2.075
+ $X2=3.665 $Y2=1.51
r110 18 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.36 $Y=2.16
+ $X2=1.275 $Y2=2.075
r111 17 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.54 $Y=2.16
+ $X2=3.665 $Y2=2.075
r112 17 18 142.225 $w=1.68e-07 $l=2.18e-06 $layer=LI1_cond $X=3.54 $Y=2.16
+ $X2=1.36 $Y2=2.16
r113 15 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.615 $Y=2.465
+ $X2=3.615 $Y2=1.675
r114 11 34 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.615 $Y=0.775
+ $X2=3.615 $Y2=1.345
r115 7 32 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.175 $Y=2.465
+ $X2=1.175 $Y2=1.675
r116 3 31 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.155 $Y=0.775
+ $X2=1.155 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_2%B 3 7 11 15 19 20 23 24 25 32 33 37
c93 32 0 8.31604e-20 $X=3.165 $Y=1.51
c94 23 0 1.78576e-19 $X=1.72 $Y=1.82
r95 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.51
+ $X2=3.165 $Y2=1.675
r96 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.51
+ $X2=3.165 $Y2=1.345
r97 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.165
+ $Y=1.51 $X2=3.165 $Y2=1.51
r98 25 33 0.961134 $w=5.58e-07 $l=4.5e-08 $layer=LI1_cond $X=3.12 $Y=1.625
+ $X2=3.165 $Y2=1.625
r99 24 25 10.2521 $w=5.58e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.625
+ $X2=3.12 $Y2=1.625
r100 24 37 8.93522 $w=5.58e-07 $l=1.2e-07 $layer=LI1_cond $X=2.64 $Y=1.625
+ $X2=2.52 $Y2=1.625
r101 23 37 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.72 $Y=1.82 $X2=2.52
+ $Y2=1.82
r102 20 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=1.51
+ $X2=1.625 $Y2=1.675
r103 20 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=1.51
+ $X2=1.625 $Y2=1.345
r104 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.51 $X2=1.625 $Y2=1.51
r105 17 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.625 $Y=1.735
+ $X2=1.72 $Y2=1.82
r106 17 19 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=1.625 $Y=1.735
+ $X2=1.625 $Y2=1.51
r107 15 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.185 $Y=2.465
+ $X2=3.185 $Y2=1.675
r108 11 34 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.145 $Y=0.775
+ $X2=3.145 $Y2=1.345
r109 7 30 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.605 $Y=2.465
+ $X2=1.605 $Y2=1.675
r110 3 29 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.585 $Y=0.775
+ $X2=1.585 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_2%A_55_155# 1 2 7 9 12 16 18 20 22 23 26 27
+ 29 36 40 45
c97 45 0 1.97015e-19 $X=2.625 $Y=1.47
c98 29 0 8.31604e-20 $X=2.185 $Y=1.47
r99 44 45 67.2922 $w=3.08e-07 $l=4.3e-07 $layer=POLY_cond $X=2.195 $Y=1.47
+ $X2=2.625 $Y2=1.47
r100 37 40 9.2607 $w=2.78e-07 $l=2.25e-07 $layer=LI1_cond $X=0.175 $Y=2.06
+ $X2=0.4 $Y2=2.06
r101 35 36 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.4 $Y=1 $X2=0.565
+ $Y2=1
r102 32 35 7.40856 $w=3.48e-07 $l=2.25e-07 $layer=LI1_cond $X=0.175 $Y=1 $X2=0.4
+ $Y2=1
r103 30 44 1.56494 $w=3.08e-07 $l=1e-08 $layer=POLY_cond $X=2.185 $Y=1.47
+ $X2=2.195 $Y2=1.47
r104 30 42 14.0844 $w=3.08e-07 $l=9e-08 $layer=POLY_cond $X=2.185 $Y=1.47
+ $X2=2.095 $Y2=1.47
r105 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.185
+ $Y=1.47 $X2=2.185 $Y2=1.47
r106 27 29 6.54797 $w=2.18e-07 $l=1.25e-07 $layer=LI1_cond $X=2.06 $Y=1.455
+ $X2=2.185 $Y2=1.455
r107 26 27 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.975 $Y=1.345
+ $X2=2.06 $Y2=1.455
r108 25 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.975 $Y=1.175
+ $X2=1.975 $Y2=1.345
r109 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.89 $Y=1.09
+ $X2=1.975 $Y2=1.175
r110 23 36 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=1.89 $Y=1.09
+ $X2=0.565 $Y2=1.09
r111 22 37 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.175 $Y=1.92
+ $X2=0.175 $Y2=2.06
r112 21 32 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.175 $Y=1.175
+ $X2=0.175 $Y2=1
r113 21 22 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.175 $Y=1.175
+ $X2=0.175 $Y2=1.92
r114 18 45 14.0844 $w=3.08e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.715 $Y=1.305
+ $X2=2.625 $Y2=1.47
r115 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.715 $Y=1.305
+ $X2=2.715 $Y2=0.775
r116 14 45 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.635
+ $X2=2.625 $Y2=1.47
r117 14 16 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.625 $Y=1.635
+ $X2=2.625 $Y2=2.465
r118 10 44 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.635
+ $X2=2.195 $Y2=1.47
r119 10 12 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.195 $Y=1.635
+ $X2=2.195 $Y2=2.465
r120 7 42 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.305
+ $X2=2.095 $Y2=1.47
r121 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.095 $Y=1.305
+ $X2=2.095 $Y2=0.775
r122 2 40 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.835 $X2=0.4 $Y2=2.035
r123 1 35 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.775 $X2=0.4 $Y2=0.99
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_2%VPWR 1 2 3 4 15 21 25 29 32 33 35 36 38 39
+ 41 42 43 59 60
r72 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 57 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r74 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r75 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r76 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r77 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r78 47 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 43 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r82 41 56 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.735 $Y=3.33
+ $X2=3.6 $Y2=3.33
r83 41 42 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.735 $Y=3.33
+ $X2=3.865 $Y2=3.33
r84 40 59 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=3.33
+ $X2=4.08 $Y2=3.33
r85 40 42 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.995 $Y=3.33
+ $X2=3.865 $Y2=3.33
r86 38 53 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 38 39 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.905 $Y2=3.33
r88 37 56 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=3.6 $Y2=3.33
r89 37 39 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=2.905 $Y2=3.33
r90 35 50 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.9 $Y2=3.33
r92 34 53 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.64 $Y2=3.33
r93 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.9 $Y2=3.33
r94 32 46 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 32 33 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.877 $Y2=3.33
r96 31 50 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.02 $Y=3.33
+ $X2=1.68 $Y2=3.33
r97 31 33 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.02 $Y=3.33
+ $X2=0.877 $Y2=3.33
r98 27 42 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=3.245
+ $X2=3.865 $Y2=3.33
r99 27 29 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=3.865 $Y=3.245
+ $X2=3.865 $Y2=2.92
r100 23 39 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=3.33
r101 23 25 11.7045 $w=3.18e-07 $l=3.25e-07 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=2.92
r102 19 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.9 $Y=3.245 $X2=1.9
+ $Y2=3.33
r103 19 21 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.9 $Y=3.245
+ $X2=1.9 $Y2=2.92
r104 15 18 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=0.877 $Y=2.085
+ $X2=0.877 $Y2=2.515
r105 13 33 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.877 $Y=3.245
+ $X2=0.877 $Y2=3.33
r106 13 18 29.5187 $w=2.83e-07 $l=7.3e-07 $layer=LI1_cond $X=0.877 $Y=3.245
+ $X2=0.877 $Y2=2.515
r107 4 29 600 $w=1.7e-07 $l=1.15288e-06 $layer=licon1_PDIFF $count=1 $X=3.69
+ $Y=1.835 $X2=3.83 $Y2=2.92
r108 3 25 600 $w=1.7e-07 $l=1.18307e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.905 $Y2=2.92
r109 2 21 600 $w=1.7e-07 $l=1.18993e-06 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.835 $X2=1.9 $Y2=2.92
r110 1 18 300 $w=1.7e-07 $l=7.88797e-07 $layer=licon1_PDIFF $count=2 $X=0.69
+ $Y=1.835 $X2=0.925 $Y2=2.515
r111 1 15 600 $w=1.7e-07 $l=3.29773e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.835 $X2=0.875 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_2%Y 1 2 3 4 15 19 21 25 28 32 34 36 38 39 40
+ 41 47 56
c89 25 0 2.4855e-20 $X=3.96 $Y=2.5
r90 47 56 0.41907 $w=2.73e-07 $l=1e-08 $layer=LI1_cond $X=4.097 $Y=2.415
+ $X2=4.097 $Y2=2.405
r91 41 47 2.80348 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.097 $Y=2.5
+ $X2=4.097 $Y2=2.415
r92 41 56 1.59247 $w=2.73e-07 $l=3.8e-08 $layer=LI1_cond $X=4.097 $Y=2.367
+ $X2=4.097 $Y2=2.405
r93 40 41 13.9131 $w=2.73e-07 $l=3.32e-07 $layer=LI1_cond $X=4.097 $Y=2.035
+ $X2=4.097 $Y2=2.367
r94 39 40 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=4.097 $Y=1.665
+ $X2=4.097 $Y2=2.035
r95 38 39 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=4.097 $Y=1.295
+ $X2=4.097 $Y2=1.665
r96 37 38 5.02884 $w=2.73e-07 $l=1.2e-07 $layer=LI1_cond $X=4.097 $Y=1.175
+ $X2=4.097 $Y2=1.295
r97 30 32 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=1.055
+ $X2=2.57 $Y2=1.055
r98 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.565 $Y=2.5 $X2=3.4
+ $Y2=2.5
r99 25 41 4.51856 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=3.96 $Y=2.5
+ $X2=4.097 $Y2=2.5
r100 25 26 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.96 $Y=2.5
+ $X2=3.565 $Y2=2.5
r101 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=2.5
+ $X2=2.41 $Y2=2.5
r102 21 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=2.5
+ $X2=3.4 $Y2=2.5
r103 21 22 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.235 $Y=2.5
+ $X2=2.575 $Y2=2.5
r104 19 37 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=3.96 $Y=1.09
+ $X2=4.097 $Y2=1.175
r105 19 32 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=3.96 $Y=1.09
+ $X2=2.57 $Y2=1.09
r106 16 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=2.5
+ $X2=1.39 $Y2=2.5
r107 15 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=2.5
+ $X2=2.41 $Y2=2.5
r108 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.245 $Y=2.5
+ $X2=1.555 $Y2=2.5
r109 4 36 300 $w=1.7e-07 $l=7.31659e-07 $layer=licon1_PDIFF $count=2 $X=3.26
+ $Y=1.835 $X2=3.4 $Y2=2.5
r110 3 34 300 $w=1.7e-07 $l=7.31659e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.5
r111 2 28 300 $w=1.7e-07 $l=7.31659e-07 $layer=licon1_PDIFF $count=2 $X=1.25
+ $Y=1.835 $X2=1.39 $Y2=2.5
r112 1 30 182 $w=1.7e-07 $l=8.03959e-07 $layer=licon1_NDIFF $count=1 $X=2.17
+ $Y=0.355 $X2=2.405 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_2%VGND 1 2 9 13 16 17 19 20 21 34 35
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r40 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r41 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r42 28 31 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r43 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r45 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 21 32 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r47 21 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r48 19 31 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.6
+ $Y2=0
r49 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.83
+ $Y2=0
r50 18 34 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=0 $X2=4.08
+ $Y2=0
r51 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.83
+ $Y2=0
r52 16 24 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.72
+ $Y2=0
r53 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.94
+ $Y2=0
r54 15 28 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.105 $Y=0 $X2=1.2
+ $Y2=0
r55 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=0.94
+ $Y2=0
r56 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0
r57 11 13 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0.72
r58 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.94 $Y=0.085 $X2=0.94
+ $Y2=0
r59 7 9 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=0.94 $Y=0.085 $X2=0.94
+ $Y2=0.705
r60 2 13 182 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=1 $X=3.69
+ $Y=0.355 $X2=3.83 $Y2=0.72
r61 1 9 182 $w=1.7e-07 $l=2.82843e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.775 $X2=0.94 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_2%A_246_71# 1 2 9 11 12 15
r27 13 15 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.38 $Y=0.425
+ $X2=3.38 $Y2=0.67
r28 11 13 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.265 $Y=0.34
+ $X2=3.38 $Y2=0.425
r29 11 12 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=3.265 $Y=0.34
+ $X2=1.535 $Y2=0.34
r30 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.405 $Y=0.425
+ $X2=1.535 $Y2=0.34
r31 7 9 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=1.405 $Y=0.425
+ $X2=1.405 $Y2=0.67
r32 2 15 182 $w=1.7e-07 $l=3.86814e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.355 $X2=3.38 $Y2=0.67
r33 1 9 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=1.23
+ $Y=0.355 $X2=1.37 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3B_2%A_332_71# 1 2 12 14 15
r20 14 15 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=0.715
+ $X2=2.765 $Y2=0.715
r21 12 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.035 $Y=0.68
+ $X2=2.765 $Y2=0.68
r22 10 12 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=0.715
+ $X2=2.035 $Y2=0.715
r23 2 14 182 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.355 $X2=2.93 $Y2=0.72
r24 1 10 182 $w=1.7e-07 $l=4.47856e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.355 $X2=1.87 $Y2=0.71
.ends

