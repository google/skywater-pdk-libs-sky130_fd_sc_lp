* File: sky130_fd_sc_lp__ebufn_1.pex.spice
* Created: Fri Aug 28 10:31:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EBUFN_1%A_105_263# 1 2 9 13 14 17 18 19 21 22 23 27
+ 30 32 34 37 39
c90 32 0 2.69861e-19 $X=0.855 $Y=1.48
r91 30 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.69 $Y=1.48
+ $X2=0.69 $Y2=1.645
r92 30 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.69 $Y=1.48
+ $X2=0.69 $Y2=1.315
r93 29 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.48
+ $X2=0.855 $Y2=1.48
r94 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.69
+ $Y=1.48 $X2=0.69 $Y2=1.48
r95 27 37 2.99104 $w=3.17e-07 $l=1.85699e-07 $layer=LI1_cond $X=3.67 $Y=2.11
+ $X2=3.522 $Y2=2.195
r96 26 34 9.10704 $w=3.55e-07 $l=3.62181e-07 $layer=LI1_cond $X=3.67 $Y=1.1
+ $X2=3.405 $Y2=0.87
r97 26 27 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.67 $Y=1.1
+ $X2=3.67 $Y2=2.11
r98 22 37 3.66292 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.29 $Y=2.195
+ $X2=3.522 $Y2=2.195
r99 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.29 $Y=2.195
+ $X2=2.62 $Y2=2.195
r100 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.535 $Y=2.28
+ $X2=2.62 $Y2=2.195
r101 20 21 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.535 $Y=2.28
+ $X2=2.535 $Y2=2.905
r102 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.45 $Y=2.99
+ $X2=2.535 $Y2=2.905
r103 18 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.45 $Y=2.99
+ $X2=1.86 $Y2=2.99
r104 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.775 $Y=2.905
+ $X2=1.86 $Y2=2.99
r105 16 17 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=1.775 $Y=1.625
+ $X2=1.775 $Y2=2.905
r106 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.69 $Y=1.54
+ $X2=1.775 $Y2=1.625
r107 14 32 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.69 $Y=1.54
+ $X2=0.855 $Y2=1.54
r108 13 39 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.78 $Y=0.785
+ $X2=0.78 $Y2=1.315
r109 9 40 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.75 $Y=2.465
+ $X2=0.75 $Y2=1.645
r110 2 37 300 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=2 $X=3.265
+ $Y=2.13 $X2=3.455 $Y2=2.275
r111 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=0.66 $X2=3.405 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_1%A_219_21# 1 2 7 9 10 11 12 14 21
c40 7 0 1.23395e-19 $X=1.17 $Y=0.255
r41 18 21 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.985 $Y=0.42
+ $X2=1.985 $Y2=0.18
r42 17 20 12.1192 $w=4.53e-07 $l=4.5e-07 $layer=LI1_cond $X=2.195 $Y=0.42
+ $X2=2.195 $Y2=0.87
r43 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.985
+ $Y=0.42 $X2=1.985 $Y2=0.42
r44 12 20 8.62573 $w=4.53e-07 $l=2.49199e-07 $layer=LI1_cond $X=2.155 $Y=1.1
+ $X2=2.195 $Y2=0.87
r45 12 14 60.849 $w=2.48e-07 $l=1.32e-06 $layer=LI1_cond $X=2.155 $Y=1.1
+ $X2=2.155 $Y2=2.42
r46 10 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=0.18
+ $X2=1.985 $Y2=0.18
r47 10 11 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.82 $Y=0.18
+ $X2=1.245 $Y2=0.18
r48 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.17 $Y=0.255
+ $X2=1.245 $Y2=0.18
r49 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.17 $Y=0.255 $X2=1.17
+ $Y2=0.785
r50 2 14 600 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=2.13 $X2=2.115 $Y2=2.42
r51 1 20 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.26
+ $Y=0.66 $X2=2.405 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_1%TE_B 3 5 6 9 13 15 18 19
c54 6 0 1.46466e-19 $X=1.215 $Y=1.63
r55 21 22 62.5979 $w=6.2e-07 $l=3.1e-07 $layer=POLY_cond $X=2.565 $Y=1.63
+ $X2=2.565 $Y2=1.94
r56 18 21 16.8275 $w=6.2e-07 $l=1.95e-07 $layer=POLY_cond $X=2.565 $Y=1.435
+ $X2=2.565 $Y2=1.63
r57 18 20 50.0851 $w=6.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.565 $Y=1.435
+ $X2=2.565 $Y2=1.27
r58 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.615
+ $Y=1.435 $X2=2.615 $Y2=1.435
r59 15 19 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.615 $Y=1.665
+ $X2=2.615 $Y2=1.435
r60 13 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.62 $Y=0.87 $X2=2.62
+ $Y2=1.27
r61 9 22 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.33 $Y=2.45 $X2=2.33
+ $Y2=1.94
r62 5 21 36.9266 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=2.255 $Y=1.63
+ $X2=2.565 $Y2=1.63
r63 5 6 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.255 $Y=1.63
+ $X2=1.215 $Y2=1.63
r64 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.14 $Y=1.705
+ $X2=1.215 $Y2=1.63
r65 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.14 $Y=1.705 $X2=1.14
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_1%A 3 7 11 12 13 16 17
r35 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.25
+ $Y=1.435 $X2=3.25 $Y2=1.435
r36 13 17 2.32075 $w=6.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=3.25 $Y2=1.605
r37 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.25 $Y=1.775
+ $X2=3.25 $Y2=1.435
r38 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.775
+ $X2=3.25 $Y2=1.94
r39 10 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.27
+ $X2=3.25 $Y2=1.435
r40 7 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.19 $Y=2.45 $X2=3.19
+ $Y2=1.94
r41 3 10 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.19 $Y=0.87 $X2=3.19
+ $Y2=1.27
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_1%Z 1 2 7 8 9 10 11 12 13 38 46 50
r25 46 47 8.29682 $w=5.73e-07 $l=1.85e-07 $layer=LI1_cond $X=0.412 $Y=2
+ $X2=0.412 $Y2=1.815
r26 28 50 1.39369 $w=5.73e-07 $l=6.7e-08 $layer=LI1_cond $X=0.412 $Y=2.102
+ $X2=0.412 $Y2=2.035
r27 13 35 3.22421 $w=5.73e-07 $l=1.55e-07 $layer=LI1_cond $X=0.412 $Y=2.775
+ $X2=0.412 $Y2=2.93
r28 12 13 7.6965 $w=5.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.412 $Y=2.405
+ $X2=0.412 $Y2=2.775
r29 11 50 0.187212 $w=5.73e-07 $l=9e-09 $layer=LI1_cond $X=0.412 $Y=2.026
+ $X2=0.412 $Y2=2.035
r30 11 46 0.540835 $w=5.73e-07 $l=2.6e-08 $layer=LI1_cond $X=0.412 $Y=2.026
+ $X2=0.412 $Y2=2
r31 11 12 6.1156 $w=5.73e-07 $l=2.94e-07 $layer=LI1_cond $X=0.412 $Y=2.111
+ $X2=0.412 $Y2=2.405
r32 11 28 0.187212 $w=5.73e-07 $l=9e-09 $layer=LI1_cond $X=0.412 $Y=2.111
+ $X2=0.412 $Y2=2.102
r33 10 47 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.815
r34 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r35 9 44 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.145
r36 8 44 9.14464 $w=6.03e-07 $l=2.2e-07 $layer=LI1_cond $X=0.427 $Y=0.925
+ $X2=0.427 $Y2=1.145
r37 7 8 7.31486 $w=6.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.427 $Y=0.555
+ $X2=0.427 $Y2=0.925
r38 7 38 0.889645 $w=6.03e-07 $l=4.5e-08 $layer=LI1_cond $X=0.427 $Y=0.555
+ $X2=0.427 $Y2=0.51
r39 2 46 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=0.39
+ $Y=1.835 $X2=0.535 $Y2=2
r40 2 35 400 $w=1.7e-07 $l=1.16525e-06 $layer=licon1_PDIFF $count=1 $X=0.39
+ $Y=1.835 $X2=0.535 $Y2=2.93
r41 1 38 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.42
+ $Y=0.365 $X2=0.565 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r40 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r41 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r42 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r43 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r46 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=3.33
+ $X2=1.355 $Y2=3.33
r48 27 29 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.52 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 25 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.19 $Y=3.33
+ $X2=1.355 $Y2=3.33
r52 22 24 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=1.19 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 20 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 20 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 18 32 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=3.33 $X2=2.64
+ $Y2=3.33
r56 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=3.33
+ $X2=2.955 $Y2=3.33
r57 17 35 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=2.955 $Y2=3.33
r59 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=2.955 $Y2=3.33
r60 13 15 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=2.955 $Y2=2.62
r61 9 12 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=1.355 $Y=1.98
+ $X2=1.355 $Y2=2.95
r62 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=3.33
r63 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=2.95
r64 2 15 600 $w=1.7e-07 $l=7.56307e-07 $layer=licon1_PDIFF $count=1 $X=2.405
+ $Y=2.13 $X2=2.955 $Y2=2.62
r65 1 12 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=1.835 $X2=1.355 $Y2=2.95
r66 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=1.835 $X2=1.355 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_1%VGND 1 2 9 13 16 17 19 20 21 37 38
r43 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r45 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r47 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r48 29 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r49 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r51 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r52 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 21 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r54 21 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r55 19 34 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.64
+ $Y2=0
r56 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.905
+ $Y2=0
r57 18 37 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=3.6
+ $Y2=0
r58 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=2.905
+ $Y2=0
r59 16 28 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.2
+ $Y2=0
r60 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.385
+ $Y2=0
r61 15 31 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=1.68
+ $Y2=0
r62 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=1.385
+ $Y2=0
r63 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=0.085
+ $X2=2.905 $Y2=0
r64 11 13 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=2.905 $Y=0.085
+ $X2=2.905 $Y2=0.87
r65 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=0.085
+ $X2=1.385 $Y2=0
r66 7 9 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.385 $Y=0.085
+ $X2=1.385 $Y2=0.51
r67 2 13 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.66 $X2=2.905 $Y2=0.87
r68 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.245
+ $Y=0.365 $X2=1.385 $Y2=0.51
.ends

