* File: sky130_fd_sc_lp__nor4bb_1.pex.spice
* Created: Wed Sep  2 10:11:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4BB_1%D_N 3 7 9 10 11 16
c33 9 0 1.68009e-19 $X=0.24 $Y=1.295
c34 7 0 1.39738e-19 $X=0.81 $Y=0.865
r35 16 19 83.6195 $w=4.85e-07 $l=5.05e-07 $layer=POLY_cond $X=0.642 $Y=1.375
+ $X2=0.642 $Y2=1.88
r36 16 18 46.1122 $w=4.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.642 $Y=1.375
+ $X2=0.642 $Y2=1.21
r37 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.565
+ $Y=1.375 $X2=0.565 $Y2=1.375
r38 10 11 7.83273 $w=5.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.367 $Y=1.665
+ $X2=0.367 $Y2=2.035
r39 10 17 6.13916 $w=5.63e-07 $l=2.9e-07 $layer=LI1_cond $X=0.367 $Y=1.665
+ $X2=0.367 $Y2=1.375
r40 9 17 1.69356 $w=5.63e-07 $l=8e-08 $layer=LI1_cond $X=0.367 $Y=1.295
+ $X2=0.367 $Y2=1.375
r41 7 18 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.81 $Y=0.865
+ $X2=0.81 $Y2=1.21
r42 3 19 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=0.475 $Y=2.75
+ $X2=0.475 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_1%A_27_508# 1 2 7 9 10 12 15 17 18 19 24 26
+ 31
c61 31 0 5.10176e-20 $X=1.26 $Y=1.35
c62 10 0 1.68009e-19 $X=1.59 $Y=1.725
r63 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.26
+ $Y=1.35 $X2=1.26 $Y2=1.35
r64 29 31 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.925 $Y=1.35
+ $X2=1.26 $Y2=1.35
r65 27 29 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=0.905 $Y=1.35
+ $X2=0.925 $Y2=1.35
r66 25 29 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=1.515
+ $X2=0.925 $Y2=1.35
r67 25 26 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=0.925 $Y=1.515
+ $X2=0.925 $Y2=2.29
r68 24 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=1.35
r69 23 24 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.905 $Y=1.035
+ $X2=0.905 $Y2=1.185
r70 19 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.82 $Y=0.87
+ $X2=0.905 $Y2=1.035
r71 19 21 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.82 $Y=0.87
+ $X2=0.595 $Y2=0.87
r72 17 26 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.82 $Y=2.375
+ $X2=0.925 $Y2=2.29
r73 17 18 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.82 $Y=2.375
+ $X2=0.355 $Y2=2.375
r74 13 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=2.46
+ $X2=0.355 $Y2=2.375
r75 13 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=2.46
+ $X2=0.225 $Y2=2.755
r76 10 32 62.1696 $w=5e-07 $l=4.68375e-07 $layer=POLY_cond $X=1.59 $Y=1.725
+ $X2=1.38 $Y2=1.35
r77 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.59 $Y=1.725
+ $X2=1.59 $Y2=2.465
r78 7 32 41.9256 $w=5e-07 $l=2.80624e-07 $layer=POLY_cond $X=1.59 $Y=1.185
+ $X2=1.38 $Y2=1.35
r79 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.59 $Y=1.185 $X2=1.59
+ $Y2=0.655
r80 2 15 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.26 $Y2=2.755
r81 1 21 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.47
+ $Y=0.655 $X2=0.595 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_1%A_375_269# 1 2 9 13 17 18 20 21 23 24 25 28
+ 32 34
c77 13 0 5.10176e-20 $X=2.02 $Y=0.655
c78 9 0 8.35911e-20 $X=1.95 $Y=2.465
r79 30 32 10.8042 $w=2.38e-07 $l=2.25e-07 $layer=LI1_cond $X=4.04 $Y=1.085
+ $X2=4.04 $Y2=0.86
r80 26 34 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=2.037
+ $X2=3.47 $Y2=2.037
r81 26 28 12.3285 $w=2.13e-07 $l=2.3e-07 $layer=LI1_cond $X=3.555 $Y=2.037
+ $X2=3.785 $Y2=2.037
r82 24 30 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.92 $Y=1.17
+ $X2=4.04 $Y2=1.085
r83 24 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.92 $Y=1.17
+ $X2=3.555 $Y2=1.17
r84 23 34 2.20034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=3.47 $Y=1.93
+ $X2=3.47 $Y2=2.037
r85 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=1.255
+ $X2=3.555 $Y2=1.17
r86 22 23 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.47 $Y=1.255
+ $X2=3.47 $Y2=1.93
r87 20 34 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=2.037
+ $X2=3.47 $Y2=2.037
r88 20 21 63.2504 $w=2.13e-07 $l=1.18e-06 $layer=LI1_cond $X=3.385 $Y=2.037
+ $X2=2.205 $Y2=2.037
r89 18 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.51
+ $X2=2.04 $Y2=1.675
r90 18 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.51
+ $X2=2.04 $Y2=1.345
r91 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.04
+ $Y=1.51 $X2=2.04 $Y2=1.51
r92 15 21 7.21882 $w=2.15e-07 $l=2.11849e-07 $layer=LI1_cond $X=2.04 $Y=1.93
+ $X2=2.205 $Y2=2.037
r93 15 17 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.04 $Y=1.93
+ $X2=2.04 $Y2=1.51
r94 13 36 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.02 $Y=0.655
+ $X2=2.02 $Y2=1.345
r95 9 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.95 $Y=2.465
+ $X2=1.95 $Y2=1.675
r96 2 28 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=3.645
+ $Y=1.835 $X2=3.785 $Y2=2.035
r97 1 32 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.655 $X2=4.015 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_1%B 3 7 9 12 13
c34 13 0 8.35911e-20 $X=2.58 $Y=1.51
c35 7 0 5.03048e-20 $X=2.555 $Y=0.655
c36 3 0 7.80666e-20 $X=2.49 $Y=2.465
r37 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.51
+ $X2=2.58 $Y2=1.675
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.51
+ $X2=2.58 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.51 $X2=2.58 $Y2=1.51
r40 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.58 $Y=1.665
+ $X2=2.58 $Y2=1.51
r41 7 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.555 $Y=0.655
+ $X2=2.555 $Y2=1.345
r42 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.49 $Y=2.465
+ $X2=2.49 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_1%A 3 6 8 9 13 15
c39 8 0 7.80666e-20 $X=3.12 $Y=1.295
r40 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.35
+ $X2=3.12 $Y2=1.515
r41 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.35
+ $X2=3.12 $Y2=1.185
r42 8 9 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.295 $X2=3.12
+ $Y2=1.665
r43 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.35 $X2=3.12 $Y2=1.35
r44 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.03 $Y=2.465
+ $X2=3.03 $Y2=1.515
r45 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.03 $Y=0.655
+ $X2=3.03 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_1%C_N 3 7 9 12
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.9
+ $Y=1.51 $X2=3.9 $Y2=1.51
r29 12 14 18.7549 $w=2.57e-07 $l=1e-07 $layer=POLY_cond $X=3.8 $Y=1.51 $X2=3.9
+ $Y2=1.51
r30 9 15 6.19223 $w=3.33e-07 $l=1.8e-07 $layer=LI1_cond $X=4.08 $Y=1.592 $X2=3.9
+ $Y2=1.592
r31 5 12 15.359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.8 $Y=1.345 $X2=3.8
+ $Y2=1.51
r32 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.8 $Y=1.345 $X2=3.8
+ $Y2=0.865
r33 1 12 43.1362 $w=2.57e-07 $l=3.01413e-07 $layer=POLY_cond $X=3.57 $Y=1.675
+ $X2=3.8 $Y2=1.51
r34 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.57 $Y=1.675 $X2=3.57
+ $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_1%VPWR 1 2 9 13 15 17 22 29 30 33 36
r39 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r43 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=3.245 $Y2=3.33
r44 27 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r48 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=3.245 $Y2=3.33
r50 22 25 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r54 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 15 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=3.245
+ $X2=3.245 $Y2=3.33
r58 11 13 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=3.245 $Y=3.245
+ $X2=3.245 $Y2=2.42
r59 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r60 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.755
r61 2 13 300 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_PDIFF $count=2 $X=3.105
+ $Y=1.835 $X2=3.245 $Y2=2.42
r62 1 9 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.54 $X2=0.69 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_1%Y 1 2 3 12 18 20 23 24 28 30 31 35
c54 35 0 1.01016e-19 $X=2.77 $Y=0.42
c55 28 0 1.90043e-19 $X=1.945 $Y=1.16
r56 30 31 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.705 $Y=0.555
+ $X2=2.705 $Y2=0.925
r57 30 35 5.18599 $w=2.98e-07 $l=1.35e-07 $layer=LI1_cond $X=2.705 $Y=0.555
+ $X2=2.705 $Y2=0.42
r58 29 31 6.14636 $w=2.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.705 $Y=1.085
+ $X2=2.705 $Y2=0.925
r59 23 24 9.42615 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.452 $Y=1.98
+ $X2=1.452 $Y2=1.815
r60 20 29 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.555 $Y=1.17
+ $X2=2.705 $Y2=1.085
r61 20 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.555 $Y=1.17
+ $X2=1.945 $Y2=1.17
r62 16 28 7.03623 $w=1.88e-07 $l=1.18e-07 $layer=LI1_cond $X=1.827 $Y=1.16
+ $X2=1.945 $Y2=1.16
r63 16 25 12.667 $w=1.88e-07 $l=2.17e-07 $layer=LI1_cond $X=1.827 $Y=1.16
+ $X2=1.61 $Y2=1.16
r64 16 18 31.6309 $w=2.33e-07 $l=6.45e-07 $layer=LI1_cond $X=1.827 $Y=1.065
+ $X2=1.827 $Y2=0.42
r65 14 25 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.61 $Y=1.255 $X2=1.61
+ $Y2=1.16
r66 14 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.61 $Y=1.255
+ $X2=1.61 $Y2=1.815
r67 10 23 1.89893 $w=4.83e-07 $l=7.7e-08 $layer=LI1_cond $X=1.452 $Y=2.057
+ $X2=1.452 $Y2=1.98
r68 10 12 21.0362 $w=4.83e-07 $l=8.53e-07 $layer=LI1_cond $X=1.452 $Y=2.057
+ $X2=1.452 $Y2=2.91
r69 3 23 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.835 $X2=1.375 $Y2=1.98
r70 3 12 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.835 $X2=1.375 $Y2=2.91
r71 2 35 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.63
+ $Y=0.235 $X2=2.77 $Y2=0.42
r72 1 18 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.665
+ $Y=0.235 $X2=1.805 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_1%VGND 1 2 3 12 16 20 22 26 31 33 40 41 44 47
+ 50
r55 51 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r56 50 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r58 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 41 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r60 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r61 38 50 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=3.415
+ $Y2=0
r62 38 40 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=4.08
+ $Y2=0
r63 36 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r64 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 33 44 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.35
+ $Y2=0
r66 33 35 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=0.24
+ $Y2=0
r67 31 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r68 31 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r69 31 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r70 26 28 8.03336 $w=6.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.415 $Y=0.38
+ $X2=3.415 $Y2=0.83
r71 24 50 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=0.085
+ $X2=3.415 $Y2=0
r72 24 26 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=0.085
+ $X2=3.415 $Y2=0.38
r73 23 47 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.25
+ $Y2=0
r74 22 50 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.415
+ $Y2=0
r75 22 23 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.385
+ $Y2=0
r76 18 47 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=0.085
+ $X2=2.25 $Y2=0
r77 18 20 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.25 $Y=0.085
+ $X2=2.25 $Y2=0.38
r78 17 44 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.54 $Y=0 $X2=1.35
+ $Y2=0
r79 16 47 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.25
+ $Y2=0
r80 16 17 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=1.54
+ $Y2=0
r81 12 14 13.0408 $w=3.78e-07 $l=4.3e-07 $layer=LI1_cond $X=1.35 $Y=0.38
+ $X2=1.35 $Y2=0.81
r82 10 44 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0
r83 10 12 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0.38
r84 3 28 182 $w=1.7e-07 $l=7.99766e-07 $layer=licon1_NDIFF $count=1 $X=3.105
+ $Y=0.235 $X2=3.585 $Y2=0.83
r85 3 28 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.105
+ $Y=0.235 $X2=3.245 $Y2=0.83
r86 3 26 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.105
+ $Y=0.235 $X2=3.245 $Y2=0.38
r87 2 20 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.095
+ $Y=0.235 $X2=2.28 $Y2=0.38
r88 1 14 182 $w=1.7e-07 $l=5.11664e-07 $layer=licon1_NDIFF $count=1 $X=0.885
+ $Y=0.655 $X2=1.325 $Y2=0.81
r89 1 12 182 $w=1.7e-07 $l=6.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.885
+ $Y=0.655 $X2=1.375 $Y2=0.38
.ends

