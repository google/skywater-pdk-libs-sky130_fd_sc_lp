* File: sky130_fd_sc_lp__nand3_lp.spice
* Created: Fri Aug 28 10:49:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand3_lp.pex.spice"
.subckt sky130_fd_sc_lp__nand3_lp  VNB VPB C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1004 A_155_47# N_C_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1005 A_233_47# N_B_M1005_g A_155_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=44.28 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g A_233_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0882 PD=1.41 PS=0.84 NRD=0 NRS=44.28 M=1 R=2.8 SA=75001.2 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.33 PD=1.28 PS=2.66 NRD=0 NRS=8.8453 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_Y_M1000_d VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000 A=0.25 P=2.5
+ MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__nand3_lp.pxi.spice"
*
.ends
*
*
