* NGSPICE file created from sky130_fd_sc_lp__buflp_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__buflp_m A VGND VNB VPB VPWR X
M1000 a_278_120# A VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.176e+11p ps=1.4e+06u
M1001 VGND a_90_94# a_120_120# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1002 a_304_490# A VPWR VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.596e+11p ps=1.6e+06u
M1003 a_120_490# a_90_94# X VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1004 a_120_120# a_90_94# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1005 a_90_94# A a_278_120# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1006 a_90_94# A a_304_490# VPB phighvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1007 VPWR a_90_94# a_120_490# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

