* File: sky130_fd_sc_lp__isolatch_lp.pxi.spice
* Created: Fri Aug 28 10:42:08 2020
* 
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%D N_D_M1001_g N_D_M1010_g N_D_c_141_n
+ N_D_c_145_n N_D_c_146_n N_D_c_147_n D D N_D_c_143_n
+ PM_SKY130_FD_SC_LP__ISOLATCH_LP%D
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_36_73# N_A_36_73#_M1018_s N_A_36_73#_M1014_d
+ N_A_36_73#_M1008_g N_A_36_73#_M1011_g N_A_36_73#_c_195_n N_A_36_73#_c_196_n
+ N_A_36_73#_c_197_n N_A_36_73#_c_201_n N_A_36_73#_c_202_n N_A_36_73#_c_198_n
+ N_A_36_73#_c_240_p N_A_36_73#_c_221_n N_A_36_73#_c_203_n N_A_36_73#_c_204_n
+ N_A_36_73#_c_205_n N_A_36_73#_c_206_n N_A_36_73#_c_199_n
+ PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_36_73#
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_21_179# N_A_21_179#_M1002_s
+ N_A_21_179#_M1006_s N_A_21_179#_c_323_n N_A_21_179#_c_324_n
+ N_A_21_179#_c_325_n N_A_21_179#_c_339_n N_A_21_179#_c_340_n
+ N_A_21_179#_M1018_g N_A_21_179#_c_327_n N_A_21_179#_c_328_n
+ N_A_21_179#_c_341_n N_A_21_179#_c_342_n N_A_21_179#_c_343_n
+ N_A_21_179#_M1019_g N_A_21_179#_M1013_g N_A_21_179#_M1014_g
+ N_A_21_179#_c_331_n N_A_21_179#_c_332_n N_A_21_179#_c_333_n
+ N_A_21_179#_c_346_n N_A_21_179#_c_347_n N_A_21_179#_c_334_n
+ N_A_21_179#_c_335_n N_A_21_179#_c_336_n N_A_21_179#_c_337_n
+ PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_21_179#
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_458_293# N_A_458_293#_M1007_d
+ N_A_458_293#_M1012_s N_A_458_293#_M1003_g N_A_458_293#_c_483_n
+ N_A_458_293#_M1015_g N_A_458_293#_c_484_n N_A_458_293#_c_485_n
+ N_A_458_293#_M1000_g N_A_458_293#_c_486_n N_A_458_293#_c_487_n
+ N_A_458_293#_c_488_n N_A_458_293#_c_489_n N_A_458_293#_c_490_n
+ N_A_458_293#_c_491_n N_A_458_293#_c_496_n N_A_458_293#_c_497_n
+ N_A_458_293#_c_498_n N_A_458_293#_c_499_n N_A_458_293#_c_500_n
+ N_A_458_293#_c_501_n N_A_458_293#_c_502_n N_A_458_293#_c_503_n
+ N_A_458_293#_c_492_n N_A_458_293#_c_505_n N_A_458_293#_c_493_n
+ PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_458_293#
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%SLEEP_B N_SLEEP_B_M1002_g N_SLEEP_B_c_632_n
+ N_SLEEP_B_c_633_n N_SLEEP_B_M1017_g N_SLEEP_B_c_635_n N_SLEEP_B_M1006_g
+ SLEEP_B PM_SKY130_FD_SC_LP__ISOLATCH_LP%SLEEP_B
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_281_535# N_A_281_535#_M1008_d
+ N_A_281_535#_M1019_d N_A_281_535#_M1016_g N_A_281_535#_M1007_g
+ N_A_281_535#_c_685_n N_A_281_535#_c_686_n N_A_281_535#_c_687_n
+ N_A_281_535#_M1012_g N_A_281_535#_c_689_n N_A_281_535#_M1004_g
+ N_A_281_535#_c_691_n N_A_281_535#_M1009_g N_A_281_535#_c_692_n
+ N_A_281_535#_c_693_n N_A_281_535#_M1005_g N_A_281_535#_c_694_n
+ N_A_281_535#_c_695_n N_A_281_535#_c_696_n N_A_281_535#_c_742_n
+ N_A_281_535#_c_697_n N_A_281_535#_c_698_n N_A_281_535#_c_699_n
+ N_A_281_535#_c_700_n N_A_281_535#_c_701_n N_A_281_535#_c_702_n
+ N_A_281_535#_c_703_n N_A_281_535#_c_704_n N_A_281_535#_c_705_n
+ N_A_281_535#_c_713_n N_A_281_535#_c_706_n N_A_281_535#_c_707_n
+ N_A_281_535#_c_708_n N_A_281_535#_c_709_n N_A_281_535#_c_710_n
+ PM_SKY130_FD_SC_LP__ISOLATCH_LP%A_281_535#
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%VPWR N_VPWR_M1001_s N_VPWR_c_871_n
+ N_VPWR_c_872_n VPWR N_VPWR_c_873_n N_VPWR_c_870_n
+ PM_SKY130_FD_SC_LP__ISOLATCH_LP%VPWR
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%KAPWR N_KAPWR_M1003_d N_KAPWR_M1006_d
+ N_KAPWR_M1012_d KAPWR N_KAPWR_c_937_n N_KAPWR_c_931_n N_KAPWR_c_932_n
+ N_KAPWR_c_933_n PM_SKY130_FD_SC_LP__ISOLATCH_LP%KAPWR
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%Q N_Q_M1005_d N_Q_M1004_d Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__ISOLATCH_LP%Q
x_PM_SKY130_FD_SC_LP__ISOLATCH_LP%VGND N_VGND_M1018_d N_VGND_M1000_d
+ N_VGND_M1017_d N_VGND_M1009_s N_VGND_c_1011_n N_VGND_c_1012_n N_VGND_c_1013_n
+ N_VGND_c_1014_n N_VGND_c_1015_n N_VGND_c_1016_n VGND N_VGND_c_1017_n
+ N_VGND_c_1018_n N_VGND_c_1019_n N_VGND_c_1020_n N_VGND_c_1021_n
+ N_VGND_c_1022_n N_VGND_c_1023_n N_VGND_c_1024_n
+ PM_SKY130_FD_SC_LP__ISOLATCH_LP%VGND
cc_1 VNB N_D_M1010_g 0.0226015f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.835
cc_2 VNB N_D_c_141_n 2.49882e-19 $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.78
cc_3 VNB D 0.0018747f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_D_c_143_n 0.0615195f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.42
cc_5 VNB N_A_36_73#_M1008_g 0.0419915f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.78
cc_6 VNB N_A_36_73#_c_195_n 0.0235012f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A_36_73#_c_196_n 0.00683539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_36_73#_c_197_n 0.00145478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_36_73#_c_198_n 0.00873857f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.515
cc_10 VNB N_A_36_73#_c_199_n 0.0293618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_21_179#_c_323_n 0.0498432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_21_179#_c_324_n 0.0234226f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.78
cc_13 VNB N_A_21_179#_c_325_n 0.0161695f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=2.185
cc_14 VNB N_A_21_179#_M1018_g 0.0160305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_21_179#_c_327_n 0.10639f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_A_21_179#_c_328_n 0.0126405f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_A_21_179#_M1013_g 0.0154886f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.517
cc_18 VNB N_A_21_179#_M1014_g 0.00277745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_21_179#_c_331_n 0.0219731f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.517
cc_20 VNB N_A_21_179#_c_332_n 0.0282782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_21_179#_c_333_n 0.0110498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_21_179#_c_334_n 0.0148136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_21_179#_c_335_n 0.0353142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_21_179#_c_336_n 0.0123141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_21_179#_c_337_n 8.10278e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_458_293#_M1003_g 0.00248794f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.78
cc_27 VNB N_A_458_293#_c_483_n 0.0171921f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=2.35
cc_28 VNB N_A_458_293#_c_484_n 0.0104651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_458_293#_c_485_n 0.018999f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_30 VNB N_A_458_293#_c_486_n 0.0448202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_458_293#_c_487_n 0.02747f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.4
cc_32 VNB N_A_458_293#_c_488_n 0.0170562f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.42
cc_33 VNB N_A_458_293#_c_489_n 0.00390043f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.42
cc_34 VNB N_A_458_293#_c_490_n 0.00412378f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.215
cc_35 VNB N_A_458_293#_c_491_n 0.039119f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.517
cc_36 VNB N_A_458_293#_c_492_n 0.00668846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_458_293#_c_493_n 0.00258424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_SLEEP_B_M1002_g 0.0312556f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.885
cc_39 VNB N_SLEEP_B_c_632_n 0.0108122f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.215
cc_40 VNB N_SLEEP_B_c_633_n 0.0100433f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.835
cc_41 VNB N_SLEEP_B_M1017_g 0.0305589f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.78
cc_42 VNB N_SLEEP_B_c_635_n 0.0273585f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=2.35
cc_43 VNB N_A_281_535#_M1016_g 0.0206524f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=1.78
cc_44 VNB N_A_281_535#_M1007_g 0.0215001f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.35
cc_45 VNB N_A_281_535#_c_685_n 0.0292187f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.35
cc_46 VNB N_A_281_535#_c_686_n 0.0150849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_281_535#_c_687_n 0.011532f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_48 VNB N_A_281_535#_M1012_g 0.00489813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_281_535#_c_689_n 0.0153893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_281_535#_M1004_g 0.00523633f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.42
cc_51 VNB N_A_281_535#_c_691_n 0.0194504f $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=1.517
cc_52 VNB N_A_281_535#_c_692_n 0.0218611f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.517
cc_53 VNB N_A_281_535#_c_693_n 0.01777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_281_535#_c_694_n 0.00723647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_281_535#_c_695_n 0.00423284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_281_535#_c_696_n 0.00621275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_281_535#_c_697_n 0.00136086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_281_535#_c_698_n 0.0073271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_281_535#_c_699_n 0.00131138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_281_535#_c_700_n 0.00938485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_281_535#_c_701_n 0.0165548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_281_535#_c_702_n 0.0034847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_281_535#_c_703_n 0.00194794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_281_535#_c_704_n 0.0179171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_281_535#_c_705_n 0.00459931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_281_535#_c_706_n 0.00204761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_281_535#_c_707_n 0.00694242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_281_535#_c_708_n 0.00675331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_281_535#_c_709_n 0.00137545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_281_535#_c_710_n 0.0322879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VPWR_c_870_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB Q 0.0675912f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.835
cc_73 VNB N_VGND_c_1011_n 0.00777968f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.35
cc_74 VNB N_VGND_c_1012_n 0.00578543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1013_n 0.016703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1014_n 0.0400191f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.42
cc_77 VNB N_VGND_c_1015_n 0.0351124f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.517
cc_78 VNB N_VGND_c_1016_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.517
cc_79 VNB N_VGND_c_1017_n 0.017915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1018_n 0.0576147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1019_n 0.0336247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1020_n 0.0272757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1021_n 0.432381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1022_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1023_n 0.00458122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1024_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VPB N_D_M1001_g 0.0287827f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.885
cc_88 VPB N_D_c_145_n 0.0117679f $X=-0.19 $Y=1.655 $X2=0.21 $Y2=2.185
cc_89 VPB N_D_c_146_n 0.0177172f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.35
cc_90 VPB N_D_c_147_n 0.0364007f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.35
cc_91 VPB D 0.00576989f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_92 VPB N_A_36_73#_M1011_g 0.0274009f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.35
cc_93 VPB N_A_36_73#_c_201_n 0.0106821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_36_73#_c_202_n 0.00544638f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.35
cc_95 VPB N_A_36_73#_c_203_n 0.0010148f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.215
cc_96 VPB N_A_36_73#_c_204_n 0.00821476f $X=-0.19 $Y=1.655 $X2=0.295 $Y2=1.517
cc_97 VPB N_A_36_73#_c_205_n 0.00222158f $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.517
cc_98 VPB N_A_36_73#_c_206_n 0.00116068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_36_73#_c_199_n 0.0506633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_21_179#_c_323_n 0.0136676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_21_179#_c_339_n 0.0422319f $X=-0.19 $Y=1.655 $X2=0.21 $Y2=2.35
cc_102 VPB N_A_21_179#_c_340_n 0.0155209f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_21_179#_c_341_n 0.0132643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_21_179#_c_342_n 0.0341039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_21_179#_c_343_n 0.0108725f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.35
cc_106 VPB N_A_21_179#_M1019_g 0.034289f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.4
cc_107 VPB N_A_21_179#_M1014_g 0.0464124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_21_179#_c_346_n 0.00240565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_21_179#_c_347_n 0.00522774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_21_179#_c_337_n 0.00856073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_458_293#_M1003_g 0.0403969f $X=-0.19 $Y=1.655 $X2=0.21 $Y2=1.78
cc_112 VPB N_A_458_293#_c_491_n 0.0090479f $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.517
cc_113 VPB N_A_458_293#_c_496_n 0.0109458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_458_293#_c_497_n 0.0733712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_458_293#_c_498_n 0.019617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_458_293#_c_499_n 0.00565612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_458_293#_c_500_n 0.00115362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_458_293#_c_501_n 0.0202206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_458_293#_c_502_n 0.0011816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_458_293#_c_503_n 0.0150474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_458_293#_c_492_n 0.00646882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_458_293#_c_505_n 0.00436141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_SLEEP_B_c_635_n 0.0165279f $X=-0.19 $Y=1.655 $X2=0.21 $Y2=2.35
cc_124 VPB N_SLEEP_B_M1006_g 0.0378746f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.35
cc_125 VPB SLEEP_B 0.00386427f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.35
cc_126 VPB N_A_281_535#_M1012_g 0.037411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_281_535#_M1004_g 0.0366806f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.42
cc_128 VPB N_A_281_535#_c_713_n 0.00255956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_281_535#_c_706_n 0.00146698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_281_535#_c_709_n 0.00329002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_281_535#_c_710_n 0.0160038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_871_n 0.0114562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_872_n 0.0118858f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=0.835
cc_134 VPB N_VPWR_c_873_n 0.175904f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.35
cc_135 VPB N_VPWR_c_870_n 0.064352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_KAPWR_c_931_n 0.0108694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_KAPWR_c_932_n 0.00799402f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.215
cc_138 VPB N_KAPWR_c_933_n 0.0613636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB Q 0.0708671f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=0.835
cc_140 N_D_M1010_g N_A_36_73#_M1008_g 0.042821f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_141 N_D_c_143_n N_A_36_73#_M1008_g 0.00465585f $X=0.66 $Y=1.42 $X2=0 $Y2=0
cc_142 N_D_M1010_g N_A_36_73#_c_196_n 0.0154645f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_143 D N_A_36_73#_c_196_n 0.0334495f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_144 N_D_c_143_n N_A_36_73#_c_196_n 0.0124036f $X=0.66 $Y=1.42 $X2=0 $Y2=0
cc_145 N_D_c_141_n N_A_36_73#_c_197_n 0.0117891f $X=0.21 $Y=1.78 $X2=0 $Y2=0
cc_146 D N_A_36_73#_c_197_n 0.010476f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_147 D N_A_36_73#_c_201_n 0.0054076f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_148 N_D_c_146_n N_A_36_73#_c_202_n 0.00960376f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_149 N_D_c_147_n N_A_36_73#_c_202_n 0.00525746f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_150 N_D_M1010_g N_A_36_73#_c_198_n 0.00535908f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_151 D N_A_36_73#_c_198_n 0.0194003f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_152 N_D_c_143_n N_A_36_73#_c_198_n 0.00212951f $X=0.66 $Y=1.42 $X2=0 $Y2=0
cc_153 N_D_M1001_g N_A_36_73#_c_221_n 0.00293823f $X=0.51 $Y=2.885 $X2=0 $Y2=0
cc_154 D N_A_36_73#_c_199_n 0.00234814f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_155 N_D_c_141_n N_A_21_179#_c_323_n 0.039021f $X=0.21 $Y=1.78 $X2=0 $Y2=0
cc_156 N_D_c_145_n N_A_21_179#_c_323_n 0.00210112f $X=0.21 $Y=2.185 $X2=0 $Y2=0
cc_157 N_D_c_143_n N_A_21_179#_c_323_n 0.0192596f $X=0.66 $Y=1.42 $X2=0 $Y2=0
cc_158 N_D_c_141_n N_A_21_179#_c_324_n 2.83068e-19 $X=0.21 $Y=1.78 $X2=0 $Y2=0
cc_159 D N_A_21_179#_c_324_n 0.00153437f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_160 N_D_c_143_n N_A_21_179#_c_324_n 0.00753298f $X=0.66 $Y=1.42 $X2=0 $Y2=0
cc_161 N_D_c_145_n N_A_21_179#_c_339_n 0.00816972f $X=0.21 $Y=2.185 $X2=0 $Y2=0
cc_162 N_D_c_146_n N_A_21_179#_c_339_n 0.00105069f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_163 N_D_c_147_n N_A_21_179#_c_339_n 0.0204884f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_164 D N_A_21_179#_c_339_n 0.0139029f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_165 N_D_c_143_n N_A_21_179#_c_339_n 0.0244079f $X=0.66 $Y=1.42 $X2=0 $Y2=0
cc_166 N_D_c_145_n N_A_21_179#_c_340_n 0.00972573f $X=0.21 $Y=2.185 $X2=0 $Y2=0
cc_167 N_D_c_146_n N_A_21_179#_c_340_n 5.44302e-19 $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_168 N_D_M1010_g N_A_21_179#_M1018_g 0.0120144f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_169 N_D_M1010_g N_A_21_179#_c_327_n 0.00870342f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_170 N_D_c_145_n N_A_21_179#_c_341_n 0.00510788f $X=0.21 $Y=2.185 $X2=0 $Y2=0
cc_171 N_D_c_143_n N_A_21_179#_c_342_n 8.12037e-19 $X=0.66 $Y=1.42 $X2=0 $Y2=0
cc_172 N_D_c_146_n N_A_21_179#_c_343_n 6.64357e-19 $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_173 N_D_c_147_n N_A_21_179#_c_343_n 0.00923361f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_174 N_D_c_147_n N_A_21_179#_M1019_g 0.0114796f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_175 N_D_M1001_g N_VPWR_c_872_n 0.0182862f $X=0.51 $Y=2.885 $X2=0 $Y2=0
cc_176 N_D_c_146_n N_VPWR_c_872_n 0.0210715f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_177 N_D_c_147_n N_VPWR_c_872_n 0.00395665f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_178 N_D_M1001_g N_VPWR_c_873_n 0.00486043f $X=0.51 $Y=2.885 $X2=0 $Y2=0
cc_179 N_D_M1001_g N_VPWR_c_870_n 0.00420493f $X=0.51 $Y=2.885 $X2=0 $Y2=0
cc_180 N_D_M1001_g N_KAPWR_c_933_n 0.00556069f $X=0.51 $Y=2.885 $X2=0 $Y2=0
cc_181 N_D_c_146_n N_KAPWR_c_933_n 0.0152169f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_182 N_D_c_147_n N_KAPWR_c_933_n 0.00479697f $X=0.42 $Y=2.35 $X2=0 $Y2=0
cc_183 N_D_M1010_g N_VGND_c_1011_n 0.00369231f $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_184 N_D_M1010_g N_VGND_c_1021_n 9.49986e-19 $X=1.085 $Y=0.835 $X2=0 $Y2=0
cc_185 N_A_36_73#_c_197_n N_A_21_179#_c_323_n 0.00343014f $X=0.41 $Y=1 $X2=0
+ $Y2=0
cc_186 N_A_36_73#_c_195_n N_A_21_179#_c_324_n 0.00413997f $X=0.325 $Y=0.575
+ $X2=0 $Y2=0
cc_187 N_A_36_73#_c_196_n N_A_21_179#_c_324_n 0.0138269f $X=1.185 $Y=1 $X2=0
+ $Y2=0
cc_188 N_A_36_73#_c_197_n N_A_21_179#_c_324_n 0.00416023f $X=0.41 $Y=1 $X2=0
+ $Y2=0
cc_189 N_A_36_73#_c_195_n N_A_21_179#_c_325_n 0.00306294f $X=0.325 $Y=0.575
+ $X2=0 $Y2=0
cc_190 N_A_36_73#_c_197_n N_A_21_179#_c_325_n 0.00685732f $X=0.41 $Y=1 $X2=0
+ $Y2=0
cc_191 N_A_36_73#_c_201_n N_A_21_179#_c_339_n 0.00772869f $X=1.24 $Y=2.12 $X2=0
+ $Y2=0
cc_192 N_A_36_73#_c_199_n N_A_21_179#_c_339_n 0.0062519f $X=1.925 $Y=1.77 $X2=0
+ $Y2=0
cc_193 N_A_36_73#_c_195_n N_A_21_179#_M1018_g 0.00544809f $X=0.325 $Y=0.575
+ $X2=0 $Y2=0
cc_194 N_A_36_73#_M1008_g N_A_21_179#_c_327_n 0.00907339f $X=1.475 $Y=0.835
+ $X2=0 $Y2=0
cc_195 N_A_36_73#_c_196_n N_A_21_179#_c_327_n 0.00588468f $X=1.185 $Y=1 $X2=0
+ $Y2=0
cc_196 N_A_36_73#_c_202_n N_A_21_179#_c_341_n 0.00177084f $X=1.24 $Y=2.905 $X2=0
+ $Y2=0
cc_197 N_A_36_73#_M1011_g N_A_21_179#_c_342_n 0.0250462f $X=1.925 $Y=2.595 $X2=0
+ $Y2=0
cc_198 N_A_36_73#_c_201_n N_A_21_179#_c_342_n 0.0024754f $X=1.24 $Y=2.12 $X2=0
+ $Y2=0
cc_199 N_A_36_73#_c_202_n N_A_21_179#_c_342_n 0.0115446f $X=1.24 $Y=2.905 $X2=0
+ $Y2=0
cc_200 N_A_36_73#_c_199_n N_A_21_179#_c_342_n 0.0120843f $X=1.925 $Y=1.77 $X2=0
+ $Y2=0
cc_201 N_A_36_73#_c_202_n N_A_21_179#_M1019_g 0.0166459f $X=1.24 $Y=2.905 $X2=0
+ $Y2=0
cc_202 N_A_36_73#_c_240_p N_A_21_179#_M1019_g 0.00637865f $X=2.175 $Y=2.99 $X2=0
+ $Y2=0
cc_203 N_A_36_73#_c_221_n N_A_21_179#_M1019_g 0.00382681f $X=1.325 $Y=2.99 $X2=0
+ $Y2=0
cc_204 N_A_36_73#_M1008_g N_A_21_179#_M1013_g 0.00598758f $X=1.475 $Y=0.835
+ $X2=0 $Y2=0
cc_205 N_A_36_73#_c_203_n N_A_21_179#_M1014_g 7.1043e-19 $X=2.26 $Y=2.905 $X2=0
+ $Y2=0
cc_206 N_A_36_73#_c_204_n N_A_21_179#_M1014_g 0.0206195f $X=3.045 $Y=1.87 $X2=0
+ $Y2=0
cc_207 N_A_36_73#_c_206_n N_A_21_179#_M1014_g 0.0194948f $X=3.21 $Y=2.22 $X2=0
+ $Y2=0
cc_208 N_A_36_73#_c_204_n N_A_21_179#_c_331_n 0.0734263f $X=3.045 $Y=1.87 $X2=0
+ $Y2=0
cc_209 N_A_36_73#_c_205_n N_A_21_179#_c_331_n 0.00832932f $X=2.345 $Y=1.87 $X2=0
+ $Y2=0
cc_210 N_A_36_73#_c_204_n N_A_21_179#_c_332_n 0.00186365f $X=3.045 $Y=1.87 $X2=0
+ $Y2=0
cc_211 N_A_36_73#_M1008_g N_A_21_179#_c_334_n 8.65923e-19 $X=1.475 $Y=0.835
+ $X2=0 $Y2=0
cc_212 N_A_36_73#_c_205_n N_A_21_179#_c_334_n 0.00658711f $X=2.345 $Y=1.87 $X2=0
+ $Y2=0
cc_213 N_A_36_73#_c_199_n N_A_21_179#_c_334_n 9.63504e-19 $X=1.925 $Y=1.77 $X2=0
+ $Y2=0
cc_214 N_A_36_73#_M1008_g N_A_21_179#_c_335_n 0.0090039f $X=1.475 $Y=0.835 $X2=0
+ $Y2=0
cc_215 N_A_36_73#_c_205_n N_A_21_179#_c_335_n 2.48408e-19 $X=2.345 $Y=1.87 $X2=0
+ $Y2=0
cc_216 N_A_36_73#_c_199_n N_A_21_179#_c_335_n 0.00554495f $X=1.925 $Y=1.77 $X2=0
+ $Y2=0
cc_217 N_A_36_73#_M1011_g N_A_458_293#_M1003_g 0.0446486f $X=1.925 $Y=2.595
+ $X2=0 $Y2=0
cc_218 N_A_36_73#_c_240_p N_A_458_293#_M1003_g 0.00518247f $X=2.175 $Y=2.99
+ $X2=0 $Y2=0
cc_219 N_A_36_73#_c_203_n N_A_458_293#_M1003_g 0.0216627f $X=2.26 $Y=2.905 $X2=0
+ $Y2=0
cc_220 N_A_36_73#_c_204_n N_A_458_293#_M1003_g 0.0155469f $X=3.045 $Y=1.87 $X2=0
+ $Y2=0
cc_221 N_A_36_73#_c_205_n N_A_458_293#_M1003_g 0.00262028f $X=2.345 $Y=1.87
+ $X2=0 $Y2=0
cc_222 N_A_36_73#_c_206_n N_A_458_293#_M1003_g 6.70548e-19 $X=3.21 $Y=2.22 $X2=0
+ $Y2=0
cc_223 N_A_36_73#_c_204_n N_A_458_293#_c_488_n 0.00171343f $X=3.045 $Y=1.87
+ $X2=0 $Y2=0
cc_224 N_A_36_73#_c_199_n N_A_458_293#_c_488_n 0.0446486f $X=1.925 $Y=1.77 $X2=0
+ $Y2=0
cc_225 N_A_36_73#_c_204_n N_A_458_293#_c_496_n 0.0117903f $X=3.045 $Y=1.87 $X2=0
+ $Y2=0
cc_226 N_A_36_73#_c_206_n N_A_458_293#_c_496_n 0.0585045f $X=3.21 $Y=2.22 $X2=0
+ $Y2=0
cc_227 N_A_36_73#_c_204_n N_A_458_293#_c_497_n 0.00151642f $X=3.045 $Y=1.87
+ $X2=0 $Y2=0
cc_228 N_A_36_73#_c_206_n N_A_458_293#_c_497_n 0.00409319f $X=3.21 $Y=2.22 $X2=0
+ $Y2=0
cc_229 N_A_36_73#_c_206_n N_A_458_293#_c_499_n 0.0114239f $X=3.21 $Y=2.22 $X2=0
+ $Y2=0
cc_230 N_A_36_73#_c_201_n N_A_281_535#_M1019_d 2.23133e-19 $X=1.24 $Y=2.12 $X2=0
+ $Y2=0
cc_231 N_A_36_73#_c_240_p N_A_281_535#_M1019_d 0.00470753f $X=2.175 $Y=2.99
+ $X2=0 $Y2=0
cc_232 N_A_36_73#_M1008_g N_A_281_535#_c_696_n 0.00602004f $X=1.475 $Y=0.835
+ $X2=0 $Y2=0
cc_233 N_A_36_73#_c_196_n N_A_281_535#_c_696_n 0.00274401f $X=1.185 $Y=1 $X2=0
+ $Y2=0
cc_234 N_A_36_73#_c_198_n N_A_281_535#_c_696_n 0.0153525f $X=1.27 $Y=1.67 $X2=0
+ $Y2=0
cc_235 N_A_36_73#_M1011_g N_A_281_535#_c_713_n 0.00886038f $X=1.925 $Y=2.595
+ $X2=0 $Y2=0
cc_236 N_A_36_73#_c_201_n N_A_281_535#_c_713_n 0.00162468f $X=1.24 $Y=2.12 $X2=0
+ $Y2=0
cc_237 N_A_36_73#_c_202_n N_A_281_535#_c_713_n 0.0332872f $X=1.24 $Y=2.905 $X2=0
+ $Y2=0
cc_238 N_A_36_73#_c_240_p N_A_281_535#_c_713_n 0.0229048f $X=2.175 $Y=2.99 $X2=0
+ $Y2=0
cc_239 N_A_36_73#_c_199_n N_A_281_535#_c_713_n 0.00606045f $X=1.925 $Y=1.77
+ $X2=0 $Y2=0
cc_240 N_A_36_73#_M1008_g N_A_281_535#_c_706_n 0.0022732f $X=1.475 $Y=0.835
+ $X2=0 $Y2=0
cc_241 N_A_36_73#_M1011_g N_A_281_535#_c_706_n 0.0113198f $X=1.925 $Y=2.595
+ $X2=0 $Y2=0
cc_242 N_A_36_73#_c_201_n N_A_281_535#_c_706_n 0.0337799f $X=1.24 $Y=2.12 $X2=0
+ $Y2=0
cc_243 N_A_36_73#_c_202_n N_A_281_535#_c_706_n 0.00687843f $X=1.24 $Y=2.905
+ $X2=0 $Y2=0
cc_244 N_A_36_73#_c_198_n N_A_281_535#_c_706_n 0.00755018f $X=1.27 $Y=1.67 $X2=0
+ $Y2=0
cc_245 N_A_36_73#_c_203_n N_A_281_535#_c_706_n 0.034234f $X=2.26 $Y=2.905 $X2=0
+ $Y2=0
cc_246 N_A_36_73#_c_205_n N_A_281_535#_c_706_n 0.00855488f $X=2.345 $Y=1.87
+ $X2=0 $Y2=0
cc_247 N_A_36_73#_c_199_n N_A_281_535#_c_706_n 0.0203542f $X=1.925 $Y=1.77 $X2=0
+ $Y2=0
cc_248 N_A_36_73#_M1008_g N_A_281_535#_c_707_n 0.0029349f $X=1.475 $Y=0.835
+ $X2=0 $Y2=0
cc_249 N_A_36_73#_M1008_g N_A_281_535#_c_708_n 0.00403458f $X=1.475 $Y=0.835
+ $X2=0 $Y2=0
cc_250 N_A_36_73#_c_198_n N_A_281_535#_c_708_n 0.0110049f $X=1.27 $Y=1.67 $X2=0
+ $Y2=0
cc_251 N_A_36_73#_c_199_n N_A_281_535#_c_708_n 0.00553757f $X=1.925 $Y=1.77
+ $X2=0 $Y2=0
cc_252 N_A_36_73#_M1011_g N_VPWR_c_873_n 0.00596462f $X=1.925 $Y=2.595 $X2=0
+ $Y2=0
cc_253 N_A_36_73#_c_240_p N_VPWR_c_873_n 0.0582113f $X=2.175 $Y=2.99 $X2=0 $Y2=0
cc_254 N_A_36_73#_c_221_n N_VPWR_c_873_n 0.00975041f $X=1.325 $Y=2.99 $X2=0
+ $Y2=0
cc_255 N_A_36_73#_c_206_n N_VPWR_c_873_n 0.0153681f $X=3.21 $Y=2.22 $X2=0 $Y2=0
cc_256 N_A_36_73#_M1014_d N_VPWR_c_870_n 0.00144002f $X=3.07 $Y=2.095 $X2=0
+ $Y2=0
cc_257 N_A_36_73#_M1011_g N_VPWR_c_870_n 0.00712108f $X=1.925 $Y=2.595 $X2=0
+ $Y2=0
cc_258 N_A_36_73#_c_240_p N_VPWR_c_870_n 0.00809996f $X=2.175 $Y=2.99 $X2=0
+ $Y2=0
cc_259 N_A_36_73#_c_221_n N_VPWR_c_870_n 0.00151197f $X=1.325 $Y=2.99 $X2=0
+ $Y2=0
cc_260 N_A_36_73#_c_206_n N_VPWR_c_870_n 0.00228685f $X=3.21 $Y=2.22 $X2=0 $Y2=0
cc_261 N_A_36_73#_c_202_n A_117_535# 0.00390173f $X=1.24 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_262 N_A_36_73#_c_221_n A_117_535# 0.00360727f $X=1.325 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_263 N_A_36_73#_c_240_p A_410_419# 0.00232806f $X=2.175 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_264 N_A_36_73#_c_203_n A_410_419# 0.0095736f $X=2.26 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_265 N_A_36_73#_M1011_g N_KAPWR_c_937_n 3.72163e-19 $X=1.925 $Y=2.595 $X2=0
+ $Y2=0
cc_266 N_A_36_73#_c_240_p N_KAPWR_c_937_n 0.0130124f $X=2.175 $Y=2.99 $X2=0
+ $Y2=0
cc_267 N_A_36_73#_c_203_n N_KAPWR_c_937_n 0.0542111f $X=2.26 $Y=2.905 $X2=0
+ $Y2=0
cc_268 N_A_36_73#_c_204_n N_KAPWR_c_937_n 0.0216087f $X=3.045 $Y=1.87 $X2=0
+ $Y2=0
cc_269 N_A_36_73#_c_206_n N_KAPWR_c_937_n 0.058567f $X=3.21 $Y=2.22 $X2=0 $Y2=0
cc_270 N_A_36_73#_M1014_d N_KAPWR_c_933_n 0.0027681f $X=3.07 $Y=2.095 $X2=0
+ $Y2=0
cc_271 N_A_36_73#_M1011_g N_KAPWR_c_933_n 0.0117926f $X=1.925 $Y=2.595 $X2=0
+ $Y2=0
cc_272 N_A_36_73#_c_201_n N_KAPWR_c_933_n 0.00616966f $X=1.24 $Y=2.12 $X2=0
+ $Y2=0
cc_273 N_A_36_73#_c_202_n N_KAPWR_c_933_n 0.0231729f $X=1.24 $Y=2.905 $X2=0
+ $Y2=0
cc_274 N_A_36_73#_c_240_p N_KAPWR_c_933_n 0.0275246f $X=2.175 $Y=2.99 $X2=0
+ $Y2=0
cc_275 N_A_36_73#_c_221_n N_KAPWR_c_933_n 0.00338685f $X=1.325 $Y=2.99 $X2=0
+ $Y2=0
cc_276 N_A_36_73#_c_203_n N_KAPWR_c_933_n 0.0220696f $X=2.26 $Y=2.905 $X2=0
+ $Y2=0
cc_277 N_A_36_73#_c_206_n N_KAPWR_c_933_n 0.0296322f $X=3.21 $Y=2.22 $X2=0 $Y2=0
cc_278 N_A_36_73#_c_196_n N_VGND_M1018_d 0.0024153f $X=1.185 $Y=1 $X2=-0.19
+ $Y2=-0.245
cc_279 N_A_36_73#_c_195_n N_VGND_c_1011_n 0.0150645f $X=0.325 $Y=0.575 $X2=0
+ $Y2=0
cc_280 N_A_36_73#_c_196_n N_VGND_c_1011_n 0.0241959f $X=1.185 $Y=1 $X2=0 $Y2=0
cc_281 N_A_36_73#_c_195_n N_VGND_c_1017_n 0.0112924f $X=0.325 $Y=0.575 $X2=0
+ $Y2=0
cc_282 N_A_36_73#_M1008_g N_VGND_c_1021_n 9.49986e-19 $X=1.475 $Y=0.835 $X2=0
+ $Y2=0
cc_283 N_A_36_73#_c_195_n N_VGND_c_1021_n 0.00918689f $X=0.325 $Y=0.575 $X2=0
+ $Y2=0
cc_284 N_A_36_73#_c_196_n A_232_125# 0.00263845f $X=1.185 $Y=1 $X2=-0.19
+ $Y2=-0.245
cc_285 N_A_21_179#_M1014_g N_A_458_293#_M1003_g 0.0299853f $X=2.945 $Y=2.595
+ $X2=0 $Y2=0
cc_286 N_A_21_179#_c_327_n N_A_458_293#_c_483_n 0.022402f $X=1.945 $Y=0.18 $X2=0
+ $Y2=0
cc_287 N_A_21_179#_c_331_n N_A_458_293#_c_484_n 0.00113471f $X=3.73 $Y=1.45
+ $X2=0 $Y2=0
cc_288 N_A_21_179#_c_332_n N_A_458_293#_c_484_n 0.018125f $X=2.985 $Y=1.45 $X2=0
+ $Y2=0
cc_289 N_A_21_179#_c_331_n N_A_458_293#_c_486_n 0.00172931f $X=3.73 $Y=1.45
+ $X2=0 $Y2=0
cc_290 N_A_21_179#_c_333_n N_A_458_293#_c_486_n 0.00662194f $X=3.895 $Y=0.76
+ $X2=0 $Y2=0
cc_291 N_A_21_179#_c_331_n N_A_458_293#_c_487_n 0.0100359f $X=3.73 $Y=1.45 $X2=0
+ $Y2=0
cc_292 N_A_21_179#_c_332_n N_A_458_293#_c_487_n 0.0207315f $X=2.985 $Y=1.45
+ $X2=0 $Y2=0
cc_293 N_A_21_179#_c_334_n N_A_458_293#_c_487_n 0.00271227f $X=2.08 $Y=1.06
+ $X2=0 $Y2=0
cc_294 N_A_21_179#_c_331_n N_A_458_293#_c_488_n 0.015262f $X=3.73 $Y=1.45 $X2=0
+ $Y2=0
cc_295 N_A_21_179#_c_334_n N_A_458_293#_c_489_n 2.54817e-19 $X=2.08 $Y=1.06
+ $X2=0 $Y2=0
cc_296 N_A_21_179#_c_335_n N_A_458_293#_c_489_n 0.020808f $X=2.08 $Y=1.06 $X2=0
+ $Y2=0
cc_297 N_A_21_179#_M1014_g N_A_458_293#_c_491_n 0.0165313f $X=2.945 $Y=2.595
+ $X2=0 $Y2=0
cc_298 N_A_21_179#_c_331_n N_A_458_293#_c_491_n 0.0219251f $X=3.73 $Y=1.45 $X2=0
+ $Y2=0
cc_299 N_A_21_179#_c_332_n N_A_458_293#_c_491_n 0.0104982f $X=2.985 $Y=1.45
+ $X2=0 $Y2=0
cc_300 N_A_21_179#_c_337_n N_A_458_293#_c_491_n 0.00332666f $X=4.14 $Y=2.055
+ $X2=0 $Y2=0
cc_301 N_A_21_179#_M1014_g N_A_458_293#_c_496_n 4.08394e-19 $X=2.945 $Y=2.595
+ $X2=0 $Y2=0
cc_302 N_A_21_179#_c_331_n N_A_458_293#_c_496_n 0.0173066f $X=3.73 $Y=1.45 $X2=0
+ $Y2=0
cc_303 N_A_21_179#_c_336_n N_A_458_293#_c_496_n 0.0101636f $X=3.855 $Y=1.45
+ $X2=0 $Y2=0
cc_304 N_A_21_179#_c_337_n N_A_458_293#_c_496_n 0.0733931f $X=4.14 $Y=2.055
+ $X2=0 $Y2=0
cc_305 N_A_21_179#_c_331_n N_A_458_293#_c_497_n 4.73499e-19 $X=3.73 $Y=1.45
+ $X2=0 $Y2=0
cc_306 N_A_21_179#_c_346_n N_A_458_293#_c_497_n 0.00328523f $X=4.14 $Y=2.18
+ $X2=0 $Y2=0
cc_307 N_A_21_179#_c_336_n N_A_458_293#_c_497_n 8.92495e-19 $X=3.855 $Y=1.45
+ $X2=0 $Y2=0
cc_308 N_A_21_179#_c_337_n N_A_458_293#_c_497_n 0.00328523f $X=4.14 $Y=2.055
+ $X2=0 $Y2=0
cc_309 N_A_21_179#_c_347_n N_A_458_293#_c_498_n 0.0179911f $X=4.18 $Y=2.22 $X2=0
+ $Y2=0
cc_310 N_A_21_179#_c_346_n N_A_458_293#_c_500_n 0.0441385f $X=4.14 $Y=2.18 $X2=0
+ $Y2=0
cc_311 N_A_21_179#_c_346_n N_A_458_293#_c_502_n 0.00527847f $X=4.14 $Y=2.18
+ $X2=0 $Y2=0
cc_312 N_A_21_179#_c_337_n N_A_458_293#_c_502_n 0.00624458f $X=4.14 $Y=2.055
+ $X2=0 $Y2=0
cc_313 N_A_21_179#_c_333_n N_SLEEP_B_M1002_g 0.00420496f $X=3.895 $Y=0.76 $X2=0
+ $Y2=0
cc_314 N_A_21_179#_c_336_n N_SLEEP_B_M1002_g 0.00552203f $X=3.855 $Y=1.45 $X2=0
+ $Y2=0
cc_315 N_A_21_179#_c_346_n N_SLEEP_B_c_632_n 0.00240272f $X=4.14 $Y=2.18 $X2=0
+ $Y2=0
cc_316 N_A_21_179#_c_336_n N_SLEEP_B_c_633_n 0.0106809f $X=3.855 $Y=1.45 $X2=0
+ $Y2=0
cc_317 N_A_21_179#_c_336_n N_SLEEP_B_c_635_n 0.00190304f $X=3.855 $Y=1.45 $X2=0
+ $Y2=0
cc_318 N_A_21_179#_c_337_n N_SLEEP_B_c_635_n 0.00175752f $X=4.14 $Y=2.055 $X2=0
+ $Y2=0
cc_319 N_A_21_179#_c_346_n N_SLEEP_B_M1006_g 0.00833797f $X=4.14 $Y=2.18 $X2=0
+ $Y2=0
cc_320 N_A_21_179#_c_337_n N_SLEEP_B_M1006_g 0.00408273f $X=4.14 $Y=2.055 $X2=0
+ $Y2=0
cc_321 N_A_21_179#_c_336_n SLEEP_B 0.013915f $X=3.855 $Y=1.45 $X2=0 $Y2=0
cc_322 N_A_21_179#_c_337_n SLEEP_B 0.0123632f $X=4.14 $Y=2.055 $X2=0 $Y2=0
cc_323 N_A_21_179#_M1013_g N_A_281_535#_c_696_n 0.00184505f $X=2.02 $Y=0.575
+ $X2=0 $Y2=0
cc_324 N_A_21_179#_c_334_n N_A_281_535#_c_696_n 0.0279232f $X=2.08 $Y=1.06 $X2=0
+ $Y2=0
cc_325 N_A_21_179#_c_335_n N_A_281_535#_c_696_n 0.00148649f $X=2.08 $Y=1.06
+ $X2=0 $Y2=0
cc_326 N_A_21_179#_M1013_g N_A_281_535#_c_742_n 0.00856795f $X=2.02 $Y=0.575
+ $X2=0 $Y2=0
cc_327 N_A_21_179#_c_331_n N_A_281_535#_c_742_n 0.00536493f $X=3.73 $Y=1.45
+ $X2=0 $Y2=0
cc_328 N_A_21_179#_c_335_n N_A_281_535#_c_742_n 9.3305e-19 $X=2.08 $Y=1.06 $X2=0
+ $Y2=0
cc_329 N_A_21_179#_M1013_g N_A_281_535#_c_697_n 0.00112728f $X=2.02 $Y=0.575
+ $X2=0 $Y2=0
cc_330 N_A_21_179#_c_334_n N_A_281_535#_c_697_n 0.00373856f $X=2.08 $Y=1.06
+ $X2=0 $Y2=0
cc_331 N_A_21_179#_c_331_n N_A_281_535#_c_698_n 0.0768788f $X=3.73 $Y=1.45 $X2=0
+ $Y2=0
cc_332 N_A_21_179#_c_332_n N_A_281_535#_c_698_n 0.00204154f $X=2.985 $Y=1.45
+ $X2=0 $Y2=0
cc_333 N_A_21_179#_c_333_n N_A_281_535#_c_698_n 0.0139293f $X=3.895 $Y=0.76
+ $X2=0 $Y2=0
cc_334 N_A_21_179#_c_331_n N_A_281_535#_c_699_n 0.0137024f $X=3.73 $Y=1.45 $X2=0
+ $Y2=0
cc_335 N_A_21_179#_c_334_n N_A_281_535#_c_699_n 0.0144066f $X=2.08 $Y=1.06 $X2=0
+ $Y2=0
cc_336 N_A_21_179#_c_335_n N_A_281_535#_c_699_n 6.41702e-19 $X=2.08 $Y=1.06
+ $X2=0 $Y2=0
cc_337 N_A_21_179#_c_333_n N_A_281_535#_c_700_n 0.0269265f $X=3.895 $Y=0.76
+ $X2=0 $Y2=0
cc_338 N_A_21_179#_c_333_n N_A_281_535#_c_701_n 0.0191962f $X=3.895 $Y=0.76
+ $X2=0 $Y2=0
cc_339 N_A_21_179#_c_333_n N_A_281_535#_c_703_n 0.0237732f $X=3.895 $Y=0.76
+ $X2=0 $Y2=0
cc_340 N_A_21_179#_c_333_n N_A_281_535#_c_705_n 0.0139713f $X=3.895 $Y=0.76
+ $X2=0 $Y2=0
cc_341 N_A_21_179#_c_336_n N_A_281_535#_c_705_n 0.00259754f $X=3.855 $Y=1.45
+ $X2=0 $Y2=0
cc_342 N_A_21_179#_c_342_n N_A_281_535#_c_713_n 0.00368305f $X=1.255 $Y=2.25
+ $X2=0 $Y2=0
cc_343 N_A_21_179#_c_342_n N_A_281_535#_c_706_n 9.80173e-19 $X=1.255 $Y=2.25
+ $X2=0 $Y2=0
cc_344 N_A_21_179#_c_334_n N_A_281_535#_c_706_n 0.00806233f $X=2.08 $Y=1.06
+ $X2=0 $Y2=0
cc_345 N_A_21_179#_c_327_n N_A_281_535#_c_707_n 0.00643781f $X=1.945 $Y=0.18
+ $X2=0 $Y2=0
cc_346 N_A_21_179#_M1013_g N_A_281_535#_c_707_n 0.00557612f $X=2.02 $Y=0.575
+ $X2=0 $Y2=0
cc_347 N_A_21_179#_c_334_n N_A_281_535#_c_707_n 0.0216022f $X=2.08 $Y=1.06 $X2=0
+ $Y2=0
cc_348 N_A_21_179#_c_334_n N_A_281_535#_c_708_n 0.0122973f $X=2.08 $Y=1.06 $X2=0
+ $Y2=0
cc_349 N_A_21_179#_M1019_g N_VPWR_c_873_n 0.0035778f $X=1.33 $Y=2.885 $X2=0
+ $Y2=0
cc_350 N_A_21_179#_M1014_g N_VPWR_c_873_n 0.00902772f $X=2.945 $Y=2.595 $X2=0
+ $Y2=0
cc_351 N_A_21_179#_M1019_g N_VPWR_c_870_n 0.00587743f $X=1.33 $Y=2.885 $X2=0
+ $Y2=0
cc_352 N_A_21_179#_M1014_g N_VPWR_c_870_n 0.00888368f $X=2.945 $Y=2.595 $X2=0
+ $Y2=0
cc_353 N_A_21_179#_M1014_g N_KAPWR_c_937_n 0.0152808f $X=2.945 $Y=2.595 $X2=0
+ $Y2=0
cc_354 N_A_21_179#_M1006_s N_KAPWR_c_933_n 0.00688115f $X=4.035 $Y=2.075 $X2=0
+ $Y2=0
cc_355 N_A_21_179#_c_343_n N_KAPWR_c_933_n 0.00828528f $X=0.945 $Y=2.25 $X2=0
+ $Y2=0
cc_356 N_A_21_179#_M1019_g N_KAPWR_c_933_n 0.00296813f $X=1.33 $Y=2.885 $X2=0
+ $Y2=0
cc_357 N_A_21_179#_M1014_g N_KAPWR_c_933_n 0.0100509f $X=2.945 $Y=2.595 $X2=0
+ $Y2=0
cc_358 N_A_21_179#_c_347_n N_KAPWR_c_933_n 0.0193038f $X=4.18 $Y=2.22 $X2=0
+ $Y2=0
cc_359 N_A_21_179#_M1018_g N_VGND_c_1011_n 0.0108093f $X=0.54 $Y=0.575 $X2=0
+ $Y2=0
cc_360 N_A_21_179#_c_327_n N_VGND_c_1011_n 0.0184206f $X=1.945 $Y=0.18 $X2=0
+ $Y2=0
cc_361 N_A_21_179#_c_328_n N_VGND_c_1011_n 0.00388727f $X=0.615 $Y=0.18 $X2=0
+ $Y2=0
cc_362 N_A_21_179#_c_328_n N_VGND_c_1017_n 0.00486043f $X=0.615 $Y=0.18 $X2=0
+ $Y2=0
cc_363 N_A_21_179#_c_327_n N_VGND_c_1018_n 0.0353793f $X=1.945 $Y=0.18 $X2=0
+ $Y2=0
cc_364 N_A_21_179#_c_327_n N_VGND_c_1021_n 0.0441359f $X=1.945 $Y=0.18 $X2=0
+ $Y2=0
cc_365 N_A_21_179#_c_328_n N_VGND_c_1021_n 0.00941964f $X=0.615 $Y=0.18 $X2=0
+ $Y2=0
cc_366 N_A_458_293#_c_486_n N_SLEEP_B_M1002_g 0.00717149f $X=3.515 $Y=0.97 $X2=0
+ $Y2=0
cc_367 N_A_458_293#_c_491_n N_SLEEP_B_c_633_n 0.00717149f $X=3.68 $Y=1.785 $X2=0
+ $Y2=0
cc_368 N_A_458_293#_c_491_n N_SLEEP_B_c_635_n 0.0032678f $X=3.68 $Y=1.785 $X2=0
+ $Y2=0
cc_369 N_A_458_293#_c_501_n N_SLEEP_B_c_635_n 5.52643e-19 $X=5.335 $Y=2.035
+ $X2=0 $Y2=0
cc_370 N_A_458_293#_c_496_n N_SLEEP_B_M1006_g 0.00122622f $X=3.68 $Y=1.95 $X2=0
+ $Y2=0
cc_371 N_A_458_293#_c_497_n N_SLEEP_B_M1006_g 0.00840084f $X=3.68 $Y=1.95 $X2=0
+ $Y2=0
cc_372 N_A_458_293#_c_500_n N_SLEEP_B_M1006_g 0.0268592f $X=4.52 $Y=2.905 $X2=0
+ $Y2=0
cc_373 N_A_458_293#_c_502_n N_SLEEP_B_M1006_g 0.00883607f $X=4.605 $Y=2.035
+ $X2=0 $Y2=0
cc_374 N_A_458_293#_c_501_n SLEEP_B 0.00592885f $X=5.335 $Y=2.035 $X2=0 $Y2=0
cc_375 N_A_458_293#_c_502_n SLEEP_B 0.0137311f $X=4.605 $Y=2.035 $X2=0 $Y2=0
cc_376 N_A_458_293#_c_492_n N_A_281_535#_M1007_g 0.00920935f $X=5.58 $Y=1.915
+ $X2=0 $Y2=0
cc_377 N_A_458_293#_c_493_n N_A_281_535#_M1007_g 5.46324e-19 $X=5.545 $Y=0.61
+ $X2=0 $Y2=0
cc_378 N_A_458_293#_c_492_n N_A_281_535#_c_685_n 0.0118516f $X=5.58 $Y=1.915
+ $X2=0 $Y2=0
cc_379 N_A_458_293#_c_493_n N_A_281_535#_c_685_n 0.00108206f $X=5.545 $Y=0.61
+ $X2=0 $Y2=0
cc_380 N_A_458_293#_c_505_n N_A_281_535#_c_686_n 0.00414139f $X=5.5 $Y=2.08
+ $X2=0 $Y2=0
cc_381 N_A_458_293#_c_492_n N_A_281_535#_c_687_n 0.00527061f $X=5.58 $Y=1.915
+ $X2=0 $Y2=0
cc_382 N_A_458_293#_c_503_n N_A_281_535#_M1012_g 0.0130656f $X=5.5 $Y=2.79 $X2=0
+ $Y2=0
cc_383 N_A_458_293#_c_492_n N_A_281_535#_M1012_g 0.0110394f $X=5.58 $Y=1.915
+ $X2=0 $Y2=0
cc_384 N_A_458_293#_c_505_n N_A_281_535#_M1012_g 0.00390926f $X=5.5 $Y=2.08
+ $X2=0 $Y2=0
cc_385 N_A_458_293#_c_503_n N_A_281_535#_M1004_g 3.10128e-19 $X=5.5 $Y=2.79
+ $X2=0 $Y2=0
cc_386 N_A_458_293#_c_492_n N_A_281_535#_M1004_g 0.00146917f $X=5.58 $Y=1.915
+ $X2=0 $Y2=0
cc_387 N_A_458_293#_c_492_n N_A_281_535#_c_691_n 5.20491e-19 $X=5.58 $Y=1.915
+ $X2=0 $Y2=0
cc_388 N_A_458_293#_c_493_n N_A_281_535#_c_691_n 9.27018e-19 $X=5.545 $Y=0.61
+ $X2=0 $Y2=0
cc_389 N_A_458_293#_c_492_n N_A_281_535#_c_694_n 0.00847731f $X=5.58 $Y=1.915
+ $X2=0 $Y2=0
cc_390 N_A_458_293#_c_483_n N_A_281_535#_c_742_n 0.0085425f $X=2.53 $Y=0.895
+ $X2=0 $Y2=0
cc_391 N_A_458_293#_c_485_n N_A_281_535#_c_742_n 5.68543e-19 $X=2.92 $Y=0.895
+ $X2=0 $Y2=0
cc_392 N_A_458_293#_c_483_n N_A_281_535#_c_697_n 0.0050071f $X=2.53 $Y=0.895
+ $X2=0 $Y2=0
cc_393 N_A_458_293#_c_485_n N_A_281_535#_c_697_n 9.11109e-19 $X=2.92 $Y=0.895
+ $X2=0 $Y2=0
cc_394 N_A_458_293#_c_489_n N_A_281_535#_c_697_n 0.00288283f $X=2.53 $Y=0.97
+ $X2=0 $Y2=0
cc_395 N_A_458_293#_c_484_n N_A_281_535#_c_698_n 0.0143579f $X=2.845 $Y=0.97
+ $X2=0 $Y2=0
cc_396 N_A_458_293#_c_486_n N_A_281_535#_c_698_n 0.0186327f $X=3.515 $Y=0.97
+ $X2=0 $Y2=0
cc_397 N_A_458_293#_c_487_n N_A_281_535#_c_698_n 0.00201986f $X=2.447 $Y=1.465
+ $X2=0 $Y2=0
cc_398 N_A_458_293#_c_489_n N_A_281_535#_c_698_n 0.00101748f $X=2.53 $Y=0.97
+ $X2=0 $Y2=0
cc_399 N_A_458_293#_c_490_n N_A_281_535#_c_698_n 0.00793019f $X=2.92 $Y=0.97
+ $X2=0 $Y2=0
cc_400 N_A_458_293#_c_491_n N_A_281_535#_c_698_n 0.0031103f $X=3.68 $Y=1.785
+ $X2=0 $Y2=0
cc_401 N_A_458_293#_c_487_n N_A_281_535#_c_699_n 0.00288523f $X=2.447 $Y=1.465
+ $X2=0 $Y2=0
cc_402 N_A_458_293#_c_488_n N_A_281_535#_c_699_n 2.00976e-19 $X=2.447 $Y=1.615
+ $X2=0 $Y2=0
cc_403 N_A_458_293#_c_489_n N_A_281_535#_c_699_n 0.00147317f $X=2.53 $Y=0.97
+ $X2=0 $Y2=0
cc_404 N_A_458_293#_c_485_n N_A_281_535#_c_700_n 0.00378091f $X=2.92 $Y=0.895
+ $X2=0 $Y2=0
cc_405 N_A_458_293#_c_486_n N_A_281_535#_c_700_n 0.00723311f $X=3.515 $Y=0.97
+ $X2=0 $Y2=0
cc_406 N_A_458_293#_c_486_n N_A_281_535#_c_701_n 0.00316633f $X=3.515 $Y=0.97
+ $X2=0 $Y2=0
cc_407 N_A_458_293#_c_485_n N_A_281_535#_c_702_n 6.49827e-19 $X=2.92 $Y=0.895
+ $X2=0 $Y2=0
cc_408 N_A_458_293#_M1003_g N_A_281_535#_c_706_n 8.26625e-19 $X=2.415 $Y=2.595
+ $X2=0 $Y2=0
cc_409 N_A_458_293#_c_488_n N_A_281_535#_c_706_n 0.0012367f $X=2.447 $Y=1.615
+ $X2=0 $Y2=0
cc_410 N_A_458_293#_c_483_n N_A_281_535#_c_707_n 9.82387e-19 $X=2.53 $Y=0.895
+ $X2=0 $Y2=0
cc_411 N_A_458_293#_c_487_n N_A_281_535#_c_708_n 4.5389e-19 $X=2.447 $Y=1.465
+ $X2=0 $Y2=0
cc_412 N_A_458_293#_c_501_n N_A_281_535#_c_709_n 0.0227189f $X=5.335 $Y=2.035
+ $X2=0 $Y2=0
cc_413 N_A_458_293#_c_492_n N_A_281_535#_c_709_n 0.0355568f $X=5.58 $Y=1.915
+ $X2=0 $Y2=0
cc_414 N_A_458_293#_c_501_n N_A_281_535#_c_710_n 0.0021942f $X=5.335 $Y=2.035
+ $X2=0 $Y2=0
cc_415 N_A_458_293#_c_492_n N_A_281_535#_c_710_n 0.0037889f $X=5.58 $Y=1.915
+ $X2=0 $Y2=0
cc_416 N_A_458_293#_M1003_g N_VPWR_c_873_n 0.0085571f $X=2.415 $Y=2.595 $X2=0
+ $Y2=0
cc_417 N_A_458_293#_c_498_n N_VPWR_c_873_n 0.0501353f $X=4.435 $Y=2.99 $X2=0
+ $Y2=0
cc_418 N_A_458_293#_c_499_n N_VPWR_c_873_n 0.0236566f $X=3.845 $Y=2.99 $X2=0
+ $Y2=0
cc_419 N_A_458_293#_c_503_n N_VPWR_c_873_n 0.0132298f $X=5.5 $Y=2.79 $X2=0 $Y2=0
cc_420 N_A_458_293#_M1003_g N_VPWR_c_870_n 0.00743141f $X=2.415 $Y=2.595 $X2=0
+ $Y2=0
cc_421 N_A_458_293#_c_498_n N_VPWR_c_870_n 0.00639426f $X=4.435 $Y=2.99 $X2=0
+ $Y2=0
cc_422 N_A_458_293#_c_499_n N_VPWR_c_870_n 0.00310102f $X=3.845 $Y=2.99 $X2=0
+ $Y2=0
cc_423 N_A_458_293#_c_503_n N_VPWR_c_870_n 0.00323356f $X=5.5 $Y=2.79 $X2=0
+ $Y2=0
cc_424 N_A_458_293#_c_501_n N_KAPWR_M1006_d 0.00661026f $X=5.335 $Y=2.035 $X2=0
+ $Y2=0
cc_425 N_A_458_293#_M1003_g N_KAPWR_c_937_n 0.0136681f $X=2.415 $Y=2.595 $X2=0
+ $Y2=0
cc_426 N_A_458_293#_c_500_n N_KAPWR_c_931_n 0.0313939f $X=4.52 $Y=2.905 $X2=0
+ $Y2=0
cc_427 N_A_458_293#_c_501_n N_KAPWR_c_931_n 0.0299249f $X=5.335 $Y=2.035 $X2=0
+ $Y2=0
cc_428 N_A_458_293#_c_503_n N_KAPWR_c_931_n 0.0468088f $X=5.5 $Y=2.79 $X2=0
+ $Y2=0
cc_429 N_A_458_293#_c_503_n N_KAPWR_c_932_n 0.0519067f $X=5.5 $Y=2.79 $X2=0
+ $Y2=0
cc_430 N_A_458_293#_c_505_n N_KAPWR_c_932_n 0.0142226f $X=5.5 $Y=2.08 $X2=0
+ $Y2=0
cc_431 N_A_458_293#_M1003_g N_KAPWR_c_933_n 0.00853161f $X=2.415 $Y=2.595 $X2=0
+ $Y2=0
cc_432 N_A_458_293#_c_496_n N_KAPWR_c_933_n 0.0252026f $X=3.68 $Y=1.95 $X2=0
+ $Y2=0
cc_433 N_A_458_293#_c_498_n N_KAPWR_c_933_n 0.0230877f $X=4.435 $Y=2.99 $X2=0
+ $Y2=0
cc_434 N_A_458_293#_c_499_n N_KAPWR_c_933_n 0.00463476f $X=3.845 $Y=2.99 $X2=0
+ $Y2=0
cc_435 N_A_458_293#_c_500_n N_KAPWR_c_933_n 0.0205382f $X=4.52 $Y=2.905 $X2=0
+ $Y2=0
cc_436 N_A_458_293#_c_501_n N_KAPWR_c_933_n 0.013107f $X=5.335 $Y=2.035 $X2=0
+ $Y2=0
cc_437 N_A_458_293#_c_503_n N_KAPWR_c_933_n 0.0365303f $X=5.5 $Y=2.79 $X2=0
+ $Y2=0
cc_438 N_A_458_293#_c_483_n N_VGND_c_1012_n 0.00221251f $X=2.53 $Y=0.895 $X2=0
+ $Y2=0
cc_439 N_A_458_293#_c_485_n N_VGND_c_1012_n 0.0124138f $X=2.92 $Y=0.895 $X2=0
+ $Y2=0
cc_440 N_A_458_293#_c_486_n N_VGND_c_1012_n 0.0045454f $X=3.515 $Y=0.97 $X2=0
+ $Y2=0
cc_441 N_A_458_293#_c_492_n N_VGND_c_1013_n 0.00202367f $X=5.58 $Y=1.915 $X2=0
+ $Y2=0
cc_442 N_A_458_293#_c_493_n N_VGND_c_1013_n 6.03896e-19 $X=5.545 $Y=0.61 $X2=0
+ $Y2=0
cc_443 N_A_458_293#_c_493_n N_VGND_c_1014_n 0.04733f $X=5.545 $Y=0.61 $X2=0
+ $Y2=0
cc_444 N_A_458_293#_c_483_n N_VGND_c_1018_n 0.00339618f $X=2.53 $Y=0.895 $X2=0
+ $Y2=0
cc_445 N_A_458_293#_c_485_n N_VGND_c_1018_n 0.00386543f $X=2.92 $Y=0.895 $X2=0
+ $Y2=0
cc_446 N_A_458_293#_c_493_n N_VGND_c_1019_n 0.00648527f $X=5.545 $Y=0.61 $X2=0
+ $Y2=0
cc_447 N_A_458_293#_c_483_n N_VGND_c_1021_n 0.00473206f $X=2.53 $Y=0.895 $X2=0
+ $Y2=0
cc_448 N_A_458_293#_c_485_n N_VGND_c_1021_n 0.00760574f $X=2.92 $Y=0.895 $X2=0
+ $Y2=0
cc_449 N_A_458_293#_c_493_n N_VGND_c_1021_n 0.0070224f $X=5.545 $Y=0.61 $X2=0
+ $Y2=0
cc_450 N_SLEEP_B_M1017_g N_A_281_535#_M1016_g 0.0131877f $X=4.47 $Y=0.675 $X2=0
+ $Y2=0
cc_451 N_SLEEP_B_c_635_n N_A_281_535#_c_686_n 0.0131877f $X=4.51 $Y=1.78 $X2=0
+ $Y2=0
cc_452 N_SLEEP_B_M1002_g N_A_281_535#_c_700_n 0.00273135f $X=4.11 $Y=0.675 $X2=0
+ $Y2=0
cc_453 N_SLEEP_B_M1002_g N_A_281_535#_c_701_n 0.0112106f $X=4.11 $Y=0.675 $X2=0
+ $Y2=0
cc_454 N_SLEEP_B_M1017_g N_A_281_535#_c_701_n 8.03883e-19 $X=4.47 $Y=0.675 $X2=0
+ $Y2=0
cc_455 N_SLEEP_B_M1002_g N_A_281_535#_c_703_n 0.0124507f $X=4.11 $Y=0.675 $X2=0
+ $Y2=0
cc_456 N_SLEEP_B_M1017_g N_A_281_535#_c_703_n 0.00727492f $X=4.47 $Y=0.675 $X2=0
+ $Y2=0
cc_457 N_SLEEP_B_M1017_g N_A_281_535#_c_704_n 0.0151372f $X=4.47 $Y=0.675 $X2=0
+ $Y2=0
cc_458 N_SLEEP_B_c_635_n N_A_281_535#_c_704_n 0.00365937f $X=4.51 $Y=1.78 $X2=0
+ $Y2=0
cc_459 SLEEP_B N_A_281_535#_c_704_n 0.0209332f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_460 N_SLEEP_B_M1002_g N_A_281_535#_c_705_n 0.00398284f $X=4.11 $Y=0.675 $X2=0
+ $Y2=0
cc_461 N_SLEEP_B_c_632_n N_A_281_535#_c_705_n 0.00139807f $X=4.355 $Y=1.375
+ $X2=0 $Y2=0
cc_462 N_SLEEP_B_M1017_g N_A_281_535#_c_709_n 8.03338e-19 $X=4.47 $Y=0.675 $X2=0
+ $Y2=0
cc_463 N_SLEEP_B_c_635_n N_A_281_535#_c_709_n 0.00163639f $X=4.51 $Y=1.78 $X2=0
+ $Y2=0
cc_464 SLEEP_B N_A_281_535#_c_709_n 0.0186952f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_465 N_SLEEP_B_c_635_n N_A_281_535#_c_710_n 0.0236505f $X=4.51 $Y=1.78 $X2=0
+ $Y2=0
cc_466 SLEEP_B N_A_281_535#_c_710_n 0.00102746f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_467 N_SLEEP_B_M1006_g N_VPWR_c_873_n 5.41636e-19 $X=4.51 $Y=2.395 $X2=0 $Y2=0
cc_468 N_SLEEP_B_M1006_g N_KAPWR_c_931_n 0.00386397f $X=4.51 $Y=2.395 $X2=0
+ $Y2=0
cc_469 N_SLEEP_B_M1006_g N_KAPWR_c_933_n 0.00273992f $X=4.51 $Y=2.395 $X2=0
+ $Y2=0
cc_470 N_SLEEP_B_M1017_g N_VGND_c_1013_n 0.00162099f $X=4.47 $Y=0.675 $X2=0
+ $Y2=0
cc_471 N_SLEEP_B_M1002_g N_VGND_c_1015_n 7.92274e-19 $X=4.11 $Y=0.675 $X2=0
+ $Y2=0
cc_472 N_SLEEP_B_M1017_g N_VGND_c_1015_n 0.00510437f $X=4.47 $Y=0.675 $X2=0
+ $Y2=0
cc_473 N_SLEEP_B_M1017_g N_VGND_c_1021_n 0.00515964f $X=4.47 $Y=0.675 $X2=0
+ $Y2=0
cc_474 N_A_281_535#_M1012_g N_VPWR_c_873_n 0.00881536f $X=5.765 $Y=2.435 $X2=0
+ $Y2=0
cc_475 N_A_281_535#_M1004_g N_VPWR_c_873_n 0.00907186f $X=6.295 $Y=2.435 $X2=0
+ $Y2=0
cc_476 N_A_281_535#_M1019_d N_VPWR_c_870_n 0.00162345f $X=1.405 $Y=2.675 $X2=0
+ $Y2=0
cc_477 N_A_281_535#_M1012_g N_VPWR_c_870_n 0.00525901f $X=5.765 $Y=2.435 $X2=0
+ $Y2=0
cc_478 N_A_281_535#_M1004_g N_VPWR_c_870_n 0.00525901f $X=6.295 $Y=2.435 $X2=0
+ $Y2=0
cc_479 N_A_281_535#_M1012_g N_KAPWR_c_932_n 0.0183771f $X=5.765 $Y=2.435 $X2=0
+ $Y2=0
cc_480 N_A_281_535#_c_689_n N_KAPWR_c_932_n 0.00207462f $X=6.17 $Y=1.5 $X2=0
+ $Y2=0
cc_481 N_A_281_535#_M1004_g N_KAPWR_c_932_n 0.0160441f $X=6.295 $Y=2.435 $X2=0
+ $Y2=0
cc_482 N_A_281_535#_M1019_d N_KAPWR_c_933_n 0.00120924f $X=1.405 $Y=2.675 $X2=0
+ $Y2=0
cc_483 N_A_281_535#_M1012_g N_KAPWR_c_933_n 0.00949503f $X=5.765 $Y=2.435 $X2=0
+ $Y2=0
cc_484 N_A_281_535#_M1004_g N_KAPWR_c_933_n 0.0113895f $X=6.295 $Y=2.435 $X2=0
+ $Y2=0
cc_485 N_A_281_535#_c_713_n N_KAPWR_c_933_n 0.0257778f $X=1.66 $Y=2.51 $X2=0
+ $Y2=0
cc_486 N_A_281_535#_M1004_g Q 0.018409f $X=6.295 $Y=2.435 $X2=0 $Y2=0
cc_487 N_A_281_535#_c_691_n Q 0.00561572f $X=6.345 $Y=1.425 $X2=0 $Y2=0
cc_488 N_A_281_535#_c_692_n Q 0.0243212f $X=6.63 $Y=1.5 $X2=0 $Y2=0
cc_489 N_A_281_535#_c_693_n Q 0.0223345f $X=6.705 $Y=1.425 $X2=0 $Y2=0
cc_490 N_A_281_535#_c_707_n N_VGND_c_1011_n 0.0106231f $X=1.97 $Y=0.535 $X2=0
+ $Y2=0
cc_491 N_A_281_535#_c_742_n N_VGND_c_1012_n 0.0068731f $X=2.415 $Y=0.64 $X2=0
+ $Y2=0
cc_492 N_A_281_535#_c_697_n N_VGND_c_1012_n 0.00179151f $X=2.5 $Y=0.945 $X2=0
+ $Y2=0
cc_493 N_A_281_535#_c_698_n N_VGND_c_1012_n 0.0169164f $X=3.39 $Y=1.03 $X2=0
+ $Y2=0
cc_494 N_A_281_535#_c_700_n N_VGND_c_1012_n 0.026606f $X=3.475 $Y=0.945 $X2=0
+ $Y2=0
cc_495 N_A_281_535#_c_702_n N_VGND_c_1012_n 0.0146589f $X=3.56 $Y=0.34 $X2=0
+ $Y2=0
cc_496 N_A_281_535#_M1016_g N_VGND_c_1013_n 0.00571646f $X=4.97 $Y=0.675 $X2=0
+ $Y2=0
cc_497 N_A_281_535#_c_701_n N_VGND_c_1013_n 0.0103973f $X=4.15 $Y=0.34 $X2=0
+ $Y2=0
cc_498 N_A_281_535#_c_703_n N_VGND_c_1013_n 0.0137617f $X=4.235 $Y=1.075 $X2=0
+ $Y2=0
cc_499 N_A_281_535#_c_704_n N_VGND_c_1013_n 0.0209461f $X=4.895 $Y=1.16 $X2=0
+ $Y2=0
cc_500 N_A_281_535#_M1007_g N_VGND_c_1014_n 0.0040687f $X=5.33 $Y=0.675 $X2=0
+ $Y2=0
cc_501 N_A_281_535#_c_685_n N_VGND_c_1014_n 0.00273805f $X=5.64 $Y=1.15 $X2=0
+ $Y2=0
cc_502 N_A_281_535#_c_689_n N_VGND_c_1014_n 0.00751391f $X=6.17 $Y=1.5 $X2=0
+ $Y2=0
cc_503 N_A_281_535#_c_691_n N_VGND_c_1014_n 0.0103735f $X=6.345 $Y=1.425 $X2=0
+ $Y2=0
cc_504 N_A_281_535#_c_693_n N_VGND_c_1014_n 4.1944e-19 $X=6.705 $Y=1.425 $X2=0
+ $Y2=0
cc_505 N_A_281_535#_c_701_n N_VGND_c_1015_n 0.0501353f $X=4.15 $Y=0.34 $X2=0
+ $Y2=0
cc_506 N_A_281_535#_c_702_n N_VGND_c_1015_n 0.0121867f $X=3.56 $Y=0.34 $X2=0
+ $Y2=0
cc_507 N_A_281_535#_c_742_n N_VGND_c_1018_n 0.0118193f $X=2.415 $Y=0.64 $X2=0
+ $Y2=0
cc_508 N_A_281_535#_c_707_n N_VGND_c_1018_n 0.0170962f $X=1.97 $Y=0.535 $X2=0
+ $Y2=0
cc_509 N_A_281_535#_M1016_g N_VGND_c_1019_n 0.00510437f $X=4.97 $Y=0.675 $X2=0
+ $Y2=0
cc_510 N_A_281_535#_M1007_g N_VGND_c_1019_n 0.00510437f $X=5.33 $Y=0.675 $X2=0
+ $Y2=0
cc_511 N_A_281_535#_c_691_n N_VGND_c_1020_n 0.00280699f $X=6.345 $Y=1.425 $X2=0
+ $Y2=0
cc_512 N_A_281_535#_c_693_n N_VGND_c_1020_n 3.9957e-19 $X=6.705 $Y=1.425 $X2=0
+ $Y2=0
cc_513 N_A_281_535#_M1016_g N_VGND_c_1021_n 0.00515964f $X=4.97 $Y=0.675 $X2=0
+ $Y2=0
cc_514 N_A_281_535#_M1007_g N_VGND_c_1021_n 0.00515964f $X=5.33 $Y=0.675 $X2=0
+ $Y2=0
cc_515 N_A_281_535#_c_691_n N_VGND_c_1021_n 0.00378994f $X=6.345 $Y=1.425 $X2=0
+ $Y2=0
cc_516 N_A_281_535#_c_742_n N_VGND_c_1021_n 0.0176535f $X=2.415 $Y=0.64 $X2=0
+ $Y2=0
cc_517 N_A_281_535#_c_701_n N_VGND_c_1021_n 0.0287839f $X=4.15 $Y=0.34 $X2=0
+ $Y2=0
cc_518 N_A_281_535#_c_702_n N_VGND_c_1021_n 0.00660921f $X=3.56 $Y=0.34 $X2=0
+ $Y2=0
cc_519 N_A_281_535#_c_707_n N_VGND_c_1021_n 0.0127183f $X=1.97 $Y=0.535 $X2=0
+ $Y2=0
cc_520 N_A_281_535#_c_742_n A_419_73# 0.00758902f $X=2.415 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_521 N_A_281_535#_c_703_n A_837_93# 0.00418617f $X=4.235 $Y=1.075 $X2=-0.19
+ $Y2=-0.245
cc_522 N_VPWR_c_870_n A_117_535# 0.00513254f $X=6.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_523 N_VPWR_c_870_n A_410_419# 9.79222e-19 $X=6.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_524 N_VPWR_c_870_n N_KAPWR_M1003_d 0.00113423f $X=6.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_525 N_VPWR_c_873_n N_KAPWR_c_937_n 0.0189236f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_526 N_VPWR_c_870_n N_KAPWR_c_937_n 0.00299499f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_527 N_VPWR_c_873_n N_KAPWR_c_931_n 0.0136983f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_528 N_VPWR_c_870_n N_KAPWR_c_931_n 0.00148031f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_529 N_VPWR_c_873_n N_KAPWR_c_932_n 0.0131608f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_530 N_VPWR_c_870_n N_KAPWR_c_932_n 0.00321285f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_531 N_VPWR_M1001_s N_KAPWR_c_933_n 0.00237027f $X=0.15 $Y=2.675 $X2=0 $Y2=0
cc_532 N_VPWR_c_871_n N_KAPWR_c_933_n 3.22928e-19 $X=0.295 $Y=3.245 $X2=0 $Y2=0
cc_533 N_VPWR_c_872_n N_KAPWR_c_933_n 0.0270423f $X=0.295 $Y=2.9 $X2=0 $Y2=0
cc_534 N_VPWR_c_873_n N_KAPWR_c_933_n 0.0153279f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_535 N_VPWR_c_870_n N_KAPWR_c_933_n 0.742869f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_536 N_VPWR_c_873_n Q 0.0256651f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_537 N_VPWR_c_870_n Q 0.00628035f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_538 A_117_535# N_KAPWR_c_933_n 0.0203066f $X=0.585 $Y=2.675 $X2=3.21 $Y2=2.22
cc_539 A_410_419# N_KAPWR_c_933_n 0.00510015f $X=2.05 $Y=2.095 $X2=3.21 $Y2=2.22
cc_540 N_KAPWR_c_933_n N_Q_M1004_d 0.00113337f $X=6 $Y=2.82 $X2=0 $Y2=0
cc_541 N_KAPWR_c_932_n Q 0.0309327f $X=6.03 $Y=2.08 $X2=0 $Y2=0
cc_542 N_KAPWR_c_933_n Q 0.0669633f $X=6 $Y=2.82 $X2=0 $Y2=0
cc_543 N_KAPWR_c_932_n N_VGND_c_1014_n 0.00934964f $X=6.03 $Y=2.08 $X2=0 $Y2=0
cc_544 Q N_VGND_c_1014_n 0.0557777f $X=6.875 $Y=0.47 $X2=0 $Y2=0
cc_545 Q N_VGND_c_1020_n 0.0206988f $X=6.875 $Y=0.47 $X2=0 $Y2=0
cc_546 Q N_VGND_c_1021_n 0.0220706f $X=6.875 $Y=0.47 $X2=0 $Y2=0
