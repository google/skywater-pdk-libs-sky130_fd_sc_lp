* NGSPICE file created from sky130_fd_sc_lp__o22a_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 X a_80_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.575e+12p ps=1.006e+07u
M1001 VGND A2 a_303_49# VNB nshort w=840000u l=150000u
+  ad=7.644e+11p pd=6.86e+06u as=7.182e+11p ps=6.75e+06u
M1002 a_303_49# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_80_23# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_566_367# A2 a_80_23# VPB phighvt w=1.26e+06u l=150000u
+  ad=5.103e+11p pd=3.33e+06u as=4.914e+11p ps=3.3e+06u
M1005 X a_80_23# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1006 VPWR A1 a_566_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_80_23# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_80_23# B1 a_303_49# VNB nshort w=840000u l=150000u
+  ad=2.52e+11p pd=2.28e+06u as=0p ps=0u
M1009 a_303_49# B2 a_80_23# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_386_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1011 a_80_23# B2 a_386_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

