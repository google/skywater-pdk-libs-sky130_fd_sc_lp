# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__and2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__and2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.190000 0.880000 2.205000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.830000 1.345000 3.215000 1.760000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 1.075000 2.310000 1.245000 ;
        RECT 1.050000 1.245000 1.285000 1.815000 ;
        RECT 1.050000 1.815000 2.300000 2.145000 ;
        RECT 1.230000 0.255000 1.450000 1.075000 ;
        RECT 2.120000 0.255000 2.310000 1.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.175000  0.720000 0.565000 1.020000 ;
      RECT 0.175000  1.020000 0.425000 2.430000 ;
      RECT 0.175000  2.430000 3.715000 2.610000 ;
      RECT 0.760000  0.085000 1.060000 0.905000 ;
      RECT 0.760000  2.780000 1.090000 3.245000 ;
      RECT 1.495000  1.415000 2.660000 1.645000 ;
      RECT 1.620000  0.085000 1.950000 0.895000 ;
      RECT 1.620000  2.780000 1.950000 3.245000 ;
      RECT 2.480000  0.995000 3.745000 1.165000 ;
      RECT 2.480000  1.165000 2.660000 1.415000 ;
      RECT 2.480000  1.645000 2.660000 1.930000 ;
      RECT 2.480000  1.930000 3.255000 2.260000 ;
      RECT 2.515000  2.780000 2.845000 3.245000 ;
      RECT 2.550000  0.085000 2.880000 0.815000 ;
      RECT 3.385000  1.375000 3.715000 1.545000 ;
      RECT 3.415000  0.255000 3.745000 0.995000 ;
      RECT 3.415000  2.780000 3.745000 3.245000 ;
      RECT 3.545000  1.545000 3.715000 2.430000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__and2b_4
END LIBRARY
