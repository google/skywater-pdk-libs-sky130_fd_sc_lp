* File: sky130_fd_sc_lp__a31oi_lp.pxi.spice
* Created: Fri Aug 28 10:00:20 2020
* 
x_PM_SKY130_FD_SC_LP__A31OI_LP%A3 N_A3_M1007_g N_A3_c_63_n N_A3_M1002_g
+ N_A3_c_64_n N_A3_c_65_n N_A3_c_66_n N_A3_c_67_n A3 A3 N_A3_c_68_n N_A3_c_69_n
+ PM_SKY130_FD_SC_LP__A31OI_LP%A3
x_PM_SKY130_FD_SC_LP__A31OI_LP%A2 N_A2_c_99_n N_A2_M1000_g N_A2_M1003_g
+ N_A2_c_101_n A2 A2 A2 A2 N_A2_c_103_n PM_SKY130_FD_SC_LP__A31OI_LP%A2
x_PM_SKY130_FD_SC_LP__A31OI_LP%A1 N_A1_M1004_g N_A1_c_149_n N_A1_M1001_g
+ N_A1_c_150_n A1 A1 N_A1_c_152_n PM_SKY130_FD_SC_LP__A31OI_LP%A1
x_PM_SKY130_FD_SC_LP__A31OI_LP%B1 N_B1_c_188_n N_B1_M1005_g N_B1_M1008_g
+ N_B1_c_189_n N_B1_M1006_g N_B1_c_190_n N_B1_c_191_n N_B1_c_192_n N_B1_c_193_n
+ B1 B1 N_B1_c_195_n PM_SKY130_FD_SC_LP__A31OI_LP%B1
x_PM_SKY130_FD_SC_LP__A31OI_LP%VPWR N_VPWR_M1007_s N_VPWR_M1000_d N_VPWR_c_238_n
+ N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n VPWR N_VPWR_c_242_n
+ N_VPWR_c_237_n N_VPWR_c_244_n PM_SKY130_FD_SC_LP__A31OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A31OI_LP%A_139_409# N_A_139_409#_M1007_d
+ N_A_139_409#_M1001_d N_A_139_409#_c_272_n N_A_139_409#_c_273_n
+ N_A_139_409#_c_274_n N_A_139_409#_c_275_n
+ PM_SKY130_FD_SC_LP__A31OI_LP%A_139_409#
x_PM_SKY130_FD_SC_LP__A31OI_LP%Y N_Y_M1004_d N_Y_M1008_d N_Y_c_314_n N_Y_c_308_n
+ N_Y_c_309_n N_Y_c_311_n N_Y_c_310_n Y Y PM_SKY130_FD_SC_LP__A31OI_LP%Y
x_PM_SKY130_FD_SC_LP__A31OI_LP%VGND N_VGND_M1002_s N_VGND_M1006_d N_VGND_c_349_n
+ N_VGND_c_350_n N_VGND_c_351_n VGND N_VGND_c_352_n N_VGND_c_353_n
+ N_VGND_c_354_n N_VGND_c_355_n PM_SKY130_FD_SC_LP__A31OI_LP%VGND
cc_1 VNB N_A3_c_63_n 0.0178258f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.73
cc_2 VNB N_A3_c_64_n 0.0197414f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.11
cc_3 VNB N_A3_c_65_n 0.027533f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.615
cc_4 VNB N_A3_c_66_n 0.00325835f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.78
cc_5 VNB N_A3_c_67_n 0.0296553f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.805
cc_6 VNB N_A3_c_68_n 0.018641f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.275
cc_7 VNB N_A3_c_69_n 0.0366214f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.275
cc_8 VNB N_A2_c_99_n 0.00193406f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.78
cc_9 VNB N_A2_M1003_g 0.0300373f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.73
cc_10 VNB N_A2_c_101_n 0.0217904f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.11
cc_11 VNB A2 0.0123076f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.615
cc_12 VNB N_A2_c_103_n 0.015746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1004_g 0.0343948f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=2.545
cc_14 VNB N_A1_c_149_n 0.00211978f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.88
cc_15 VNB N_A1_c_150_n 0.0238828f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.11
cc_16 VNB A1 0.00171029f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.615
cc_17 VNB N_A1_c_152_n 0.0167674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_188_n 0.0135266f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.78
cc_19 VNB N_B1_c_189_n 0.0177624f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.275
cc_20 VNB N_B1_c_190_n 0.023666f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.805
cc_21 VNB N_B1_c_191_n 0.0153942f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_B1_c_192_n 0.023974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_c_193_n 0.00212787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB B1 0.00489144f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.275
cc_25 VNB N_B1_c_195_n 0.0137645f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.295
cc_26 VNB N_VPWR_c_237_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.295
cc_27 VNB N_Y_c_308_n 0.0210079f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.11
cc_28 VNB N_Y_c_309_n 0.00620767f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.615
cc_29 VNB N_Y_c_310_n 0.0340953f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_VGND_c_349_n 0.0221946f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.445
cc_31 VNB N_VGND_c_350_n 0.011456f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.11
cc_32 VNB N_VGND_c_351_n 0.0162633f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.78
cc_33 VNB N_VGND_c_352_n 0.0155085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_353_n 0.045485f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.275
cc_35 VNB N_VGND_c_354_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_355_n 0.182076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A3_M1007_g 0.0416537f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.545
cc_38 VPB N_A3_c_66_n 0.0124658f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.78
cc_39 VPB N_A3_c_69_n 0.00912507f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.275
cc_40 VPB N_A2_c_99_n 0.0109595f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.78
cc_41 VPB N_A2_M1000_g 0.0316344f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=2.545
cc_42 VPB A2 0.00208375f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.615
cc_43 VPB N_A1_c_149_n 0.0117652f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=0.88
cc_44 VPB N_A1_M1001_g 0.0320833f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.73
cc_45 VPB A1 7.45984e-19 $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.615
cc_46 VPB N_B1_M1008_g 0.0359925f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.445
cc_47 VPB N_B1_c_193_n 0.0118303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB B1 0.00200558f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.275
cc_49 VPB N_VPWR_c_238_n 0.0121543f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.73
cc_50 VPB N_VPWR_c_239_n 0.0471248f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.445
cc_51 VPB N_VPWR_c_240_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.78
cc_52 VPB N_VPWR_c_241_n 0.00416546f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_242_n 0.0378977f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_237_n 0.0546255f $X=-0.19 $Y=1.655 $X2=0.41 $Y2=1.295
cc_55 VPB N_VPWR_c_244_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_139_409#_c_272_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.445
cc_57 VPB N_A_139_409#_c_273_n 0.0166938f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.78
cc_58 VPB N_A_139_409#_c_274_n 0.0100597f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=0.805
cc_59 VPB N_A_139_409#_c_275_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_Y_c_311_n 0.018013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_Y_c_310_n 0.0181461f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_62 VPB Y 0.0390561f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_63 N_A3_c_66_n N_A2_c_99_n 0.0115383f $X=0.53 $Y=1.78 $X2=-0.19 $Y2=-0.245
cc_64 N_A3_M1007_g N_A2_M1000_g 0.0196643f $X=0.57 $Y=2.545 $X2=0 $Y2=0
cc_65 N_A3_c_63_n N_A2_M1003_g 0.0407168f $X=0.8 $Y=0.73 $X2=0 $Y2=0
cc_66 N_A3_c_64_n N_A2_M1003_g 0.00553506f $X=0.53 $Y=1.11 $X2=0 $Y2=0
cc_67 N_A3_c_65_n N_A2_c_101_n 0.0115383f $X=0.53 $Y=1.615 $X2=0 $Y2=0
cc_68 N_A3_c_63_n A2 0.00736312f $X=0.8 $Y=0.73 $X2=0 $Y2=0
cc_69 N_A3_c_64_n A2 0.00548279f $X=0.53 $Y=1.11 $X2=0 $Y2=0
cc_70 N_A3_c_68_n A2 0.00248585f $X=0.53 $Y=1.275 $X2=0 $Y2=0
cc_71 N_A3_c_69_n A2 0.0401731f $X=0.53 $Y=1.275 $X2=0 $Y2=0
cc_72 N_A3_c_68_n N_A2_c_103_n 0.0115383f $X=0.53 $Y=1.275 $X2=0 $Y2=0
cc_73 N_A3_c_69_n N_A2_c_103_n 0.00241663f $X=0.53 $Y=1.275 $X2=0 $Y2=0
cc_74 N_A3_M1007_g N_VPWR_c_239_n 0.023763f $X=0.57 $Y=2.545 $X2=0 $Y2=0
cc_75 N_A3_c_66_n N_VPWR_c_239_n 6.00125e-19 $X=0.53 $Y=1.78 $X2=0 $Y2=0
cc_76 N_A3_c_69_n N_VPWR_c_239_n 0.0231278f $X=0.53 $Y=1.275 $X2=0 $Y2=0
cc_77 N_A3_M1007_g N_VPWR_c_240_n 0.00769046f $X=0.57 $Y=2.545 $X2=0 $Y2=0
cc_78 N_A3_M1007_g N_VPWR_c_241_n 8.63241e-19 $X=0.57 $Y=2.545 $X2=0 $Y2=0
cc_79 N_A3_M1007_g N_VPWR_c_237_n 0.0134474f $X=0.57 $Y=2.545 $X2=0 $Y2=0
cc_80 N_A3_M1007_g N_A_139_409#_c_272_n 0.016587f $X=0.57 $Y=2.545 $X2=0 $Y2=0
cc_81 N_A3_M1007_g N_A_139_409#_c_274_n 0.00598056f $X=0.57 $Y=2.545 $X2=0 $Y2=0
cc_82 N_A3_c_69_n N_A_139_409#_c_274_n 0.0018544f $X=0.53 $Y=1.275 $X2=0 $Y2=0
cc_83 N_A3_c_63_n N_VGND_c_349_n 0.0140804f $X=0.8 $Y=0.73 $X2=0 $Y2=0
cc_84 N_A3_c_67_n N_VGND_c_349_n 0.00684764f $X=0.8 $Y=0.805 $X2=0 $Y2=0
cc_85 N_A3_c_68_n N_VGND_c_349_n 8.52482e-19 $X=0.53 $Y=1.275 $X2=0 $Y2=0
cc_86 N_A3_c_69_n N_VGND_c_349_n 0.0119821f $X=0.53 $Y=1.275 $X2=0 $Y2=0
cc_87 N_A3_c_63_n N_VGND_c_353_n 0.00486043f $X=0.8 $Y=0.73 $X2=0 $Y2=0
cc_88 N_A3_c_63_n N_VGND_c_355_n 0.00827383f $X=0.8 $Y=0.73 $X2=0 $Y2=0
cc_89 N_A2_M1003_g N_A1_M1004_g 0.0220003f $X=1.19 $Y=0.445 $X2=0 $Y2=0
cc_90 A2 N_A1_M1004_g 0.0109467f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_91 N_A2_c_99_n N_A1_c_149_n 0.0220003f $X=1.1 $Y=1.79 $X2=0 $Y2=0
cc_92 N_A2_M1000_g N_A1_M1001_g 0.0270132f $X=1.1 $Y=2.545 $X2=0 $Y2=0
cc_93 N_A2_c_101_n N_A1_c_150_n 0.0220003f $X=1.1 $Y=1.625 $X2=0 $Y2=0
cc_94 A2 A1 0.0492677f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_95 N_A2_c_103_n A1 7.73334e-19 $X=1.1 $Y=1.285 $X2=0 $Y2=0
cc_96 N_A2_c_103_n N_A1_c_152_n 0.0220003f $X=1.1 $Y=1.285 $X2=0 $Y2=0
cc_97 N_A2_M1000_g N_VPWR_c_239_n 9.45246e-19 $X=1.1 $Y=2.545 $X2=0 $Y2=0
cc_98 N_A2_M1000_g N_VPWR_c_240_n 0.00769046f $X=1.1 $Y=2.545 $X2=0 $Y2=0
cc_99 N_A2_M1000_g N_VPWR_c_241_n 0.0175124f $X=1.1 $Y=2.545 $X2=0 $Y2=0
cc_100 N_A2_M1000_g N_VPWR_c_237_n 0.0134474f $X=1.1 $Y=2.545 $X2=0 $Y2=0
cc_101 N_A2_M1000_g N_A_139_409#_c_272_n 0.016703f $X=1.1 $Y=2.545 $X2=0 $Y2=0
cc_102 N_A2_c_99_n N_A_139_409#_c_273_n 2.74849e-19 $X=1.1 $Y=1.79 $X2=0 $Y2=0
cc_103 N_A2_M1000_g N_A_139_409#_c_273_n 0.0180783f $X=1.1 $Y=2.545 $X2=0 $Y2=0
cc_104 A2 N_A_139_409#_c_273_n 0.0233693f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_105 N_A2_c_99_n N_A_139_409#_c_274_n 3.03142e-19 $X=1.1 $Y=1.79 $X2=0 $Y2=0
cc_106 N_A2_M1000_g N_A_139_409#_c_274_n 0.00163378f $X=1.1 $Y=2.545 $X2=0 $Y2=0
cc_107 A2 N_A_139_409#_c_274_n 0.00534949f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_108 N_A2_M1000_g N_A_139_409#_c_275_n 9.22077e-19 $X=1.1 $Y=2.545 $X2=0 $Y2=0
cc_109 N_A2_M1003_g N_Y_c_314_n 0.00119561f $X=1.19 $Y=0.445 $X2=0 $Y2=0
cc_110 A2 N_Y_c_314_n 0.0106926f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_111 A2 N_Y_c_309_n 0.00907994f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_112 N_A2_M1003_g N_VGND_c_349_n 0.00228773f $X=1.19 $Y=0.445 $X2=0 $Y2=0
cc_113 A2 N_VGND_c_349_n 0.0173098f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_114 N_A2_M1003_g N_VGND_c_353_n 0.00393362f $X=1.19 $Y=0.445 $X2=0 $Y2=0
cc_115 A2 N_VGND_c_353_n 0.0101611f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_116 N_A2_M1003_g N_VGND_c_355_n 0.00544199f $X=1.19 $Y=0.445 $X2=0 $Y2=0
cc_117 A2 N_VGND_c_355_n 0.0124321f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_118 A2 A_175_47# 0.0035472f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_119 N_A1_M1004_g N_B1_c_188_n 0.0186671f $X=1.58 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A1_M1001_g N_B1_M1008_g 0.0197364f $X=1.67 $Y=2.545 $X2=0 $Y2=0
cc_121 N_A1_M1004_g N_B1_c_191_n 0.00782887f $X=1.58 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A1_c_150_n N_B1_c_192_n 0.0118172f $X=1.67 $Y=1.625 $X2=0 $Y2=0
cc_123 N_A1_c_149_n N_B1_c_193_n 0.0118172f $X=1.67 $Y=1.79 $X2=0 $Y2=0
cc_124 A1 B1 0.0455282f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A1_c_152_n B1 0.0041102f $X=1.67 $Y=1.285 $X2=0 $Y2=0
cc_126 A1 N_B1_c_195_n 8.06741e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A1_c_152_n N_B1_c_195_n 0.0118172f $X=1.67 $Y=1.285 $X2=0 $Y2=0
cc_128 N_A1_M1001_g N_VPWR_c_241_n 0.00313212f $X=1.67 $Y=2.545 $X2=0 $Y2=0
cc_129 N_A1_M1001_g N_VPWR_c_242_n 0.0086001f $X=1.67 $Y=2.545 $X2=0 $Y2=0
cc_130 N_A1_M1001_g N_VPWR_c_237_n 0.0156334f $X=1.67 $Y=2.545 $X2=0 $Y2=0
cc_131 N_A1_M1001_g N_A_139_409#_c_272_n 8.74142e-19 $X=1.67 $Y=2.545 $X2=0
+ $Y2=0
cc_132 N_A1_c_149_n N_A_139_409#_c_273_n 5.7112e-19 $X=1.67 $Y=1.79 $X2=0 $Y2=0
cc_133 N_A1_M1001_g N_A_139_409#_c_273_n 0.0204363f $X=1.67 $Y=2.545 $X2=0 $Y2=0
cc_134 A1 N_A_139_409#_c_273_n 0.0246384f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_135 N_A1_M1001_g N_A_139_409#_c_275_n 0.0146952f $X=1.67 $Y=2.545 $X2=0 $Y2=0
cc_136 N_A1_M1004_g N_Y_c_314_n 0.00911841f $X=1.58 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A1_M1004_g N_Y_c_309_n 0.00486439f $X=1.58 $Y=0.445 $X2=0 $Y2=0
cc_138 A1 N_Y_c_309_n 0.0172717f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A1_c_152_n N_Y_c_309_n 0.00138198f $X=1.67 $Y=1.285 $X2=0 $Y2=0
cc_140 N_A1_M1001_g N_Y_c_311_n 2.76452e-19 $X=1.67 $Y=2.545 $X2=0 $Y2=0
cc_141 N_A1_M1004_g N_VGND_c_353_n 0.00549284f $X=1.58 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A1_M1004_g N_VGND_c_355_n 0.0100377f $X=1.58 $Y=0.445 $X2=0 $Y2=0
cc_143 N_B1_M1008_g N_VPWR_c_242_n 0.00826654f $X=2.2 $Y=2.545 $X2=0 $Y2=0
cc_144 N_B1_M1008_g N_VPWR_c_237_n 0.0156146f $X=2.2 $Y=2.545 $X2=0 $Y2=0
cc_145 N_B1_M1008_g N_A_139_409#_c_273_n 0.00446471f $X=2.2 $Y=2.545 $X2=0 $Y2=0
cc_146 B1 N_A_139_409#_c_273_n 0.00462379f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_147 N_B1_M1008_g N_A_139_409#_c_275_n 0.016587f $X=2.2 $Y=2.545 $X2=0 $Y2=0
cc_148 N_B1_c_188_n N_Y_c_314_n 0.00876976f $X=2.01 $Y=0.73 $X2=0 $Y2=0
cc_149 N_B1_c_189_n N_Y_c_314_n 0.00158177f $X=2.37 $Y=0.73 $X2=0 $Y2=0
cc_150 N_B1_c_190_n N_Y_c_314_n 0.00230187f $X=2.37 $Y=0.805 $X2=0 $Y2=0
cc_151 N_B1_c_190_n N_Y_c_308_n 0.0206836f $X=2.37 $Y=0.805 $X2=0 $Y2=0
cc_152 N_B1_c_191_n N_Y_c_308_n 0.00516508f $X=2.24 $Y=1.12 $X2=0 $Y2=0
cc_153 B1 N_Y_c_308_n 0.0269266f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_154 N_B1_c_195_n N_Y_c_308_n 5.44711e-19 $X=2.24 $Y=1.285 $X2=0 $Y2=0
cc_155 N_B1_c_190_n N_Y_c_309_n 0.00194918f $X=2.37 $Y=0.805 $X2=0 $Y2=0
cc_156 N_B1_M1008_g N_Y_c_311_n 0.00467277f $X=2.2 $Y=2.545 $X2=0 $Y2=0
cc_157 N_B1_c_193_n N_Y_c_311_n 5.95422e-19 $X=2.24 $Y=1.79 $X2=0 $Y2=0
cc_158 B1 N_Y_c_311_n 0.00707451f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_159 N_B1_M1008_g N_Y_c_310_n 0.0071198f $X=2.2 $Y=2.545 $X2=0 $Y2=0
cc_160 N_B1_c_191_n N_Y_c_310_n 0.00500796f $X=2.24 $Y=1.12 $X2=0 $Y2=0
cc_161 B1 N_Y_c_310_n 0.0484816f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B1_c_195_n N_Y_c_310_n 0.0148853f $X=2.24 $Y=1.285 $X2=0 $Y2=0
cc_163 N_B1_M1008_g Y 0.0143689f $X=2.2 $Y=2.545 $X2=0 $Y2=0
cc_164 N_B1_c_188_n N_VGND_c_351_n 0.00216659f $X=2.01 $Y=0.73 $X2=0 $Y2=0
cc_165 N_B1_c_189_n N_VGND_c_351_n 0.0119191f $X=2.37 $Y=0.73 $X2=0 $Y2=0
cc_166 N_B1_c_188_n N_VGND_c_353_n 0.00549284f $X=2.01 $Y=0.73 $X2=0 $Y2=0
cc_167 N_B1_c_189_n N_VGND_c_353_n 0.00486043f $X=2.37 $Y=0.73 $X2=0 $Y2=0
cc_168 N_B1_c_190_n N_VGND_c_353_n 6.21075e-19 $X=2.37 $Y=0.805 $X2=0 $Y2=0
cc_169 N_B1_c_188_n N_VGND_c_355_n 0.00601009f $X=2.01 $Y=0.73 $X2=0 $Y2=0
cc_170 N_B1_c_189_n N_VGND_c_355_n 0.00426155f $X=2.37 $Y=0.73 $X2=0 $Y2=0
cc_171 N_B1_c_190_n N_VGND_c_355_n 8.18184e-19 $X=2.37 $Y=0.805 $X2=0 $Y2=0
cc_172 N_VPWR_c_239_n N_A_139_409#_c_272_n 0.0609159f $X=0.305 $Y=2.19 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_240_n N_A_139_409#_c_272_n 0.021949f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_174 N_VPWR_c_241_n N_A_139_409#_c_272_n 0.0490886f $X=1.365 $Y=2.485 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_237_n N_A_139_409#_c_272_n 0.0124703f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_176 N_VPWR_M1000_d N_A_139_409#_c_273_n 0.00224299f $X=1.225 $Y=2.045 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_241_n N_A_139_409#_c_273_n 0.017764f $X=1.365 $Y=2.485 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_239_n N_A_139_409#_c_274_n 0.00805415f $X=0.305 $Y=2.19 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_241_n N_A_139_409#_c_275_n 0.0218428f $X=1.365 $Y=2.485 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_242_n N_A_139_409#_c_275_n 0.021949f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_181 N_VPWR_c_237_n N_A_139_409#_c_275_n 0.0124703f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_242_n Y 0.0304602f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_237_n Y 0.0174175f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_184 N_A_139_409#_c_273_n N_Y_c_311_n 0.00824572f $X=1.77 $Y=2.055 $X2=0 $Y2=0
cc_185 N_A_139_409#_c_275_n N_Y_c_311_n 0.0624161f $X=1.935 $Y=2.19 $X2=0 $Y2=0
cc_186 N_A_139_409#_c_273_n N_Y_c_310_n 0.00196599f $X=1.77 $Y=2.055 $X2=0 $Y2=0
cc_187 N_Y_c_314_n N_VGND_c_351_n 0.0108736f $X=1.795 $Y=0.47 $X2=0 $Y2=0
cc_188 N_Y_c_308_n N_VGND_c_351_n 0.0238292f $X=2.585 $Y=0.855 $X2=0 $Y2=0
cc_189 N_Y_c_314_n N_VGND_c_353_n 0.0178485f $X=1.795 $Y=0.47 $X2=0 $Y2=0
cc_190 N_Y_M1004_d N_VGND_c_355_n 0.0022543f $X=1.655 $Y=0.235 $X2=0 $Y2=0
cc_191 N_Y_c_314_n N_VGND_c_355_n 0.0124677f $X=1.795 $Y=0.47 $X2=0 $Y2=0
cc_192 N_Y_c_308_n N_VGND_c_355_n 0.0159072f $X=2.585 $Y=0.855 $X2=0 $Y2=0
cc_193 N_VGND_c_355_n A_175_47# 0.00424617f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_194 N_VGND_c_355_n A_253_47# 0.00862756f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_195 N_VGND_c_355_n A_417_47# 0.00286135f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
