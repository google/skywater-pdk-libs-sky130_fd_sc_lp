* File: sky130_fd_sc_lp__srdlrtp_1.pxi.spice
* Created: Wed Sep  2 10:38:27 2020
* 
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%D N_D_M1005_g N_D_M1032_g D N_D_c_213_n
+ PM_SKY130_FD_SC_LP__SRDLRTP_1%D
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%RESET_B N_RESET_B_M1030_g N_RESET_B_M1031_g
+ N_RESET_B_M1022_g N_RESET_B_c_233_n N_RESET_B_M1014_g N_RESET_B_c_234_n
+ N_RESET_B_c_235_n N_RESET_B_c_241_n N_RESET_B_c_242_n RESET_B
+ N_RESET_B_c_243_n N_RESET_B_c_244_n N_RESET_B_c_236_n N_RESET_B_c_237_n
+ PM_SKY130_FD_SC_LP__SRDLRTP_1%RESET_B
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%A_27_97# N_A_27_97#_M1005_s N_A_27_97#_M1032_d
+ N_A_27_97#_M1025_g N_A_27_97#_M1008_g N_A_27_97#_c_389_n N_A_27_97#_c_390_n
+ N_A_27_97#_c_391_n N_A_27_97#_c_392_n N_A_27_97#_c_400_n N_A_27_97#_c_393_n
+ N_A_27_97#_c_394_n N_A_27_97#_c_395_n N_A_27_97#_c_396_n N_A_27_97#_c_397_n
+ N_A_27_97#_c_403_n N_A_27_97#_c_404_n PM_SKY130_FD_SC_LP__SRDLRTP_1%A_27_97#
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%A_336_71# N_A_336_71#_M1006_d
+ N_A_336_71#_M1033_s N_A_336_71#_M1002_g N_A_336_71#_c_481_n
+ N_A_336_71#_c_482_n N_A_336_71#_M1010_g N_A_336_71#_M1027_g
+ N_A_336_71#_c_485_n N_A_336_71#_c_486_n N_A_336_71#_c_515_p
+ N_A_336_71#_c_487_n N_A_336_71#_c_488_n N_A_336_71#_c_489_n
+ N_A_336_71#_c_490_n N_A_336_71#_c_491_n N_A_336_71#_c_492_n
+ N_A_336_71#_c_493_n N_A_336_71#_c_494_n N_A_336_71#_c_495_n
+ N_A_336_71#_c_496_n N_A_336_71#_c_497_n N_A_336_71#_c_498_n
+ N_A_336_71#_c_504_n N_A_336_71#_c_499_n N_A_336_71#_c_500_n
+ N_A_336_71#_c_501_n PM_SKY130_FD_SC_LP__SRDLRTP_1%A_336_71#
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%A_612_71# N_A_612_71#_M1013_d
+ N_A_612_71#_M1014_d N_A_612_71#_M1026_g N_A_612_71#_M1015_g
+ N_A_612_71#_M1028_g N_A_612_71#_c_680_n N_A_612_71#_c_689_n
+ N_A_612_71#_c_690_n N_A_612_71#_c_691_n N_A_612_71#_c_692_n
+ N_A_612_71#_c_693_n N_A_612_71#_c_749_p N_A_612_71#_c_694_n
+ N_A_612_71#_c_695_n N_A_612_71#_c_696_n N_A_612_71#_c_729_n
+ N_A_612_71#_c_708_n N_A_612_71#_c_713_n N_A_612_71#_c_681_n
+ N_A_612_71#_c_682_n N_A_612_71#_c_683_n N_A_612_71#_c_684_n
+ N_A_612_71#_c_732_n N_A_612_71#_c_718_n N_A_612_71#_c_685_n
+ N_A_612_71#_c_686_n PM_SKY130_FD_SC_LP__SRDLRTP_1%A_612_71#
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%A_393_335# N_A_393_335#_M1019_s
+ N_A_393_335#_M1000_d N_A_393_335#_M1018_g N_A_393_335#_c_888_n
+ N_A_393_335#_c_889_n N_A_393_335#_M1021_g N_A_393_335#_c_891_n
+ N_A_393_335#_M1024_g N_A_393_335#_c_893_n N_A_393_335#_c_880_n
+ N_A_393_335#_M1033_g N_A_393_335#_M1006_g N_A_393_335#_c_895_n
+ N_A_393_335#_c_896_n N_A_393_335#_c_882_n N_A_393_335#_c_897_n
+ N_A_393_335#_c_883_n N_A_393_335#_c_884_n N_A_393_335#_c_885_n
+ N_A_393_335#_c_886_n PM_SKY130_FD_SC_LP__SRDLRTP_1%A_393_335#
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%GATE N_GATE_M1000_g N_GATE_M1019_g GATE
+ N_GATE_c_1004_n PM_SKY130_FD_SC_LP__SRDLRTP_1%GATE
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%SLEEP_B N_SLEEP_B_M1020_g N_SLEEP_B_M1035_g
+ N_SLEEP_B_M1001_g N_SLEEP_B_M1023_g N_SLEEP_B_M1003_g N_SLEEP_B_c_1047_n
+ N_SLEEP_B_c_1048_n N_SLEEP_B_M1029_g SLEEP_B SLEEP_B
+ PM_SKY130_FD_SC_LP__SRDLRTP_1%SLEEP_B
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%A_1324_394# N_A_1324_394#_M1029_d
+ N_A_1324_394#_M1023_d N_A_1324_394#_M1007_g N_A_1324_394#_c_1133_n
+ N_A_1324_394#_M1009_g N_A_1324_394#_c_1135_n N_A_1324_394#_c_1156_n
+ N_A_1324_394#_c_1136_n N_A_1324_394#_c_1137_n N_A_1324_394#_c_1140_n
+ PM_SKY130_FD_SC_LP__SRDLRTP_1%A_1324_394#
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%A_438_97# N_A_438_97#_M1010_d
+ N_A_438_97#_M1021_d N_A_438_97#_M1027_s N_A_438_97#_M1011_g
+ N_A_438_97#_M1013_g N_A_438_97#_M1004_g N_A_438_97#_c_1221_n
+ N_A_438_97#_c_1222_n N_A_438_97#_M1017_g N_A_438_97#_M1034_g
+ N_A_438_97#_c_1225_n N_A_438_97#_c_1236_n N_A_438_97#_c_1237_n
+ N_A_438_97#_c_1226_n N_A_438_97#_c_1227_n N_A_438_97#_c_1238_n
+ N_A_438_97#_c_1239_n N_A_438_97#_c_1240_n N_A_438_97#_c_1228_n
+ N_A_438_97#_c_1406_p N_A_438_97#_c_1241_n N_A_438_97#_c_1259_n
+ N_A_438_97#_c_1242_n N_A_438_97#_c_1260_n N_A_438_97#_c_1288_n
+ N_A_438_97#_c_1229_n N_A_438_97#_c_1230_n N_A_438_97#_c_1231_n
+ N_A_438_97#_c_1245_n N_A_438_97#_c_1232_n N_A_438_97#_c_1233_n
+ PM_SKY130_FD_SC_LP__SRDLRTP_1%A_438_97#
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%A_2120_55# N_A_2120_55#_M1017_s
+ N_A_2120_55#_M1034_s N_A_2120_55#_M1016_g N_A_2120_55#_M1012_g
+ N_A_2120_55#_c_1446_n N_A_2120_55#_c_1451_n N_A_2120_55#_c_1447_n
+ N_A_2120_55#_c_1448_n N_A_2120_55#_c_1449_n
+ PM_SKY130_FD_SC_LP__SRDLRTP_1%A_2120_55#
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%VPWR N_VPWR_M1032_s N_VPWR_M1031_d
+ N_VPWR_M1033_d N_VPWR_M1034_d N_VPWR_c_1495_n N_VPWR_c_1496_n N_VPWR_c_1497_n
+ N_VPWR_c_1498_n N_VPWR_c_1499_n VPWR N_VPWR_c_1500_n N_VPWR_c_1501_n
+ N_VPWR_c_1502_n N_VPWR_c_1494_n N_VPWR_c_1504_n N_VPWR_c_1505_n
+ N_VPWR_c_1506_n PM_SKY130_FD_SC_LP__SRDLRTP_1%VPWR
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%A_280_97# N_A_280_97#_M1025_d
+ N_A_280_97#_M1008_d N_A_280_97#_c_1616_n N_A_280_97#_c_1617_n
+ N_A_280_97#_c_1614_n N_A_280_97#_c_1615_n
+ PM_SKY130_FD_SC_LP__SRDLRTP_1%A_280_97#
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%KAPWR N_KAPWR_M1000_s N_KAPWR_M1035_d
+ N_KAPWR_M1028_d N_KAPWR_M1004_d KAPWR N_KAPWR_c_1660_n N_KAPWR_c_1661_n
+ N_KAPWR_c_1666_n N_KAPWR_c_1662_n N_KAPWR_c_1663_n
+ PM_SKY130_FD_SC_LP__SRDLRTP_1%KAPWR
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%Q N_Q_M1016_d N_Q_M1012_d N_Q_c_1777_n
+ N_Q_c_1778_n N_Q_c_1774_n Q Q N_Q_c_1776_n Q PM_SKY130_FD_SC_LP__SRDLRTP_1%Q
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%VGND N_VGND_M1030_d N_VGND_M1015_d
+ N_VGND_M1001_d N_VGND_M1007_d N_VGND_M1017_d N_VGND_c_1799_n N_VGND_c_1800_n
+ N_VGND_c_1801_n N_VGND_c_1802_n N_VGND_c_1803_n N_VGND_c_1804_n
+ N_VGND_c_1805_n N_VGND_c_1806_n N_VGND_c_1807_n VGND N_VGND_c_1808_n
+ N_VGND_c_1809_n N_VGND_c_1810_n N_VGND_c_1811_n N_VGND_c_1812_n
+ N_VGND_c_1813_n PM_SKY130_FD_SC_LP__SRDLRTP_1%VGND
x_PM_SKY130_FD_SC_LP__SRDLRTP_1%A_1624_47# N_A_1624_47#_M1007_s
+ N_A_1624_47#_M1022_d N_A_1624_47#_c_1932_n N_A_1624_47#_c_1929_n
+ N_A_1624_47#_c_1930_n N_A_1624_47#_c_1931_n
+ PM_SKY130_FD_SC_LP__SRDLRTP_1%A_1624_47#
cc_1 VNB N_D_M1005_g 0.0275463f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.695
cc_2 VNB N_D_M1032_g 0.0193156f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.755
cc_3 VNB D 0.01487f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_D_c_213_n 0.0571862f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.245
cc_5 VNB N_RESET_B_M1030_g 0.0468127f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.695
cc_6 VNB N_RESET_B_c_233_n 0.0335245f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.245
cc_7 VNB N_RESET_B_c_234_n 0.0174603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_RESET_B_c_235_n 0.0110407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_RESET_B_c_236_n 0.0126718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_RESET_B_c_237_n 0.00503495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_97#_c_389_n 0.0173017f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.245
cc_12 VNB N_A_27_97#_c_390_n 0.02684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_97#_c_391_n 0.0192729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_97#_c_392_n 0.0113867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_97#_c_393_n 0.00717989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_97#_c_394_n 0.00342539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_97#_c_395_n 0.0163484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_97#_c_396_n 0.023752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_97#_c_397_n 8.03993e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_336_71#_M1002_g 0.0183206f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_21 VNB N_A_336_71#_c_481_n 0.0121167f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.245
cc_22 VNB N_A_336_71#_c_482_n 0.00808919f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.245
cc_23 VNB N_A_336_71#_M1010_g 0.0204622f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.245
cc_24 VNB N_A_336_71#_M1027_g 0.0868811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_336_71#_c_485_n 0.0119492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_336_71#_c_486_n 0.00610625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_336_71#_c_487_n 0.0134679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_336_71#_c_488_n 0.0131843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_336_71#_c_489_n 0.0272609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_336_71#_c_490_n 5.38139e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_336_71#_c_491_n 0.00655005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_336_71#_c_492_n 0.00363795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_336_71#_c_493_n 4.43157e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_336_71#_c_494_n 0.0124592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_336_71#_c_495_n 0.00303305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_336_71#_c_496_n 0.00392484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_336_71#_c_497_n 0.00162134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_336_71#_c_498_n 0.00432058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_336_71#_c_499_n 0.00342822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_336_71#_c_500_n 0.0416763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_336_71#_c_501_n 0.0317632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_612_71#_M1026_g 0.0194963f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_43 VNB N_A_612_71#_M1015_g 0.0225882f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.245
cc_44 VNB N_A_612_71#_c_680_n 0.00391367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_612_71#_c_681_n 0.0174435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_612_71#_c_682_n 0.00254381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_612_71#_c_683_n 0.00112679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_612_71#_c_684_n 0.0116041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_612_71#_c_685_n 0.010102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_612_71#_c_686_n 0.0372197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_393_335#_M1024_g 0.0509017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_393_335#_c_880_n 0.0733265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_393_335#_M1006_g 0.0270501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_393_335#_c_882_n 0.00302669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_393_335#_c_883_n 0.0059243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_393_335#_c_884_n 0.0100022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_393_335#_c_885_n 0.00455433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_393_335#_c_886_n 0.0142127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_GATE_M1019_g 0.0227698f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.755
cc_60 VNB GATE 0.00657653f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_61 VNB N_GATE_c_1004_n 0.0252355f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.245
cc_62 VNB N_SLEEP_B_M1020_g 0.0206104f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.695
cc_63 VNB N_SLEEP_B_M1001_g 0.0228234f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.245
cc_64 VNB N_SLEEP_B_M1003_g 0.0234003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_SLEEP_B_c_1047_n 0.01957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_SLEEP_B_c_1048_n 0.0517399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_SLEEP_B_M1029_g 0.0233041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1324_394#_M1007_g 0.0261351f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_69 VNB N_A_1324_394#_c_1133_n 0.0515123f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.245
cc_70 VNB N_A_1324_394#_M1009_g 0.0261047f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.245
cc_71 VNB N_A_1324_394#_c_1135_n 0.00163005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1324_394#_c_1136_n 0.0160277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1324_394#_c_1137_n 0.0253413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_438_97#_M1011_g 0.0285303f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.245
cc_75 VNB N_A_438_97#_M1013_g 0.0329815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_438_97#_M1004_g 0.0215025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_438_97#_c_1221_n 0.0646062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_438_97#_c_1222_n 0.038592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_438_97#_M1017_g 0.0469723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_438_97#_M1034_g 0.0175593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_438_97#_c_1225_n 0.00574765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_438_97#_c_1226_n 0.00637298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_438_97#_c_1227_n 0.00665884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_438_97#_c_1228_n 0.00613465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_438_97#_c_1229_n 0.00450394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_438_97#_c_1230_n 0.00657999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_438_97#_c_1231_n 0.00294655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_438_97#_c_1232_n 0.0179625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_438_97#_c_1233_n 0.00671908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2120_55#_M1016_g 0.027575f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_91 VNB N_A_2120_55#_M1012_g 5.51802e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.245
cc_92 VNB N_A_2120_55#_c_1446_n 0.0125939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2120_55#_c_1447_n 0.0093588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2120_55#_c_1448_n 0.0353978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2120_55#_c_1449_n 0.00336498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VPWR_c_1494_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_280_97#_c_1614_n 0.00298751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_280_97#_c_1615_n 0.00932818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_Q_c_1774_n 0.0244783f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.245
cc_100 VNB Q 0.00971172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_Q_c_1776_n 0.0301057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1799_n 0.0180334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1800_n 0.0117751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1801_n 0.00838292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1802_n 0.0289671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1803_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1804_n 0.0151292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1805_n 0.0624918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1806_n 0.0508852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1807_n 0.00632327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1808_n 0.053829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1809_n 0.0583191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1810_n 0.0185363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1811_n 0.654882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1812_n 0.0109039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1813_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_1624_47#_c_1929_n 0.00454708f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.245
cc_118 VNB N_A_1624_47#_c_1930_n 0.0027632f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.245
cc_119 VNB N_A_1624_47#_c_1931_n 0.00332489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VPB N_D_M1032_g 0.0764439f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.755
cc_121 VPB N_RESET_B_M1030_g 0.0147977f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.695
cc_122 VPB N_RESET_B_M1031_g 0.0231033f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.755
cc_123 VPB N_RESET_B_M1014_g 0.0254486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_RESET_B_c_241_n 0.0746693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_RESET_B_c_242_n 0.00304991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_RESET_B_c_243_n 0.0430607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_RESET_B_c_244_n 0.00448239f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_RESET_B_c_236_n 0.0311418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_27_97#_M1008_g 0.0501393f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.245
cc_130 VPB N_A_27_97#_c_391_n 0.0120709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_27_97#_c_400_n 0.00171751f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_27_97#_c_393_n 0.00457896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_27_97#_c_397_n 0.00101839f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_27_97#_c_403_n 0.0137263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_27_97#_c_404_n 0.00161401f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_336_71#_M1027_g 0.0520955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_336_71#_c_488_n 0.00133307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_336_71#_c_504_n 0.00113418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_612_71#_M1028_g 0.0234533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_612_71#_c_680_n 0.0204318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_612_71#_c_689_n 0.0264312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_612_71#_c_690_n 0.00306263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_612_71#_c_691_n 0.00250607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_612_71#_c_692_n 0.00744448f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_612_71#_c_693_n 0.00208089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_612_71#_c_694_n 0.00974687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_612_71#_c_695_n 8.37163e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_612_71#_c_696_n 9.14535e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_612_71#_c_681_n 0.00909277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_612_71#_c_683_n 0.00499144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_612_71#_c_684_n 0.0177343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_393_335#_M1018_g 0.0388136f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_153 VPB N_A_393_335#_c_888_n 0.0081647f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.245
cc_154 VPB N_A_393_335#_c_889_n 0.00837111f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.245
cc_155 VPB N_A_393_335#_M1021_g 0.0457005f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.245
cc_156 VPB N_A_393_335#_c_891_n 0.0144336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_393_335#_M1024_g 0.00125789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_393_335#_c_893_n 0.0759691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_393_335#_c_880_n 0.0533232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_393_335#_c_895_n 0.0104023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_393_335#_c_896_n 0.00741022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_393_335#_c_897_n 0.00128662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_393_335#_c_883_n 0.00747577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_GATE_M1000_g 0.0799373f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.695
cc_165 VPB GATE 0.00261172f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_166 VPB N_GATE_c_1004_n 0.00533921f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.245
cc_167 VPB N_SLEEP_B_M1035_g 0.0663813f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.755
cc_168 VPB N_SLEEP_B_M1023_g 0.0586233f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.245
cc_169 VPB N_SLEEP_B_c_1048_n 0.0205483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_1324_394#_M1009_g 0.0404612f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.245
cc_171 VPB N_A_1324_394#_c_1135_n 0.00510288f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_1324_394#_c_1140_n 0.00438429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_438_97#_M1004_g 0.0471973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_438_97#_M1034_g 0.0284303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_438_97#_c_1236_n 0.00213543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_438_97#_c_1237_n 0.0101486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_438_97#_c_1238_n 0.00970918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_438_97#_c_1239_n 0.00391778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_438_97#_c_1240_n 0.00396974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_438_97#_c_1241_n 0.0219773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_438_97#_c_1242_n 0.00808942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_438_97#_c_1230_n 0.0138789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_438_97#_c_1231_n 2.75787e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_438_97#_c_1245_n 0.00398462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_2120_55#_M1012_g 0.028321f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.245
cc_186 VPB N_A_2120_55#_c_1451_n 0.0127054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1495_n 0.0111279f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.245
cc_188 VPB N_VPWR_c_1496_n 0.0113222f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.245
cc_189 VPB N_VPWR_c_1497_n 0.018502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1498_n 0.00976484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1499_n 0.0202297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1500_n 0.0754428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1501_n 0.171114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1502_n 0.0185366f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1494_n 0.0735944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1504_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1505_n 0.017235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1506_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_280_97#_c_1616_n 0.00204432f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_200 VPB N_A_280_97#_c_1617_n 0.00120814f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.245
cc_201 VPB N_A_280_97#_c_1615_n 0.00747475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_KAPWR_c_1660_n 0.00514394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_KAPWR_c_1661_n 0.0033174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_KAPWR_c_1662_n 0.0153539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_KAPWR_c_1663_n 0.0643793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_Q_c_1777_n 0.0362634f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_207 VPB N_Q_c_1778_n 0.00971172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_Q_c_1774_n 0.00773243f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.245
cc_209 N_D_M1005_g N_RESET_B_M1030_g 0.0480533f $X=0.495 $Y=0.695 $X2=0 $Y2=0
cc_210 N_D_M1032_g N_RESET_B_c_243_n 0.0286762f $X=0.495 $Y=2.755 $X2=0 $Y2=0
cc_211 N_D_c_213_n N_RESET_B_c_243_n 0.0480533f $X=0.495 $Y=1.245 $X2=0 $Y2=0
cc_212 N_D_M1005_g N_A_27_97#_c_392_n 0.0103449f $X=0.495 $Y=0.695 $X2=0 $Y2=0
cc_213 D N_A_27_97#_c_392_n 0.024798f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_214 N_D_M1032_g N_A_27_97#_c_400_n 0.00338179f $X=0.495 $Y=2.755 $X2=0 $Y2=0
cc_215 N_D_M1005_g N_A_27_97#_c_396_n 0.0186778f $X=0.495 $Y=0.695 $X2=0 $Y2=0
cc_216 D N_A_27_97#_c_396_n 0.0260514f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_217 N_D_c_213_n N_A_27_97#_c_396_n 0.00231791f $X=0.495 $Y=1.245 $X2=0 $Y2=0
cc_218 N_D_M1032_g N_A_27_97#_c_397_n 0.00534437f $X=0.495 $Y=2.755 $X2=0 $Y2=0
cc_219 N_D_M1032_g N_A_27_97#_c_403_n 0.0176056f $X=0.495 $Y=2.755 $X2=0 $Y2=0
cc_220 N_D_M1032_g N_VPWR_c_1496_n 0.00894485f $X=0.495 $Y=2.755 $X2=0 $Y2=0
cc_221 N_D_M1032_g N_VPWR_c_1497_n 0.00469214f $X=0.495 $Y=2.755 $X2=0 $Y2=0
cc_222 N_D_M1032_g N_VPWR_c_1494_n 0.00373058f $X=0.495 $Y=2.755 $X2=0 $Y2=0
cc_223 N_D_M1032_g N_KAPWR_c_1663_n 0.0101068f $X=0.495 $Y=2.755 $X2=0 $Y2=0
cc_224 N_D_M1005_g N_VGND_c_1802_n 0.00386132f $X=0.495 $Y=0.695 $X2=0 $Y2=0
cc_225 N_D_M1005_g N_VGND_c_1811_n 0.00509887f $X=0.495 $Y=0.695 $X2=0 $Y2=0
cc_226 N_RESET_B_M1030_g N_A_27_97#_M1008_g 0.00508923f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_227 N_RESET_B_M1031_g N_A_27_97#_M1008_g 0.0217263f $X=0.995 $Y=2.755 $X2=0
+ $Y2=0
cc_228 N_RESET_B_c_241_n N_A_27_97#_M1008_g 0.0108383f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_229 N_RESET_B_c_242_n N_A_27_97#_M1008_g 0.00135047f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_230 N_RESET_B_c_243_n N_A_27_97#_M1008_g 0.0159562f $X=0.995 $Y=2.09 $X2=0
+ $Y2=0
cc_231 N_RESET_B_c_244_n N_A_27_97#_M1008_g 0.00205759f $X=1.11 $Y=2.09 $X2=0
+ $Y2=0
cc_232 N_RESET_B_M1030_g N_A_27_97#_c_389_n 0.010322f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_233 N_RESET_B_c_241_n N_A_27_97#_c_391_n 0.00129059f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_234 N_RESET_B_c_243_n N_A_27_97#_c_391_n 0.00745317f $X=0.995 $Y=2.09 $X2=0
+ $Y2=0
cc_235 N_RESET_B_c_244_n N_A_27_97#_c_391_n 5.17957e-19 $X=1.11 $Y=2.09 $X2=0
+ $Y2=0
cc_236 N_RESET_B_M1030_g N_A_27_97#_c_392_n 0.00799575f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_237 N_RESET_B_M1031_g N_A_27_97#_c_400_n 0.00621615f $X=0.995 $Y=2.755 $X2=0
+ $Y2=0
cc_238 N_RESET_B_M1030_g N_A_27_97#_c_393_n 0.0158223f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_239 N_RESET_B_c_241_n N_A_27_97#_c_393_n 0.00409371f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_240 N_RESET_B_c_242_n N_A_27_97#_c_393_n 0.00841911f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_241 N_RESET_B_c_243_n N_A_27_97#_c_393_n 0.00233841f $X=0.995 $Y=2.09 $X2=0
+ $Y2=0
cc_242 N_RESET_B_c_244_n N_A_27_97#_c_393_n 0.0273278f $X=1.11 $Y=2.09 $X2=0
+ $Y2=0
cc_243 N_RESET_B_M1030_g N_A_27_97#_c_394_n 0.00192836f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_244 N_RESET_B_M1030_g N_A_27_97#_c_395_n 0.0403486f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_245 N_RESET_B_M1030_g N_A_27_97#_c_396_n 0.00149664f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_246 N_RESET_B_M1030_g N_A_27_97#_c_403_n 0.00534751f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_247 N_RESET_B_c_242_n N_A_27_97#_c_403_n 0.00127867f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_248 N_RESET_B_c_243_n N_A_27_97#_c_403_n 0.00509567f $X=0.995 $Y=2.09 $X2=0
+ $Y2=0
cc_249 N_RESET_B_c_244_n N_A_27_97#_c_403_n 0.0241429f $X=1.11 $Y=2.09 $X2=0
+ $Y2=0
cc_250 N_RESET_B_M1031_g N_A_27_97#_c_404_n 0.0041896f $X=0.995 $Y=2.755 $X2=0
+ $Y2=0
cc_251 N_RESET_B_c_243_n N_A_27_97#_c_404_n 0.0037912f $X=0.995 $Y=2.09 $X2=0
+ $Y2=0
cc_252 N_RESET_B_c_241_n N_A_336_71#_M1027_g 0.0051188f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_253 N_RESET_B_c_241_n N_A_336_71#_c_488_n 0.00463621f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_254 N_RESET_B_c_241_n N_A_336_71#_c_496_n 0.0100595f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_255 N_RESET_B_c_241_n N_A_336_71#_c_504_n 0.0205884f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_256 RESET_B N_A_612_71#_M1014_d 0.00114225f $X=9.275 $Y=1.95 $X2=0 $Y2=0
cc_257 N_RESET_B_c_237_n N_A_612_71#_M1014_d 0.0035607f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_258 N_RESET_B_c_241_n N_A_612_71#_M1028_g 0.00454477f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_259 N_RESET_B_c_241_n N_A_612_71#_c_680_n 0.0176234f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_260 N_RESET_B_c_241_n N_A_612_71#_c_689_n 0.00807173f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_261 N_RESET_B_c_241_n N_A_612_71#_c_692_n 0.0134352f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_262 N_RESET_B_c_241_n N_A_612_71#_c_693_n 0.00127682f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_263 N_RESET_B_c_241_n N_A_612_71#_c_696_n 0.0183696f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_264 N_RESET_B_M1014_g N_A_612_71#_c_708_n 0.0163285f $X=9.16 $Y=2.595 $X2=0
+ $Y2=0
cc_265 N_RESET_B_c_241_n N_A_612_71#_c_708_n 0.0399952f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_266 RESET_B N_A_612_71#_c_708_n 9.32318e-19 $X=9.275 $Y=1.95 $X2=0 $Y2=0
cc_267 N_RESET_B_c_236_n N_A_612_71#_c_708_n 3.00716e-19 $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_268 N_RESET_B_c_237_n N_A_612_71#_c_708_n 0.00675061f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_269 N_RESET_B_c_237_n N_A_612_71#_c_713_n 0.0140944f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_270 N_RESET_B_c_237_n N_A_612_71#_c_681_n 0.0476584f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_271 N_RESET_B_c_241_n N_A_612_71#_c_682_n 0.00553691f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_272 N_RESET_B_c_241_n N_A_612_71#_c_683_n 0.0105806f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_273 N_RESET_B_c_241_n N_A_612_71#_c_684_n 0.00209789f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_274 N_RESET_B_M1014_g N_A_612_71#_c_718_n 0.0153975f $X=9.16 $Y=2.595 $X2=0
+ $Y2=0
cc_275 RESET_B N_A_612_71#_c_718_n 7.04285e-19 $X=9.275 $Y=1.95 $X2=0 $Y2=0
cc_276 N_RESET_B_c_236_n N_A_612_71#_c_718_n 8.7245e-19 $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_277 N_RESET_B_c_237_n N_A_612_71#_c_718_n 0.0267201f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_278 N_RESET_B_c_241_n N_A_393_335#_M1000_d 0.00225499f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_279 N_RESET_B_c_241_n N_A_393_335#_M1018_g 0.0105814f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_280 N_RESET_B_c_241_n N_A_393_335#_c_888_n 6.4692e-19 $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_281 N_RESET_B_c_241_n N_A_393_335#_M1021_g 0.0141001f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_282 N_RESET_B_c_241_n N_A_393_335#_c_880_n 0.0233236f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_283 N_RESET_B_c_241_n N_A_393_335#_c_896_n 0.0123968f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_284 N_RESET_B_c_241_n N_A_393_335#_c_897_n 0.0131379f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_285 N_RESET_B_c_241_n N_A_393_335#_c_883_n 0.0214327f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_286 N_RESET_B_c_241_n N_GATE_M1000_g 0.00173607f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_287 N_RESET_B_c_241_n N_SLEEP_B_M1035_g 0.00394222f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_288 N_RESET_B_c_241_n N_SLEEP_B_M1023_g 0.0043417f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_289 N_RESET_B_c_241_n N_SLEEP_B_c_1048_n 0.00672995f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_290 N_RESET_B_c_241_n SLEEP_B 0.013437f $X=9.215 $Y=2.035 $X2=0 $Y2=0
cc_291 N_RESET_B_c_241_n N_A_1324_394#_M1023_d 0.00225499f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_292 N_RESET_B_c_234_n N_A_1324_394#_M1007_g 0.0189512f $X=9.09 $Y=0.765 $X2=0
+ $Y2=0
cc_293 N_RESET_B_c_233_n N_A_1324_394#_c_1133_n 0.0797643f $X=9.11 $Y=1.605
+ $X2=0 $Y2=0
cc_294 N_RESET_B_c_235_n N_A_1324_394#_c_1133_n 0.00401446f $X=9.09 $Y=0.915
+ $X2=0 $Y2=0
cc_295 N_RESET_B_c_241_n N_A_1324_394#_M1009_g 0.00880874f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_296 RESET_B N_A_1324_394#_M1009_g 3.98422e-19 $X=9.275 $Y=1.95 $X2=0 $Y2=0
cc_297 N_RESET_B_c_236_n N_A_1324_394#_M1009_g 0.0701235f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_298 N_RESET_B_c_237_n N_A_1324_394#_M1009_g 0.00334072f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_299 N_RESET_B_c_233_n N_A_1324_394#_c_1137_n 8.13733e-19 $X=9.11 $Y=1.605
+ $X2=0 $Y2=0
cc_300 N_RESET_B_c_235_n N_A_1324_394#_c_1137_n 2.4449e-19 $X=9.09 $Y=0.915
+ $X2=0 $Y2=0
cc_301 N_RESET_B_c_241_n N_A_1324_394#_c_1140_n 0.00846276f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_302 N_RESET_B_c_234_n N_A_438_97#_M1011_g 0.0129517f $X=9.09 $Y=0.765 $X2=0
+ $Y2=0
cc_303 N_RESET_B_c_235_n N_A_438_97#_M1011_g 0.0162787f $X=9.09 $Y=0.915 $X2=0
+ $Y2=0
cc_304 N_RESET_B_c_233_n N_A_438_97#_M1004_g 0.00540022f $X=9.11 $Y=1.605 $X2=0
+ $Y2=0
cc_305 N_RESET_B_M1014_g N_A_438_97#_M1004_g 0.0278708f $X=9.16 $Y=2.595 $X2=0
+ $Y2=0
cc_306 N_RESET_B_c_236_n N_A_438_97#_M1004_g 0.0181679f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_307 N_RESET_B_c_237_n N_A_438_97#_M1004_g 0.032214f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_308 N_RESET_B_c_233_n N_A_438_97#_c_1222_n 0.0162787f $X=9.11 $Y=1.605 $X2=0
+ $Y2=0
cc_309 N_RESET_B_c_236_n N_A_438_97#_c_1222_n 0.00671841f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_310 N_RESET_B_c_237_n N_A_438_97#_c_1222_n 0.00777955f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_311 N_RESET_B_c_241_n N_A_438_97#_c_1236_n 0.00205789f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_312 N_RESET_B_c_241_n N_A_438_97#_c_1238_n 0.0104053f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_313 N_RESET_B_c_241_n N_A_438_97#_c_1239_n 0.0155137f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_314 N_RESET_B_c_241_n N_A_438_97#_c_1241_n 0.105135f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_315 N_RESET_B_c_241_n N_A_438_97#_c_1259_n 0.00866278f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_316 N_RESET_B_c_241_n N_A_438_97#_c_1260_n 0.00974163f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_317 N_RESET_B_c_233_n N_A_438_97#_c_1229_n 0.0132222f $X=9.11 $Y=1.605 $X2=0
+ $Y2=0
cc_318 N_RESET_B_c_241_n N_A_438_97#_c_1229_n 0.00416495f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_319 RESET_B N_A_438_97#_c_1229_n 0.00139998f $X=9.275 $Y=1.95 $X2=0 $Y2=0
cc_320 N_RESET_B_c_236_n N_A_438_97#_c_1229_n 0.00314453f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_321 N_RESET_B_c_237_n N_A_438_97#_c_1229_n 0.0423181f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_322 N_RESET_B_c_241_n N_A_438_97#_c_1230_n 0.0333509f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_323 N_RESET_B_c_241_n N_A_438_97#_c_1231_n 0.00630652f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_324 N_RESET_B_c_241_n N_A_438_97#_c_1245_n 0.0391277f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_325 N_RESET_B_c_241_n N_A_438_97#_c_1232_n 0.0274478f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_326 N_RESET_B_c_233_n N_A_438_97#_c_1233_n 0.00994234f $X=9.11 $Y=1.605 $X2=0
+ $Y2=0
cc_327 N_RESET_B_c_235_n N_A_438_97#_c_1233_n 0.00123929f $X=9.09 $Y=0.915 $X2=0
+ $Y2=0
cc_328 N_RESET_B_c_241_n N_VPWR_M1033_d 0.00483465f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_329 N_RESET_B_M1031_g N_VPWR_c_1496_n 0.00107912f $X=0.995 $Y=2.755 $X2=0
+ $Y2=0
cc_330 N_RESET_B_M1031_g N_VPWR_c_1497_n 0.00529818f $X=0.995 $Y=2.755 $X2=0
+ $Y2=0
cc_331 N_RESET_B_M1031_g N_VPWR_c_1498_n 0.00879363f $X=0.995 $Y=2.755 $X2=0
+ $Y2=0
cc_332 N_RESET_B_c_241_n N_VPWR_c_1498_n 0.00446587f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_333 N_RESET_B_c_242_n N_VPWR_c_1498_n 0.0011714f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_334 N_RESET_B_c_243_n N_VPWR_c_1498_n 0.0026557f $X=0.995 $Y=2.09 $X2=0 $Y2=0
cc_335 N_RESET_B_c_244_n N_VPWR_c_1498_n 0.0115637f $X=1.11 $Y=2.09 $X2=0 $Y2=0
cc_336 N_RESET_B_M1014_g N_VPWR_c_1501_n 0.00975641f $X=9.16 $Y=2.595 $X2=0
+ $Y2=0
cc_337 N_RESET_B_M1031_g N_VPWR_c_1494_n 0.00560347f $X=0.995 $Y=2.755 $X2=0
+ $Y2=0
cc_338 N_RESET_B_M1014_g N_VPWR_c_1494_n 0.0078066f $X=9.16 $Y=2.595 $X2=0 $Y2=0
cc_339 N_RESET_B_c_241_n N_A_280_97#_c_1616_n 0.00708898f $X=9.215 $Y=2.035
+ $X2=0 $Y2=0
cc_340 N_RESET_B_M1031_g N_A_280_97#_c_1615_n 9.3735e-19 $X=0.995 $Y=2.755 $X2=0
+ $Y2=0
cc_341 N_RESET_B_c_241_n N_A_280_97#_c_1615_n 0.0264906f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_342 N_RESET_B_c_242_n N_A_280_97#_c_1615_n 0.00233076f $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_343 N_RESET_B_c_243_n N_A_280_97#_c_1615_n 4.25244e-19 $X=0.995 $Y=2.09 $X2=0
+ $Y2=0
cc_344 N_RESET_B_c_244_n N_A_280_97#_c_1615_n 0.0118662f $X=1.11 $Y=2.09 $X2=0
+ $Y2=0
cc_345 N_RESET_B_c_241_n N_KAPWR_M1028_d 0.00240778f $X=9.215 $Y=2.035 $X2=0
+ $Y2=0
cc_346 N_RESET_B_M1014_g N_KAPWR_c_1666_n 0.00252581f $X=9.16 $Y=2.595 $X2=0
+ $Y2=0
cc_347 N_RESET_B_M1031_g N_KAPWR_c_1663_n 0.00503971f $X=0.995 $Y=2.755 $X2=0
+ $Y2=0
cc_348 N_RESET_B_M1014_g N_KAPWR_c_1663_n 0.0108012f $X=9.16 $Y=2.595 $X2=0
+ $Y2=0
cc_349 N_RESET_B_c_242_n N_KAPWR_c_1663_n 0.0127877f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_350 RESET_B N_KAPWR_c_1663_n 0.0128099f $X=9.275 $Y=1.95 $X2=0 $Y2=0
cc_351 N_RESET_B_c_243_n N_KAPWR_c_1663_n 0.00135801f $X=0.995 $Y=2.09 $X2=0
+ $Y2=0
cc_352 N_RESET_B_c_244_n N_KAPWR_c_1663_n 0.00640821f $X=1.11 $Y=2.09 $X2=0
+ $Y2=0
cc_353 N_RESET_B_c_237_n N_KAPWR_c_1663_n 0.00144507f $X=9.39 $Y=1.77 $X2=0
+ $Y2=0
cc_354 N_RESET_B_c_241_n A_1565_419# 0.0040317f $X=9.215 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_355 N_RESET_B_c_241_n A_1765_419# 0.00174357f $X=9.215 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_356 N_RESET_B_M1030_g N_VGND_c_1799_n 0.00329625f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_357 N_RESET_B_M1030_g N_VGND_c_1802_n 0.00497279f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_358 N_RESET_B_c_234_n N_VGND_c_1809_n 0.00404211f $X=9.09 $Y=0.765 $X2=0
+ $Y2=0
cc_359 N_RESET_B_M1030_g N_VGND_c_1811_n 0.00509887f $X=0.855 $Y=0.695 $X2=0
+ $Y2=0
cc_360 N_RESET_B_c_234_n N_VGND_c_1811_n 0.00605843f $X=9.09 $Y=0.765 $X2=0
+ $Y2=0
cc_361 N_RESET_B_c_234_n N_VGND_c_1812_n 0.00392695f $X=9.09 $Y=0.765 $X2=0
+ $Y2=0
cc_362 N_RESET_B_c_234_n N_A_1624_47#_c_1932_n 7.9013e-19 $X=9.09 $Y=0.765 $X2=0
+ $Y2=0
cc_363 N_RESET_B_c_234_n N_A_1624_47#_c_1929_n 0.0102024f $X=9.09 $Y=0.765 $X2=0
+ $Y2=0
cc_364 N_RESET_B_c_234_n N_A_1624_47#_c_1931_n 0.00674093f $X=9.09 $Y=0.765
+ $X2=0 $Y2=0
cc_365 N_RESET_B_c_235_n N_A_1624_47#_c_1931_n 0.00133922f $X=9.09 $Y=0.915
+ $X2=0 $Y2=0
cc_366 N_A_27_97#_c_389_n N_A_336_71#_M1002_g 0.0124145f $X=1.305 $Y=1.015 $X2=0
+ $Y2=0
cc_367 N_A_27_97#_c_394_n N_A_336_71#_M1002_g 2.76524e-19 $X=1.305 $Y=1.18 $X2=0
+ $Y2=0
cc_368 N_A_27_97#_c_395_n N_A_336_71#_M1002_g 0.0071867f $X=1.305 $Y=1.18 $X2=0
+ $Y2=0
cc_369 N_A_27_97#_c_390_n N_A_336_71#_c_482_n 0.0071867f $X=1.305 $Y=1.535 $X2=0
+ $Y2=0
cc_370 N_A_27_97#_c_391_n N_A_336_71#_c_482_n 2.18762e-19 $X=1.61 $Y=1.61 $X2=0
+ $Y2=0
cc_371 N_A_27_97#_c_390_n N_A_336_71#_c_501_n 0.00278537f $X=1.305 $Y=1.535
+ $X2=0 $Y2=0
cc_372 N_A_27_97#_M1008_g N_A_393_335#_M1018_g 0.0251097f $X=1.61 $Y=2.755 $X2=0
+ $Y2=0
cc_373 N_A_27_97#_c_391_n N_A_393_335#_c_889_n 0.0251097f $X=1.61 $Y=1.61 $X2=0
+ $Y2=0
cc_374 N_A_27_97#_c_400_n N_VPWR_c_1496_n 0.013992f $X=0.78 $Y=2.75 $X2=0 $Y2=0
cc_375 N_A_27_97#_c_400_n N_VPWR_c_1497_n 0.0206168f $X=0.78 $Y=2.75 $X2=0 $Y2=0
cc_376 N_A_27_97#_M1008_g N_VPWR_c_1498_n 0.00761183f $X=1.61 $Y=2.755 $X2=0
+ $Y2=0
cc_377 N_A_27_97#_c_393_n N_VPWR_c_1498_n 0.0020928f $X=1.14 $Y=1.665 $X2=0
+ $Y2=0
cc_378 N_A_27_97#_c_404_n N_VPWR_c_1498_n 0.0388066f $X=0.775 $Y=2.595 $X2=0
+ $Y2=0
cc_379 N_A_27_97#_M1008_g N_VPWR_c_1500_n 0.00529818f $X=1.61 $Y=2.755 $X2=0
+ $Y2=0
cc_380 N_A_27_97#_M1008_g N_VPWR_c_1494_n 0.00533311f $X=1.61 $Y=2.755 $X2=0
+ $Y2=0
cc_381 N_A_27_97#_c_400_n N_VPWR_c_1494_n 0.00304853f $X=0.78 $Y=2.75 $X2=0
+ $Y2=0
cc_382 N_A_27_97#_M1008_g N_A_280_97#_c_1616_n 0.00340479f $X=1.61 $Y=2.755
+ $X2=0 $Y2=0
cc_383 N_A_27_97#_M1008_g N_A_280_97#_c_1617_n 0.00596204f $X=1.61 $Y=2.755
+ $X2=0 $Y2=0
cc_384 N_A_27_97#_c_389_n N_A_280_97#_c_1614_n 0.00481772f $X=1.305 $Y=1.015
+ $X2=0 $Y2=0
cc_385 N_A_27_97#_c_391_n N_A_280_97#_c_1614_n 0.00429858f $X=1.61 $Y=1.61 $X2=0
+ $Y2=0
cc_386 N_A_27_97#_c_394_n N_A_280_97#_c_1614_n 0.00537787f $X=1.305 $Y=1.18
+ $X2=0 $Y2=0
cc_387 N_A_27_97#_c_395_n N_A_280_97#_c_1614_n 3.61461e-19 $X=1.305 $Y=1.18
+ $X2=0 $Y2=0
cc_388 N_A_27_97#_M1008_g N_A_280_97#_c_1615_n 0.0200324f $X=1.61 $Y=2.755 $X2=0
+ $Y2=0
cc_389 N_A_27_97#_c_389_n N_A_280_97#_c_1615_n 0.00217723f $X=1.305 $Y=1.015
+ $X2=0 $Y2=0
cc_390 N_A_27_97#_c_391_n N_A_280_97#_c_1615_n 0.00550818f $X=1.61 $Y=1.61 $X2=0
+ $Y2=0
cc_391 N_A_27_97#_c_393_n N_A_280_97#_c_1615_n 0.0121057f $X=1.14 $Y=1.665 $X2=0
+ $Y2=0
cc_392 N_A_27_97#_c_394_n N_A_280_97#_c_1615_n 0.038781f $X=1.305 $Y=1.18 $X2=0
+ $Y2=0
cc_393 N_A_27_97#_c_395_n N_A_280_97#_c_1615_n 0.00524606f $X=1.305 $Y=1.18
+ $X2=0 $Y2=0
cc_394 N_A_27_97#_M1032_d N_KAPWR_c_1663_n 0.00173511f $X=0.57 $Y=2.435 $X2=0
+ $Y2=0
cc_395 N_A_27_97#_M1008_g N_KAPWR_c_1663_n 0.00875171f $X=1.61 $Y=2.755 $X2=0
+ $Y2=0
cc_396 N_A_27_97#_c_400_n N_KAPWR_c_1663_n 0.0346362f $X=0.78 $Y=2.75 $X2=0
+ $Y2=0
cc_397 N_A_27_97#_c_404_n N_KAPWR_c_1663_n 3.51259e-19 $X=0.775 $Y=2.595 $X2=0
+ $Y2=0
cc_398 N_A_27_97#_c_396_n A_114_97# 0.00196091f $X=0.28 $Y=0.685 $X2=-0.19
+ $Y2=-0.245
cc_399 N_A_27_97#_c_389_n N_VGND_c_1799_n 0.0030567f $X=1.305 $Y=1.015 $X2=0
+ $Y2=0
cc_400 N_A_27_97#_c_394_n N_VGND_c_1799_n 0.00458736f $X=1.305 $Y=1.18 $X2=0
+ $Y2=0
cc_401 N_A_27_97#_c_395_n N_VGND_c_1799_n 4.11901e-19 $X=1.305 $Y=1.18 $X2=0
+ $Y2=0
cc_402 N_A_27_97#_c_396_n N_VGND_c_1799_n 0.00464705f $X=0.28 $Y=0.685 $X2=0
+ $Y2=0
cc_403 N_A_27_97#_c_396_n N_VGND_c_1802_n 0.0136054f $X=0.28 $Y=0.685 $X2=0
+ $Y2=0
cc_404 N_A_27_97#_c_389_n N_VGND_c_1805_n 0.00475526f $X=1.305 $Y=1.015 $X2=0
+ $Y2=0
cc_405 N_A_27_97#_c_389_n N_VGND_c_1811_n 0.00509887f $X=1.305 $Y=1.015 $X2=0
+ $Y2=0
cc_406 N_A_27_97#_c_396_n N_VGND_c_1811_n 0.0199511f $X=0.28 $Y=0.685 $X2=0
+ $Y2=0
cc_407 N_A_336_71#_c_515_p N_A_612_71#_M1026_g 0.00875001f $X=3.9 $Y=0.61 $X2=0
+ $Y2=0
cc_408 N_A_336_71#_c_498_n N_A_612_71#_M1026_g 0.00311173f $X=2.925 $Y=0.34
+ $X2=0 $Y2=0
cc_409 N_A_336_71#_c_515_p N_A_612_71#_M1015_g 0.0112328f $X=3.9 $Y=0.61 $X2=0
+ $Y2=0
cc_410 N_A_336_71#_c_487_n N_A_612_71#_M1015_g 0.00500501f $X=3.985 $Y=0.925
+ $X2=0 $Y2=0
cc_411 N_A_336_71#_c_488_n N_A_612_71#_M1015_g 0.00137376f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_412 N_A_336_71#_M1027_g N_A_612_71#_c_694_n 0.0146972f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_413 N_A_336_71#_M1027_g N_A_612_71#_c_696_n 0.00206757f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_414 N_A_336_71#_M1027_g N_A_612_71#_c_729_n 0.00437666f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_415 N_A_336_71#_M1027_g N_A_612_71#_c_683_n 0.00184322f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_416 N_A_336_71#_M1027_g N_A_612_71#_c_684_n 0.103228f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_417 N_A_336_71#_M1027_g N_A_612_71#_c_732_n 0.00115219f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_418 N_A_336_71#_c_481_n N_A_393_335#_c_889_n 0.00150571f $X=2 $Y=1.17 $X2=0
+ $Y2=0
cc_419 N_A_336_71#_c_496_n N_A_393_335#_c_889_n 0.00242362f $X=2.165 $Y=1.26
+ $X2=0 $Y2=0
cc_420 N_A_336_71#_c_501_n N_A_393_335#_c_889_n 0.0176029f $X=2.165 $Y=1.17
+ $X2=0 $Y2=0
cc_421 N_A_336_71#_M1010_g N_A_393_335#_M1024_g 0.0123467f $X=2.115 $Y=0.695
+ $X2=0 $Y2=0
cc_422 N_A_336_71#_c_485_n N_A_393_335#_M1024_g 0.00783646f $X=2.84 $Y=0.34
+ $X2=0 $Y2=0
cc_423 N_A_336_71#_c_496_n N_A_393_335#_M1024_g 3.14634e-19 $X=2.165 $Y=1.26
+ $X2=0 $Y2=0
cc_424 N_A_336_71#_c_497_n N_A_393_335#_M1024_g 9.00903e-19 $X=2.165 $Y=1.095
+ $X2=0 $Y2=0
cc_425 N_A_336_71#_c_498_n N_A_393_335#_M1024_g 0.00685868f $X=2.925 $Y=0.34
+ $X2=0 $Y2=0
cc_426 N_A_336_71#_c_501_n N_A_393_335#_M1024_g 0.00981078f $X=2.165 $Y=1.17
+ $X2=0 $Y2=0
cc_427 N_A_336_71#_c_488_n N_A_393_335#_c_893_n 0.0079637f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_428 N_A_336_71#_c_504_n N_A_393_335#_c_893_n 0.00831564f $X=3.985 $Y=2.04
+ $X2=0 $Y2=0
cc_429 N_A_336_71#_c_487_n N_A_393_335#_c_880_n 0.00815795f $X=3.985 $Y=0.925
+ $X2=0 $Y2=0
cc_430 N_A_336_71#_c_488_n N_A_393_335#_c_880_n 0.0106398f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_431 N_A_336_71#_c_489_n N_A_393_335#_c_880_n 0.00201723f $X=5.805 $Y=0.34
+ $X2=0 $Y2=0
cc_432 N_A_336_71#_c_504_n N_A_393_335#_c_880_n 0.0054935f $X=3.985 $Y=2.04
+ $X2=0 $Y2=0
cc_433 N_A_336_71#_c_487_n N_A_393_335#_M1006_g 0.0289516f $X=3.985 $Y=0.925
+ $X2=0 $Y2=0
cc_434 N_A_336_71#_c_488_n N_A_393_335#_M1006_g 0.0156012f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_435 N_A_336_71#_c_488_n N_A_393_335#_c_897_n 0.00822976f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_436 N_A_336_71#_c_487_n N_A_393_335#_c_884_n 0.0135922f $X=3.985 $Y=0.925
+ $X2=0 $Y2=0
cc_437 N_A_336_71#_c_488_n N_A_393_335#_c_884_n 0.0267457f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_438 N_A_336_71#_c_487_n N_A_393_335#_c_885_n 4.19909e-19 $X=3.985 $Y=0.925
+ $X2=0 $Y2=0
cc_439 N_A_336_71#_c_488_n N_A_393_335#_c_885_n 0.00532095f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_440 N_A_336_71#_c_487_n N_A_393_335#_c_886_n 0.0295372f $X=3.985 $Y=0.925
+ $X2=0 $Y2=0
cc_441 N_A_336_71#_c_489_n N_A_393_335#_c_886_n 0.0356462f $X=5.805 $Y=0.34
+ $X2=0 $Y2=0
cc_442 N_A_336_71#_c_490_n N_A_393_335#_c_886_n 0.00587052f $X=5.89 $Y=0.8 $X2=0
+ $Y2=0
cc_443 N_A_336_71#_c_492_n N_A_393_335#_c_886_n 0.00385662f $X=5.975 $Y=0.885
+ $X2=0 $Y2=0
cc_444 N_A_336_71#_c_487_n N_GATE_M1019_g 0.00368199f $X=3.985 $Y=0.925 $X2=0
+ $Y2=0
cc_445 N_A_336_71#_c_489_n N_GATE_M1019_g 0.00971062f $X=5.805 $Y=0.34 $X2=0
+ $Y2=0
cc_446 N_A_336_71#_c_489_n GATE 0.0112188f $X=5.805 $Y=0.34 $X2=0 $Y2=0
cc_447 N_A_336_71#_c_489_n N_GATE_c_1004_n 4.57251e-19 $X=5.805 $Y=0.34 $X2=0
+ $Y2=0
cc_448 N_A_336_71#_c_489_n N_SLEEP_B_M1020_g 0.0106006f $X=5.805 $Y=0.34 $X2=0
+ $Y2=0
cc_449 N_A_336_71#_c_490_n N_SLEEP_B_M1020_g 0.00603882f $X=5.89 $Y=0.8 $X2=0
+ $Y2=0
cc_450 N_A_336_71#_c_492_n N_SLEEP_B_M1020_g 0.00319622f $X=5.975 $Y=0.885 $X2=0
+ $Y2=0
cc_451 N_A_336_71#_c_489_n N_SLEEP_B_M1001_g 0.001894f $X=5.805 $Y=0.34 $X2=0
+ $Y2=0
cc_452 N_A_336_71#_c_490_n N_SLEEP_B_M1001_g 0.00765891f $X=5.89 $Y=0.8 $X2=0
+ $Y2=0
cc_453 N_A_336_71#_c_491_n N_SLEEP_B_M1001_g 0.00903966f $X=6.83 $Y=0.885 $X2=0
+ $Y2=0
cc_454 N_A_336_71#_c_492_n N_SLEEP_B_M1001_g 0.00183577f $X=5.975 $Y=0.885 $X2=0
+ $Y2=0
cc_455 N_A_336_71#_c_490_n N_SLEEP_B_M1003_g 8.00397e-19 $X=5.89 $Y=0.8 $X2=0
+ $Y2=0
cc_456 N_A_336_71#_c_491_n N_SLEEP_B_M1003_g 0.0155734f $X=6.83 $Y=0.885 $X2=0
+ $Y2=0
cc_457 N_A_336_71#_c_493_n N_SLEEP_B_M1003_g 0.00517788f $X=6.915 $Y=0.8 $X2=0
+ $Y2=0
cc_458 N_A_336_71#_c_495_n N_SLEEP_B_M1003_g 6.63377e-19 $X=7 $Y=0.34 $X2=0
+ $Y2=0
cc_459 N_A_336_71#_M1027_g N_SLEEP_B_c_1047_n 0.00830726f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_460 N_A_336_71#_c_491_n N_SLEEP_B_c_1047_n 7.41461e-19 $X=6.83 $Y=0.885 $X2=0
+ $Y2=0
cc_461 N_A_336_71#_c_491_n N_SLEEP_B_c_1048_n 0.00740205f $X=6.83 $Y=0.885 $X2=0
+ $Y2=0
cc_462 N_A_336_71#_c_492_n N_SLEEP_B_c_1048_n 0.00145041f $X=5.975 $Y=0.885
+ $X2=0 $Y2=0
cc_463 N_A_336_71#_c_491_n N_SLEEP_B_M1029_g 0.00485865f $X=6.83 $Y=0.885 $X2=0
+ $Y2=0
cc_464 N_A_336_71#_c_493_n N_SLEEP_B_M1029_g 0.00818401f $X=6.915 $Y=0.8 $X2=0
+ $Y2=0
cc_465 N_A_336_71#_c_494_n N_SLEEP_B_M1029_g 0.00649418f $X=7.59 $Y=0.34 $X2=0
+ $Y2=0
cc_466 N_A_336_71#_c_495_n N_SLEEP_B_M1029_g 0.00190259f $X=7 $Y=0.34 $X2=0
+ $Y2=0
cc_467 N_A_336_71#_c_499_n N_SLEEP_B_M1029_g 6.30759e-19 $X=7.755 $Y=0.34 $X2=0
+ $Y2=0
cc_468 N_A_336_71#_c_500_n N_SLEEP_B_M1029_g 0.00830726f $X=7.755 $Y=0.42 $X2=0
+ $Y2=0
cc_469 N_A_336_71#_c_491_n SLEEP_B 0.0460233f $X=6.83 $Y=0.885 $X2=0 $Y2=0
cc_470 N_A_336_71#_c_492_n SLEEP_B 0.00748683f $X=5.975 $Y=0.885 $X2=0 $Y2=0
cc_471 N_A_336_71#_M1027_g N_A_1324_394#_M1007_g 0.00486868f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_472 N_A_336_71#_c_500_n N_A_1324_394#_M1007_g 0.00327491f $X=7.755 $Y=0.42
+ $X2=0 $Y2=0
cc_473 N_A_336_71#_M1027_g N_A_1324_394#_c_1133_n 0.0102991f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_474 N_A_336_71#_M1027_g N_A_1324_394#_c_1135_n 0.0053446f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_475 N_A_336_71#_M1027_g N_A_1324_394#_c_1156_n 0.00713715f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_476 N_A_336_71#_c_491_n N_A_1324_394#_c_1156_n 0.0060189f $X=6.83 $Y=0.885
+ $X2=0 $Y2=0
cc_477 N_A_336_71#_c_493_n N_A_1324_394#_c_1156_n 0.0148007f $X=6.915 $Y=0.8
+ $X2=0 $Y2=0
cc_478 N_A_336_71#_c_494_n N_A_1324_394#_c_1156_n 0.0192796f $X=7.59 $Y=0.34
+ $X2=0 $Y2=0
cc_479 N_A_336_71#_M1027_g N_A_1324_394#_c_1136_n 0.00529099f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_480 N_A_336_71#_c_491_n N_A_1324_394#_c_1136_n 0.0194466f $X=6.83 $Y=0.885
+ $X2=0 $Y2=0
cc_481 N_A_336_71#_M1027_g N_A_1324_394#_c_1137_n 0.0237075f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_482 N_A_336_71#_c_494_n N_A_1324_394#_c_1137_n 0.00651649f $X=7.59 $Y=0.34
+ $X2=0 $Y2=0
cc_483 N_A_336_71#_c_499_n N_A_1324_394#_c_1137_n 0.0162095f $X=7.755 $Y=0.34
+ $X2=0 $Y2=0
cc_484 N_A_336_71#_c_500_n N_A_1324_394#_c_1137_n 6.19373e-19 $X=7.755 $Y=0.42
+ $X2=0 $Y2=0
cc_485 N_A_336_71#_M1027_g N_A_1324_394#_c_1140_n 0.00281591f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_486 N_A_336_71#_c_491_n N_A_1324_394#_c_1140_n 0.00449564f $X=6.83 $Y=0.885
+ $X2=0 $Y2=0
cc_487 N_A_336_71#_M1010_g N_A_438_97#_c_1226_n 0.00374709f $X=2.115 $Y=0.695
+ $X2=0 $Y2=0
cc_488 N_A_336_71#_c_485_n N_A_438_97#_c_1226_n 0.0253087f $X=2.84 $Y=0.34 $X2=0
+ $Y2=0
cc_489 N_A_336_71#_c_497_n N_A_438_97#_c_1226_n 0.0281427f $X=2.165 $Y=1.095
+ $X2=0 $Y2=0
cc_490 N_A_336_71#_c_485_n N_A_438_97#_c_1227_n 0.0018681f $X=2.84 $Y=0.34 $X2=0
+ $Y2=0
cc_491 N_A_336_71#_c_515_p N_A_438_97#_c_1227_n 0.0355121f $X=3.9 $Y=0.61 $X2=0
+ $Y2=0
cc_492 N_A_336_71#_c_487_n N_A_438_97#_c_1227_n 0.0054524f $X=3.985 $Y=0.925
+ $X2=0 $Y2=0
cc_493 N_A_336_71#_c_488_n N_A_438_97#_c_1227_n 0.00925191f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_494 N_A_336_71#_c_498_n N_A_438_97#_c_1227_n 0.0082023f $X=2.925 $Y=0.34
+ $X2=0 $Y2=0
cc_495 N_A_336_71#_c_488_n N_A_438_97#_c_1238_n 0.00635341f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_496 N_A_336_71#_c_504_n N_A_438_97#_c_1238_n 0.0123605f $X=3.985 $Y=2.04
+ $X2=0 $Y2=0
cc_497 N_A_336_71#_M1033_s N_A_438_97#_c_1239_n 0.00837825f $X=3.66 $Y=1.9 $X2=0
+ $Y2=0
cc_498 N_A_336_71#_c_504_n N_A_438_97#_c_1239_n 0.0238059f $X=3.985 $Y=2.04
+ $X2=0 $Y2=0
cc_499 N_A_336_71#_c_488_n N_A_438_97#_c_1228_n 0.0436331f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_500 N_A_336_71#_c_504_n N_A_438_97#_c_1259_n 0.00642428f $X=3.985 $Y=2.04
+ $X2=0 $Y2=0
cc_501 N_A_336_71#_M1027_g N_A_438_97#_c_1242_n 0.0187782f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_502 N_A_336_71#_M1027_g N_A_438_97#_c_1260_n 0.0261457f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_503 N_A_336_71#_M1027_g N_A_438_97#_c_1288_n 0.00763143f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_504 N_A_336_71#_M1010_g N_A_438_97#_c_1230_n 4.58063e-19 $X=2.115 $Y=0.695
+ $X2=0 $Y2=0
cc_505 N_A_336_71#_c_496_n N_A_438_97#_c_1230_n 0.0257787f $X=2.165 $Y=1.26
+ $X2=0 $Y2=0
cc_506 N_A_336_71#_c_497_n N_A_438_97#_c_1230_n 0.00268801f $X=2.165 $Y=1.095
+ $X2=0 $Y2=0
cc_507 N_A_336_71#_c_501_n N_A_438_97#_c_1230_n 0.0026255f $X=2.165 $Y=1.17
+ $X2=0 $Y2=0
cc_508 N_A_336_71#_c_488_n N_A_438_97#_c_1231_n 0.0127934f $X=3.985 $Y=1.955
+ $X2=0 $Y2=0
cc_509 N_A_336_71#_c_504_n N_A_438_97#_c_1231_n 0.00577892f $X=3.985 $Y=2.04
+ $X2=0 $Y2=0
cc_510 N_A_336_71#_M1027_g N_A_438_97#_c_1245_n 0.00808057f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_511 N_A_336_71#_M1027_g N_A_438_97#_c_1232_n 0.00739365f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_512 N_A_336_71#_M1027_g N_VPWR_c_1501_n 0.00596462f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_513 N_A_336_71#_M1027_g N_VPWR_c_1494_n 0.00815384f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_514 N_A_336_71#_M1002_g N_A_280_97#_c_1614_n 0.00786993f $X=1.755 $Y=0.695
+ $X2=0 $Y2=0
cc_515 N_A_336_71#_M1010_g N_A_280_97#_c_1614_n 4.39797e-19 $X=2.115 $Y=0.695
+ $X2=0 $Y2=0
cc_516 N_A_336_71#_c_497_n N_A_280_97#_c_1614_n 0.0156587f $X=2.165 $Y=1.095
+ $X2=0 $Y2=0
cc_517 N_A_336_71#_M1002_g N_A_280_97#_c_1615_n 0.00618205f $X=1.755 $Y=0.695
+ $X2=0 $Y2=0
cc_518 N_A_336_71#_c_482_n N_A_280_97#_c_1615_n 0.00810302f $X=1.83 $Y=1.17
+ $X2=0 $Y2=0
cc_519 N_A_336_71#_M1010_g N_A_280_97#_c_1615_n 2.92571e-19 $X=2.115 $Y=0.695
+ $X2=0 $Y2=0
cc_520 N_A_336_71#_c_497_n N_A_280_97#_c_1615_n 0.039754f $X=2.165 $Y=1.095
+ $X2=0 $Y2=0
cc_521 N_A_336_71#_c_501_n N_A_280_97#_c_1615_n 0.00163593f $X=2.165 $Y=1.17
+ $X2=0 $Y2=0
cc_522 N_A_336_71#_M1027_g N_KAPWR_c_1666_n 2.4832e-19 $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_523 N_A_336_71#_M1027_g N_KAPWR_c_1663_n 0.00675355f $X=7.7 $Y=2.595 $X2=0
+ $Y2=0
cc_524 N_A_336_71#_c_515_p N_VGND_M1015_d 0.0117984f $X=3.9 $Y=0.61 $X2=0 $Y2=0
cc_525 N_A_336_71#_c_487_n N_VGND_M1015_d 0.00443551f $X=3.985 $Y=0.925 $X2=0
+ $Y2=0
cc_526 N_A_336_71#_c_491_n N_VGND_M1001_d 0.00473966f $X=6.83 $Y=0.885 $X2=0
+ $Y2=0
cc_527 N_A_336_71#_c_489_n N_VGND_c_1800_n 0.0144113f $X=5.805 $Y=0.34 $X2=0
+ $Y2=0
cc_528 N_A_336_71#_c_490_n N_VGND_c_1800_n 0.00915958f $X=5.89 $Y=0.8 $X2=0
+ $Y2=0
cc_529 N_A_336_71#_c_491_n N_VGND_c_1800_n 0.0260356f $X=6.83 $Y=0.885 $X2=0
+ $Y2=0
cc_530 N_A_336_71#_c_493_n N_VGND_c_1800_n 0.00936377f $X=6.915 $Y=0.8 $X2=0
+ $Y2=0
cc_531 N_A_336_71#_c_495_n N_VGND_c_1800_n 0.00909341f $X=7 $Y=0.34 $X2=0 $Y2=0
cc_532 N_A_336_71#_c_515_p N_VGND_c_1804_n 0.0175214f $X=3.9 $Y=0.61 $X2=0 $Y2=0
cc_533 N_A_336_71#_c_487_n N_VGND_c_1804_n 0.014731f $X=3.985 $Y=0.925 $X2=0
+ $Y2=0
cc_534 N_A_336_71#_c_498_n N_VGND_c_1804_n 0.00311108f $X=2.925 $Y=0.34 $X2=0
+ $Y2=0
cc_535 N_A_336_71#_M1002_g N_VGND_c_1805_n 0.00366761f $X=1.755 $Y=0.695 $X2=0
+ $Y2=0
cc_536 N_A_336_71#_M1010_g N_VGND_c_1805_n 7.52598e-19 $X=2.115 $Y=0.695 $X2=0
+ $Y2=0
cc_537 N_A_336_71#_c_485_n N_VGND_c_1805_n 0.0431311f $X=2.84 $Y=0.34 $X2=0
+ $Y2=0
cc_538 N_A_336_71#_c_486_n N_VGND_c_1805_n 0.0121867f $X=2.17 $Y=0.34 $X2=0
+ $Y2=0
cc_539 N_A_336_71#_c_515_p N_VGND_c_1805_n 0.0122771f $X=3.9 $Y=0.61 $X2=0 $Y2=0
cc_540 N_A_336_71#_c_498_n N_VGND_c_1805_n 0.011658f $X=2.925 $Y=0.34 $X2=0
+ $Y2=0
cc_541 N_A_336_71#_c_487_n N_VGND_c_1806_n 0.0280429f $X=3.985 $Y=0.925 $X2=0
+ $Y2=0
cc_542 N_A_336_71#_c_489_n N_VGND_c_1806_n 0.0939863f $X=5.805 $Y=0.34 $X2=0
+ $Y2=0
cc_543 N_A_336_71#_c_494_n N_VGND_c_1808_n 0.037934f $X=7.59 $Y=0.34 $X2=0 $Y2=0
cc_544 N_A_336_71#_c_495_n N_VGND_c_1808_n 0.0122334f $X=7 $Y=0.34 $X2=0 $Y2=0
cc_545 N_A_336_71#_c_499_n N_VGND_c_1808_n 0.0212434f $X=7.755 $Y=0.34 $X2=0
+ $Y2=0
cc_546 N_A_336_71#_c_500_n N_VGND_c_1808_n 0.0025639f $X=7.755 $Y=0.42 $X2=0
+ $Y2=0
cc_547 N_A_336_71#_M1002_g N_VGND_c_1811_n 0.00509887f $X=1.755 $Y=0.695 $X2=0
+ $Y2=0
cc_548 N_A_336_71#_c_485_n N_VGND_c_1811_n 0.0251865f $X=2.84 $Y=0.34 $X2=0
+ $Y2=0
cc_549 N_A_336_71#_c_486_n N_VGND_c_1811_n 0.00660921f $X=2.17 $Y=0.34 $X2=0
+ $Y2=0
cc_550 N_A_336_71#_c_515_p N_VGND_c_1811_n 0.0212981f $X=3.9 $Y=0.61 $X2=0 $Y2=0
cc_551 N_A_336_71#_c_487_n N_VGND_c_1811_n 0.0202776f $X=3.985 $Y=0.925 $X2=0
+ $Y2=0
cc_552 N_A_336_71#_c_489_n N_VGND_c_1811_n 0.0543592f $X=5.805 $Y=0.34 $X2=0
+ $Y2=0
cc_553 N_A_336_71#_c_491_n N_VGND_c_1811_n 0.0190297f $X=6.83 $Y=0.885 $X2=0
+ $Y2=0
cc_554 N_A_336_71#_c_494_n N_VGND_c_1811_n 0.0221702f $X=7.59 $Y=0.34 $X2=0
+ $Y2=0
cc_555 N_A_336_71#_c_495_n N_VGND_c_1811_n 0.00661802f $X=7 $Y=0.34 $X2=0 $Y2=0
cc_556 N_A_336_71#_c_498_n N_VGND_c_1811_n 0.00645941f $X=2.925 $Y=0.34 $X2=0
+ $Y2=0
cc_557 N_A_336_71#_c_499_n N_VGND_c_1811_n 0.0123341f $X=7.755 $Y=0.34 $X2=0
+ $Y2=0
cc_558 N_A_336_71#_c_500_n N_VGND_c_1811_n 6.09111e-19 $X=7.755 $Y=0.42 $X2=0
+ $Y2=0
cc_559 N_A_336_71#_c_498_n A_570_97# 0.00105092f $X=2.925 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_560 N_A_336_71#_c_515_p A_642_97# 0.00243339f $X=3.9 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_561 N_A_336_71#_c_490_n A_1147_97# 0.00398124f $X=5.89 $Y=0.8 $X2=-0.19
+ $Y2=-0.245
cc_562 N_A_336_71#_c_492_n A_1147_97# 0.00149572f $X=5.975 $Y=0.885 $X2=-0.19
+ $Y2=-0.245
cc_563 N_A_336_71#_c_491_n A_1344_97# 0.00100952f $X=6.83 $Y=0.885 $X2=-0.19
+ $Y2=-0.245
cc_564 N_A_336_71#_c_493_n A_1344_97# 0.00349699f $X=6.915 $Y=0.8 $X2=-0.19
+ $Y2=-0.245
cc_565 N_A_336_71#_c_499_n N_A_1624_47#_c_1932_n 0.0153317f $X=7.755 $Y=0.34
+ $X2=0 $Y2=0
cc_566 N_A_336_71#_c_500_n N_A_1624_47#_c_1932_n 0.00236469f $X=7.755 $Y=0.42
+ $X2=0 $Y2=0
cc_567 N_A_336_71#_M1027_g N_A_1624_47#_c_1930_n 0.00298044f $X=7.7 $Y=2.595
+ $X2=0 $Y2=0
cc_568 N_A_336_71#_c_499_n N_A_1624_47#_c_1930_n 0.00297857f $X=7.755 $Y=0.34
+ $X2=0 $Y2=0
cc_569 N_A_336_71#_c_500_n N_A_1624_47#_c_1930_n 4.63853e-19 $X=7.755 $Y=0.42
+ $X2=0 $Y2=0
cc_570 N_A_612_71#_c_692_n N_A_393_335#_M1000_d 0.00854189f $X=6.565 $Y=2.405
+ $X2=0 $Y2=0
cc_571 N_A_612_71#_c_680_n N_A_393_335#_M1021_g 6.04997e-19 $X=3.045 $Y=2.635
+ $X2=0 $Y2=0
cc_572 N_A_612_71#_M1026_g N_A_393_335#_M1024_g 0.0682847f $X=3.135 $Y=0.695
+ $X2=0 $Y2=0
cc_573 N_A_612_71#_c_680_n N_A_393_335#_M1024_g 0.0044277f $X=3.045 $Y=2.635
+ $X2=0 $Y2=0
cc_574 N_A_612_71#_c_682_n N_A_393_335#_M1024_g 0.00145964f $X=3.225 $Y=1.3
+ $X2=0 $Y2=0
cc_575 N_A_612_71#_c_680_n N_A_393_335#_c_893_n 0.0130636f $X=3.045 $Y=2.635
+ $X2=0 $Y2=0
cc_576 N_A_612_71#_c_682_n N_A_393_335#_c_893_n 0.00163889f $X=3.225 $Y=1.3
+ $X2=0 $Y2=0
cc_577 N_A_612_71#_c_686_n N_A_393_335#_c_893_n 0.0337359f $X=3.495 $Y=1.3 $X2=0
+ $Y2=0
cc_578 N_A_612_71#_c_689_n N_A_393_335#_c_880_n 0.0086871f $X=4.6 $Y=2.72 $X2=0
+ $Y2=0
cc_579 N_A_612_71#_c_691_n N_A_393_335#_c_880_n 0.00390453f $X=4.685 $Y=2.635
+ $X2=0 $Y2=0
cc_580 N_A_612_71#_c_693_n N_A_393_335#_c_880_n 0.00152869f $X=4.77 $Y=2.405
+ $X2=0 $Y2=0
cc_581 N_A_612_71#_c_686_n N_A_393_335#_c_880_n 0.0103892f $X=3.495 $Y=1.3 $X2=0
+ $Y2=0
cc_582 N_A_612_71#_M1015_g N_A_393_335#_M1006_g 0.0103892f $X=3.495 $Y=0.695
+ $X2=0 $Y2=0
cc_583 N_A_612_71#_c_691_n N_GATE_M1000_g 0.00381776f $X=4.685 $Y=2.635 $X2=0
+ $Y2=0
cc_584 N_A_612_71#_c_692_n N_GATE_M1000_g 0.0131944f $X=6.565 $Y=2.405 $X2=0
+ $Y2=0
cc_585 N_A_612_71#_c_692_n N_SLEEP_B_M1035_g 0.0120631f $X=6.565 $Y=2.405 $X2=0
+ $Y2=0
cc_586 N_A_612_71#_c_749_p N_SLEEP_B_M1035_g 8.95396e-19 $X=6.65 $Y=2.905 $X2=0
+ $Y2=0
cc_587 N_A_612_71#_c_695_n N_SLEEP_B_M1035_g 4.09993e-19 $X=6.735 $Y=2.99 $X2=0
+ $Y2=0
cc_588 N_A_612_71#_c_692_n N_SLEEP_B_M1023_g 0.0156333f $X=6.565 $Y=2.405 $X2=0
+ $Y2=0
cc_589 N_A_612_71#_c_749_p N_SLEEP_B_M1023_g 0.01388f $X=6.65 $Y=2.905 $X2=0
+ $Y2=0
cc_590 N_A_612_71#_c_695_n N_SLEEP_B_M1023_g 0.0080338f $X=6.735 $Y=2.99 $X2=0
+ $Y2=0
cc_591 N_A_612_71#_c_692_n N_A_1324_394#_M1023_d 0.0039285f $X=6.565 $Y=2.405
+ $X2=0 $Y2=0
cc_592 N_A_612_71#_c_749_p N_A_1324_394#_M1023_d 0.00702999f $X=6.65 $Y=2.905
+ $X2=0 $Y2=0
cc_593 N_A_612_71#_c_694_n N_A_1324_394#_M1023_d 0.00561815f $X=7.93 $Y=2.99
+ $X2=0 $Y2=0
cc_594 N_A_612_71#_M1028_g N_A_1324_394#_M1009_g 0.0427093f $X=8.16 $Y=2.595
+ $X2=0 $Y2=0
cc_595 N_A_612_71#_c_696_n N_A_1324_394#_M1009_g 0.00204915f $X=8.015 $Y=2.32
+ $X2=0 $Y2=0
cc_596 N_A_612_71#_c_729_n N_A_1324_394#_M1009_g 9.12121e-19 $X=8.015 $Y=2.905
+ $X2=0 $Y2=0
cc_597 N_A_612_71#_c_708_n N_A_1324_394#_M1009_g 0.0154866f $X=9.375 $Y=2.405
+ $X2=0 $Y2=0
cc_598 N_A_612_71#_c_683_n N_A_1324_394#_M1009_g 0.00200113f $X=8.2 $Y=1.77
+ $X2=0 $Y2=0
cc_599 N_A_612_71#_c_684_n N_A_1324_394#_M1009_g 0.0208121f $X=8.2 $Y=1.77 $X2=0
+ $Y2=0
cc_600 N_A_612_71#_c_694_n N_A_438_97#_M1027_s 0.00419191f $X=7.93 $Y=2.99 $X2=0
+ $Y2=0
cc_601 N_A_612_71#_c_685_n N_A_438_97#_M1011_g 0.00114528f $X=10.085 $Y=0.465
+ $X2=0 $Y2=0
cc_602 N_A_612_71#_c_681_n N_A_438_97#_M1013_g 0.0158226f $X=10.21 $Y=2.32 $X2=0
+ $Y2=0
cc_603 N_A_612_71#_c_685_n N_A_438_97#_M1013_g 0.00881901f $X=10.085 $Y=0.465
+ $X2=0 $Y2=0
cc_604 N_A_612_71#_c_713_n N_A_438_97#_M1004_g 0.0202968f $X=10.125 $Y=2.405
+ $X2=0 $Y2=0
cc_605 N_A_612_71#_c_718_n N_A_438_97#_M1004_g 0.00947416f $X=9.54 $Y=2.485
+ $X2=0 $Y2=0
cc_606 N_A_612_71#_c_681_n N_A_438_97#_c_1221_n 0.016062f $X=10.21 $Y=2.32 $X2=0
+ $Y2=0
cc_607 N_A_612_71#_c_681_n N_A_438_97#_c_1222_n 0.0292653f $X=10.21 $Y=2.32
+ $X2=0 $Y2=0
cc_608 N_A_612_71#_c_685_n N_A_438_97#_c_1222_n 0.0028563f $X=10.085 $Y=0.465
+ $X2=0 $Y2=0
cc_609 N_A_612_71#_c_685_n N_A_438_97#_M1017_g 0.00275571f $X=10.085 $Y=0.465
+ $X2=0 $Y2=0
cc_610 N_A_612_71#_c_713_n N_A_438_97#_M1034_g 4.22095e-19 $X=10.125 $Y=2.405
+ $X2=0 $Y2=0
cc_611 N_A_612_71#_c_681_n N_A_438_97#_M1034_g 0.00263529f $X=10.21 $Y=2.32
+ $X2=0 $Y2=0
cc_612 N_A_612_71#_c_690_n N_A_438_97#_c_1237_n 0.0123945f $X=3.13 $Y=2.72 $X2=0
+ $Y2=0
cc_613 N_A_612_71#_M1026_g N_A_438_97#_c_1227_n 0.00943164f $X=3.135 $Y=0.695
+ $X2=0 $Y2=0
cc_614 N_A_612_71#_M1015_g N_A_438_97#_c_1227_n 0.0110228f $X=3.495 $Y=0.695
+ $X2=0 $Y2=0
cc_615 N_A_612_71#_c_682_n N_A_438_97#_c_1227_n 0.0313849f $X=3.225 $Y=1.3 $X2=0
+ $Y2=0
cc_616 N_A_612_71#_c_686_n N_A_438_97#_c_1227_n 7.30626e-19 $X=3.495 $Y=1.3
+ $X2=0 $Y2=0
cc_617 N_A_612_71#_c_680_n N_A_438_97#_c_1238_n 0.0373989f $X=3.045 $Y=2.635
+ $X2=0 $Y2=0
cc_618 N_A_612_71#_c_689_n N_A_438_97#_c_1239_n 0.0593484f $X=4.6 $Y=2.72 $X2=0
+ $Y2=0
cc_619 N_A_612_71#_c_693_n N_A_438_97#_c_1239_n 0.0130734f $X=4.77 $Y=2.405
+ $X2=0 $Y2=0
cc_620 N_A_612_71#_c_680_n N_A_438_97#_c_1240_n 0.0143583f $X=3.045 $Y=2.635
+ $X2=0 $Y2=0
cc_621 N_A_612_71#_c_689_n N_A_438_97#_c_1240_n 0.01259f $X=4.6 $Y=2.72 $X2=0
+ $Y2=0
cc_622 N_A_612_71#_M1026_g N_A_438_97#_c_1228_n 4.83662e-19 $X=3.135 $Y=0.695
+ $X2=0 $Y2=0
cc_623 N_A_612_71#_M1015_g N_A_438_97#_c_1228_n 0.00264807f $X=3.495 $Y=0.695
+ $X2=0 $Y2=0
cc_624 N_A_612_71#_c_680_n N_A_438_97#_c_1228_n 0.00658989f $X=3.045 $Y=2.635
+ $X2=0 $Y2=0
cc_625 N_A_612_71#_c_682_n N_A_438_97#_c_1228_n 0.0174543f $X=3.225 $Y=1.3 $X2=0
+ $Y2=0
cc_626 N_A_612_71#_c_686_n N_A_438_97#_c_1228_n 0.010934f $X=3.495 $Y=1.3 $X2=0
+ $Y2=0
cc_627 N_A_612_71#_c_689_n N_A_438_97#_c_1241_n 0.00351116f $X=4.6 $Y=2.72 $X2=0
+ $Y2=0
cc_628 N_A_612_71#_c_692_n N_A_438_97#_c_1241_n 0.118663f $X=6.565 $Y=2.405
+ $X2=0 $Y2=0
cc_629 N_A_612_71#_c_693_n N_A_438_97#_c_1241_n 0.0122461f $X=4.77 $Y=2.405
+ $X2=0 $Y2=0
cc_630 N_A_612_71#_M1028_g N_A_438_97#_c_1242_n 5.71437e-19 $X=8.16 $Y=2.595
+ $X2=0 $Y2=0
cc_631 N_A_612_71#_c_692_n N_A_438_97#_c_1242_n 0.00664512f $X=6.565 $Y=2.405
+ $X2=0 $Y2=0
cc_632 N_A_612_71#_c_749_p N_A_438_97#_c_1242_n 0.00770551f $X=6.65 $Y=2.905
+ $X2=0 $Y2=0
cc_633 N_A_612_71#_c_694_n N_A_438_97#_c_1242_n 0.0315411f $X=7.93 $Y=2.99 $X2=0
+ $Y2=0
cc_634 N_A_612_71#_c_696_n N_A_438_97#_c_1242_n 0.0128736f $X=8.015 $Y=2.32
+ $X2=0 $Y2=0
cc_635 N_A_612_71#_c_729_n N_A_438_97#_c_1242_n 0.018087f $X=8.015 $Y=2.905
+ $X2=0 $Y2=0
cc_636 N_A_612_71#_c_732_n N_A_438_97#_c_1242_n 0.014438f $X=8.015 $Y=2.405
+ $X2=0 $Y2=0
cc_637 N_A_612_71#_c_696_n N_A_438_97#_c_1260_n 0.00312887f $X=8.015 $Y=2.32
+ $X2=0 $Y2=0
cc_638 N_A_612_71#_c_683_n N_A_438_97#_c_1260_n 0.0223623f $X=8.2 $Y=1.77 $X2=0
+ $Y2=0
cc_639 N_A_612_71#_c_684_n N_A_438_97#_c_1260_n 5.18756e-19 $X=8.2 $Y=1.77 $X2=0
+ $Y2=0
cc_640 N_A_612_71#_c_681_n N_A_438_97#_c_1229_n 0.0143217f $X=10.21 $Y=2.32
+ $X2=0 $Y2=0
cc_641 N_A_612_71#_M1026_g N_A_438_97#_c_1230_n 0.00100884f $X=3.135 $Y=0.695
+ $X2=0 $Y2=0
cc_642 N_A_612_71#_c_680_n N_A_438_97#_c_1230_n 0.0862829f $X=3.045 $Y=2.635
+ $X2=0 $Y2=0
cc_643 N_A_612_71#_c_682_n N_A_438_97#_c_1230_n 0.0183011f $X=3.225 $Y=1.3 $X2=0
+ $Y2=0
cc_644 N_A_612_71#_c_686_n N_A_438_97#_c_1230_n 2.37058e-19 $X=3.495 $Y=1.3
+ $X2=0 $Y2=0
cc_645 N_A_612_71#_c_680_n N_A_438_97#_c_1231_n 0.0127936f $X=3.045 $Y=2.635
+ $X2=0 $Y2=0
cc_646 N_A_612_71#_c_682_n N_A_438_97#_c_1231_n 0.00639139f $X=3.225 $Y=1.3
+ $X2=0 $Y2=0
cc_647 N_A_612_71#_c_686_n N_A_438_97#_c_1231_n 0.00233469f $X=3.495 $Y=1.3
+ $X2=0 $Y2=0
cc_648 N_A_612_71#_M1028_g N_A_438_97#_c_1245_n 2.27384e-19 $X=8.16 $Y=2.595
+ $X2=0 $Y2=0
cc_649 N_A_612_71#_c_696_n N_A_438_97#_c_1245_n 0.0120938f $X=8.015 $Y=2.32
+ $X2=0 $Y2=0
cc_650 N_A_612_71#_c_683_n N_A_438_97#_c_1232_n 0.0315967f $X=8.2 $Y=1.77 $X2=0
+ $Y2=0
cc_651 N_A_612_71#_c_684_n N_A_438_97#_c_1232_n 0.00878396f $X=8.2 $Y=1.77 $X2=0
+ $Y2=0
cc_652 N_A_612_71#_c_685_n N_A_2120_55#_c_1446_n 0.0590104f $X=10.085 $Y=0.465
+ $X2=0 $Y2=0
cc_653 N_A_612_71#_c_713_n N_A_2120_55#_c_1451_n 0.0101643f $X=10.125 $Y=2.405
+ $X2=0 $Y2=0
cc_654 N_A_612_71#_c_681_n N_A_2120_55#_c_1451_n 0.0370019f $X=10.21 $Y=2.32
+ $X2=0 $Y2=0
cc_655 N_A_612_71#_c_681_n N_A_2120_55#_c_1449_n 0.0192646f $X=10.21 $Y=2.32
+ $X2=0 $Y2=0
cc_656 N_A_612_71#_c_689_n N_VPWR_M1033_d 0.00741996f $X=4.6 $Y=2.72 $X2=0 $Y2=0
cc_657 N_A_612_71#_c_691_n N_VPWR_M1033_d 0.00206629f $X=4.685 $Y=2.635 $X2=0
+ $Y2=0
cc_658 N_A_612_71#_c_693_n N_VPWR_M1033_d 0.00195856f $X=4.77 $Y=2.405 $X2=0
+ $Y2=0
cc_659 N_A_612_71#_c_689_n N_VPWR_c_1500_n 0.030817f $X=4.6 $Y=2.72 $X2=0 $Y2=0
cc_660 N_A_612_71#_c_690_n N_VPWR_c_1500_n 0.00459235f $X=3.13 $Y=2.72 $X2=0
+ $Y2=0
cc_661 N_A_612_71#_M1028_g N_VPWR_c_1501_n 0.0085571f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_662 N_A_612_71#_c_689_n N_VPWR_c_1501_n 0.00376167f $X=4.6 $Y=2.72 $X2=0
+ $Y2=0
cc_663 N_A_612_71#_c_694_n N_VPWR_c_1501_n 0.0823483f $X=7.93 $Y=2.99 $X2=0
+ $Y2=0
cc_664 N_A_612_71#_c_695_n N_VPWR_c_1501_n 0.0119935f $X=6.735 $Y=2.99 $X2=0
+ $Y2=0
cc_665 N_A_612_71#_c_718_n N_VPWR_c_1501_n 0.0230625f $X=9.54 $Y=2.485 $X2=0
+ $Y2=0
cc_666 N_A_612_71#_M1014_d N_VPWR_c_1494_n 0.00249245f $X=9.285 $Y=2.095 $X2=0
+ $Y2=0
cc_667 N_A_612_71#_M1028_g N_VPWR_c_1494_n 0.00716339f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_668 N_A_612_71#_c_689_n N_VPWR_c_1494_n 0.00461658f $X=4.6 $Y=2.72 $X2=0
+ $Y2=0
cc_669 N_A_612_71#_c_690_n N_VPWR_c_1494_n 5.55225e-19 $X=3.13 $Y=2.72 $X2=0
+ $Y2=0
cc_670 N_A_612_71#_c_694_n N_VPWR_c_1494_n 0.0109778f $X=7.93 $Y=2.99 $X2=0
+ $Y2=0
cc_671 N_A_612_71#_c_695_n N_VPWR_c_1494_n 0.00153814f $X=6.735 $Y=2.99 $X2=0
+ $Y2=0
cc_672 N_A_612_71#_c_718_n N_VPWR_c_1494_n 0.00308223f $X=9.54 $Y=2.485 $X2=0
+ $Y2=0
cc_673 N_A_612_71#_c_689_n N_VPWR_c_1505_n 0.0221823f $X=4.6 $Y=2.72 $X2=0 $Y2=0
cc_674 N_A_612_71#_c_692_n N_KAPWR_M1000_s 0.00334554f $X=6.565 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_675 N_A_612_71#_c_692_n N_KAPWR_M1035_d 0.00529017f $X=6.565 $Y=2.405 $X2=0
+ $Y2=0
cc_676 N_A_612_71#_c_708_n N_KAPWR_M1028_d 0.00401588f $X=9.375 $Y=2.405 $X2=0
+ $Y2=0
cc_677 N_A_612_71#_c_713_n N_KAPWR_M1004_d 0.00555959f $X=10.125 $Y=2.405 $X2=0
+ $Y2=0
cc_678 N_A_612_71#_c_681_n N_KAPWR_M1004_d 0.00612077f $X=10.21 $Y=2.32 $X2=0
+ $Y2=0
cc_679 N_A_612_71#_c_689_n N_KAPWR_c_1660_n 0.0107872f $X=4.6 $Y=2.72 $X2=0
+ $Y2=0
cc_680 N_A_612_71#_c_692_n N_KAPWR_c_1660_n 0.0384825f $X=6.565 $Y=2.405 $X2=0
+ $Y2=0
cc_681 N_A_612_71#_c_692_n N_KAPWR_c_1661_n 0.0261615f $X=6.565 $Y=2.405 $X2=0
+ $Y2=0
cc_682 N_A_612_71#_c_749_p N_KAPWR_c_1661_n 0.0161017f $X=6.65 $Y=2.905 $X2=0
+ $Y2=0
cc_683 N_A_612_71#_c_695_n N_KAPWR_c_1661_n 0.00630246f $X=6.735 $Y=2.99 $X2=0
+ $Y2=0
cc_684 N_A_612_71#_M1028_g N_KAPWR_c_1666_n 0.00506519f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_685 N_A_612_71#_c_694_n N_KAPWR_c_1666_n 0.0130124f $X=7.93 $Y=2.99 $X2=0
+ $Y2=0
cc_686 N_A_612_71#_c_729_n N_KAPWR_c_1666_n 0.0160054f $X=8.015 $Y=2.905 $X2=0
+ $Y2=0
cc_687 N_A_612_71#_c_708_n N_KAPWR_c_1666_n 0.014634f $X=9.375 $Y=2.405 $X2=0
+ $Y2=0
cc_688 N_A_612_71#_c_713_n N_KAPWR_c_1662_n 0.0165226f $X=10.125 $Y=2.405 $X2=0
+ $Y2=0
cc_689 N_A_612_71#_c_718_n N_KAPWR_c_1662_n 0.0163158f $X=9.54 $Y=2.485 $X2=0
+ $Y2=0
cc_690 N_A_612_71#_M1014_d N_KAPWR_c_1663_n 0.00230074f $X=9.285 $Y=2.095 $X2=0
+ $Y2=0
cc_691 N_A_612_71#_M1028_g N_KAPWR_c_1663_n 0.00267193f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_692 N_A_612_71#_c_689_n N_KAPWR_c_1663_n 0.0710112f $X=4.6 $Y=2.72 $X2=0
+ $Y2=0
cc_693 N_A_612_71#_c_690_n N_KAPWR_c_1663_n 0.0155657f $X=3.13 $Y=2.72 $X2=0
+ $Y2=0
cc_694 N_A_612_71#_c_692_n N_KAPWR_c_1663_n 0.0350258f $X=6.565 $Y=2.405 $X2=0
+ $Y2=0
cc_695 N_A_612_71#_c_749_p N_KAPWR_c_1663_n 0.0161479f $X=6.65 $Y=2.905 $X2=0
+ $Y2=0
cc_696 N_A_612_71#_c_694_n N_KAPWR_c_1663_n 0.0410344f $X=7.93 $Y=2.99 $X2=0
+ $Y2=0
cc_697 N_A_612_71#_c_695_n N_KAPWR_c_1663_n 0.00249295f $X=6.735 $Y=2.99 $X2=0
+ $Y2=0
cc_698 N_A_612_71#_c_729_n N_KAPWR_c_1663_n 0.0216791f $X=8.015 $Y=2.905 $X2=0
+ $Y2=0
cc_699 N_A_612_71#_c_708_n N_KAPWR_c_1663_n 0.0401332f $X=9.375 $Y=2.405 $X2=0
+ $Y2=0
cc_700 N_A_612_71#_c_713_n N_KAPWR_c_1663_n 0.0154364f $X=10.125 $Y=2.405 $X2=0
+ $Y2=0
cc_701 N_A_612_71#_c_718_n N_KAPWR_c_1663_n 0.0320764f $X=9.54 $Y=2.485 $X2=0
+ $Y2=0
cc_702 N_A_612_71#_c_694_n A_1565_419# 0.00170171f $X=7.93 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_703 N_A_612_71#_c_696_n A_1565_419# 0.00180385f $X=8.015 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_704 N_A_612_71#_c_729_n A_1565_419# 0.00467504f $X=8.015 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_705 N_A_612_71#_c_732_n A_1565_419# 0.00145348f $X=8.015 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_706 N_A_612_71#_c_708_n A_1765_419# 0.00256529f $X=9.375 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_707 N_A_612_71#_M1026_g N_VGND_c_1805_n 0.00372253f $X=3.135 $Y=0.695 $X2=0
+ $Y2=0
cc_708 N_A_612_71#_M1015_g N_VGND_c_1805_n 0.00372253f $X=3.495 $Y=0.695 $X2=0
+ $Y2=0
cc_709 N_A_612_71#_c_685_n N_VGND_c_1809_n 0.0239268f $X=10.085 $Y=0.465 $X2=0
+ $Y2=0
cc_710 N_A_612_71#_M1013_d N_VGND_c_1811_n 0.00232718f $X=9.945 $Y=0.235 $X2=0
+ $Y2=0
cc_711 N_A_612_71#_M1026_g N_VGND_c_1811_n 0.00509887f $X=3.135 $Y=0.695 $X2=0
+ $Y2=0
cc_712 N_A_612_71#_M1015_g N_VGND_c_1811_n 0.00509887f $X=3.495 $Y=0.695 $X2=0
+ $Y2=0
cc_713 N_A_612_71#_c_685_n N_VGND_c_1811_n 0.0142953f $X=10.085 $Y=0.465 $X2=0
+ $Y2=0
cc_714 N_A_612_71#_c_681_n N_A_1624_47#_c_1931_n 7.69019e-19 $X=10.21 $Y=2.32
+ $X2=0 $Y2=0
cc_715 N_A_612_71#_c_685_n N_A_1624_47#_c_1931_n 0.0140597f $X=10.085 $Y=0.465
+ $X2=0 $Y2=0
cc_716 N_A_393_335#_c_880_n N_GATE_M1000_g 0.008872f $X=4.135 $Y=1.825 $X2=0
+ $Y2=0
cc_717 N_A_393_335#_c_882_n N_GATE_M1000_g 0.00517994f $X=4.625 $Y=1.64 $X2=0
+ $Y2=0
cc_718 N_A_393_335#_c_883_n N_GATE_M1000_g 0.0122445f $X=5.57 $Y=1.725 $X2=0
+ $Y2=0
cc_719 N_A_393_335#_c_885_n N_GATE_M1019_g 0.0049454f $X=4.625 $Y=1.105 $X2=0
+ $Y2=0
cc_720 N_A_393_335#_c_886_n N_GATE_M1019_g 0.00683718f $X=5.055 $Y=0.715 $X2=0
+ $Y2=0
cc_721 N_A_393_335#_c_880_n GATE 3.05276e-19 $X=4.135 $Y=1.825 $X2=0 $Y2=0
cc_722 N_A_393_335#_c_883_n GATE 0.0346198f $X=5.57 $Y=1.725 $X2=0 $Y2=0
cc_723 N_A_393_335#_c_885_n GATE 0.027941f $X=4.625 $Y=1.105 $X2=0 $Y2=0
cc_724 N_A_393_335#_c_886_n GATE 0.0137304f $X=5.055 $Y=0.715 $X2=0 $Y2=0
cc_725 N_A_393_335#_c_880_n N_GATE_c_1004_n 0.0111281f $X=4.135 $Y=1.825 $X2=0
+ $Y2=0
cc_726 N_A_393_335#_c_883_n N_GATE_c_1004_n 0.00401567f $X=5.57 $Y=1.725 $X2=0
+ $Y2=0
cc_727 N_A_393_335#_c_885_n N_GATE_c_1004_n 0.0013302f $X=4.625 $Y=1.105 $X2=0
+ $Y2=0
cc_728 N_A_393_335#_c_886_n N_GATE_c_1004_n 0.0035342f $X=5.055 $Y=0.715 $X2=0
+ $Y2=0
cc_729 N_A_393_335#_c_886_n N_SLEEP_B_M1020_g 9.54032e-19 $X=5.055 $Y=0.715
+ $X2=0 $Y2=0
cc_730 N_A_393_335#_c_883_n N_SLEEP_B_M1035_g 0.00552863f $X=5.57 $Y=1.725 $X2=0
+ $Y2=0
cc_731 N_A_393_335#_c_883_n N_SLEEP_B_c_1048_n 0.0036751f $X=5.57 $Y=1.725 $X2=0
+ $Y2=0
cc_732 N_A_393_335#_M1018_g N_A_438_97#_c_1236_n 0.00193636f $X=2.04 $Y=2.755
+ $X2=0 $Y2=0
cc_733 N_A_393_335#_M1021_g N_A_438_97#_c_1236_n 0.00587306f $X=2.4 $Y=2.755
+ $X2=0 $Y2=0
cc_734 N_A_393_335#_M1021_g N_A_438_97#_c_1237_n 0.00970222f $X=2.4 $Y=2.755
+ $X2=0 $Y2=0
cc_735 N_A_393_335#_M1024_g N_A_438_97#_c_1226_n 0.00555448f $X=2.775 $Y=0.695
+ $X2=0 $Y2=0
cc_736 N_A_393_335#_M1024_g N_A_438_97#_c_1227_n 0.00708869f $X=2.775 $Y=0.695
+ $X2=0 $Y2=0
cc_737 N_A_393_335#_c_893_n N_A_438_97#_c_1227_n 6.77846e-19 $X=4.06 $Y=1.75
+ $X2=0 $Y2=0
cc_738 N_A_393_335#_c_893_n N_A_438_97#_c_1238_n 0.00653988f $X=4.06 $Y=1.75
+ $X2=0 $Y2=0
cc_739 N_A_393_335#_c_880_n N_A_438_97#_c_1238_n 0.0047896f $X=4.135 $Y=1.825
+ $X2=0 $Y2=0
cc_740 N_A_393_335#_c_893_n N_A_438_97#_c_1239_n 0.00299511f $X=4.06 $Y=1.75
+ $X2=0 $Y2=0
cc_741 N_A_393_335#_c_880_n N_A_438_97#_c_1239_n 0.0139067f $X=4.135 $Y=1.825
+ $X2=0 $Y2=0
cc_742 N_A_393_335#_c_893_n N_A_438_97#_c_1228_n 0.00139136f $X=4.06 $Y=1.75
+ $X2=0 $Y2=0
cc_743 N_A_393_335#_M1000_d N_A_438_97#_c_1241_n 0.00579882f $X=5.315 $Y=2.33
+ $X2=0 $Y2=0
cc_744 N_A_393_335#_c_880_n N_A_438_97#_c_1241_n 0.00724431f $X=4.135 $Y=1.825
+ $X2=0 $Y2=0
cc_745 N_A_393_335#_c_897_n N_A_438_97#_c_1241_n 0.0314028f $X=4.875 $Y=1.725
+ $X2=0 $Y2=0
cc_746 N_A_393_335#_c_883_n N_A_438_97#_c_1241_n 0.0549492f $X=5.57 $Y=1.725
+ $X2=0 $Y2=0
cc_747 N_A_393_335#_c_880_n N_A_438_97#_c_1259_n 0.00922054f $X=4.135 $Y=1.825
+ $X2=0 $Y2=0
cc_748 N_A_393_335#_c_897_n N_A_438_97#_c_1259_n 0.00384769f $X=4.875 $Y=1.725
+ $X2=0 $Y2=0
cc_749 N_A_393_335#_M1021_g N_A_438_97#_c_1230_n 0.0172336f $X=2.4 $Y=2.755
+ $X2=0 $Y2=0
cc_750 N_A_393_335#_c_891_n N_A_438_97#_c_1230_n 0.014793f $X=2.7 $Y=1.75 $X2=0
+ $Y2=0
cc_751 N_A_393_335#_M1024_g N_A_438_97#_c_1230_n 0.019089f $X=2.775 $Y=0.695
+ $X2=0 $Y2=0
cc_752 N_A_393_335#_c_896_n N_A_438_97#_c_1230_n 0.00524843f $X=2.775 $Y=1.75
+ $X2=0 $Y2=0
cc_753 N_A_393_335#_c_893_n N_A_438_97#_c_1231_n 0.0140755f $X=4.06 $Y=1.75
+ $X2=0 $Y2=0
cc_754 N_A_393_335#_M1018_g N_VPWR_c_1500_n 0.00529818f $X=2.04 $Y=2.755 $X2=0
+ $Y2=0
cc_755 N_A_393_335#_M1021_g N_VPWR_c_1500_n 0.00529818f $X=2.4 $Y=2.755 $X2=0
+ $Y2=0
cc_756 N_A_393_335#_c_880_n N_VPWR_c_1500_n 5.53268e-19 $X=4.135 $Y=1.825 $X2=0
+ $Y2=0
cc_757 N_A_393_335#_M1018_g N_VPWR_c_1494_n 0.00492443f $X=2.04 $Y=2.755 $X2=0
+ $Y2=0
cc_758 N_A_393_335#_M1021_g N_VPWR_c_1494_n 0.00610075f $X=2.4 $Y=2.755 $X2=0
+ $Y2=0
cc_759 N_A_393_335#_M1018_g N_A_280_97#_c_1616_n 0.00472269f $X=2.04 $Y=2.755
+ $X2=0 $Y2=0
cc_760 N_A_393_335#_M1021_g N_A_280_97#_c_1616_n 0.00193636f $X=2.4 $Y=2.755
+ $X2=0 $Y2=0
cc_761 N_A_393_335#_M1018_g N_A_280_97#_c_1617_n 0.00855185f $X=2.04 $Y=2.755
+ $X2=0 $Y2=0
cc_762 N_A_393_335#_c_889_n N_A_280_97#_c_1615_n 0.00818565f $X=2.115 $Y=1.75
+ $X2=0 $Y2=0
cc_763 N_A_393_335#_M1000_d N_KAPWR_c_1660_n 0.00731249f $X=5.315 $Y=2.33 $X2=0
+ $Y2=0
cc_764 N_A_393_335#_M1000_d N_KAPWR_c_1663_n 0.00294035f $X=5.315 $Y=2.33 $X2=0
+ $Y2=0
cc_765 N_A_393_335#_M1018_g N_KAPWR_c_1663_n 0.00781454f $X=2.04 $Y=2.755 $X2=0
+ $Y2=0
cc_766 N_A_393_335#_M1021_g N_KAPWR_c_1663_n 0.00781454f $X=2.4 $Y=2.755 $X2=0
+ $Y2=0
cc_767 N_A_393_335#_M1024_g N_VGND_c_1805_n 7.30437e-19 $X=2.775 $Y=0.695 $X2=0
+ $Y2=0
cc_768 N_A_393_335#_M1006_g N_VGND_c_1806_n 0.00322375f $X=4.155 $Y=0.695 $X2=0
+ $Y2=0
cc_769 N_A_393_335#_M1006_g N_VGND_c_1811_n 0.00424906f $X=4.155 $Y=0.695 $X2=0
+ $Y2=0
cc_770 N_GATE_M1019_g N_SLEEP_B_M1020_g 0.0388178f $X=5.27 $Y=0.695 $X2=0 $Y2=0
cc_771 GATE N_SLEEP_B_M1020_g 0.00289335f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_772 N_GATE_c_1004_n N_SLEEP_B_M1020_g 0.0129767f $X=5.21 $Y=1.255 $X2=0 $Y2=0
cc_773 GATE N_SLEEP_B_M1001_g 2.51836e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_774 N_GATE_M1000_g N_SLEEP_B_c_1048_n 0.0404391f $X=5.24 $Y=2.65 $X2=0 $Y2=0
cc_775 GATE N_SLEEP_B_c_1048_n 0.00697257f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_776 N_GATE_c_1004_n N_SLEEP_B_c_1048_n 0.00300408f $X=5.21 $Y=1.255 $X2=0
+ $Y2=0
cc_777 N_GATE_M1000_g SLEEP_B 2.31646e-19 $X=5.24 $Y=2.65 $X2=0 $Y2=0
cc_778 GATE SLEEP_B 0.0177025f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_779 N_GATE_M1000_g N_A_438_97#_c_1241_n 0.0125818f $X=5.24 $Y=2.65 $X2=0
+ $Y2=0
cc_780 N_GATE_M1000_g N_VPWR_c_1501_n 0.00295805f $X=5.24 $Y=2.65 $X2=0 $Y2=0
cc_781 N_GATE_M1000_g N_VPWR_c_1494_n 0.00333824f $X=5.24 $Y=2.65 $X2=0 $Y2=0
cc_782 N_GATE_M1000_g N_VPWR_c_1505_n 0.00271737f $X=5.24 $Y=2.65 $X2=0 $Y2=0
cc_783 N_GATE_M1000_g N_KAPWR_c_1660_n 0.0133229f $X=5.24 $Y=2.65 $X2=0 $Y2=0
cc_784 N_GATE_M1000_g N_KAPWR_c_1661_n 3.58969e-19 $X=5.24 $Y=2.65 $X2=0 $Y2=0
cc_785 N_GATE_M1019_g N_VGND_c_1806_n 7.35405e-19 $X=5.27 $Y=0.695 $X2=0 $Y2=0
cc_786 N_SLEEP_B_M1023_g N_A_1324_394#_c_1135_n 0.00564979f $X=6.495 $Y=2.47
+ $X2=0 $Y2=0
cc_787 N_SLEEP_B_c_1048_n N_A_1324_394#_c_1135_n 0.00452499f $X=6.72 $Y=1.215
+ $X2=0 $Y2=0
cc_788 SLEEP_B N_A_1324_394#_c_1135_n 0.00884506f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_789 N_SLEEP_B_M1029_g N_A_1324_394#_c_1156_n 0.00256406f $X=7.005 $Y=0.695
+ $X2=0 $Y2=0
cc_790 N_SLEEP_B_c_1047_n N_A_1324_394#_c_1136_n 0.0175872f $X=6.93 $Y=1.215
+ $X2=0 $Y2=0
cc_791 N_SLEEP_B_c_1048_n N_A_1324_394#_c_1136_n 5.86572e-19 $X=6.72 $Y=1.215
+ $X2=0 $Y2=0
cc_792 N_SLEEP_B_M1029_g N_A_1324_394#_c_1136_n 0.00647688f $X=7.005 $Y=0.695
+ $X2=0 $Y2=0
cc_793 SLEEP_B N_A_1324_394#_c_1136_n 0.00967384f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_794 N_SLEEP_B_M1023_g N_A_1324_394#_c_1140_n 0.00719436f $X=6.495 $Y=2.47
+ $X2=0 $Y2=0
cc_795 N_SLEEP_B_c_1047_n N_A_1324_394#_c_1140_n 0.00408067f $X=6.93 $Y=1.215
+ $X2=0 $Y2=0
cc_796 N_SLEEP_B_c_1048_n N_A_1324_394#_c_1140_n 3.12848e-19 $X=6.72 $Y=1.215
+ $X2=0 $Y2=0
cc_797 N_SLEEP_B_M1035_g N_A_438_97#_c_1241_n 0.0130671f $X=5.9 $Y=2.65 $X2=0
+ $Y2=0
cc_798 N_SLEEP_B_M1023_g N_A_438_97#_c_1241_n 0.0186832f $X=6.495 $Y=2.47 $X2=0
+ $Y2=0
cc_799 N_SLEEP_B_c_1047_n N_A_438_97#_c_1241_n 2.09814e-19 $X=6.93 $Y=1.215
+ $X2=0 $Y2=0
cc_800 N_SLEEP_B_c_1048_n N_A_438_97#_c_1241_n 0.00760096f $X=6.72 $Y=1.215
+ $X2=0 $Y2=0
cc_801 SLEEP_B N_A_438_97#_c_1241_n 0.012396f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_802 N_SLEEP_B_M1023_g N_A_438_97#_c_1242_n 0.00629125f $X=6.495 $Y=2.47 $X2=0
+ $Y2=0
cc_803 N_SLEEP_B_M1035_g N_VPWR_c_1501_n 0.0036535f $X=5.9 $Y=2.65 $X2=0 $Y2=0
cc_804 N_SLEEP_B_M1023_g N_VPWR_c_1501_n 0.00685476f $X=6.495 $Y=2.47 $X2=0
+ $Y2=0
cc_805 N_SLEEP_B_M1035_g N_VPWR_c_1494_n 0.00334423f $X=5.9 $Y=2.65 $X2=0 $Y2=0
cc_806 N_SLEEP_B_M1023_g N_VPWR_c_1494_n 0.00562956f $X=6.495 $Y=2.47 $X2=0
+ $Y2=0
cc_807 N_SLEEP_B_M1035_g N_KAPWR_c_1660_n 0.00244001f $X=5.9 $Y=2.65 $X2=0 $Y2=0
cc_808 N_SLEEP_B_M1035_g N_KAPWR_c_1661_n 0.0115429f $X=5.9 $Y=2.65 $X2=0 $Y2=0
cc_809 N_SLEEP_B_M1023_g N_KAPWR_c_1661_n 0.00444653f $X=6.495 $Y=2.47 $X2=0
+ $Y2=0
cc_810 N_SLEEP_B_M1035_g N_KAPWR_c_1663_n 0.00359064f $X=5.9 $Y=2.65 $X2=0 $Y2=0
cc_811 N_SLEEP_B_M1023_g N_KAPWR_c_1663_n 0.00265631f $X=6.495 $Y=2.47 $X2=0
+ $Y2=0
cc_812 N_SLEEP_B_M1001_g N_VGND_c_1800_n 0.00223712f $X=6.02 $Y=0.695 $X2=0
+ $Y2=0
cc_813 N_SLEEP_B_M1003_g N_VGND_c_1800_n 0.00326f $X=6.645 $Y=0.695 $X2=0 $Y2=0
cc_814 N_SLEEP_B_M1020_g N_VGND_c_1806_n 7.35405e-19 $X=5.66 $Y=0.695 $X2=0
+ $Y2=0
cc_815 N_SLEEP_B_M1001_g N_VGND_c_1806_n 0.0041251f $X=6.02 $Y=0.695 $X2=0 $Y2=0
cc_816 N_SLEEP_B_M1003_g N_VGND_c_1808_n 0.00497279f $X=6.645 $Y=0.695 $X2=0
+ $Y2=0
cc_817 N_SLEEP_B_M1029_g N_VGND_c_1808_n 7.53033e-19 $X=7.005 $Y=0.695 $X2=0
+ $Y2=0
cc_818 N_SLEEP_B_M1001_g N_VGND_c_1811_n 0.00407909f $X=6.02 $Y=0.695 $X2=0
+ $Y2=0
cc_819 N_SLEEP_B_M1003_g N_VGND_c_1811_n 0.00509887f $X=6.645 $Y=0.695 $X2=0
+ $Y2=0
cc_820 N_A_1324_394#_M1023_d N_A_438_97#_c_1241_n 0.0100498f $X=6.62 $Y=1.97
+ $X2=0 $Y2=0
cc_821 N_A_1324_394#_c_1136_n N_A_438_97#_c_1241_n 0.00533101f $X=7.42 $Y=1.005
+ $X2=0 $Y2=0
cc_822 N_A_1324_394#_c_1140_n N_A_438_97#_c_1241_n 0.0210478f $X=6.875 $Y=1.725
+ $X2=0 $Y2=0
cc_823 N_A_1324_394#_c_1135_n N_A_438_97#_c_1260_n 0.00486929f $X=6.955 $Y=1.64
+ $X2=0 $Y2=0
cc_824 N_A_1324_394#_c_1140_n N_A_438_97#_c_1260_n 0.00527768f $X=6.875 $Y=1.725
+ $X2=0 $Y2=0
cc_825 N_A_1324_394#_c_1135_n N_A_438_97#_c_1288_n 0.00537905f $X=6.955 $Y=1.64
+ $X2=0 $Y2=0
cc_826 N_A_1324_394#_c_1136_n N_A_438_97#_c_1288_n 4.38412e-19 $X=7.42 $Y=1.005
+ $X2=0 $Y2=0
cc_827 N_A_1324_394#_c_1137_n N_A_438_97#_c_1288_n 0.0133403f $X=8.55 $Y=1.005
+ $X2=0 $Y2=0
cc_828 N_A_1324_394#_c_1136_n N_A_438_97#_c_1245_n 0.00383156f $X=7.42 $Y=1.005
+ $X2=0 $Y2=0
cc_829 N_A_1324_394#_c_1133_n N_A_438_97#_c_1232_n 0.00601522f $X=8.7 $Y=1.305
+ $X2=0 $Y2=0
cc_830 N_A_1324_394#_M1009_g N_A_438_97#_c_1232_n 0.0191462f $X=8.7 $Y=2.595
+ $X2=0 $Y2=0
cc_831 N_A_1324_394#_c_1137_n N_A_438_97#_c_1232_n 0.0719246f $X=8.55 $Y=1.005
+ $X2=0 $Y2=0
cc_832 N_A_1324_394#_c_1133_n N_A_438_97#_c_1233_n 0.00606197f $X=8.7 $Y=1.305
+ $X2=0 $Y2=0
cc_833 N_A_1324_394#_c_1137_n N_A_438_97#_c_1233_n 0.00873702f $X=8.55 $Y=1.005
+ $X2=0 $Y2=0
cc_834 N_A_1324_394#_M1009_g N_VPWR_c_1501_n 0.00939206f $X=8.7 $Y=2.595 $X2=0
+ $Y2=0
cc_835 N_A_1324_394#_M1009_g N_VPWR_c_1494_n 0.0072846f $X=8.7 $Y=2.595 $X2=0
+ $Y2=0
cc_836 N_A_1324_394#_M1009_g N_KAPWR_c_1666_n 0.00982282f $X=8.7 $Y=2.595 $X2=0
+ $Y2=0
cc_837 N_A_1324_394#_M1023_d N_KAPWR_c_1663_n 0.00450206f $X=6.62 $Y=1.97 $X2=0
+ $Y2=0
cc_838 N_A_1324_394#_M1009_g N_KAPWR_c_1663_n 0.00639118f $X=8.7 $Y=2.595 $X2=0
+ $Y2=0
cc_839 N_A_1324_394#_M1007_g N_VGND_c_1808_n 0.0040248f $X=8.48 $Y=0.445 $X2=0
+ $Y2=0
cc_840 N_A_1324_394#_M1007_g N_VGND_c_1811_n 0.0073925f $X=8.48 $Y=0.445 $X2=0
+ $Y2=0
cc_841 N_A_1324_394#_M1007_g N_VGND_c_1812_n 0.00392695f $X=8.48 $Y=0.445 $X2=0
+ $Y2=0
cc_842 N_A_1324_394#_M1007_g N_A_1624_47#_c_1932_n 0.00495662f $X=8.48 $Y=0.445
+ $X2=0 $Y2=0
cc_843 N_A_1324_394#_M1007_g N_A_1624_47#_c_1929_n 0.00883768f $X=8.48 $Y=0.445
+ $X2=0 $Y2=0
cc_844 N_A_1324_394#_c_1133_n N_A_1624_47#_c_1929_n 0.00686592f $X=8.7 $Y=1.305
+ $X2=0 $Y2=0
cc_845 N_A_1324_394#_c_1137_n N_A_1624_47#_c_1929_n 0.0205336f $X=8.55 $Y=1.005
+ $X2=0 $Y2=0
cc_846 N_A_1324_394#_M1007_g N_A_1624_47#_c_1930_n 0.00143065f $X=8.48 $Y=0.445
+ $X2=0 $Y2=0
cc_847 N_A_1324_394#_c_1133_n N_A_1624_47#_c_1930_n 5.13598e-19 $X=8.7 $Y=1.305
+ $X2=0 $Y2=0
cc_848 N_A_1324_394#_c_1137_n N_A_1624_47#_c_1930_n 0.0207616f $X=8.55 $Y=1.005
+ $X2=0 $Y2=0
cc_849 N_A_1324_394#_M1007_g N_A_1624_47#_c_1931_n 8.64736e-19 $X=8.48 $Y=0.445
+ $X2=0 $Y2=0
cc_850 N_A_438_97#_M1017_g N_A_2120_55#_M1016_g 0.0218676f $X=10.96 $Y=0.485
+ $X2=0 $Y2=0
cc_851 N_A_438_97#_M1034_g N_A_2120_55#_M1012_g 0.0149717f $X=10.96 $Y=2.155
+ $X2=0 $Y2=0
cc_852 N_A_438_97#_M1013_g N_A_2120_55#_c_1446_n 8.19022e-19 $X=9.87 $Y=0.445
+ $X2=0 $Y2=0
cc_853 N_A_438_97#_c_1221_n N_A_2120_55#_c_1446_n 0.011239f $X=10.885 $Y=1.26
+ $X2=0 $Y2=0
cc_854 N_A_438_97#_M1017_g N_A_2120_55#_c_1446_n 0.0235315f $X=10.96 $Y=0.485
+ $X2=0 $Y2=0
cc_855 N_A_438_97#_c_1225_n N_A_2120_55#_c_1446_n 0.00258935f $X=10.96 $Y=1.26
+ $X2=0 $Y2=0
cc_856 N_A_438_97#_M1004_g N_A_2120_55#_c_1451_n 0.00215709f $X=9.92 $Y=2.595
+ $X2=0 $Y2=0
cc_857 N_A_438_97#_M1034_g N_A_2120_55#_c_1451_n 0.0155216f $X=10.96 $Y=2.155
+ $X2=0 $Y2=0
cc_858 N_A_438_97#_M1034_g N_A_2120_55#_c_1447_n 0.0122767f $X=10.96 $Y=2.155
+ $X2=0 $Y2=0
cc_859 N_A_438_97#_c_1225_n N_A_2120_55#_c_1447_n 0.00631774f $X=10.96 $Y=1.26
+ $X2=0 $Y2=0
cc_860 N_A_438_97#_c_1225_n N_A_2120_55#_c_1448_n 0.0213254f $X=10.96 $Y=1.26
+ $X2=0 $Y2=0
cc_861 N_A_438_97#_c_1221_n N_A_2120_55#_c_1449_n 0.00613583f $X=10.885 $Y=1.26
+ $X2=0 $Y2=0
cc_862 N_A_438_97#_M1034_g N_A_2120_55#_c_1449_n 0.00697028f $X=10.96 $Y=2.155
+ $X2=0 $Y2=0
cc_863 N_A_438_97#_c_1239_n N_VPWR_M1033_d 0.00475226f $X=4.26 $Y=2.38 $X2=0
+ $Y2=0
cc_864 N_A_438_97#_c_1406_p N_VPWR_M1033_d 0.00576493f $X=4.345 $Y=2.295 $X2=0
+ $Y2=0
cc_865 N_A_438_97#_c_1241_n N_VPWR_M1033_d 0.0053941f $X=7.27 $Y=2.065 $X2=0
+ $Y2=0
cc_866 N_A_438_97#_c_1259_n N_VPWR_M1033_d 0.0033171f $X=4.43 $Y=2.065 $X2=0
+ $Y2=0
cc_867 N_A_438_97#_M1034_g N_VPWR_c_1499_n 0.00890208f $X=10.96 $Y=2.155 $X2=0
+ $Y2=0
cc_868 N_A_438_97#_c_1237_n N_VPWR_c_1500_n 0.0210483f $X=2.615 $Y=2.745 $X2=0
+ $Y2=0
cc_869 N_A_438_97#_M1004_g N_VPWR_c_1501_n 0.00937723f $X=9.92 $Y=2.595 $X2=0
+ $Y2=0
cc_870 N_A_438_97#_M1034_g N_VPWR_c_1501_n 0.00312414f $X=10.96 $Y=2.155 $X2=0
+ $Y2=0
cc_871 N_A_438_97#_M1027_s N_VPWR_c_1494_n 0.00119816f $X=7.29 $Y=2.095 $X2=0
+ $Y2=0
cc_872 N_A_438_97#_M1004_g N_VPWR_c_1494_n 0.00934125f $X=9.92 $Y=2.595 $X2=0
+ $Y2=0
cc_873 N_A_438_97#_c_1237_n N_VPWR_c_1494_n 0.00305483f $X=2.615 $Y=2.745 $X2=0
+ $Y2=0
cc_874 N_A_438_97#_c_1236_n N_A_280_97#_c_1616_n 0.00894451f $X=2.615 $Y=2.58
+ $X2=0 $Y2=0
cc_875 N_A_438_97#_c_1237_n N_A_280_97#_c_1617_n 0.00894451f $X=2.615 $Y=2.745
+ $X2=0 $Y2=0
cc_876 N_A_438_97#_c_1230_n N_A_280_97#_c_1615_n 0.0266129f $X=2.615 $Y=2.415
+ $X2=0 $Y2=0
cc_877 N_A_438_97#_c_1241_n N_KAPWR_M1035_d 0.00531266f $X=7.27 $Y=2.065 $X2=0
+ $Y2=0
cc_878 N_A_438_97#_M1004_g N_KAPWR_c_1662_n 0.0067579f $X=9.92 $Y=2.595 $X2=0
+ $Y2=0
cc_879 N_A_438_97#_M1004_g N_KAPWR_c_1663_n 0.00758846f $X=9.92 $Y=2.595 $X2=0
+ $Y2=0
cc_880 N_A_438_97#_M1034_g N_KAPWR_c_1663_n 0.00480838f $X=10.96 $Y=2.155 $X2=0
+ $Y2=0
cc_881 N_A_438_97#_c_1237_n N_KAPWR_c_1663_n 0.0422338f $X=2.615 $Y=2.745 $X2=0
+ $Y2=0
cc_882 N_A_438_97#_c_1239_n N_KAPWR_c_1663_n 0.00655371f $X=4.26 $Y=2.38 $X2=0
+ $Y2=0
cc_883 N_A_438_97#_c_1240_n N_KAPWR_c_1663_n 0.00129886f $X=3.47 $Y=2.38 $X2=0
+ $Y2=0
cc_884 N_A_438_97#_c_1241_n N_KAPWR_c_1663_n 0.0209708f $X=7.27 $Y=2.065 $X2=0
+ $Y2=0
cc_885 N_A_438_97#_c_1242_n N_KAPWR_c_1663_n 0.0373154f $X=7.435 $Y=2.405 $X2=0
+ $Y2=0
cc_886 N_A_438_97#_M1017_g N_Q_c_1776_n 6.86967e-19 $X=10.96 $Y=0.485 $X2=0
+ $Y2=0
cc_887 N_A_438_97#_c_1227_n N_VGND_M1015_d 0.00150181f $X=3.56 $Y=0.95 $X2=0
+ $Y2=0
cc_888 N_A_438_97#_M1017_g N_VGND_c_1801_n 0.0085758f $X=10.96 $Y=0.485 $X2=0
+ $Y2=0
cc_889 N_A_438_97#_M1011_g N_VGND_c_1809_n 0.0055654f $X=9.51 $Y=0.445 $X2=0
+ $Y2=0
cc_890 N_A_438_97#_M1013_g N_VGND_c_1809_n 0.0054895f $X=9.87 $Y=0.445 $X2=0
+ $Y2=0
cc_891 N_A_438_97#_M1017_g N_VGND_c_1809_n 0.00511358f $X=10.96 $Y=0.485 $X2=0
+ $Y2=0
cc_892 N_A_438_97#_M1011_g N_VGND_c_1811_n 0.0101191f $X=9.51 $Y=0.445 $X2=0
+ $Y2=0
cc_893 N_A_438_97#_M1013_g N_VGND_c_1811_n 0.0112803f $X=9.87 $Y=0.445 $X2=0
+ $Y2=0
cc_894 N_A_438_97#_M1017_g N_VGND_c_1811_n 0.0108382f $X=10.96 $Y=0.485 $X2=0
+ $Y2=0
cc_895 N_A_438_97#_c_1227_n A_570_97# 0.0010205f $X=3.56 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_896 N_A_438_97#_c_1227_n A_642_97# 0.00102299f $X=3.56 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_897 N_A_438_97#_c_1232_n N_A_1624_47#_c_1929_n 0.00489506f $X=8.885 $Y=1.255
+ $X2=0 $Y2=0
cc_898 N_A_438_97#_c_1233_n N_A_1624_47#_c_1929_n 0.0113083f $X=9.055 $Y=1.255
+ $X2=0 $Y2=0
cc_899 N_A_438_97#_M1011_g N_A_1624_47#_c_1931_n 0.00845674f $X=9.51 $Y=0.445
+ $X2=0 $Y2=0
cc_900 N_A_438_97#_M1013_g N_A_1624_47#_c_1931_n 0.00122391f $X=9.87 $Y=0.445
+ $X2=0 $Y2=0
cc_901 N_A_438_97#_c_1229_n N_A_1624_47#_c_1931_n 0.0172111f $X=9.6 $Y=1.2 $X2=0
+ $Y2=0
cc_902 N_A_2120_55#_M1012_g N_VPWR_c_1499_n 0.0071691f $X=11.505 $Y=2.465 $X2=0
+ $Y2=0
cc_903 N_A_2120_55#_c_1451_n N_VPWR_c_1499_n 0.0428704f $X=10.745 $Y=1.98 $X2=0
+ $Y2=0
cc_904 N_A_2120_55#_c_1447_n N_VPWR_c_1499_n 0.0214059f $X=11.41 $Y=1.48 $X2=0
+ $Y2=0
cc_905 N_A_2120_55#_c_1448_n N_VPWR_c_1499_n 0.00300514f $X=11.41 $Y=1.48 $X2=0
+ $Y2=0
cc_906 N_A_2120_55#_M1012_g N_VPWR_c_1502_n 0.0054895f $X=11.505 $Y=2.465 $X2=0
+ $Y2=0
cc_907 N_A_2120_55#_M1012_g N_VPWR_c_1494_n 0.0072954f $X=11.505 $Y=2.465 $X2=0
+ $Y2=0
cc_908 N_A_2120_55#_M1012_g N_KAPWR_c_1663_n 0.00753768f $X=11.505 $Y=2.465
+ $X2=0 $Y2=0
cc_909 N_A_2120_55#_c_1451_n N_KAPWR_c_1663_n 0.0179077f $X=10.745 $Y=1.98 $X2=0
+ $Y2=0
cc_910 N_A_2120_55#_M1012_g N_Q_c_1777_n 0.0137945f $X=11.505 $Y=2.465 $X2=0
+ $Y2=0
cc_911 N_A_2120_55#_M1012_g N_Q_c_1778_n 0.00270591f $X=11.505 $Y=2.465 $X2=0
+ $Y2=0
cc_912 N_A_2120_55#_c_1447_n N_Q_c_1778_n 0.00151667f $X=11.41 $Y=1.48 $X2=0
+ $Y2=0
cc_913 N_A_2120_55#_M1016_g N_Q_c_1774_n 0.0160633f $X=11.505 $Y=0.695 $X2=0
+ $Y2=0
cc_914 N_A_2120_55#_c_1447_n N_Q_c_1774_n 0.0262122f $X=11.41 $Y=1.48 $X2=0
+ $Y2=0
cc_915 N_A_2120_55#_M1016_g Q 0.00430192f $X=11.505 $Y=0.695 $X2=0 $Y2=0
cc_916 N_A_2120_55#_c_1446_n Q 0.00422903f $X=10.745 $Y=0.485 $X2=0 $Y2=0
cc_917 N_A_2120_55#_c_1447_n Q 0.00144832f $X=11.41 $Y=1.48 $X2=0 $Y2=0
cc_918 N_A_2120_55#_M1016_g N_Q_c_1776_n 0.0112457f $X=11.505 $Y=0.695 $X2=0
+ $Y2=0
cc_919 N_A_2120_55#_M1016_g N_VGND_c_1801_n 0.00268481f $X=11.505 $Y=0.695 $X2=0
+ $Y2=0
cc_920 N_A_2120_55#_c_1446_n N_VGND_c_1801_n 0.0454719f $X=10.745 $Y=0.485 $X2=0
+ $Y2=0
cc_921 N_A_2120_55#_c_1447_n N_VGND_c_1801_n 0.0122725f $X=11.41 $Y=1.48 $X2=0
+ $Y2=0
cc_922 N_A_2120_55#_c_1448_n N_VGND_c_1801_n 0.00269229f $X=11.41 $Y=1.48 $X2=0
+ $Y2=0
cc_923 N_A_2120_55#_c_1446_n N_VGND_c_1809_n 0.0234289f $X=10.745 $Y=0.485 $X2=0
+ $Y2=0
cc_924 N_A_2120_55#_M1016_g N_VGND_c_1810_n 0.00511358f $X=11.505 $Y=0.695 $X2=0
+ $Y2=0
cc_925 N_A_2120_55#_M1016_g N_VGND_c_1811_n 0.0104744f $X=11.505 $Y=0.695 $X2=0
+ $Y2=0
cc_926 N_A_2120_55#_c_1446_n N_VGND_c_1811_n 0.0126421f $X=10.745 $Y=0.485 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1498_n N_A_280_97#_c_1616_n 0.0282666f $X=1.325 $Y=2.59 $X2=0
+ $Y2=0
cc_928 N_VPWR_c_1500_n N_A_280_97#_c_1617_n 0.0189735f $X=4.3 $Y=3.33 $X2=0
+ $Y2=0
cc_929 N_VPWR_c_1494_n N_A_280_97#_c_1617_n 0.00302557f $X=11.76 $Y=3.33 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1494_n N_KAPWR_M1028_d 0.00118319f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_931 N_VPWR_c_1494_n N_KAPWR_M1004_d 0.00119816f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_932 N_VPWR_c_1501_n N_KAPWR_c_1660_n 0.0301317f $X=11.125 $Y=3.33 $X2=0 $Y2=0
cc_933 N_VPWR_c_1494_n N_KAPWR_c_1660_n 0.00607782f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_934 N_VPWR_c_1505_n N_KAPWR_c_1660_n 8.16568e-19 $X=4.465 $Y=3.06 $X2=0 $Y2=0
cc_935 N_VPWR_c_1501_n N_KAPWR_c_1661_n 0.0220975f $X=11.125 $Y=3.33 $X2=0 $Y2=0
cc_936 N_VPWR_c_1494_n N_KAPWR_c_1661_n 0.00445397f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_937 N_VPWR_c_1501_n N_KAPWR_c_1666_n 0.0184875f $X=11.125 $Y=3.33 $X2=0 $Y2=0
cc_938 N_VPWR_c_1494_n N_KAPWR_c_1666_n 0.00288279f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_939 N_VPWR_c_1501_n N_KAPWR_c_1662_n 0.0262182f $X=11.125 $Y=3.33 $X2=0 $Y2=0
cc_940 N_VPWR_c_1494_n N_KAPWR_c_1662_n 0.00367312f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_941 N_VPWR_M1032_s N_KAPWR_c_1663_n 0.0115361f $X=0.135 $Y=2.435 $X2=0 $Y2=0
cc_942 N_VPWR_M1031_d N_KAPWR_c_1663_n 0.00323939f $X=1.07 $Y=2.435 $X2=0 $Y2=0
cc_943 N_VPWR_M1033_d N_KAPWR_c_1663_n 0.0015771f $X=4.21 $Y=1.935 $X2=0 $Y2=0
cc_944 N_VPWR_M1034_d N_KAPWR_c_1663_n 0.00244555f $X=11.035 $Y=1.835 $X2=0
+ $Y2=0
cc_945 N_VPWR_c_1495_n N_KAPWR_c_1663_n 2.42196e-19 $X=0.28 $Y=3.245 $X2=0 $Y2=0
cc_946 N_VPWR_c_1496_n N_KAPWR_c_1663_n 0.0234704f $X=0.28 $Y=2.93 $X2=0 $Y2=0
cc_947 N_VPWR_c_1497_n N_KAPWR_c_1663_n 0.00218028f $X=1.16 $Y=3.33 $X2=0 $Y2=0
cc_948 N_VPWR_c_1498_n N_KAPWR_c_1663_n 0.0310158f $X=1.325 $Y=2.59 $X2=0 $Y2=0
cc_949 N_VPWR_c_1499_n N_KAPWR_c_1663_n 0.0369087f $X=11.29 $Y=1.98 $X2=0 $Y2=0
cc_950 N_VPWR_c_1500_n N_KAPWR_c_1663_n 0.00862591f $X=4.3 $Y=3.33 $X2=0 $Y2=0
cc_951 N_VPWR_c_1501_n N_KAPWR_c_1663_n 0.0164436f $X=11.125 $Y=3.33 $X2=0 $Y2=0
cc_952 N_VPWR_c_1502_n N_KAPWR_c_1663_n 0.00124399f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_953 N_VPWR_c_1494_n N_KAPWR_c_1663_n 1.25077f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_954 N_VPWR_c_1505_n N_KAPWR_c_1663_n 0.00267734f $X=4.465 $Y=3.06 $X2=0 $Y2=0
cc_955 N_VPWR_c_1494_n A_1565_419# 8.56818e-19 $X=11.76 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_956 N_VPWR_c_1494_n A_1765_419# 0.00128775f $X=11.76 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_957 N_VPWR_c_1494_n N_Q_M1012_d 0.00119401f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_958 N_VPWR_c_1502_n N_Q_c_1777_n 0.0231698f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_959 N_VPWR_c_1494_n N_Q_c_1777_n 0.00332052f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_960 N_VPWR_c_1499_n N_Q_c_1778_n 0.0494754f $X=11.29 $Y=1.98 $X2=0 $Y2=0
cc_961 N_A_280_97#_c_1617_n N_KAPWR_c_1663_n 0.0376925f $X=1.825 $Y=2.745 $X2=0
+ $Y2=0
cc_962 N_A_280_97#_c_1614_n N_VGND_c_1799_n 0.0149959f $X=1.745 $Y=0.655 $X2=0
+ $Y2=0
cc_963 N_A_280_97#_c_1614_n N_VGND_c_1805_n 0.0128163f $X=1.745 $Y=0.655 $X2=0
+ $Y2=0
cc_964 N_A_280_97#_c_1614_n N_VGND_c_1811_n 0.0150619f $X=1.745 $Y=0.655 $X2=0
+ $Y2=0
cc_965 A_423_487# N_KAPWR_c_1663_n 0.00952953f $X=2.115 $Y=2.435 $X2=10.32
+ $Y2=2.82
cc_966 N_KAPWR_c_1663_n A_1565_419# 0.0042906f $X=10.32 $Y=2.82 $X2=-0.19
+ $Y2=1.655
cc_967 N_KAPWR_c_1663_n A_1765_419# 0.00282253f $X=10.32 $Y=2.82 $X2=-0.19
+ $Y2=1.655
cc_968 N_KAPWR_c_1663_n N_Q_c_1777_n 0.041515f $X=10.32 $Y=2.82 $X2=0 $Y2=0
cc_969 N_Q_c_1776_n N_VGND_c_1801_n 0.0264802f $X=11.72 $Y=0.42 $X2=0 $Y2=0
cc_970 N_Q_c_1776_n N_VGND_c_1810_n 0.0255795f $X=11.72 $Y=0.42 $X2=0 $Y2=0
cc_971 N_Q_c_1776_n N_VGND_c_1811_n 0.0138084f $X=11.72 $Y=0.42 $X2=0 $Y2=0
cc_972 N_VGND_c_1811_n N_A_1624_47#_M1007_s 0.00444922f $X=11.76 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_973 N_VGND_c_1811_n N_A_1624_47#_M1022_d 0.00233209f $X=11.76 $Y=0 $X2=0
+ $Y2=0
cc_974 N_VGND_c_1808_n N_A_1624_47#_c_1932_n 0.0150075f $X=8.61 $Y=0 $X2=0 $Y2=0
cc_975 N_VGND_c_1811_n N_A_1624_47#_c_1932_n 0.0094309f $X=11.76 $Y=0 $X2=0
+ $Y2=0
cc_976 N_VGND_M1007_d N_A_1624_47#_c_1929_n 0.00378274f $X=8.555 $Y=0.235 $X2=0
+ $Y2=0
cc_977 N_VGND_c_1808_n N_A_1624_47#_c_1929_n 0.00330923f $X=8.61 $Y=0 $X2=0
+ $Y2=0
cc_978 N_VGND_c_1809_n N_A_1624_47#_c_1929_n 0.00342183f $X=11.125 $Y=0 $X2=0
+ $Y2=0
cc_979 N_VGND_c_1811_n N_A_1624_47#_c_1929_n 0.0117739f $X=11.76 $Y=0 $X2=0
+ $Y2=0
cc_980 N_VGND_c_1812_n N_A_1624_47#_c_1929_n 0.0239935f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_981 N_VGND_c_1809_n N_A_1624_47#_c_1931_n 0.0185707f $X=11.125 $Y=0 $X2=0
+ $Y2=0
cc_982 N_VGND_c_1811_n N_A_1624_47#_c_1931_n 0.0124445f $X=11.76 $Y=0 $X2=0
+ $Y2=0
cc_983 N_VGND_c_1811_n A_1917_47# 0.00899413f $X=11.76 $Y=0 $X2=-0.19 $Y2=-0.245
