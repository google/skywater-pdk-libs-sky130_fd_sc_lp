* File: sky130_fd_sc_lp__a221o_lp.spice
* Created: Fri Aug 28 09:52:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a221o_lp.pex.spice"
.subckt sky130_fd_sc_lp__a221o_lp  VNB VPB A2 A1 B1 B2 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1010 A_162_66# N_A_96_183#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_96_183#_M1013_g A_162_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0441 PD=0.78 PS=0.63 NRD=22.848 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1004 A_336_66# N_A2_M1004_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.1 SB=75002.7
+ A=0.063 P=1.14 MULT=1
MM1011 N_A_96_183#_M1011_d N_A1_M1011_g A_336_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.1449 AS=0.0504 PD=1.11 PS=0.66 NRD=117.132 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1000 A_582_66# N_B1_M1000_g N_A_96_183#_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1449 PD=0.66 PS=1.11 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_B2_M1001_g A_582_66# VNB NSHORT L=0.15 W=0.42 AD=0.0777
+ AS=0.0504 PD=0.79 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.7 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1007 A_764_66# N_C1_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0777 PD=0.63 PS=0.79 NRD=14.28 NRS=25.704 M=1 R=2.8 SA=75003.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_96_183#_M1008_d N_C1_M1008_g A_764_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_96_183#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.275 AS=0.285 PD=1.55 PS=2.57 NRD=45.2903 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1005 N_A_322_419#_M1005_d N_A2_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.275 PD=1.28 PS=1.55 NRD=0 NRS=7.8603 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g N_A_322_419#_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1009 N_A_322_419#_M1009_d N_B1_M1009_g N_A_545_400#_M1009_s VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1006 N_A_545_400#_M1006_d N_B2_M1006_g N_A_322_419#_M1009_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1002 N_A_96_183#_M1002_d N_C1_M1002_g N_A_545_400#_M1006_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__a221o_lp.pxi.spice"
*
.ends
*
*
