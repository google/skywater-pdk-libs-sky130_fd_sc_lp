* File: sky130_fd_sc_lp__o22a_2.pex.spice
* Created: Fri Aug 28 11:09:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22A_2%A_80_23# 1 2 9 13 17 21 26 28 29 30 31 34 36
+ 38 45
r89 44 45 16.3786 $w=3.09e-07 $l=1.05e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=1.01 $Y2=1.41
r90 43 44 50.6958 $w=3.09e-07 $l=3.25e-07 $layer=POLY_cond $X=0.58 $Y=1.41
+ $X2=0.905 $Y2=1.41
r91 36 41 2.61083 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.417 $Y=2.1
+ $X2=2.417 $Y2=2.015
r92 36 38 27.0574 $w=3.43e-07 $l=8.1e-07 $layer=LI1_cond $X=2.417 $Y=2.1
+ $X2=2.417 $Y2=2.91
r93 32 34 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.09 $Y=1.075
+ $X2=2.09 $Y2=0.76
r94 30 41 5.28309 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.245 $Y=2.015
+ $X2=2.417 $Y2=2.015
r95 30 31 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.245 $Y=2.015 $X2=1.31
+ $Y2=2.015
r96 28 32 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.975 $Y=1.16
+ $X2=2.09 $Y2=1.075
r97 28 29 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.975 $Y=1.16
+ $X2=1.31 $Y2=1.16
r98 27 45 21.0583 $w=3.09e-07 $l=1.35e-07 $layer=POLY_cond $X=1.145 $Y=1.41
+ $X2=1.01 $Y2=1.41
r99 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.145
+ $Y=1.41 $X2=1.145 $Y2=1.41
r100 24 31 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.18 $Y=1.93
+ $X2=1.31 $Y2=2.015
r101 24 26 23.0489 $w=2.58e-07 $l=5.2e-07 $layer=LI1_cond $X=1.18 $Y=1.93
+ $X2=1.18 $Y2=1.41
r102 23 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.18 $Y=1.245
+ $X2=1.31 $Y2=1.16
r103 23 26 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.18 $Y=1.245
+ $X2=1.18 $Y2=1.41
r104 19 45 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.575
+ $X2=1.01 $Y2=1.41
r105 19 21 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.01 $Y=1.575
+ $X2=1.01 $Y2=2.465
r106 15 44 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.245
+ $X2=0.905 $Y2=1.41
r107 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.905 $Y=1.245
+ $X2=0.905 $Y2=0.665
r108 11 43 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.575
+ $X2=0.58 $Y2=1.41
r109 11 13 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.58 $Y=1.575
+ $X2=0.58 $Y2=2.465
r110 7 43 16.3786 $w=3.09e-07 $l=2.11069e-07 $layer=POLY_cond $X=0.475 $Y=1.245
+ $X2=0.58 $Y2=1.41
r111 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.475 $Y=1.245
+ $X2=0.475 $Y2=0.665
r112 2 41 400 $w=1.7e-07 $l=3.42053e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.48 $Y2=2.095
r113 2 38 400 $w=1.7e-07 $l=1.16614e-06 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.48 $Y2=2.91
r114 1 34 182 $w=1.7e-07 $l=5.89597e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.245 $X2=2.09 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_2%B1 3 7 9 12 13
c38 3 0 8.31843e-20 $X=1.855 $Y=0.665
r39 12 15 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.747 $Y=1.51
+ $X2=1.747 $Y2=1.675
r40 12 14 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.747 $Y=1.51
+ $X2=1.747 $Y2=1.345
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.51 $X2=1.73 $Y2=1.51
r42 9 13 4.30431 $w=4.13e-07 $l=1.55e-07 $layer=LI1_cond $X=1.687 $Y=1.665
+ $X2=1.687 $Y2=1.51
r43 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.855 $Y=2.465
+ $X2=1.855 $Y2=1.675
r44 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.855 $Y=0.665
+ $X2=1.855 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_2%B2 3 7 9 12 13
c40 7 0 6.40318e-20 $X=2.305 $Y=0.665
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.51
+ $X2=2.305 $Y2=1.675
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.305
+ $Y=1.51 $X2=2.305 $Y2=1.51
r43 9 13 4.52224 $w=3.93e-07 $l=1.55e-07 $layer=LI1_cond $X=2.272 $Y=1.665
+ $X2=2.272 $Y2=1.51
r44 5 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.345
+ $X2=2.305 $Y2=1.51
r45 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.305 $Y=1.345
+ $X2=2.305 $Y2=0.665
r46 3 14 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.215 $Y=2.465
+ $X2=2.215 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_2%A2 3 7 9 10 11 12 18 19
c38 18 0 1.7958e-19 $X=2.845 $Y=1.51
r39 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.51
+ $X2=2.845 $Y2=1.675
r40 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.51
+ $X2=2.845 $Y2=1.345
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.51 $X2=2.845 $Y2=1.51
r42 11 12 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.982 $Y=2.405
+ $X2=2.982 $Y2=2.775
r43 10 11 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.982 $Y=2.035
+ $X2=2.982 $Y2=2.405
r44 9 10 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.982 $Y=1.665
+ $X2=2.982 $Y2=2.035
r45 9 19 4.01413 $w=4.43e-07 $l=1.55e-07 $layer=LI1_cond $X=2.982 $Y=1.665
+ $X2=2.982 $Y2=1.51
r46 7 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.78 $Y=0.665
+ $X2=2.78 $Y2=1.345
r47 3 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.755 $Y=2.465
+ $X2=2.755 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_2%A1 3 7 9 14 15
c23 15 0 1.7958e-19 $X=3.55 $Y=1.46
r24 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.46 $X2=3.55 $Y2=1.46
r25 11 14 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.31 $Y=1.46
+ $X2=3.55 $Y2=1.46
r26 9 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.46
r27 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.625
+ $X2=3.31 $Y2=1.46
r28 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.31 $Y=1.625 $X2=3.31
+ $Y2=2.465
r29 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.295
+ $X2=3.31 $Y2=1.46
r30 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.31 $Y=1.295 $X2=3.31
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_2%VPWR 1 2 3 10 12 18 20 22 26 28 33 45 49
r49 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 40 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r53 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r56 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 34 45 14.1136 $w=1.7e-07 $l=3.73e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.432 $Y2=3.33
r58 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 33 48 4.52193 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.607 $Y2=3.33
r60 33 39 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 32 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 32 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 29 42 3.92003 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.225 $Y2=3.33
r65 29 31 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=3.33 $X2=0.72
+ $Y2=3.33
r66 28 45 14.1136 $w=1.7e-07 $l=3.72e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=1.432 $Y2=3.33
r67 28 31 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 26 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 26 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 22 25 31.6465 $w=3.13e-07 $l=8.65e-07 $layer=LI1_cond $X=3.532 $Y=2.085
+ $X2=3.532 $Y2=2.95
r71 20 48 3.11857 $w=3.15e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.532 $Y=3.245
+ $X2=3.607 $Y2=3.33
r72 20 25 10.7927 $w=3.13e-07 $l=2.95e-07 $layer=LI1_cond $X=3.532 $Y=3.245
+ $X2=3.532 $Y2=2.95
r73 16 45 2.99104 $w=7.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.432 $Y=3.245
+ $X2=1.432 $Y2=3.33
r74 16 18 13.9676 $w=7.43e-07 $l=8.7e-07 $layer=LI1_cond $X=1.432 $Y=3.245
+ $X2=1.432 $Y2=2.375
r75 12 15 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.325 $Y=2.16
+ $X2=0.325 $Y2=2.95
r76 10 42 3.22313 $w=2.5e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.325 $Y=3.245
+ $X2=0.225 $Y2=3.33
r77 10 15 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.325 $Y=3.245
+ $X2=0.325 $Y2=2.95
r78 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.835 $X2=3.525 $Y2=2.95
r79 3 22 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.835 $X2=3.525 $Y2=2.085
r80 2 18 150 $w=1.7e-07 $l=7.79567e-07 $layer=licon1_PDIFF $count=4 $X=1.085
+ $Y=1.835 $X2=1.64 $Y2=2.375
r81 1 15 400 $w=1.7e-07 $l=1.18763e-06 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.365 $Y2=2.95
r82 1 12 400 $w=1.7e-07 $l=3.92906e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.365 $Y2=2.16
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_2%X 1 2 9 11 12 13 14 15 26 43
c20 13 0 5.82976e-20 $X=0.72 $Y=2.035
r21 24 43 0.40085 $w=3.43e-07 $l=1.2e-08 $layer=LI1_cond $X=0.707 $Y=1.653
+ $X2=0.707 $Y2=1.665
r22 23 26 1.6034 $w=3.43e-07 $l=4.8e-08 $layer=LI1_cond $X=0.707 $Y=1.247
+ $X2=0.707 $Y2=1.295
r23 15 38 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.75 $Y=2.775
+ $X2=0.75 $Y2=2.91
r24 14 15 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.75 $Y=2.405
+ $X2=0.75 $Y2=2.775
r25 13 14 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=0.75 $Y=1.98
+ $X2=0.75 $Y2=2.405
r26 13 45 6.87033 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.75 $Y=1.98
+ $X2=0.75 $Y2=1.825
r27 12 45 4.86827 $w=3.43e-07 $l=1.24e-07 $layer=LI1_cond $X=0.707 $Y=1.701
+ $X2=0.707 $Y2=1.825
r28 12 43 1.20255 $w=3.43e-07 $l=3.6e-08 $layer=LI1_cond $X=0.707 $Y=1.701
+ $X2=0.707 $Y2=1.665
r29 12 24 1.23595 $w=3.43e-07 $l=3.7e-08 $layer=LI1_cond $X=0.707 $Y=1.616
+ $X2=0.707 $Y2=1.653
r30 11 23 0.634679 $w=3.43e-07 $l=1.9e-08 $layer=LI1_cond $X=0.707 $Y=1.228
+ $X2=0.707 $Y2=1.247
r31 11 41 6.19006 $w=3.43e-07 $l=1.53e-07 $layer=LI1_cond $X=0.707 $Y=1.228
+ $X2=0.707 $Y2=1.075
r32 11 12 10.1215 $w=3.43e-07 $l=3.03e-07 $layer=LI1_cond $X=0.707 $Y=1.313
+ $X2=0.707 $Y2=1.616
r33 11 26 0.601275 $w=3.43e-07 $l=1.8e-08 $layer=LI1_cond $X=0.707 $Y=1.313
+ $X2=0.707 $Y2=1.295
r34 9 41 31.4521 $w=2.38e-07 $l=6.55e-07 $layer=LI1_cond $X=0.655 $Y=0.42
+ $X2=0.655 $Y2=1.075
r35 2 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=1.835 $X2=0.795 $Y2=2.91
r36 2 13 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=1.835 $X2=0.795 $Y2=1.98
r37 1 9 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.245 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
r50 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r54 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.04
+ $Y2=0
r56 37 39 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.6
+ $Y2=0
r57 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r58 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r59 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r60 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r61 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r62 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r63 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.68
+ $Y2=0
r64 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=3.04
+ $Y2=0
r65 29 35 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.64
+ $Y2=0
r66 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r67 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r68 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 25 43 4.21867 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r70 25 27 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r71 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r72 24 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.72
+ $Y2=0
r73 22 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r74 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r75 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0
r76 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.04 $Y=0.085
+ $X2=3.04 $Y2=0.37
r77 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r78 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.39
r79 10 43 3.06603 $w=2.7e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.182 $Y2=0
r80 10 12 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.23 $Y2=0.39
r81 3 20 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=2.855
+ $Y=0.245 $X2=3.04 $Y2=0.37
r82 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.245 $X2=1.12 $Y2=0.39
r83 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.245 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_2%A_303_49# 1 2 3 12 14 15 16 17 20 23
c44 17 0 8.31843e-20 $X=2.705 $Y=1.08
c45 14 0 6.40318e-20 $X=2.54 $Y=0.425
r46 18 20 21.0367 $w=3.13e-07 $l=5.75e-07 $layer=LI1_cond $X=3.532 $Y=0.995
+ $X2=3.532 $Y2=0.42
r47 16 18 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=3.375 $Y=1.08
+ $X2=3.532 $Y2=0.995
r48 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.375 $Y=1.08
+ $X2=2.705 $Y2=1.08
r49 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.54 $Y=0.995
+ $X2=2.705 $Y2=1.08
r50 14 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.425 $X2=2.54
+ $Y2=0.34
r51 14 15 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=2.54 $Y=0.425
+ $X2=2.54 $Y2=0.995
r52 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0.34
+ $X2=1.64 $Y2=0.34
r53 12 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0.34
+ $X2=2.54 $Y2=0.34
r54 12 13 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.375 $Y=0.34
+ $X2=1.805 $Y2=0.34
r55 3 20 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.245 $X2=3.525 $Y2=0.42
r56 2 25 91 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_NDIFF $count=2 $X=2.38
+ $Y=0.245 $X2=2.54 $Y2=0.42
r57 1 23 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.245 $X2=1.64 $Y2=0.39
.ends

