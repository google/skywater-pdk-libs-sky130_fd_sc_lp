* File: sky130_fd_sc_lp__o211a_2.spice
* Created: Fri Aug 28 11:02:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o211a_2.pex.spice"
.subckt sky130_fd_sc_lp__o211a_2  VNB VPB C1 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1006 A_110_47# N_C1_M1006_g N_A_27_47#_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1000 N_A_182_47#_M1000_d N_B1_M1000_g A_110_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_182_47#_M1004_d N_A2_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A1_M1011_g N_A_182_47#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1011_d N_A_27_47#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A_27_47#_M1008_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.3276 AS=0.1176 PD=2.46 PS=1.12 NRD=8.928 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1010 N_VPWR_M1010_d N_C1_M1010_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.3339 PD=1.58 PS=3.05 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1007 N_A_27_47#_M1007_d N_B1_M1007_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3276 AS=0.2016 PD=1.78 PS=1.58 NRD=12.4898 NRS=3.1126 M=1 R=8.4
+ SA=75000.7 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1003 A_372_367# N_A2_M1003_g N_A_27_47#_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3276 PD=1.47 PS=1.78 NRD=7.8012 NRS=24.9993 M=1 R=8.4
+ SA=75001.3 SB=75001.8 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g A_372_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.1323 PD=1.88 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.7
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3906 PD=1.54 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_X_M1001_d N_A_27_47#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o211a_2.pxi.spice"
*
.ends
*
*
