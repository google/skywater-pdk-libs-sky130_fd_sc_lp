* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
X0 VPWR a_1046_367# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_453_480# a_27_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND GATE a_279_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR CLK a_1046_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_437_81# a_27_367# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_321_55# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_27_367# a_80_269# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_27_367# a_80_269# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_1046_367# a_27_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VGND CLK a_1002_79# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_279_81# a_321_55# a_80_269# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND a_321_55# a_315_382# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_80_269# a_321_55# a_453_480# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_321_55# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_321_55# a_315_382# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_1002_79# a_27_367# a_1046_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR GATE a_273_480# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_273_480# a_315_382# a_80_269# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_80_269# a_315_382# a_437_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_1046_367# GCLK VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
