* File: sky130_fd_sc_lp__and4_0.pex.spice
* Created: Wed Sep  2 09:32:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4_0%A 3 7 9 10 12 13 14 15 16 22
c38 13 0 9.5044e-20 $X=0.24 $Y=0.925
r39 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.35
+ $Y=1.005 $X2=0.35 $Y2=1.005
r40 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.035
r41 14 15 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r42 14 23 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.005
r43 13 23 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=0.925 $X2=0.26
+ $Y2=1.005
r44 11 22 33.2483 $w=4.6e-07 $l=2.75e-07 $layer=POLY_cond $X=0.415 $Y=1.28
+ $X2=0.415 $Y2=1.005
r45 11 12 55.0748 $w=4.6e-07 $l=2.3e-07 $layer=POLY_cond $X=0.415 $Y=1.28
+ $X2=0.415 $Y2=1.51
r46 10 22 4.23161 $w=4.6e-07 $l=3.5e-08 $layer=POLY_cond $X=0.415 $Y=0.97
+ $X2=0.415 $Y2=1.005
r47 9 10 45.4026 $w=4.6e-07 $l=1.5e-07 $layer=POLY_cond $X=0.51 $Y=0.82 $X2=0.51
+ $Y2=0.97
r48 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.76 $Y=0.5 $X2=0.76
+ $Y2=0.82
r49 3 12 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=0.57 $Y=2.6 $X2=0.57
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_0%B 3 7 11 12 13 14 18
c43 7 0 9.5044e-20 $X=1.12 $Y=0.5
r44 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.03
+ $Y=1.375 $X2=1.03 $Y2=1.375
r45 14 19 8.56945 $w=3.88e-07 $l=2.9e-07 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.375
r46 13 19 2.36399 $w=3.88e-07 $l=8e-08 $layer=LI1_cond $X=1.14 $Y=1.295 $X2=1.14
+ $Y2=1.375
r47 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.03 $Y=1.715
+ $X2=1.03 $Y2=1.375
r48 11 12 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.715
+ $X2=1.03 $Y2=1.88
r49 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.21
+ $X2=1.03 $Y2=1.375
r50 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.12 $Y=0.5 $X2=1.12
+ $Y2=1.21
r51 3 12 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1 $Y=2.6 $X2=1
+ $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_0%C 3 6 9 11 12 13 17
c40 3 0 3.59751e-20 $X=1.48 $Y=0.5
r41 17 19 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.335
+ $X2=1.58 $Y2=1.17
r42 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.59
+ $Y=1.335 $X2=1.59 $Y2=1.335
r43 13 18 11.8846 $w=3.18e-07 $l=3.3e-07 $layer=LI1_cond $X=1.665 $Y=1.665
+ $X2=1.665 $Y2=1.335
r44 12 18 1.44055 $w=3.18e-07 $l=4e-08 $layer=LI1_cond $X=1.665 $Y=1.295
+ $X2=1.665 $Y2=1.335
r45 9 11 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.48 $Y=2.6 $X2=1.48
+ $Y2=1.84
r46 6 11 48.0802 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.58 $Y=1.665
+ $X2=1.58 $Y2=1.84
r47 5 17 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=1.58 $Y=1.345 $X2=1.58
+ $Y2=1.335
r48 5 6 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.58 $Y=1.345 $X2=1.58
+ $Y2=1.665
r49 3 19 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.48 $Y=0.5 $X2=1.48
+ $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_0%D 1 3 6 12 15 16 18 19 20 21 26
c49 19 0 3.59751e-20 $X=2.16 $Y=1.295
c50 15 0 1.73574e-19 $X=2.08 $Y=2.08
r51 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=2.035
r52 20 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.16
+ $Y=1.725 $X2=2.16 $Y2=1.725
r53 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.665
r54 18 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.56
+ $X2=2.16 $Y2=1.725
r55 15 26 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.16 $Y=2.08
+ $X2=2.16 $Y2=1.725
r56 15 16 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.08 $Y=2.08
+ $X2=2.08 $Y2=2.23
r57 10 12 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.84 $Y=0.885
+ $X2=2.07 $Y2=0.885
r58 8 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.07 $Y=0.96 $X2=2.07
+ $Y2=0.885
r59 8 18 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.07 $Y=0.96 $X2=2.07
+ $Y2=1.56
r60 6 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.91 $Y=2.6 $X2=1.91
+ $Y2=2.23
r61 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=0.81 $X2=1.84
+ $Y2=0.885
r62 1 3 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.84 $Y=0.81 $X2=1.84
+ $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_0%A_84_58# 1 2 3 12 15 18 19 21 23 25 28 30 32
+ 36 43 45 46 48 49
c95 32 0 1.73574e-19 $X=1.555 $Y=2.162
r96 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.73
+ $Y=0.985 $X2=2.73 $Y2=0.985
r97 41 43 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.545 $Y=0.495
+ $X2=0.695 $Y2=0.495
r98 34 36 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.69 $Y=2.265
+ $X2=1.69 $Y2=2.575
r99 33 46 1.51462 $w=2.05e-07 $l=1.55e-07 $layer=LI1_cond $X=0.915 $Y=2.162
+ $X2=0.76 $Y2=2.162
r100 32 34 6.98383 $w=2.05e-07 $l=1.79248e-07 $layer=LI1_cond $X=1.555 $Y=2.162
+ $X2=1.69 $Y2=2.265
r101 32 33 34.6253 $w=2.03e-07 $l=6.4e-07 $layer=LI1_cond $X=1.555 $Y=2.162
+ $X2=0.915 $Y2=2.162
r102 31 45 1.44715 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.785 $Y=0.905
+ $X2=0.695 $Y2=0.905
r103 30 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.565 $Y=0.905
+ $X2=2.69 $Y2=0.905
r104 30 31 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=2.565 $Y=0.905
+ $X2=0.785 $Y2=0.905
r105 26 46 4.96437 $w=2.15e-07 $l=1.14822e-07 $layer=LI1_cond $X=0.785 $Y=2.265
+ $X2=0.76 $Y2=2.162
r106 26 28 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=0.785 $Y=2.265
+ $X2=0.785 $Y2=2.6
r107 25 46 4.96437 $w=2.15e-07 $l=1.32454e-07 $layer=LI1_cond $X=0.69 $Y=2.06
+ $X2=0.76 $Y2=2.162
r108 24 45 5.04255 $w=1.75e-07 $l=8.74643e-08 $layer=LI1_cond $X=0.69 $Y=0.99
+ $X2=0.695 $Y2=0.905
r109 24 25 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=0.69 $Y=0.99
+ $X2=0.69 $Y2=2.06
r110 23 45 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.82
+ $X2=0.695 $Y2=0.905
r111 22 43 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=0.66
+ $X2=0.695 $Y2=0.495
r112 22 23 9.85859 $w=1.78e-07 $l=1.6e-07 $layer=LI1_cond $X=0.695 $Y=0.66
+ $X2=0.695 $Y2=0.82
r113 20 49 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=0.985
r114 20 21 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=1.49
r115 19 49 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.73 $Y=0.97
+ $X2=2.73 $Y2=0.985
r116 18 19 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.715 $Y=0.82
+ $X2=2.715 $Y2=0.97
r117 15 21 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.745 $Y=2.71
+ $X2=2.745 $Y2=1.49
r118 12 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.61 $Y=0.5
+ $X2=2.61 $Y2=0.82
r119 3 36 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=1.555
+ $Y=2.39 $X2=1.695 $Y2=2.575
r120 2 28 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=2.39 $X2=0.785 $Y2=2.6
r121 1 41 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.42
+ $Y=0.29 $X2=0.545 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_0%VPWR 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r38 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 37 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 34 46 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.332 $Y2=3.33
r44 34 36 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 30 43 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.235 $Y2=3.33
r46 30 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 29 46 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.332 $Y2=3.33
r48 29 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 25 40 4.2956 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.242 $Y2=3.33
r53 25 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 24 43 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=1.235 $Y2=3.33
r55 24 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 22 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 22 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 22 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 18 46 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.332 $Y=3.245
+ $X2=2.332 $Y2=3.33
r60 18 20 12.4038 $w=6.73e-07 $l=7e-07 $layer=LI1_cond $X=2.332 $Y=3.245
+ $X2=2.332 $Y2=2.545
r61 14 43 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=3.33
r62 14 16 24.7775 $w=2.98e-07 $l=6.45e-07 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=2.6
r63 10 40 3.18193 $w=2.95e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.337 $Y=3.245
+ $X2=0.242 $Y2=3.33
r64 10 12 25.1975 $w=2.93e-07 $l=6.45e-07 $layer=LI1_cond $X=0.337 $Y=3.245
+ $X2=0.337 $Y2=2.6
r65 3 20 200 $w=1.7e-07 $l=6.17657e-07 $layer=licon1_PDIFF $count=3 $X=1.985
+ $Y=2.39 $X2=2.53 $Y2=2.545
r66 2 16 600 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=2.39 $X2=1.23 $Y2=2.6
r67 1 12 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.23
+ $Y=2.39 $X2=0.355 $Y2=2.6
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_0%X 1 2 7 8 9 10 11 12 13 42 45
r18 45 46 2.21075 $w=4.33e-07 $l=3.5e-08 $layer=LI1_cond $X=3.057 $Y=2.405
+ $X2=3.057 $Y2=2.37
r19 33 49 1.37763 $w=4.33e-07 $l=5.2e-08 $layer=LI1_cond $X=3.057 $Y=2.587
+ $X2=3.057 $Y2=2.535
r20 22 42 1.49285 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=0.65
+ $X2=3.13 $Y2=0.485
r21 13 33 4.98067 $w=4.33e-07 $l=1.88e-07 $layer=LI1_cond $X=3.057 $Y=2.775
+ $X2=3.057 $Y2=2.587
r22 12 49 2.78176 $w=4.33e-07 $l=1.05e-07 $layer=LI1_cond $X=3.057 $Y=2.43
+ $X2=3.057 $Y2=2.535
r23 12 45 0.662324 $w=4.33e-07 $l=2.5e-08 $layer=LI1_cond $X=3.057 $Y=2.43
+ $X2=3.057 $Y2=2.405
r24 12 46 0.993485 $w=2.88e-07 $l=2.5e-08 $layer=LI1_cond $X=3.13 $Y=2.345
+ $X2=3.13 $Y2=2.37
r25 11 12 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=3.13 $Y=2.035
+ $X2=3.13 $Y2=2.345
r26 10 11 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=1.665
+ $X2=3.13 $Y2=2.035
r27 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=1.295
+ $X2=3.13 $Y2=1.665
r28 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=0.925 $X2=3.13
+ $Y2=1.295
r29 8 22 10.9283 $w=2.88e-07 $l=2.75e-07 $layer=LI1_cond $X=3.13 $Y=0.925
+ $X2=3.13 $Y2=0.65
r30 7 42 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=3.12 $Y=0.485 $X2=3.13
+ $Y2=0.485
r31 7 38 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.12 $Y=0.485
+ $X2=2.825 $Y2=0.485
r32 2 49 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.82
+ $Y=2.39 $X2=2.96 $Y2=2.535
r33 1 38 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.685
+ $Y=0.29 $X2=2.825 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_0%VGND 1 4 6 16 17
r24 17 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r25 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r26 14 16 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.525 $Y=0 $X2=3.12
+ $Y2=0
r27 8 12 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r28 8 9 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 6 24 9.1354 $w=6.33e-07 $l=4.85e-07 $layer=LI1_cond $X=2.207 $Y=0 $X2=2.207
+ $Y2=0.485
r30 6 14 8.68381 $w=1.7e-07 $l=3.18e-07 $layer=LI1_cond $X=2.207 $Y=0 $X2=2.525
+ $Y2=0
r31 6 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r32 6 12 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.68
+ $Y2=0
r33 4 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r34 4 9 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r35 4 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r36 1 24 91 $w=1.7e-07 $l=5.6921e-07 $layer=licon1_NDIFF $count=2 $X=1.915
+ $Y=0.29 $X2=2.395 $Y2=0.485
.ends

