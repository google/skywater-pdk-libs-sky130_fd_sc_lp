* File: sky130_fd_sc_lp__a21boi_1.pex.spice
* Created: Fri Aug 28 09:49:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BOI_1%B1_N 2 5 7 8 11 15 18 20 21 22 23 29
r40 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r41 22 23 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=2.035
r42 21 22 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.665
r43 21 30 7.46954 $w=2.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.12
r44 20 30 8.3232 $w=2.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.22 $Y=0.925
+ $X2=0.22 $Y2=1.12
r45 16 18 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=0.36 $Y=1.99
+ $X2=0.475 $Y2=1.99
r46 14 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.27 $Y2=1.12
r47 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.27 $Y2=1.625
r48 13 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.105
+ $X2=0.27 $Y2=1.12
r49 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.805 $Y=0.955
+ $X2=0.805 $Y2=0.445
r50 8 13 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=1.03
+ $X2=0.27 $Y2=1.105
r51 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.73 $Y=1.03
+ $X2=0.805 $Y2=0.955
r52 7 8 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.73 $Y=1.03
+ $X2=0.435 $Y2=1.03
r53 3 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.065
+ $X2=0.475 $Y2=1.99
r54 3 5 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.475 $Y=2.065
+ $X2=0.475 $Y2=2.75
r55 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=1.915
+ $X2=0.36 $Y2=1.99
r56 2 15 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.36 $Y=1.915
+ $X2=0.36 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_1%A_27_508# 1 2 7 11 15 18 22 24 25 28 31 36
+ 38 39
c72 39 0 1.74246e-19 $X=0.84 $Y=1.42
c73 18 0 1.41666e-19 $X=1.435 $Y=1.42
c74 11 0 1.04703e-19 $X=1.33 $Y=0.655
r75 34 36 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=0.59 $Y=0.445
+ $X2=0.745 $Y2=0.445
r76 32 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.84 $Y=1.51 $X2=0.84
+ $Y2=1.42
r77 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.84
+ $Y=1.51 $X2=0.84 $Y2=1.51
r78 29 31 34.3558 $w=2.63e-07 $l=7.9e-07 $layer=LI1_cond $X=0.792 $Y=2.3
+ $X2=0.792 $Y2=1.51
r79 28 38 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=0.792 $Y=1.477
+ $X2=0.792 $Y2=1.345
r80 28 31 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=0.792 $Y=1.477
+ $X2=0.792 $Y2=1.51
r81 26 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.745 $Y=0.61
+ $X2=0.745 $Y2=0.445
r82 26 38 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.745 $Y=0.61
+ $X2=0.745 $Y2=1.345
r83 24 29 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=0.66 $Y=2.385
+ $X2=0.792 $Y2=2.3
r84 24 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.66 $Y=2.385
+ $X2=0.355 $Y2=2.385
r85 20 25 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=2.47
+ $X2=0.355 $Y2=2.385
r86 20 22 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=0.225 $Y=2.47
+ $X2=0.225 $Y2=2.75
r87 17 18 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=1.33 $Y=1.42
+ $X2=1.435 $Y2=1.42
r88 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.435 $Y=1.495
+ $X2=1.435 $Y2=1.42
r89 13 15 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=1.435 $Y=1.495
+ $X2=1.435 $Y2=2.465
r90 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.33 $Y=1.345
+ $X2=1.33 $Y2=1.42
r91 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.33 $Y=1.345
+ $X2=1.33 $Y2=0.655
r92 8 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.42
+ $X2=0.84 $Y2=1.42
r93 7 17 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.255 $Y=1.42
+ $X2=1.33 $Y2=1.42
r94 7 8 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.255 $Y=1.42
+ $X2=1.005 $Y2=1.42
r95 2 22 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.26 $Y2=2.75
r96 1 34 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.465
+ $Y=0.235 $X2=0.59 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_1%A1 3 6 8 9 10 15 17
c36 10 0 2.46369e-19 $X=2.16 $Y=1.295
r37 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.35
+ $X2=1.915 $Y2=1.515
r38 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.35
+ $X2=1.915 $Y2=1.185
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.35 $X2=1.915 $Y2=1.35
r40 10 16 1.4914 $w=4.23e-07 $l=5.5e-08 $layer=LI1_cond $X=2.042 $Y=1.295
+ $X2=2.042 $Y2=1.35
r41 10 29 7.59257 $w=4.23e-07 $l=2.8e-07 $layer=LI1_cond $X=2.042 $Y=1.295
+ $X2=2.042 $Y2=1.015
r42 9 29 2.33078 $w=4.43e-07 $l=9e-08 $layer=LI1_cond $X=2.052 $Y=0.925
+ $X2=2.052 $Y2=1.015
r43 8 9 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.052 $Y=0.555
+ $X2=2.052 $Y2=0.925
r44 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.865 $Y=2.465
+ $X2=1.865 $Y2=1.515
r45 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.825 $Y=0.655
+ $X2=1.825 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_1%A2 3 6 8 11 13
r23 11 14 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=2.497 $Y=1.35
+ $X2=2.497 $Y2=1.515
r24 11 13 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=2.497 $Y=1.35
+ $X2=2.497 $Y2=1.185
r25 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.35 $X2=2.51 $Y2=1.35
r26 8 12 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=1.35 $X2=2.51
+ $Y2=1.35
r27 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.395 $Y=2.465
+ $X2=2.395 $Y2=1.515
r28 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.395 $Y=0.655
+ $X2=2.395 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_1%VPWR 1 2 9 13 17 19 24 31 32 35 38
r37 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.135 $Y2=3.33
r42 29 31 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.3 $Y=3.33 $X2=2.64
+ $Y2=3.33
r43 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 25 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r46 25 27 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=2.135 $Y2=3.33
r48 24 27 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 19 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r52 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 17 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 17 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 13 16 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.135 $Y=2.11
+ $X2=2.135 $Y2=2.95
r56 11 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=3.33
r57 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=2.95
r58 7 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r59 7 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.765
r60 2 16 400 $w=1.7e-07 $l=1.20857e-06 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.135 $Y2=2.95
r61 2 13 400 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.135 $Y2=2.11
r62 1 9 600 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.54 $X2=0.69 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_1%Y 1 2 7 9 11 12 13 14 15
c33 7 0 1.74246e-19 $X=1.537 $Y=1.21
r34 21 37 1.67288 $w=2.6e-07 $l=1.53e-07 $layer=LI1_cond $X=1.225 $Y=1.515
+ $X2=1.225 $Y2=1.362
r35 15 32 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=1.225 $Y=2.775
+ $X2=1.225 $Y2=2.91
r36 14 15 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.225 $Y=2.405
+ $X2=1.225 $Y2=2.775
r37 13 14 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=1.225 $Y=1.98
+ $X2=1.225 $Y2=2.405
r38 12 13 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.225 $Y=1.665
+ $X2=1.225 $Y2=1.98
r39 12 21 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.225 $Y=1.665
+ $X2=1.225 $Y2=1.515
r40 11 37 0.944625 $w=3.03e-07 $l=2.5e-08 $layer=LI1_cond $X=1.2 $Y=1.362
+ $X2=1.225 $Y2=1.362
r41 7 37 11.7889 $w=3.03e-07 $l=3.12e-07 $layer=LI1_cond $X=1.537 $Y=1.362
+ $X2=1.225 $Y2=1.362
r42 7 9 37.1604 $w=2.43e-07 $l=7.9e-07 $layer=LI1_cond $X=1.537 $Y=1.21
+ $X2=1.537 $Y2=0.42
r43 2 32 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.835 $X2=1.22 $Y2=2.91
r44 2 13 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.835 $X2=1.22 $Y2=1.98
r45 1 9 91 $w=1.7e-07 $l=2.56271e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.235 $X2=1.575 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_1%A_302_367# 1 2 9 13 14 17
r25 17 19 35.1401 $w=3.03e-07 $l=9.3e-07 $layer=LI1_cond $X=2.622 $Y=1.98
+ $X2=2.622 $Y2=2.91
r26 15 17 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=2.622 $Y=1.855
+ $X2=2.622 $Y2=1.98
r27 13 15 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=2.47 $Y=1.77
+ $X2=2.622 $Y2=1.855
r28 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.47 $Y=1.77 $X2=1.8
+ $Y2=1.77
r29 9 11 38.9735 $w=2.73e-07 $l=9.3e-07 $layer=LI1_cond $X=1.662 $Y=1.98
+ $X2=1.662 $Y2=2.91
r30 7 14 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=1.662 $Y=1.855
+ $X2=1.8 $Y2=1.77
r31 7 9 5.23838 $w=2.73e-07 $l=1.25e-07 $layer=LI1_cond $X=1.662 $Y=1.855
+ $X2=1.662 $Y2=1.98
r32 2 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.835 $X2=2.61 $Y2=2.91
r33 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.835 $X2=2.61 $Y2=1.98
r34 1 11 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.835 $X2=1.65 $Y2=2.91
r35 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.835 $X2=1.65 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_1%VGND 1 2 9 11 13 15 17 22 28 32
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r37 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r39 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r40 23 28 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.122
+ $Y2=0
r41 23 25 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=2.16
+ $Y2=0
r42 22 31 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.662
+ $Y2=0
r43 22 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.16
+ $Y2=0
r44 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r45 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 17 28 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=1 $Y=0 $X2=1.122
+ $Y2=0
r47 17 19 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.72
+ $Y2=0
r48 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r49 15 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r50 11 31 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.662 $Y2=0
r51 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.38
r52 7 28 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.122 $Y=0.085
+ $X2=1.122 $Y2=0
r53 7 9 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=1.122 $Y=0.085
+ $X2=1.122 $Y2=0.38
r54 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.47
+ $Y=0.235 $X2=2.61 $Y2=0.38
r55 1 9 91 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=2 $X=0.88
+ $Y=0.235 $X2=1.115 $Y2=0.38
.ends

