* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrbp_1 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_626_119# a_218_483# a_773_525# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1000_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_373_481# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 Q_N a_1187_131# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR a_49_93# a_218_483# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VGND a_776_93# a_1187_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_49_93# a_218_483# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_776_93# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR a_626_119# a_776_93# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR a_776_93# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND a_373_481# a_554_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_626_119# a_49_93# a_734_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_776_93# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_373_481# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_773_525# a_776_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_49_93# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 a_554_119# a_218_483# a_626_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_734_119# a_776_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_776_93# a_626_119# a_1000_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VPWR a_373_481# a_596_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_596_481# a_49_93# a_626_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VPWR a_776_93# a_1187_131# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 Q_N a_1187_131# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_49_93# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
