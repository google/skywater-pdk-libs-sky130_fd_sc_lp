* File: sky130_fd_sc_lp__iso1p_lp2.pxi.spice
* Created: Wed Sep  2 09:58:15 2020
* 
x_PM_SKY130_FD_SC_LP__ISO1P_LP2%A N_A_M1006_g N_A_c_54_n N_A_M1003_g N_A_M1000_g
+ N_A_c_55_n A A N_A_c_52_n N_A_c_53_n PM_SKY130_FD_SC_LP__ISO1P_LP2%A
x_PM_SKY130_FD_SC_LP__ISO1P_LP2%SLEEP N_SLEEP_M1007_g N_SLEEP_c_90_n
+ N_SLEEP_M1004_g N_SLEEP_c_91_n N_SLEEP_M1008_g N_SLEEP_c_96_n SLEEP SLEEP
+ PM_SKY130_FD_SC_LP__ISO1P_LP2%SLEEP
x_PM_SKY130_FD_SC_LP__ISO1P_LP2%A_137_409# N_A_137_409#_M1000_d
+ N_A_137_409#_M1003_s N_A_137_409#_M1001_g N_A_137_409#_M1005_g
+ N_A_137_409#_M1002_g N_A_137_409#_c_142_n N_A_137_409#_c_143_n
+ N_A_137_409#_c_151_n N_A_137_409#_c_144_n N_A_137_409#_c_145_n
+ N_A_137_409#_c_146_n N_A_137_409#_c_147_n N_A_137_409#_c_148_n
+ N_A_137_409#_c_153_n N_A_137_409#_c_149_n
+ PM_SKY130_FD_SC_LP__ISO1P_LP2%A_137_409#
x_PM_SKY130_FD_SC_LP__ISO1P_LP2%KAPWR N_KAPWR_M1004_d KAPWR N_KAPWR_c_228_n
+ N_KAPWR_c_226_n N_KAPWR_c_227_n PM_SKY130_FD_SC_LP__ISO1P_LP2%KAPWR
x_PM_SKY130_FD_SC_LP__ISO1P_LP2%X N_X_M1002_d N_X_M1005_d N_X_c_258_n X X X X X
+ X N_X_c_257_n PM_SKY130_FD_SC_LP__ISO1P_LP2%X
x_PM_SKY130_FD_SC_LP__ISO1P_LP2%VGND N_VGND_M1006_s N_VGND_M1008_d
+ N_VGND_c_278_n N_VGND_c_279_n N_VGND_c_280_n N_VGND_c_281_n VGND
+ N_VGND_c_282_n N_VGND_c_283_n N_VGND_c_284_n N_VGND_c_285_n
+ PM_SKY130_FD_SC_LP__ISO1P_LP2%VGND
x_PM_SKY130_FD_SC_LP__ISO1P_LP2%VPWR VPWR N_VPWR_c_316_n VPWR
+ PM_SKY130_FD_SC_LP__ISO1P_LP2%VPWR
cc_1 VNB N_A_M1006_g 0.0355136f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.495
cc_2 VNB N_A_M1000_g 0.0241568f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=0.495
cc_3 VNB N_A_c_52_n 0.0677891f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.17
cc_4 VNB N_A_c_53_n 0.0429613f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.17
cc_5 VNB N_SLEEP_M1007_g 0.0305305f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.495
cc_6 VNB N_SLEEP_c_90_n 0.0215092f $X=-0.19 $Y=-0.245 $X2=1.037 $Y2=1.915
cc_7 VNB N_SLEEP_c_91_n 0.0262562f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=0.495
cc_8 VNB N_SLEEP_M1008_g 0.0309151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB SLEEP 0.00352148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_137_409#_M1001_g 0.0180448f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=2.545
cc_11 VNB N_A_137_409#_M1005_g 0.00927166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_137_409#_M1002_g 0.0229269f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_A_137_409#_c_142_n 0.0274427f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.17
cc_14 VNB N_A_137_409#_c_143_n 0.016656f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.675
cc_15 VNB N_A_137_409#_c_144_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_137_409#_c_145_n 0.00464655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_137_409#_c_146_n 0.0213231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_137_409#_c_147_n 0.00124064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_137_409#_c_148_n 0.0278529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_137_409#_c_149_n 0.00549821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_257_n 0.0813828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_278_n 0.0255778f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=2.545
cc_23 VNB N_VGND_c_279_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_280_n 0.0110534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_281_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_26 VNB N_VGND_c_282_n 0.0362073f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.17
cc_27 VNB N_VGND_c_283_n 0.0328777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_284_n 0.219229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_285_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB VPWR 0.143779f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.005
cc_31 VPB N_A_c_54_n 0.0308788f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=2.04
cc_32 VPB N_A_c_55_n 0.0163225f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=1.915
cc_33 VPB N_A_c_52_n 0.0124157f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.17
cc_34 VPB N_A_c_53_n 0.0310389f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.17
cc_35 VPB N_SLEEP_c_90_n 6.8022e-19 $X=-0.19 $Y=1.655 $X2=1.037 $Y2=1.915
cc_36 VPB N_SLEEP_M1004_g 0.0324556f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=2.545
cc_37 VPB N_SLEEP_c_96_n 0.0147539f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_38 VPB SLEEP 0.00371997f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_137_409#_M1005_g 0.0510103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_137_409#_c_151_n 0.0304728f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_137_409#_c_145_n 0.003116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_137_409#_c_153_n 0.00993551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_KAPWR_c_226_n 0.020402f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=0.495
cc_44 VPB N_KAPWR_c_227_n 0.0545402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_X_c_258_n 0.0173753f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=2.545
cc_46 VPB X 0.0466135f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=0.495
cc_47 VPB N_X_c_257_n 0.0184503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB VPWR 0.0571699f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.005
cc_49 VPB N_VPWR_c_316_n 0.0968731f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=2.545
cc_50 N_A_M1000_g N_SLEEP_M1007_g 0.0182874f $X=1.05 $Y=0.495 $X2=0 $Y2=0
cc_51 N_A_c_52_n N_SLEEP_c_90_n 0.0114152f $X=0.75 $Y=1.17 $X2=0 $Y2=0
cc_52 N_A_c_54_n N_SLEEP_M1004_g 0.0808369f $X=1.075 $Y=2.04 $X2=0 $Y2=0
cc_53 N_A_c_52_n N_SLEEP_c_91_n 0.0182874f $X=0.75 $Y=1.17 $X2=0 $Y2=0
cc_54 N_A_c_55_n N_SLEEP_c_96_n 0.0114152f $X=1.075 $Y=1.915 $X2=0 $Y2=0
cc_55 N_A_c_52_n SLEEP 6.16949e-19 $X=0.75 $Y=1.17 $X2=0 $Y2=0
cc_56 N_A_c_54_n N_A_137_409#_c_151_n 0.01732f $X=1.075 $Y=2.04 $X2=0 $Y2=0
cc_57 N_A_M1006_g N_A_137_409#_c_144_n 0.00177001f $X=0.66 $Y=0.495 $X2=0 $Y2=0
cc_58 N_A_M1000_g N_A_137_409#_c_144_n 0.0114071f $X=1.05 $Y=0.495 $X2=0 $Y2=0
cc_59 N_A_c_54_n N_A_137_409#_c_145_n 0.00782483f $X=1.075 $Y=2.04 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_A_137_409#_c_145_n 3.10823e-19 $X=1.05 $Y=0.495 $X2=0 $Y2=0
cc_61 N_A_c_55_n N_A_137_409#_c_145_n 0.00845693f $X=1.075 $Y=1.915 $X2=0 $Y2=0
cc_62 N_A_c_52_n N_A_137_409#_c_145_n 0.0159626f $X=0.75 $Y=1.17 $X2=0 $Y2=0
cc_63 N_A_c_53_n N_A_137_409#_c_145_n 0.0554449f $X=0.75 $Y=1.17 $X2=0 $Y2=0
cc_64 N_A_c_54_n N_A_137_409#_c_153_n 0.0166607f $X=1.075 $Y=2.04 $X2=0 $Y2=0
cc_65 N_A_c_52_n N_A_137_409#_c_153_n 0.00259263f $X=0.75 $Y=1.17 $X2=0 $Y2=0
cc_66 N_A_c_53_n N_A_137_409#_c_153_n 0.0176002f $X=0.75 $Y=1.17 $X2=0 $Y2=0
cc_67 N_A_M1006_g N_A_137_409#_c_149_n 8.3456e-19 $X=0.66 $Y=0.495 $X2=0 $Y2=0
cc_68 N_A_M1000_g N_A_137_409#_c_149_n 0.00525549f $X=1.05 $Y=0.495 $X2=0 $Y2=0
cc_69 N_A_c_54_n N_KAPWR_c_228_n 0.00143422f $X=1.075 $Y=2.04 $X2=0 $Y2=0
cc_70 N_A_c_54_n N_KAPWR_c_226_n 0.00182597f $X=1.075 $Y=2.04 $X2=0 $Y2=0
cc_71 N_A_c_54_n N_KAPWR_c_227_n 0.00702466f $X=1.075 $Y=2.04 $X2=0 $Y2=0
cc_72 N_A_M1006_g N_VGND_c_278_n 0.014477f $X=0.66 $Y=0.495 $X2=0 $Y2=0
cc_73 N_A_M1000_g N_VGND_c_278_n 0.00213234f $X=1.05 $Y=0.495 $X2=0 $Y2=0
cc_74 N_A_c_53_n N_VGND_c_278_n 0.0213781f $X=0.75 $Y=1.17 $X2=0 $Y2=0
cc_75 N_A_M1006_g N_VGND_c_282_n 0.00445056f $X=0.66 $Y=0.495 $X2=0 $Y2=0
cc_76 N_A_M1000_g N_VGND_c_282_n 0.00502664f $X=1.05 $Y=0.495 $X2=0 $Y2=0
cc_77 N_A_M1006_g N_VGND_c_284_n 0.00802306f $X=0.66 $Y=0.495 $X2=0 $Y2=0
cc_78 N_A_M1000_g N_VGND_c_284_n 0.00948105f $X=1.05 $Y=0.495 $X2=0 $Y2=0
cc_79 N_A_c_54_n VPWR 0.00834414f $X=1.075 $Y=2.04 $X2=-0.19 $Y2=-0.245
cc_80 N_A_c_54_n N_VPWR_c_316_n 0.0086001f $X=1.075 $Y=2.04 $X2=0 $Y2=0
cc_81 N_SLEEP_M1008_g N_A_137_409#_M1001_g 0.0193087f $X=1.84 $Y=0.495 $X2=0
+ $Y2=0
cc_82 N_SLEEP_c_90_n N_A_137_409#_M1005_g 0.00510685f $X=1.575 $Y=1.665 $X2=0
+ $Y2=0
cc_83 N_SLEEP_M1004_g N_A_137_409#_M1005_g 0.00784066f $X=1.535 $Y=2.545 $X2=0
+ $Y2=0
cc_84 SLEEP N_A_137_409#_M1005_g 0.00539226f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_85 N_SLEEP_c_91_n N_A_137_409#_c_142_n 0.0193087f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_86 N_SLEEP_M1004_g N_A_137_409#_c_151_n 0.00204468f $X=1.535 $Y=2.545 $X2=0
+ $Y2=0
cc_87 N_SLEEP_M1007_g N_A_137_409#_c_144_n 0.0111815f $X=1.48 $Y=0.495 $X2=0
+ $Y2=0
cc_88 N_SLEEP_M1008_g N_A_137_409#_c_144_n 0.00192036f $X=1.84 $Y=0.495 $X2=0
+ $Y2=0
cc_89 N_SLEEP_M1007_g N_A_137_409#_c_145_n 0.00516537f $X=1.48 $Y=0.495 $X2=0
+ $Y2=0
cc_90 N_SLEEP_c_90_n N_A_137_409#_c_145_n 0.00739372f $X=1.575 $Y=1.665 $X2=0
+ $Y2=0
cc_91 SLEEP N_A_137_409#_c_145_n 0.0453483f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_92 N_SLEEP_M1007_g N_A_137_409#_c_146_n 0.00909887f $X=1.48 $Y=0.495 $X2=0
+ $Y2=0
cc_93 N_SLEEP_c_91_n N_A_137_409#_c_146_n 2.08789e-19 $X=1.84 $Y=1.16 $X2=0
+ $Y2=0
cc_94 N_SLEEP_M1008_g N_A_137_409#_c_146_n 0.0144162f $X=1.84 $Y=0.495 $X2=0
+ $Y2=0
cc_95 SLEEP N_A_137_409#_c_146_n 0.0257428f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_96 N_SLEEP_M1008_g N_A_137_409#_c_147_n 0.00197081f $X=1.84 $Y=0.495 $X2=0
+ $Y2=0
cc_97 SLEEP N_A_137_409#_c_147_n 0.0148177f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_98 N_SLEEP_c_90_n N_A_137_409#_c_148_n 0.00386246f $X=1.575 $Y=1.665 $X2=0
+ $Y2=0
cc_99 SLEEP N_A_137_409#_c_148_n 0.00195827f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_100 N_SLEEP_M1004_g N_A_137_409#_c_153_n 0.00156068f $X=1.535 $Y=2.545 $X2=0
+ $Y2=0
cc_101 N_SLEEP_M1007_g N_A_137_409#_c_149_n 0.00366045f $X=1.48 $Y=0.495 $X2=0
+ $Y2=0
cc_102 N_SLEEP_M1004_g N_KAPWR_c_228_n 0.0137081f $X=1.535 $Y=2.545 $X2=0 $Y2=0
cc_103 N_SLEEP_M1004_g N_KAPWR_c_226_n 0.0183009f $X=1.535 $Y=2.545 $X2=0 $Y2=0
cc_104 N_SLEEP_c_91_n N_KAPWR_c_226_n 0.00370206f $X=1.84 $Y=1.16 $X2=0 $Y2=0
cc_105 N_SLEEP_c_96_n N_KAPWR_c_226_n 6.15373e-19 $X=1.575 $Y=1.83 $X2=0 $Y2=0
cc_106 SLEEP N_KAPWR_c_226_n 0.0128211f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_107 N_SLEEP_M1004_g N_KAPWR_c_227_n 0.0113013f $X=1.535 $Y=2.545 $X2=0 $Y2=0
cc_108 N_SLEEP_M1007_g N_VGND_c_279_n 0.00188065f $X=1.48 $Y=0.495 $X2=0 $Y2=0
cc_109 N_SLEEP_M1008_g N_VGND_c_279_n 0.0105659f $X=1.84 $Y=0.495 $X2=0 $Y2=0
cc_110 N_SLEEP_M1007_g N_VGND_c_282_n 0.00502664f $X=1.48 $Y=0.495 $X2=0 $Y2=0
cc_111 N_SLEEP_M1008_g N_VGND_c_282_n 0.00445056f $X=1.84 $Y=0.495 $X2=0 $Y2=0
cc_112 N_SLEEP_M1007_g N_VGND_c_284_n 0.00562693f $X=1.48 $Y=0.495 $X2=0 $Y2=0
cc_113 N_SLEEP_M1008_g N_VGND_c_284_n 0.00418511f $X=1.84 $Y=0.495 $X2=0 $Y2=0
cc_114 N_SLEEP_M1004_g VPWR 0.00699111f $X=1.535 $Y=2.545 $X2=-0.19 $Y2=-0.245
cc_115 N_SLEEP_M1004_g N_VPWR_c_316_n 0.00591772f $X=1.535 $Y=2.545 $X2=0 $Y2=0
cc_116 N_A_137_409#_c_153_n A_240_409# 0.00199525f $X=1.185 $Y=2.11 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_137_409#_c_151_n N_KAPWR_c_228_n 0.00635454f $X=0.81 $Y=2.9 $X2=0
+ $Y2=0
cc_118 N_A_137_409#_M1005_g N_KAPWR_c_226_n 0.0212932f $X=2.405 $Y=2.545 $X2=0
+ $Y2=0
cc_119 N_A_137_409#_c_143_n N_KAPWR_c_226_n 5.61113e-19 $X=2.362 $Y=1.535 $X2=0
+ $Y2=0
cc_120 N_A_137_409#_c_151_n N_KAPWR_c_226_n 0.0164244f $X=0.81 $Y=2.9 $X2=0
+ $Y2=0
cc_121 N_A_137_409#_c_147_n N_KAPWR_c_226_n 0.0053106f $X=2.36 $Y=1.03 $X2=0
+ $Y2=0
cc_122 N_A_137_409#_c_153_n N_KAPWR_c_226_n 0.00810268f $X=1.185 $Y=2.11 $X2=0
+ $Y2=0
cc_123 N_A_137_409#_M1005_g N_KAPWR_c_227_n 0.00860102f $X=2.405 $Y=2.545 $X2=0
+ $Y2=0
cc_124 N_A_137_409#_c_151_n N_KAPWR_c_227_n 0.0295961f $X=0.81 $Y=2.9 $X2=0
+ $Y2=0
cc_125 N_A_137_409#_c_153_n N_KAPWR_c_227_n 0.0097815f $X=1.185 $Y=2.11 $X2=0
+ $Y2=0
cc_126 N_A_137_409#_M1005_g N_X_c_258_n 0.007909f $X=2.405 $Y=2.545 $X2=0 $Y2=0
cc_127 N_A_137_409#_M1005_g X 0.0170239f $X=2.405 $Y=2.545 $X2=0 $Y2=0
cc_128 N_A_137_409#_c_147_n X 7.88315e-19 $X=2.36 $Y=1.03 $X2=0 $Y2=0
cc_129 N_A_137_409#_M1001_g N_X_c_257_n 0.00197815f $X=2.27 $Y=0.495 $X2=0 $Y2=0
cc_130 N_A_137_409#_M1002_g N_X_c_257_n 0.0149277f $X=2.66 $Y=0.495 $X2=0 $Y2=0
cc_131 N_A_137_409#_c_142_n N_X_c_257_n 0.0065668f $X=2.66 $Y=0.94 $X2=0 $Y2=0
cc_132 N_A_137_409#_c_146_n N_X_c_257_n 0.0132836f $X=2.195 $Y=0.905 $X2=0 $Y2=0
cc_133 N_A_137_409#_c_147_n N_X_c_257_n 0.0418161f $X=2.36 $Y=1.03 $X2=0 $Y2=0
cc_134 N_A_137_409#_c_148_n N_X_c_257_n 0.0277138f $X=2.36 $Y=1.03 $X2=0 $Y2=0
cc_135 N_A_137_409#_c_144_n N_VGND_c_278_n 0.0145731f $X=1.265 $Y=0.495 $X2=0
+ $Y2=0
cc_136 N_A_137_409#_M1001_g N_VGND_c_279_n 0.0108205f $X=2.27 $Y=0.495 $X2=0
+ $Y2=0
cc_137 N_A_137_409#_M1002_g N_VGND_c_279_n 0.00189174f $X=2.66 $Y=0.495 $X2=0
+ $Y2=0
cc_138 N_A_137_409#_c_144_n N_VGND_c_279_n 0.0125465f $X=1.265 $Y=0.495 $X2=0
+ $Y2=0
cc_139 N_A_137_409#_c_146_n N_VGND_c_279_n 0.020143f $X=2.195 $Y=0.905 $X2=0
+ $Y2=0
cc_140 N_A_137_409#_c_144_n N_VGND_c_282_n 0.021949f $X=1.265 $Y=0.495 $X2=0
+ $Y2=0
cc_141 N_A_137_409#_M1001_g N_VGND_c_283_n 0.00445056f $X=2.27 $Y=0.495 $X2=0
+ $Y2=0
cc_142 N_A_137_409#_M1002_g N_VGND_c_283_n 0.00502664f $X=2.66 $Y=0.495 $X2=0
+ $Y2=0
cc_143 N_A_137_409#_M1001_g N_VGND_c_284_n 0.00424333f $X=2.27 $Y=0.495 $X2=0
+ $Y2=0
cc_144 N_A_137_409#_M1002_g N_VGND_c_284_n 0.0102162f $X=2.66 $Y=0.495 $X2=0
+ $Y2=0
cc_145 N_A_137_409#_c_144_n N_VGND_c_284_n 0.0124703f $X=1.265 $Y=0.495 $X2=0
+ $Y2=0
cc_146 N_A_137_409#_c_146_n N_VGND_c_284_n 0.0268598f $X=2.195 $Y=0.905 $X2=0
+ $Y2=0
cc_147 N_A_137_409#_M1005_g VPWR 0.00866127f $X=2.405 $Y=2.545 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A_137_409#_c_151_n VPWR 0.00355217f $X=0.81 $Y=2.9 $X2=-0.19 $Y2=-0.245
cc_149 N_A_137_409#_M1005_g N_VPWR_c_316_n 0.00784959f $X=2.405 $Y=2.545 $X2=0
+ $Y2=0
cc_150 N_A_137_409#_c_151_n N_VPWR_c_316_n 0.0220321f $X=0.81 $Y=2.9 $X2=0 $Y2=0
cc_151 A_240_409# N_KAPWR_c_228_n 0.00232299f $X=1.2 $Y=2.045 $X2=0 $Y2=0
cc_152 A_240_409# N_KAPWR_c_227_n 0.00500544f $X=1.2 $Y=2.045 $X2=2.66 $Y2=0.495
cc_153 N_KAPWR_c_227_n N_X_c_258_n 0.0399757f $X=2.2 $Y=2.775 $X2=0 $Y2=0
cc_154 N_KAPWR_c_226_n X 0.0816843f $X=1.8 $Y=2.19 $X2=0 $Y2=0
cc_155 N_KAPWR_c_227_n X 0.0226011f $X=2.2 $Y=2.775 $X2=0 $Y2=0
cc_156 N_KAPWR_c_228_n VPWR 0.00172069f $X=1.635 $Y=2.775 $X2=-0.19 $Y2=1.655
cc_157 N_KAPWR_c_226_n VPWR 0.00752488f $X=1.8 $Y=2.19 $X2=-0.19 $Y2=1.655
cc_158 N_KAPWR_c_227_n VPWR 0.293573f $X=2.2 $Y=2.775 $X2=-0.19 $Y2=1.655
cc_159 N_KAPWR_c_228_n N_VPWR_c_316_n 0.00854674f $X=1.635 $Y=2.775 $X2=0 $Y2=0
cc_160 N_KAPWR_c_226_n N_VPWR_c_316_n 0.0467922f $X=1.8 $Y=2.19 $X2=0 $Y2=0
cc_161 N_KAPWR_c_227_n N_VPWR_c_316_n 0.0100763f $X=2.2 $Y=2.775 $X2=0 $Y2=0
cc_162 N_X_c_257_n N_VGND_c_279_n 0.0123173f $X=2.875 $Y=0.495 $X2=0 $Y2=0
cc_163 N_X_c_257_n N_VGND_c_283_n 0.0351799f $X=2.875 $Y=0.495 $X2=0 $Y2=0
cc_164 N_X_c_257_n N_VGND_c_284_n 0.020126f $X=2.875 $Y=0.495 $X2=0 $Y2=0
cc_165 N_X_c_258_n VPWR 0.00355217f $X=2.67 $Y=2.9 $X2=-0.19 $Y2=-0.245
cc_166 N_X_c_258_n N_VPWR_c_316_n 0.0220321f $X=2.67 $Y=2.9 $X2=0 $Y2=0
