* NGSPICE file created from sky130_fd_sc_lp__a21bo_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 VPWR a_188_315# X VPB phighvt w=1.26e+06u l=150000u
+  ad=1.7955e+12p pd=1.545e+07u as=7.056e+11p ps=6.16e+06u
M1001 X a_188_315# VGND VNB nshort w=840000u l=150000u
+  ad=4.788e+11p pd=4.5e+06u as=1.9152e+12p ps=1.296e+07u
M1002 a_908_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1003 X a_188_315# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_188_315# a_42_47# a_645_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.3734e+12p ps=1.226e+07u
M1005 a_188_315# a_42_47# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1006 a_645_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_908_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A2 a_645_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_188_315# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_645_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_188_315# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_188_315# A1 a_908_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND B1_N a_42_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1014 a_908_47# A1 a_188_315# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A1 a_645_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_188_315# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_645_367# a_42_47# a_188_315# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_188_315# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_188_315# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_42_47# a_188_315# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR B1_N a_42_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

