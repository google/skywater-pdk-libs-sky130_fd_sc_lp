# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__clkbuflp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__clkbuflp_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.384000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.140000 0.715000 1.565000 ;
        RECT 0.125000 1.565000 0.425000 1.880000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.428000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745000 1.705000 6.735000 1.790000 ;
        RECT 2.745000 1.790000 5.195000 1.875000 ;
        RECT 2.745000 1.875000 4.135000 1.885000 ;
        RECT 2.745000 1.885000 3.075000 3.075000 ;
        RECT 3.005000 0.345000 3.335000 0.775000 ;
        RECT 3.005000 0.775000 4.960000 1.035000 ;
        RECT 3.805000 1.885000 4.135000 3.075000 ;
        RECT 4.100000 1.035000 4.960000 1.170000 ;
        RECT 4.100000 1.170000 6.735000 1.705000 ;
        RECT 4.585000 0.345000 4.960000 0.775000 ;
        RECT 4.865000 1.875000 5.195000 3.075000 ;
        RECT 5.875000 0.265000 6.735000 1.170000 ;
        RECT 5.925000 1.790000 6.255000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.095000  2.065000 0.425000 3.245000 ;
      RECT 0.125000  0.085000 0.425000 0.890000 ;
      RECT 0.625000  1.770000 1.995000 1.940000 ;
      RECT 0.625000  1.940000 0.955000 3.075000 ;
      RECT 0.885000  0.255000 1.230000 0.985000 ;
      RECT 0.955000  0.985000 1.230000 1.205000 ;
      RECT 0.955000  1.205000 3.870000 1.535000 ;
      RECT 0.955000  1.535000 1.995000 1.770000 ;
      RECT 1.155000  2.110000 1.485000 3.245000 ;
      RECT 1.660000  1.940000 1.995000 3.075000 ;
      RECT 1.675000  0.085000 2.550000 0.875000 ;
      RECT 2.215000  2.085000 2.545000 3.245000 ;
      RECT 3.275000  2.085000 3.605000 3.245000 ;
      RECT 3.795000  0.085000 4.125000 0.605000 ;
      RECT 4.335000  2.085000 4.665000 3.245000 ;
      RECT 5.375000  0.085000 5.705000 0.675000 ;
      RECT 5.395000  2.085000 5.725000 3.245000 ;
      RECT 6.455000  2.085000 6.785000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_lp__clkbuflp_8
END LIBRARY
