* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__ha_0 A B VGND VNB VPB VPWR COUT SUM
X0 a_80_60# a_204_315# a_307_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_307_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR a_204_315# a_80_60# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR a_204_315# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_204_315# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR B a_204_315# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND a_204_315# COUT VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND A a_307_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_687_135# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_393_491# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_204_315# B a_687_135# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 SUM a_80_60# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_80_60# B a_393_491# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 SUM a_80_60# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
