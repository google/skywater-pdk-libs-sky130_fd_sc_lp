* File: sky130_fd_sc_lp__o2111ai_2.pex.spice
* Created: Fri Aug 28 11:01:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111AI_2%D1 1 3 6 8 10 13 15 16 24
r42 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.555 $Y=1.46
+ $X2=0.985 $Y2=1.46
r43 20 23 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.34 $Y=1.46
+ $X2=0.555 $Y2=1.46
r44 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.46 $X2=0.34 $Y2=1.46
r45 16 21 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=1.46
r46 15 21 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.46
r47 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.625
+ $X2=0.985 $Y2=1.46
r48 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.985 $Y=1.625
+ $X2=0.985 $Y2=2.465
r49 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.295
+ $X2=0.985 $Y2=1.46
r50 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.985 $Y=1.295
+ $X2=0.985 $Y2=0.765
r51 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.625
+ $X2=0.555 $Y2=1.46
r52 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.555 $Y=1.625
+ $X2=0.555 $Y2=2.465
r53 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.295
+ $X2=0.555 $Y2=1.46
r54 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.555 $Y=1.295
+ $X2=0.555 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%C1 1 3 6 8 10 13 15 16 25 27 33
c60 25 0 1.86523e-19 $X=1.845 $Y=1.46
c61 1 0 6.1024e-20 $X=1.415 $Y=1.295
r62 27 33 3.58273 $w=3.35e-07 $l=7.2e-08 $layer=LI1_cond $X=1.608 $Y=1.377
+ $X2=1.68 $Y2=1.377
r63 23 25 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.825 $Y=1.46
+ $X2=1.845 $Y2=1.46
r64 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.825
+ $Y=1.46 $X2=1.825 $Y2=1.46
r65 20 23 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.415 $Y=1.46
+ $X2=1.825 $Y2=1.46
r66 16 24 7.00744 $w=2.42e-07 $l=1.39e-07 $layer=LI1_cond $X=1.686 $Y=1.377
+ $X2=1.825 $Y2=1.377
r67 16 33 0.302479 $w=2.42e-07 $l=6e-09 $layer=LI1_cond $X=1.686 $Y=1.377
+ $X2=1.68 $Y2=1.377
r68 16 27 0.240809 $w=3.33e-07 $l=7e-09 $layer=LI1_cond $X=1.601 $Y=1.377
+ $X2=1.608 $Y2=1.377
r69 15 16 13.7949 $w=3.33e-07 $l=4.01e-07 $layer=LI1_cond $X=1.2 $Y=1.377
+ $X2=1.601 $Y2=1.377
r70 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.625
+ $X2=1.845 $Y2=1.46
r71 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.845 $Y=1.625
+ $X2=1.845 $Y2=2.465
r72 8 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.295
+ $X2=1.845 $Y2=1.46
r73 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.845 $Y=1.295
+ $X2=1.845 $Y2=0.765
r74 4 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.625
+ $X2=1.415 $Y2=1.46
r75 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.415 $Y=1.625
+ $X2=1.415 $Y2=2.465
r76 1 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.295
+ $X2=1.415 $Y2=1.46
r77 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.415 $Y=1.295
+ $X2=1.415 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%B1 3 7 9 11 12 14 15 16 17 28
c51 28 0 1.74432e-19 $X=3.29 $Y=1.35
c52 12 0 1.79774e-20 $X=3.38 $Y=1.185
r53 28 30 14.223 $w=3.05e-07 $l=9e-08 $layer=POLY_cond $X=3.29 $Y=1.35 $X2=3.38
+ $Y2=1.35
r54 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.29
+ $Y=1.35 $X2=3.29 $Y2=1.35
r55 26 28 53.7311 $w=3.05e-07 $l=3.4e-07 $layer=POLY_cond $X=2.95 $Y=1.35
+ $X2=3.29 $Y2=1.35
r56 25 26 38.718 $w=3.05e-07 $l=2.45e-07 $layer=POLY_cond $X=2.705 $Y=1.35
+ $X2=2.95 $Y2=1.35
r57 23 25 15.0131 $w=3.05e-07 $l=9.5e-08 $layer=POLY_cond $X=2.61 $Y=1.35
+ $X2=2.705 $Y2=1.35
r58 17 29 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.6 $Y=1.35 $X2=3.29
+ $Y2=1.35
r59 16 29 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.12 $Y=1.35
+ $X2=3.29 $Y2=1.35
r60 15 16 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.61 $Y=1.35
+ $X2=3.12 $Y2=1.35
r61 15 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.35 $X2=2.61 $Y2=1.35
r62 12 30 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.185
+ $X2=3.38 $Y2=1.35
r63 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.38 $Y=1.185
+ $X2=3.38 $Y2=0.655
r64 9 26 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.185
+ $X2=2.95 $Y2=1.35
r65 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.95 $Y=1.185
+ $X2=2.95 $Y2=0.655
r66 5 25 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.515
+ $X2=2.705 $Y2=1.35
r67 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.705 $Y=1.515
+ $X2=2.705 $Y2=2.465
r68 1 23 52.941 $w=3.05e-07 $l=4.09268e-07 $layer=POLY_cond $X=2.275 $Y=1.515
+ $X2=2.61 $Y2=1.35
r69 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.275 $Y=1.515
+ $X2=2.275 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%A2 1 3 6 8 10 13 15 16 24
c48 24 0 1.29415e-19 $X=4.24 $Y=1.35
c49 16 0 1.74432e-19 $X=4.56 $Y=1.295
r50 22 24 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.03 $Y=1.35
+ $X2=4.24 $Y2=1.35
r51 19 22 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.81 $Y=1.35
+ $X2=4.03 $Y2=1.35
r52 15 16 24.4318 $w=2.48e-07 $l=5.3e-07 $layer=LI1_cond $X=4.03 $Y=1.31
+ $X2=4.56 $Y2=1.31
r53 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.35 $X2=4.03 $Y2=1.35
r54 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.24 $Y=1.515
+ $X2=4.24 $Y2=1.35
r55 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.24 $Y=1.515
+ $X2=4.24 $Y2=2.465
r56 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.24 $Y=1.185
+ $X2=4.24 $Y2=1.35
r57 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.24 $Y=1.185
+ $X2=4.24 $Y2=0.655
r58 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.515
+ $X2=3.81 $Y2=1.35
r59 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.81 $Y=1.515 $X2=3.81
+ $Y2=2.465
r60 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.185
+ $X2=3.81 $Y2=1.35
r61 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.81 $Y=1.185 $X2=3.81
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%A1 1 3 6 8 10 13 15 16 24
c37 16 0 1.29415e-19 $X=5.52 $Y=1.295
c38 6 0 8.95735e-20 $X=4.67 $Y=2.465
r39 22 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.01 $Y=1.35 $X2=5.1
+ $Y2=1.35
r40 19 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.67 $Y=1.35
+ $X2=5.01 $Y2=1.35
r41 15 16 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=5.01 $Y=1.31
+ $X2=5.52 $Y2=1.31
r42 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.01
+ $Y=1.35 $X2=5.01 $Y2=1.35
r43 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.1 $Y=1.515
+ $X2=5.1 $Y2=1.35
r44 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.1 $Y=1.515 $X2=5.1
+ $Y2=2.465
r45 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.1 $Y=1.185 $X2=5.1
+ $Y2=1.35
r46 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.1 $Y=1.185 $X2=5.1
+ $Y2=0.655
r47 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.67 $Y=1.515
+ $X2=4.67 $Y2=1.35
r48 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.67 $Y=1.515 $X2=4.67
+ $Y2=2.465
r49 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.67 $Y=1.185
+ $X2=4.67 $Y2=1.35
r50 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.67 $Y=1.185 $X2=4.67
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%VPWR 1 2 3 4 5 16 18 24 30 36 42 47 48 50
+ 51 53 54 55 57 76 77 83
r84 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r85 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r86 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r87 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r88 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r89 71 74 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 70 73 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r93 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r95 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r96 62 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.2 $Y2=3.33
r97 62 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.68 $Y2=3.33
r98 61 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r99 61 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r100 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 58 80 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r102 58 60 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 57 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.2 $Y2=3.33
r104 57 60 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.72 $Y2=3.33
r105 55 71 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 55 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 53 73 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.72 $Y=3.33
+ $X2=4.56 $Y2=3.33
r108 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.72 $Y=3.33
+ $X2=4.885 $Y2=3.33
r109 52 76 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.05 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.05 $Y=3.33
+ $X2=4.885 $Y2=3.33
r111 50 67 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.92 $Y2=3.33
r113 49 70 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=2.92 $Y2=3.33
r115 47 64 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=2.06 $Y2=3.33
r117 46 67 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.06 $Y2=3.33
r119 42 45 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=4.885 $Y=2.03
+ $X2=4.885 $Y2=2.95
r120 40 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=3.245
+ $X2=4.885 $Y2=3.33
r121 40 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.885 $Y=3.245
+ $X2=4.885 $Y2=2.95
r122 36 39 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.92 $Y=2.11
+ $X2=2.92 $Y2=2.95
r123 34 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=3.33
r124 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=2.95
r125 30 33 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.06 $Y=2.18
+ $X2=2.06 $Y2=2.95
r126 28 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=3.245
+ $X2=2.06 $Y2=3.33
r127 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.06 $Y=3.245
+ $X2=2.06 $Y2=2.95
r128 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.2 $Y=2.18 $X2=1.2
+ $Y2=2.95
r129 22 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=3.245 $X2=1.2
+ $Y2=3.33
r130 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=3.245
+ $X2=1.2 $Y2=2.95
r131 18 21 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=0.3 $Y=2.09 $X2=0.3
+ $Y2=2.95
r132 16 80 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.212 $Y2=3.33
r133 16 21 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.3 $Y2=2.95
r134 5 45 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.835 $X2=4.885 $Y2=2.95
r135 5 42 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=4.745
+ $Y=1.835 $X2=4.885 $Y2=2.03
r136 4 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.835 $X2=2.92 $Y2=2.95
r137 4 36 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=1.835 $X2=2.92 $Y2=2.11
r138 3 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=2.95
r139 3 30 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=2.18
r140 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.835 $X2=1.2 $Y2=2.95
r141 2 24 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.835 $X2=1.2 $Y2=2.18
r142 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.95
r143 1 18 400 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.09
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%Y 1 2 3 4 5 18 24 26 30 34 38 42 46 51 52
+ 53 54 55 66
c69 54 0 2.47547e-19 $X=0.635 $Y=1.21
c70 42 0 8.95735e-20 $X=3.86 $Y=1.77
r71 59 66 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=0.765 $Y=1.335
+ $X2=0.765 $Y2=1.295
r72 54 66 0.779594 $w=3.38e-07 $l=2.3e-08 $layer=LI1_cond $X=0.765 $Y=1.272
+ $X2=0.765 $Y2=1.295
r73 54 64 3.62681 $w=3.38e-07 $l=1.07e-07 $layer=LI1_cond $X=0.765 $Y=1.272
+ $X2=0.765 $Y2=1.165
r74 54 55 10.4398 $w=3.38e-07 $l=3.08e-07 $layer=LI1_cond $X=0.765 $Y=1.357
+ $X2=0.765 $Y2=1.665
r75 54 59 0.745698 $w=3.38e-07 $l=2.2e-08 $layer=LI1_cond $X=0.765 $Y=1.357
+ $X2=0.765 $Y2=1.335
r76 50 55 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=0.765 $Y=1.755
+ $X2=0.765 $Y2=1.665
r77 50 51 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=1.755
+ $X2=0.765 $Y2=1.84
r78 46 48 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.025 $Y=1.97
+ $X2=4.025 $Y2=2.65
r79 44 46 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.025 $Y=1.855
+ $X2=4.025 $Y2=1.97
r80 43 53 5.41628 $w=1.7e-07 $l=1.11131e-07 $layer=LI1_cond $X=2.575 $Y=1.77
+ $X2=2.48 $Y2=1.805
r81 42 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.86 $Y=1.77
+ $X2=4.025 $Y2=1.855
r82 42 43 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=3.86 $Y=1.77
+ $X2=2.575 $Y2=1.77
r83 38 40 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=2.485 $Y=1.98
+ $X2=2.485 $Y2=2.91
r84 36 53 1.13756 $w=1.8e-07 $l=1.22474e-07 $layer=LI1_cond $X=2.485 $Y=1.925
+ $X2=2.48 $Y2=1.805
r85 36 38 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=2.485 $Y=1.925
+ $X2=2.485 $Y2=1.98
r86 35 52 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.725 $Y=1.84
+ $X2=1.63 $Y2=1.84
r87 34 53 5.41628 $w=1.7e-07 $l=1.11131e-07 $layer=LI1_cond $X=2.385 $Y=1.84
+ $X2=2.48 $Y2=1.805
r88 34 35 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.385 $Y=1.84
+ $X2=1.725 $Y2=1.84
r89 30 32 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.63 $Y=1.98
+ $X2=1.63 $Y2=2.91
r90 28 52 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=1.925
+ $X2=1.63 $Y2=1.84
r91 28 30 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.63 $Y=1.925
+ $X2=1.63 $Y2=1.98
r92 27 51 3.51065 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.935 $Y=1.84
+ $X2=0.765 $Y2=1.84
r93 26 52 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.535 $Y=1.84
+ $X2=1.63 $Y2=1.84
r94 26 27 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.535 $Y=1.84
+ $X2=0.935 $Y2=1.84
r95 24 64 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=0.77 $Y=0.68
+ $X2=0.77 $Y2=1.165
r96 18 20 39.6953 $w=2.68e-07 $l=9.3e-07 $layer=LI1_cond $X=0.73 $Y=1.98
+ $X2=0.73 $Y2=2.91
r97 16 51 3.10218 $w=3.05e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.73 $Y=1.925
+ $X2=0.765 $Y2=1.84
r98 16 18 2.34757 $w=2.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.73 $Y=1.925
+ $X2=0.73 $Y2=1.98
r99 5 48 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.835 $X2=4.025 $Y2=2.65
r100 5 46 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.835 $X2=4.025 $Y2=1.97
r101 4 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.835 $X2=2.49 $Y2=2.91
r102 4 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.35
+ $Y=1.835 $X2=2.49 $Y2=1.98
r103 3 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.835 $X2=1.63 $Y2=2.91
r104 3 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.835 $X2=1.63 $Y2=1.98
r105 2 20 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=2.91
r106 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=1.98
r107 1 24 91 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.345 $X2=0.77 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%A_694_367# 1 2 3 10 12 14 17 19 20 21 24
r42 24 26 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=5.35 $Y=1.98 $X2=5.35
+ $Y2=2.91
r43 22 24 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=5.35 $Y=1.775
+ $X2=5.35 $Y2=1.98
r44 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.22 $Y=1.69
+ $X2=5.35 $Y2=1.775
r45 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.22 $Y=1.69
+ $X2=4.55 $Y2=1.69
r46 17 31 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=2.905
+ $X2=4.455 $Y2=2.99
r47 17 19 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=4.455 $Y=2.905
+ $X2=4.455 $Y2=1.98
r48 16 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.455 $Y=1.775
+ $X2=4.55 $Y2=1.69
r49 16 19 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=4.455 $Y=1.775
+ $X2=4.455 $Y2=1.98
r50 15 29 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.69 $Y=2.99 $X2=3.56
+ $Y2=2.99
r51 14 31 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.36 $Y=2.99
+ $X2=4.455 $Y2=2.99
r52 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.36 $Y=2.99
+ $X2=3.69 $Y2=2.99
r53 10 29 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=2.905
+ $X2=3.56 $Y2=2.99
r54 10 12 31.6922 $w=2.58e-07 $l=7.15e-07 $layer=LI1_cond $X=3.56 $Y=2.905
+ $X2=3.56 $Y2=2.19
r55 3 26 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.175
+ $Y=1.835 $X2=5.315 $Y2=2.91
r56 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.175
+ $Y=1.835 $X2=5.315 $Y2=1.98
r57 2 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=1.835 $X2=4.455 $Y2=2.91
r58 2 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=1.835 $X2=4.455 $Y2=1.98
r59 1 29 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.835 $X2=3.595 $Y2=2.91
r60 1 12 400 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.835 $X2=3.595 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%A_43_69# 1 2 3 12 14 15 20 21 23
r36 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.11 $Y=0.68
+ $X2=2.11 $Y2=0.955
r37 20 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0.955
+ $X2=2.11 $Y2=0.955
r38 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.945 $Y=0.955
+ $X2=1.335 $Y2=0.955
r39 17 21 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.225 $Y=0.87
+ $X2=1.335 $Y2=0.955
r40 17 19 19.9058 $w=2.18e-07 $l=3.8e-07 $layer=LI1_cond $X=1.225 $Y=0.87
+ $X2=1.225 $Y2=0.49
r41 16 19 3.40495 $w=2.18e-07 $l=6.5e-08 $layer=LI1_cond $X=1.225 $Y=0.425
+ $X2=1.225 $Y2=0.49
r42 14 16 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.115 $Y=0.34
+ $X2=1.225 $Y2=0.425
r43 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.115 $Y=0.34
+ $X2=0.435 $Y2=0.34
r44 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.305 $Y=0.425
+ $X2=0.435 $Y2=0.34
r45 10 12 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.305 $Y=0.425
+ $X2=0.305 $Y2=0.49
r46 3 23 91 $w=1.7e-07 $l=4.19375e-07 $layer=licon1_NDIFF $count=2 $X=1.92
+ $Y=0.345 $X2=2.11 $Y2=0.68
r47 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.06
+ $Y=0.345 $X2=1.2 $Y2=0.49
r48 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.215
+ $Y=0.345 $X2=0.34 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%A_298_69# 1 2 9 11 12 13
c26 11 0 1.79774e-20 $X=3 $Y=0.34
r27 13 16 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.165 $Y=0.34
+ $X2=3.165 $Y2=0.48
r28 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3 $Y=0.34 $X2=3.165
+ $Y2=0.34
r29 11 12 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=3 $Y=0.34
+ $X2=1.775 $Y2=0.34
r30 7 12 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.64 $Y=0.425
+ $X2=1.775 $Y2=0.34
r31 7 9 4.69514 $w=2.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.64 $Y=0.425 $X2=1.64
+ $Y2=0.535
r32 2 16 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.235 $X2=3.165 $Y2=0.48
r33 1 9 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.345 $X2=1.63 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%A_522_47# 1 2 3 4 13 19 21 25 27 29 31 34
+ 36
r43 29 38 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.35 $Y=0.845
+ $X2=5.35 $Y2=0.93
r44 29 31 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=5.35 $Y=0.845
+ $X2=5.35 $Y2=0.42
r45 28 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.55 $Y=0.93
+ $X2=4.455 $Y2=0.93
r46 27 38 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.22 $Y=0.93 $X2=5.35
+ $Y2=0.93
r47 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.22 $Y=0.93
+ $X2=4.55 $Y2=0.93
r48 23 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=0.845
+ $X2=4.455 $Y2=0.93
r49 23 25 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=4.455 $Y=0.845
+ $X2=4.455 $Y2=0.42
r50 22 34 4.84724 $w=2.05e-07 $l=1.11131e-07 $layer=LI1_cond $X=3.69 $Y=0.93
+ $X2=3.595 $Y2=0.895
r51 21 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.36 $Y=0.93
+ $X2=4.455 $Y2=0.93
r52 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.36 $Y=0.93
+ $X2=3.69 $Y2=0.93
r53 17 34 1.61756 $w=1.9e-07 $l=1.2e-07 $layer=LI1_cond $X=3.595 $Y=0.775
+ $X2=3.595 $Y2=0.895
r54 17 19 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=3.595 $Y=0.775
+ $X2=3.595 $Y2=0.42
r55 13 34 4.84724 $w=2.05e-07 $l=9.5e-08 $layer=LI1_cond $X=3.5 $Y=0.895
+ $X2=3.595 $Y2=0.895
r56 13 15 36.7341 $w=2.38e-07 $l=7.65e-07 $layer=LI1_cond $X=3.5 $Y=0.895
+ $X2=2.735 $Y2=0.895
r57 4 38 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=5.175
+ $Y=0.235 $X2=5.315 $Y2=0.93
r58 4 31 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.175
+ $Y=0.235 $X2=5.315 $Y2=0.42
r59 3 36 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=4.315
+ $Y=0.235 $X2=4.455 $Y2=0.93
r60 3 25 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.315
+ $Y=0.235 $X2=4.455 $Y2=0.42
r61 2 34 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.235 $X2=3.595 $Y2=0.93
r62 2 19 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.235 $X2=3.595 $Y2=0.42
r63 1 15 182 $w=1.7e-07 $l=7.04734e-07 $layer=licon1_NDIFF $count=1 $X=2.61
+ $Y=0.235 $X2=2.735 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_2%VGND 1 2 9 13 16 17 18 20 33 34 37
r63 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r64 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r65 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r66 31 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r67 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r68 28 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=4.025
+ $Y2=0
r69 28 30 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.19 $Y=0 $X2=4.56
+ $Y2=0
r70 27 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r71 26 27 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r72 22 26 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r73 22 23 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r74 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.86 $Y=0 $X2=4.025
+ $Y2=0
r75 20 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.86 $Y=0 $X2=3.6
+ $Y2=0
r76 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r77 18 23 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=0.24
+ $Y2=0
r78 16 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.72 $Y=0 $X2=4.56
+ $Y2=0
r79 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.72 $Y=0 $X2=4.885
+ $Y2=0
r80 15 33 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.05 $Y=0 $X2=5.52
+ $Y2=0
r81 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.05 $Y=0 $X2=4.885
+ $Y2=0
r82 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.885 $Y=0.085
+ $X2=4.885 $Y2=0
r83 11 13 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.885 $Y=0.085
+ $X2=4.885 $Y2=0.55
r84 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.025 $Y=0.085
+ $X2=4.025 $Y2=0
r85 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.025 $Y=0.085
+ $X2=4.025 $Y2=0.55
r86 2 13 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=4.745
+ $Y=0.235 $X2=4.885 $Y2=0.55
r87 1 9 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.025 $Y2=0.55
.ends

