* File: sky130_fd_sc_lp__nand4b_2.spice
* Created: Wed Sep  2 10:06:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4b_2.pex.spice"
.subckt sky130_fd_sc_lp__nand4b_2  VNB VPB A_N B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_N_M1013_g N_A_27_51#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_217_65#_M1002_d N_A_27_51#_M1002_g N_Y_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1009 N_A_217_65#_M1009_d N_A_27_51#_M1009_g N_Y_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_486_65#_M1000_d N_B_M1000_g N_A_217_65#_M1009_d VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1016 N_A_486_65#_M1000_d N_B_M1016_g N_A_217_65#_M1016_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.2226 PD=1.19 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_A_486_65#_M1006_d N_C_M1006_g N_A_697_69#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2898 PD=1.12 PS=2.37 NRD=0 NRS=11.424 M=1 R=5.6
+ SA=75000.3 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1012 N_A_486_65#_M1006_d N_C_M1012_g N_A_697_69#_M1012_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_D_M1005_g N_A_697_69#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1218 AS=0.1176 PD=1.13 PS=1.12 NRD=1.428 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1005_d N_D_M1014_g N_A_697_69#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1218 AS=0.2226 PD=1.13 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VPWR_M1010_d N_A_N_M1010_g N_A_27_51#_M1010_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.109725 AS=0.1113 PD=0.8675 PS=1.37 NRD=11.7215 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75004.6 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A_27_51#_M1003_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.329175 PD=1.54 PS=2.6025 NRD=0 NRS=8.8453 M=1 R=8.4 SA=75000.4
+ SB=75004 A=0.189 P=2.82 MULT=1
MM1015 N_Y_M1003_d N_A_27_51#_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2205 PD=1.54 PS=1.61 NRD=0 NRS=5.4569 M=1 R=8.4 SA=75000.8
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1827 AS=0.2205 PD=1.55 PS=1.61 NRD=1.5563 NRS=5.4569 M=1 R=8.4 SA=75001.3
+ SB=75003 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1001_d N_B_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1827 AS=0.6048 PD=1.55 PS=2.22 NRD=0 NRS=0 M=1 R=8.4 SA=75001.8
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1008_s N_C_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.6048 AS=0.1764 PD=2.22 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_C_M1011_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1011_d N_D_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_D_M1017_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__nand4b_2.pxi.spice"
*
.ends
*
*
