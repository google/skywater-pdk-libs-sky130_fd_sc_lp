* File: sky130_fd_sc_lp__dlclkp_4.pxi.spice
* Created: Wed Sep  2 09:45:54 2020
* 
x_PM_SKY130_FD_SC_LP__DLCLKP_4%A_73_269# N_A_73_269#_M1001_d N_A_73_269#_M1020_d
+ N_A_73_269#_M1025_g N_A_73_269#_M1022_g N_A_73_269#_c_170_n
+ N_A_73_269#_c_178_n N_A_73_269#_c_171_n N_A_73_269#_c_180_n
+ N_A_73_269#_c_187_p N_A_73_269#_c_172_n N_A_73_269#_c_173_n
+ N_A_73_269#_c_174_n N_A_73_269#_c_191_p N_A_73_269#_c_175_n
+ N_A_73_269#_c_183_n PM_SKY130_FD_SC_LP__DLCLKP_4%A_73_269#
x_PM_SKY130_FD_SC_LP__DLCLKP_4%GATE N_GATE_M1006_g N_GATE_M1009_g GATE
+ N_GATE_c_282_n PM_SKY130_FD_SC_LP__DLCLKP_4%GATE
x_PM_SKY130_FD_SC_LP__DLCLKP_4%A_277_367# N_A_277_367#_M1008_d
+ N_A_277_367#_M1021_d N_A_277_367#_M1020_g N_A_277_367#_M1014_g
+ N_A_277_367#_c_340_n N_A_277_367#_c_341_n N_A_277_367#_c_333_n
+ N_A_277_367#_c_334_n N_A_277_367#_c_343_n N_A_277_367#_c_335_n
+ N_A_277_367#_c_344_n N_A_277_367#_c_336_n N_A_277_367#_c_346_n
+ N_A_277_367#_c_337_n N_A_277_367#_c_347_n N_A_277_367#_c_338_n
+ PM_SKY130_FD_SC_LP__DLCLKP_4%A_277_367#
x_PM_SKY130_FD_SC_LP__DLCLKP_4%A_295_55# N_A_295_55#_M1024_s N_A_295_55#_M1012_s
+ N_A_295_55#_M1001_g N_A_295_55#_c_463_n N_A_295_55#_c_464_n
+ N_A_295_55#_M1007_g N_A_295_55#_M1008_g N_A_295_55#_c_466_n
+ N_A_295_55#_M1021_g N_A_295_55#_c_468_n N_A_295_55#_c_469_n
+ N_A_295_55#_c_470_n N_A_295_55#_c_471_n N_A_295_55#_c_472_n
+ N_A_295_55#_c_543_p N_A_295_55#_c_473_n N_A_295_55#_c_474_n
+ N_A_295_55#_c_475_n PM_SKY130_FD_SC_LP__DLCLKP_4%A_295_55#
x_PM_SKY130_FD_SC_LP__DLCLKP_4%A_27_367# N_A_27_367#_M1022_s N_A_27_367#_M1025_s
+ N_A_27_367#_M1011_g N_A_27_367#_M1010_g N_A_27_367#_c_590_n
+ N_A_27_367#_c_591_n N_A_27_367#_c_576_n N_A_27_367#_M1002_g
+ N_A_27_367#_M1017_g N_A_27_367#_c_577_n N_A_27_367#_c_610_n
+ N_A_27_367#_c_578_n N_A_27_367#_c_618_n N_A_27_367#_c_579_n
+ N_A_27_367#_c_580_n N_A_27_367#_c_593_n N_A_27_367#_c_594_n
+ N_A_27_367#_c_595_n N_A_27_367#_c_596_n N_A_27_367#_c_581_n
+ N_A_27_367#_c_672_n N_A_27_367#_c_597_n N_A_27_367#_c_598_n
+ N_A_27_367#_c_599_n N_A_27_367#_c_582_n N_A_27_367#_c_600_n
+ N_A_27_367#_c_583_n N_A_27_367#_c_602_n N_A_27_367#_c_603_n
+ N_A_27_367#_c_604_n N_A_27_367#_c_584_n N_A_27_367#_c_585_n
+ N_A_27_367#_c_605_n N_A_27_367#_c_606_n N_A_27_367#_c_607_n
+ N_A_27_367#_c_586_n N_A_27_367#_c_587_n N_A_27_367#_c_588_n
+ PM_SKY130_FD_SC_LP__DLCLKP_4%A_27_367#
x_PM_SKY130_FD_SC_LP__DLCLKP_4%CLK N_CLK_c_822_n N_CLK_M1024_g N_CLK_M1012_g
+ N_CLK_c_824_n N_CLK_c_825_n N_CLK_M1005_g N_CLK_M1000_g N_CLK_c_827_n CLK
+ N_CLK_c_828_n N_CLK_c_829_n PM_SKY130_FD_SC_LP__DLCLKP_4%CLK
x_PM_SKY130_FD_SC_LP__DLCLKP_4%A_1078_367# N_A_1078_367#_M1002_d
+ N_A_1078_367#_M1000_d N_A_1078_367#_M1003_g N_A_1078_367#_M1004_g
+ N_A_1078_367#_M1016_g N_A_1078_367#_M1013_g N_A_1078_367#_M1018_g
+ N_A_1078_367#_M1015_g N_A_1078_367#_M1023_g N_A_1078_367#_M1019_g
+ N_A_1078_367#_c_902_n N_A_1078_367#_c_903_n N_A_1078_367#_c_904_n
+ N_A_1078_367#_c_905_n N_A_1078_367#_c_968_p N_A_1078_367#_c_906_n
+ N_A_1078_367#_c_918_n N_A_1078_367#_c_907_n
+ PM_SKY130_FD_SC_LP__DLCLKP_4%A_1078_367#
x_PM_SKY130_FD_SC_LP__DLCLKP_4%VPWR N_VPWR_M1025_d N_VPWR_M1011_d N_VPWR_M1012_d
+ N_VPWR_M1017_d N_VPWR_M1016_d N_VPWR_M1023_d N_VPWR_c_1018_n N_VPWR_c_1019_n
+ N_VPWR_c_1020_n N_VPWR_c_1021_n N_VPWR_c_1022_n N_VPWR_c_1023_n
+ N_VPWR_c_1024_n N_VPWR_c_1025_n VPWR N_VPWR_c_1026_n N_VPWR_c_1027_n
+ N_VPWR_c_1028_n N_VPWR_c_1029_n N_VPWR_c_1030_n N_VPWR_c_1031_n
+ N_VPWR_c_1032_n N_VPWR_c_1033_n N_VPWR_c_1034_n N_VPWR_c_1017_n
+ PM_SKY130_FD_SC_LP__DLCLKP_4%VPWR
x_PM_SKY130_FD_SC_LP__DLCLKP_4%GCLK N_GCLK_M1004_d N_GCLK_M1015_d N_GCLK_M1003_s
+ N_GCLK_M1018_s N_GCLK_c_1134_n N_GCLK_c_1168_n N_GCLK_c_1178_p N_GCLK_c_1135_n
+ N_GCLK_c_1130_n N_GCLK_c_1131_n GCLK GCLK GCLK GCLK GCLK GCLK GCLK
+ N_GCLK_c_1179_p GCLK GCLK PM_SKY130_FD_SC_LP__DLCLKP_4%GCLK
x_PM_SKY130_FD_SC_LP__DLCLKP_4%VGND N_VGND_M1022_d N_VGND_M1010_d N_VGND_M1024_d
+ N_VGND_M1004_s N_VGND_M1013_s N_VGND_M1019_s N_VGND_c_1184_n N_VGND_c_1185_n
+ N_VGND_c_1186_n N_VGND_c_1187_n N_VGND_c_1188_n N_VGND_c_1189_n
+ N_VGND_c_1190_n N_VGND_c_1191_n N_VGND_c_1192_n N_VGND_c_1193_n
+ N_VGND_c_1194_n VGND N_VGND_c_1195_n N_VGND_c_1196_n N_VGND_c_1197_n
+ N_VGND_c_1198_n N_VGND_c_1199_n N_VGND_c_1200_n N_VGND_c_1201_n
+ N_VGND_c_1202_n PM_SKY130_FD_SC_LP__DLCLKP_4%VGND
cc_1 VNB N_A_73_269#_M1022_g 0.0328734f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_2 VNB N_A_73_269#_c_170_n 0.00371539f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.645
cc_3 VNB N_A_73_269#_c_171_n 0.00649833f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.645
cc_4 VNB N_A_73_269#_c_172_n 0.00527326f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=1.56
cc_5 VNB N_A_73_269#_c_173_n 0.0013439f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.51
cc_6 VNB N_A_73_269#_c_174_n 0.0287634f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.51
cc_7 VNB N_A_73_269#_c_175_n 0.00318387f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.7
cc_8 VNB N_GATE_M1006_g 0.0103457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_GATE_M1009_g 0.0272293f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.675
cc_10 VNB GATE 0.00708601f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_11 VNB N_GATE_c_282_n 0.0299915f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_12 VNB N_A_277_367#_c_333_n 0.0093868f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=2.365
cc_13 VNB N_A_277_367#_c_334_n 0.0307991f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=2.365
cc_14 VNB N_A_277_367#_c_335_n 0.024912f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.51
cc_15 VNB N_A_277_367#_c_336_n 0.00376562f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.645
cc_16 VNB N_A_277_367#_c_337_n 0.00754367f $X=-0.19 $Y=-0.245 $X2=1.765
+ $Y2=0.725
cc_17 VNB N_A_277_367#_c_338_n 0.0158201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_295_55#_M1001_g 0.0411015f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_19 VNB N_A_295_55#_c_463_n 0.0186698f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.345
cc_20 VNB N_A_295_55#_c_464_n 0.00658555f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_21 VNB N_A_295_55#_M1008_g 0.0267819f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.645
cc_22 VNB N_A_295_55#_c_466_n 0.0352379f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=2.365
cc_23 VNB N_A_295_55#_M1021_g 4.71742e-19 $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.51
cc_24 VNB N_A_295_55#_c_468_n 0.00524433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_295_55#_c_469_n 0.0185878f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.645
cc_26 VNB N_A_295_55#_c_470_n 0.00803153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_295_55#_c_471_n 0.0293998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_295_55#_c_472_n 0.00456253f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.7
cc_29 VNB N_A_295_55#_c_473_n 0.0235859f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.365
cc_30 VNB N_A_295_55#_c_474_n 0.00818795f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.345
cc_31 VNB N_A_295_55#_c_475_n 0.0198518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_367#_c_576_n 0.0188874f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.645
cc_33 VNB N_A_27_367#_c_577_n 0.022836f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.51
cc_34 VNB N_A_27_367#_c_578_n 0.00592274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_367#_c_579_n 0.00941734f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.365
cc_36 VNB N_A_27_367#_c_580_n 0.00226982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_367#_c_581_n 0.00195788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_367#_c_582_n 0.0153942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_367#_c_583_n 0.026445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_367#_c_584_n 0.00347572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_367#_c_585_n 0.0332952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_367#_c_586_n 0.00394158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_367#_c_587_n 0.0170569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_367#_c_588_n 0.0544988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_CLK_c_822_n 0.0182783f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=0.405
cc_46 VNB N_CLK_M1024_g 0.044696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_CLK_c_824_n 0.00582738f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.345
cc_48 VNB N_CLK_c_825_n 0.00555802f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_49 VNB N_CLK_M1005_g 0.0370948f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.645
cc_50 VNB N_CLK_c_827_n 0.0154747f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=1.56
cc_51 VNB N_CLK_c_828_n 0.0278177f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.645
cc_52 VNB N_CLK_c_829_n 0.00590275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1078_367#_M1004_g 0.0265717f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_54 VNB N_A_1078_367#_M1013_g 0.0221671f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=2.365
cc_55 VNB N_A_1078_367#_M1015_g 0.0221495f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.645
cc_56 VNB N_A_1078_367#_M1019_g 0.033551f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.365
cc_57 VNB N_A_1078_367#_c_902_n 0.00403192f $X=-0.19 $Y=-0.245 $X2=1.675
+ $Y2=2.57
cc_58 VNB N_A_1078_367#_c_903_n 0.00849941f $X=-0.19 $Y=-0.245 $X2=0.53
+ $Y2=1.345
cc_59 VNB N_A_1078_367#_c_904_n 0.0129573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1078_367#_c_905_n 9.81998e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1078_367#_c_906_n 9.62967e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1078_367#_c_907_n 0.0942101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VPWR_c_1017_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_GCLK_c_1130_n 0.00883403f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=0.845
cc_65 VNB N_GCLK_c_1131_n 0.00270021f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=1.56
cc_66 VNB GCLK 0.00202901f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.645
cc_67 VNB GCLK 0.00162609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1184_n 0.00498979f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=2.365
cc_69 VNB N_VGND_c_1185_n 0.00737153f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.51
cc_70 VNB N_VGND_c_1186_n 0.011127f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.645
cc_71 VNB N_VGND_c_1187_n 0.0091336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1188_n 3.15212e-19 $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.365
cc_73 VNB N_VGND_c_1189_n 0.0118625f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.57
cc_74 VNB N_VGND_c_1190_n 0.0496322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1191_n 0.0436536f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.675
cc_76 VNB N_VGND_c_1192_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1193_n 0.0474805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1194_n 0.00510065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1195_n 0.0159362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1196_n 0.0265259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1197_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1198_n 0.0151004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1199_n 0.00532666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1200_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1201_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1202_n 0.440151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VPB N_A_73_269#_M1025_g 0.0256927f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_88 VPB N_A_73_269#_c_170_n 0.0117834f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=1.645
cc_89 VPB N_A_73_269#_c_178_n 0.00524258f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.28
cc_90 VPB N_A_73_269#_c_171_n 0.00448359f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=1.645
cc_91 VPB N_A_73_269#_c_180_n 0.00239821f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=2.365
cc_92 VPB N_A_73_269#_c_173_n 0.00520645f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.51
cc_93 VPB N_A_73_269#_c_174_n 0.0064633f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.51
cc_94 VPB N_A_73_269#_c_183_n 0.00243281f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=2.365
cc_95 VPB N_GATE_M1006_g 0.0491402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_277_367#_M1020_g 0.0206495f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_97 VPB N_A_277_367#_c_340_n 0.00369331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_277_367#_c_341_n 0.0303421f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=1.73
cc_99 VPB N_A_277_367#_c_333_n 0.00607322f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=2.365
cc_100 VPB N_A_277_367#_c_343_n 0.0170156f $X=-0.19 $Y=1.655 $X2=1.57 $Y2=1.56
cc_101 VPB N_A_277_367#_c_344_n 0.013976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_277_367#_c_336_n 8.49111e-19 $X=-0.19 $Y=1.655 $X2=1.12 $Y2=1.645
cc_103 VPB N_A_277_367#_c_346_n 0.00569004f $X=-0.19 $Y=1.655 $X2=1.57 $Y2=0.725
cc_104 VPB N_A_277_367#_c_347_n 0.0136545f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=2.57
cc_105 VPB N_A_295_55#_M1007_g 0.0412229f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=1.645
cc_106 VPB N_A_295_55#_M1021_g 0.0451233f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.51
cc_107 VPB N_A_295_55#_c_468_n 0.00666874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_295_55#_c_470_n 0.00423362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_295_55#_c_471_n 0.0270967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_295_55#_c_474_n 0.009112f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.345
cc_111 VPB N_A_27_367#_M1011_g 0.0307828f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_112 VPB N_A_27_367#_c_590_n 0.0958705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_27_367#_c_591_n 0.012806f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=1.645
cc_114 VPB N_A_27_367#_M1017_g 0.0191284f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=2.365
cc_115 VPB N_A_27_367#_c_593_n 0.0118667f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=2.57
cc_116 VPB N_A_27_367#_c_594_n 0.00153612f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.51
cc_117 VPB N_A_27_367#_c_595_n 0.0014437f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.345
cc_118 VPB N_A_27_367#_c_596_n 8.23242e-19 $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.675
cc_119 VPB N_A_27_367#_c_597_n 0.00136158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_27_367#_c_598_n 0.00597134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_27_367#_c_599_n 0.00171165f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_27_367#_c_600_n 0.00638732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_27_367#_c_583_n 0.011126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_27_367#_c_602_n 0.0175711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_27_367#_c_603_n 0.0217943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_27_367#_c_604_n 9.93719e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_27_367#_c_605_n 0.0579381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_27_367#_c_606_n 0.0117437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_27_367#_c_607_n 0.0227564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_27_367#_c_586_n 2.77223e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_27_367#_c_588_n 0.00677073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_CLK_c_822_n 0.0228082f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=0.405
cc_133 VPB N_CLK_M1012_g 0.0213344f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_134 VPB N_CLK_c_824_n 0.00428214f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.345
cc_135 VPB N_CLK_c_825_n 0.00880555f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.655
cc_136 VPB N_CLK_M1000_g 0.0206911f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=1.645
cc_137 VPB N_CLK_c_827_n 0.00881687f $X=-0.19 $Y=1.655 $X2=1.57 $Y2=1.56
cc_138 VPB N_CLK_c_828_n 0.0112695f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.645
cc_139 VPB N_CLK_c_829_n 0.00620348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_1078_367#_M1003_g 0.0199827f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=2.465
cc_141 VPB N_A_1078_367#_M1016_g 0.0188338f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=1.73
cc_142 VPB N_A_1078_367#_M1018_g 0.0188073f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.51
cc_143 VPB N_A_1078_367#_M1023_g 0.0256595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_1078_367#_c_902_n 0.00144814f $X=-0.19 $Y=1.655 $X2=1.675
+ $Y2=2.57
cc_145 VPB N_A_1078_367#_c_907_n 0.00999708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_1018_n 0.00448502f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=2.365
cc_147 VPB N_VPWR_c_1019_n 0.00824156f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.51
cc_148 VPB N_VPWR_c_1020_n 0.00210998f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.645
cc_149 VPB N_VPWR_c_1021_n 4.06069e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_1022_n 0.0135196f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=2.365
cc_151 VPB N_VPWR_c_1023_n 0.0625673f $X=-0.19 $Y=1.655 $X2=1.675 $Y2=2.57
cc_152 VPB N_VPWR_c_1024_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.675
cc_153 VPB N_VPWR_c_1025_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_1026_n 0.0171749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_1027_n 0.0381674f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_1028_n 0.0463348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_1029_n 0.0160917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_1030_n 0.0171979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_1031_n 0.0120341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_1032_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1033_n 0.00631534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1034_n 0.00510217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1017_n 0.0671343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_GCLK_c_1134_n 0.0022405f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.655
cc_165 VPB N_GCLK_c_1135_n 0.00353551f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=2.365
cc_166 VPB GCLK 0.00163723f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=1.645
cc_167 VPB GCLK 0.00147694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 N_A_73_269#_M1025_g N_GATE_M1006_g 0.0311052f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_73_269#_c_170_n N_GATE_M1006_g 0.0029792f $X=1.035 $Y=1.645 $X2=0
+ $Y2=0
cc_170 N_A_73_269#_c_178_n N_GATE_M1006_g 0.0175803f $X=1.12 $Y=2.28 $X2=0 $Y2=0
cc_171 N_A_73_269#_c_187_p N_GATE_M1006_g 0.00820898f $X=1.205 $Y=2.365 $X2=0
+ $Y2=0
cc_172 N_A_73_269#_c_172_n N_GATE_M1006_g 6.00478e-19 $X=1.57 $Y=1.56 $X2=0
+ $Y2=0
cc_173 N_A_73_269#_c_173_n N_GATE_M1006_g 7.16539e-19 $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_174 N_A_73_269#_c_174_n N_GATE_M1006_g 0.00821482f $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_175 N_A_73_269#_c_191_p N_GATE_M1006_g 0.00741923f $X=1.12 $Y=1.645 $X2=0
+ $Y2=0
cc_176 N_A_73_269#_c_183_n N_GATE_M1006_g 0.00107299f $X=1.675 $Y=2.365 $X2=0
+ $Y2=0
cc_177 N_A_73_269#_M1022_g N_GATE_M1009_g 0.0120262f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_178 N_A_73_269#_c_172_n N_GATE_M1009_g 0.0016161f $X=1.57 $Y=1.56 $X2=0 $Y2=0
cc_179 N_A_73_269#_c_175_n N_GATE_M1009_g 7.28749e-19 $X=1.765 $Y=0.7 $X2=0
+ $Y2=0
cc_180 N_A_73_269#_M1022_g GATE 0.00174603f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_181 N_A_73_269#_c_170_n GATE 0.013362f $X=1.035 $Y=1.645 $X2=0 $Y2=0
cc_182 N_A_73_269#_c_171_n GATE 0.00817592f $X=1.485 $Y=1.645 $X2=0 $Y2=0
cc_183 N_A_73_269#_c_172_n GATE 0.0170086f $X=1.57 $Y=1.56 $X2=0 $Y2=0
cc_184 N_A_73_269#_c_173_n GATE 0.00352441f $X=0.53 $Y=1.51 $X2=0 $Y2=0
cc_185 N_A_73_269#_c_174_n GATE 2.79937e-19 $X=0.53 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A_73_269#_c_191_p GATE 0.0133189f $X=1.12 $Y=1.645 $X2=0 $Y2=0
cc_187 N_A_73_269#_M1022_g N_GATE_c_282_n 0.00678312f $X=0.5 $Y=0.655 $X2=0
+ $Y2=0
cc_188 N_A_73_269#_c_170_n N_GATE_c_282_n 0.00219188f $X=1.035 $Y=1.645 $X2=0
+ $Y2=0
cc_189 N_A_73_269#_c_171_n N_GATE_c_282_n 0.0017138f $X=1.485 $Y=1.645 $X2=0
+ $Y2=0
cc_190 N_A_73_269#_c_172_n N_GATE_c_282_n 7.42469e-19 $X=1.57 $Y=1.56 $X2=0
+ $Y2=0
cc_191 N_A_73_269#_c_173_n N_GATE_c_282_n 5.33158e-19 $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_192 N_A_73_269#_c_174_n N_GATE_c_282_n 0.00649561f $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_193 N_A_73_269#_c_191_p N_GATE_c_282_n 8.88538e-19 $X=1.12 $Y=1.645 $X2=0
+ $Y2=0
cc_194 N_A_73_269#_c_180_n N_A_277_367#_M1020_g 0.00862793f $X=1.51 $Y=2.365
+ $X2=0 $Y2=0
cc_195 N_A_73_269#_c_183_n N_A_277_367#_M1020_g 0.00702773f $X=1.675 $Y=2.365
+ $X2=0 $Y2=0
cc_196 N_A_73_269#_c_178_n N_A_277_367#_c_340_n 0.0159151f $X=1.12 $Y=2.28 $X2=0
+ $Y2=0
cc_197 N_A_73_269#_c_171_n N_A_277_367#_c_340_n 0.0211323f $X=1.485 $Y=1.645
+ $X2=0 $Y2=0
cc_198 N_A_73_269#_c_180_n N_A_277_367#_c_340_n 0.00861249f $X=1.51 $Y=2.365
+ $X2=0 $Y2=0
cc_199 N_A_73_269#_c_183_n N_A_277_367#_c_340_n 0.0259437f $X=1.675 $Y=2.365
+ $X2=0 $Y2=0
cc_200 N_A_73_269#_c_178_n N_A_277_367#_c_341_n 0.0046394f $X=1.12 $Y=2.28 $X2=0
+ $Y2=0
cc_201 N_A_73_269#_c_171_n N_A_277_367#_c_341_n 0.00384696f $X=1.485 $Y=1.645
+ $X2=0 $Y2=0
cc_202 N_A_73_269#_c_183_n N_A_277_367#_c_341_n 0.00442109f $X=1.675 $Y=2.365
+ $X2=0 $Y2=0
cc_203 N_A_73_269#_c_178_n N_A_277_367#_c_333_n 0.00534813f $X=1.12 $Y=2.28
+ $X2=0 $Y2=0
cc_204 N_A_73_269#_c_171_n N_A_277_367#_c_333_n 0.0138732f $X=1.485 $Y=1.645
+ $X2=0 $Y2=0
cc_205 N_A_73_269#_c_172_n N_A_277_367#_c_333_n 0.0397522f $X=1.57 $Y=1.56 $X2=0
+ $Y2=0
cc_206 N_A_73_269#_c_175_n N_A_277_367#_c_333_n 0.00760456f $X=1.765 $Y=0.7
+ $X2=0 $Y2=0
cc_207 N_A_73_269#_c_172_n N_A_277_367#_c_334_n 0.00293536f $X=1.57 $Y=1.56
+ $X2=0 $Y2=0
cc_208 N_A_73_269#_c_175_n N_A_277_367#_c_334_n 0.00175689f $X=1.765 $Y=0.7
+ $X2=0 $Y2=0
cc_209 N_A_73_269#_c_172_n N_A_277_367#_c_338_n 0.00168714f $X=1.57 $Y=1.56
+ $X2=0 $Y2=0
cc_210 N_A_73_269#_c_175_n N_A_277_367#_c_338_n 0.00454263f $X=1.765 $Y=0.7
+ $X2=0 $Y2=0
cc_211 N_A_73_269#_c_172_n N_A_295_55#_M1001_g 0.0178635f $X=1.57 $Y=1.56 $X2=0
+ $Y2=0
cc_212 N_A_73_269#_c_175_n N_A_295_55#_M1001_g 0.00718883f $X=1.765 $Y=0.7 $X2=0
+ $Y2=0
cc_213 N_A_73_269#_c_171_n N_A_295_55#_c_463_n 0.00127817f $X=1.485 $Y=1.645
+ $X2=0 $Y2=0
cc_214 N_A_73_269#_c_172_n N_A_295_55#_c_463_n 0.00206217f $X=1.57 $Y=1.56 $X2=0
+ $Y2=0
cc_215 N_A_73_269#_c_175_n N_A_295_55#_c_463_n 0.00407379f $X=1.765 $Y=0.7 $X2=0
+ $Y2=0
cc_216 N_A_73_269#_c_171_n N_A_295_55#_c_464_n 0.00278327f $X=1.485 $Y=1.645
+ $X2=0 $Y2=0
cc_217 N_A_73_269#_c_172_n N_A_295_55#_c_464_n 0.00220328f $X=1.57 $Y=1.56 $X2=0
+ $Y2=0
cc_218 N_A_73_269#_c_183_n N_A_295_55#_M1007_g 0.00385189f $X=1.675 $Y=2.365
+ $X2=0 $Y2=0
cc_219 N_A_73_269#_c_171_n N_A_295_55#_c_468_n 6.5424e-19 $X=1.485 $Y=1.645
+ $X2=0 $Y2=0
cc_220 N_A_73_269#_M1025_g N_A_27_367#_c_610_n 0.0124839f $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_221 N_A_73_269#_c_187_p N_A_27_367#_c_610_n 0.0058194f $X=1.205 $Y=2.365
+ $X2=0 $Y2=0
cc_222 N_A_73_269#_M1022_g N_A_27_367#_c_578_n 0.0108351f $X=0.5 $Y=0.655 $X2=0
+ $Y2=0
cc_223 N_A_73_269#_c_170_n N_A_27_367#_c_578_n 0.005326f $X=1.035 $Y=1.645 $X2=0
+ $Y2=0
cc_224 N_A_73_269#_c_172_n N_A_27_367#_c_578_n 0.0085263f $X=1.57 $Y=1.56 $X2=0
+ $Y2=0
cc_225 N_A_73_269#_c_173_n N_A_27_367#_c_578_n 0.00864524f $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_226 N_A_73_269#_c_174_n N_A_27_367#_c_578_n 7.34064e-19 $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_227 N_A_73_269#_c_175_n N_A_27_367#_c_578_n 8.27727e-19 $X=1.765 $Y=0.7 $X2=0
+ $Y2=0
cc_228 N_A_73_269#_M1022_g N_A_27_367#_c_618_n 3.7394e-19 $X=0.5 $Y=0.655 $X2=0
+ $Y2=0
cc_229 N_A_73_269#_c_175_n N_A_27_367#_c_618_n 0.0118715f $X=1.765 $Y=0.7 $X2=0
+ $Y2=0
cc_230 N_A_73_269#_M1001_d N_A_27_367#_c_579_n 0.00174403f $X=1.625 $Y=0.405
+ $X2=0 $Y2=0
cc_231 N_A_73_269#_c_175_n N_A_27_367#_c_579_n 0.0224021f $X=1.765 $Y=0.7 $X2=0
+ $Y2=0
cc_232 N_A_73_269#_M1022_g N_A_27_367#_c_580_n 3.03248e-19 $X=0.5 $Y=0.655 $X2=0
+ $Y2=0
cc_233 N_A_73_269#_M1020_d N_A_27_367#_c_593_n 0.00248866f $X=1.535 $Y=2.325
+ $X2=0 $Y2=0
cc_234 N_A_73_269#_c_180_n N_A_27_367#_c_593_n 0.00532413f $X=1.51 $Y=2.365
+ $X2=0 $Y2=0
cc_235 N_A_73_269#_c_183_n N_A_27_367#_c_593_n 0.0199075f $X=1.675 $Y=2.365
+ $X2=0 $Y2=0
cc_236 N_A_73_269#_c_183_n N_A_27_367#_c_594_n 0.0201471f $X=1.675 $Y=2.365
+ $X2=0 $Y2=0
cc_237 N_A_73_269#_c_183_n N_A_27_367#_c_596_n 0.0134678f $X=1.675 $Y=2.365
+ $X2=0 $Y2=0
cc_238 N_A_73_269#_c_175_n N_A_27_367#_c_581_n 0.00492705f $X=1.765 $Y=0.7 $X2=0
+ $Y2=0
cc_239 N_A_73_269#_M1022_g N_A_27_367#_c_582_n 0.00471714f $X=0.5 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_73_269#_c_173_n N_A_27_367#_c_582_n 7.18885e-19 $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_241 N_A_73_269#_c_174_n N_A_27_367#_c_582_n 0.00233386f $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_242 N_A_73_269#_M1025_g N_A_27_367#_c_600_n 0.00437955f $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_243 N_A_73_269#_c_178_n N_A_27_367#_c_600_n 0.00939037f $X=1.12 $Y=2.28 $X2=0
+ $Y2=0
cc_244 N_A_73_269#_M1025_g N_A_27_367#_c_583_n 0.00508114f $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_245 N_A_73_269#_M1022_g N_A_27_367#_c_583_n 0.00499736f $X=0.5 $Y=0.655 $X2=0
+ $Y2=0
cc_246 N_A_73_269#_c_173_n N_A_27_367#_c_583_n 0.0282952f $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_247 N_A_73_269#_c_174_n N_A_27_367#_c_583_n 0.00803689f $X=0.53 $Y=1.51 $X2=0
+ $Y2=0
cc_248 N_A_73_269#_M1025_g N_A_27_367#_c_602_n 0.0075038f $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_249 N_A_73_269#_M1025_g N_A_27_367#_c_603_n 0.0128688f $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_250 N_A_73_269#_c_187_p N_A_27_367#_c_603_n 0.00456298f $X=1.205 $Y=2.365
+ $X2=0 $Y2=0
cc_251 N_A_73_269#_M1025_g N_A_27_367#_c_604_n 9.11509e-19 $X=0.475 $Y=2.465
+ $X2=0 $Y2=0
cc_252 N_A_73_269#_c_180_n N_A_27_367#_c_604_n 0.00391728f $X=1.51 $Y=2.365
+ $X2=0 $Y2=0
cc_253 N_A_73_269#_c_187_p N_A_27_367#_c_604_n 0.00461904f $X=1.205 $Y=2.365
+ $X2=0 $Y2=0
cc_254 N_A_73_269#_c_183_n N_A_27_367#_c_604_n 0.00624844f $X=1.675 $Y=2.365
+ $X2=0 $Y2=0
cc_255 N_A_73_269#_c_175_n N_A_27_367#_c_587_n 2.45633e-19 $X=1.765 $Y=0.7 $X2=0
+ $Y2=0
cc_256 N_A_73_269#_M1025_g N_VPWR_c_1026_n 0.00398394f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_A_73_269#_M1025_g N_VPWR_c_1031_n 0.00539556f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_258 N_A_73_269#_M1025_g N_VPWR_c_1017_n 0.00776348f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_259 N_A_73_269#_c_180_n A_235_465# 0.00130477f $X=1.51 $Y=2.365 $X2=-0.19
+ $Y2=-0.245
cc_260 N_A_73_269#_M1022_g N_VGND_c_1184_n 0.0129971f $X=0.5 $Y=0.655 $X2=0
+ $Y2=0
cc_261 N_A_73_269#_M1022_g N_VGND_c_1195_n 0.00486043f $X=0.5 $Y=0.655 $X2=0
+ $Y2=0
cc_262 N_A_73_269#_M1022_g N_VGND_c_1202_n 0.00545913f $X=0.5 $Y=0.655 $X2=0
+ $Y2=0
cc_263 N_GATE_M1006_g N_A_277_367#_c_340_n 2.46589e-19 $X=1.1 $Y=2.645 $X2=0
+ $Y2=0
cc_264 N_GATE_M1006_g N_A_277_367#_c_341_n 0.0780801f $X=1.1 $Y=2.645 $X2=0
+ $Y2=0
cc_265 N_GATE_M1006_g N_A_277_367#_c_333_n 9.06719e-19 $X=1.1 $Y=2.645 $X2=0
+ $Y2=0
cc_266 N_GATE_M1006_g N_A_295_55#_M1001_g 0.00735403f $X=1.1 $Y=2.645 $X2=0
+ $Y2=0
cc_267 N_GATE_M1009_g N_A_295_55#_M1001_g 0.0698816f $X=1.19 $Y=0.615 $X2=0
+ $Y2=0
cc_268 GATE N_A_295_55#_M1001_g 0.00118502f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_269 N_GATE_M1006_g N_A_27_367#_c_610_n 0.00795544f $X=1.1 $Y=2.645 $X2=0
+ $Y2=0
cc_270 N_GATE_M1009_g N_A_27_367#_c_578_n 0.00783094f $X=1.19 $Y=0.615 $X2=0
+ $Y2=0
cc_271 GATE N_A_27_367#_c_578_n 0.0286498f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_272 N_GATE_c_282_n N_A_27_367#_c_578_n 0.00465049f $X=1.1 $Y=1.295 $X2=0
+ $Y2=0
cc_273 N_GATE_M1009_g N_A_27_367#_c_618_n 0.0116422f $X=1.19 $Y=0.615 $X2=0
+ $Y2=0
cc_274 N_GATE_M1009_g N_A_27_367#_c_579_n 0.00391181f $X=1.19 $Y=0.615 $X2=0
+ $Y2=0
cc_275 N_GATE_M1009_g N_A_27_367#_c_580_n 0.00485951f $X=1.19 $Y=0.615 $X2=0
+ $Y2=0
cc_276 N_GATE_M1009_g N_A_27_367#_c_582_n 4.83753e-19 $X=1.19 $Y=0.615 $X2=0
+ $Y2=0
cc_277 N_GATE_M1006_g N_A_27_367#_c_600_n 0.00247507f $X=1.1 $Y=2.645 $X2=0
+ $Y2=0
cc_278 GATE N_A_27_367#_c_583_n 0.00592038f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_279 N_GATE_M1006_g N_A_27_367#_c_602_n 8.66486e-19 $X=1.1 $Y=2.645 $X2=0
+ $Y2=0
cc_280 N_GATE_M1006_g N_A_27_367#_c_604_n 0.009875f $X=1.1 $Y=2.645 $X2=0 $Y2=0
cc_281 N_GATE_M1006_g N_VPWR_c_1027_n 0.00303969f $X=1.1 $Y=2.645 $X2=0 $Y2=0
cc_282 N_GATE_M1006_g N_VPWR_c_1031_n 0.00148161f $X=1.1 $Y=2.645 $X2=0 $Y2=0
cc_283 N_GATE_M1006_g N_VPWR_c_1017_n 0.00384886f $X=1.1 $Y=2.645 $X2=0 $Y2=0
cc_284 N_GATE_M1009_g N_VGND_c_1184_n 0.00142593f $X=1.19 $Y=0.615 $X2=0 $Y2=0
cc_285 N_GATE_M1009_g N_VGND_c_1191_n 9.47364e-19 $X=1.19 $Y=0.615 $X2=0 $Y2=0
cc_286 N_A_277_367#_c_335_n N_A_295_55#_M1024_s 0.00534304f $X=4.7 $Y=0.71
+ $X2=-0.19 $Y2=-0.245
cc_287 N_A_277_367#_c_344_n N_A_295_55#_M1012_s 0.00923189f $X=4.7 $Y=2.25 $X2=0
+ $Y2=0
cc_288 N_A_277_367#_c_333_n N_A_295_55#_M1001_g 0.00173547f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_289 N_A_277_367#_c_334_n N_A_295_55#_M1001_g 0.0205745f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_290 N_A_277_367#_c_338_n N_A_295_55#_M1001_g 0.0151544f $X=2 $Y=0.935 $X2=0
+ $Y2=0
cc_291 N_A_277_367#_c_340_n N_A_295_55#_c_463_n 0.00409274f $X=1.835 $Y=2.005
+ $X2=0 $Y2=0
cc_292 N_A_277_367#_c_333_n N_A_295_55#_c_463_n 0.0061032f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_293 N_A_277_367#_c_334_n N_A_295_55#_c_463_n 0.0214155f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_294 N_A_277_367#_c_341_n N_A_295_55#_c_464_n 0.0152711f $X=1.55 $Y=2 $X2=0
+ $Y2=0
cc_295 N_A_277_367#_M1020_g N_A_295_55#_M1007_g 0.0140791f $X=1.46 $Y=2.645
+ $X2=0 $Y2=0
cc_296 N_A_277_367#_c_341_n N_A_295_55#_M1007_g 0.0214576f $X=1.55 $Y=2 $X2=0
+ $Y2=0
cc_297 N_A_277_367#_c_333_n N_A_295_55#_M1007_g 0.00352149f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_298 N_A_277_367#_c_346_n N_A_295_55#_M1007_g 0.0153905f $X=2 $Y=2.005 $X2=0
+ $Y2=0
cc_299 N_A_277_367#_c_343_n N_A_295_55#_M1021_g 0.0175757f $X=3.365 $Y=2.02
+ $X2=0 $Y2=0
cc_300 N_A_277_367#_c_347_n N_A_295_55#_M1021_g 0.0129603f $X=3.53 $Y=2.25 $X2=0
+ $Y2=0
cc_301 N_A_277_367#_c_333_n N_A_295_55#_c_468_n 0.008915f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_302 N_A_277_367#_c_343_n N_A_295_55#_c_469_n 0.00109587f $X=3.365 $Y=2.02
+ $X2=0 $Y2=0
cc_303 N_A_277_367#_c_333_n N_A_295_55#_c_470_n 0.0215724f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_304 N_A_277_367#_c_343_n N_A_295_55#_c_470_n 0.0693268f $X=3.365 $Y=2.02
+ $X2=0 $Y2=0
cc_305 N_A_277_367#_c_333_n N_A_295_55#_c_471_n 0.0114779f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_306 N_A_277_367#_c_343_n N_A_295_55#_c_471_n 0.0126257f $X=3.365 $Y=2.02
+ $X2=0 $Y2=0
cc_307 N_A_277_367#_c_337_n N_A_295_55#_c_472_n 0.00951179f $X=3.21 $Y=0.63
+ $X2=0 $Y2=0
cc_308 N_A_277_367#_c_335_n N_A_295_55#_c_473_n 0.0848087f $X=4.7 $Y=0.71 $X2=0
+ $Y2=0
cc_309 N_A_277_367#_c_336_n N_A_295_55#_c_473_n 0.0193359f $X=4.89 $Y=2.16 $X2=0
+ $Y2=0
cc_310 N_A_277_367#_c_337_n N_A_295_55#_c_473_n 0.0115259f $X=3.21 $Y=0.63 $X2=0
+ $Y2=0
cc_311 N_A_277_367#_c_344_n N_A_295_55#_c_474_n 0.0268479f $X=4.7 $Y=2.25 $X2=0
+ $Y2=0
cc_312 N_A_277_367#_c_336_n N_A_295_55#_c_474_n 0.0626286f $X=4.89 $Y=2.16 $X2=0
+ $Y2=0
cc_313 N_A_277_367#_c_347_n N_A_295_55#_c_474_n 0.00249179f $X=3.53 $Y=2.25
+ $X2=0 $Y2=0
cc_314 N_A_277_367#_c_337_n N_A_295_55#_c_475_n 0.00116001f $X=3.21 $Y=0.63
+ $X2=0 $Y2=0
cc_315 N_A_277_367#_c_343_n N_A_27_367#_M1011_g 0.00152701f $X=3.365 $Y=2.02
+ $X2=0 $Y2=0
cc_316 N_A_277_367#_c_335_n N_A_27_367#_c_576_n 5.20381e-19 $X=4.7 $Y=0.71 $X2=0
+ $Y2=0
cc_317 N_A_277_367#_c_336_n N_A_27_367#_c_576_n 0.00108963f $X=4.89 $Y=2.16
+ $X2=0 $Y2=0
cc_318 N_A_277_367#_c_333_n N_A_27_367#_c_579_n 0.00587057f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_319 N_A_277_367#_c_334_n N_A_27_367#_c_579_n 0.00177277f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_320 N_A_277_367#_c_338_n N_A_27_367#_c_579_n 0.0119541f $X=2 $Y=0.935 $X2=0
+ $Y2=0
cc_321 N_A_277_367#_M1020_g N_A_27_367#_c_593_n 0.0110858f $X=1.46 $Y=2.645
+ $X2=0 $Y2=0
cc_322 N_A_277_367#_M1020_g N_A_27_367#_c_594_n 0.00133769f $X=1.46 $Y=2.645
+ $X2=0 $Y2=0
cc_323 N_A_277_367#_c_343_n N_A_27_367#_c_595_n 0.070112f $X=3.365 $Y=2.02 $X2=0
+ $Y2=0
cc_324 N_A_277_367#_c_347_n N_A_27_367#_c_595_n 0.0142237f $X=3.53 $Y=2.25 $X2=0
+ $Y2=0
cc_325 N_A_277_367#_c_343_n N_A_27_367#_c_596_n 0.0020816f $X=3.365 $Y=2.02
+ $X2=0 $Y2=0
cc_326 N_A_277_367#_c_346_n N_A_27_367#_c_596_n 0.0130885f $X=2 $Y=2.005 $X2=0
+ $Y2=0
cc_327 N_A_277_367#_c_334_n N_A_27_367#_c_581_n 0.0016138f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_328 N_A_277_367#_c_338_n N_A_27_367#_c_581_n 0.00295333f $X=2 $Y=0.935 $X2=0
+ $Y2=0
cc_329 N_A_277_367#_c_347_n N_A_27_367#_c_672_n 0.00618661f $X=3.53 $Y=2.25
+ $X2=0 $Y2=0
cc_330 N_A_277_367#_c_344_n N_A_27_367#_c_598_n 0.0280546f $X=4.7 $Y=2.25 $X2=0
+ $Y2=0
cc_331 N_A_277_367#_M1020_g N_A_27_367#_c_604_n 0.00454354f $X=1.46 $Y=2.645
+ $X2=0 $Y2=0
cc_332 N_A_277_367#_c_333_n N_A_27_367#_c_584_n 0.0190208f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_333 N_A_277_367#_c_334_n N_A_27_367#_c_584_n 0.00141712f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_334 N_A_277_367#_c_333_n N_A_27_367#_c_585_n 2.92426e-19 $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_335 N_A_277_367#_c_334_n N_A_27_367#_c_585_n 0.0206819f $X=2 $Y=1.1 $X2=0
+ $Y2=0
cc_336 N_A_277_367#_c_344_n N_A_27_367#_c_605_n 0.00128606f $X=4.7 $Y=2.25 $X2=0
+ $Y2=0
cc_337 N_A_277_367#_c_343_n N_A_27_367#_c_606_n 0.00368364f $X=3.365 $Y=2.02
+ $X2=0 $Y2=0
cc_338 N_A_277_367#_c_344_n N_A_27_367#_c_606_n 0.00458552f $X=4.7 $Y=2.25 $X2=0
+ $Y2=0
cc_339 N_A_277_367#_c_347_n N_A_27_367#_c_606_n 0.0200558f $X=3.53 $Y=2.25 $X2=0
+ $Y2=0
cc_340 N_A_277_367#_c_344_n N_A_27_367#_c_607_n 0.0699027f $X=4.7 $Y=2.25 $X2=0
+ $Y2=0
cc_341 N_A_277_367#_c_347_n N_A_27_367#_c_607_n 0.00206778f $X=3.53 $Y=2.25
+ $X2=0 $Y2=0
cc_342 N_A_277_367#_c_338_n N_A_27_367#_c_587_n 0.0234317f $X=2 $Y=0.935 $X2=0
+ $Y2=0
cc_343 N_A_277_367#_c_344_n N_CLK_c_822_n 0.00121884f $X=4.7 $Y=2.25 $X2=-0.19
+ $Y2=-0.245
cc_344 N_A_277_367#_c_335_n N_CLK_M1024_g 0.0151873f $X=4.7 $Y=0.71 $X2=0 $Y2=0
cc_345 N_A_277_367#_c_336_n N_CLK_M1024_g 0.00920987f $X=4.89 $Y=2.16 $X2=0
+ $Y2=0
cc_346 N_A_277_367#_c_344_n N_CLK_M1012_g 0.0149077f $X=4.7 $Y=2.25 $X2=0 $Y2=0
cc_347 N_A_277_367#_c_336_n N_CLK_M1012_g 0.0186872f $X=4.89 $Y=2.16 $X2=0 $Y2=0
cc_348 N_A_277_367#_c_336_n N_CLK_c_824_n 0.00869799f $X=4.89 $Y=2.16 $X2=0
+ $Y2=0
cc_349 N_A_277_367#_c_344_n N_CLK_c_825_n 0.00205033f $X=4.7 $Y=2.25 $X2=0 $Y2=0
cc_350 N_A_277_367#_c_336_n N_CLK_c_825_n 0.00483548f $X=4.89 $Y=2.16 $X2=0
+ $Y2=0
cc_351 N_A_277_367#_c_335_n N_CLK_M1005_g 0.00802582f $X=4.7 $Y=0.71 $X2=0 $Y2=0
cc_352 N_A_277_367#_c_336_n N_CLK_M1005_g 0.0218995f $X=4.89 $Y=2.16 $X2=0 $Y2=0
cc_353 N_A_277_367#_c_344_n N_CLK_M1000_g 0.00153751f $X=4.7 $Y=2.25 $X2=0 $Y2=0
cc_354 N_A_277_367#_c_336_n N_CLK_M1000_g 0.00373484f $X=4.89 $Y=2.16 $X2=0
+ $Y2=0
cc_355 N_A_277_367#_c_336_n N_CLK_c_827_n 0.00575194f $X=4.89 $Y=2.16 $X2=0
+ $Y2=0
cc_356 N_A_277_367#_c_344_n N_CLK_c_828_n 0.0096866f $X=4.7 $Y=2.25 $X2=0 $Y2=0
cc_357 N_A_277_367#_c_347_n N_CLK_c_828_n 0.00113653f $X=3.53 $Y=2.25 $X2=0
+ $Y2=0
cc_358 N_A_277_367#_c_344_n N_CLK_c_829_n 0.00687881f $X=4.7 $Y=2.25 $X2=0 $Y2=0
cc_359 N_A_277_367#_c_347_n N_CLK_c_829_n 0.0260679f $X=3.53 $Y=2.25 $X2=0 $Y2=0
cc_360 N_A_277_367#_c_336_n N_A_1078_367#_c_902_n 0.0580703f $X=4.89 $Y=2.16
+ $X2=0 $Y2=0
cc_361 N_A_277_367#_c_335_n N_A_1078_367#_c_903_n 0.00701093f $X=4.7 $Y=0.71
+ $X2=0 $Y2=0
cc_362 N_A_277_367#_c_336_n N_A_1078_367#_c_903_n 0.0105706f $X=4.89 $Y=2.16
+ $X2=0 $Y2=0
cc_363 N_A_277_367#_c_336_n N_A_1078_367#_c_906_n 0.014458f $X=4.89 $Y=2.16
+ $X2=0 $Y2=0
cc_364 N_A_277_367#_c_344_n N_A_1078_367#_c_918_n 0.0149894f $X=4.7 $Y=2.25
+ $X2=0 $Y2=0
cc_365 N_A_277_367#_c_336_n N_A_1078_367#_c_918_n 0.0118213f $X=4.89 $Y=2.16
+ $X2=0 $Y2=0
cc_366 N_A_277_367#_c_343_n N_VPWR_M1011_d 0.00591796f $X=3.365 $Y=2.02 $X2=0
+ $Y2=0
cc_367 N_A_277_367#_c_344_n N_VPWR_M1012_d 0.00553698f $X=4.7 $Y=2.25 $X2=0
+ $Y2=0
cc_368 N_A_277_367#_c_336_n N_VPWR_M1012_d 0.00464539f $X=4.89 $Y=2.16 $X2=0
+ $Y2=0
cc_369 N_A_277_367#_M1020_g N_VPWR_c_1027_n 0.0028086f $X=1.46 $Y=2.645 $X2=0
+ $Y2=0
cc_370 N_A_277_367#_M1020_g N_VPWR_c_1017_n 0.0037128f $X=1.46 $Y=2.645 $X2=0
+ $Y2=0
cc_371 N_A_277_367#_c_335_n N_VGND_M1024_d 0.00487126f $X=4.7 $Y=0.71 $X2=0
+ $Y2=0
cc_372 N_A_277_367#_c_336_n N_VGND_M1024_d 0.00386648f $X=4.89 $Y=2.16 $X2=0
+ $Y2=0
cc_373 N_A_277_367#_c_335_n N_VGND_c_1186_n 0.0224106f $X=4.7 $Y=0.71 $X2=0
+ $Y2=0
cc_374 N_A_277_367#_c_338_n N_VGND_c_1191_n 9.29198e-19 $X=2 $Y=0.935 $X2=0
+ $Y2=0
cc_375 N_A_277_367#_c_335_n N_VGND_c_1193_n 0.0239195f $X=4.7 $Y=0.71 $X2=0
+ $Y2=0
cc_376 N_A_277_367#_c_337_n N_VGND_c_1193_n 0.0071156f $X=3.21 $Y=0.63 $X2=0
+ $Y2=0
cc_377 N_A_277_367#_c_335_n N_VGND_c_1196_n 0.00136551f $X=4.7 $Y=0.71 $X2=0
+ $Y2=0
cc_378 N_A_277_367#_c_335_n N_VGND_c_1202_n 0.0409344f $X=4.7 $Y=0.71 $X2=0
+ $Y2=0
cc_379 N_A_277_367#_c_337_n N_VGND_c_1202_n 0.00860093f $X=3.21 $Y=0.63 $X2=0
+ $Y2=0
cc_380 N_A_295_55#_M1007_g N_A_27_367#_M1011_g 0.0413462f $X=2 $Y=2.535 $X2=0
+ $Y2=0
cc_381 N_A_295_55#_M1021_g N_A_27_367#_M1011_g 0.00760229f $X=3.205 $Y=2.415
+ $X2=0 $Y2=0
cc_382 N_A_295_55#_c_471_n N_A_27_367#_M1011_g 0.00388244f $X=2.51 $Y=1.64 $X2=0
+ $Y2=0
cc_383 N_A_295_55#_M1021_g N_A_27_367#_c_590_n 0.00920339f $X=3.205 $Y=2.415
+ $X2=0 $Y2=0
cc_384 N_A_295_55#_M1001_g N_A_27_367#_c_578_n 4.93129e-19 $X=1.55 $Y=0.615
+ $X2=0 $Y2=0
cc_385 N_A_295_55#_M1001_g N_A_27_367#_c_618_n 0.00170147f $X=1.55 $Y=0.615
+ $X2=0 $Y2=0
cc_386 N_A_295_55#_M1001_g N_A_27_367#_c_579_n 0.00996442f $X=1.55 $Y=0.615
+ $X2=0 $Y2=0
cc_387 N_A_295_55#_M1007_g N_A_27_367#_c_593_n 0.00457473f $X=2 $Y=2.535 $X2=0
+ $Y2=0
cc_388 N_A_295_55#_M1007_g N_A_27_367#_c_594_n 0.00951605f $X=2 $Y=2.535 $X2=0
+ $Y2=0
cc_389 N_A_295_55#_M1021_g N_A_27_367#_c_595_n 0.00673163f $X=3.205 $Y=2.415
+ $X2=0 $Y2=0
cc_390 N_A_295_55#_M1007_g N_A_27_367#_c_596_n 0.00445753f $X=2 $Y=2.535 $X2=0
+ $Y2=0
cc_391 N_A_295_55#_c_471_n N_A_27_367#_c_596_n 4.22682e-19 $X=2.51 $Y=1.64 $X2=0
+ $Y2=0
cc_392 N_A_295_55#_M1008_g N_A_27_367#_c_581_n 9.47157e-19 $X=2.995 $Y=0.615
+ $X2=0 $Y2=0
cc_393 N_A_295_55#_c_472_n N_A_27_367#_c_581_n 0.00186536f $X=3.075 $Y=1.195
+ $X2=0 $Y2=0
cc_394 N_A_295_55#_M1021_g N_A_27_367#_c_672_n 0.0106359f $X=3.205 $Y=2.415
+ $X2=0 $Y2=0
cc_395 N_A_295_55#_M1021_g N_A_27_367#_c_597_n 0.00249323f $X=3.205 $Y=2.415
+ $X2=0 $Y2=0
cc_396 N_A_295_55#_c_466_n N_A_27_367#_c_584_n 2.4706e-19 $X=3.1 $Y=1.465 $X2=0
+ $Y2=0
cc_397 N_A_295_55#_c_470_n N_A_27_367#_c_584_n 0.0223307f $X=2.92 $Y=1.617 $X2=0
+ $Y2=0
cc_398 N_A_295_55#_c_471_n N_A_27_367#_c_584_n 0.00170816f $X=2.51 $Y=1.64 $X2=0
+ $Y2=0
cc_399 N_A_295_55#_c_472_n N_A_27_367#_c_584_n 0.0119192f $X=3.075 $Y=1.195
+ $X2=0 $Y2=0
cc_400 N_A_295_55#_c_543_p N_A_27_367#_c_584_n 0.00428673f $X=3.075 $Y=1.475
+ $X2=0 $Y2=0
cc_401 N_A_295_55#_c_475_n N_A_27_367#_c_584_n 2.2593e-19 $X=3.085 $Y=1.14 $X2=0
+ $Y2=0
cc_402 N_A_295_55#_M1008_g N_A_27_367#_c_585_n 0.0205909f $X=2.995 $Y=0.615
+ $X2=0 $Y2=0
cc_403 N_A_295_55#_c_470_n N_A_27_367#_c_585_n 0.00179318f $X=2.92 $Y=1.617
+ $X2=0 $Y2=0
cc_404 N_A_295_55#_c_471_n N_A_27_367#_c_585_n 0.0188545f $X=2.51 $Y=1.64 $X2=0
+ $Y2=0
cc_405 N_A_295_55#_c_472_n N_A_27_367#_c_585_n 4.29341e-19 $X=3.075 $Y=1.195
+ $X2=0 $Y2=0
cc_406 N_A_295_55#_M1021_g N_A_27_367#_c_605_n 0.00153497f $X=3.205 $Y=2.415
+ $X2=0 $Y2=0
cc_407 N_A_295_55#_M1021_g N_A_27_367#_c_606_n 0.00569306f $X=3.205 $Y=2.415
+ $X2=0 $Y2=0
cc_408 N_A_295_55#_M1021_g N_A_27_367#_c_607_n 0.00387387f $X=3.205 $Y=2.415
+ $X2=0 $Y2=0
cc_409 N_A_295_55#_M1008_g N_A_27_367#_c_587_n 0.0118852f $X=2.995 $Y=0.615
+ $X2=0 $Y2=0
cc_410 N_A_295_55#_c_473_n N_CLK_c_822_n 0.0102272f $X=4.2 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_411 N_A_295_55#_c_474_n N_CLK_c_822_n 0.0164913f $X=4.365 $Y=1.895 $X2=-0.19
+ $Y2=-0.245
cc_412 N_A_295_55#_c_473_n N_CLK_M1024_g 0.0103834f $X=4.2 $Y=1.08 $X2=0 $Y2=0
cc_413 N_A_295_55#_c_474_n N_CLK_M1024_g 0.0110429f $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_414 N_A_295_55#_c_474_n N_CLK_M1012_g 0.00630655f $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_415 N_A_295_55#_c_474_n N_CLK_c_825_n 0.00532568f $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_416 N_A_295_55#_c_474_n N_CLK_M1005_g 2.79513e-19 $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_417 N_A_295_55#_c_466_n N_CLK_c_828_n 0.0171945f $X=3.1 $Y=1.465 $X2=0 $Y2=0
cc_418 N_A_295_55#_c_470_n N_CLK_c_828_n 2.02477e-19 $X=2.92 $Y=1.617 $X2=0
+ $Y2=0
cc_419 N_A_295_55#_c_473_n N_CLK_c_828_n 0.00237107f $X=4.2 $Y=1.08 $X2=0 $Y2=0
cc_420 N_A_295_55#_c_474_n N_CLK_c_828_n 0.00160326f $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_421 N_A_295_55#_c_466_n N_CLK_c_829_n 0.00360511f $X=3.1 $Y=1.465 $X2=0 $Y2=0
cc_422 N_A_295_55#_c_470_n N_CLK_c_829_n 0.0244437f $X=2.92 $Y=1.617 $X2=0 $Y2=0
cc_423 N_A_295_55#_c_543_p N_CLK_c_829_n 0.00881075f $X=3.075 $Y=1.475 $X2=0
+ $Y2=0
cc_424 N_A_295_55#_c_473_n N_CLK_c_829_n 0.0356038f $X=4.2 $Y=1.08 $X2=0 $Y2=0
cc_425 N_A_295_55#_c_474_n N_CLK_c_829_n 0.0183376f $X=4.365 $Y=1.895 $X2=0
+ $Y2=0
cc_426 N_A_295_55#_M1021_g N_VPWR_c_1018_n 8.65752e-19 $X=3.205 $Y=2.415 $X2=0
+ $Y2=0
cc_427 N_A_295_55#_M1007_g N_VPWR_c_1027_n 3.27402e-19 $X=2 $Y=2.535 $X2=0 $Y2=0
cc_428 N_A_295_55#_M1008_g N_VGND_c_1185_n 0.0139287f $X=2.995 $Y=0.615 $X2=0
+ $Y2=0
cc_429 N_A_295_55#_c_472_n N_VGND_c_1185_n 0.00185745f $X=3.075 $Y=1.195 $X2=0
+ $Y2=0
cc_430 N_A_295_55#_M1001_g N_VGND_c_1191_n 9.29198e-19 $X=1.55 $Y=0.615 $X2=0
+ $Y2=0
cc_431 N_A_295_55#_M1008_g N_VGND_c_1193_n 0.0045897f $X=2.995 $Y=0.615 $X2=0
+ $Y2=0
cc_432 N_A_295_55#_M1008_g N_VGND_c_1202_n 0.0044912f $X=2.995 $Y=0.615 $X2=0
+ $Y2=0
cc_433 N_A_27_367#_c_598_n N_CLK_M1012_g 0.00960813f $X=5.795 $Y=2.595 $X2=0
+ $Y2=0
cc_434 N_A_27_367#_c_576_n N_CLK_M1005_g 0.0724447f $X=5.415 $Y=1.185 $X2=0
+ $Y2=0
cc_435 N_A_27_367#_c_588_n N_CLK_M1005_g 0.00385913f $X=5.745 $Y=1.425 $X2=0
+ $Y2=0
cc_436 N_A_27_367#_c_598_n N_CLK_M1000_g 0.0135905f $X=5.795 $Y=2.595 $X2=0
+ $Y2=0
cc_437 N_A_27_367#_c_599_n N_CLK_M1000_g 7.71267e-19 $X=5.885 $Y=2.51 $X2=0
+ $Y2=0
cc_438 N_A_27_367#_c_607_n N_CLK_M1000_g 0.00450842f $X=4.54 $Y=2.792 $X2=0
+ $Y2=0
cc_439 N_A_27_367#_M1017_g N_CLK_c_827_n 0.0523997f $X=5.745 $Y=2.465 $X2=0
+ $Y2=0
cc_440 N_A_27_367#_c_599_n N_CLK_c_827_n 3.45306e-19 $X=5.885 $Y=2.51 $X2=0
+ $Y2=0
cc_441 N_A_27_367#_c_588_n N_CLK_c_827_n 0.0110929f $X=5.745 $Y=1.425 $X2=0
+ $Y2=0
cc_442 N_A_27_367#_c_598_n N_A_1078_367#_M1000_d 0.00470942f $X=5.795 $Y=2.595
+ $X2=0 $Y2=0
cc_443 N_A_27_367#_M1017_g N_A_1078_367#_M1003_g 0.0425874f $X=5.745 $Y=2.465
+ $X2=0 $Y2=0
cc_444 N_A_27_367#_c_598_n N_A_1078_367#_M1003_g 0.00157399f $X=5.795 $Y=2.595
+ $X2=0 $Y2=0
cc_445 N_A_27_367#_c_599_n N_A_1078_367#_M1003_g 0.00860656f $X=5.885 $Y=2.51
+ $X2=0 $Y2=0
cc_446 N_A_27_367#_c_588_n N_A_1078_367#_M1004_g 0.00480498f $X=5.745 $Y=1.425
+ $X2=0 $Y2=0
cc_447 N_A_27_367#_M1017_g N_A_1078_367#_c_902_n 0.00154611f $X=5.745 $Y=2.465
+ $X2=0 $Y2=0
cc_448 N_A_27_367#_c_599_n N_A_1078_367#_c_902_n 0.00990203f $X=5.885 $Y=2.51
+ $X2=0 $Y2=0
cc_449 N_A_27_367#_c_586_n N_A_1078_367#_c_902_n 0.0188423f $X=5.885 $Y=1.535
+ $X2=0 $Y2=0
cc_450 N_A_27_367#_c_588_n N_A_1078_367#_c_902_n 0.0089442f $X=5.745 $Y=1.425
+ $X2=0 $Y2=0
cc_451 N_A_27_367#_c_576_n N_A_1078_367#_c_903_n 0.0151367f $X=5.415 $Y=1.185
+ $X2=0 $Y2=0
cc_452 N_A_27_367#_c_586_n N_A_1078_367#_c_904_n 0.0129265f $X=5.885 $Y=1.535
+ $X2=0 $Y2=0
cc_453 N_A_27_367#_c_588_n N_A_1078_367#_c_904_n 0.00539944f $X=5.745 $Y=1.425
+ $X2=0 $Y2=0
cc_454 N_A_27_367#_c_586_n N_A_1078_367#_c_905_n 0.0151309f $X=5.885 $Y=1.535
+ $X2=0 $Y2=0
cc_455 N_A_27_367#_c_588_n N_A_1078_367#_c_905_n 0.00286363f $X=5.745 $Y=1.425
+ $X2=0 $Y2=0
cc_456 N_A_27_367#_c_576_n N_A_1078_367#_c_906_n 0.0109108f $X=5.415 $Y=1.185
+ $X2=0 $Y2=0
cc_457 N_A_27_367#_c_586_n N_A_1078_367#_c_906_n 0.0153021f $X=5.885 $Y=1.535
+ $X2=0 $Y2=0
cc_458 N_A_27_367#_c_588_n N_A_1078_367#_c_906_n 0.0204094f $X=5.745 $Y=1.425
+ $X2=0 $Y2=0
cc_459 N_A_27_367#_c_598_n N_A_1078_367#_c_918_n 0.0226087f $X=5.795 $Y=2.595
+ $X2=0 $Y2=0
cc_460 N_A_27_367#_c_586_n N_A_1078_367#_c_918_n 8.22615e-19 $X=5.885 $Y=1.535
+ $X2=0 $Y2=0
cc_461 N_A_27_367#_c_588_n N_A_1078_367#_c_918_n 0.00447339f $X=5.745 $Y=1.425
+ $X2=0 $Y2=0
cc_462 N_A_27_367#_c_586_n N_A_1078_367#_c_907_n 0.00308875f $X=5.885 $Y=1.535
+ $X2=0 $Y2=0
cc_463 N_A_27_367#_c_588_n N_A_1078_367#_c_907_n 0.022298f $X=5.745 $Y=1.425
+ $X2=0 $Y2=0
cc_464 N_A_27_367#_c_610_n N_VPWR_M1025_d 0.0186075f $X=1.115 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_465 N_A_27_367#_c_595_n N_VPWR_M1011_d 0.0158736f $X=3.025 $Y=2.365 $X2=0
+ $Y2=0
cc_466 N_A_27_367#_c_672_n N_VPWR_M1011_d 0.00420986f $X=3.11 $Y=2.765 $X2=0
+ $Y2=0
cc_467 N_A_27_367#_c_597_n N_VPWR_M1011_d 0.00156804f $X=3.195 $Y=2.92 $X2=0
+ $Y2=0
cc_468 N_A_27_367#_c_598_n N_VPWR_M1012_d 0.0102596f $X=5.795 $Y=2.595 $X2=0
+ $Y2=0
cc_469 N_A_27_367#_c_598_n N_VPWR_M1017_d 0.00295499f $X=5.795 $Y=2.595 $X2=0
+ $Y2=0
cc_470 N_A_27_367#_c_599_n N_VPWR_M1017_d 0.00729317f $X=5.885 $Y=2.51 $X2=0
+ $Y2=0
cc_471 N_A_27_367#_M1011_g N_VPWR_c_1018_n 0.00837549f $X=2.36 $Y=2.535 $X2=0
+ $Y2=0
cc_472 N_A_27_367#_c_590_n N_VPWR_c_1018_n 0.0250323f $X=3.815 $Y=3.15 $X2=0
+ $Y2=0
cc_473 N_A_27_367#_c_593_n N_VPWR_c_1018_n 0.00935401f $X=2.02 $Y=2.99 $X2=0
+ $Y2=0
cc_474 N_A_27_367#_c_594_n N_VPWR_c_1018_n 0.0136805f $X=2.105 $Y=2.905 $X2=0
+ $Y2=0
cc_475 N_A_27_367#_c_595_n N_VPWR_c_1018_n 0.0266856f $X=3.025 $Y=2.365 $X2=0
+ $Y2=0
cc_476 N_A_27_367#_c_672_n N_VPWR_c_1018_n 0.0110448f $X=3.11 $Y=2.765 $X2=0
+ $Y2=0
cc_477 N_A_27_367#_c_597_n N_VPWR_c_1018_n 0.0269118f $X=3.195 $Y=2.92 $X2=0
+ $Y2=0
cc_478 N_A_27_367#_c_598_n N_VPWR_c_1019_n 0.0252356f $X=5.795 $Y=2.595 $X2=0
+ $Y2=0
cc_479 N_A_27_367#_c_605_n N_VPWR_c_1019_n 0.00276509f $X=3.98 $Y=2.94 $X2=0
+ $Y2=0
cc_480 N_A_27_367#_c_607_n N_VPWR_c_1019_n 0.01334f $X=4.54 $Y=2.792 $X2=0 $Y2=0
cc_481 N_A_27_367#_M1017_g N_VPWR_c_1020_n 0.00870662f $X=5.745 $Y=2.465 $X2=0
+ $Y2=0
cc_482 N_A_27_367#_c_598_n N_VPWR_c_1020_n 0.0101142f $X=5.795 $Y=2.595 $X2=0
+ $Y2=0
cc_483 N_A_27_367#_c_610_n N_VPWR_c_1026_n 0.00314202f $X=1.115 $Y=2.715 $X2=0
+ $Y2=0
cc_484 N_A_27_367#_c_602_n N_VPWR_c_1026_n 0.02171f $X=0.265 $Y=2.715 $X2=0
+ $Y2=0
cc_485 N_A_27_367#_c_591_n N_VPWR_c_1027_n 0.00932713f $X=2.435 $Y=3.15 $X2=0
+ $Y2=0
cc_486 N_A_27_367#_c_610_n N_VPWR_c_1027_n 0.00338574f $X=1.115 $Y=2.715 $X2=0
+ $Y2=0
cc_487 N_A_27_367#_c_593_n N_VPWR_c_1027_n 0.0590684f $X=2.02 $Y=2.99 $X2=0
+ $Y2=0
cc_488 N_A_27_367#_c_604_n N_VPWR_c_1027_n 0.0114718f $X=1.2 $Y=2.715 $X2=0
+ $Y2=0
cc_489 N_A_27_367#_c_590_n N_VPWR_c_1028_n 0.0296784f $X=3.815 $Y=3.15 $X2=0
+ $Y2=0
cc_490 N_A_27_367#_c_597_n N_VPWR_c_1028_n 0.0115893f $X=3.195 $Y=2.92 $X2=0
+ $Y2=0
cc_491 N_A_27_367#_c_598_n N_VPWR_c_1028_n 0.00528231f $X=5.795 $Y=2.595 $X2=0
+ $Y2=0
cc_492 N_A_27_367#_c_606_n N_VPWR_c_1028_n 0.0914052f $X=3.805 $Y=2.792 $X2=0
+ $Y2=0
cc_493 N_A_27_367#_M1017_g N_VPWR_c_1029_n 0.00355356f $X=5.745 $Y=2.465 $X2=0
+ $Y2=0
cc_494 N_A_27_367#_c_598_n N_VPWR_c_1029_n 0.00894688f $X=5.795 $Y=2.595 $X2=0
+ $Y2=0
cc_495 N_A_27_367#_c_610_n N_VPWR_c_1031_n 0.0240513f $X=1.115 $Y=2.715 $X2=0
+ $Y2=0
cc_496 N_A_27_367#_c_604_n N_VPWR_c_1031_n 0.00759507f $X=1.2 $Y=2.715 $X2=0
+ $Y2=0
cc_497 N_A_27_367#_M1025_s N_VPWR_c_1017_n 0.00215158f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_498 N_A_27_367#_c_590_n N_VPWR_c_1017_n 0.0328122f $X=3.815 $Y=3.15 $X2=0
+ $Y2=0
cc_499 N_A_27_367#_c_591_n N_VPWR_c_1017_n 0.0115794f $X=2.435 $Y=3.15 $X2=0
+ $Y2=0
cc_500 N_A_27_367#_M1017_g N_VPWR_c_1017_n 0.00423632f $X=5.745 $Y=2.465 $X2=0
+ $Y2=0
cc_501 N_A_27_367#_c_610_n N_VPWR_c_1017_n 0.011672f $X=1.115 $Y=2.715 $X2=0
+ $Y2=0
cc_502 N_A_27_367#_c_593_n N_VPWR_c_1017_n 0.033557f $X=2.02 $Y=2.99 $X2=0 $Y2=0
cc_503 N_A_27_367#_c_597_n N_VPWR_c_1017_n 0.00583135f $X=3.195 $Y=2.92 $X2=0
+ $Y2=0
cc_504 N_A_27_367#_c_598_n N_VPWR_c_1017_n 0.0271222f $X=5.795 $Y=2.595 $X2=0
+ $Y2=0
cc_505 N_A_27_367#_c_602_n N_VPWR_c_1017_n 0.0129082f $X=0.265 $Y=2.715 $X2=0
+ $Y2=0
cc_506 N_A_27_367#_c_604_n N_VPWR_c_1017_n 0.00619154f $X=1.2 $Y=2.715 $X2=0
+ $Y2=0
cc_507 N_A_27_367#_c_605_n N_VPWR_c_1017_n 0.0101219f $X=3.98 $Y=2.94 $X2=0
+ $Y2=0
cc_508 N_A_27_367#_c_606_n N_VPWR_c_1017_n 0.0476445f $X=3.805 $Y=2.792 $X2=0
+ $Y2=0
cc_509 N_A_27_367#_c_593_n A_235_465# 8.78902e-19 $X=2.02 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_510 N_A_27_367#_c_604_n A_235_465# 0.00359192f $X=1.2 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_511 N_A_27_367#_c_594_n A_415_465# 0.00323238f $X=2.105 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_512 N_A_27_367#_c_595_n A_415_465# 0.00141176f $X=3.025 $Y=2.365 $X2=-0.19
+ $Y2=-0.245
cc_513 N_A_27_367#_c_599_n N_GCLK_c_1134_n 0.00451666f $X=5.885 $Y=2.51 $X2=0
+ $Y2=0
cc_514 N_A_27_367#_c_578_n N_VGND_M1022_d 0.00649064f $X=1.06 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_515 N_A_27_367#_c_578_n N_VGND_c_1184_n 0.0222397f $X=1.06 $Y=0.915 $X2=0
+ $Y2=0
cc_516 N_A_27_367#_c_580_n N_VGND_c_1184_n 0.0135766f $X=1.23 $Y=0.35 $X2=0
+ $Y2=0
cc_517 N_A_27_367#_c_579_n N_VGND_c_1185_n 0.0140159f $X=2.345 $Y=0.35 $X2=0
+ $Y2=0
cc_518 N_A_27_367#_c_581_n N_VGND_c_1185_n 0.02501f $X=2.43 $Y=1.015 $X2=0 $Y2=0
cc_519 N_A_27_367#_c_584_n N_VGND_c_1185_n 0.00119981f $X=2.54 $Y=1.1 $X2=0
+ $Y2=0
cc_520 N_A_27_367#_c_585_n N_VGND_c_1185_n 4.71302e-19 $X=2.54 $Y=1.1 $X2=0
+ $Y2=0
cc_521 N_A_27_367#_c_587_n N_VGND_c_1185_n 0.00356708f $X=2.54 $Y=0.935 $X2=0
+ $Y2=0
cc_522 N_A_27_367#_c_576_n N_VGND_c_1186_n 0.0017762f $X=5.415 $Y=1.185 $X2=0
+ $Y2=0
cc_523 N_A_27_367#_c_576_n N_VGND_c_1187_n 0.00357683f $X=5.415 $Y=1.185 $X2=0
+ $Y2=0
cc_524 N_A_27_367#_c_579_n N_VGND_c_1191_n 0.0790151f $X=2.345 $Y=0.35 $X2=0
+ $Y2=0
cc_525 N_A_27_367#_c_580_n N_VGND_c_1191_n 0.0114622f $X=1.23 $Y=0.35 $X2=0
+ $Y2=0
cc_526 N_A_27_367#_c_587_n N_VGND_c_1191_n 0.00123424f $X=2.54 $Y=0.935 $X2=0
+ $Y2=0
cc_527 N_A_27_367#_c_577_n N_VGND_c_1195_n 0.0196033f $X=0.285 $Y=0.42 $X2=0
+ $Y2=0
cc_528 N_A_27_367#_c_576_n N_VGND_c_1196_n 0.0054895f $X=5.415 $Y=1.185 $X2=0
+ $Y2=0
cc_529 N_A_27_367#_M1022_s N_VGND_c_1202_n 0.00242815f $X=0.16 $Y=0.235 $X2=0
+ $Y2=0
cc_530 N_A_27_367#_c_576_n N_VGND_c_1202_n 0.0111524f $X=5.415 $Y=1.185 $X2=0
+ $Y2=0
cc_531 N_A_27_367#_c_577_n N_VGND_c_1202_n 0.0110024f $X=0.285 $Y=0.42 $X2=0
+ $Y2=0
cc_532 N_A_27_367#_c_578_n N_VGND_c_1202_n 0.00983314f $X=1.06 $Y=0.915 $X2=0
+ $Y2=0
cc_533 N_A_27_367#_c_579_n N_VGND_c_1202_n 0.0482406f $X=2.345 $Y=0.35 $X2=0
+ $Y2=0
cc_534 N_A_27_367#_c_580_n N_VGND_c_1202_n 0.00657784f $X=1.23 $Y=0.35 $X2=0
+ $Y2=0
cc_535 N_A_27_367#_c_582_n N_VGND_c_1202_n 0.00226556f $X=0.272 $Y=0.915 $X2=0
+ $Y2=0
cc_536 N_A_27_367#_c_587_n N_VGND_c_1202_n 3.56444e-19 $X=2.54 $Y=0.935 $X2=0
+ $Y2=0
cc_537 N_A_27_367#_c_579_n A_253_81# 0.00366293f $X=2.345 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_538 N_A_27_367#_c_579_n A_411_81# 0.00668369f $X=2.345 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_539 N_CLK_M1012_g N_A_1078_367#_c_902_n 2.61113e-19 $X=4.695 $Y=2.155 $X2=0
+ $Y2=0
cc_540 N_CLK_M1005_g N_A_1078_367#_c_902_n 0.00223487f $X=5.055 $Y=0.655 $X2=0
+ $Y2=0
cc_541 N_CLK_M1000_g N_A_1078_367#_c_902_n 0.00716145f $X=5.315 $Y=2.465 $X2=0
+ $Y2=0
cc_542 N_CLK_c_827_n N_A_1078_367#_c_902_n 0.00683095f $X=5.315 $Y=1.62 $X2=0
+ $Y2=0
cc_543 N_CLK_M1005_g N_A_1078_367#_c_903_n 0.00254104f $X=5.055 $Y=0.655 $X2=0
+ $Y2=0
cc_544 N_CLK_M1005_g N_A_1078_367#_c_906_n 0.00105747f $X=5.055 $Y=0.655 $X2=0
+ $Y2=0
cc_545 N_CLK_M1012_g N_A_1078_367#_c_918_n 2.73647e-19 $X=4.695 $Y=2.155 $X2=0
+ $Y2=0
cc_546 N_CLK_M1000_g N_A_1078_367#_c_918_n 0.00823358f $X=5.315 $Y=2.465 $X2=0
+ $Y2=0
cc_547 N_CLK_M1000_g N_VPWR_c_1019_n 0.00994467f $X=5.315 $Y=2.465 $X2=0 $Y2=0
cc_548 N_CLK_M1000_g N_VPWR_c_1020_n 0.00121197f $X=5.315 $Y=2.465 $X2=0 $Y2=0
cc_549 N_CLK_M1012_g N_VPWR_c_1028_n 5.01637e-19 $X=4.695 $Y=2.155 $X2=0 $Y2=0
cc_550 N_CLK_M1000_g N_VPWR_c_1029_n 0.00427295f $X=5.315 $Y=2.465 $X2=0 $Y2=0
cc_551 N_CLK_M1000_g N_VPWR_c_1017_n 0.00740863f $X=5.315 $Y=2.465 $X2=0 $Y2=0
cc_552 N_CLK_M1005_g N_VGND_c_1186_n 0.00974209f $X=5.055 $Y=0.655 $X2=0 $Y2=0
cc_553 N_CLK_M1024_g N_VGND_c_1193_n 0.00309082f $X=4.51 $Y=0.865 $X2=0 $Y2=0
cc_554 N_CLK_M1005_g N_VGND_c_1196_n 0.00406161f $X=5.055 $Y=0.655 $X2=0 $Y2=0
cc_555 N_CLK_M1024_g N_VGND_c_1202_n 0.0046122f $X=4.51 $Y=0.865 $X2=0 $Y2=0
cc_556 N_CLK_M1005_g N_VGND_c_1202_n 0.00566259f $X=5.055 $Y=0.655 $X2=0 $Y2=0
cc_557 N_A_1078_367#_M1003_g N_VPWR_c_1020_n 0.00166734f $X=6.215 $Y=2.465 $X2=0
+ $Y2=0
cc_558 N_A_1078_367#_M1003_g N_VPWR_c_1021_n 7.23592e-19 $X=6.215 $Y=2.465 $X2=0
+ $Y2=0
cc_559 N_A_1078_367#_M1016_g N_VPWR_c_1021_n 0.0136135f $X=6.645 $Y=2.465 $X2=0
+ $Y2=0
cc_560 N_A_1078_367#_M1018_g N_VPWR_c_1021_n 0.0147143f $X=7.075 $Y=2.465 $X2=0
+ $Y2=0
cc_561 N_A_1078_367#_M1023_g N_VPWR_c_1021_n 0.0014178f $X=7.505 $Y=2.465 $X2=0
+ $Y2=0
cc_562 N_A_1078_367#_M1023_g N_VPWR_c_1023_n 0.0302457f $X=7.505 $Y=2.465 $X2=0
+ $Y2=0
cc_563 N_A_1078_367#_c_907_n N_VPWR_c_1023_n 9.792e-19 $X=7.505 $Y=1.5 $X2=0
+ $Y2=0
cc_564 N_A_1078_367#_M1003_g N_VPWR_c_1024_n 0.00585385f $X=6.215 $Y=2.465 $X2=0
+ $Y2=0
cc_565 N_A_1078_367#_M1016_g N_VPWR_c_1024_n 0.00486043f $X=6.645 $Y=2.465 $X2=0
+ $Y2=0
cc_566 N_A_1078_367#_M1018_g N_VPWR_c_1030_n 0.00486043f $X=7.075 $Y=2.465 $X2=0
+ $Y2=0
cc_567 N_A_1078_367#_M1023_g N_VPWR_c_1030_n 0.00427501f $X=7.505 $Y=2.465 $X2=0
+ $Y2=0
cc_568 N_A_1078_367#_M1000_d N_VPWR_c_1017_n 0.00331682f $X=5.39 $Y=1.835 $X2=0
+ $Y2=0
cc_569 N_A_1078_367#_M1003_g N_VPWR_c_1017_n 0.0106551f $X=6.215 $Y=2.465 $X2=0
+ $Y2=0
cc_570 N_A_1078_367#_M1016_g N_VPWR_c_1017_n 0.00824727f $X=6.645 $Y=2.465 $X2=0
+ $Y2=0
cc_571 N_A_1078_367#_M1018_g N_VPWR_c_1017_n 0.00824727f $X=7.075 $Y=2.465 $X2=0
+ $Y2=0
cc_572 N_A_1078_367#_M1023_g N_VPWR_c_1017_n 0.00820182f $X=7.505 $Y=2.465 $X2=0
+ $Y2=0
cc_573 N_A_1078_367#_M1003_g N_GCLK_c_1134_n 2.36962e-19 $X=6.215 $Y=2.465 $X2=0
+ $Y2=0
cc_574 N_A_1078_367#_c_905_n N_GCLK_c_1134_n 0.00136166f $X=6.23 $Y=1.415 $X2=0
+ $Y2=0
cc_575 N_A_1078_367#_c_968_p N_GCLK_c_1134_n 0.0135016f $X=6.99 $Y=1.5 $X2=0
+ $Y2=0
cc_576 N_A_1078_367#_c_907_n N_GCLK_c_1134_n 0.00289076f $X=7.505 $Y=1.5 $X2=0
+ $Y2=0
cc_577 N_A_1078_367#_M1016_g N_GCLK_c_1135_n 0.0128211f $X=6.645 $Y=2.465 $X2=0
+ $Y2=0
cc_578 N_A_1078_367#_M1018_g N_GCLK_c_1135_n 0.0128097f $X=7.075 $Y=2.465 $X2=0
+ $Y2=0
cc_579 N_A_1078_367#_c_968_p N_GCLK_c_1135_n 0.0347798f $X=6.99 $Y=1.5 $X2=0
+ $Y2=0
cc_580 N_A_1078_367#_c_907_n N_GCLK_c_1135_n 0.00277043f $X=7.505 $Y=1.5 $X2=0
+ $Y2=0
cc_581 N_A_1078_367#_M1013_g N_GCLK_c_1130_n 0.0138436f $X=6.795 $Y=0.655 $X2=0
+ $Y2=0
cc_582 N_A_1078_367#_M1015_g N_GCLK_c_1130_n 0.0154528f $X=7.225 $Y=0.655 $X2=0
+ $Y2=0
cc_583 N_A_1078_367#_c_968_p N_GCLK_c_1130_n 0.0337166f $X=6.99 $Y=1.5 $X2=0
+ $Y2=0
cc_584 N_A_1078_367#_c_907_n N_GCLK_c_1130_n 0.00289453f $X=7.505 $Y=1.5 $X2=0
+ $Y2=0
cc_585 N_A_1078_367#_M1004_g N_GCLK_c_1131_n 0.00139496f $X=6.365 $Y=0.655 $X2=0
+ $Y2=0
cc_586 N_A_1078_367#_c_904_n N_GCLK_c_1131_n 0.0142158f $X=6.145 $Y=1.15 $X2=0
+ $Y2=0
cc_587 N_A_1078_367#_c_905_n N_GCLK_c_1131_n 7.72657e-19 $X=6.23 $Y=1.415 $X2=0
+ $Y2=0
cc_588 N_A_1078_367#_c_968_p N_GCLK_c_1131_n 0.0153308f $X=6.99 $Y=1.5 $X2=0
+ $Y2=0
cc_589 N_A_1078_367#_c_907_n N_GCLK_c_1131_n 0.00299787f $X=7.505 $Y=1.5 $X2=0
+ $Y2=0
cc_590 N_A_1078_367#_M1019_g GCLK 0.00498038f $X=7.655 $Y=0.655 $X2=0 $Y2=0
cc_591 N_A_1078_367#_M1023_g GCLK 0.00294385f $X=7.505 $Y=2.465 $X2=0 $Y2=0
cc_592 N_A_1078_367#_c_907_n GCLK 0.00338141f $X=7.505 $Y=1.5 $X2=0 $Y2=0
cc_593 N_A_1078_367#_M1018_g GCLK 0.00298602f $X=7.075 $Y=2.465 $X2=0 $Y2=0
cc_594 N_A_1078_367#_M1015_g GCLK 0.00214724f $X=7.225 $Y=0.655 $X2=0 $Y2=0
cc_595 N_A_1078_367#_M1023_g GCLK 0.00776117f $X=7.505 $Y=2.465 $X2=0 $Y2=0
cc_596 N_A_1078_367#_M1019_g GCLK 0.00217473f $X=7.655 $Y=0.655 $X2=0 $Y2=0
cc_597 N_A_1078_367#_c_968_p GCLK 0.0112725f $X=6.99 $Y=1.5 $X2=0 $Y2=0
cc_598 N_A_1078_367#_c_907_n GCLK 0.0303556f $X=7.505 $Y=1.5 $X2=0 $Y2=0
cc_599 N_A_1078_367#_M1023_g GCLK 0.019635f $X=7.505 $Y=2.465 $X2=0 $Y2=0
cc_600 N_A_1078_367#_c_904_n N_VGND_M1004_s 0.00223089f $X=6.145 $Y=1.15 $X2=0
+ $Y2=0
cc_601 N_A_1078_367#_c_903_n N_VGND_c_1186_n 0.00669147f $X=5.63 $Y=0.42 $X2=0
+ $Y2=0
cc_602 N_A_1078_367#_M1004_g N_VGND_c_1187_n 0.0126571f $X=6.365 $Y=0.655 $X2=0
+ $Y2=0
cc_603 N_A_1078_367#_M1013_g N_VGND_c_1187_n 6.30983e-19 $X=6.795 $Y=0.655 $X2=0
+ $Y2=0
cc_604 N_A_1078_367#_c_903_n N_VGND_c_1187_n 0.0492815f $X=5.63 $Y=0.42 $X2=0
+ $Y2=0
cc_605 N_A_1078_367#_c_904_n N_VGND_c_1187_n 0.0227487f $X=6.145 $Y=1.15 $X2=0
+ $Y2=0
cc_606 N_A_1078_367#_c_907_n N_VGND_c_1187_n 5.47574e-19 $X=7.505 $Y=1.5 $X2=0
+ $Y2=0
cc_607 N_A_1078_367#_M1004_g N_VGND_c_1188_n 6.33812e-19 $X=6.365 $Y=0.655 $X2=0
+ $Y2=0
cc_608 N_A_1078_367#_M1013_g N_VGND_c_1188_n 0.0114862f $X=6.795 $Y=0.655 $X2=0
+ $Y2=0
cc_609 N_A_1078_367#_M1015_g N_VGND_c_1188_n 0.0115088f $X=7.225 $Y=0.655 $X2=0
+ $Y2=0
cc_610 N_A_1078_367#_M1019_g N_VGND_c_1188_n 6.48031e-19 $X=7.655 $Y=0.655 $X2=0
+ $Y2=0
cc_611 N_A_1078_367#_M1019_g N_VGND_c_1190_n 0.00708988f $X=7.655 $Y=0.655 $X2=0
+ $Y2=0
cc_612 N_A_1078_367#_c_903_n N_VGND_c_1196_n 0.0210467f $X=5.63 $Y=0.42 $X2=0
+ $Y2=0
cc_613 N_A_1078_367#_M1004_g N_VGND_c_1197_n 0.00486043f $X=6.365 $Y=0.655 $X2=0
+ $Y2=0
cc_614 N_A_1078_367#_M1013_g N_VGND_c_1197_n 0.00486043f $X=6.795 $Y=0.655 $X2=0
+ $Y2=0
cc_615 N_A_1078_367#_M1015_g N_VGND_c_1198_n 0.00486043f $X=7.225 $Y=0.655 $X2=0
+ $Y2=0
cc_616 N_A_1078_367#_M1019_g N_VGND_c_1198_n 0.00585385f $X=7.655 $Y=0.655 $X2=0
+ $Y2=0
cc_617 N_A_1078_367#_M1002_d N_VGND_c_1202_n 0.00215158f $X=5.49 $Y=0.235 $X2=0
+ $Y2=0
cc_618 N_A_1078_367#_M1004_g N_VGND_c_1202_n 0.00824727f $X=6.365 $Y=0.655 $X2=0
+ $Y2=0
cc_619 N_A_1078_367#_M1013_g N_VGND_c_1202_n 0.00824727f $X=6.795 $Y=0.655 $X2=0
+ $Y2=0
cc_620 N_A_1078_367#_M1015_g N_VGND_c_1202_n 0.00824727f $X=7.225 $Y=0.655 $X2=0
+ $Y2=0
cc_621 N_A_1078_367#_M1019_g N_VGND_c_1202_n 0.0114822f $X=7.655 $Y=0.655 $X2=0
+ $Y2=0
cc_622 N_A_1078_367#_c_903_n N_VGND_c_1202_n 0.0125689f $X=5.63 $Y=0.42 $X2=0
+ $Y2=0
cc_623 N_A_1078_367#_c_906_n A_1026_47# 0.00157447f $X=5.522 $Y=1.15 $X2=-0.19
+ $Y2=-0.245
cc_624 N_VPWR_c_1017_n N_GCLK_M1003_s 0.00397496f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_625 N_VPWR_c_1017_n N_GCLK_M1018_s 0.00380103f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_626 N_VPWR_c_1024_n N_GCLK_c_1168_n 0.0138717f $X=6.695 $Y=3.33 $X2=0 $Y2=0
cc_627 N_VPWR_c_1017_n N_GCLK_c_1168_n 0.00886411f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_628 N_VPWR_M1016_d N_GCLK_c_1135_n 0.00180746f $X=6.72 $Y=1.835 $X2=0 $Y2=0
cc_629 N_VPWR_c_1021_n N_GCLK_c_1135_n 0.0163515f $X=6.86 $Y=2.27 $X2=0 $Y2=0
cc_630 N_VPWR_c_1023_n GCLK 0.013759f $X=7.79 $Y=1.98 $X2=0 $Y2=0
cc_631 N_VPWR_c_1023_n GCLK 0.0829857f $X=7.79 $Y=1.98 $X2=0 $Y2=0
cc_632 N_VPWR_c_1030_n GCLK 0.0211418f $X=7.705 $Y=3.33 $X2=0 $Y2=0
cc_633 N_VPWR_c_1017_n GCLK 0.0125916f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_634 N_GCLK_c_1130_n N_VGND_c_1188_n 0.0216087f $X=7.345 $Y=1.16 $X2=0 $Y2=0
cc_635 GCLK N_VGND_c_1190_n 0.00145953f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_636 N_GCLK_c_1178_p N_VGND_c_1197_n 0.0124525f $X=6.58 $Y=0.42 $X2=0 $Y2=0
cc_637 N_GCLK_c_1179_p N_VGND_c_1198_n 0.0124525f $X=7.44 $Y=0.42 $X2=0 $Y2=0
cc_638 N_GCLK_M1004_d N_VGND_c_1202_n 0.00536646f $X=6.44 $Y=0.235 $X2=0 $Y2=0
cc_639 N_GCLK_M1015_d N_VGND_c_1202_n 0.00536646f $X=7.3 $Y=0.235 $X2=0 $Y2=0
cc_640 N_GCLK_c_1178_p N_VGND_c_1202_n 0.00730901f $X=6.58 $Y=0.42 $X2=0 $Y2=0
cc_641 N_GCLK_c_1179_p N_VGND_c_1202_n 0.00730901f $X=7.44 $Y=0.42 $X2=0 $Y2=0
cc_642 N_VGND_c_1202_n A_1026_47# 0.00899413f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
