* File: sky130_fd_sc_lp__and4bb_lp.pxi.spice
* Created: Fri Aug 28 10:09:35 2020
* 
x_PM_SKY130_FD_SC_LP__AND4BB_LP%A_N N_A_N_c_109_n N_A_N_M1009_g N_A_N_M1012_g
+ N_A_N_c_111_n N_A_N_M1002_g A_N N_A_N_c_113_n
+ PM_SKY130_FD_SC_LP__AND4BB_LP%A_N
x_PM_SKY130_FD_SC_LP__AND4BB_LP%B_N N_B_N_M1010_g N_B_N_c_148_n N_B_N_c_149_n
+ N_B_N_M1011_g N_B_N_M1003_g B_N N_B_N_c_153_n
+ PM_SKY130_FD_SC_LP__AND4BB_LP%B_N
x_PM_SKY130_FD_SC_LP__AND4BB_LP%A_27_51# N_A_27_51#_M1009_s N_A_27_51#_M1012_s
+ N_A_27_51#_c_196_n N_A_27_51#_M1013_g N_A_27_51#_M1014_g N_A_27_51#_c_198_n
+ N_A_27_51#_c_199_n N_A_27_51#_c_200_n N_A_27_51#_c_201_n N_A_27_51#_c_208_n
+ N_A_27_51#_c_202_n N_A_27_51#_c_203_n N_A_27_51#_c_204_n N_A_27_51#_c_205_n
+ PM_SKY130_FD_SC_LP__AND4BB_LP%A_27_51#
x_PM_SKY130_FD_SC_LP__AND4BB_LP%A_291_409# N_A_291_409#_M1011_d
+ N_A_291_409#_M1003_s N_A_291_409#_M1005_g N_A_291_409#_M1006_g
+ N_A_291_409#_c_276_n N_A_291_409#_c_284_n N_A_291_409#_c_285_n
+ N_A_291_409#_c_277_n N_A_291_409#_c_286_n N_A_291_409#_c_287_n
+ N_A_291_409#_c_278_n N_A_291_409#_c_279_n N_A_291_409#_c_288_n
+ N_A_291_409#_c_318_n N_A_291_409#_c_280_n N_A_291_409#_c_281_n
+ PM_SKY130_FD_SC_LP__AND4BB_LP%A_291_409#
x_PM_SKY130_FD_SC_LP__AND4BB_LP%C N_C_M1007_g N_C_c_376_n N_C_M1004_g
+ N_C_c_377_n C C N_C_c_379_n PM_SKY130_FD_SC_LP__AND4BB_LP%C
x_PM_SKY130_FD_SC_LP__AND4BB_LP%D N_D_c_429_n N_D_M1008_g N_D_M1001_g
+ N_D_c_430_n N_D_c_431_n N_D_c_432_n N_D_c_433_n D D N_D_c_435_n
+ PM_SKY130_FD_SC_LP__AND4BB_LP%D
x_PM_SKY130_FD_SC_LP__AND4BB_LP%A_461_47# N_A_461_47#_M1014_s
+ N_A_461_47#_M1013_d N_A_461_47#_M1004_d N_A_461_47#_c_485_n
+ N_A_461_47#_M1016_g N_A_461_47#_M1015_g N_A_461_47#_c_487_n
+ N_A_461_47#_M1000_g N_A_461_47#_c_488_n N_A_461_47#_c_489_n
+ N_A_461_47#_c_490_n N_A_461_47#_c_515_n N_A_461_47#_c_491_n
+ N_A_461_47#_c_492_n N_A_461_47#_c_493_n N_A_461_47#_c_521_n
+ N_A_461_47#_c_500_n N_A_461_47#_c_501_n N_A_461_47#_c_502_n
+ N_A_461_47#_c_494_n N_A_461_47#_c_495_n N_A_461_47#_c_496_n
+ N_A_461_47#_c_504_n N_A_461_47#_c_544_n N_A_461_47#_c_497_n
+ N_A_461_47#_c_498_n PM_SKY130_FD_SC_LP__AND4BB_LP%A_461_47#
x_PM_SKY130_FD_SC_LP__AND4BB_LP%VPWR N_VPWR_M1012_d N_VPWR_M1003_d
+ N_VPWR_M1005_d N_VPWR_M1001_d N_VPWR_c_623_n N_VPWR_c_624_n N_VPWR_c_625_n
+ N_VPWR_c_626_n N_VPWR_c_627_n N_VPWR_c_628_n VPWR N_VPWR_c_629_n
+ N_VPWR_c_630_n N_VPWR_c_631_n N_VPWR_c_622_n N_VPWR_c_633_n N_VPWR_c_634_n
+ N_VPWR_c_635_n PM_SKY130_FD_SC_LP__AND4BB_LP%VPWR
x_PM_SKY130_FD_SC_LP__AND4BB_LP%X N_X_M1000_d N_X_M1015_d N_X_c_689_n X X X
+ N_X_c_690_n X PM_SKY130_FD_SC_LP__AND4BB_LP%X
x_PM_SKY130_FD_SC_LP__AND4BB_LP%VGND N_VGND_M1002_d N_VGND_M1008_d
+ N_VGND_c_714_n N_VGND_c_715_n VGND N_VGND_c_716_n N_VGND_c_717_n
+ N_VGND_c_718_n N_VGND_c_719_n N_VGND_c_720_n N_VGND_c_721_n
+ PM_SKY130_FD_SC_LP__AND4BB_LP%VGND
cc_1 VNB N_A_N_c_109_n 0.0194751f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.785
cc_2 VNB N_A_N_M1012_g 0.0204172f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.505
cc_3 VNB N_A_N_c_111_n 0.0154981f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.785
cc_4 VNB A_N 0.00702815f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.84
cc_5 VNB N_A_N_c_113_n 0.0765408f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.95
cc_6 VNB N_B_N_M1010_g 0.0307631f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.465
cc_7 VNB N_B_N_c_148_n 0.0116307f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.505
cc_8 VNB N_B_N_c_149_n 0.00856639f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.505
cc_9 VNB N_B_N_M1011_g 0.0399399f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.465
cc_10 VNB N_B_N_M1003_g 0.0181433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB B_N 0.00310011f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.95
cc_12 VNB N_B_N_c_153_n 0.0340804f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.12
cc_13 VNB N_A_27_51#_c_196_n 8.733e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_51#_M1014_g 0.0233685f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.95
cc_15 VNB N_A_27_51#_c_198_n 0.0110193f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.455
cc_16 VNB N_A_27_51#_c_199_n 0.0237245f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.12
cc_17 VNB N_A_27_51#_c_200_n 0.0256961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_51#_c_201_n 0.0558479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_51#_c_202_n 0.0175309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_51#_c_203_n 0.0017465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_51#_c_204_n 0.0179131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_51#_c_205_n 9.07016e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_291_409#_M1006_g 0.0401436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_291_409#_c_276_n 0.0193765f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.95
cc_25 VNB N_A_291_409#_c_277_n 0.00613482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_291_409#_c_278_n 0.0202749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_291_409#_c_279_n 0.0056059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_291_409#_c_280_n 0.0167483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_291_409#_c_281_n 0.00489168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_M1007_g 0.0328533f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.465
cc_31 VNB N_C_c_376_n 0.00193406f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.505
cc_32 VNB N_C_c_377_n 0.0217904f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.84
cc_33 VNB C 0.00551176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_C_c_379_n 0.0157831f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.95
cc_35 VNB N_D_c_429_n 0.0151828f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.785
cc_36 VNB N_D_c_430_n 0.0188943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_D_c_431_n 0.0144854f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.95
cc_38 VNB N_D_c_432_n 0.0239185f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.95
cc_39 VNB N_D_c_433_n 0.00219364f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.95
cc_40 VNB D 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.455
cc_41 VNB N_D_c_435_n 0.0167682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_461_47#_c_485_n 0.0149541f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.465
cc_43 VNB N_A_461_47#_M1015_g 0.00284729f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.95
cc_44 VNB N_A_461_47#_c_487_n 0.0168724f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.95
cc_45 VNB N_A_461_47#_c_488_n 0.0201418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_461_47#_c_489_n 0.0139578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_461_47#_c_490_n 0.00324064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_461_47#_c_491_n 0.00110171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_461_47#_c_492_n 0.0231166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_461_47#_c_493_n 0.00378385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_461_47#_c_494_n 0.00418802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_461_47#_c_495_n 0.00173165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_461_47#_c_496_n 2.70146e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_461_47#_c_497_n 0.0423078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_461_47#_c_498_n 0.00138065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VPWR_c_622_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_X_c_689_n 0.0243953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_X_c_690_n 0.0469837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_714_n 0.00100404f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.465
cc_60 VNB N_VGND_c_715_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_716_n 0.0270011f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.95
cc_62 VNB N_VGND_c_717_n 0.0682705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_718_n 0.0325773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_719_n 0.290508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_720_n 0.00461329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_721_n 0.00510817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VPB N_A_N_M1012_g 0.0537073f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.505
cc_68 VPB N_B_N_M1003_g 0.0493619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_27_51#_c_196_n 0.0110163f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_27_51#_M1013_g 0.0302046f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.465
cc_71 VPB N_A_27_51#_c_208_n 0.049552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_27_51#_c_202_n 0.0294937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_27_51#_c_205_n 0.00680262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_291_409#_M1005_g 0.0256392f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.465
cc_75 VPB N_A_291_409#_c_276_n 0.00452586f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.95
cc_76 VPB N_A_291_409#_c_284_n 0.0121925f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.455
cc_77 VPB N_A_291_409#_c_285_n 0.0157931f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.12
cc_78 VPB N_A_291_409#_c_286_n 0.0109485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_291_409#_c_287_n 0.00534976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_291_409#_c_288_n 0.00523124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_C_c_376_n 0.010958f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.505
cc_82 VPB N_C_M1004_g 0.0328034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB C 0.00204589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_D_M1001_g 0.0324055f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.785
cc_85 VPB N_D_c_433_n 0.0121263f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.95
cc_86 VPB D 7.56276e-19 $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.455
cc_87 VPB N_A_461_47#_M1015_g 0.0454945f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=0.95
cc_88 VPB N_A_461_47#_c_500_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_461_47#_c_501_n 0.00673628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_461_47#_c_502_n 0.00958881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_461_47#_c_496_n 0.00267143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_461_47#_c_504_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_623_n 0.0236575f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.95
cc_94 VPB N_VPWR_c_624_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_625_n 0.00417575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_626_n 0.00418937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_627_n 0.0219685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_628_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_629_n 0.0276965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_630_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_631_n 0.023544f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_622_n 0.0791326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_633_n 0.0251939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_634_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_635_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB X 0.0576042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_X_c_690_n 0.0128754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 N_A_N_c_111_n N_B_N_M1010_g 0.0144633f $X=0.855 $Y=0.785 $X2=0 $Y2=0
cc_109 A_N N_B_N_M1010_g 0.0138745f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_110 N_A_N_c_113_n N_B_N_M1010_g 0.0250083f $X=0.79 $Y=0.95 $X2=0 $Y2=0
cc_111 A_N N_B_N_c_149_n 0.00764542f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_112 A_N N_B_N_M1011_g 0.0015474f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_113 A_N B_N 0.0204582f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_114 N_A_N_c_113_n B_N 2.12773e-19 $X=0.79 $Y=0.95 $X2=0 $Y2=0
cc_115 A_N N_B_N_c_153_n 8.99517e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_116 N_A_N_c_113_n N_B_N_c_153_n 0.00244257f $X=0.79 $Y=0.95 $X2=0 $Y2=0
cc_117 N_A_N_c_109_n N_A_27_51#_c_201_n 0.0113092f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_118 N_A_N_M1012_g N_A_27_51#_c_201_n 0.0115416f $X=0.545 $Y=2.505 $X2=0 $Y2=0
cc_119 N_A_N_c_111_n N_A_27_51#_c_201_n 0.00182322f $X=0.855 $Y=0.785 $X2=0
+ $Y2=0
cc_120 A_N N_A_27_51#_c_201_n 0.0509798f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_121 N_A_N_c_113_n N_A_27_51#_c_201_n 0.0247054f $X=0.79 $Y=0.95 $X2=0 $Y2=0
cc_122 N_A_N_M1012_g N_A_27_51#_c_208_n 0.0307921f $X=0.545 $Y=2.505 $X2=0 $Y2=0
cc_123 N_A_N_M1012_g N_A_27_51#_c_202_n 0.0253819f $X=0.545 $Y=2.505 $X2=0 $Y2=0
cc_124 A_N N_A_27_51#_c_202_n 0.0539787f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_125 N_A_N_c_113_n N_A_27_51#_c_202_n 0.00744212f $X=0.79 $Y=0.95 $X2=0 $Y2=0
cc_126 N_A_N_M1012_g N_A_27_51#_c_205_n 0.00383478f $X=0.545 $Y=2.505 $X2=0
+ $Y2=0
cc_127 A_N N_A_291_409#_c_279_n 0.00658732f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_128 N_A_N_M1012_g N_VPWR_c_623_n 0.0258594f $X=0.545 $Y=2.505 $X2=0 $Y2=0
cc_129 N_A_N_M1012_g N_VPWR_c_622_n 0.0135501f $X=0.545 $Y=2.505 $X2=0 $Y2=0
cc_130 N_A_N_M1012_g N_VPWR_c_633_n 0.00717535f $X=0.545 $Y=2.505 $X2=0 $Y2=0
cc_131 N_A_N_c_109_n N_VGND_c_714_n 0.0020386f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_132 N_A_N_c_111_n N_VGND_c_714_n 0.0106393f $X=0.855 $Y=0.785 $X2=0 $Y2=0
cc_133 A_N N_VGND_c_714_n 0.0223243f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_134 N_A_N_c_109_n N_VGND_c_716_n 0.00530134f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_135 N_A_N_c_111_n N_VGND_c_716_n 0.00469214f $X=0.855 $Y=0.785 $X2=0 $Y2=0
cc_136 N_A_N_c_109_n N_VGND_c_719_n 0.0105687f $X=0.495 $Y=0.785 $X2=0 $Y2=0
cc_137 N_A_N_c_111_n N_VGND_c_719_n 0.00422139f $X=0.855 $Y=0.785 $X2=0 $Y2=0
cc_138 A_N N_VGND_c_719_n 0.0140272f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_139 N_A_N_c_113_n N_VGND_c_719_n 7.86289e-19 $X=0.79 $Y=0.95 $X2=0 $Y2=0
cc_140 N_B_N_M1003_g N_A_27_51#_c_196_n 0.0138901f $X=1.865 $Y=2.545 $X2=0 $Y2=0
cc_141 N_B_N_M1003_g N_A_27_51#_M1013_g 0.0314405f $X=1.865 $Y=2.545 $X2=0 $Y2=0
cc_142 B_N N_A_27_51#_c_199_n 4.71756e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_143 N_B_N_c_153_n N_A_27_51#_c_199_n 0.0138901f $X=1.725 $Y=1.29 $X2=0 $Y2=0
cc_144 N_B_N_M1011_g N_A_27_51#_c_200_n 0.0054956f $X=1.675 $Y=0.465 $X2=0 $Y2=0
cc_145 N_B_N_c_149_n N_A_27_51#_c_202_n 0.00838933f $X=1.36 $Y=1.2 $X2=0 $Y2=0
cc_146 N_B_N_M1003_g N_A_27_51#_c_202_n 0.0194538f $X=1.865 $Y=2.545 $X2=0 $Y2=0
cc_147 B_N N_A_27_51#_c_202_n 0.0231899f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_148 N_B_N_c_153_n N_A_27_51#_c_202_n 0.00471135f $X=1.725 $Y=1.29 $X2=0 $Y2=0
cc_149 B_N N_A_27_51#_c_203_n 0.013752f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_150 N_B_N_c_153_n N_A_27_51#_c_203_n 0.00204863f $X=1.725 $Y=1.29 $X2=0 $Y2=0
cc_151 B_N N_A_27_51#_c_204_n 6.94223e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_152 N_B_N_c_153_n N_A_27_51#_c_204_n 0.00586059f $X=1.725 $Y=1.29 $X2=0 $Y2=0
cc_153 N_B_N_M1003_g N_A_291_409#_c_285_n 0.0164265f $X=1.865 $Y=2.545 $X2=0
+ $Y2=0
cc_154 N_B_N_M1010_g N_A_291_409#_c_277_n 0.00180211f $X=1.285 $Y=0.465 $X2=0
+ $Y2=0
cc_155 N_B_N_M1011_g N_A_291_409#_c_277_n 0.011207f $X=1.675 $Y=0.465 $X2=0
+ $Y2=0
cc_156 N_B_N_M1003_g N_A_291_409#_c_286_n 0.0178604f $X=1.865 $Y=2.545 $X2=0
+ $Y2=0
cc_157 N_B_N_M1003_g N_A_291_409#_c_287_n 0.00195515f $X=1.865 $Y=2.545 $X2=0
+ $Y2=0
cc_158 N_B_N_M1010_g N_A_291_409#_c_279_n 4.83953e-19 $X=1.285 $Y=0.465 $X2=0
+ $Y2=0
cc_159 N_B_N_M1011_g N_A_291_409#_c_279_n 0.00662164f $X=1.675 $Y=0.465 $X2=0
+ $Y2=0
cc_160 B_N N_A_291_409#_c_279_n 0.0132149f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_161 N_B_N_c_153_n N_A_291_409#_c_279_n 0.00771406f $X=1.725 $Y=1.29 $X2=0
+ $Y2=0
cc_162 N_B_N_M1011_g N_A_461_47#_c_490_n 7.21241e-19 $X=1.675 $Y=0.465 $X2=0
+ $Y2=0
cc_163 N_B_N_M1003_g N_VPWR_c_624_n 0.0181825f $X=1.865 $Y=2.545 $X2=0 $Y2=0
cc_164 N_B_N_M1003_g N_VPWR_c_629_n 0.00769046f $X=1.865 $Y=2.545 $X2=0 $Y2=0
cc_165 N_B_N_M1003_g N_VPWR_c_622_n 0.0143431f $X=1.865 $Y=2.545 $X2=0 $Y2=0
cc_166 N_B_N_M1010_g N_VGND_c_714_n 0.0108718f $X=1.285 $Y=0.465 $X2=0 $Y2=0
cc_167 N_B_N_M1011_g N_VGND_c_714_n 0.00203639f $X=1.675 $Y=0.465 $X2=0 $Y2=0
cc_168 N_B_N_M1010_g N_VGND_c_717_n 0.00469214f $X=1.285 $Y=0.465 $X2=0 $Y2=0
cc_169 N_B_N_M1011_g N_VGND_c_717_n 0.00530134f $X=1.675 $Y=0.465 $X2=0 $Y2=0
cc_170 N_B_N_M1010_g N_VGND_c_719_n 0.00567722f $X=1.285 $Y=0.465 $X2=0 $Y2=0
cc_171 N_B_N_M1011_g N_VGND_c_719_n 0.010971f $X=1.675 $Y=0.465 $X2=0 $Y2=0
cc_172 N_A_27_51#_M1014_g N_A_291_409#_M1006_g 0.0471814f $X=2.665 $Y=0.445
+ $X2=0 $Y2=0
cc_173 N_A_27_51#_c_198_n N_A_291_409#_M1006_g 0.00481692f $X=2.395 $Y=1.135
+ $X2=0 $Y2=0
cc_174 N_A_27_51#_c_199_n N_A_291_409#_c_276_n 0.010283f $X=2.395 $Y=1.64 $X2=0
+ $Y2=0
cc_175 N_A_27_51#_c_202_n N_A_291_409#_c_276_n 3.08664e-19 $X=2.23 $Y=1.72 $X2=0
+ $Y2=0
cc_176 N_A_27_51#_c_196_n N_A_291_409#_c_284_n 0.010283f $X=2.395 $Y=1.805 $X2=0
+ $Y2=0
cc_177 N_A_27_51#_M1013_g N_A_291_409#_c_284_n 0.0305364f $X=2.395 $Y=2.545
+ $X2=0 $Y2=0
cc_178 N_A_27_51#_M1013_g N_A_291_409#_c_285_n 9.07377e-19 $X=2.395 $Y=2.545
+ $X2=0 $Y2=0
cc_179 N_A_27_51#_M1014_g N_A_291_409#_c_277_n 0.00421377f $X=2.665 $Y=0.445
+ $X2=0 $Y2=0
cc_180 N_A_27_51#_c_196_n N_A_291_409#_c_286_n 5.50032e-19 $X=2.395 $Y=1.805
+ $X2=0 $Y2=0
cc_181 N_A_27_51#_M1013_g N_A_291_409#_c_286_n 0.0209996f $X=2.395 $Y=2.545
+ $X2=0 $Y2=0
cc_182 N_A_27_51#_c_202_n N_A_291_409#_c_286_n 0.0561346f $X=2.23 $Y=1.72 $X2=0
+ $Y2=0
cc_183 N_A_27_51#_c_202_n N_A_291_409#_c_287_n 0.0265555f $X=2.23 $Y=1.72 $X2=0
+ $Y2=0
cc_184 N_A_27_51#_M1014_g N_A_291_409#_c_278_n 0.00433158f $X=2.665 $Y=0.445
+ $X2=0 $Y2=0
cc_185 N_A_27_51#_c_200_n N_A_291_409#_c_278_n 0.0185593f $X=2.665 $Y=0.9 $X2=0
+ $Y2=0
cc_186 N_A_27_51#_c_203_n N_A_291_409#_c_278_n 0.0234949f $X=2.395 $Y=1.3 $X2=0
+ $Y2=0
cc_187 N_A_27_51#_c_204_n N_A_291_409#_c_278_n 0.00121645f $X=2.395 $Y=1.3 $X2=0
+ $Y2=0
cc_188 N_A_27_51#_M1013_g N_A_291_409#_c_288_n 0.00119013f $X=2.395 $Y=2.545
+ $X2=0 $Y2=0
cc_189 N_A_27_51#_c_199_n N_A_291_409#_c_288_n 8.78698e-19 $X=2.395 $Y=1.64
+ $X2=0 $Y2=0
cc_190 N_A_27_51#_c_202_n N_A_291_409#_c_288_n 0.0102464f $X=2.23 $Y=1.72 $X2=0
+ $Y2=0
cc_191 N_A_27_51#_c_204_n N_A_291_409#_c_318_n 7.71269e-19 $X=2.395 $Y=1.3 $X2=0
+ $Y2=0
cc_192 N_A_27_51#_c_203_n N_A_291_409#_c_280_n 0.0015419f $X=2.395 $Y=1.3 $X2=0
+ $Y2=0
cc_193 N_A_27_51#_c_204_n N_A_291_409#_c_280_n 0.010283f $X=2.395 $Y=1.3 $X2=0
+ $Y2=0
cc_194 N_A_27_51#_c_198_n N_A_291_409#_c_281_n 0.00383847f $X=2.395 $Y=1.135
+ $X2=0 $Y2=0
cc_195 N_A_27_51#_c_200_n N_A_291_409#_c_281_n 6.97324e-19 $X=2.665 $Y=0.9 $X2=0
+ $Y2=0
cc_196 N_A_27_51#_c_203_n N_A_291_409#_c_281_n 0.0284581f $X=2.395 $Y=1.3 $X2=0
+ $Y2=0
cc_197 N_A_27_51#_M1014_g N_A_461_47#_c_490_n 0.0114538f $X=2.665 $Y=0.445 $X2=0
+ $Y2=0
cc_198 N_A_27_51#_c_200_n N_A_461_47#_c_490_n 0.00101421f $X=2.665 $Y=0.9 $X2=0
+ $Y2=0
cc_199 N_A_27_51#_M1013_g N_A_461_47#_c_504_n 0.0131865f $X=2.395 $Y=2.545 $X2=0
+ $Y2=0
cc_200 N_A_27_51#_c_208_n N_VPWR_c_623_n 0.0685263f $X=0.28 $Y=2.15 $X2=0 $Y2=0
cc_201 N_A_27_51#_c_202_n N_VPWR_c_623_n 0.0264016f $X=2.23 $Y=1.72 $X2=0 $Y2=0
cc_202 N_A_27_51#_M1013_g N_VPWR_c_624_n 0.0171369f $X=2.395 $Y=2.545 $X2=0
+ $Y2=0
cc_203 N_A_27_51#_M1013_g N_VPWR_c_625_n 7.73692e-19 $X=2.395 $Y=2.545 $X2=0
+ $Y2=0
cc_204 N_A_27_51#_M1013_g N_VPWR_c_630_n 0.00769046f $X=2.395 $Y=2.545 $X2=0
+ $Y2=0
cc_205 N_A_27_51#_M1013_g N_VPWR_c_622_n 0.0134474f $X=2.395 $Y=2.545 $X2=0
+ $Y2=0
cc_206 N_A_27_51#_c_208_n N_VPWR_c_622_n 0.0123184f $X=0.28 $Y=2.15 $X2=0 $Y2=0
cc_207 N_A_27_51#_c_208_n N_VPWR_c_633_n 0.0177662f $X=0.28 $Y=2.15 $X2=0 $Y2=0
cc_208 N_A_27_51#_c_201_n N_VGND_c_714_n 0.0113755f $X=0.28 $Y=0.48 $X2=0 $Y2=0
cc_209 N_A_27_51#_c_201_n N_VGND_c_716_n 0.0197885f $X=0.28 $Y=0.48 $X2=0 $Y2=0
cc_210 N_A_27_51#_M1014_g N_VGND_c_717_n 0.00359964f $X=2.665 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_A_27_51#_M1014_g N_VGND_c_719_n 0.00657133f $X=2.665 $Y=0.445 $X2=0
+ $Y2=0
cc_212 N_A_27_51#_c_201_n N_VGND_c_719_n 0.0125808f $X=0.28 $Y=0.48 $X2=0 $Y2=0
cc_213 N_A_291_409#_M1006_g N_C_M1007_g 0.0222252f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A_291_409#_c_284_n N_C_c_376_n 0.0222252f $X=2.965 $Y=1.885 $X2=0 $Y2=0
cc_215 N_A_291_409#_c_288_n N_C_c_376_n 2.5809e-19 $X=2.965 $Y=1.72 $X2=0 $Y2=0
cc_216 N_A_291_409#_M1005_g N_C_M1004_g 0.0369201f $X=2.925 $Y=2.545 $X2=0 $Y2=0
cc_217 N_A_291_409#_c_284_n N_C_M1004_g 0.00408524f $X=2.965 $Y=1.885 $X2=0
+ $Y2=0
cc_218 N_A_291_409#_c_288_n N_C_M1004_g 0.00177498f $X=2.965 $Y=1.72 $X2=0 $Y2=0
cc_219 N_A_291_409#_c_276_n N_C_c_377_n 0.0222252f $X=2.965 $Y=1.72 $X2=0 $Y2=0
cc_220 N_A_291_409#_c_288_n N_C_c_377_n 9.25891e-19 $X=2.965 $Y=1.72 $X2=0 $Y2=0
cc_221 N_A_291_409#_M1006_g C 0.00218582f $X=3.055 $Y=0.445 $X2=0 $Y2=0
cc_222 N_A_291_409#_c_288_n C 0.00401677f $X=2.965 $Y=1.72 $X2=0 $Y2=0
cc_223 N_A_291_409#_c_318_n C 0.0287541f $X=2.965 $Y=1.38 $X2=0 $Y2=0
cc_224 N_A_291_409#_c_281_n C 0.00374847f $X=2.965 $Y=1.215 $X2=0 $Y2=0
cc_225 N_A_291_409#_c_318_n N_C_c_379_n 9.25891e-19 $X=2.965 $Y=1.38 $X2=0 $Y2=0
cc_226 N_A_291_409#_c_280_n N_C_c_379_n 0.0222252f $X=2.965 $Y=1.38 $X2=0 $Y2=0
cc_227 N_A_291_409#_c_286_n N_A_461_47#_M1013_d 0.00180746f $X=2.8 $Y=2.07 $X2=0
+ $Y2=0
cc_228 N_A_291_409#_M1006_g N_A_461_47#_c_490_n 0.016933f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_229 N_A_291_409#_c_277_n N_A_461_47#_c_490_n 0.0234648f $X=1.89 $Y=0.48 $X2=0
+ $Y2=0
cc_230 N_A_291_409#_c_278_n N_A_461_47#_c_490_n 0.0435154f $X=2.8 $Y=0.86 $X2=0
+ $Y2=0
cc_231 N_A_291_409#_c_318_n N_A_461_47#_c_490_n 0.00419127f $X=2.965 $Y=1.38
+ $X2=0 $Y2=0
cc_232 N_A_291_409#_c_280_n N_A_461_47#_c_490_n 4.53216e-19 $X=2.965 $Y=1.38
+ $X2=0 $Y2=0
cc_233 N_A_291_409#_M1005_g N_A_461_47#_c_515_n 0.0147863f $X=2.925 $Y=2.545
+ $X2=0 $Y2=0
cc_234 N_A_291_409#_c_284_n N_A_461_47#_c_515_n 2.67759e-19 $X=2.965 $Y=1.885
+ $X2=0 $Y2=0
cc_235 N_A_291_409#_c_288_n N_A_461_47#_c_515_n 0.0152047f $X=2.965 $Y=1.72
+ $X2=0 $Y2=0
cc_236 N_A_291_409#_M1006_g N_A_461_47#_c_491_n 0.00346628f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_237 N_A_291_409#_M1006_g N_A_461_47#_c_493_n 0.00152461f $X=3.055 $Y=0.445
+ $X2=0 $Y2=0
cc_238 N_A_291_409#_c_278_n N_A_461_47#_c_493_n 0.00949973f $X=2.8 $Y=0.86 $X2=0
+ $Y2=0
cc_239 N_A_291_409#_M1005_g N_A_461_47#_c_521_n 8.00952e-19 $X=2.925 $Y=2.545
+ $X2=0 $Y2=0
cc_240 N_A_291_409#_c_288_n N_A_461_47#_c_521_n 3.6965e-19 $X=2.965 $Y=1.72
+ $X2=0 $Y2=0
cc_241 N_A_291_409#_M1005_g N_A_461_47#_c_500_n 8.64184e-19 $X=2.925 $Y=2.545
+ $X2=0 $Y2=0
cc_242 N_A_291_409#_M1005_g N_A_461_47#_c_502_n 4.85655e-19 $X=2.925 $Y=2.545
+ $X2=0 $Y2=0
cc_243 N_A_291_409#_c_288_n N_A_461_47#_c_502_n 0.00453365f $X=2.965 $Y=1.72
+ $X2=0 $Y2=0
cc_244 N_A_291_409#_M1005_g N_A_461_47#_c_504_n 0.0115522f $X=2.925 $Y=2.545
+ $X2=0 $Y2=0
cc_245 N_A_291_409#_c_286_n N_A_461_47#_c_504_n 0.0147186f $X=2.8 $Y=2.07 $X2=0
+ $Y2=0
cc_246 N_A_291_409#_c_288_n N_A_461_47#_c_504_n 0.00197994f $X=2.965 $Y=1.72
+ $X2=0 $Y2=0
cc_247 N_A_291_409#_c_286_n N_VPWR_M1003_d 0.00180746f $X=2.8 $Y=2.07 $X2=0
+ $Y2=0
cc_248 N_A_291_409#_c_285_n N_VPWR_c_623_n 0.0380652f $X=1.6 $Y=2.19 $X2=0 $Y2=0
cc_249 N_A_291_409#_c_287_n N_VPWR_c_623_n 0.00753858f $X=1.765 $Y=2.07 $X2=0
+ $Y2=0
cc_250 N_A_291_409#_M1005_g N_VPWR_c_624_n 8.62694e-19 $X=2.925 $Y=2.545 $X2=0
+ $Y2=0
cc_251 N_A_291_409#_c_285_n N_VPWR_c_624_n 0.0481002f $X=1.6 $Y=2.19 $X2=0 $Y2=0
cc_252 N_A_291_409#_c_286_n N_VPWR_c_624_n 0.0163515f $X=2.8 $Y=2.07 $X2=0 $Y2=0
cc_253 N_A_291_409#_M1005_g N_VPWR_c_625_n 0.011221f $X=2.925 $Y=2.545 $X2=0
+ $Y2=0
cc_254 N_A_291_409#_c_285_n N_VPWR_c_629_n 0.0220321f $X=1.6 $Y=2.19 $X2=0 $Y2=0
cc_255 N_A_291_409#_M1005_g N_VPWR_c_630_n 0.00769046f $X=2.925 $Y=2.545 $X2=0
+ $Y2=0
cc_256 N_A_291_409#_M1005_g N_VPWR_c_622_n 0.00739173f $X=2.925 $Y=2.545 $X2=0
+ $Y2=0
cc_257 N_A_291_409#_c_285_n N_VPWR_c_622_n 0.0125808f $X=1.6 $Y=2.19 $X2=0 $Y2=0
cc_258 N_A_291_409#_c_277_n N_VGND_c_714_n 0.0107714f $X=1.89 $Y=0.48 $X2=0
+ $Y2=0
cc_259 N_A_291_409#_M1006_g N_VGND_c_717_n 0.00359964f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_260 N_A_291_409#_c_277_n N_VGND_c_717_n 0.0197885f $X=1.89 $Y=0.48 $X2=0
+ $Y2=0
cc_261 N_A_291_409#_M1006_g N_VGND_c_719_n 0.00526116f $X=3.055 $Y=0.445 $X2=0
+ $Y2=0
cc_262 N_A_291_409#_c_277_n N_VGND_c_719_n 0.0125808f $X=1.89 $Y=0.48 $X2=0
+ $Y2=0
cc_263 N_A_291_409#_c_278_n N_VGND_c_719_n 0.00919746f $X=2.8 $Y=0.86 $X2=0
+ $Y2=0
cc_264 N_C_M1007_g N_D_c_429_n 0.040473f $X=3.445 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_265 N_C_M1004_g N_D_M1001_g 0.0196512f $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_266 N_C_M1007_g N_D_c_431_n 0.00783362f $X=3.445 $Y=0.445 $X2=0 $Y2=0
cc_267 N_C_c_377_n N_D_c_432_n 0.0118516f $X=3.535 $Y=1.625 $X2=0 $Y2=0
cc_268 N_C_c_376_n N_D_c_433_n 0.0118516f $X=3.535 $Y=1.79 $X2=0 $Y2=0
cc_269 C D 0.0431061f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_270 N_C_c_379_n D 8.31475e-19 $X=3.535 $Y=1.285 $X2=0 $Y2=0
cc_271 C N_D_c_435_n 0.00409697f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_272 N_C_c_379_n N_D_c_435_n 0.0118516f $X=3.535 $Y=1.285 $X2=0 $Y2=0
cc_273 N_C_M1007_g N_A_461_47#_c_490_n 0.0112434f $X=3.445 $Y=0.445 $X2=0 $Y2=0
cc_274 N_C_M1004_g N_A_461_47#_c_515_n 0.0169168f $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_275 C N_A_461_47#_c_515_n 0.00717689f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_276 N_C_M1007_g N_A_461_47#_c_491_n 0.00468984f $X=3.445 $Y=0.445 $X2=0 $Y2=0
cc_277 N_C_M1007_g N_A_461_47#_c_492_n 0.00406237f $X=3.445 $Y=0.445 $X2=0 $Y2=0
cc_278 C N_A_461_47#_c_492_n 0.0177641f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_279 N_C_c_379_n N_A_461_47#_c_492_n 0.00123716f $X=3.535 $Y=1.285 $X2=0 $Y2=0
cc_280 N_C_M1007_g N_A_461_47#_c_493_n 0.00405072f $X=3.445 $Y=0.445 $X2=0 $Y2=0
cc_281 C N_A_461_47#_c_493_n 0.00879384f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_282 N_C_M1004_g N_A_461_47#_c_521_n 0.00416508f $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_283 N_C_M1004_g N_A_461_47#_c_500_n 0.0100273f $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_284 N_C_c_376_n N_A_461_47#_c_502_n 3.10915e-19 $X=3.535 $Y=1.79 $X2=0 $Y2=0
cc_285 N_C_M1004_g N_A_461_47#_c_502_n 0.00506276f $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_286 C N_A_461_47#_c_502_n 0.00668688f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_287 N_C_M1004_g N_A_461_47#_c_504_n 8.38826e-19 $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_288 N_C_M1004_g N_A_461_47#_c_544_n 3.84191e-19 $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_289 N_C_M1004_g N_VPWR_c_625_n 0.00496936f $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_290 N_C_M1004_g N_VPWR_c_626_n 8.63039e-19 $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_291 N_C_M1004_g N_VPWR_c_627_n 0.0086001f $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_292 N_C_M1004_g N_VPWR_c_622_n 0.00903025f $X=3.535 $Y=2.545 $X2=0 $Y2=0
cc_293 N_C_M1007_g N_VGND_c_715_n 0.00211602f $X=3.445 $Y=0.445 $X2=0 $Y2=0
cc_294 N_C_M1007_g N_VGND_c_717_n 0.00419924f $X=3.445 $Y=0.445 $X2=0 $Y2=0
cc_295 N_C_M1007_g N_VGND_c_719_n 0.00551032f $X=3.445 $Y=0.445 $X2=0 $Y2=0
cc_296 N_D_c_429_n N_A_461_47#_c_485_n 0.0120131f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_297 N_D_M1001_g N_A_461_47#_M1015_g 0.0281008f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_298 N_D_c_432_n N_A_461_47#_M1015_g 0.00687047f $X=4.105 $Y=1.625 $X2=0 $Y2=0
cc_299 N_D_c_430_n N_A_461_47#_c_488_n 0.00879872f $X=4.015 $Y=0.805 $X2=0 $Y2=0
cc_300 N_D_c_432_n N_A_461_47#_c_489_n 0.012903f $X=4.105 $Y=1.625 $X2=0 $Y2=0
cc_301 N_D_c_429_n N_A_461_47#_c_490_n 0.00108063f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_302 N_D_c_429_n N_A_461_47#_c_491_n 0.00105416f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_303 N_D_c_430_n N_A_461_47#_c_492_n 0.0126085f $X=4.015 $Y=0.805 $X2=0 $Y2=0
cc_304 N_D_c_431_n N_A_461_47#_c_492_n 0.0047468f $X=4.105 $Y=1.12 $X2=0 $Y2=0
cc_305 D N_A_461_47#_c_492_n 0.0245051f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_306 N_D_c_435_n N_A_461_47#_c_492_n 0.00123061f $X=4.105 $Y=1.285 $X2=0 $Y2=0
cc_307 N_D_M1001_g N_A_461_47#_c_521_n 0.00415929f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_308 N_D_M1001_g N_A_461_47#_c_500_n 0.00990719f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_309 N_D_M1001_g N_A_461_47#_c_501_n 0.0184003f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_310 N_D_c_433_n N_A_461_47#_c_501_n 5.43485e-19 $X=4.105 $Y=1.79 $X2=0 $Y2=0
cc_311 D N_A_461_47#_c_501_n 0.0223517f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_312 N_D_M1001_g N_A_461_47#_c_502_n 0.00161889f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_313 D N_A_461_47#_c_502_n 0.00193735f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_314 N_D_c_431_n N_A_461_47#_c_494_n 0.00369602f $X=4.105 $Y=1.12 $X2=0 $Y2=0
cc_315 D N_A_461_47#_c_494_n 0.00115784f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_316 D N_A_461_47#_c_495_n 0.0492653f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_317 N_D_c_435_n N_A_461_47#_c_495_n 0.00135938f $X=4.105 $Y=1.285 $X2=0 $Y2=0
cc_318 N_D_M1001_g N_A_461_47#_c_496_n 0.00356794f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_319 N_D_c_433_n N_A_461_47#_c_496_n 0.00135938f $X=4.105 $Y=1.79 $X2=0 $Y2=0
cc_320 N_D_M1001_g N_A_461_47#_c_544_n 0.00297707f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_321 N_D_c_431_n N_A_461_47#_c_497_n 0.00584957f $X=4.105 $Y=1.12 $X2=0 $Y2=0
cc_322 D N_A_461_47#_c_497_n 5.58507e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_323 N_D_c_435_n N_A_461_47#_c_497_n 0.012903f $X=4.105 $Y=1.285 $X2=0 $Y2=0
cc_324 N_D_c_432_n N_A_461_47#_c_498_n 0.00135938f $X=4.105 $Y=1.625 $X2=0 $Y2=0
cc_325 N_D_M1001_g N_VPWR_c_626_n 0.0177086f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_326 N_D_M1001_g N_VPWR_c_627_n 0.00769046f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_327 N_D_M1001_g N_VPWR_c_622_n 0.0134474f $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_328 N_D_M1001_g X 9.22088e-19 $X=4.065 $Y=2.545 $X2=0 $Y2=0
cc_329 N_D_c_429_n N_VGND_c_715_n 0.0107519f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_330 N_D_c_430_n N_VGND_c_715_n 0.00468659f $X=4.015 $Y=0.805 $X2=0 $Y2=0
cc_331 N_D_c_429_n N_VGND_c_717_n 0.00486043f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_332 N_D_c_429_n N_VGND_c_719_n 0.00439113f $X=3.835 $Y=0.73 $X2=0 $Y2=0
cc_333 N_A_461_47#_c_515_n N_VPWR_M1005_d 0.0114735f $X=3.635 $Y=2.42 $X2=0
+ $Y2=0
cc_334 N_A_461_47#_c_501_n N_VPWR_M1001_d 0.00391101f $X=4.45 $Y=2.055 $X2=0
+ $Y2=0
cc_335 N_A_461_47#_c_504_n N_VPWR_c_624_n 0.048772f $X=2.66 $Y=2.5 $X2=0 $Y2=0
cc_336 N_A_461_47#_c_515_n N_VPWR_c_625_n 0.0203106f $X=3.635 $Y=2.42 $X2=0
+ $Y2=0
cc_337 N_A_461_47#_c_500_n N_VPWR_c_625_n 0.0101276f $X=3.8 $Y=2.9 $X2=0 $Y2=0
cc_338 N_A_461_47#_c_504_n N_VPWR_c_625_n 0.0250385f $X=2.66 $Y=2.5 $X2=0 $Y2=0
cc_339 N_A_461_47#_M1015_g N_VPWR_c_626_n 0.0108204f $X=4.7 $Y=2.545 $X2=0 $Y2=0
cc_340 N_A_461_47#_c_521_n N_VPWR_c_626_n 9.55415e-19 $X=3.8 $Y=2.19 $X2=0 $Y2=0
cc_341 N_A_461_47#_c_500_n N_VPWR_c_626_n 0.0368658f $X=3.8 $Y=2.9 $X2=0 $Y2=0
cc_342 N_A_461_47#_c_501_n N_VPWR_c_626_n 0.0212953f $X=4.45 $Y=2.055 $X2=0
+ $Y2=0
cc_343 N_A_461_47#_c_544_n N_VPWR_c_626_n 0.0119061f $X=3.8 $Y=2.42 $X2=0 $Y2=0
cc_344 N_A_461_47#_c_500_n N_VPWR_c_627_n 0.021949f $X=3.8 $Y=2.9 $X2=0 $Y2=0
cc_345 N_A_461_47#_c_504_n N_VPWR_c_630_n 0.0219185f $X=2.66 $Y=2.5 $X2=0 $Y2=0
cc_346 N_A_461_47#_M1015_g N_VPWR_c_631_n 0.0086001f $X=4.7 $Y=2.545 $X2=0 $Y2=0
cc_347 N_A_461_47#_M1015_g N_VPWR_c_622_n 0.0165658f $X=4.7 $Y=2.545 $X2=0 $Y2=0
cc_348 N_A_461_47#_c_515_n N_VPWR_c_622_n 0.0148815f $X=3.635 $Y=2.42 $X2=0
+ $Y2=0
cc_349 N_A_461_47#_c_500_n N_VPWR_c_622_n 0.0124703f $X=3.8 $Y=2.9 $X2=0 $Y2=0
cc_350 N_A_461_47#_c_504_n N_VPWR_c_622_n 0.0124654f $X=2.66 $Y=2.5 $X2=0 $Y2=0
cc_351 N_A_461_47#_c_485_n N_X_c_689_n 0.00137089f $X=4.405 $Y=0.73 $X2=0 $Y2=0
cc_352 N_A_461_47#_c_487_n N_X_c_689_n 0.00861434f $X=4.765 $Y=0.73 $X2=0 $Y2=0
cc_353 N_A_461_47#_c_494_n N_X_c_689_n 0.00141803f $X=4.645 $Y=1.135 $X2=0 $Y2=0
cc_354 N_A_461_47#_M1015_g X 0.0230055f $X=4.7 $Y=2.545 $X2=0 $Y2=0
cc_355 N_A_461_47#_c_501_n X 0.0130802f $X=4.45 $Y=2.055 $X2=0 $Y2=0
cc_356 N_A_461_47#_c_496_n X 0.00342469f $X=4.535 $Y=1.97 $X2=0 $Y2=0
cc_357 N_A_461_47#_c_498_n X 0.00204411f $X=4.645 $Y=1.61 $X2=0 $Y2=0
cc_358 N_A_461_47#_M1015_g N_X_c_690_n 0.00709538f $X=4.7 $Y=2.545 $X2=0 $Y2=0
cc_359 N_A_461_47#_c_487_n N_X_c_690_n 0.00780981f $X=4.765 $Y=0.73 $X2=0 $Y2=0
cc_360 N_A_461_47#_c_494_n N_X_c_690_n 0.021384f $X=4.645 $Y=1.135 $X2=0 $Y2=0
cc_361 N_A_461_47#_c_495_n N_X_c_690_n 0.034525f $X=4.645 $Y=1.415 $X2=0 $Y2=0
cc_362 N_A_461_47#_c_496_n N_X_c_690_n 0.0116742f $X=4.535 $Y=1.97 $X2=0 $Y2=0
cc_363 N_A_461_47#_c_497_n N_X_c_690_n 0.011919f $X=4.675 $Y=1.105 $X2=0 $Y2=0
cc_364 N_A_461_47#_c_485_n N_VGND_c_715_n 0.00790169f $X=4.405 $Y=0.73 $X2=0
+ $Y2=0
cc_365 N_A_461_47#_c_490_n N_VGND_c_715_n 0.0128489f $X=3.31 $Y=0.43 $X2=0 $Y2=0
cc_366 N_A_461_47#_c_492_n N_VGND_c_715_n 0.0218449f $X=4.45 $Y=0.855 $X2=0
+ $Y2=0
cc_367 N_A_461_47#_c_490_n N_VGND_c_717_n 0.0658094f $X=3.31 $Y=0.43 $X2=0 $Y2=0
cc_368 N_A_461_47#_c_485_n N_VGND_c_718_n 0.00585385f $X=4.405 $Y=0.73 $X2=0
+ $Y2=0
cc_369 N_A_461_47#_c_487_n N_VGND_c_718_n 0.00547815f $X=4.765 $Y=0.73 $X2=0
+ $Y2=0
cc_370 N_A_461_47#_c_488_n N_VGND_c_718_n 6.21075e-19 $X=4.765 $Y=0.805 $X2=0
+ $Y2=0
cc_371 N_A_461_47#_M1014_s N_VGND_c_719_n 0.00232217f $X=2.305 $Y=0.235 $X2=0
+ $Y2=0
cc_372 N_A_461_47#_c_485_n N_VGND_c_719_n 0.00649787f $X=4.405 $Y=0.73 $X2=0
+ $Y2=0
cc_373 N_A_461_47#_c_487_n N_VGND_c_719_n 0.0108866f $X=4.765 $Y=0.73 $X2=0
+ $Y2=0
cc_374 N_A_461_47#_c_488_n N_VGND_c_719_n 8.18184e-19 $X=4.765 $Y=0.805 $X2=0
+ $Y2=0
cc_375 N_A_461_47#_c_490_n N_VGND_c_719_n 0.0435153f $X=3.31 $Y=0.43 $X2=0 $Y2=0
cc_376 N_A_461_47#_c_492_n N_VGND_c_719_n 0.0226213f $X=4.45 $Y=0.855 $X2=0
+ $Y2=0
cc_377 N_A_461_47#_c_494_n N_VGND_c_719_n 0.00634285f $X=4.645 $Y=1.135 $X2=0
+ $Y2=0
cc_378 N_A_461_47#_c_490_n A_548_47# 0.00247906f $X=3.31 $Y=0.43 $X2=-0.19
+ $Y2=-0.245
cc_379 N_A_461_47#_c_490_n A_626_47# 0.00623866f $X=3.31 $Y=0.43 $X2=-0.19
+ $Y2=-0.245
cc_380 N_A_461_47#_c_491_n A_626_47# 6.88945e-19 $X=3.395 $Y=0.77 $X2=-0.19
+ $Y2=-0.245
cc_381 N_VPWR_c_626_n X 0.0374288f $X=4.33 $Y=2.485 $X2=0 $Y2=0
cc_382 N_VPWR_c_631_n X 0.0260776f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_383 N_VPWR_c_622_n X 0.0149024f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_384 N_X_c_689_n N_VGND_c_715_n 0.00940253f $X=5.105 $Y=0.47 $X2=0 $Y2=0
cc_385 N_X_c_689_n N_VGND_c_718_n 0.0220603f $X=5.105 $Y=0.47 $X2=0 $Y2=0
cc_386 N_X_M1000_d N_VGND_c_719_n 0.00233022f $X=4.84 $Y=0.235 $X2=0 $Y2=0
cc_387 N_X_c_689_n N_VGND_c_719_n 0.014194f $X=5.105 $Y=0.47 $X2=0 $Y2=0
cc_388 N_VGND_c_719_n A_548_47# 0.00193256f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
cc_389 N_VGND_c_719_n A_626_47# 0.00193248f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
cc_390 N_VGND_c_719_n A_704_47# 0.00327011f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
cc_391 N_VGND_c_719_n A_896_47# 0.00490351f $X=5.04 $Y=0 $X2=-0.19 $Y2=-0.245
