* File: sky130_fd_sc_lp__fa_lp.spice
* Created: Fri Aug 28 10:35:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__fa_lp.pex.spice"
.subckt sky130_fd_sc_lp__fa_lp  VNB VPB B CIN A COUT VPWR SUM VGND
* 
* VGND	VGND
* SUM	SUM
* VPWR	VPWR
* COUT	COUT
* A	A
* CIN	CIN
* B	B
* VPB	VPB
* VNB	VNB
MM1018 A_134_85# N_A_84_209#_M1018_g N_COUT_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_84_209#_M1005_g A_134_85# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_M1019_g N_A_355_141#_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.09345 AS=0.1533 PD=0.865 PS=1.57 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.3
+ SB=75006.9 A=0.063 P=1.14 MULT=1
MM1020 A_577_141# N_A_M1020_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.09345 PD=0.66 PS=0.865 NRD=18.564 NRS=47.136 M=1 R=2.8 SA=75000.9
+ SB=75006.3 A=0.063 P=1.14 MULT=1
MM1007 N_A_84_209#_M1007_d N_B_M1007_g A_577_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.3
+ SB=75005.9 A=0.063 P=1.14 MULT=1
MM1002 N_A_355_141#_M1002_d N_CIN_M1002_g N_A_84_209#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.145325 AS=0.0882 PD=1.225 PS=0.84 NRD=83.136 NRS=39.996 M=1 R=2.8
+ SA=75001.8 SB=75005.3 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_B_M1015_g N_A_355_141#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.145325 AS=0.145325 PD=1.225 PS=1.225 NRD=83.136 NRS=83.136 M=1 R=2.8
+ SA=75002.4 SB=75004.7 A=0.063 P=1.14 MULT=1
MM1024 N_A_1005_141#_M1024_d N_B_M1024_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.42
+ AD=0.145325 AS=0.145325 PD=1.225 PS=1.225 NRD=83.136 NRS=83.136 M=1 R=2.8
+ SA=75003 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_CIN_M1004_g N_A_1005_141#_M1024_d VNB NSHORT L=0.15
+ W=0.42 AD=0.35175 AS=0.145325 PD=2.095 PS=1.225 NRD=0 NRS=83.136 M=1 R=2.8
+ SA=75003.6 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1008 N_A_1005_141#_M1008_d N_A_M1008_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.35175 PD=0.7 PS=2.095 NRD=0 NRS=398.568 M=1 R=2.8 SA=75005.4
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1010 N_A_1574_141#_M1010_d N_A_84_209#_M1010_g N_A_1005_141#_M1008_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.0861 AS=0.0588 PD=0.83 PS=0.7 NRD=37.14 NRS=0 M=1
+ R=2.8 SA=75005.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1022 A_1686_141# N_CIN_M1022_g N_A_1574_141#_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0861 PD=0.66 PS=0.83 NRD=18.564 NRS=0 M=1 R=2.8 SA=75006.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1012 A_1764_141# N_B_M1012_g A_1686_141# VNB NSHORT L=0.15 W=0.42 AD=0.101062
+ AS=0.0504 PD=1.12 PS=0.66 NRD=53.028 NRS=18.564 M=1 R=2.8 SA=75006.8
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g A_1764_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.101062 PD=0.755 PS=1.12 NRD=0 NRS=53.028 M=1 R=2.8 SA=75000.9
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 A_1956_66# N_A_1574_141#_M1006_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.07035 PD=0.63 PS=0.755 NRD=14.28 NRS=15.708 M=1 R=2.8
+ SA=75001.4 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1026 N_SUM_M1026_d N_A_1574_141#_M1026_g A_1956_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_84_209#_M1014_g N_COUT_M1014_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1029 N_VPWR_M1029_d N_A_M1029_g N_A_245_409#_M1029_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1021 N_A_458_409#_M1021_d N_A_M1021_g N_VPWR_M1029_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1011 N_A_84_209#_M1011_d N_B_M1011_g N_A_245_409#_M1011_s VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.46 PD=1.28 PS=2.92 NRD=0 NRS=34.4553 M=1 R=4 SA=125000
+ SB=125007 A=0.25 P=2.5 MULT=1
MM1027 N_A_458_409#_M1027_d N_CIN_M1027_g N_A_84_209#_M1011_d VPB PHIGHVT L=0.25
+ W=1 AD=0.19 AS=0.14 PD=1.38 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125006
+ A=0.25 P=2.5 MULT=1
MM1016 N_VPWR_M1016_d N_B_M1016_g N_A_458_409#_M1027_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.19 PD=1.28 PS=1.38 NRD=0 NRS=19.7 M=1 R=4 SA=125001 SB=125006
+ A=0.25 P=2.5 MULT=1
MM1000 N_A_1049_419#_M1000_d N_B_M1000_g N_VPWR_M1016_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125005 A=0.25
+ P=2.5 MULT=1
MM1028 N_VPWR_M1028_d N_CIN_M1028_g N_A_1049_419#_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.7575 AS=0.14 PD=2.515 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125005
+ A=0.25 P=2.5 MULT=1
MM1003 N_A_1049_419#_M1003_d N_A_M1003_g N_VPWR_M1028_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.7575 PD=1.28 PS=2.515 NRD=0 NRS=243.275 M=1 R=4 SA=125004
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1023 N_A_1574_141#_M1023_d N_A_84_209#_M1023_g N_A_1049_419#_M1003_d VPB
+ PHIGHVT L=0.25 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4
+ SA=125005 SB=125002 A=0.25 P=2.5 MULT=1
MM1009 A_1720_419# N_CIN_M1009_g N_A_1574_141#_M1023_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.14 PD=1.24 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125005 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1025 A_1818_419# N_B_M1025_g A_1720_419# VPB PHIGHVT L=0.25 W=1 AD=0.135
+ AS=0.12 PD=1.27 PS=1.24 NRD=15.7403 NRS=12.7853 M=1 R=4 SA=125006 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1017 N_VPWR_M1017_d N_A_M1017_g A_1818_419# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.135 PD=1.28 PS=1.27 NRD=0 NRS=15.7403 M=1 R=4 SA=125006 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1001 N_SUM_M1001_d N_A_1574_141#_M1001_g N_VPWR_M1017_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125007 SB=125000
+ A=0.25 P=2.5 MULT=1
DX30_noxref VNB VPB NWDIODE A=20.4031 P=25.61
*
.include "sky130_fd_sc_lp__fa_lp.pxi.spice"
*
.ends
*
*
