* File: sky130_fd_sc_lp__buflp_0.pxi.spice
* Created: Wed Sep  2 09:36:21 2020
* 
x_PM_SKY130_FD_SC_LP__BUFLP_0%A N_A_M1007_g N_A_M1006_g N_A_M1003_g N_A_M1000_g
+ A A A A N_A_c_41_n PM_SKY130_FD_SC_LP__BUFLP_0%A
x_PM_SKY130_FD_SC_LP__BUFLP_0%A_36_120# N_A_36_120#_M1007_s N_A_36_120#_M1006_s
+ N_A_36_120#_M1002_g N_A_36_120#_M1004_g N_A_36_120#_M1005_g
+ N_A_36_120#_M1001_g N_A_36_120#_c_81_n N_A_36_120#_c_90_n N_A_36_120#_c_82_n
+ N_A_36_120#_c_83_n N_A_36_120#_c_84_n N_A_36_120#_c_85_n N_A_36_120#_c_86_n
+ N_A_36_120#_c_87_n PM_SKY130_FD_SC_LP__BUFLP_0%A_36_120#
x_PM_SKY130_FD_SC_LP__BUFLP_0%VPWR N_VPWR_M1000_d N_VPWR_c_141_n VPWR
+ N_VPWR_c_142_n N_VPWR_c_143_n N_VPWR_c_140_n N_VPWR_c_145_n
+ PM_SKY130_FD_SC_LP__BUFLP_0%VPWR
x_PM_SKY130_FD_SC_LP__BUFLP_0%X N_X_M1005_d N_X_M1001_d X X X X X X X
+ PM_SKY130_FD_SC_LP__BUFLP_0%X
x_PM_SKY130_FD_SC_LP__BUFLP_0%VGND N_VGND_M1003_d N_VGND_c_181_n VGND
+ N_VGND_c_182_n N_VGND_c_183_n N_VGND_c_184_n N_VGND_c_185_n
+ PM_SKY130_FD_SC_LP__BUFLP_0%VGND
cc_1 VNB N_A_M1007_g 0.0466811f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.81
cc_2 VNB N_A_M1003_g 0.0369896f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.81
cc_3 VNB A 0.00225372f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_c_41_n 0.00718801f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.765
cc_5 VNB N_A_36_120#_M1002_g 0.0197921f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.6
cc_6 VNB N_A_36_120#_M1005_g 0.0236954f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_7 VNB N_A_36_120#_M1001_g 0.0164857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_36_120#_c_81_n 0.0279118f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.665
cc_9 VNB N_A_36_120#_c_82_n 0.0284375f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.405
cc_10 VNB N_A_36_120#_c_83_n 0.013969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_36_120#_c_84_n 0.0206657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_36_120#_c_85_n 0.00893146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_36_120#_c_86_n 0.00248963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_36_120#_c_87_n 0.0199719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_140_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_16 VNB X 0.0617467f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.66
cc_17 VNB N_VGND_c_181_n 0.0251566f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.66
cc_18 VNB N_VGND_c_182_n 0.0317002f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.81
cc_19 VNB N_VGND_c_183_n 0.0337328f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_20 VNB N_VGND_c_184_n 0.188179f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_21 VNB N_VGND_c_185_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_A_M1006_g 0.0224434f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.66
cc_23 VPB N_A_M1000_g 0.0200132f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.66
cc_24 VPB A 0.00239195f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_25 VPB N_A_c_41_n 0.0686462f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.765
cc_26 VPB N_A_36_120#_M1004_g 0.0296211f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=2.27
cc_27 VPB N_A_36_120#_M1001_g 0.0460288f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_A_36_120#_c_90_n 0.0164185f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.765
cc_29 VPB N_A_36_120#_c_83_n 0.0611351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_A_36_120#_c_86_n 0.00218298f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_A_36_120#_c_87_n 0.00404413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_141_n 0.022142f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.66
cc_33 VPB N_VPWR_c_142_n 0.0338496f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.81
cc_34 VPB N_VPWR_c_143_n 0.0292778f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_35 VPB N_VPWR_c_140_n 0.0788362f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_36 VPB N_VPWR_c_145_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB X 0.0603456f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.66
cc_38 N_A_M1003_g N_A_36_120#_M1002_g 0.0167142f $X=0.93 $Y=0.81 $X2=0 $Y2=0
cc_39 A N_A_36_120#_M1004_g 0.00182354f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_40 N_A_c_41_n N_A_36_120#_M1004_g 0.0218336f $X=0.77 $Y=1.765 $X2=0 $Y2=0
cc_41 N_A_M1003_g N_A_36_120#_c_81_n 0.0182642f $X=0.93 $Y=0.81 $X2=0 $Y2=0
cc_42 N_A_M1007_g N_A_36_120#_c_82_n 0.015833f $X=0.54 $Y=0.81 $X2=0 $Y2=0
cc_43 N_A_M1003_g N_A_36_120#_c_82_n 0.00214178f $X=0.93 $Y=0.81 $X2=0 $Y2=0
cc_44 N_A_M1007_g N_A_36_120#_c_83_n 0.0281953f $X=0.54 $Y=0.81 $X2=0 $Y2=0
cc_45 N_A_M1006_g N_A_36_120#_c_83_n 0.0050011f $X=0.565 $Y=2.66 $X2=0 $Y2=0
cc_46 A N_A_36_120#_c_83_n 0.0873586f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_47 N_A_M1007_g N_A_36_120#_c_84_n 0.0144017f $X=0.54 $Y=0.81 $X2=0 $Y2=0
cc_48 N_A_M1003_g N_A_36_120#_c_84_n 0.0159121f $X=0.93 $Y=0.81 $X2=0 $Y2=0
cc_49 A N_A_36_120#_c_84_n 0.0269732f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_50 N_A_c_41_n N_A_36_120#_c_84_n 3.63979e-19 $X=0.77 $Y=1.765 $X2=0 $Y2=0
cc_51 N_A_M1007_g N_A_36_120#_c_85_n 0.00513266f $X=0.54 $Y=0.81 $X2=0 $Y2=0
cc_52 N_A_M1003_g N_A_36_120#_c_86_n 0.00243994f $X=0.93 $Y=0.81 $X2=0 $Y2=0
cc_53 A N_A_36_120#_c_86_n 0.0152668f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_54 A N_A_36_120#_c_87_n 0.00108855f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_55 N_A_c_41_n N_A_36_120#_c_87_n 0.0182642f $X=0.77 $Y=1.765 $X2=0 $Y2=0
cc_56 A N_VPWR_c_141_n 0.0498171f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_57 N_A_c_41_n N_VPWR_c_141_n 0.00890612f $X=0.77 $Y=1.765 $X2=0 $Y2=0
cc_58 N_A_M1006_g N_VPWR_c_142_n 0.00482473f $X=0.565 $Y=2.66 $X2=0 $Y2=0
cc_59 N_A_M1000_g N_VPWR_c_142_n 0.00464052f $X=0.955 $Y=2.66 $X2=0 $Y2=0
cc_60 A N_VPWR_c_142_n 0.0104923f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_61 N_A_M1006_g N_VPWR_c_140_n 0.00517496f $X=0.565 $Y=2.66 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_VPWR_c_140_n 0.00517496f $X=0.955 $Y=2.66 $X2=0 $Y2=0
cc_63 A N_VPWR_c_140_n 0.0113503f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_64 N_A_M1007_g N_VGND_c_181_n 0.0018473f $X=0.54 $Y=0.81 $X2=0 $Y2=0
cc_65 N_A_M1003_g N_VGND_c_181_n 0.0125894f $X=0.93 $Y=0.81 $X2=0 $Y2=0
cc_66 N_A_M1007_g N_VGND_c_182_n 0.00412501f $X=0.54 $Y=0.81 $X2=0 $Y2=0
cc_67 N_A_M1003_g N_VGND_c_182_n 0.00356352f $X=0.93 $Y=0.81 $X2=0 $Y2=0
cc_68 N_A_M1007_g N_VGND_c_184_n 0.00476395f $X=0.54 $Y=0.81 $X2=0 $Y2=0
cc_69 N_A_M1003_g N_VGND_c_184_n 0.00400172f $X=0.93 $Y=0.81 $X2=0 $Y2=0
cc_70 N_A_36_120#_M1004_g N_VPWR_c_141_n 0.0143841f $X=1.5 $Y=2.55 $X2=0 $Y2=0
cc_71 N_A_36_120#_M1001_g N_VPWR_c_141_n 0.00125969f $X=1.89 $Y=2.55 $X2=0 $Y2=0
cc_72 N_A_36_120#_c_90_n N_VPWR_c_141_n 0.00129266f $X=1.41 $Y=1.88 $X2=0 $Y2=0
cc_73 N_A_36_120#_c_86_n N_VPWR_c_141_n 0.0108833f $X=1.41 $Y=1.375 $X2=0 $Y2=0
cc_74 N_A_36_120#_c_83_n N_VPWR_c_142_n 0.00892695f $X=0.35 $Y=2.66 $X2=0 $Y2=0
cc_75 N_A_36_120#_M1004_g N_VPWR_c_143_n 0.00426961f $X=1.5 $Y=2.55 $X2=0 $Y2=0
cc_76 N_A_36_120#_M1001_g N_VPWR_c_143_n 0.00375632f $X=1.89 $Y=2.55 $X2=0 $Y2=0
cc_77 N_A_36_120#_M1004_g N_VPWR_c_140_n 0.00434697f $X=1.5 $Y=2.55 $X2=0 $Y2=0
cc_78 N_A_36_120#_M1001_g N_VPWR_c_140_n 0.00517496f $X=1.89 $Y=2.55 $X2=0 $Y2=0
cc_79 N_A_36_120#_c_83_n N_VPWR_c_140_n 0.00951858f $X=0.35 $Y=2.66 $X2=0 $Y2=0
cc_80 N_A_36_120#_M1002_g X 0.00244234f $X=1.36 $Y=0.81 $X2=0 $Y2=0
cc_81 N_A_36_120#_M1005_g X 0.0206271f $X=1.75 $Y=0.81 $X2=0 $Y2=0
cc_82 N_A_36_120#_M1001_g X 0.0449164f $X=1.89 $Y=2.55 $X2=0 $Y2=0
cc_83 N_A_36_120#_c_81_n X 0.0113602f $X=1.89 $Y=1.285 $X2=0 $Y2=0
cc_84 N_A_36_120#_c_86_n X 0.0441875f $X=1.41 $Y=1.375 $X2=0 $Y2=0
cc_85 N_A_36_120#_c_87_n X 0.0128971f $X=1.41 $Y=1.375 $X2=0 $Y2=0
cc_86 N_A_36_120#_M1002_g N_VGND_c_181_n 0.0124649f $X=1.36 $Y=0.81 $X2=0 $Y2=0
cc_87 N_A_36_120#_M1005_g N_VGND_c_181_n 0.0016134f $X=1.75 $Y=0.81 $X2=0 $Y2=0
cc_88 N_A_36_120#_c_81_n N_VGND_c_181_n 3.13156e-19 $X=1.89 $Y=1.285 $X2=0 $Y2=0
cc_89 N_A_36_120#_c_82_n N_VGND_c_181_n 0.0145731f $X=0.325 $Y=0.81 $X2=0 $Y2=0
cc_90 N_A_36_120#_c_84_n N_VGND_c_181_n 0.0220609f $X=1.245 $Y=1.295 $X2=0 $Y2=0
cc_91 N_A_36_120#_c_86_n N_VGND_c_181_n 0.0055918f $X=1.41 $Y=1.375 $X2=0 $Y2=0
cc_92 N_A_36_120#_c_82_n N_VGND_c_182_n 0.00742154f $X=0.325 $Y=0.81 $X2=0 $Y2=0
cc_93 N_A_36_120#_M1002_g N_VGND_c_183_n 0.00356352f $X=1.36 $Y=0.81 $X2=0 $Y2=0
cc_94 N_A_36_120#_M1005_g N_VGND_c_183_n 0.00371425f $X=1.75 $Y=0.81 $X2=0 $Y2=0
cc_95 N_A_36_120#_M1002_g N_VGND_c_184_n 0.00400172f $X=1.36 $Y=0.81 $X2=0 $Y2=0
cc_96 N_A_36_120#_M1005_g N_VGND_c_184_n 0.00400172f $X=1.75 $Y=0.81 $X2=0 $Y2=0
cc_97 N_A_36_120#_c_82_n N_VGND_c_184_n 0.0103348f $X=0.325 $Y=0.81 $X2=0 $Y2=0
cc_98 N_VPWR_c_141_n X 0.0153089f $X=1.285 $Y=2.375 $X2=0 $Y2=0
cc_99 N_VPWR_c_143_n X 0.0150695f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_100 N_VPWR_c_140_n X 0.0163455f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_101 X N_VGND_c_181_n 0.0198105f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_102 X N_VGND_c_183_n 0.0154668f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_103 X N_VGND_c_184_n 0.0164919f $X=2.075 $Y=0.47 $X2=0 $Y2=0
