* File: sky130_fd_sc_lp__and3_lp.pxi.spice
* Created: Fri Aug 28 10:06:22 2020
* 
x_PM_SKY130_FD_SC_LP__AND3_LP%A N_A_c_63_n N_A_c_64_n N_A_c_65_n N_A_M1003_g
+ N_A_M1006_g A A N_A_c_68_n N_A_c_69_n PM_SKY130_FD_SC_LP__AND3_LP%A
x_PM_SKY130_FD_SC_LP__AND3_LP%B N_B_c_107_n N_B_M1000_g N_B_M1007_g N_B_c_104_n
+ B N_B_c_105_n N_B_c_106_n PM_SKY130_FD_SC_LP__AND3_LP%B
x_PM_SKY130_FD_SC_LP__AND3_LP%C N_C_c_149_n N_C_M1001_g N_C_M1008_g N_C_c_150_n
+ N_C_c_151_n N_C_c_152_n N_C_c_157_n C N_C_c_153_n N_C_c_154_n
+ PM_SKY130_FD_SC_LP__AND3_LP%C
x_PM_SKY130_FD_SC_LP__AND3_LP%A_38_416# N_A_38_416#_M1006_s N_A_38_416#_M1003_s
+ N_A_38_416#_M1000_d N_A_38_416#_M1002_g N_A_38_416#_M1005_g
+ N_A_38_416#_M1004_g N_A_38_416#_c_201_n N_A_38_416#_c_202_n
+ N_A_38_416#_c_211_n N_A_38_416#_c_203_n N_A_38_416#_c_204_n
+ N_A_38_416#_c_205_n N_A_38_416#_c_213_n N_A_38_416#_c_214_n
+ N_A_38_416#_c_225_n N_A_38_416#_c_206_n N_A_38_416#_c_207_n
+ N_A_38_416#_c_208_n N_A_38_416#_c_209_n PM_SKY130_FD_SC_LP__AND3_LP%A_38_416#
x_PM_SKY130_FD_SC_LP__AND3_LP%VPWR N_VPWR_M1003_d N_VPWR_M1008_d N_VPWR_c_301_n
+ N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_304_n VPWR N_VPWR_c_305_n
+ N_VPWR_c_300_n N_VPWR_c_307_n PM_SKY130_FD_SC_LP__AND3_LP%VPWR
x_PM_SKY130_FD_SC_LP__AND3_LP%X N_X_M1004_d N_X_M1005_d N_X_c_337_n N_X_c_340_n
+ N_X_c_338_n X X N_X_c_339_n PM_SKY130_FD_SC_LP__AND3_LP%X
x_PM_SKY130_FD_SC_LP__AND3_LP%VGND N_VGND_M1001_d N_VGND_c_368_n VGND
+ N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n N_VGND_c_372_n
+ PM_SKY130_FD_SC_LP__AND3_LP%VGND
cc_1 VNB N_A_c_63_n 0.0190737f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.885
cc_2 VNB N_A_c_64_n 0.0255813f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.885
cc_3 VNB N_A_c_65_n 0.0363052f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.525
cc_4 VNB N_A_M1003_g 0.00780336f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.58
cc_5 VNB N_A_M1006_g 0.0217028f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.445
cc_6 VNB N_A_c_68_n 0.0428289f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_7 VNB N_A_c_69_n 0.00561744f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_8 VNB N_B_M1007_g 0.0402066f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.81
cc_9 VNB N_B_c_104_n 0.0186773f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.96
cc_10 VNB N_B_c_105_n 0.0170399f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.45
cc_11 VNB N_B_c_106_n 0.00497282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C_c_149_n 0.0146996f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.885
cc_13 VNB N_C_c_150_n 0.0160561f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.45
cc_14 VNB N_C_c_151_n 0.0176042f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.45
cc_15 VNB N_C_c_152_n 0.0204533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C_c_153_n 0.0167748f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_17 VNB N_C_c_154_n 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_18 VNB N_A_38_416#_M1002_g 0.0183478f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.45
cc_19 VNB N_A_38_416#_M1005_g 0.00926592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_38_416#_M1004_g 0.0209791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_38_416#_c_201_n 0.020168f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_22 VNB N_A_38_416#_c_202_n 0.0149889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_38_416#_c_203_n 0.00642878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_38_416#_c_204_n 0.00749687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_38_416#_c_205_n 0.0352864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_38_416#_c_206_n 0.0191587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_38_416#_c_207_n 5.74534e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_38_416#_c_208_n 0.00284241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_38_416#_c_209_n 0.0318227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_300_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_337_n 0.0180081f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.445
cc_32 VNB N_X_c_338_n 0.0471496f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.375
cc_33 VNB N_X_c_339_n 0.00873257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_368_n 0.00510506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_369_n 0.0456898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_370_n 0.0276259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_371_n 0.172135f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_38 VNB N_VGND_c_372_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_39 VPB N_A_M1003_g 0.0515468f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.58
cc_40 VPB N_A_c_69_n 0.0118607f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.02
cc_41 VPB N_B_c_107_n 0.0128851f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.885
cc_42 VPB N_B_M1000_g 0.0285344f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.525
cc_43 VPB N_B_c_104_n 0.00315682f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.96
cc_44 VPB N_B_c_106_n 0.00239121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_C_M1008_g 0.029187f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.445
cc_46 VPB N_C_c_152_n 0.00347176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_C_c_157_n 0.0139455f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_48 VPB N_C_c_154_n 7.69351e-19 $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.02
cc_49 VPB N_A_38_416#_M1005_g 0.0485626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_38_416#_c_211_n 0.0322735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_38_416#_c_204_n 0.00328099f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_38_416#_c_213_n 0.0158556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_38_416#_c_214_n 0.010077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_301_n 8.75318e-19 $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.96
cc_55 VPB N_VPWR_c_302_n 0.0131183f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.45
cc_56 VPB N_VPWR_c_303_n 0.0182443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_304_n 0.00522215f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.02
cc_58 VPB N_VPWR_c_305_n 0.0231034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_300_n 0.055148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_307_n 0.0249964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_X_c_340_n 0.0536999f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.45
cc_62 VPB N_X_c_338_n 0.0205479f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.375
cc_63 N_A_M1003_g N_B_c_107_n 0.0130365f $X=0.6 $Y=2.58 $X2=-0.19 $Y2=-0.245
cc_64 N_A_M1003_g N_B_M1000_g 0.0280896f $X=0.6 $Y=2.58 $X2=0 $Y2=0
cc_65 N_A_M1006_g N_B_M1007_g 0.0449482f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_66 N_A_c_68_n N_B_M1007_g 0.00188467f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_67 N_A_c_69_n N_B_M1007_g 2.22046e-19 $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_68 N_A_c_65_n N_B_c_104_n 0.0130365f $X=0.6 $Y=1.525 $X2=0 $Y2=0
cc_69 N_A_c_68_n N_B_c_105_n 0.00131516f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_70 N_A_c_65_n N_B_c_106_n 5.59077e-19 $X=0.6 $Y=1.525 $X2=0 $Y2=0
cc_71 N_A_M1003_g N_A_38_416#_c_211_n 0.0208373f $X=0.6 $Y=2.58 $X2=0 $Y2=0
cc_72 N_A_c_63_n N_A_38_416#_c_203_n 0.00252951f $X=0.63 $Y=0.885 $X2=0 $Y2=0
cc_73 N_A_M1006_g N_A_38_416#_c_203_n 0.00497114f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A_c_65_n N_A_38_416#_c_204_n 0.00599269f $X=0.6 $Y=1.525 $X2=0 $Y2=0
cc_75 N_A_M1003_g N_A_38_416#_c_204_n 0.0205916f $X=0.6 $Y=2.58 $X2=0 $Y2=0
cc_76 N_A_c_68_n N_A_38_416#_c_204_n 0.00220637f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_77 N_A_c_69_n N_A_38_416#_c_204_n 0.0541297f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_78 N_A_c_65_n N_A_38_416#_c_214_n 0.0020006f $X=0.6 $Y=1.525 $X2=0 $Y2=0
cc_79 N_A_M1003_g N_A_38_416#_c_214_n 0.0222226f $X=0.6 $Y=2.58 $X2=0 $Y2=0
cc_80 N_A_c_69_n N_A_38_416#_c_214_n 0.0161393f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_81 N_A_M1003_g N_A_38_416#_c_225_n 7.1089e-19 $X=0.6 $Y=2.58 $X2=0 $Y2=0
cc_82 N_A_c_64_n N_A_38_416#_c_206_n 0.0102583f $X=0.435 $Y=0.885 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_A_38_416#_c_206_n 0.00893076f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A_c_69_n N_A_38_416#_c_206_n 0.00866343f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_85 N_A_c_63_n N_A_38_416#_c_207_n 0.00779463f $X=0.63 $Y=0.885 $X2=0 $Y2=0
cc_86 N_A_c_69_n N_A_38_416#_c_207_n 0.012816f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_87 N_A_M1003_g N_VPWR_c_301_n 0.017713f $X=0.6 $Y=2.58 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_VPWR_c_300_n 0.0145382f $X=0.6 $Y=2.58 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_VPWR_c_307_n 0.00818185f $X=0.6 $Y=2.58 $X2=0 $Y2=0
cc_90 N_A_M1006_g N_VGND_c_369_n 0.00359964f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_c_64_n N_VGND_c_371_n 0.00572104f $X=0.435 $Y=0.885 $X2=0 $Y2=0
cc_92 N_A_M1006_g N_VGND_c_371_n 0.00651574f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_c_69_n N_VGND_c_371_n 0.00783511f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_94 N_B_M1007_g N_C_c_149_n 0.0419203f $X=1.095 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_95 N_B_M1000_g N_C_M1008_g 0.0306971f $X=1.13 $Y=2.58 $X2=0 $Y2=0
cc_96 N_B_M1007_g N_C_c_151_n 0.0115744f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_97 N_B_c_104_n N_C_c_152_n 0.01184f $X=1.13 $Y=1.705 $X2=0 $Y2=0
cc_98 N_B_c_107_n N_C_c_157_n 0.01184f $X=1.13 $Y=1.87 $X2=0 $Y2=0
cc_99 N_B_c_105_n N_C_c_153_n 0.01184f $X=1.13 $Y=1.365 $X2=0 $Y2=0
cc_100 N_B_c_106_n N_C_c_153_n 0.00410205f $X=1.13 $Y=1.365 $X2=0 $Y2=0
cc_101 N_B_c_105_n N_C_c_154_n 8.23261e-19 $X=1.13 $Y=1.365 $X2=0 $Y2=0
cc_102 N_B_c_106_n N_C_c_154_n 0.0438819f $X=1.13 $Y=1.365 $X2=0 $Y2=0
cc_103 N_B_M1000_g N_A_38_416#_c_211_n 7.1315e-19 $X=1.13 $Y=2.58 $X2=0 $Y2=0
cc_104 N_B_M1007_g N_A_38_416#_c_203_n 0.00326198f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_105 N_B_M1000_g N_A_38_416#_c_204_n 0.00356753f $X=1.13 $Y=2.58 $X2=0 $Y2=0
cc_106 N_B_M1007_g N_A_38_416#_c_204_n 0.00419164f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_107 N_B_c_105_n N_A_38_416#_c_204_n 0.00556031f $X=1.13 $Y=1.365 $X2=0 $Y2=0
cc_108 N_B_c_106_n N_A_38_416#_c_204_n 0.0483771f $X=1.13 $Y=1.365 $X2=0 $Y2=0
cc_109 N_B_M1007_g N_A_38_416#_c_205_n 0.0127513f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_110 N_B_c_105_n N_A_38_416#_c_205_n 0.00123061f $X=1.13 $Y=1.365 $X2=0 $Y2=0
cc_111 N_B_c_106_n N_A_38_416#_c_205_n 0.0261169f $X=1.13 $Y=1.365 $X2=0 $Y2=0
cc_112 N_B_c_107_n N_A_38_416#_c_213_n 5.79218e-19 $X=1.13 $Y=1.87 $X2=0 $Y2=0
cc_113 N_B_M1000_g N_A_38_416#_c_213_n 0.0189516f $X=1.13 $Y=2.58 $X2=0 $Y2=0
cc_114 N_B_c_106_n N_A_38_416#_c_213_n 0.0264309f $X=1.13 $Y=1.365 $X2=0 $Y2=0
cc_115 N_B_M1000_g N_A_38_416#_c_225_n 0.0183428f $X=1.13 $Y=2.58 $X2=0 $Y2=0
cc_116 N_B_M1007_g N_A_38_416#_c_206_n 0.00141412f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_117 N_B_M1000_g N_VPWR_c_301_n 0.016723f $X=1.13 $Y=2.58 $X2=0 $Y2=0
cc_118 N_B_M1000_g N_VPWR_c_302_n 0.00122348f $X=1.13 $Y=2.58 $X2=0 $Y2=0
cc_119 N_B_M1000_g N_VPWR_c_303_n 0.00818185f $X=1.13 $Y=2.58 $X2=0 $Y2=0
cc_120 N_B_M1000_g N_VPWR_c_300_n 0.0136091f $X=1.13 $Y=2.58 $X2=0 $Y2=0
cc_121 N_B_M1007_g N_VGND_c_368_n 0.00324405f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_122 N_B_M1007_g N_VGND_c_369_n 0.00585385f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_123 N_B_M1007_g N_VGND_c_371_n 0.00639597f $X=1.095 $Y=0.445 $X2=0 $Y2=0
cc_124 N_C_c_149_n N_A_38_416#_M1002_g 0.0127817f $X=1.485 $Y=0.73 $X2=0 $Y2=0
cc_125 N_C_c_150_n N_A_38_416#_M1002_g 0.00679169f $X=1.61 $Y=0.805 $X2=0 $Y2=0
cc_126 N_C_M1008_g N_A_38_416#_M1005_g 0.0151677f $X=1.66 $Y=2.58 $X2=0 $Y2=0
cc_127 N_C_c_157_n N_A_38_416#_M1005_g 0.0122196f $X=1.7 $Y=1.87 $X2=0 $Y2=0
cc_128 N_C_c_151_n N_A_38_416#_c_201_n 0.00679169f $X=1.7 $Y=1.2 $X2=0 $Y2=0
cc_129 N_C_c_152_n N_A_38_416#_c_202_n 0.0122196f $X=1.7 $Y=1.705 $X2=0 $Y2=0
cc_130 N_C_c_150_n N_A_38_416#_c_205_n 0.00795162f $X=1.61 $Y=0.805 $X2=0 $Y2=0
cc_131 N_C_c_151_n N_A_38_416#_c_205_n 0.00776128f $X=1.7 $Y=1.2 $X2=0 $Y2=0
cc_132 N_C_c_153_n N_A_38_416#_c_205_n 0.00123061f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_133 N_C_c_154_n N_A_38_416#_c_205_n 0.0245051f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_134 N_C_M1008_g N_A_38_416#_c_213_n 0.00370641f $X=1.66 $Y=2.58 $X2=0 $Y2=0
cc_135 N_C_c_154_n N_A_38_416#_c_213_n 0.00193735f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_136 N_C_M1008_g N_A_38_416#_c_225_n 0.0177953f $X=1.66 $Y=2.58 $X2=0 $Y2=0
cc_137 N_C_c_151_n N_A_38_416#_c_208_n 0.00101368f $X=1.7 $Y=1.2 $X2=0 $Y2=0
cc_138 N_C_c_153_n N_A_38_416#_c_208_n 0.00117439f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_139 N_C_c_154_n N_A_38_416#_c_208_n 0.0181736f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_140 N_C_c_151_n N_A_38_416#_c_209_n 0.00718191f $X=1.7 $Y=1.2 $X2=0 $Y2=0
cc_141 N_C_c_153_n N_A_38_416#_c_209_n 0.0122196f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_142 N_C_c_154_n N_A_38_416#_c_209_n 0.00354526f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_143 N_C_M1008_g N_VPWR_c_301_n 0.00113006f $X=1.66 $Y=2.58 $X2=0 $Y2=0
cc_144 N_C_M1008_g N_VPWR_c_302_n 0.0226026f $X=1.66 $Y=2.58 $X2=0 $Y2=0
cc_145 N_C_c_157_n N_VPWR_c_302_n 6.10059e-19 $X=1.7 $Y=1.87 $X2=0 $Y2=0
cc_146 N_C_c_154_n N_VPWR_c_302_n 0.00832065f $X=1.7 $Y=1.365 $X2=0 $Y2=0
cc_147 N_C_M1008_g N_VPWR_c_303_n 0.00818185f $X=1.66 $Y=2.58 $X2=0 $Y2=0
cc_148 N_C_M1008_g N_VPWR_c_300_n 0.0136091f $X=1.66 $Y=2.58 $X2=0 $Y2=0
cc_149 N_C_M1008_g N_X_c_340_n 2.80395e-19 $X=1.66 $Y=2.58 $X2=0 $Y2=0
cc_150 N_C_c_149_n N_VGND_c_368_n 0.0134783f $X=1.485 $Y=0.73 $X2=0 $Y2=0
cc_151 N_C_c_150_n N_VGND_c_368_n 0.00391262f $X=1.61 $Y=0.805 $X2=0 $Y2=0
cc_152 N_C_c_149_n N_VGND_c_369_n 0.00486043f $X=1.485 $Y=0.73 $X2=0 $Y2=0
cc_153 N_C_c_149_n N_VGND_c_371_n 0.00455901f $X=1.485 $Y=0.73 $X2=0 $Y2=0
cc_154 N_A_38_416#_c_213_n N_VPWR_M1003_d 0.00176391f $X=1.23 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_38_416#_c_211_n N_VPWR_c_301_n 0.0438173f $X=0.335 $Y=2.225 $X2=0
+ $Y2=0
cc_156 N_A_38_416#_c_214_n N_VPWR_c_301_n 0.0163165f $X=0.785 $Y=2.135 $X2=0
+ $Y2=0
cc_157 N_A_38_416#_c_225_n N_VPWR_c_301_n 0.0438173f $X=1.395 $Y=2.225 $X2=0
+ $Y2=0
cc_158 N_A_38_416#_M1005_g N_VPWR_c_302_n 0.00336873f $X=2.23 $Y=2.58 $X2=0
+ $Y2=0
cc_159 N_A_38_416#_c_213_n N_VPWR_c_302_n 0.0112058f $X=1.23 $Y=2.135 $X2=0
+ $Y2=0
cc_160 N_A_38_416#_c_225_n N_VPWR_c_302_n 0.0556447f $X=1.395 $Y=2.225 $X2=0
+ $Y2=0
cc_161 N_A_38_416#_c_225_n N_VPWR_c_303_n 0.0177952f $X=1.395 $Y=2.225 $X2=0
+ $Y2=0
cc_162 N_A_38_416#_M1005_g N_VPWR_c_305_n 0.00914935f $X=2.23 $Y=2.58 $X2=0
+ $Y2=0
cc_163 N_A_38_416#_M1005_g N_VPWR_c_300_n 0.0169988f $X=2.23 $Y=2.58 $X2=0 $Y2=0
cc_164 N_A_38_416#_c_211_n N_VPWR_c_300_n 0.0125705f $X=0.335 $Y=2.225 $X2=0
+ $Y2=0
cc_165 N_A_38_416#_c_225_n N_VPWR_c_300_n 0.0124497f $X=1.395 $Y=2.225 $X2=0
+ $Y2=0
cc_166 N_A_38_416#_c_211_n N_VPWR_c_307_n 0.019758f $X=0.335 $Y=2.225 $X2=0
+ $Y2=0
cc_167 N_A_38_416#_M1005_g N_X_c_340_n 0.0217278f $X=2.23 $Y=2.58 $X2=0 $Y2=0
cc_168 N_A_38_416#_c_202_n N_X_c_340_n 5.13283e-19 $X=2.27 $Y=1.52 $X2=0 $Y2=0
cc_169 N_A_38_416#_c_208_n N_X_c_340_n 0.00371773f $X=2.27 $Y=1.015 $X2=0 $Y2=0
cc_170 N_A_38_416#_M1005_g N_X_c_338_n 0.0177781f $X=2.23 $Y=2.58 $X2=0 $Y2=0
cc_171 N_A_38_416#_M1004_g N_X_c_338_n 0.00627787f $X=2.36 $Y=0.445 $X2=0 $Y2=0
cc_172 N_A_38_416#_c_201_n N_X_c_338_n 0.00117327f $X=2.36 $Y=0.885 $X2=0 $Y2=0
cc_173 N_A_38_416#_c_208_n N_X_c_338_n 0.0488899f $X=2.27 $Y=1.015 $X2=0 $Y2=0
cc_174 N_A_38_416#_c_209_n N_X_c_338_n 0.0111183f $X=2.27 $Y=1.015 $X2=0 $Y2=0
cc_175 N_A_38_416#_M1002_g N_X_c_339_n 0.00873631f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_176 N_A_38_416#_M1004_g N_X_c_339_n 0.0131518f $X=2.36 $Y=0.445 $X2=0 $Y2=0
cc_177 N_A_38_416#_c_201_n N_X_c_339_n 8.38438e-19 $X=2.36 $Y=0.885 $X2=0 $Y2=0
cc_178 N_A_38_416#_c_205_n N_X_c_339_n 0.0041488f $X=2.105 $Y=0.935 $X2=0 $Y2=0
cc_179 N_A_38_416#_c_208_n N_X_c_339_n 0.0255299f $X=2.27 $Y=1.015 $X2=0 $Y2=0
cc_180 N_A_38_416#_M1002_g N_VGND_c_368_n 0.00722724f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_181 N_A_38_416#_c_205_n N_VGND_c_368_n 0.025292f $X=2.105 $Y=0.935 $X2=0
+ $Y2=0
cc_182 N_A_38_416#_c_206_n N_VGND_c_369_n 0.0269861f $X=0.7 $Y=0.47 $X2=0 $Y2=0
cc_183 N_A_38_416#_M1002_g N_VGND_c_370_n 0.00540301f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_38_416#_M1004_g N_VGND_c_370_n 0.00359964f $X=2.36 $Y=0.445 $X2=0
+ $Y2=0
cc_185 N_A_38_416#_M1006_s N_VGND_c_371_n 0.00233022f $X=0.345 $Y=0.235 $X2=0
+ $Y2=0
cc_186 N_A_38_416#_M1002_g N_VGND_c_371_n 0.00624732f $X=2 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A_38_416#_M1004_g N_VGND_c_371_n 0.00626011f $X=2.36 $Y=0.445 $X2=0
+ $Y2=0
cc_188 N_A_38_416#_c_205_n N_VGND_c_371_n 0.030162f $X=2.105 $Y=0.935 $X2=0
+ $Y2=0
cc_189 N_A_38_416#_c_206_n N_VGND_c_371_n 0.0168622f $X=0.7 $Y=0.47 $X2=0 $Y2=0
cc_190 N_VPWR_c_302_n N_X_c_340_n 0.030661f $X=1.925 $Y=2.225 $X2=0 $Y2=0
cc_191 N_VPWR_c_305_n N_X_c_340_n 0.0281861f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_192 N_VPWR_c_300_n N_X_c_340_n 0.0174072f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_193 N_X_c_339_n N_VGND_c_368_n 0.0317851f $X=2.615 $Y=0.467 $X2=0 $Y2=0
cc_194 N_X_c_337_n N_VGND_c_370_n 0.0113194f $X=2.7 $Y=0.67 $X2=0 $Y2=0
cc_195 N_X_c_339_n N_VGND_c_370_n 0.030545f $X=2.615 $Y=0.467 $X2=0 $Y2=0
cc_196 N_X_M1004_d N_VGND_c_371_n 0.00233008f $X=2.435 $Y=0.235 $X2=0 $Y2=0
cc_197 N_X_c_337_n N_VGND_c_371_n 0.00657784f $X=2.7 $Y=0.67 $X2=0 $Y2=0
cc_198 N_X_c_339_n N_VGND_c_371_n 0.0209098f $X=2.615 $Y=0.467 $X2=0 $Y2=0
cc_199 N_X_c_339_n A_415_47# 9.46545e-19 $X=2.615 $Y=0.467 $X2=-0.19 $Y2=-0.245
cc_200 A_156_47# N_VGND_c_371_n 0.00348365f $X=0.78 $Y=0.235 $X2=2.64 $Y2=0
cc_201 A_234_47# N_VGND_c_371_n 0.00355777f $X=1.17 $Y=0.235 $X2=2.64 $Y2=0
cc_202 N_VGND_c_371_n A_415_47# 0.00169099f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
