* File: sky130_fd_sc_lp__o311ai_lp.pxi.spice
* Created: Wed Sep  2 10:24:06 2020
* 
x_PM_SKY130_FD_SC_LP__O311AI_LP%A1 N_A1_M1008_g N_A1_M1009_g A1 N_A1_c_57_n
+ N_A1_c_58_n PM_SKY130_FD_SC_LP__O311AI_LP%A1
x_PM_SKY130_FD_SC_LP__O311AI_LP%A2 N_A2_M1003_g N_A2_M1000_g A2 A2 A2
+ N_A2_c_84_n N_A2_c_85_n PM_SKY130_FD_SC_LP__O311AI_LP%A2
x_PM_SKY130_FD_SC_LP__O311AI_LP%A3 N_A3_c_120_n N_A3_M1001_g N_A3_M1004_g A3 A3
+ N_A3_c_124_n PM_SKY130_FD_SC_LP__O311AI_LP%A3
x_PM_SKY130_FD_SC_LP__O311AI_LP%B1 N_B1_M1006_g N_B1_M1007_g B1 B1 N_B1_c_158_n
+ PM_SKY130_FD_SC_LP__O311AI_LP%B1
x_PM_SKY130_FD_SC_LP__O311AI_LP%C1 N_C1_M1005_g N_C1_M1002_g C1 N_C1_c_197_n
+ N_C1_c_198_n PM_SKY130_FD_SC_LP__O311AI_LP%C1
x_PM_SKY130_FD_SC_LP__O311AI_LP%VPWR N_VPWR_M1009_s N_VPWR_M1006_d
+ N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n
+ VPWR N_VPWR_c_239_n N_VPWR_c_233_n PM_SKY130_FD_SC_LP__O311AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O311AI_LP%Y N_Y_M1005_d N_Y_M1001_d N_Y_M1002_d
+ N_Y_c_288_n N_Y_c_284_n Y Y Y Y Y Y Y Y PM_SKY130_FD_SC_LP__O311AI_LP%Y
x_PM_SKY130_FD_SC_LP__O311AI_LP%VGND N_VGND_M1008_s N_VGND_M1003_d
+ N_VGND_c_326_n N_VGND_c_327_n N_VGND_c_328_n VGND N_VGND_c_329_n
+ N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n
+ PM_SKY130_FD_SC_LP__O311AI_LP%VGND
x_PM_SKY130_FD_SC_LP__O311AI_LP%A_114_148# N_A_114_148#_M1008_d
+ N_A_114_148#_M1004_d N_A_114_148#_c_360_n N_A_114_148#_c_361_n
+ N_A_114_148#_c_362_n N_A_114_148#_c_363_n
+ PM_SKY130_FD_SC_LP__O311AI_LP%A_114_148#
cc_1 VNB N_A1_M1008_g 0.0243903f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_2 VNB N_A1_c_57_n 0.00400656f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.46
cc_3 VNB N_A1_c_58_n 0.0639633f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.522
cc_4 VNB N_A2_M1003_g 0.0376835f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_5 VNB N_A2_c_84_n 0.00830366f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.46
cc_6 VNB N_A2_c_85_n 0.00304966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A3_c_120_n 0.0106667f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.295
cc_8 VNB N_A3_M1001_g 0.0168433f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_9 VNB N_A3_M1004_g 0.0150303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A3 0.0239255f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.522
cc_11 VNB N_A3_c_124_n 0.0461743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_M1007_g 0.0358454f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_13 VNB B1 0.00339328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_158_n 0.00914984f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.522
cc_15 VNB N_C1_M1005_g 0.0244814f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_16 VNB N_C1_c_197_n 0.0272693f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.46
cc_17 VNB N_C1_c_198_n 0.00171579f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.46
cc_18 VNB N_VPWR_c_233_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB Y 0.0226071f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.46
cc_20 VNB Y 0.0402885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB Y 0.0256949f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_22 VNB N_VGND_c_326_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_23 VNB N_VGND_c_327_n 0.0470797f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_VGND_c_328_n 0.0226342f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.46
cc_25 VNB N_VGND_c_329_n 0.0184158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_330_n 0.0558399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_331_n 0.231209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_332_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_114_148#_c_360_n 0.00606357f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_30 VNB N_A_114_148#_c_361_n 0.0213826f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.522
cc_31 VNB N_A_114_148#_c_362_n 0.0105431f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.46
cc_32 VNB N_A_114_148#_c_363_n 0.00252423f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=1.522
cc_33 VPB N_A1_M1009_g 0.0480492f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_34 VPB N_A1_c_57_n 0.00816414f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.46
cc_35 VPB N_A1_c_58_n 0.00680297f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.522
cc_36 VPB N_A2_M1000_g 0.0232262f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_37 VPB N_A2_c_84_n 0.0195933f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.46
cc_38 VPB N_A2_c_85_n 0.00468283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A3_M1001_g 0.0402619f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.95
cc_40 VPB N_B1_M1006_g 0.0239407f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.95
cc_41 VPB B1 0.00451125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_B1_c_158_n 0.0187776f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.522
cc_43 VPB N_C1_M1002_g 0.0457746f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_44 VPB N_C1_c_197_n 0.00528043f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.46
cc_45 VPB N_C1_c_198_n 0.00240449f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.46
cc_46 VPB N_VPWR_c_234_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_47 VPB N_VPWR_c_235_n 0.0440356f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_48 VPB N_VPWR_c_236_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.522
cc_49 VPB N_VPWR_c_237_n 0.0470343f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.665
cc_50 VPB N_VPWR_c_238_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_239_n 0.0236177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_233_n 0.0475443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB Y 0.0224287f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.665
cc_54 VPB Y 0.028708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB Y 0.0277948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 N_A1_M1008_g N_A2_M1003_g 0.0117807f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_57 N_A1_c_57_n N_A2_M1003_g 0.00141327f $X=0.28 $Y=1.46 $X2=0 $Y2=0
cc_58 N_A1_M1009_g N_A2_M1000_g 0.0695181f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_59 N_A1_c_58_n N_A2_c_84_n 0.0316841f $X=0.495 $Y=1.522 $X2=0 $Y2=0
cc_60 N_A1_M1009_g N_A2_c_85_n 0.00588081f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_61 N_A1_c_57_n N_A2_c_85_n 0.00625527f $X=0.28 $Y=1.46 $X2=0 $Y2=0
cc_62 N_A1_c_58_n N_A2_c_85_n 0.00176131f $X=0.495 $Y=1.522 $X2=0 $Y2=0
cc_63 N_A1_M1009_g N_VPWR_c_235_n 0.0256381f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_64 N_A1_c_57_n N_VPWR_c_235_n 0.020151f $X=0.28 $Y=1.46 $X2=0 $Y2=0
cc_65 N_A1_c_58_n N_VPWR_c_235_n 0.00167176f $X=0.495 $Y=1.522 $X2=0 $Y2=0
cc_66 N_A1_M1009_g N_VPWR_c_237_n 0.008763f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_67 N_A1_M1009_g N_VPWR_c_233_n 0.0144563f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_68 N_A1_M1008_g N_VGND_c_327_n 0.00982452f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_69 N_A1_c_57_n N_VGND_c_327_n 0.0242582f $X=0.28 $Y=1.46 $X2=0 $Y2=0
cc_70 N_A1_c_58_n N_VGND_c_327_n 0.00220957f $X=0.495 $Y=1.522 $X2=0 $Y2=0
cc_71 N_A1_M1008_g N_VGND_c_329_n 0.00298903f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_72 N_A1_M1008_g N_VGND_c_331_n 0.00368577f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_73 N_A1_M1008_g N_A_114_148#_c_360_n 0.00272581f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_74 N_A1_M1008_g N_A_114_148#_c_362_n 0.00257765f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_75 N_A1_c_57_n N_A_114_148#_c_362_n 0.0104995f $X=0.28 $Y=1.46 $X2=0 $Y2=0
cc_76 N_A1_c_58_n N_A_114_148#_c_362_n 0.00210312f $X=0.495 $Y=1.522 $X2=0 $Y2=0
cc_77 N_A2_M1003_g N_A3_c_120_n 0.0109118f $X=0.955 $Y=0.95 $X2=-0.19 $Y2=-0.245
cc_78 N_A2_M1000_g N_A3_M1001_g 0.062353f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_79 N_A2_c_84_n N_A3_M1001_g 0.020056f $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_80 N_A2_c_85_n N_A3_M1001_g 0.0146348f $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_81 N_A2_M1003_g N_A3_c_124_n 0.00893002f $X=0.955 $Y=0.95 $X2=0 $Y2=0
cc_82 N_A2_c_84_n B1 2.79131e-19 $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_83 N_A2_c_85_n B1 0.0348426f $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_84 N_A2_M1000_g N_VPWR_c_235_n 0.00252625f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_85 N_A2_c_85_n N_VPWR_c_235_n 0.0147315f $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_86 N_A2_M1000_g N_VPWR_c_237_n 0.00655603f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_87 N_A2_c_85_n N_VPWR_c_237_n 0.0120368f $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_88 N_A2_M1000_g N_VPWR_c_233_n 0.00810006f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_89 N_A2_c_85_n N_VPWR_c_233_n 0.0138515f $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_90 N_A2_c_85_n A_232_419# 0.010357f $X=1.045 $Y=1.77 $X2=-0.19 $Y2=-0.245
cc_91 N_A2_M1000_g N_Y_c_284_n 0.0010528f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_92 N_A2_c_85_n N_Y_c_284_n 0.0271513f $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_93 N_A2_M1003_g N_VGND_c_327_n 4.45872e-19 $X=0.955 $Y=0.95 $X2=0 $Y2=0
cc_94 N_A2_M1003_g N_VGND_c_328_n 0.00211768f $X=0.955 $Y=0.95 $X2=0 $Y2=0
cc_95 N_A2_M1003_g N_VGND_c_329_n 0.00359559f $X=0.955 $Y=0.95 $X2=0 $Y2=0
cc_96 N_A2_M1003_g N_VGND_c_331_n 0.00438782f $X=0.955 $Y=0.95 $X2=0 $Y2=0
cc_97 N_A2_M1003_g N_A_114_148#_c_360_n 0.00291944f $X=0.955 $Y=0.95 $X2=0 $Y2=0
cc_98 N_A2_M1003_g N_A_114_148#_c_361_n 0.0152194f $X=0.955 $Y=0.95 $X2=0 $Y2=0
cc_99 N_A2_c_84_n N_A_114_148#_c_361_n 0.00124137f $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_100 N_A2_c_85_n N_A_114_148#_c_361_n 0.0330463f $X=1.045 $Y=1.77 $X2=0 $Y2=0
cc_101 N_A3_M1001_g N_B1_M1006_g 0.0247463f $X=1.545 $Y=2.595 $X2=0 $Y2=0
cc_102 N_A3_M1004_g N_B1_M1007_g 0.0239829f $X=1.595 $Y=0.95 $X2=0 $Y2=0
cc_103 A3 N_B1_M1007_g 0.0120447f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_104 N_A3_c_124_n N_B1_M1007_g 0.00125607f $X=1.73 $Y=0.465 $X2=0 $Y2=0
cc_105 N_A3_M1001_g B1 0.0229761f $X=1.545 $Y=2.595 $X2=0 $Y2=0
cc_106 N_A3_M1001_g N_B1_c_158_n 0.0164234f $X=1.545 $Y=2.595 $X2=0 $Y2=0
cc_107 A3 N_C1_M1005_g 0.00152975f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_108 N_A3_M1001_g N_VPWR_c_236_n 0.00103917f $X=1.545 $Y=2.595 $X2=0 $Y2=0
cc_109 N_A3_M1001_g N_VPWR_c_237_n 0.00939541f $X=1.545 $Y=2.595 $X2=0 $Y2=0
cc_110 N_A3_M1001_g N_VPWR_c_233_n 0.0162077f $X=1.545 $Y=2.595 $X2=0 $Y2=0
cc_111 N_A3_M1001_g N_Y_c_284_n 0.0131949f $X=1.545 $Y=2.595 $X2=0 $Y2=0
cc_112 A3 N_VGND_c_328_n 0.029626f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_113 N_A3_c_124_n N_VGND_c_328_n 0.0154353f $X=1.73 $Y=0.465 $X2=0 $Y2=0
cc_114 A3 N_VGND_c_330_n 0.0366812f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_115 N_A3_c_124_n N_VGND_c_330_n 0.00898392f $X=1.73 $Y=0.465 $X2=0 $Y2=0
cc_116 A3 N_VGND_c_331_n 0.026263f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_117 N_A3_c_124_n N_VGND_c_331_n 0.0122736f $X=1.73 $Y=0.465 $X2=0 $Y2=0
cc_118 N_A3_c_120_n N_A_114_148#_c_361_n 0.00815086f $X=1.545 $Y=1.415 $X2=0
+ $Y2=0
cc_119 N_A3_M1001_g N_A_114_148#_c_361_n 0.00832156f $X=1.545 $Y=2.595 $X2=0
+ $Y2=0
cc_120 N_A3_M1004_g N_A_114_148#_c_361_n 0.00634631f $X=1.595 $Y=0.95 $X2=0
+ $Y2=0
cc_121 A3 N_A_114_148#_c_361_n 0.00457812f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_122 N_A3_c_124_n N_A_114_148#_c_361_n 2.61807e-19 $X=1.73 $Y=0.465 $X2=0
+ $Y2=0
cc_123 N_A3_M1004_g N_A_114_148#_c_363_n 0.00463411f $X=1.595 $Y=0.95 $X2=0
+ $Y2=0
cc_124 A3 N_A_114_148#_c_363_n 0.0263086f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_125 N_A3_c_124_n N_A_114_148#_c_363_n 0.0011707f $X=1.73 $Y=0.465 $X2=0 $Y2=0
cc_126 N_B1_M1007_g N_C1_M1005_g 0.0329975f $X=2.185 $Y=0.95 $X2=0 $Y2=0
cc_127 N_B1_M1006_g N_C1_M1002_g 0.0378479f $X=2.075 $Y=2.595 $X2=0 $Y2=0
cc_128 B1 N_C1_M1002_g 0.00873238f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_129 N_B1_c_158_n N_C1_M1002_g 0.0127258f $X=2.095 $Y=1.77 $X2=0 $Y2=0
cc_130 B1 N_C1_c_197_n 5.5354e-19 $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_131 N_B1_c_158_n N_C1_c_197_n 0.0329975f $X=2.095 $Y=1.77 $X2=0 $Y2=0
cc_132 N_B1_M1007_g N_C1_c_198_n 0.00141699f $X=2.185 $Y=0.95 $X2=0 $Y2=0
cc_133 B1 N_C1_c_198_n 0.0136401f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_134 N_B1_c_158_n N_C1_c_198_n 3.95969e-19 $X=2.095 $Y=1.77 $X2=0 $Y2=0
cc_135 B1 N_VPWR_M1006_d 9.31012e-19 $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_136 N_B1_M1006_g N_VPWR_c_236_n 0.0128016f $X=2.075 $Y=2.595 $X2=0 $Y2=0
cc_137 N_B1_M1006_g N_VPWR_c_237_n 0.00840199f $X=2.075 $Y=2.595 $X2=0 $Y2=0
cc_138 N_B1_M1006_g N_VPWR_c_233_n 0.00756435f $X=2.075 $Y=2.595 $X2=0 $Y2=0
cc_139 B1 N_Y_M1001_d 0.00187356f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_140 N_B1_M1006_g N_Y_c_288_n 0.0139016f $X=2.075 $Y=2.595 $X2=0 $Y2=0
cc_141 B1 N_Y_c_288_n 0.0173306f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_142 N_B1_M1006_g N_Y_c_284_n 0.0112789f $X=2.075 $Y=2.595 $X2=0 $Y2=0
cc_143 B1 N_Y_c_284_n 0.0179173f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_144 N_B1_M1007_g Y 0.00157319f $X=2.185 $Y=0.95 $X2=0 $Y2=0
cc_145 N_B1_M1006_g Y 0.00166818f $X=2.075 $Y=2.595 $X2=0 $Y2=0
cc_146 B1 Y 0.00301122f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_147 N_B1_M1007_g N_VGND_c_330_n 4.51359e-19 $X=2.185 $Y=0.95 $X2=0 $Y2=0
cc_148 N_B1_M1007_g N_A_114_148#_c_361_n 0.00457809f $X=2.185 $Y=0.95 $X2=0
+ $Y2=0
cc_149 B1 N_A_114_148#_c_361_n 0.0399407f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_150 N_B1_c_158_n N_A_114_148#_c_361_n 0.00328776f $X=2.095 $Y=1.77 $X2=0
+ $Y2=0
cc_151 N_B1_M1007_g N_A_114_148#_c_363_n 0.0043789f $X=2.185 $Y=0.95 $X2=0 $Y2=0
cc_152 N_C1_M1002_g N_VPWR_c_236_n 0.0121063f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_153 N_C1_M1002_g N_VPWR_c_239_n 0.0091825f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_154 N_C1_M1002_g N_VPWR_c_233_n 0.00925362f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_155 N_C1_M1002_g N_Y_c_288_n 0.0173139f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_156 N_C1_c_198_n N_Y_c_288_n 0.00681033f $X=2.635 $Y=1.53 $X2=0 $Y2=0
cc_157 N_C1_M1002_g N_Y_c_284_n 8.70102e-19 $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_158 N_C1_M1005_g Y 0.00310799f $X=2.545 $Y=0.95 $X2=0 $Y2=0
cc_159 N_C1_M1005_g Y 0.010515f $X=2.545 $Y=0.95 $X2=0 $Y2=0
cc_160 N_C1_c_197_n Y 0.0013327f $X=2.635 $Y=1.53 $X2=0 $Y2=0
cc_161 N_C1_c_198_n Y 0.0157803f $X=2.635 $Y=1.53 $X2=0 $Y2=0
cc_162 N_C1_M1005_g Y 0.00521362f $X=2.545 $Y=0.95 $X2=0 $Y2=0
cc_163 N_C1_M1002_g Y 0.0106237f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_164 N_C1_c_197_n Y 0.0072883f $X=2.635 $Y=1.53 $X2=0 $Y2=0
cc_165 N_C1_c_198_n Y 0.0281023f $X=2.635 $Y=1.53 $X2=0 $Y2=0
cc_166 N_C1_M1002_g Y 0.00852888f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_167 N_C1_c_197_n Y 3.0636e-19 $X=2.635 $Y=1.53 $X2=0 $Y2=0
cc_168 N_C1_c_198_n Y 0.00426389f $X=2.635 $Y=1.53 $X2=0 $Y2=0
cc_169 N_C1_M1002_g Y 0.0155094f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_170 N_C1_M1005_g N_VGND_c_330_n 0.00346978f $X=2.545 $Y=0.95 $X2=0 $Y2=0
cc_171 N_C1_M1005_g N_VGND_c_331_n 0.00438782f $X=2.545 $Y=0.95 $X2=0 $Y2=0
cc_172 N_C1_c_198_n N_A_114_148#_c_361_n 0.00259503f $X=2.635 $Y=1.53 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_233_n A_134_419# 0.00930162f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_174 N_VPWR_c_233_n A_232_419# 0.00594533f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_175 N_VPWR_c_233_n N_Y_M1001_d 0.00223819f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_176 N_VPWR_c_233_n N_Y_M1002_d 0.0023218f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_177 N_VPWR_M1006_d N_Y_c_288_n 0.00856907f $X=2.2 $Y=2.095 $X2=0 $Y2=0
cc_178 N_VPWR_c_236_n N_Y_c_288_n 0.0160925f $X=2.34 $Y=2.895 $X2=0 $Y2=0
cc_179 N_VPWR_c_233_n N_Y_c_288_n 0.0127514f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_180 N_VPWR_c_236_n N_Y_c_284_n 0.0253679f $X=2.34 $Y=2.895 $X2=0 $Y2=0
cc_181 N_VPWR_c_237_n N_Y_c_284_n 0.0177952f $X=2.175 $Y=3.33 $X2=0 $Y2=0
cc_182 N_VPWR_c_233_n N_Y_c_284_n 0.0123247f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_236_n Y 0.0243195f $X=2.34 $Y=2.895 $X2=0 $Y2=0
cc_184 N_VPWR_c_239_n Y 0.0318944f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_185 N_VPWR_c_233_n Y 0.0194728f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_186 Y N_VGND_c_330_n 0.00700678f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_187 Y N_VGND_c_330_n 0.00677452f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_188 Y N_VGND_c_331_n 0.00769349f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_189 Y N_VGND_c_331_n 0.0114827f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_190 Y N_A_114_148#_c_363_n 0.00563544f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_191 N_VGND_c_327_n N_A_114_148#_c_360_n 0.0148853f $X=0.28 $Y=0.915 $X2=0
+ $Y2=0
cc_192 N_VGND_c_328_n N_A_114_148#_c_360_n 0.00148713f $X=1.22 $Y=0.895 $X2=0
+ $Y2=0
cc_193 N_VGND_c_329_n N_A_114_148#_c_360_n 0.00426279f $X=1.055 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_c_331_n N_A_114_148#_c_360_n 0.00707958f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_c_328_n N_A_114_148#_c_361_n 0.0246804f $X=1.22 $Y=0.895 $X2=0
+ $Y2=0
