* File: sky130_fd_sc_lp__inv_8.spice
* Created: Wed Sep  2 09:56:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__inv_8.pex.spice"
.subckt sky130_fd_sc_lp__inv_8  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84 AD=0.2394
+ AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75003.2 A=0.126
+ P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6 SB=75002.8 A=0.126
+ P=1.98 MULT=1
MM1005 N_VGND_M1004_d N_A_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1 SB=75002.4 A=0.126
+ P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5 SB=75001.9 A=0.126
+ P=1.98 MULT=1
MM1010 N_VGND_M1007_d N_A_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9 SB=75001.5 A=0.126
+ P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A_M1012_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4 SB=75001.1 A=0.126
+ P=1.98 MULT=1
MM1013 N_VGND_M1012_d N_A_M1013_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8 SB=75000.6 A=0.126
+ P=1.98 MULT=1
MM1014 N_VGND_M1014_d N_A_M1014_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.84 AD=0.2394
+ AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1002_d N_A_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_Y_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1006_d N_A_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1009_d N_A_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__inv_8.pxi.spice"
*
.ends
*
*
