* File: sky130_fd_sc_lp__a22oi_0.pex.spice
* Created: Wed Sep  2 09:22:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22OI_0%B2 5 9 11 12 13 14 15 20
r34 20 23 77.6472 $w=4.9e-07 $l=5.05e-07 $layer=POLY_cond $X=0.36 $Y=1.005
+ $X2=0.36 $Y2=1.51
r35 20 22 46.2534 $w=4.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.36 $Y=1.005
+ $X2=0.36 $Y2=0.84
r36 14 15 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.665
r37 13 14 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=0.925
+ $X2=0.23 $Y2=1.295
r38 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.28
+ $Y=1.005 $X2=0.28 $Y2=1.005
r39 11 12 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.55 $Y=1.725
+ $X2=0.55 $Y2=1.875
r40 11 23 83.5726 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=0.515 $Y=1.725
+ $X2=0.515 $Y2=1.51
r41 9 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.6 $Y=2.345 $X2=0.6
+ $Y2=1.875
r42 5 22 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.53 $Y=0.445
+ $X2=0.53 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_0%B1 3 7 11 12 13 14 18
r36 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.98
+ $Y=0.98 $X2=0.98 $Y2=0.98
r37 14 19 9.07549 $w=3.98e-07 $l=3.15e-07 $layer=LI1_cond $X=1.095 $Y=1.295
+ $X2=1.095 $Y2=0.98
r38 13 19 1.58461 $w=3.98e-07 $l=5.5e-08 $layer=LI1_cond $X=1.095 $Y=0.925
+ $X2=1.095 $Y2=0.98
r39 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.98 $Y=1.32
+ $X2=0.98 $Y2=0.98
r40 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.32
+ $X2=0.98 $Y2=1.485
r41 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=0.815
+ $X2=0.98 $Y2=0.98
r42 7 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.03 $Y=2.345
+ $X2=1.03 $Y2=1.485
r43 3 10 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.89 $Y=0.445
+ $X2=0.89 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_0%A1 3 7 9 10 11 16
c38 7 0 1.1168e-19 $X=1.46 $Y=2.345
r39 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.32
+ $X2=1.55 $Y2=1.485
r40 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.32
+ $X2=1.55 $Y2=1.155
r41 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.32 $X2=1.55 $Y2=1.32
r42 11 17 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=1.62 $Y=1.295
+ $X2=1.62 $Y2=1.32
r43 10 11 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.62 $Y=0.925
+ $X2=1.62 $Y2=1.295
r44 9 10 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.62 $Y=0.555 $X2=1.62
+ $Y2=0.925
r45 7 19 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.46 $Y=2.345
+ $X2=1.46 $Y2=1.485
r46 3 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.46 $Y=0.445
+ $X2=1.46 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_0%A2 1 3 6 9 13 17 20 21 22 26
c38 13 0 3.34511e-20 $X=2.12 $Y=0.915
r39 21 22 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.13 $Y=0.925
+ $X2=2.13 $Y2=1.295
r40 21 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.12
+ $Y=0.98 $X2=2.12 $Y2=0.98
r41 19 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.12 $Y=1.32
+ $X2=2.12 $Y2=0.98
r42 19 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.12 $Y=1.32
+ $X2=2.12 $Y2=1.485
r43 15 17 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.89 $Y=1.8 $X2=2.03
+ $Y2=1.8
r44 13 26 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=2.12 $Y=0.915
+ $X2=2.12 $Y2=0.98
r45 10 13 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.82 $Y=0.84 $X2=2.12
+ $Y2=0.84
r46 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.03 $Y=1.725
+ $X2=2.03 $Y2=1.8
r47 9 20 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.03 $Y=1.725
+ $X2=2.03 $Y2=1.485
r48 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.89 $Y=1.875
+ $X2=1.89 $Y2=1.8
r49 4 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.89 $Y=1.875 $X2=1.89
+ $Y2=2.345
r50 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.82 $Y=0.765
+ $X2=1.82 $Y2=0.84
r51 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.82 $Y=0.765 $X2=1.82
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_0%A_45_405# 1 2 3 12 14 15 19 20 21 24
c41 24 0 1.1168e-19 $X=2.105 $Y=2.17
r42 22 24 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.125 $Y=1.835
+ $X2=2.125 $Y2=2.17
r43 20 22 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=1.98 $Y=1.75
+ $X2=2.125 $Y2=1.835
r44 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.98 $Y=1.75
+ $X2=1.37 $Y2=1.75
r45 17 19 30.9578 $w=2.53e-07 $l=6.85e-07 $layer=LI1_cond $X=1.242 $Y=2.855
+ $X2=1.242 $Y2=2.17
r46 16 21 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=1.242 $Y=1.835
+ $X2=1.37 $Y2=1.75
r47 16 19 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=1.242 $Y=1.835
+ $X2=1.242 $Y2=2.17
r48 14 17 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.115 $Y=2.94
+ $X2=1.242 $Y2=2.855
r49 14 15 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.115 $Y=2.94
+ $X2=0.455 $Y2=2.94
r50 10 15 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.32 $Y=2.855
+ $X2=0.455 $Y2=2.94
r51 10 12 29.2379 $w=2.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.32 $Y=2.855
+ $X2=0.32 $Y2=2.17
r52 3 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.965
+ $Y=2.025 $X2=2.105 $Y2=2.17
r53 2 19 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.105
+ $Y=2.025 $X2=1.245 $Y2=2.17
r54 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.025 $X2=0.35 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_0%Y 1 2 9 11 14 15 16 17
c36 14 0 9.10919e-20 $X=0.745 $Y=1.665
r37 17 23 8.46325 $w=3.18e-07 $l=2.35e-07 $layer=LI1_cond $X=0.785 $Y=2.405
+ $X2=0.785 $Y2=2.17
r38 16 23 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=0.785 $Y=2.035
+ $X2=0.785 $Y2=2.17
r39 15 16 7.20277 $w=3.18e-07 $l=2e-07 $layer=LI1_cond $X=0.785 $Y=1.835
+ $X2=0.785 $Y2=2.035
r40 14 15 8.64032 $w=3.18e-07 $l=1.7e-07 $layer=LI1_cond $X=0.745 $Y=1.665
+ $X2=0.745 $Y2=1.835
r41 9 11 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.715 $Y=0.43
+ $X2=1.13 $Y2=0.43
r42 7 9 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.63 $Y=0.595
+ $X2=0.715 $Y2=0.43
r43 7 14 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=0.63 $Y=0.595
+ $X2=0.63 $Y2=1.665
r44 2 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.675
+ $Y=2.025 $X2=0.815 $Y2=2.17
r45 1 11 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.235 $X2=1.13 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_0%VPWR 1 6 8 10 20 21 24
r22 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r23 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r24 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r25 18 24 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.675 $Y2=3.33
r26 18 20 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 12 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r28 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 10 24 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.675 $Y2=3.33
r30 10 16 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.54 $Y=3.33 $X2=1.2
+ $Y2=3.33
r31 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r32 8 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.24
+ $Y2=3.33
r33 8 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r34 4 24 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=3.245
+ $X2=1.675 $Y2=3.33
r35 4 6 45.8843 $w=2.68e-07 $l=1.075e-06 $layer=LI1_cond $X=1.675 $Y=3.245
+ $X2=1.675 $Y2=2.17
r36 1 6 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=2.025 $X2=1.675 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_0%VGND 1 2 7 9 11 13 15 17 30
c36 11 0 3.34511e-20 $X=2.11 $Y=0.085
r37 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r40 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r41 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r42 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r43 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 18 26 3.99677 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0 $X2=0.187
+ $Y2=0
r45 18 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.375 $Y=0 $X2=0.72
+ $Y2=0
r46 17 29 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.172
+ $Y2=0
r47 17 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.68
+ $Y2=0
r48 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r49 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r50 11 29 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.172 $Y2=0
r51 11 13 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.43
r52 7 26 3.14639 $w=2.5e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.25 $Y=0.085
+ $X2=0.187 $Y2=0
r53 7 9 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=0.25 $Y=0.085
+ $X2=0.25 $Y2=0.43
r54 2 13 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.035 $Y2=0.43
r55 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.43
.ends

