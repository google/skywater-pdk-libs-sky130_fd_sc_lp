* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
X0 VGND D a_671_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 X a_254_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_851_47# a_929_21# a_254_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_254_21# a_929_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND a_254_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR D a_254_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 X a_254_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_49_131# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_49_131# a_254_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_254_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_49_131# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VPWR a_254_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND a_254_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 X a_254_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VPWR A_N a_929_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 a_671_47# C a_743_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_743_47# a_49_131# a_851_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VPWR a_254_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 X a_254_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VGND A_N a_929_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
