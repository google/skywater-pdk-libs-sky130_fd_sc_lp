* File: sky130_fd_sc_lp__mux4_1.pxi.spice
* Created: Wed Sep  2 10:01:52 2020
* 
x_PM_SKY130_FD_SC_LP__MUX4_1%A1 N_A1_c_219_n N_A1_M1000_g N_A1_M1014_g
+ N_A1_c_225_n A1 A1 A1 N_A1_c_222_n PM_SKY130_FD_SC_LP__MUX4_1%A1
x_PM_SKY130_FD_SC_LP__MUX4_1%A0 N_A0_M1013_g N_A0_M1008_g N_A0_c_259_n
+ N_A0_c_260_n A0 A0 A0 N_A0_c_257_n PM_SKY130_FD_SC_LP__MUX4_1%A0
x_PM_SKY130_FD_SC_LP__MUX4_1%A_254_55# N_A_254_55#_M1011_s N_A_254_55#_M1021_s
+ N_A_254_55#_M1009_g N_A_254_55#_c_301_n N_A_254_55#_c_302_n
+ N_A_254_55#_M1005_g N_A_254_55#_c_304_n N_A_254_55#_c_313_n
+ N_A_254_55#_M1007_g N_A_254_55#_M1024_g N_A_254_55#_c_306_n
+ N_A_254_55#_c_307_n N_A_254_55#_c_315_n N_A_254_55#_c_316_n
+ N_A_254_55#_c_317_n N_A_254_55#_c_318_n N_A_254_55#_c_308_n
+ N_A_254_55#_c_309_n N_A_254_55#_c_310_n N_A_254_55#_c_311_n
+ PM_SKY130_FD_SC_LP__MUX4_1%A_254_55#
x_PM_SKY130_FD_SC_LP__MUX4_1%S0 N_S0_M1018_g N_S0_c_451_n N_S0_c_452_n
+ N_S0_c_461_n N_S0_M1023_g N_S0_c_462_n N_S0_c_463_n N_S0_c_453_n N_S0_M1011_g
+ N_S0_c_454_n N_S0_c_455_n N_S0_c_465_n N_S0_M1021_g N_S0_c_467_n N_S0_c_468_n
+ N_S0_c_469_n N_S0_M1016_g N_S0_c_470_n N_S0_M1003_g N_S0_c_457_n N_S0_c_471_n
+ N_S0_c_458_n N_S0_c_459_n S0 N_S0_c_460_n N_S0_c_473_n
+ PM_SKY130_FD_SC_LP__MUX4_1%S0
x_PM_SKY130_FD_SC_LP__MUX4_1%A3 N_A3_M1019_g N_A3_M1012_g N_A3_c_562_n
+ N_A3_c_563_n N_A3_c_564_n N_A3_c_565_n N_A3_c_566_n A3 A3 N_A3_c_567_n
+ N_A3_c_568_n PM_SKY130_FD_SC_LP__MUX4_1%A3
x_PM_SKY130_FD_SC_LP__MUX4_1%A2 N_A2_M1025_g N_A2_M1015_g N_A2_c_617_n
+ N_A2_c_622_n A2 A2 N_A2_c_619_n PM_SKY130_FD_SC_LP__MUX4_1%A2
x_PM_SKY130_FD_SC_LP__MUX4_1%S1 N_S1_M1004_g N_S1_M1010_g N_S1_c_662_n
+ N_S1_c_663_n N_S1_M1001_g N_S1_M1017_g N_S1_c_665_n N_S1_c_670_n N_S1_c_666_n
+ S1 N_S1_c_667_n N_S1_c_673_p PM_SKY130_FD_SC_LP__MUX4_1%S1
x_PM_SKY130_FD_SC_LP__MUX4_1%A_1245_21# N_A_1245_21#_M1004_d
+ N_A_1245_21#_M1010_d N_A_1245_21#_c_744_n N_A_1245_21#_c_730_n
+ N_A_1245_21#_c_731_n N_A_1245_21#_c_745_n N_A_1245_21#_c_746_n
+ N_A_1245_21#_c_732_n N_A_1245_21#_M1006_g N_A_1245_21#_M1022_g
+ N_A_1245_21#_c_734_n N_A_1245_21#_c_735_n N_A_1245_21#_c_736_n
+ N_A_1245_21#_c_737_n N_A_1245_21#_c_738_n N_A_1245_21#_c_739_n
+ N_A_1245_21#_c_757_n N_A_1245_21#_c_740_n N_A_1245_21#_c_741_n
+ N_A_1245_21#_c_742_n N_A_1245_21#_c_749_n N_A_1245_21#_c_743_n
+ N_A_1245_21#_c_750_n N_A_1245_21#_c_751_n N_A_1245_21#_c_752_n
+ PM_SKY130_FD_SC_LP__MUX4_1%A_1245_21#
x_PM_SKY130_FD_SC_LP__MUX4_1%A_1635_149# N_A_1635_149#_M1001_d
+ N_A_1635_149#_M1017_d N_A_1635_149#_M1020_g N_A_1635_149#_M1002_g
+ N_A_1635_149#_c_860_n N_A_1635_149#_c_866_n N_A_1635_149#_c_861_n
+ N_A_1635_149#_c_862_n N_A_1635_149#_c_863_n N_A_1635_149#_c_864_n
+ PM_SKY130_FD_SC_LP__MUX4_1%A_1635_149#
x_PM_SKY130_FD_SC_LP__MUX4_1%A_27_519# N_A_27_519#_M1000_s N_A_27_519#_M1005_s
+ N_A_27_519#_c_902_n N_A_27_519#_c_903_n N_A_27_519#_c_904_n
+ N_A_27_519#_c_905_n PM_SKY130_FD_SC_LP__MUX4_1%A_27_519#
x_PM_SKY130_FD_SC_LP__MUX4_1%VPWR N_VPWR_M1000_d N_VPWR_M1021_d N_VPWR_M1019_d
+ N_VPWR_M1010_s N_VPWR_M1002_s N_VPWR_c_924_n N_VPWR_c_925_n N_VPWR_c_926_n
+ N_VPWR_c_927_n N_VPWR_c_928_n N_VPWR_c_929_n VPWR N_VPWR_c_930_n
+ N_VPWR_c_931_n N_VPWR_c_932_n N_VPWR_c_933_n N_VPWR_c_934_n N_VPWR_c_923_n
+ N_VPWR_c_936_n N_VPWR_c_937_n N_VPWR_c_938_n N_VPWR_c_939_n N_VPWR_c_940_n
+ PM_SKY130_FD_SC_LP__MUX4_1%VPWR
x_PM_SKY130_FD_SC_LP__MUX4_1%A_196_519# N_A_196_519#_M1013_d
+ N_A_196_519#_M1023_d N_A_196_519#_c_1021_n N_A_196_519#_c_1022_n
+ N_A_196_519#_c_1023_n PM_SKY130_FD_SC_LP__MUX4_1%A_196_519#
x_PM_SKY130_FD_SC_LP__MUX4_1%A_284_81# N_A_284_81#_M1009_d N_A_284_81#_M1006_d
+ N_A_284_81#_M1005_d N_A_284_81#_M1017_s N_A_284_81#_c_1044_n
+ N_A_284_81#_c_1063_n N_A_284_81#_c_1045_n N_A_284_81#_c_1046_n
+ N_A_284_81#_c_1047_n N_A_284_81#_c_1048_n N_A_284_81#_c_1051_n
+ N_A_284_81#_c_1052_n N_A_284_81#_c_1053_n N_A_284_81#_c_1115_n
+ N_A_284_81#_c_1116_n N_A_284_81#_c_1049_n N_A_284_81#_c_1050_n
+ PM_SKY130_FD_SC_LP__MUX4_1%A_284_81#
x_PM_SKY130_FD_SC_LP__MUX4_1%A_799_501# N_A_799_501#_M1003_s
+ N_A_799_501#_M1025_d N_A_799_501#_c_1179_n N_A_799_501#_c_1180_n
+ N_A_799_501#_c_1181_n N_A_799_501#_c_1182_n N_A_799_501#_c_1183_n
+ N_A_799_501#_c_1184_n N_A_799_501#_c_1185_n
+ PM_SKY130_FD_SC_LP__MUX4_1%A_799_501#
x_PM_SKY130_FD_SC_LP__MUX4_1%A_793_117# N_A_793_117#_M1016_d
+ N_A_793_117#_M1001_s N_A_793_117#_M1003_d N_A_793_117#_M1022_d
+ N_A_793_117#_c_1243_n N_A_793_117#_c_1226_n N_A_793_117#_c_1227_n
+ N_A_793_117#_c_1228_n N_A_793_117#_c_1232_n N_A_793_117#_c_1233_n
+ N_A_793_117#_c_1234_n N_A_793_117#_c_1229_n N_A_793_117#_c_1236_n
+ N_A_793_117#_c_1237_n N_A_793_117#_c_1238_n N_A_793_117#_c_1239_n
+ N_A_793_117#_c_1256_n N_A_793_117#_c_1240_n N_A_793_117#_c_1241_n
+ N_A_793_117#_c_1230_n N_A_793_117#_c_1242_n
+ PM_SKY130_FD_SC_LP__MUX4_1%A_793_117#
x_PM_SKY130_FD_SC_LP__MUX4_1%X N_X_M1020_d N_X_M1002_d X X X X X X X
+ PM_SKY130_FD_SC_LP__MUX4_1%X
x_PM_SKY130_FD_SC_LP__MUX4_1%A_33_81# N_A_33_81#_M1014_s N_A_33_81#_M1018_d
+ N_A_33_81#_c_1372_n N_A_33_81#_c_1373_n N_A_33_81#_c_1374_n
+ N_A_33_81#_c_1383_n N_A_33_81#_c_1375_n N_A_33_81#_c_1376_n
+ N_A_33_81#_c_1377_n PM_SKY130_FD_SC_LP__MUX4_1%A_33_81#
x_PM_SKY130_FD_SC_LP__MUX4_1%VGND N_VGND_M1014_d N_VGND_M1011_d N_VGND_M1012_d
+ N_VGND_M1004_s N_VGND_M1020_s N_VGND_c_1416_n N_VGND_c_1417_n N_VGND_c_1418_n
+ N_VGND_c_1419_n N_VGND_c_1420_n N_VGND_c_1421_n N_VGND_c_1422_n VGND
+ N_VGND_c_1423_n N_VGND_c_1424_n N_VGND_c_1425_n N_VGND_c_1426_n
+ N_VGND_c_1427_n N_VGND_c_1428_n N_VGND_c_1429_n N_VGND_c_1430_n
+ N_VGND_c_1431_n N_VGND_c_1432_n PM_SKY130_FD_SC_LP__MUX4_1%VGND
x_PM_SKY130_FD_SC_LP__MUX4_1%A_710_117# N_A_710_117#_M1016_s
+ N_A_710_117#_M1012_s N_A_710_117#_c_1520_n N_A_710_117#_c_1521_n
+ N_A_710_117#_c_1522_n N_A_710_117#_c_1523_n
+ PM_SKY130_FD_SC_LP__MUX4_1%A_710_117#
x_PM_SKY130_FD_SC_LP__MUX4_1%A_879_117# N_A_879_117#_M1007_d
+ N_A_879_117#_M1015_d N_A_879_117#_c_1546_n N_A_879_117#_c_1547_n
+ N_A_879_117#_c_1548_n PM_SKY130_FD_SC_LP__MUX4_1%A_879_117#
cc_1 VNB N_A1_c_219_n 0.0230424f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.7
cc_2 VNB N_A1_M1014_g 0.0415114f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.615
cc_3 VNB A1 0.0238805f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_222_n 0.0218472f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_5 VNB N_A0_M1008_g 0.0469803f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.21
cc_6 VNB A0 0.011364f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A0_c_257_n 0.0104186f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_8 VNB N_A_254_55#_M1009_g 0.0295538f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.615
cc_9 VNB N_A_254_55#_c_301_n 0.0298594f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.88
cc_10 VNB N_A_254_55#_c_302_n 0.00819143f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A_254_55#_M1005_g 0.0179225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_254_55#_c_304_n 0.0131286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_254_55#_M1007_g 0.0361936f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.375
cc_14 VNB N_A_254_55#_c_306_n 0.00580412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_254_55#_c_307_n 0.0121968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_254_55#_c_308_n 0.00103372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_254_55#_c_309_n 0.0409604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_254_55#_c_310_n 0.0183133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_254_55#_c_311_n 0.0459148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_S0_M1018_g 0.0186717f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.88
cc_21 VNB N_S0_c_451_n 0.165287f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.805
cc_22 VNB N_S0_c_452_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_S0_c_453_n 0.0210117f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_24 VNB N_S0_c_454_n 0.019237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_S0_c_455_n 0.0211934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_S0_M1016_g 0.0250414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_S0_c_457_n 0.00576509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_S0_c_458_n 0.0366418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_S0_c_459_n 0.00193429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_S0_c_460_n 0.0260831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A3_c_562_n 0.0122753f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.88
cc_32 VNB N_A3_c_563_n 0.022675f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_33 VNB N_A3_c_564_n 0.00440602f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_34 VNB N_A3_c_565_n 0.0206271f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_35 VNB N_A3_c_566_n 0.0145484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A3_c_567_n 0.0179616f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.21
cc_37 VNB N_A3_c_568_n 0.00612591f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_38 VNB N_A2_M1015_g 0.0398587f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.21
cc_39 VNB N_A2_c_617_n 0.0225311f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.88
cc_40 VNB A2 0.00454201f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_41 VNB N_A2_c_619_n 0.0168097f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.375
cc_42 VNB N_S1_M1004_g 0.028548f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.88
cc_43 VNB N_S1_c_662_n 0.0647667f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.615
cc_44 VNB N_S1_c_663_n 0.0174201f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.88
cc_45 VNB N_S1_M1017_g 0.0145132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_S1_c_665_n 0.0102428f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_47 VNB N_S1_c_666_n 0.00534064f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_48 VNB N_S1_c_667_n 0.0181719f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_49 VNB N_A_1245_21#_c_730_n 0.205408f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.88
cc_50 VNB N_A_1245_21#_c_731_n 0.0101178f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_51 VNB N_A_1245_21#_c_732_n 0.0176952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1245_21#_M1022_g 0.0121546f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.375
cc_53 VNB N_A_1245_21#_c_734_n 0.0278393f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_54 VNB N_A_1245_21#_c_735_n 0.0586656f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.375
cc_55 VNB N_A_1245_21#_c_736_n 0.0517797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1245_21#_c_737_n 0.025269f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=2.035
cc_57 VNB N_A_1245_21#_c_738_n 0.0018683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1245_21#_c_739_n 0.00481183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1245_21#_c_740_n 0.0167672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1245_21#_c_741_n 0.017278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1245_21#_c_742_n 0.00735904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1245_21#_c_743_n 0.00547222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1635_149#_c_860_n 0.00300439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1635_149#_c_861_n 0.00657903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1635_149#_c_862_n 0.0312684f $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.375
cc_66 VNB N_A_1635_149#_c_863_n 0.00235884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1635_149#_c_864_n 0.0206946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VPWR_c_923_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_284_81#_c_1044_n 0.00645808f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_70 VNB N_A_284_81#_c_1045_n 0.0134015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_284_81#_c_1046_n 0.0106266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_284_81#_c_1047_n 0.00605847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_284_81#_c_1048_n 0.00328112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_284_81#_c_1049_n 0.00611023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_284_81#_c_1050_n 0.0061322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_793_117#_c_1226_n 0.00914154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_793_117#_c_1227_n 0.0102848f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.375
cc_78 VNB N_A_793_117#_c_1228_n 0.00463359f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.375
cc_79 VNB N_A_793_117#_c_1229_n 0.0066642f $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=2.035
cc_80 VNB N_A_793_117#_c_1230_n 0.00358286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB X 0.0576438f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.21
cc_82 VNB N_A_33_81#_c_1372_n 0.0140933f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.615
cc_83 VNB N_A_33_81#_c_1373_n 0.0118732f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.88
cc_84 VNB N_A_33_81#_c_1374_n 0.00958375f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_85 VNB N_A_33_81#_c_1375_n 0.00415427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_33_81#_c_1376_n 0.00135468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_33_81#_c_1377_n 0.0142347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1416_n 0.00822758f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.375
cc_89 VNB N_VGND_c_1417_n 0.0152212f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_90 VNB N_VGND_c_1418_n 0.00283848f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_91 VNB N_VGND_c_1419_n 0.0140823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1420_n 0.0151332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1421_n 0.0191722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1422_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1423_n 0.0181485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1424_n 0.0539614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1425_n 0.0477026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1426_n 0.0668973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1427_n 0.0168564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1428_n 0.502866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1429_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1430_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1431_n 0.00515773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1432_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_710_117#_c_1520_n 0.00657455f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=0.615
cc_106 VNB N_A_710_117#_c_1521_n 0.00273273f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_107 VNB N_A_710_117#_c_1522_n 0.00161387f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_108 VNB N_A_710_117#_c_1523_n 0.0211055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_879_117#_c_1546_n 0.030822f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.21
cc_110 VNB N_A_879_117#_c_1547_n 0.00352702f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.88
cc_111 VNB N_A_879_117#_c_1548_n 0.00135821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VPB N_A1_c_219_n 0.00374385f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.7
cc_113 VPB N_A1_M1000_g 0.061061f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.805
cc_114 VPB N_A1_c_225_n 0.0214234f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.88
cc_115 VPB A1 0.024006f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_116 VPB N_A0_M1013_g 0.0357365f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.88
cc_117 VPB N_A0_c_259_n 0.0258817f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.88
cc_118 VPB N_A0_c_260_n 0.0178713f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_119 VPB A0 0.00961334f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_120 VPB N_A0_c_257_n 0.00720605f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.375
cc_121 VPB N_A_254_55#_M1005_g 0.0537339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_254_55#_c_313_n 0.0573496f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.295
cc_123 VPB N_A_254_55#_M1024_g 0.0273974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_254_55#_c_315_n 0.00481843f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_254_55#_c_316_n 0.0107321f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_254_55#_c_317_n 0.0178257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_254_55#_c_318_n 0.0015284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_254_55#_c_309_n 6.93452e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_254_55#_c_310_n 0.00371999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_254_55#_c_311_n 0.0126477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_S0_c_461_n 0.0173547f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.21
cc_132 VPB N_S0_c_462_n 0.0350551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_S0_c_463_n 0.0062736f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.88
cc_134 VPB N_S0_c_454_n 0.0211875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_S0_c_465_n 0.0186473f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.375
cc_136 VPB N_S0_M1021_g 0.0299699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_S0_c_467_n 0.0261228f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_138 VPB N_S0_c_468_n 0.0448278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_S0_c_469_n 0.0111315f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=2.035
cc_140 VPB N_S0_c_470_n 0.020683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_S0_c_471_n 0.00723013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_S0_c_459_n 0.0155186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_S0_c_473_n 0.00230021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A3_M1019_g 0.0469788f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.88
cc_145 VPB N_A3_c_564_n 0.0109439f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_146 VPB N_A3_c_568_n 0.00179458f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.295
cc_147 VPB N_A2_M1025_g 0.0518176f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.88
cc_148 VPB N_A2_c_617_n 6.16351e-19 $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.88
cc_149 VPB N_A2_c_622_n 0.016628f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_150 VPB A2 0.00180465f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_151 VPB N_S1_M1010_g 0.0292243f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.21
cc_152 VPB N_S1_M1017_g 0.0234575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_S1_c_670_n 0.0186067f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.21
cc_154 VPB N_S1_c_667_n 0.00984191f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_155 VPB N_A_1245_21#_c_744_n 0.075989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_1245_21#_c_745_n 0.0658518f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_157 VPB N_A_1245_21#_c_746_n 0.0123046f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_158 VPB N_A_1245_21#_M1022_g 0.0255239f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.375
cc_159 VPB N_A_1245_21#_c_738_n 0.0150435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_1245_21#_c_749_n 0.00923287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_1245_21#_c_750_n 0.00154748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_1245_21#_c_751_n 0.0130191f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_1245_21#_c_752_n 0.0490604f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_1635_149#_M1002_g 0.0284848f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_165 VPB N_A_1635_149#_c_866_n 0.00265899f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.375
cc_166 VPB N_A_1635_149#_c_861_n 0.0179384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_1635_149#_c_862_n 0.00714818f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.375
cc_168 VPB N_A_1635_149#_c_863_n 3.55821e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_27_519#_c_902_n 0.0184203f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.615
cc_170 VPB N_A_27_519#_c_903_n 0.024448f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.88
cc_171 VPB N_A_27_519#_c_904_n 0.00983105f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_172 VPB N_A_27_519#_c_905_n 0.0048195f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_173 VPB N_VPWR_c_924_n 0.00254872f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.375
cc_174 VPB N_VPWR_c_925_n 0.0182982f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.295
cc_175 VPB N_VPWR_c_926_n 0.00990536f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_176 VPB N_VPWR_c_927_n 0.0254135f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=2.035
cc_177 VPB N_VPWR_c_928_n 0.0127605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_929_n 0.031411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_930_n 0.0163534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_931_n 0.0626318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_932_n 0.0412183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_933_n 0.0665837f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_934_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_923_n 0.150767f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_936_n 0.00534513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_937_n 0.00574453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_938_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_939_n 0.00563364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_940_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_196_519#_c_1021_n 0.0356347f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.21
cc_191 VPB N_A_196_519#_c_1022_n 0.00774918f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.88
cc_192 VPB N_A_196_519#_c_1023_n 0.00651684f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_193 VPB N_A_284_81#_c_1051_n 0.0614623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_284_81#_c_1052_n 0.00547051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_284_81#_c_1053_n 0.00308231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_284_81#_c_1049_n 0.00317872f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_284_81#_c_1050_n 0.00199603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_799_501#_c_1179_n 0.00417365f $X=-0.19 $Y=1.655 $X2=0.505
+ $Y2=0.615
cc_199 VPB N_A_799_501#_c_1180_n 0.00667271f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.88
cc_200 VPB N_A_799_501#_c_1181_n 0.00427344f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.21
cc_201 VPB N_A_799_501#_c_1182_n 3.4571e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_202 VPB N_A_799_501#_c_1183_n 0.0127213f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_799_501#_c_1184_n 0.00169815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_799_501#_c_1185_n 0.00533818f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.375
cc_205 VPB N_A_793_117#_c_1228_n 0.00243788f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.375
cc_206 VPB N_A_793_117#_c_1232_n 0.00633292f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.295
cc_207 VPB N_A_793_117#_c_1233_n 0.0337521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_793_117#_c_1234_n 0.0168043f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.375
cc_209 VPB N_A_793_117#_c_1229_n 0.00862127f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=2.035
cc_210 VPB N_A_793_117#_c_1236_n 0.00523761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_793_117#_c_1237_n 0.0323783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_793_117#_c_1238_n 0.00404339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_793_117#_c_1239_n 0.00274232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_793_117#_c_1240_n 2.3787e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_793_117#_c_1241_n 0.00726622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_793_117#_c_1242_n 0.00197718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB X 0.057609f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.21
cc_218 N_A1_M1014_g N_A0_M1008_g 0.0358823f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_219 A1 N_A0_M1008_g 5.62311e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A1_M1000_g N_A0_c_259_n 0.0393416f $X=0.475 $Y=2.805 $X2=0 $Y2=0
cc_221 N_A1_c_225_n N_A0_c_259_n 0.00733406f $X=0.4 $Y=1.88 $X2=0 $Y2=0
cc_222 N_A1_c_219_n A0 0.0011345f $X=0.4 $Y=1.7 $X2=0 $Y2=0
cc_223 N_A1_M1000_g A0 9.83175e-19 $X=0.475 $Y=2.805 $X2=0 $Y2=0
cc_224 N_A1_M1014_g A0 0.00326057f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_225 A1 A0 0.0560031f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_226 N_A1_c_219_n N_A0_c_257_n 0.00733406f $X=0.4 $Y=1.7 $X2=0 $Y2=0
cc_227 A1 N_A0_c_257_n 0.00218958f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_228 N_A1_M1000_g N_A_27_519#_c_902_n 0.00354946f $X=0.475 $Y=2.805 $X2=0
+ $Y2=0
cc_229 N_A1_M1000_g N_A_27_519#_c_903_n 0.0129354f $X=0.475 $Y=2.805 $X2=0 $Y2=0
cc_230 N_A1_c_225_n N_A_27_519#_c_903_n 0.00107561f $X=0.4 $Y=1.88 $X2=0 $Y2=0
cc_231 A1 N_A_27_519#_c_903_n 0.015113f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_232 N_A1_c_225_n N_A_27_519#_c_904_n 5.51034e-19 $X=0.4 $Y=1.88 $X2=0 $Y2=0
cc_233 A1 N_A_27_519#_c_904_n 0.0242089f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_234 N_A1_M1000_g N_VPWR_c_924_n 0.0118175f $X=0.475 $Y=2.805 $X2=0 $Y2=0
cc_235 N_A1_M1000_g N_VPWR_c_930_n 0.00422142f $X=0.475 $Y=2.805 $X2=0 $Y2=0
cc_236 N_A1_M1000_g N_VPWR_c_923_n 0.00458201f $X=0.475 $Y=2.805 $X2=0 $Y2=0
cc_237 N_A1_M1014_g N_A_33_81#_c_1373_n 0.0141489f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_238 A1 N_A_33_81#_c_1373_n 0.0128273f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_239 N_A1_c_222_n N_A_33_81#_c_1373_n 2.67499e-19 $X=0.385 $Y=1.375 $X2=0
+ $Y2=0
cc_240 A1 N_A_33_81#_c_1374_n 0.0239312f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_241 N_A1_c_222_n N_A_33_81#_c_1374_n 0.00108709f $X=0.385 $Y=1.375 $X2=0
+ $Y2=0
cc_242 N_A1_M1014_g N_A_33_81#_c_1383_n 3.36945e-19 $X=0.505 $Y=0.615 $X2=0
+ $Y2=0
cc_243 N_A1_M1014_g N_VGND_c_1416_n 0.012006f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_244 N_A1_M1014_g N_VGND_c_1423_n 0.0045897f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_245 N_A1_M1014_g N_VGND_c_1428_n 0.0044912f $X=0.505 $Y=0.615 $X2=0 $Y2=0
cc_246 N_A0_M1008_g N_A_254_55#_M1009_g 0.0657f $X=0.985 $Y=0.615 $X2=0 $Y2=0
cc_247 A0 N_A_254_55#_M1009_g 0.00760203f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_248 A0 N_A_254_55#_c_301_n 0.00520956f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_249 A0 N_A_254_55#_c_302_n 0.00726614f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_250 N_A0_M1008_g N_A_254_55#_M1005_g 0.00216684f $X=0.985 $Y=0.615 $X2=0
+ $Y2=0
cc_251 A0 N_A_254_55#_M1005_g 0.00857487f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_252 N_A0_c_257_n N_A_254_55#_M1005_g 0.00930365f $X=0.995 $Y=1.75 $X2=0 $Y2=0
cc_253 N_A0_M1013_g N_A_27_519#_c_903_n 0.013331f $X=0.905 $Y=2.805 $X2=0 $Y2=0
cc_254 N_A0_c_260_n N_A_27_519#_c_903_n 0.00516471f $X=0.995 $Y=2.255 $X2=0
+ $Y2=0
cc_255 A0 N_A_27_519#_c_903_n 0.0501427f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_256 N_A0_M1013_g N_A_27_519#_c_905_n 0.00427872f $X=0.905 $Y=2.805 $X2=0
+ $Y2=0
cc_257 N_A0_M1013_g N_VPWR_c_924_n 0.00968429f $X=0.905 $Y=2.805 $X2=0 $Y2=0
cc_258 N_A0_M1013_g N_VPWR_c_931_n 0.00422142f $X=0.905 $Y=2.805 $X2=0 $Y2=0
cc_259 N_A0_M1013_g N_VPWR_c_923_n 0.00475143f $X=0.905 $Y=2.805 $X2=0 $Y2=0
cc_260 N_A0_M1013_g N_A_196_519#_c_1023_n 4.46816e-19 $X=0.905 $Y=2.805 $X2=0
+ $Y2=0
cc_261 N_A0_M1008_g N_A_284_81#_c_1048_n 3.85956e-19 $X=0.985 $Y=0.615 $X2=0
+ $Y2=0
cc_262 A0 N_A_284_81#_c_1048_n 0.00455704f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_263 A0 N_A_284_81#_c_1052_n 0.00150746f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_264 A0 N_A_284_81#_c_1049_n 0.0364488f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_265 N_A0_M1008_g N_A_33_81#_c_1373_n 0.011003f $X=0.985 $Y=0.615 $X2=0 $Y2=0
cc_266 A0 N_A_33_81#_c_1373_n 0.0309681f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_267 N_A0_c_257_n N_A_33_81#_c_1373_n 5.81761e-19 $X=0.995 $Y=1.75 $X2=0 $Y2=0
cc_268 N_A0_M1008_g N_A_33_81#_c_1383_n 0.00726643f $X=0.985 $Y=0.615 $X2=0
+ $Y2=0
cc_269 N_A0_M1008_g N_A_33_81#_c_1376_n 0.00293487f $X=0.985 $Y=0.615 $X2=0
+ $Y2=0
cc_270 N_A0_M1008_g N_VGND_c_1416_n 0.00111447f $X=0.985 $Y=0.615 $X2=0 $Y2=0
cc_271 N_A0_M1008_g N_VGND_c_1424_n 0.00537026f $X=0.985 $Y=0.615 $X2=0 $Y2=0
cc_272 N_A0_M1008_g N_VGND_c_1428_n 0.00516844f $X=0.985 $Y=0.615 $X2=0 $Y2=0
cc_273 N_A_254_55#_M1009_g N_S0_M1018_g 0.0159778f $X=1.345 $Y=0.615 $X2=0 $Y2=0
cc_274 N_A_254_55#_c_301_n N_S0_M1018_g 0.00795185f $X=1.78 $Y=1.27 $X2=0 $Y2=0
cc_275 N_A_254_55#_c_307_n N_S0_c_451_n 0.00491825f $X=2.725 $Y=0.805 $X2=0
+ $Y2=0
cc_276 N_A_254_55#_c_316_n N_S0_c_461_n 0.00293965f $X=3.05 $Y=2.68 $X2=0 $Y2=0
cc_277 N_A_254_55#_c_315_n N_S0_c_462_n 0.00145489f $X=2.735 $Y=1.975 $X2=0
+ $Y2=0
cc_278 N_A_254_55#_c_318_n N_S0_c_462_n 0.0147239f $X=3.175 $Y=2.06 $X2=0 $Y2=0
cc_279 N_A_254_55#_c_310_n N_S0_c_462_n 0.00271358f $X=2.34 $Y=1.265 $X2=0 $Y2=0
cc_280 N_A_254_55#_M1005_g N_S0_c_463_n 0.0191335f $X=1.855 $Y=2.505 $X2=0 $Y2=0
cc_281 N_A_254_55#_c_310_n N_S0_c_463_n 0.00100277f $X=2.34 $Y=1.265 $X2=0 $Y2=0
cc_282 N_A_254_55#_c_311_n N_S0_c_463_n 0.0150626f $X=2.34 $Y=1.265 $X2=0 $Y2=0
cc_283 N_A_254_55#_c_307_n N_S0_c_453_n 0.0062427f $X=2.725 $Y=0.805 $X2=0 $Y2=0
cc_284 N_A_254_55#_c_311_n N_S0_c_453_n 0.00985214f $X=2.34 $Y=1.265 $X2=0 $Y2=0
cc_285 N_A_254_55#_c_315_n N_S0_c_454_n 0.0062427f $X=2.735 $Y=1.975 $X2=0 $Y2=0
cc_286 N_A_254_55#_c_318_n N_S0_c_454_n 0.00510872f $X=3.175 $Y=2.06 $X2=0 $Y2=0
cc_287 N_A_254_55#_c_316_n N_S0_c_465_n 0.00370529f $X=3.05 $Y=2.68 $X2=0 $Y2=0
cc_288 N_A_254_55#_c_317_n N_S0_c_465_n 0.0125017f $X=4.175 $Y=2.06 $X2=0 $Y2=0
cc_289 N_A_254_55#_c_318_n N_S0_c_465_n 0.0045553f $X=3.175 $Y=2.06 $X2=0 $Y2=0
cc_290 N_A_254_55#_c_316_n N_S0_M1021_g 0.0125838f $X=3.05 $Y=2.68 $X2=0 $Y2=0
cc_291 N_A_254_55#_c_316_n N_S0_c_467_n 2.08187e-19 $X=3.05 $Y=2.68 $X2=0 $Y2=0
cc_292 N_A_254_55#_c_317_n N_S0_c_467_n 0.0154194f $X=4.175 $Y=2.06 $X2=0 $Y2=0
cc_293 N_A_254_55#_c_313_n N_S0_c_468_n 0.0148643f $X=4.472 $Y=1.99 $X2=0 $Y2=0
cc_294 N_A_254_55#_M1024_g N_S0_c_468_n 0.0214622f $X=4.765 $Y=2.715 $X2=0 $Y2=0
cc_295 N_A_254_55#_c_317_n N_S0_c_468_n 0.0195031f $X=4.175 $Y=2.06 $X2=0 $Y2=0
cc_296 N_A_254_55#_M1007_g N_S0_M1016_g 0.0194434f $X=4.32 $Y=0.795 $X2=0 $Y2=0
cc_297 N_A_254_55#_c_310_n N_S0_c_457_n 0.0062427f $X=2.34 $Y=1.265 $X2=0 $Y2=0
cc_298 N_A_254_55#_c_311_n N_S0_c_457_n 0.00985214f $X=2.34 $Y=1.265 $X2=0 $Y2=0
cc_299 N_A_254_55#_c_316_n N_S0_c_471_n 0.00504898f $X=3.05 $Y=2.68 $X2=0 $Y2=0
cc_300 N_A_254_55#_c_318_n N_S0_c_471_n 0.00272314f $X=3.175 $Y=2.06 $X2=0 $Y2=0
cc_301 N_A_254_55#_c_313_n N_S0_c_459_n 0.00914152f $X=4.472 $Y=1.99 $X2=0 $Y2=0
cc_302 N_A_254_55#_c_317_n N_S0_c_459_n 0.00455213f $X=4.175 $Y=2.06 $X2=0 $Y2=0
cc_303 N_A_254_55#_c_308_n N_S0_c_460_n 0.00288626f $X=4.34 $Y=1.53 $X2=0 $Y2=0
cc_304 N_A_254_55#_c_309_n N_S0_c_460_n 0.00914152f $X=4.34 $Y=1.53 $X2=0 $Y2=0
cc_305 N_A_254_55#_M1007_g N_S0_c_473_n 0.00148858f $X=4.32 $Y=0.795 $X2=0 $Y2=0
cc_306 N_A_254_55#_c_318_n N_S0_c_473_n 0.0439658f $X=3.175 $Y=2.06 $X2=0 $Y2=0
cc_307 N_A_254_55#_c_308_n N_S0_c_473_n 0.0132754f $X=4.34 $Y=1.53 $X2=0 $Y2=0
cc_308 N_A_254_55#_c_309_n N_S0_c_473_n 0.00180911f $X=4.34 $Y=1.53 $X2=0 $Y2=0
cc_309 N_A_254_55#_c_310_n N_S0_c_473_n 0.0580212f $X=2.34 $Y=1.265 $X2=0 $Y2=0
cc_310 N_A_254_55#_c_311_n N_S0_c_473_n 4.3714e-19 $X=2.34 $Y=1.265 $X2=0 $Y2=0
cc_311 N_A_254_55#_c_313_n N_A3_M1019_g 0.074468f $X=4.472 $Y=1.99 $X2=0 $Y2=0
cc_312 N_A_254_55#_c_309_n N_A3_c_563_n 0.0124961f $X=4.34 $Y=1.53 $X2=0 $Y2=0
cc_313 N_A_254_55#_c_313_n N_A3_c_564_n 0.0124961f $X=4.472 $Y=1.99 $X2=0 $Y2=0
cc_314 N_A_254_55#_M1007_g N_A3_c_567_n 0.00385617f $X=4.32 $Y=0.795 $X2=0 $Y2=0
cc_315 N_A_254_55#_M1007_g N_A3_c_568_n 4.17491e-19 $X=4.32 $Y=0.795 $X2=0 $Y2=0
cc_316 N_A_254_55#_c_309_n N_A3_c_568_n 0.00126698f $X=4.34 $Y=1.53 $X2=0 $Y2=0
cc_317 N_A_254_55#_c_317_n N_VPWR_c_925_n 0.0104895f $X=4.175 $Y=2.06 $X2=0
+ $Y2=0
cc_318 N_A_254_55#_c_316_n N_VPWR_c_931_n 0.00751229f $X=3.05 $Y=2.68 $X2=0
+ $Y2=0
cc_319 N_A_254_55#_M1024_g N_VPWR_c_932_n 9.15902e-19 $X=4.765 $Y=2.715 $X2=0
+ $Y2=0
cc_320 N_A_254_55#_c_316_n N_VPWR_c_923_n 0.00974862f $X=3.05 $Y=2.68 $X2=0
+ $Y2=0
cc_321 N_A_254_55#_M1005_g N_A_196_519#_c_1021_n 0.00692651f $X=1.855 $Y=2.505
+ $X2=0 $Y2=0
cc_322 N_A_254_55#_c_316_n N_A_196_519#_c_1022_n 0.0341482f $X=3.05 $Y=2.68
+ $X2=0 $Y2=0
cc_323 N_A_254_55#_c_318_n N_A_196_519#_c_1022_n 8.92347e-19 $X=3.175 $Y=2.06
+ $X2=0 $Y2=0
cc_324 N_A_254_55#_c_310_n N_A_196_519#_c_1022_n 0.00356589f $X=2.34 $Y=1.265
+ $X2=0 $Y2=0
cc_325 N_A_254_55#_M1005_g N_A_196_519#_c_1023_n 0.00385782f $X=1.855 $Y=2.505
+ $X2=0 $Y2=0
cc_326 N_A_254_55#_M1009_g N_A_284_81#_c_1044_n 2.41076e-19 $X=1.345 $Y=0.615
+ $X2=0 $Y2=0
cc_327 N_A_254_55#_c_301_n N_A_284_81#_c_1044_n 0.00476906f $X=1.78 $Y=1.27
+ $X2=0 $Y2=0
cc_328 N_A_254_55#_c_307_n N_A_284_81#_c_1044_n 0.00678258f $X=2.725 $Y=0.805
+ $X2=0 $Y2=0
cc_329 N_A_254_55#_M1005_g N_A_284_81#_c_1063_n 0.0126989f $X=1.855 $Y=2.505
+ $X2=0 $Y2=0
cc_330 N_A_254_55#_c_316_n N_A_284_81#_c_1063_n 0.00471989f $X=3.05 $Y=2.68
+ $X2=0 $Y2=0
cc_331 N_A_254_55#_M1009_g N_A_284_81#_c_1048_n 0.00721333f $X=1.345 $Y=0.615
+ $X2=0 $Y2=0
cc_332 N_A_254_55#_c_301_n N_A_284_81#_c_1048_n 0.0100875f $X=1.78 $Y=1.27 $X2=0
+ $Y2=0
cc_333 N_A_254_55#_c_313_n N_A_284_81#_c_1051_n 0.0113502f $X=4.472 $Y=1.99
+ $X2=0 $Y2=0
cc_334 N_A_254_55#_c_315_n N_A_284_81#_c_1051_n 0.00967835f $X=2.735 $Y=1.975
+ $X2=0 $Y2=0
cc_335 N_A_254_55#_c_316_n N_A_284_81#_c_1051_n 0.00350532f $X=3.05 $Y=2.68
+ $X2=0 $Y2=0
cc_336 N_A_254_55#_c_317_n N_A_284_81#_c_1051_n 0.0572963f $X=4.175 $Y=2.06
+ $X2=0 $Y2=0
cc_337 N_A_254_55#_c_318_n N_A_284_81#_c_1051_n 0.0251261f $X=3.175 $Y=2.06
+ $X2=0 $Y2=0
cc_338 N_A_254_55#_c_308_n N_A_284_81#_c_1051_n 0.0143698f $X=4.34 $Y=1.53 $X2=0
+ $Y2=0
cc_339 N_A_254_55#_c_310_n N_A_284_81#_c_1051_n 0.0124747f $X=2.34 $Y=1.265
+ $X2=0 $Y2=0
cc_340 N_A_254_55#_c_315_n N_A_284_81#_c_1052_n 0.00120021f $X=2.735 $Y=1.975
+ $X2=0 $Y2=0
cc_341 N_A_254_55#_c_318_n N_A_284_81#_c_1052_n 8.71255e-19 $X=3.175 $Y=2.06
+ $X2=0 $Y2=0
cc_342 N_A_254_55#_c_310_n N_A_284_81#_c_1052_n 0.00142058f $X=2.34 $Y=1.265
+ $X2=0 $Y2=0
cc_343 N_A_254_55#_c_311_n N_A_284_81#_c_1052_n 0.00175479f $X=2.34 $Y=1.265
+ $X2=0 $Y2=0
cc_344 N_A_254_55#_M1005_g N_A_284_81#_c_1053_n 0.00770286f $X=1.855 $Y=2.505
+ $X2=0 $Y2=0
cc_345 N_A_254_55#_c_315_n N_A_284_81#_c_1053_n 0.00117599f $X=2.735 $Y=1.975
+ $X2=0 $Y2=0
cc_346 N_A_254_55#_c_316_n N_A_284_81#_c_1053_n 6.16221e-19 $X=3.05 $Y=2.68
+ $X2=0 $Y2=0
cc_347 N_A_254_55#_c_318_n N_A_284_81#_c_1053_n 0.00528212f $X=3.175 $Y=2.06
+ $X2=0 $Y2=0
cc_348 N_A_254_55#_c_310_n N_A_284_81#_c_1053_n 0.00336576f $X=2.34 $Y=1.265
+ $X2=0 $Y2=0
cc_349 N_A_254_55#_c_311_n N_A_284_81#_c_1053_n 0.00244698f $X=2.34 $Y=1.265
+ $X2=0 $Y2=0
cc_350 N_A_254_55#_M1009_g N_A_284_81#_c_1049_n 0.0042738f $X=1.345 $Y=0.615
+ $X2=0 $Y2=0
cc_351 N_A_254_55#_M1005_g N_A_284_81#_c_1049_n 0.01625f $X=1.855 $Y=2.505 $X2=0
+ $Y2=0
cc_352 N_A_254_55#_c_304_n N_A_284_81#_c_1049_n 0.00843661f $X=2.175 $Y=1.27
+ $X2=0 $Y2=0
cc_353 N_A_254_55#_c_306_n N_A_284_81#_c_1049_n 0.00436997f $X=1.855 $Y=1.27
+ $X2=0 $Y2=0
cc_354 N_A_254_55#_c_307_n N_A_284_81#_c_1049_n 0.00354257f $X=2.725 $Y=0.805
+ $X2=0 $Y2=0
cc_355 N_A_254_55#_c_315_n N_A_284_81#_c_1049_n 0.0051568f $X=2.735 $Y=1.975
+ $X2=0 $Y2=0
cc_356 N_A_254_55#_c_310_n N_A_284_81#_c_1049_n 0.0496803f $X=2.34 $Y=1.265
+ $X2=0 $Y2=0
cc_357 N_A_254_55#_c_311_n N_A_284_81#_c_1049_n 0.00518821f $X=2.34 $Y=1.265
+ $X2=0 $Y2=0
cc_358 N_A_254_55#_c_317_n N_A_799_501#_c_1179_n 0.00899061f $X=4.175 $Y=2.06
+ $X2=0 $Y2=0
cc_359 N_A_254_55#_M1024_g N_A_799_501#_c_1180_n 0.0113365f $X=4.765 $Y=2.715
+ $X2=0 $Y2=0
cc_360 N_A_254_55#_M1024_g N_A_799_501#_c_1182_n 0.00524618f $X=4.765 $Y=2.715
+ $X2=0 $Y2=0
cc_361 N_A_254_55#_M1024_g N_A_799_501#_c_1184_n 0.00109046f $X=4.765 $Y=2.715
+ $X2=0 $Y2=0
cc_362 N_A_254_55#_M1007_g N_A_793_117#_c_1243_n 2.98514e-19 $X=4.32 $Y=0.795
+ $X2=0 $Y2=0
cc_363 N_A_254_55#_M1007_g N_A_793_117#_c_1226_n 0.0126624f $X=4.32 $Y=0.795
+ $X2=0 $Y2=0
cc_364 N_A_254_55#_c_308_n N_A_793_117#_c_1226_n 0.0173024f $X=4.34 $Y=1.53
+ $X2=0 $Y2=0
cc_365 N_A_254_55#_c_309_n N_A_793_117#_c_1226_n 0.00751325f $X=4.34 $Y=1.53
+ $X2=0 $Y2=0
cc_366 N_A_254_55#_c_308_n N_A_793_117#_c_1227_n 0.00201896f $X=4.34 $Y=1.53
+ $X2=0 $Y2=0
cc_367 N_A_254_55#_c_313_n N_A_793_117#_c_1228_n 0.00854312f $X=4.472 $Y=1.99
+ $X2=0 $Y2=0
cc_368 N_A_254_55#_M1007_g N_A_793_117#_c_1228_n 0.00400936f $X=4.32 $Y=0.795
+ $X2=0 $Y2=0
cc_369 N_A_254_55#_c_308_n N_A_793_117#_c_1228_n 0.039834f $X=4.34 $Y=1.53 $X2=0
+ $Y2=0
cc_370 N_A_254_55#_c_309_n N_A_793_117#_c_1228_n 0.0124307f $X=4.34 $Y=1.53
+ $X2=0 $Y2=0
cc_371 N_A_254_55#_c_313_n N_A_793_117#_c_1232_n 0.00290642f $X=4.472 $Y=1.99
+ $X2=0 $Y2=0
cc_372 N_A_254_55#_M1024_g N_A_793_117#_c_1232_n 0.00963241f $X=4.765 $Y=2.715
+ $X2=0 $Y2=0
cc_373 N_A_254_55#_c_317_n N_A_793_117#_c_1232_n 0.00333992f $X=4.175 $Y=2.06
+ $X2=0 $Y2=0
cc_374 N_A_254_55#_c_313_n N_A_793_117#_c_1233_n 0.00422861f $X=4.472 $Y=1.99
+ $X2=0 $Y2=0
cc_375 N_A_254_55#_c_313_n N_A_793_117#_c_1256_n 0.00361972f $X=4.472 $Y=1.99
+ $X2=0 $Y2=0
cc_376 N_A_254_55#_M1024_g N_A_793_117#_c_1256_n 0.00431376f $X=4.765 $Y=2.715
+ $X2=0 $Y2=0
cc_377 N_A_254_55#_c_317_n N_A_793_117#_c_1256_n 0.00162135f $X=4.175 $Y=2.06
+ $X2=0 $Y2=0
cc_378 N_A_254_55#_c_313_n N_A_793_117#_c_1240_n 0.00560036f $X=4.472 $Y=1.99
+ $X2=0 $Y2=0
cc_379 N_A_254_55#_c_317_n N_A_793_117#_c_1240_n 0.00921915f $X=4.175 $Y=2.06
+ $X2=0 $Y2=0
cc_380 N_A_254_55#_c_308_n N_A_793_117#_c_1240_n 0.00297955f $X=4.34 $Y=1.53
+ $X2=0 $Y2=0
cc_381 N_A_254_55#_M1009_g N_A_33_81#_c_1373_n 0.00119278f $X=1.345 $Y=0.615
+ $X2=0 $Y2=0
cc_382 N_A_254_55#_M1009_g N_A_33_81#_c_1375_n 0.0135297f $X=1.345 $Y=0.615
+ $X2=0 $Y2=0
cc_383 N_A_254_55#_c_304_n N_A_33_81#_c_1377_n 0.00305881f $X=2.175 $Y=1.27
+ $X2=0 $Y2=0
cc_384 N_A_254_55#_c_306_n N_A_33_81#_c_1377_n 5.88112e-19 $X=1.855 $Y=1.27
+ $X2=0 $Y2=0
cc_385 N_A_254_55#_c_307_n N_A_33_81#_c_1377_n 0.00127885f $X=2.725 $Y=0.805
+ $X2=0 $Y2=0
cc_386 N_A_254_55#_c_311_n N_A_33_81#_c_1377_n 0.00166541f $X=2.34 $Y=1.265
+ $X2=0 $Y2=0
cc_387 N_A_254_55#_M1009_g N_VGND_c_1424_n 9.29198e-19 $X=1.345 $Y=0.615 $X2=0
+ $Y2=0
cc_388 N_A_254_55#_c_307_n N_VGND_c_1424_n 0.00485084f $X=2.725 $Y=0.805 $X2=0
+ $Y2=0
cc_389 N_A_254_55#_c_307_n N_VGND_c_1428_n 0.00678661f $X=2.725 $Y=0.805 $X2=0
+ $Y2=0
cc_390 N_A_254_55#_M1007_g N_A_710_117#_c_1522_n 5.02084e-19 $X=4.32 $Y=0.795
+ $X2=0 $Y2=0
cc_391 N_A_254_55#_M1007_g N_A_710_117#_c_1523_n 0.00549226f $X=4.32 $Y=0.795
+ $X2=0 $Y2=0
cc_392 N_A_254_55#_M1007_g N_A_879_117#_c_1548_n 0.00293961f $X=4.32 $Y=0.795
+ $X2=0 $Y2=0
cc_393 N_A_254_55#_c_309_n N_A_879_117#_c_1548_n 7.58531e-19 $X=4.34 $Y=1.53
+ $X2=0 $Y2=0
cc_394 N_S0_M1021_g N_VPWR_c_925_n 0.00598921f $X=3.265 $Y=2.68 $X2=0 $Y2=0
cc_395 N_S0_c_469_n N_VPWR_c_925_n 0.00206689f $X=3.73 $Y=2.32 $X2=0 $Y2=0
cc_396 N_S0_c_470_n N_VPWR_c_925_n 0.00166852f $X=4.335 $Y=2.395 $X2=0 $Y2=0
cc_397 N_S0_M1021_g N_VPWR_c_931_n 0.00527445f $X=3.265 $Y=2.68 $X2=0 $Y2=0
cc_398 N_S0_c_470_n N_VPWR_c_932_n 9.15902e-19 $X=4.335 $Y=2.395 $X2=0 $Y2=0
cc_399 N_S0_M1021_g N_VPWR_c_923_n 0.00523671f $X=3.265 $Y=2.68 $X2=0 $Y2=0
cc_400 N_S0_c_461_n N_A_196_519#_c_1021_n 0.00692651f $X=2.285 $Y=2.185 $X2=0
+ $Y2=0
cc_401 N_S0_M1021_g N_A_196_519#_c_1021_n 0.00427842f $X=3.265 $Y=2.68 $X2=0
+ $Y2=0
cc_402 N_S0_c_461_n N_A_196_519#_c_1022_n 0.00563562f $X=2.285 $Y=2.185 $X2=0
+ $Y2=0
cc_403 N_S0_c_462_n N_A_196_519#_c_1022_n 0.00551314f $X=2.865 $Y=2.11 $X2=0
+ $Y2=0
cc_404 N_S0_M1018_g N_A_284_81#_c_1044_n 0.00715325f $X=1.775 $Y=0.615 $X2=0
+ $Y2=0
cc_405 N_S0_c_461_n N_A_284_81#_c_1063_n 0.00858916f $X=2.285 $Y=2.185 $X2=0
+ $Y2=0
cc_406 N_S0_c_463_n N_A_284_81#_c_1063_n 6.09752e-19 $X=2.36 $Y=2.11 $X2=0 $Y2=0
cc_407 N_S0_M1018_g N_A_284_81#_c_1048_n 0.010511f $X=1.775 $Y=0.615 $X2=0 $Y2=0
cc_408 N_S0_c_462_n N_A_284_81#_c_1051_n 0.00582099f $X=2.865 $Y=2.11 $X2=0
+ $Y2=0
cc_409 N_S0_c_463_n N_A_284_81#_c_1051_n 0.00225339f $X=2.36 $Y=2.11 $X2=0 $Y2=0
cc_410 N_S0_c_454_n N_A_284_81#_c_1051_n 0.00552643f $X=2.94 $Y=2.035 $X2=0
+ $Y2=0
cc_411 N_S0_c_467_n N_A_284_81#_c_1051_n 0.00418f $X=3.655 $Y=2.245 $X2=0 $Y2=0
cc_412 N_S0_c_459_n N_A_284_81#_c_1051_n 0.00494548f $X=3.565 $Y=1.795 $X2=0
+ $Y2=0
cc_413 N_S0_c_473_n N_A_284_81#_c_1051_n 0.0168815f $X=3.565 $Y=1.29 $X2=0 $Y2=0
cc_414 N_S0_c_463_n N_A_284_81#_c_1052_n 5.37321e-19 $X=2.36 $Y=2.11 $X2=0 $Y2=0
cc_415 N_S0_c_463_n N_A_284_81#_c_1053_n 0.00857702f $X=2.36 $Y=2.11 $X2=0 $Y2=0
cc_416 N_S0_c_454_n N_A_284_81#_c_1053_n 2.61282e-19 $X=2.94 $Y=2.035 $X2=0
+ $Y2=0
cc_417 N_S0_c_468_n N_A_799_501#_c_1179_n 0.005854f $X=4.26 $Y=2.32 $X2=0 $Y2=0
cc_418 N_S0_c_470_n N_A_799_501#_c_1180_n 0.0146835f $X=4.335 $Y=2.395 $X2=0
+ $Y2=0
cc_419 N_S0_M1016_g N_A_793_117#_c_1243_n 3.15041e-19 $X=3.89 $Y=0.795 $X2=0
+ $Y2=0
cc_420 N_S0_M1016_g N_A_793_117#_c_1227_n 0.00472475f $X=3.89 $Y=0.795 $X2=0
+ $Y2=0
cc_421 N_S0_c_473_n N_A_793_117#_c_1227_n 0.00322444f $X=3.565 $Y=1.29 $X2=0
+ $Y2=0
cc_422 N_S0_c_468_n N_A_793_117#_c_1232_n 0.00575527f $X=4.26 $Y=2.32 $X2=0
+ $Y2=0
cc_423 N_S0_c_470_n N_A_793_117#_c_1256_n 0.00360831f $X=4.335 $Y=2.395 $X2=0
+ $Y2=0
cc_424 N_S0_M1018_g N_A_33_81#_c_1375_n 0.0113762f $X=1.775 $Y=0.615 $X2=0 $Y2=0
cc_425 N_S0_M1018_g N_A_33_81#_c_1377_n 0.00165341f $X=1.775 $Y=0.615 $X2=0
+ $Y2=0
cc_426 N_S0_c_451_n N_A_33_81#_c_1377_n 0.00683623f $X=3.815 $Y=0.18 $X2=0 $Y2=0
cc_427 N_S0_c_453_n N_A_33_81#_c_1377_n 0.00373331f $X=2.94 $Y=1.125 $X2=0 $Y2=0
cc_428 N_S0_c_451_n N_VGND_c_1417_n 0.0256263f $X=3.815 $Y=0.18 $X2=0 $Y2=0
cc_429 N_S0_c_453_n N_VGND_c_1417_n 0.0144348f $X=2.94 $Y=1.125 $X2=0 $Y2=0
cc_430 N_S0_c_455_n N_VGND_c_1417_n 0.00433746f $X=3.4 $Y=1.2 $X2=0 $Y2=0
cc_431 N_S0_M1016_g N_VGND_c_1417_n 0.0011921f $X=3.89 $Y=0.795 $X2=0 $Y2=0
cc_432 N_S0_c_473_n N_VGND_c_1417_n 0.02586f $X=3.565 $Y=1.29 $X2=0 $Y2=0
cc_433 N_S0_c_452_n N_VGND_c_1424_n 0.0357798f $X=1.85 $Y=0.18 $X2=0 $Y2=0
cc_434 N_S0_c_451_n N_VGND_c_1425_n 0.0167179f $X=3.815 $Y=0.18 $X2=0 $Y2=0
cc_435 N_S0_c_451_n N_VGND_c_1428_n 0.0638433f $X=3.815 $Y=0.18 $X2=0 $Y2=0
cc_436 N_S0_c_452_n N_VGND_c_1428_n 0.00603775f $X=1.85 $Y=0.18 $X2=0 $Y2=0
cc_437 N_S0_c_453_n N_VGND_c_1428_n 7.88961e-19 $X=2.94 $Y=1.125 $X2=0 $Y2=0
cc_438 N_S0_c_453_n N_A_710_117#_c_1520_n 0.00108271f $X=2.94 $Y=1.125 $X2=0
+ $Y2=0
cc_439 N_S0_M1016_g N_A_710_117#_c_1520_n 0.00625614f $X=3.89 $Y=0.795 $X2=0
+ $Y2=0
cc_440 N_S0_c_458_n N_A_710_117#_c_1520_n 0.00737373f $X=3.89 $Y=1.2 $X2=0 $Y2=0
cc_441 N_S0_c_473_n N_A_710_117#_c_1520_n 0.0121734f $X=3.565 $Y=1.29 $X2=0
+ $Y2=0
cc_442 N_S0_c_451_n N_A_710_117#_c_1521_n 0.00760194f $X=3.815 $Y=0.18 $X2=0
+ $Y2=0
cc_443 N_S0_M1016_g N_A_710_117#_c_1523_n 0.01729f $X=3.89 $Y=0.795 $X2=0 $Y2=0
cc_444 N_A3_c_562_n N_A2_M1015_g 0.00862847f $X=5.145 $Y=1.08 $X2=0 $Y2=0
cc_445 N_A3_c_565_n N_A2_M1015_g 0.0215136f $X=5.252 $Y=0.77 $X2=0 $Y2=0
cc_446 N_A3_c_568_n N_A2_M1015_g 3.97493e-19 $X=5.145 $Y=1.245 $X2=0 $Y2=0
cc_447 N_A3_c_563_n N_A2_c_617_n 0.010339f $X=5.145 $Y=1.585 $X2=0 $Y2=0
cc_448 N_A3_M1019_g N_A2_c_622_n 0.0338025f $X=5.125 $Y=2.715 $X2=0 $Y2=0
cc_449 N_A3_c_564_n N_A2_c_622_n 0.010339f $X=5.145 $Y=1.75 $X2=0 $Y2=0
cc_450 N_A3_c_567_n A2 0.00396779f $X=5.145 $Y=1.245 $X2=0 $Y2=0
cc_451 N_A3_c_568_n A2 0.0447878f $X=5.145 $Y=1.245 $X2=0 $Y2=0
cc_452 N_A3_c_567_n N_A2_c_619_n 0.010339f $X=5.145 $Y=1.245 $X2=0 $Y2=0
cc_453 N_A3_c_568_n N_A2_c_619_n 7.53056e-19 $X=5.145 $Y=1.245 $X2=0 $Y2=0
cc_454 N_A3_M1019_g N_VPWR_c_926_n 0.00187706f $X=5.125 $Y=2.715 $X2=0 $Y2=0
cc_455 N_A3_M1019_g N_VPWR_c_932_n 0.00352627f $X=5.125 $Y=2.715 $X2=0 $Y2=0
cc_456 N_A3_M1019_g N_VPWR_c_923_n 0.00302978f $X=5.125 $Y=2.715 $X2=0 $Y2=0
cc_457 N_A3_M1019_g N_A_284_81#_c_1051_n 0.00134062f $X=5.125 $Y=2.715 $X2=0
+ $Y2=0
cc_458 N_A3_c_568_n N_A_284_81#_c_1051_n 0.0022033f $X=5.145 $Y=1.245 $X2=0
+ $Y2=0
cc_459 N_A3_M1019_g N_A_799_501#_c_1180_n 0.00422754f $X=5.125 $Y=2.715 $X2=0
+ $Y2=0
cc_460 N_A3_M1019_g N_A_799_501#_c_1182_n 0.00943643f $X=5.125 $Y=2.715 $X2=0
+ $Y2=0
cc_461 N_A3_M1019_g N_A_799_501#_c_1183_n 0.00834596f $X=5.125 $Y=2.715 $X2=0
+ $Y2=0
cc_462 N_A3_M1019_g N_A_799_501#_c_1184_n 0.00270904f $X=5.125 $Y=2.715 $X2=0
+ $Y2=0
cc_463 N_A3_c_562_n N_A_793_117#_c_1226_n 0.00211385f $X=5.145 $Y=1.08 $X2=0
+ $Y2=0
cc_464 N_A3_c_567_n N_A_793_117#_c_1226_n 4.63259e-19 $X=5.145 $Y=1.245 $X2=0
+ $Y2=0
cc_465 N_A3_c_568_n N_A_793_117#_c_1226_n 0.00919045f $X=5.145 $Y=1.245 $X2=0
+ $Y2=0
cc_466 N_A3_M1019_g N_A_793_117#_c_1228_n 0.00311965f $X=5.125 $Y=2.715 $X2=0
+ $Y2=0
cc_467 N_A3_c_567_n N_A_793_117#_c_1228_n 0.00168105f $X=5.145 $Y=1.245 $X2=0
+ $Y2=0
cc_468 N_A3_c_568_n N_A_793_117#_c_1228_n 0.0454039f $X=5.145 $Y=1.245 $X2=0
+ $Y2=0
cc_469 N_A3_M1019_g N_A_793_117#_c_1232_n 0.00120726f $X=5.125 $Y=2.715 $X2=0
+ $Y2=0
cc_470 N_A3_M1019_g N_A_793_117#_c_1233_n 0.00954074f $X=5.125 $Y=2.715 $X2=0
+ $Y2=0
cc_471 N_A3_c_564_n N_A_793_117#_c_1233_n 0.00396785f $X=5.145 $Y=1.75 $X2=0
+ $Y2=0
cc_472 N_A3_c_568_n N_A_793_117#_c_1233_n 0.0204612f $X=5.145 $Y=1.245 $X2=0
+ $Y2=0
cc_473 N_A3_c_565_n N_VGND_c_1418_n 0.00435875f $X=5.252 $Y=0.77 $X2=0 $Y2=0
cc_474 N_A3_c_565_n N_VGND_c_1425_n 0.00415117f $X=5.252 $Y=0.77 $X2=0 $Y2=0
cc_475 N_A3_c_565_n N_VGND_c_1428_n 0.00724772f $X=5.252 $Y=0.77 $X2=0 $Y2=0
cc_476 N_A3_c_565_n N_A_710_117#_c_1522_n 0.0027795f $X=5.252 $Y=0.77 $X2=0
+ $Y2=0
cc_477 N_A3_c_565_n N_A_879_117#_c_1546_n 0.00968327f $X=5.252 $Y=0.77 $X2=0
+ $Y2=0
cc_478 N_A3_c_566_n N_A_879_117#_c_1546_n 0.0108393f $X=5.252 $Y=0.92 $X2=0
+ $Y2=0
cc_479 N_A3_c_567_n N_A_879_117#_c_1546_n 0.00118952f $X=5.145 $Y=1.245 $X2=0
+ $Y2=0
cc_480 N_A3_c_568_n N_A_879_117#_c_1546_n 0.0178225f $X=5.145 $Y=1.245 $X2=0
+ $Y2=0
cc_481 N_A3_c_565_n N_A_879_117#_c_1548_n 7.66338e-19 $X=5.252 $Y=0.77 $X2=0
+ $Y2=0
cc_482 N_A2_M1025_g N_A_1245_21#_c_744_n 0.021166f $X=5.625 $Y=2.715 $X2=0 $Y2=0
cc_483 N_A2_M1015_g N_A_1245_21#_c_731_n 0.0264549f $X=5.78 $Y=0.445 $X2=0 $Y2=0
cc_484 N_A2_c_617_n N_A_1245_21#_c_737_n 0.00771985f $X=5.715 $Y=1.665 $X2=0
+ $Y2=0
cc_485 N_A2_c_622_n N_A_1245_21#_c_738_n 0.00771985f $X=5.715 $Y=1.83 $X2=0
+ $Y2=0
cc_486 A2 N_A_1245_21#_c_757_n 0.0242214f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_487 N_A2_c_619_n N_A_1245_21#_c_757_n 0.0024337f $X=5.715 $Y=1.325 $X2=0
+ $Y2=0
cc_488 A2 N_A_1245_21#_c_740_n 0.0022699f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_489 N_A2_c_619_n N_A_1245_21#_c_740_n 0.00771985f $X=5.715 $Y=1.325 $X2=0
+ $Y2=0
cc_490 N_A2_M1015_g N_A_1245_21#_c_742_n 8.3801e-19 $X=5.78 $Y=0.445 $X2=0 $Y2=0
cc_491 N_A2_M1025_g N_VPWR_c_926_n 0.00361744f $X=5.625 $Y=2.715 $X2=0 $Y2=0
cc_492 N_A2_M1025_g N_VPWR_c_927_n 0.00552345f $X=5.625 $Y=2.715 $X2=0 $Y2=0
cc_493 N_A2_M1025_g N_VPWR_c_923_n 0.00534666f $X=5.625 $Y=2.715 $X2=0 $Y2=0
cc_494 N_A2_M1025_g N_A_284_81#_c_1051_n 0.00134123f $X=5.625 $Y=2.715 $X2=0
+ $Y2=0
cc_495 A2 N_A_284_81#_c_1051_n 0.00361615f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_496 N_A2_M1025_g N_A_799_501#_c_1182_n 5.64248e-19 $X=5.625 $Y=2.715 $X2=0
+ $Y2=0
cc_497 N_A2_M1025_g N_A_799_501#_c_1183_n 0.0155792f $X=5.625 $Y=2.715 $X2=0
+ $Y2=0
cc_498 N_A2_M1025_g N_A_799_501#_c_1185_n 0.00117516f $X=5.625 $Y=2.715 $X2=0
+ $Y2=0
cc_499 N_A2_M1025_g N_A_793_117#_c_1233_n 0.010925f $X=5.625 $Y=2.715 $X2=0
+ $Y2=0
cc_500 N_A2_c_622_n N_A_793_117#_c_1233_n 0.00511977f $X=5.715 $Y=1.83 $X2=0
+ $Y2=0
cc_501 A2 N_A_793_117#_c_1233_n 0.0341254f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_502 N_A2_M1015_g N_VGND_c_1418_n 0.00742172f $X=5.78 $Y=0.445 $X2=0 $Y2=0
cc_503 N_A2_M1015_g N_VGND_c_1419_n 7.53527e-19 $X=5.78 $Y=0.445 $X2=0 $Y2=0
cc_504 N_A2_M1015_g N_VGND_c_1421_n 0.0038319f $X=5.78 $Y=0.445 $X2=0 $Y2=0
cc_505 N_A2_M1015_g N_VGND_c_1428_n 0.00473239f $X=5.78 $Y=0.445 $X2=0 $Y2=0
cc_506 N_A2_M1015_g N_A_879_117#_c_1546_n 0.0145216f $X=5.78 $Y=0.445 $X2=0
+ $Y2=0
cc_507 A2 N_A_879_117#_c_1546_n 0.0215251f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_508 N_A2_c_619_n N_A_879_117#_c_1546_n 0.00434694f $X=5.715 $Y=1.325 $X2=0
+ $Y2=0
cc_509 N_S1_c_670_n N_A_1245_21#_c_744_n 0.0250966f $X=6.96 $Y=1.945 $X2=0 $Y2=0
cc_510 N_S1_c_673_p N_A_1245_21#_c_744_n 3.93386e-19 $X=6.96 $Y=1.44 $X2=0 $Y2=0
cc_511 N_S1_M1004_g N_A_1245_21#_c_730_n 0.0103107f $X=6.87 $Y=0.805 $X2=0 $Y2=0
cc_512 N_S1_c_663_n N_A_1245_21#_c_730_n 0.004313f $X=8.1 $Y=1.275 $X2=0 $Y2=0
cc_513 N_S1_M1010_g N_A_1245_21#_c_745_n 0.0104426f $X=6.87 $Y=2.435 $X2=0 $Y2=0
cc_514 N_S1_c_663_n N_A_1245_21#_c_732_n 0.0132093f $X=8.1 $Y=1.275 $X2=0 $Y2=0
cc_515 N_S1_M1017_g N_A_1245_21#_M1022_g 0.0132093f $X=8.1 $Y=2.045 $X2=0 $Y2=0
cc_516 N_S1_M1004_g N_A_1245_21#_c_736_n 0.0114353f $X=6.87 $Y=0.805 $X2=0 $Y2=0
cc_517 N_S1_c_665_n N_A_1245_21#_c_737_n 0.0121181f $X=6.96 $Y=1.35 $X2=0 $Y2=0
cc_518 N_S1_c_673_p N_A_1245_21#_c_737_n 0.00171118f $X=6.96 $Y=1.44 $X2=0 $Y2=0
cc_519 N_S1_c_667_n N_A_1245_21#_c_738_n 0.0121181f $X=6.96 $Y=1.44 $X2=0 $Y2=0
cc_520 N_S1_c_666_n N_A_1245_21#_c_739_n 0.0132093f $X=8.1 $Y=1.35 $X2=0 $Y2=0
cc_521 N_S1_M1004_g N_A_1245_21#_c_757_n 0.00272563f $X=6.87 $Y=0.805 $X2=0
+ $Y2=0
cc_522 N_S1_c_673_p N_A_1245_21#_c_757_n 0.023301f $X=6.96 $Y=1.44 $X2=0 $Y2=0
cc_523 N_S1_M1004_g N_A_1245_21#_c_740_n 0.0121181f $X=6.87 $Y=0.805 $X2=0 $Y2=0
cc_524 N_S1_M1004_g N_A_1245_21#_c_741_n 0.0157395f $X=6.87 $Y=0.805 $X2=0 $Y2=0
cc_525 N_S1_c_665_n N_A_1245_21#_c_741_n 0.00875173f $X=6.96 $Y=1.35 $X2=0 $Y2=0
cc_526 N_S1_c_673_p N_A_1245_21#_c_741_n 0.0259822f $X=6.96 $Y=1.44 $X2=0 $Y2=0
cc_527 N_S1_M1010_g N_A_1245_21#_c_749_n 0.00728803f $X=6.87 $Y=2.435 $X2=0
+ $Y2=0
cc_528 N_S1_c_663_n N_A_1635_149#_c_860_n 0.00150194f $X=8.1 $Y=1.275 $X2=0
+ $Y2=0
cc_529 N_S1_M1017_g N_A_1635_149#_c_866_n 0.00122787f $X=8.1 $Y=2.045 $X2=0
+ $Y2=0
cc_530 N_S1_c_666_n N_A_1635_149#_c_863_n 0.002866f $X=8.1 $Y=1.35 $X2=0 $Y2=0
cc_531 N_S1_M1010_g N_VPWR_c_928_n 0.00285881f $X=6.87 $Y=2.435 $X2=0 $Y2=0
cc_532 N_S1_M1010_g N_VPWR_c_923_n 7.01701e-19 $X=6.87 $Y=2.435 $X2=0 $Y2=0
cc_533 N_S1_c_663_n N_A_284_81#_c_1045_n 0.00706359f $X=8.1 $Y=1.275 $X2=0 $Y2=0
cc_534 N_S1_c_663_n N_A_284_81#_c_1046_n 3.56349e-19 $X=8.1 $Y=1.275 $X2=0 $Y2=0
cc_535 N_S1_M1010_g N_A_284_81#_c_1051_n 0.00299124f $X=6.87 $Y=2.435 $X2=0
+ $Y2=0
cc_536 N_S1_c_662_n N_A_284_81#_c_1051_n 0.00667791f $X=8.025 $Y=1.35 $X2=0
+ $Y2=0
cc_537 N_S1_c_670_n N_A_284_81#_c_1051_n 0.00544277f $X=6.96 $Y=1.945 $X2=0
+ $Y2=0
cc_538 N_S1_c_673_p N_A_284_81#_c_1051_n 0.00849114f $X=6.96 $Y=1.44 $X2=0 $Y2=0
cc_539 N_S1_M1017_g N_A_284_81#_c_1115_n 0.00275504f $X=8.1 $Y=2.045 $X2=0 $Y2=0
cc_540 N_S1_c_662_n N_A_284_81#_c_1116_n 0.00272508f $X=8.025 $Y=1.35 $X2=0
+ $Y2=0
cc_541 N_S1_M1017_g N_A_284_81#_c_1116_n 0.00292665f $X=8.1 $Y=2.045 $X2=0 $Y2=0
cc_542 N_S1_c_662_n N_A_284_81#_c_1050_n 0.0073082f $X=8.025 $Y=1.35 $X2=0 $Y2=0
cc_543 N_S1_c_663_n N_A_284_81#_c_1050_n 0.0192326f $X=8.1 $Y=1.275 $X2=0 $Y2=0
cc_544 N_S1_M1017_g N_A_284_81#_c_1050_n 0.0119108f $X=8.1 $Y=2.045 $X2=0 $Y2=0
cc_545 N_S1_c_666_n N_A_284_81#_c_1050_n 0.00152009f $X=8.1 $Y=1.35 $X2=0 $Y2=0
cc_546 N_S1_M1010_g N_A_793_117#_c_1234_n 0.0149494f $X=6.87 $Y=2.435 $X2=0
+ $Y2=0
cc_547 N_S1_c_662_n N_A_793_117#_c_1234_n 0.00364684f $X=8.025 $Y=1.35 $X2=0
+ $Y2=0
cc_548 N_S1_c_670_n N_A_793_117#_c_1234_n 0.00510425f $X=6.96 $Y=1.945 $X2=0
+ $Y2=0
cc_549 N_S1_c_673_p N_A_793_117#_c_1234_n 0.0216611f $X=6.96 $Y=1.44 $X2=0 $Y2=0
cc_550 N_S1_M1004_g N_A_793_117#_c_1229_n 0.00244974f $X=6.87 $Y=0.805 $X2=0
+ $Y2=0
cc_551 N_S1_M1010_g N_A_793_117#_c_1229_n 0.00156093f $X=6.87 $Y=2.435 $X2=0
+ $Y2=0
cc_552 N_S1_c_662_n N_A_793_117#_c_1229_n 0.0167715f $X=8.025 $Y=1.35 $X2=0
+ $Y2=0
cc_553 N_S1_c_663_n N_A_793_117#_c_1229_n 7.44344e-19 $X=8.1 $Y=1.275 $X2=0
+ $Y2=0
cc_554 N_S1_M1017_g N_A_793_117#_c_1229_n 0.00229716f $X=8.1 $Y=2.045 $X2=0
+ $Y2=0
cc_555 N_S1_c_667_n N_A_793_117#_c_1229_n 0.0115404f $X=6.96 $Y=1.44 $X2=0 $Y2=0
cc_556 N_S1_c_673_p N_A_793_117#_c_1229_n 0.0244684f $X=6.96 $Y=1.44 $X2=0 $Y2=0
cc_557 N_S1_M1010_g N_A_793_117#_c_1236_n 0.00307615f $X=6.87 $Y=2.435 $X2=0
+ $Y2=0
cc_558 N_S1_M1017_g N_A_793_117#_c_1236_n 0.00404557f $X=8.1 $Y=2.045 $X2=0
+ $Y2=0
cc_559 N_S1_M1017_g N_A_793_117#_c_1237_n 0.00851776f $X=8.1 $Y=2.045 $X2=0
+ $Y2=0
cc_560 N_S1_M1010_g N_A_793_117#_c_1241_n 2.27062e-19 $X=6.87 $Y=2.435 $X2=0
+ $Y2=0
cc_561 N_S1_c_670_n N_A_793_117#_c_1241_n 0.00187279f $X=6.96 $Y=1.945 $X2=0
+ $Y2=0
cc_562 N_S1_M1004_g N_A_793_117#_c_1230_n 7.31873e-19 $X=6.87 $Y=0.805 $X2=0
+ $Y2=0
cc_563 N_S1_c_662_n N_A_793_117#_c_1230_n 0.00506739f $X=8.025 $Y=1.35 $X2=0
+ $Y2=0
cc_564 N_S1_c_663_n N_A_793_117#_c_1230_n 0.00170863f $X=8.1 $Y=1.275 $X2=0
+ $Y2=0
cc_565 N_S1_M1004_g N_VGND_c_1419_n 0.0121055f $X=6.87 $Y=0.805 $X2=0 $Y2=0
cc_566 N_S1_M1004_g N_VGND_c_1428_n 7.88961e-19 $X=6.87 $Y=0.805 $X2=0 $Y2=0
cc_567 N_A_1245_21#_c_732_n N_A_1635_149#_c_860_n 0.00494679f $X=8.53 $Y=1.275
+ $X2=0 $Y2=0
cc_568 N_A_1245_21#_M1022_g N_A_1635_149#_c_866_n 0.00424555f $X=8.53 $Y=2.045
+ $X2=0 $Y2=0
cc_569 N_A_1245_21#_M1022_g N_A_1635_149#_c_861_n 0.0180879f $X=8.53 $Y=2.045
+ $X2=0 $Y2=0
cc_570 N_A_1245_21#_c_734_n N_A_1635_149#_c_861_n 0.0265891f $X=8.945 $Y=1.35
+ $X2=0 $Y2=0
cc_571 N_A_1245_21#_c_739_n N_A_1635_149#_c_861_n 0.00901112f $X=8.53 $Y=1.35
+ $X2=0 $Y2=0
cc_572 N_A_1245_21#_M1022_g N_A_1635_149#_c_862_n 0.0024289f $X=8.53 $Y=2.045
+ $X2=0 $Y2=0
cc_573 N_A_1245_21#_c_734_n N_A_1635_149#_c_862_n 0.0052232f $X=8.945 $Y=1.35
+ $X2=0 $Y2=0
cc_574 N_A_1245_21#_c_735_n N_A_1635_149#_c_864_n 0.0165468f $X=9.02 $Y=1.275
+ $X2=0 $Y2=0
cc_575 N_A_1245_21#_c_744_n N_VPWR_c_926_n 0.00185439f $X=6.3 $Y=2.985 $X2=0
+ $Y2=0
cc_576 N_A_1245_21#_c_746_n N_VPWR_c_927_n 0.00612772f $X=6.375 $Y=3.06 $X2=0
+ $Y2=0
cc_577 N_A_1245_21#_c_744_n N_VPWR_c_928_n 0.0127161f $X=6.3 $Y=2.985 $X2=0
+ $Y2=0
cc_578 N_A_1245_21#_c_745_n N_VPWR_c_928_n 0.0262563f $X=7.32 $Y=3.06 $X2=0
+ $Y2=0
cc_579 N_A_1245_21#_c_738_n N_VPWR_c_928_n 2.52772e-19 $X=6.39 $Y=1.795 $X2=0
+ $Y2=0
cc_580 N_A_1245_21#_c_749_n N_VPWR_c_928_n 0.020776f $X=7.085 $Y=2.48 $X2=0
+ $Y2=0
cc_581 N_A_1245_21#_c_750_n N_VPWR_c_928_n 0.025373f $X=7.25 $Y=2.927 $X2=0
+ $Y2=0
cc_582 N_A_1245_21#_c_752_n N_VPWR_c_928_n 6.6504e-19 $X=7.485 $Y=2.945 $X2=0
+ $Y2=0
cc_583 N_A_1245_21#_M1022_g N_VPWR_c_929_n 0.00168884f $X=8.53 $Y=2.045 $X2=0
+ $Y2=0
cc_584 N_A_1245_21#_c_745_n N_VPWR_c_933_n 0.0183215f $X=7.32 $Y=3.06 $X2=0
+ $Y2=0
cc_585 N_A_1245_21#_c_750_n N_VPWR_c_933_n 0.0225443f $X=7.25 $Y=2.927 $X2=0
+ $Y2=0
cc_586 N_A_1245_21#_c_751_n N_VPWR_c_933_n 0.0254727f $X=7.485 $Y=2.945 $X2=0
+ $Y2=0
cc_587 N_A_1245_21#_c_745_n N_VPWR_c_923_n 0.0180856f $X=7.32 $Y=3.06 $X2=0
+ $Y2=0
cc_588 N_A_1245_21#_c_746_n N_VPWR_c_923_n 0.00998482f $X=6.375 $Y=3.06 $X2=0
+ $Y2=0
cc_589 N_A_1245_21#_c_750_n N_VPWR_c_923_n 0.0113294f $X=7.25 $Y=2.927 $X2=0
+ $Y2=0
cc_590 N_A_1245_21#_c_751_n N_VPWR_c_923_n 0.01336f $X=7.485 $Y=2.945 $X2=0
+ $Y2=0
cc_591 N_A_1245_21#_c_752_n N_VPWR_c_923_n 0.00867605f $X=7.485 $Y=2.945 $X2=0
+ $Y2=0
cc_592 N_A_1245_21#_c_730_n N_A_284_81#_c_1045_n 0.0142686f $X=8.945 $Y=0.18
+ $X2=0 $Y2=0
cc_593 N_A_1245_21#_c_732_n N_A_284_81#_c_1045_n 0.00854467f $X=8.53 $Y=1.275
+ $X2=0 $Y2=0
cc_594 N_A_1245_21#_c_735_n N_A_284_81#_c_1045_n 0.00604384f $X=9.02 $Y=1.275
+ $X2=0 $Y2=0
cc_595 N_A_1245_21#_c_730_n N_A_284_81#_c_1046_n 0.0036023f $X=8.945 $Y=0.18
+ $X2=0 $Y2=0
cc_596 N_A_1245_21#_c_732_n N_A_284_81#_c_1047_n 0.00194992f $X=8.53 $Y=1.275
+ $X2=0 $Y2=0
cc_597 N_A_1245_21#_c_734_n N_A_284_81#_c_1047_n 0.00340068f $X=8.945 $Y=1.35
+ $X2=0 $Y2=0
cc_598 N_A_1245_21#_c_735_n N_A_284_81#_c_1047_n 0.00543761f $X=9.02 $Y=1.275
+ $X2=0 $Y2=0
cc_599 N_A_1245_21#_c_744_n N_A_284_81#_c_1051_n 0.00616318f $X=6.3 $Y=2.985
+ $X2=0 $Y2=0
cc_600 N_A_1245_21#_c_757_n N_A_284_81#_c_1051_n 0.00246552f $X=6.39 $Y=1.29
+ $X2=0 $Y2=0
cc_601 N_A_1245_21#_c_749_n N_A_284_81#_c_1051_n 0.00221311f $X=7.085 $Y=2.48
+ $X2=0 $Y2=0
cc_602 N_A_1245_21#_c_732_n N_A_284_81#_c_1050_n 6.0711e-19 $X=8.53 $Y=1.275
+ $X2=0 $Y2=0
cc_603 N_A_1245_21#_M1022_g N_A_284_81#_c_1050_n 2.36695e-19 $X=8.53 $Y=2.045
+ $X2=0 $Y2=0
cc_604 N_A_1245_21#_c_739_n N_A_284_81#_c_1050_n 2.40763e-19 $X=8.53 $Y=1.35
+ $X2=0 $Y2=0
cc_605 N_A_1245_21#_c_743_n N_A_284_81#_c_1050_n 0.0046335f $X=7.085 $Y=0.805
+ $X2=0 $Y2=0
cc_606 N_A_1245_21#_c_744_n N_A_799_501#_c_1183_n 0.0036015f $X=6.3 $Y=2.985
+ $X2=0 $Y2=0
cc_607 N_A_1245_21#_c_744_n N_A_799_501#_c_1185_n 0.00440422f $X=6.3 $Y=2.985
+ $X2=0 $Y2=0
cc_608 N_A_1245_21#_c_744_n N_A_793_117#_c_1233_n 0.0124f $X=6.3 $Y=2.985 $X2=0
+ $Y2=0
cc_609 N_A_1245_21#_c_738_n N_A_793_117#_c_1233_n 0.0018813f $X=6.39 $Y=1.795
+ $X2=0 $Y2=0
cc_610 N_A_1245_21#_c_757_n N_A_793_117#_c_1233_n 0.0153173f $X=6.39 $Y=1.29
+ $X2=0 $Y2=0
cc_611 N_A_1245_21#_c_749_n N_A_793_117#_c_1234_n 0.022684f $X=7.085 $Y=2.48
+ $X2=0 $Y2=0
cc_612 N_A_1245_21#_c_751_n N_A_793_117#_c_1234_n 0.0055892f $X=7.485 $Y=2.945
+ $X2=0 $Y2=0
cc_613 N_A_1245_21#_c_752_n N_A_793_117#_c_1234_n 0.00182841f $X=7.485 $Y=2.945
+ $X2=0 $Y2=0
cc_614 N_A_1245_21#_c_741_n N_A_793_117#_c_1229_n 0.00527179f $X=7 $Y=1.1 $X2=0
+ $Y2=0
cc_615 N_A_1245_21#_c_749_n N_A_793_117#_c_1236_n 3.44607e-19 $X=7.085 $Y=2.48
+ $X2=0 $Y2=0
cc_616 N_A_1245_21#_M1022_g N_A_793_117#_c_1237_n 0.00975286f $X=8.53 $Y=2.045
+ $X2=0 $Y2=0
cc_617 N_A_1245_21#_c_751_n N_A_793_117#_c_1237_n 0.00362542f $X=7.485 $Y=2.945
+ $X2=0 $Y2=0
cc_618 N_A_1245_21#_c_752_n N_A_793_117#_c_1237_n 0.00114358f $X=7.485 $Y=2.945
+ $X2=0 $Y2=0
cc_619 N_A_1245_21#_c_749_n N_A_793_117#_c_1238_n 0.0195377f $X=7.085 $Y=2.48
+ $X2=0 $Y2=0
cc_620 N_A_1245_21#_c_751_n N_A_793_117#_c_1238_n 0.0135346f $X=7.485 $Y=2.945
+ $X2=0 $Y2=0
cc_621 N_A_1245_21#_c_752_n N_A_793_117#_c_1238_n 0.00401199f $X=7.485 $Y=2.945
+ $X2=0 $Y2=0
cc_622 N_A_1245_21#_M1022_g N_A_793_117#_c_1239_n 0.00560037f $X=8.53 $Y=2.045
+ $X2=0 $Y2=0
cc_623 N_A_1245_21#_c_734_n N_A_793_117#_c_1239_n 9.91663e-19 $X=8.945 $Y=1.35
+ $X2=0 $Y2=0
cc_624 N_A_1245_21#_c_744_n N_A_793_117#_c_1241_n 0.00294528f $X=6.3 $Y=2.985
+ $X2=0 $Y2=0
cc_625 N_A_1245_21#_c_738_n N_A_793_117#_c_1241_n 0.00297768f $X=6.39 $Y=1.795
+ $X2=0 $Y2=0
cc_626 N_A_1245_21#_c_757_n N_A_793_117#_c_1241_n 0.00817467f $X=6.39 $Y=1.29
+ $X2=0 $Y2=0
cc_627 N_A_1245_21#_c_730_n N_A_793_117#_c_1230_n 0.00709325f $X=8.945 $Y=0.18
+ $X2=0 $Y2=0
cc_628 N_A_1245_21#_c_741_n N_A_793_117#_c_1230_n 0.00877079f $X=7 $Y=1.1 $X2=0
+ $Y2=0
cc_629 N_A_1245_21#_c_743_n N_A_793_117#_c_1230_n 0.017366f $X=7.085 $Y=0.805
+ $X2=0 $Y2=0
cc_630 N_A_1245_21#_c_742_n N_VGND_M1004_s 2.76656e-19 $X=6.555 $Y=1.1 $X2=0
+ $Y2=0
cc_631 N_A_1245_21#_c_731_n N_VGND_c_1418_n 0.00117161f $X=6.375 $Y=0.18 $X2=0
+ $Y2=0
cc_632 N_A_1245_21#_c_730_n N_VGND_c_1419_n 0.0248713f $X=8.945 $Y=0.18 $X2=0
+ $Y2=0
cc_633 N_A_1245_21#_c_736_n N_VGND_c_1419_n 0.00913038f $X=6.39 $Y=1.125 $X2=0
+ $Y2=0
cc_634 N_A_1245_21#_c_740_n N_VGND_c_1419_n 3.80919e-19 $X=6.39 $Y=1.29 $X2=0
+ $Y2=0
cc_635 N_A_1245_21#_c_741_n N_VGND_c_1419_n 0.0190355f $X=7 $Y=1.1 $X2=0 $Y2=0
cc_636 N_A_1245_21#_c_742_n N_VGND_c_1419_n 0.00590791f $X=6.555 $Y=1.1 $X2=0
+ $Y2=0
cc_637 N_A_1245_21#_c_730_n N_VGND_c_1420_n 0.0178829f $X=8.945 $Y=0.18 $X2=0
+ $Y2=0
cc_638 N_A_1245_21#_c_731_n N_VGND_c_1421_n 0.0102096f $X=6.375 $Y=0.18 $X2=0
+ $Y2=0
cc_639 N_A_1245_21#_c_730_n N_VGND_c_1426_n 0.0647193f $X=8.945 $Y=0.18 $X2=0
+ $Y2=0
cc_640 N_A_1245_21#_c_743_n N_VGND_c_1426_n 0.00467787f $X=7.085 $Y=0.805 $X2=0
+ $Y2=0
cc_641 N_A_1245_21#_c_730_n N_VGND_c_1428_n 0.0857915f $X=8.945 $Y=0.18 $X2=0
+ $Y2=0
cc_642 N_A_1245_21#_c_731_n N_VGND_c_1428_n 0.0103883f $X=6.375 $Y=0.18 $X2=0
+ $Y2=0
cc_643 N_A_1245_21#_c_743_n N_VGND_c_1428_n 0.00643971f $X=7.085 $Y=0.805 $X2=0
+ $Y2=0
cc_644 N_A_1245_21#_c_736_n N_A_879_117#_c_1546_n 0.00241888f $X=6.39 $Y=1.125
+ $X2=0 $Y2=0
cc_645 N_A_1245_21#_c_736_n N_A_879_117#_c_1547_n 0.00395609f $X=6.39 $Y=1.125
+ $X2=0 $Y2=0
cc_646 N_A_1635_149#_M1002_g N_VPWR_c_929_n 0.0237794f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_647 N_A_1635_149#_c_861_n N_VPWR_c_929_n 0.0248138f $X=9.47 $Y=1.51 $X2=0
+ $Y2=0
cc_648 N_A_1635_149#_c_862_n N_VPWR_c_929_n 0.00506784f $X=9.47 $Y=1.51 $X2=0
+ $Y2=0
cc_649 N_A_1635_149#_M1002_g N_VPWR_c_934_n 0.00486043f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_650 N_A_1635_149#_M1002_g N_VPWR_c_923_n 0.00917987f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_651 N_A_1635_149#_c_860_n N_A_284_81#_c_1045_n 0.0158362f $X=8.315 $Y=0.955
+ $X2=0 $Y2=0
cc_652 N_A_1635_149#_c_861_n N_A_284_81#_c_1047_n 0.0178926f $X=9.47 $Y=1.51
+ $X2=0 $Y2=0
cc_653 N_A_1635_149#_c_866_n N_A_284_81#_c_1115_n 0.0064667f $X=8.315 $Y=2.045
+ $X2=0 $Y2=0
cc_654 N_A_1635_149#_c_860_n N_A_284_81#_c_1050_n 0.0257635f $X=8.315 $Y=0.955
+ $X2=0 $Y2=0
cc_655 N_A_1635_149#_c_866_n N_A_284_81#_c_1050_n 0.0242257f $X=8.315 $Y=2.045
+ $X2=0 $Y2=0
cc_656 N_A_1635_149#_c_863_n N_A_284_81#_c_1050_n 0.0265873f $X=8.332 $Y=1.51
+ $X2=0 $Y2=0
cc_657 N_A_1635_149#_c_866_n N_A_793_117#_c_1237_n 0.0160798f $X=8.315 $Y=2.045
+ $X2=0 $Y2=0
cc_658 N_A_1635_149#_M1002_g N_A_793_117#_c_1239_n 0.00115982f $X=9.605 $Y=2.465
+ $X2=0 $Y2=0
cc_659 N_A_1635_149#_c_861_n N_A_793_117#_c_1239_n 0.0160202f $X=9.47 $Y=1.51
+ $X2=0 $Y2=0
cc_660 N_A_1635_149#_c_861_n X 0.0271104f $X=9.47 $Y=1.51 $X2=0 $Y2=0
cc_661 N_A_1635_149#_c_864_n X 0.0265179f $X=9.492 $Y=1.345 $X2=0 $Y2=0
cc_662 N_A_1635_149#_c_861_n N_VGND_c_1420_n 0.0248138f $X=9.47 $Y=1.51 $X2=0
+ $Y2=0
cc_663 N_A_1635_149#_c_862_n N_VGND_c_1420_n 0.00506784f $X=9.47 $Y=1.51 $X2=0
+ $Y2=0
cc_664 N_A_1635_149#_c_864_n N_VGND_c_1420_n 0.0180198f $X=9.492 $Y=1.345 $X2=0
+ $Y2=0
cc_665 N_A_1635_149#_c_864_n N_VGND_c_1427_n 0.00465077f $X=9.492 $Y=1.345 $X2=0
+ $Y2=0
cc_666 N_A_1635_149#_c_864_n N_VGND_c_1428_n 0.00451796f $X=9.492 $Y=1.345 $X2=0
+ $Y2=0
cc_667 N_A_27_519#_c_903_n N_VPWR_c_924_n 0.0209198f $X=1.475 $Y=2.43 $X2=0
+ $Y2=0
cc_668 N_A_27_519#_c_902_n N_VPWR_c_930_n 0.0105318f $X=0.26 $Y=2.805 $X2=0
+ $Y2=0
cc_669 N_A_27_519#_c_902_n N_VPWR_c_923_n 0.00944361f $X=0.26 $Y=2.805 $X2=0
+ $Y2=0
cc_670 N_A_27_519#_c_903_n N_VPWR_c_923_n 0.0123129f $X=1.475 $Y=2.43 $X2=0
+ $Y2=0
cc_671 N_A_27_519#_c_903_n N_A_196_519#_c_1021_n 0.00763428f $X=1.475 $Y=2.43
+ $X2=0 $Y2=0
cc_672 N_A_27_519#_c_905_n N_A_196_519#_c_1021_n 0.0171104f $X=1.605 $Y=2.43
+ $X2=0 $Y2=0
cc_673 N_A_27_519#_c_903_n N_A_196_519#_c_1023_n 0.0193364f $X=1.475 $Y=2.43
+ $X2=0 $Y2=0
cc_674 N_VPWR_c_931_n N_A_196_519#_c_1021_n 0.0725786f $X=3.345 $Y=3.33 $X2=0
+ $Y2=0
cc_675 N_VPWR_c_923_n N_A_196_519#_c_1021_n 0.0509917f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_924_n N_A_196_519#_c_1023_n 0.0138953f $X=0.69 $Y=2.805 $X2=0
+ $Y2=0
cc_677 N_VPWR_c_931_n N_A_196_519#_c_1023_n 0.0140542f $X=3.345 $Y=3.33 $X2=0
+ $Y2=0
cc_678 N_VPWR_c_923_n N_A_196_519#_c_1023_n 0.00964728f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_679 N_VPWR_c_925_n N_A_284_81#_c_1051_n 0.00230201f $X=3.48 $Y=2.68 $X2=0
+ $Y2=0
cc_680 N_VPWR_c_928_n N_A_284_81#_c_1051_n 0.00292759f $X=6.585 $Y=2.48 $X2=0
+ $Y2=0
cc_681 N_VPWR_c_925_n N_A_799_501#_c_1179_n 0.0191949f $X=3.48 $Y=2.68 $X2=0
+ $Y2=0
cc_682 N_VPWR_c_926_n N_A_799_501#_c_1180_n 0.0140344f $X=5.385 $Y=2.78 $X2=0
+ $Y2=0
cc_683 N_VPWR_c_932_n N_A_799_501#_c_1180_n 0.0597618f $X=5.285 $Y=3.33 $X2=0
+ $Y2=0
cc_684 N_VPWR_c_923_n N_A_799_501#_c_1180_n 0.0344183f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_685 N_VPWR_c_925_n N_A_799_501#_c_1181_n 0.00983147f $X=3.48 $Y=2.68 $X2=0
+ $Y2=0
cc_686 N_VPWR_c_932_n N_A_799_501#_c_1181_n 0.0175915f $X=5.285 $Y=3.33 $X2=0
+ $Y2=0
cc_687 N_VPWR_c_923_n N_A_799_501#_c_1181_n 0.00965744f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_688 N_VPWR_c_926_n N_A_799_501#_c_1182_n 0.0209516f $X=5.385 $Y=2.78 $X2=0
+ $Y2=0
cc_689 N_VPWR_c_926_n N_A_799_501#_c_1183_n 0.0180403f $X=5.385 $Y=2.78 $X2=0
+ $Y2=0
cc_690 N_VPWR_c_928_n N_A_799_501#_c_1183_n 0.00338276f $X=6.585 $Y=2.48 $X2=0
+ $Y2=0
cc_691 N_VPWR_c_927_n N_A_799_501#_c_1185_n 0.00839504f $X=6.41 $Y=3.33 $X2=0
+ $Y2=0
cc_692 N_VPWR_c_928_n N_A_799_501#_c_1185_n 0.0196727f $X=6.585 $Y=2.48 $X2=0
+ $Y2=0
cc_693 N_VPWR_c_923_n N_A_799_501#_c_1185_n 0.0102726f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_694 N_VPWR_c_928_n N_A_793_117#_c_1233_n 0.001569f $X=6.585 $Y=2.48 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_928_n N_A_793_117#_c_1234_n 0.00976926f $X=6.585 $Y=2.48 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_929_n N_A_793_117#_c_1237_n 0.01175f $X=9.39 $Y=1.98 $X2=0 $Y2=0
cc_697 N_VPWR_c_933_n N_A_793_117#_c_1237_n 0.0191817f $X=9.225 $Y=3.33 $X2=0
+ $Y2=0
cc_698 N_VPWR_c_923_n N_A_793_117#_c_1237_n 0.0329256f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_699 N_VPWR_c_929_n N_A_793_117#_c_1239_n 0.0229123f $X=9.39 $Y=1.98 $X2=0
+ $Y2=0
cc_700 N_VPWR_c_928_n N_A_793_117#_c_1241_n 0.0133207f $X=6.585 $Y=2.48 $X2=0
+ $Y2=0
cc_701 N_VPWR_c_923_n N_X_M1002_d 0.00371702f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_702 N_VPWR_c_934_n X 0.018528f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_703 N_VPWR_c_923_n X 0.0104192f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_704 N_A_196_519#_c_1021_n N_A_284_81#_c_1063_n 0.0186346f $X=2.405 $Y=2.95
+ $X2=0 $Y2=0
cc_705 N_A_196_519#_c_1022_n N_A_284_81#_c_1051_n 0.00672729f $X=2.5 $Y=2.505
+ $X2=0 $Y2=0
cc_706 N_A_284_81#_c_1051_n N_A_799_501#_c_1179_n 0.00183788f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_707 N_A_284_81#_c_1051_n N_A_799_501#_c_1183_n 0.0217211f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_708 N_A_284_81#_c_1051_n N_A_799_501#_c_1184_n 0.00416872f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_709 N_A_284_81#_c_1050_n N_A_793_117#_M1001_s 0.00502816f $X=7.915 $Y=1.88
+ $X2=0 $Y2=0
cc_710 N_A_284_81#_c_1051_n N_A_793_117#_c_1233_n 0.0745108f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_711 N_A_284_81#_c_1051_n N_A_793_117#_c_1234_n 0.0393819f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_712 N_A_284_81#_c_1051_n N_A_793_117#_c_1229_n 0.0092236f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_713 N_A_284_81#_c_1115_n N_A_793_117#_c_1229_n 0.00128795f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_714 N_A_284_81#_c_1116_n N_A_793_117#_c_1229_n 0.0102938f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_715 N_A_284_81#_c_1050_n N_A_793_117#_c_1229_n 0.0390789f $X=7.915 $Y=1.88
+ $X2=0 $Y2=0
cc_716 N_A_284_81#_c_1116_n N_A_793_117#_c_1236_n 3.31159e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_717 N_A_284_81#_c_1051_n N_A_793_117#_c_1237_n 0.00734222f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_718 N_A_284_81#_c_1115_n N_A_793_117#_c_1237_n 0.00266409f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_719 N_A_284_81#_c_1116_n N_A_793_117#_c_1237_n 0.017701f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_720 N_A_284_81#_c_1051_n N_A_793_117#_c_1256_n 0.00693504f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_721 N_A_284_81#_c_1051_n N_A_793_117#_c_1240_n 0.0158485f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_722 N_A_284_81#_c_1051_n N_A_793_117#_c_1241_n 0.0108238f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_723 N_A_284_81#_c_1050_n N_A_793_117#_c_1230_n 0.0248702f $X=7.915 $Y=1.88
+ $X2=0 $Y2=0
cc_724 N_A_284_81#_c_1051_n N_A_793_117#_c_1242_n 0.010455f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_725 N_A_284_81#_c_1115_n N_A_793_117#_c_1242_n 0.00133146f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_726 N_A_284_81#_c_1116_n N_A_793_117#_c_1242_n 0.0123634f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_727 N_A_284_81#_c_1048_n N_A_33_81#_c_1373_n 0.0138216f $X=1.56 $Y=0.7 $X2=0
+ $Y2=0
cc_728 N_A_284_81#_M1009_d N_A_33_81#_c_1375_n 0.00180746f $X=1.42 $Y=0.405
+ $X2=0 $Y2=0
cc_729 N_A_284_81#_c_1044_n N_A_33_81#_c_1375_n 0.00433484f $X=1.905 $Y=0.92
+ $X2=0 $Y2=0
cc_730 N_A_284_81#_c_1048_n N_A_33_81#_c_1375_n 0.0146114f $X=1.56 $Y=0.7 $X2=0
+ $Y2=0
cc_731 N_A_284_81#_c_1044_n N_A_33_81#_c_1377_n 0.0145734f $X=1.905 $Y=0.92
+ $X2=0 $Y2=0
cc_732 N_A_284_81#_c_1045_n N_VGND_c_1420_n 0.0132082f $X=8.615 $Y=0.505 $X2=0
+ $Y2=0
cc_733 N_A_284_81#_c_1047_n N_VGND_c_1420_n 0.0268278f $X=8.745 $Y=0.955 $X2=0
+ $Y2=0
cc_734 N_A_284_81#_c_1045_n N_VGND_c_1426_n 0.0313323f $X=8.615 $Y=0.505 $X2=0
+ $Y2=0
cc_735 N_A_284_81#_c_1046_n N_VGND_c_1426_n 0.00652607f $X=8.05 $Y=0.505 $X2=0
+ $Y2=0
cc_736 N_A_284_81#_c_1044_n N_VGND_c_1428_n 4.88312e-19 $X=1.905 $Y=0.92 $X2=0
+ $Y2=0
cc_737 N_A_284_81#_c_1045_n N_VGND_c_1428_n 0.0267735f $X=8.615 $Y=0.505 $X2=0
+ $Y2=0
cc_738 N_A_284_81#_c_1046_n N_VGND_c_1428_n 0.00544303f $X=8.05 $Y=0.505 $X2=0
+ $Y2=0
cc_739 N_A_799_501#_c_1180_n N_A_793_117#_M1003_d 0.00176891f $X=4.945 $Y=2.99
+ $X2=0 $Y2=0
cc_740 N_A_799_501#_c_1182_n N_A_793_117#_c_1232_n 0.00565754f $X=5.03 $Y=2.905
+ $X2=0 $Y2=0
cc_741 N_A_799_501#_c_1184_n N_A_793_117#_c_1232_n 0.0137149f $X=5.115 $Y=2.36
+ $X2=0 $Y2=0
cc_742 N_A_799_501#_c_1183_n N_A_793_117#_c_1233_n 0.0591959f $X=5.705 $Y=2.36
+ $X2=0 $Y2=0
cc_743 N_A_799_501#_c_1184_n N_A_793_117#_c_1233_n 0.0120129f $X=5.115 $Y=2.36
+ $X2=0 $Y2=0
cc_744 N_A_799_501#_c_1180_n N_A_793_117#_c_1256_n 0.0185491f $X=4.945 $Y=2.99
+ $X2=0 $Y2=0
cc_745 N_A_799_501#_c_1182_n N_A_793_117#_c_1256_n 0.0156377f $X=5.03 $Y=2.905
+ $X2=0 $Y2=0
cc_746 N_A_799_501#_c_1180_n A_968_501# 0.00179331f $X=4.945 $Y=2.99 $X2=-0.19
+ $Y2=1.655
cc_747 N_A_799_501#_c_1182_n A_968_501# 0.00376962f $X=5.03 $Y=2.905 $X2=-0.19
+ $Y2=1.655
cc_748 N_A_793_117#_c_1230_n N_VGND_c_1428_n 0.00967032f $X=7.615 $Y=0.955 $X2=0
+ $Y2=0
cc_749 N_A_793_117#_c_1243_n N_A_710_117#_c_1523_n 0.0143371f $X=4.105 $Y=0.79
+ $X2=0 $Y2=0
cc_750 N_A_793_117#_c_1226_n N_A_710_117#_c_1523_n 0.00506028f $X=4.605 $Y=1.1
+ $X2=0 $Y2=0
cc_751 N_A_793_117#_c_1226_n N_A_879_117#_c_1548_n 0.0298633f $X=4.605 $Y=1.1
+ $X2=0 $Y2=0
cc_752 X N_VGND_c_1420_n 0.0307847f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_753 X N_VGND_c_1427_n 0.0108661f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_754 X N_VGND_c_1428_n 0.00974763f $X=9.755 $Y=0.47 $X2=0 $Y2=0
cc_755 N_A_33_81#_c_1373_n N_VGND_M1014_d 0.00226049f $X=1.055 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_756 N_A_33_81#_c_1373_n N_VGND_c_1416_n 0.0188922f $X=1.055 $Y=0.9 $X2=0
+ $Y2=0
cc_757 N_A_33_81#_c_1376_n N_VGND_c_1416_n 0.0130139f $X=1.225 $Y=0.35 $X2=0
+ $Y2=0
cc_758 N_A_33_81#_c_1372_n N_VGND_c_1423_n 0.00767437f $X=0.29 $Y=0.615 $X2=0
+ $Y2=0
cc_759 N_A_33_81#_c_1375_n N_VGND_c_1424_n 0.0401682f $X=1.895 $Y=0.35 $X2=0
+ $Y2=0
cc_760 N_A_33_81#_c_1376_n N_VGND_c_1424_n 0.0115119f $X=1.225 $Y=0.35 $X2=0
+ $Y2=0
cc_761 N_A_33_81#_c_1377_n N_VGND_c_1424_n 0.0212546f $X=2.06 $Y=0.35 $X2=0
+ $Y2=0
cc_762 N_A_33_81#_c_1372_n N_VGND_c_1428_n 0.00885121f $X=0.29 $Y=0.615 $X2=0
+ $Y2=0
cc_763 N_A_33_81#_c_1373_n N_VGND_c_1428_n 0.0122144f $X=1.055 $Y=0.9 $X2=0
+ $Y2=0
cc_764 N_A_33_81#_c_1375_n N_VGND_c_1428_n 0.0241404f $X=1.895 $Y=0.35 $X2=0
+ $Y2=0
cc_765 N_A_33_81#_c_1376_n N_VGND_c_1428_n 0.00658819f $X=1.225 $Y=0.35 $X2=0
+ $Y2=0
cc_766 N_A_33_81#_c_1377_n N_VGND_c_1428_n 0.0112078f $X=2.06 $Y=0.35 $X2=0
+ $Y2=0
cc_767 N_VGND_c_1428_n N_A_710_117#_M1012_s 0.00215176f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_768 N_VGND_c_1417_n N_A_710_117#_c_1520_n 0.038903f $X=3.155 $Y=0.805 $X2=0
+ $Y2=0
cc_769 N_VGND_c_1417_n N_A_710_117#_c_1521_n 0.0155356f $X=3.155 $Y=0.805 $X2=0
+ $Y2=0
cc_770 N_VGND_c_1425_n N_A_710_117#_c_1521_n 0.0201532f $X=5.39 $Y=0 $X2=0 $Y2=0
cc_771 N_VGND_c_1428_n N_A_710_117#_c_1521_n 0.0101278f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_772 N_VGND_c_1425_n N_A_710_117#_c_1523_n 0.089516f $X=5.39 $Y=0 $X2=0 $Y2=0
cc_773 N_VGND_c_1428_n N_A_710_117#_c_1523_n 0.0524213f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_774 N_VGND_c_1428_n N_A_879_117#_M1015_d 0.00224755f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_775 N_VGND_M1012_d N_A_879_117#_c_1546_n 0.0025308f $X=5.345 $Y=0.235 $X2=0
+ $Y2=0
cc_776 N_VGND_c_1418_n N_A_879_117#_c_1546_n 0.0199842f $X=5.555 $Y=0.36 $X2=0
+ $Y2=0
cc_777 N_VGND_c_1419_n N_A_879_117#_c_1546_n 0.0111203f $X=6.655 $Y=0.76 $X2=0
+ $Y2=0
cc_778 N_VGND_c_1421_n N_A_879_117#_c_1546_n 0.00250027f $X=6.49 $Y=0 $X2=0
+ $Y2=0
cc_779 N_VGND_c_1425_n N_A_879_117#_c_1546_n 0.00243439f $X=5.39 $Y=0 $X2=0
+ $Y2=0
cc_780 N_VGND_c_1428_n N_A_879_117#_c_1546_n 0.0109239f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_781 N_VGND_c_1419_n N_A_879_117#_c_1547_n 0.0190898f $X=6.655 $Y=0.76 $X2=0
+ $Y2=0
cc_782 N_VGND_c_1421_n N_A_879_117#_c_1547_n 0.0159076f $X=6.49 $Y=0 $X2=0 $Y2=0
cc_783 N_VGND_c_1428_n N_A_879_117#_c_1547_n 0.0102681f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_784 N_A_710_117#_M1012_s N_A_879_117#_c_1546_n 0.00216977f $X=4.93 $Y=0.235
+ $X2=0 $Y2=0
cc_785 N_A_710_117#_c_1522_n N_A_879_117#_c_1546_n 0.019398f $X=5.055 $Y=0.38
+ $X2=0 $Y2=0
cc_786 N_A_710_117#_c_1523_n N_A_879_117#_c_1546_n 0.012046f $X=4.89 $Y=0.365
+ $X2=0 $Y2=0
cc_787 N_A_710_117#_c_1523_n N_A_879_117#_c_1548_n 0.0218248f $X=4.89 $Y=0.365
+ $X2=0 $Y2=0
