# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__bufkapwr_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.440000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.345000 1.015000 1.750000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.445200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.300000 0.430000 0.635000 ;
        RECT 0.085000 0.635000 0.255000 1.525000 ;
        RECT 0.085000 1.525000 0.395000 3.075000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.690000 1.370000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.440000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.440000 0.085000 ;
      RECT 0.000000  3.245000 1.440000 3.415000 ;
      RECT 0.425000  0.805000 1.355000 1.135000 ;
      RECT 0.565000  1.920000 0.825000 3.075000 ;
      RECT 0.600000  0.085000 0.875000 0.635000 ;
      RECT 0.995000  1.920000 1.355000 3.075000 ;
      RECT 1.045000  0.300000 1.355000 0.805000 ;
      RECT 1.185000  1.135000 1.355000 1.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.615000  2.725000 0.785000 2.895000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
  END
END sky130_fd_sc_lp__bufkapwr_1
END LIBRARY
