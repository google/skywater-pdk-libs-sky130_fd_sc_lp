# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__sdfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.015000 1.530000 2.255000 1.840000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.925000 0.325000 14.315000 1.125000 ;
        RECT 14.035000 1.850000 14.315000 3.075000 ;
        RECT 14.065000 1.125000 14.315000 1.850000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.170000 0.620000 1.840000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.430000 0.265000 3.275000 0.640000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.835000 0.265000 10.620000 0.640000 ;
        RECT 10.450000 0.640000 10.620000 1.585000 ;
        RECT 10.450000 1.585000 11.660000 1.765000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.950000 0.780000 4.285000 1.825000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.095000  2.010000  2.185000 2.180000 ;
      RECT  0.095000  2.180000  0.390000 2.700000 ;
      RECT  0.165000  0.085000  0.495000 1.000000 ;
      RECT  0.560000  2.350000  0.855000 3.245000 ;
      RECT  0.955000  0.685000  1.285000 1.190000 ;
      RECT  0.955000  1.190000  2.595000 1.360000 ;
      RECT  1.370000  2.350000  1.700000 2.450000 ;
      RECT  1.370000  2.450000  3.055000 2.640000 ;
      RECT  1.745000  0.085000  2.015000 1.015000 ;
      RECT  1.855000  2.180000  2.185000 2.280000 ;
      RECT  2.215000  0.810000  3.025000 1.020000 ;
      RECT  2.375000  2.810000  2.705000 3.245000 ;
      RECT  2.425000  1.360000  2.595000 2.450000 ;
      RECT  2.765000  1.020000  3.025000 1.620000 ;
      RECT  2.765000  1.620000  3.440000 1.790000 ;
      RECT  2.885000  2.640000  3.055000 2.895000 ;
      RECT  2.885000  2.895000  4.060000 3.065000 ;
      RECT  3.225000  1.790000  3.440000 2.725000 ;
      RECT  3.470000  0.280000  3.780000 0.610000 ;
      RECT  3.610000  0.610000  3.780000 1.995000 ;
      RECT  3.610000  1.995000  4.835000 2.185000 ;
      RECT  3.610000  2.185000  4.025000 2.315000 ;
      RECT  3.890000  2.495000  5.550000 2.525000 ;
      RECT  3.890000  2.525000  4.570000 2.665000 ;
      RECT  3.890000  2.665000  4.060000 2.895000 ;
      RECT  3.950000  0.085000  4.200000 0.610000 ;
      RECT  4.240000  2.845000  4.570000 3.245000 ;
      RECT  4.370000  0.265000  5.550000 0.435000 ;
      RECT  4.370000  0.435000  4.660000 0.610000 ;
      RECT  4.400000  2.355000  5.550000 2.495000 ;
      RECT  4.740000  2.695000  5.000000 2.865000 ;
      RECT  4.740000  2.865000  6.250000 3.035000 ;
      RECT  4.870000  0.605000  5.200000 0.805000 ;
      RECT  5.030000  0.805000  5.200000 2.295000 ;
      RECT  5.030000  2.295000  5.550000 2.355000 ;
      RECT  5.200000  2.525000  5.550000 2.690000 ;
      RECT  5.370000  0.435000  5.550000 1.845000 ;
      RECT  5.720000  0.325000  5.920000 0.725000 ;
      RECT  5.720000  0.725000  5.900000 1.245000 ;
      RECT  5.720000  1.245000  8.695000 1.425000 ;
      RECT  5.720000  1.425000  5.900000 2.690000 ;
      RECT  6.080000  1.595000  6.410000 1.945000 ;
      RECT  6.080000  1.945000  7.060000 2.115000 ;
      RECT  6.080000  2.115000  6.250000 2.865000 ;
      RECT  6.440000  0.085000  6.770000 0.665000 ;
      RECT  6.440000  2.370000  6.720000 3.245000 ;
      RECT  6.470000  0.835000  7.315000 1.075000 ;
      RECT  6.620000  1.595000  7.460000 1.775000 ;
      RECT  6.890000  2.115000  7.060000 2.840000 ;
      RECT  6.890000  2.840000  7.800000 3.010000 ;
      RECT  7.055000  0.660000  7.315000 0.835000 ;
      RECT  7.230000  1.775000  7.460000 2.670000 ;
      RECT  7.485000  0.085000  7.655000 0.820000 ;
      RECT  7.485000  0.820000  8.855000 1.010000 ;
      RECT  7.630000  1.815000  9.470000 1.985000 ;
      RECT  7.630000  1.985000  7.800000 2.840000 ;
      RECT  7.970000  2.155000  8.310000 3.245000 ;
      RECT  8.365000  1.425000  8.695000 1.645000 ;
      RECT  8.490000  2.155000  8.820000 2.285000 ;
      RECT  8.490000  2.285000 10.410000 2.455000 ;
      RECT  8.490000  2.455000  8.820000 2.755000 ;
      RECT  9.010000  2.625000  9.340000 2.795000 ;
      RECT  9.010000  2.795000 10.920000 2.965000 ;
      RECT  9.140000  1.985000  9.470000 2.105000 ;
      RECT  9.640000  0.810000 10.280000 1.935000 ;
      RECT  9.640000  1.935000 12.340000 2.115000 ;
      RECT 10.080000  2.455000 10.410000 2.625000 ;
      RECT 10.630000  2.465000 10.920000 2.795000 ;
      RECT 10.790000  1.235000 12.770000 1.415000 ;
      RECT 11.090000  2.465000 11.350000 3.245000 ;
      RECT 11.495000  0.085000 11.825000 0.995000 ;
      RECT 11.520000  2.115000 12.340000 2.255000 ;
      RECT 11.520000  2.255000 11.760000 2.795000 ;
      RECT 11.995000  0.665000 12.325000 1.235000 ;
      RECT 12.010000  2.465000 12.340000 3.245000 ;
      RECT 12.090000  1.585000 12.340000 1.935000 ;
      RECT 12.510000  1.415000 12.770000 2.795000 ;
      RECT 12.950000  0.810000 13.230000 1.295000 ;
      RECT 12.950000  1.295000 13.895000 1.625000 ;
      RECT 12.950000  1.625000 13.255000 2.495000 ;
      RECT 13.400000  0.085000 13.755000 1.125000 ;
      RECT 13.425000  1.815000 13.865000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfstp_1
END LIBRARY
