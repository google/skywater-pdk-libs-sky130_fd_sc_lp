* File: sky130_fd_sc_lp__a211oi_1.pxi.spice
* Created: Fri Aug 28 09:48:16 2020
* 
x_PM_SKY130_FD_SC_LP__A211OI_1%A2 N_A2_c_48_n N_A2_M1002_g N_A2_M1006_g A2 A2
+ N_A2_c_51_n PM_SKY130_FD_SC_LP__A211OI_1%A2
x_PM_SKY130_FD_SC_LP__A211OI_1%A1 N_A1_M1007_g N_A1_M1000_g A1 A1 A1 A1
+ N_A1_c_78_n N_A1_c_79_n PM_SKY130_FD_SC_LP__A211OI_1%A1
x_PM_SKY130_FD_SC_LP__A211OI_1%B1 N_B1_M1001_g N_B1_M1003_g B1 N_B1_c_117_n
+ PM_SKY130_FD_SC_LP__A211OI_1%B1
x_PM_SKY130_FD_SC_LP__A211OI_1%C1 N_C1_M1005_g N_C1_M1004_g C1 N_C1_c_151_n
+ N_C1_c_152_n PM_SKY130_FD_SC_LP__A211OI_1%C1
x_PM_SKY130_FD_SC_LP__A211OI_1%A_27_367# N_A_27_367#_M1006_s N_A_27_367#_M1000_d
+ N_A_27_367#_c_177_n N_A_27_367#_c_178_n N_A_27_367#_c_183_n
+ N_A_27_367#_c_189_n N_A_27_367#_c_194_p PM_SKY130_FD_SC_LP__A211OI_1%A_27_367#
x_PM_SKY130_FD_SC_LP__A211OI_1%VPWR N_VPWR_M1006_d N_VPWR_c_200_n VPWR
+ N_VPWR_c_201_n N_VPWR_c_202_n N_VPWR_c_199_n N_VPWR_c_204_n
+ PM_SKY130_FD_SC_LP__A211OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A211OI_1%Y N_Y_M1007_d N_Y_M1005_d N_Y_M1004_d N_Y_c_228_n
+ N_Y_c_238_n N_Y_c_229_n N_Y_c_230_n N_Y_c_231_n Y Y Y N_Y_c_233_n N_Y_c_232_n
+ PM_SKY130_FD_SC_LP__A211OI_1%Y
x_PM_SKY130_FD_SC_LP__A211OI_1%VGND N_VGND_M1002_s N_VGND_M1001_d N_VGND_c_272_n
+ N_VGND_c_273_n N_VGND_c_274_n VGND N_VGND_c_275_n N_VGND_c_276_n
+ N_VGND_c_277_n N_VGND_c_278_n PM_SKY130_FD_SC_LP__A211OI_1%VGND
cc_1 VNB N_A2_c_48_n 0.0219236f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.21
cc_2 VNB N_A2_M1006_g 0.00763498f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB A2 0.0194233f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A2_c_51_n 0.0447002f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.375
cc_5 VNB N_A1_M1000_g 0.00703869f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_6 VNB A1 0.00102607f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB A1 0.00835749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A1_c_78_n 0.0307167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_c_79_n 0.0162041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_M1001_g 0.0257721f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.665
cc_11 VNB B1 0.00604739f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_B1_c_117_n 0.0217959f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.375
cc_13 VNB N_C1_M1005_g 0.0272173f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.665
cc_14 VNB N_C1_M1004_g 0.00176076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_C1_c_151_n 0.0473945f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.375
cc_16 VNB N_C1_c_152_n 0.0030216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_199_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.665
cc_18 VNB N_Y_c_228_n 0.0045273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_229_n 0.0242382f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.295
cc_20 VNB N_Y_c_230_n 0.00429407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_231_n 0.0453703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_232_n 0.0276036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_272_n 0.0104415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_273_n 0.0342756f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_25 VNB N_VGND_c_274_n 0.00319039f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.375
cc_26 VNB N_VGND_c_275_n 0.0287086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_276_n 0.0313707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_277_n 0.188336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_278_n 0.00529002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_A2_M1006_g 0.0273657f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_31 VPB A2 0.00693541f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_32 VPB N_A1_M1000_g 0.0227225f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_33 VPB A1 0.00452104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_B1_M1003_g 0.0187037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB B1 0.0107494f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_36 VPB N_B1_c_117_n 0.00624595f $X=-0.19 $Y=1.655 $X2=0.3 $Y2=1.375
cc_37 VPB N_C1_M1004_g 0.0239008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_C1_c_152_n 0.00387157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_367#_c_177_n 0.00754068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_27_367#_c_178_n 0.0377822f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_41 VPB N_VPWR_c_200_n 0.0055721f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_42 VPB N_VPWR_c_201_n 0.0175363f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_202_n 0.053924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_199_n 0.0488467f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.665
cc_45 VPB N_VPWR_c_204_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_Y_c_233_n 0.0814687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_Y_c_232_n 0.0157833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 N_A2_c_51_n N_A1_M1000_g 0.0271003f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_49 N_A2_c_48_n A1 0.00505292f $X=0.475 $Y=1.21 $X2=0 $Y2=0
cc_50 N_A2_c_48_n A1 0.0049398f $X=0.475 $Y=1.21 $X2=0 $Y2=0
cc_51 A2 A1 0.0439193f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_52 A2 N_A1_c_78_n 2.39011e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_53 N_A2_c_51_n N_A1_c_78_n 0.0424086f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_54 N_A2_c_48_n N_A1_c_79_n 0.0424086f $X=0.475 $Y=1.21 $X2=0 $Y2=0
cc_55 N_A2_M1006_g N_A_27_367#_c_177_n 2.7414e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_56 A2 N_A_27_367#_c_177_n 0.0257895f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_A2_c_51_n N_A_27_367#_c_177_n 0.00115827f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_58 N_A2_M1006_g N_A_27_367#_c_178_n 0.0130023f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A2_M1006_g N_A_27_367#_c_183_n 0.0166238f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_60 A2 N_A_27_367#_c_183_n 0.00101367f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_A2_M1006_g N_VPWR_c_200_n 0.00419107f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_62 N_A2_M1006_g N_VPWR_c_201_n 0.00571722f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_63 N_A2_M1006_g N_VPWR_c_199_n 0.0114807f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A2_c_48_n N_VGND_c_273_n 0.0184296f $X=0.475 $Y=1.21 $X2=0 $Y2=0
cc_65 A2 N_VGND_c_273_n 0.0257902f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A2_c_51_n N_VGND_c_273_n 0.00192467f $X=0.475 $Y=1.375 $X2=0 $Y2=0
cc_67 N_A2_c_48_n N_VGND_c_275_n 0.00477554f $X=0.475 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A2_c_48_n N_VGND_c_277_n 0.00814835f $X=0.475 $Y=1.21 $X2=0 $Y2=0
cc_69 A1 N_B1_M1001_g 4.40849e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_70 A1 N_B1_M1001_g 8.30097e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_71 N_A1_c_78_n N_B1_M1001_g 0.0149167f $X=0.925 $Y=1.36 $X2=0 $Y2=0
cc_72 N_A1_c_79_n N_B1_M1001_g 0.0179793f $X=0.925 $Y=1.195 $X2=0 $Y2=0
cc_73 N_A1_M1000_g N_B1_M1003_g 0.0260856f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_74 A1 B1 0.0224004f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_75 N_A1_c_78_n B1 0.00341332f $X=0.925 $Y=1.36 $X2=0 $Y2=0
cc_76 N_A1_M1000_g N_B1_c_117_n 0.0149167f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A1_M1000_g N_A_27_367#_c_178_n 7.67736e-19 $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A1_M1000_g N_A_27_367#_c_183_n 0.0189093f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_79 A1 N_A_27_367#_c_183_n 0.0266579f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_80 N_A1_c_78_n N_A_27_367#_c_183_n 6.66716e-19 $X=0.925 $Y=1.36 $X2=0 $Y2=0
cc_81 N_A1_M1000_g N_VPWR_c_200_n 0.00419107f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A1_M1000_g N_VPWR_c_202_n 0.00585385f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A1_M1000_g N_VPWR_c_199_n 0.0112404f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_84 A1 N_Y_c_228_n 0.0229057f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_85 N_A1_c_78_n N_Y_c_228_n 0.00339685f $X=0.925 $Y=1.36 $X2=0 $Y2=0
cc_86 N_A1_c_79_n N_Y_c_228_n 0.00305175f $X=0.925 $Y=1.195 $X2=0 $Y2=0
cc_87 A1 N_Y_c_238_n 0.0317914f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_88 N_A1_c_79_n N_Y_c_238_n 0.00503521f $X=0.925 $Y=1.195 $X2=0 $Y2=0
cc_89 N_A1_c_79_n N_VGND_c_273_n 0.00201933f $X=0.925 $Y=1.195 $X2=0 $Y2=0
cc_90 A1 N_VGND_c_275_n 0.00821604f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_91 N_A1_c_79_n N_VGND_c_275_n 0.00463154f $X=0.925 $Y=1.195 $X2=0 $Y2=0
cc_92 A1 N_VGND_c_277_n 0.00858173f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_93 N_A1_c_79_n N_VGND_c_277_n 0.00792059f $X=0.925 $Y=1.195 $X2=0 $Y2=0
cc_94 A1 A_110_49# 0.00120322f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_95 N_B1_M1001_g N_C1_M1005_g 0.0252441f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_96 N_B1_M1003_g N_C1_M1004_g 0.0562297f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_97 B1 N_C1_c_151_n 0.00339844f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_98 N_B1_c_117_n N_C1_c_151_n 0.0562297f $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_99 B1 N_C1_c_152_n 0.0333955f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_100 N_B1_c_117_n N_C1_c_152_n 3.01852e-19 $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_101 B1 N_A_27_367#_c_189_n 0.015315f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_102 N_B1_c_117_n N_A_27_367#_c_189_n 8.9513e-19 $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_103 N_B1_M1003_g N_VPWR_c_202_n 0.00585385f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_104 N_B1_M1003_g N_VPWR_c_199_n 0.0109726f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_105 N_B1_M1001_g N_Y_c_228_n 0.00721761f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_106 B1 N_Y_c_228_n 0.00720625f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_107 N_B1_M1001_g N_Y_c_238_n 0.00688678f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_108 N_B1_M1001_g N_Y_c_230_n 0.00796116f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_109 B1 N_Y_c_230_n 0.0352623f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_110 N_B1_c_117_n N_Y_c_230_n 0.00463193f $X=1.465 $Y=1.51 $X2=0 $Y2=0
cc_111 N_B1_M1003_g N_Y_c_233_n 0.00320795f $X=1.555 $Y=2.465 $X2=0 $Y2=0
cc_112 N_B1_M1001_g N_VGND_c_274_n 0.0080598f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_113 N_B1_M1001_g N_VGND_c_275_n 0.00501942f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_114 N_B1_M1001_g N_VGND_c_277_n 0.00950163f $X=1.375 $Y=0.665 $X2=0 $Y2=0
cc_115 N_C1_M1004_g N_VPWR_c_202_n 0.0054895f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_116 N_C1_M1004_g N_VPWR_c_199_n 0.0111524f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_117 N_C1_M1005_g N_Y_c_228_n 2.83863e-19 $X=1.915 $Y=0.665 $X2=0 $Y2=0
cc_118 N_C1_M1005_g N_Y_c_230_n 0.0188767f $X=1.915 $Y=0.665 $X2=0 $Y2=0
cc_119 N_C1_c_151_n N_Y_c_230_n 0.00748166f $X=2.135 $Y=1.46 $X2=0 $Y2=0
cc_120 N_C1_c_152_n N_Y_c_230_n 0.0267705f $X=2.135 $Y=1.46 $X2=0 $Y2=0
cc_121 N_C1_M1004_g N_Y_c_233_n 0.0238722f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_122 N_C1_c_151_n N_Y_c_233_n 0.00166713f $X=2.135 $Y=1.46 $X2=0 $Y2=0
cc_123 N_C1_c_152_n N_Y_c_233_n 0.0262213f $X=2.135 $Y=1.46 $X2=0 $Y2=0
cc_124 N_C1_M1005_g N_Y_c_232_n 0.00304964f $X=1.915 $Y=0.665 $X2=0 $Y2=0
cc_125 N_C1_M1004_g N_Y_c_232_n 0.00385685f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_126 N_C1_c_151_n N_Y_c_232_n 0.00396834f $X=2.135 $Y=1.46 $X2=0 $Y2=0
cc_127 N_C1_c_152_n N_Y_c_232_n 0.0303187f $X=2.135 $Y=1.46 $X2=0 $Y2=0
cc_128 N_C1_M1005_g N_VGND_c_274_n 0.0105132f $X=1.915 $Y=0.665 $X2=0 $Y2=0
cc_129 N_C1_M1005_g N_VGND_c_276_n 0.0053507f $X=1.915 $Y=0.665 $X2=0 $Y2=0
cc_130 N_C1_M1005_g N_VGND_c_277_n 0.0104858f $X=1.915 $Y=0.665 $X2=0 $Y2=0
cc_131 N_A_27_367#_c_183_n N_VPWR_M1006_d 0.00599733f $X=1.125 $Y=2.015
+ $X2=-0.19 $Y2=1.655
cc_132 N_A_27_367#_c_183_n N_VPWR_c_200_n 0.022455f $X=1.125 $Y=2.015 $X2=0
+ $Y2=0
cc_133 N_A_27_367#_c_178_n N_VPWR_c_201_n 0.0200241f $X=0.26 $Y=2.91 $X2=0 $Y2=0
cc_134 N_A_27_367#_c_194_p N_VPWR_c_202_n 0.0212513f $X=1.29 $Y=2.455 $X2=0
+ $Y2=0
cc_135 N_A_27_367#_M1006_s N_VPWR_c_199_n 0.00215158f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_136 N_A_27_367#_M1000_d N_VPWR_c_199_n 0.00526034f $X=1.09 $Y=1.835 $X2=0
+ $Y2=0
cc_137 N_A_27_367#_c_178_n N_VPWR_c_199_n 0.0120544f $X=0.26 $Y=2.91 $X2=0 $Y2=0
cc_138 N_A_27_367#_c_194_p N_VPWR_c_199_n 0.0127519f $X=1.29 $Y=2.455 $X2=0
+ $Y2=0
cc_139 N_VPWR_c_199_n A_326_367# 0.00899413f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_140 N_VPWR_c_199_n N_Y_M1004_d 0.00215158f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_141 N_VPWR_c_202_n N_Y_c_233_n 0.0561732f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_142 N_VPWR_c_199_n N_Y_c_233_n 0.031619f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_143 N_Y_c_230_n N_VGND_M1001_d 0.0034757f $X=2.02 $Y=1.03 $X2=0 $Y2=0
cc_144 N_Y_c_238_n N_VGND_c_273_n 0.00364535f $X=1.13 $Y=0.42 $X2=0 $Y2=0
cc_145 N_Y_c_228_n N_VGND_c_274_n 0.00210872f $X=1.182 $Y=0.798 $X2=0 $Y2=0
cc_146 N_Y_c_238_n N_VGND_c_274_n 0.0421595f $X=1.13 $Y=0.42 $X2=0 $Y2=0
cc_147 N_Y_c_230_n N_VGND_c_274_n 0.0220444f $X=2.02 $Y=1.03 $X2=0 $Y2=0
cc_148 N_Y_c_238_n N_VGND_c_275_n 0.0213278f $X=1.13 $Y=0.42 $X2=0 $Y2=0
cc_149 N_Y_c_229_n N_VGND_c_276_n 0.0182456f $X=2.13 $Y=0.42 $X2=0 $Y2=0
cc_150 N_Y_M1007_d N_VGND_c_277_n 0.00681569f $X=0.91 $Y=0.245 $X2=0 $Y2=0
cc_151 N_Y_M1005_d N_VGND_c_277_n 0.00316663f $X=1.99 $Y=0.245 $X2=0 $Y2=0
cc_152 N_Y_c_238_n N_VGND_c_277_n 0.0126562f $X=1.13 $Y=0.42 $X2=0 $Y2=0
cc_153 N_Y_c_229_n N_VGND_c_277_n 0.0105923f $X=2.13 $Y=0.42 $X2=0 $Y2=0
cc_154 N_VGND_c_277_n A_110_49# 0.00337783f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
