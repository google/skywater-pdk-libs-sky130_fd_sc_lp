* File: sky130_fd_sc_lp__ha_0.pex.spice
* Created: Fri Aug 28 10:36:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__HA_0%A_80_60# 1 2 9 12 15 17 19 21 22 24 28 29 34
c68 28 0 6.17501e-20 $X=0.59 $Y=1.76
c69 19 0 7.08146e-21 $X=1.06 $Y=1.595
r70 31 34 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=0.445
+ $X2=1.225 $Y2=0.445
r71 28 37 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.76
+ $X2=0.577 $Y2=1.595
r72 27 29 11.0058 $w=5.21e-07 $l=4.7e-07 $layer=LI1_cond $X=0.59 $Y=1.93
+ $X2=1.06 $Y2=1.93
r73 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.76 $X2=0.59 $Y2=1.76
r74 22 24 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=1.415 $Y=2.665
+ $X2=1.675 $Y2=2.665
r75 21 22 7.01204 $w=3.3e-07 $l=2.17991e-07 $layer=LI1_cond $X=1.292 $Y=2.5
+ $X2=1.415 $Y2=2.665
r76 20 29 5.43263 $w=5.21e-07 $l=4.35827e-07 $layer=LI1_cond $X=1.292 $Y=2.265
+ $X2=1.06 $Y2=1.93
r77 20 21 11.054 $w=2.43e-07 $l=2.35e-07 $layer=LI1_cond $X=1.292 $Y=2.265
+ $X2=1.292 $Y2=2.5
r78 19 29 7.41575 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.06 $Y=1.595
+ $X2=1.06 $Y2=1.93
r79 18 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=0.61
+ $X2=1.06 $Y2=0.445
r80 18 19 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=1.06 $Y=0.61
+ $X2=1.06 $Y2=1.595
r81 15 17 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.57 $Y=2.775
+ $X2=0.57 $Y2=2.265
r82 12 17 38.9865 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.577 $Y=2.088
+ $X2=0.577 $Y2=2.265
r83 11 28 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.577 $Y=1.772
+ $X2=0.577 $Y2=1.76
r84 11 12 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.577 $Y=1.772
+ $X2=0.577 $Y2=2.088
r85 9 37 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=0.475 $Y=0.64
+ $X2=0.475 $Y2=1.595
r86 2 24 300 $w=1.7e-07 $l=6.00895e-07 $layer=licon1_PDIFF $count=2 $X=1.17
+ $Y=2.455 $X2=1.675 $Y2=2.665
r87 1 34 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.235 $X2=1.225 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__HA_0%A_204_315# 1 2 9 13 16 19 23 28 32 35 36 38 39
+ 42 47 50 52 53
c109 39 0 6.17501e-20 $X=1.575 $Y=1.65
c110 36 0 1.08071e-19 $X=1.41 $Y=1.22
r111 52 53 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.48 $Y=2.665
+ $X2=3.48 $Y2=2.5
r112 50 57 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=4.202 $Y=1.76
+ $X2=4.202 $Y2=1.595
r113 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.17
+ $Y=1.76 $X2=4.17 $Y2=1.76
r114 47 49 15.6753 $w=5.02e-07 $l=6.45e-07 $layer=LI1_cond $X=3.525 $Y=1.915
+ $X2=4.17 $Y2=1.915
r115 44 47 7.18174 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=3.525 $Y=2.265
+ $X2=3.525 $Y2=1.915
r116 44 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.525 $Y=2.265
+ $X2=3.525 $Y2=2.5
r117 40 47 5.2251 $w=5.02e-07 $l=4.44691e-07 $layer=LI1_cond $X=3.31 $Y=1.565
+ $X2=3.525 $Y2=1.915
r118 40 42 13.5556 $w=5.98e-07 $l=6.8e-07 $layer=LI1_cond $X=3.31 $Y=1.565
+ $X2=3.31 $Y2=0.885
r119 38 40 13.0009 $w=5.02e-07 $l=3.39853e-07 $layer=LI1_cond $X=3.01 $Y=1.65
+ $X2=3.31 $Y2=1.565
r120 38 39 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=3.01 $Y=1.65
+ $X2=1.575 $Y2=1.65
r121 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.41
+ $Y=1.22 $X2=1.41 $Y2=1.22
r122 33 39 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.445 $Y=1.565
+ $X2=1.575 $Y2=1.65
r123 33 35 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=1.445 $Y=1.565
+ $X2=1.445 $Y2=1.22
r124 31 36 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.055
+ $X2=1.41 $Y2=1.22
r125 28 36 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.41 $Y=1.575
+ $X2=1.41 $Y2=1.22
r126 25 28 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.095 $Y=1.65
+ $X2=1.41 $Y2=1.65
r127 23 57 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.325 $Y=0.885
+ $X2=4.325 $Y2=1.595
r128 19 32 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.205 $Y=2.775
+ $X2=4.205 $Y2=2.265
r129 16 32 39.0652 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=4.202 $Y=2.068
+ $X2=4.202 $Y2=2.265
r130 15 50 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=4.202 $Y=1.792
+ $X2=4.202 $Y2=1.76
r131 15 16 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=4.202 $Y=1.792
+ $X2=4.202 $Y2=2.068
r132 13 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.46 $Y=0.445
+ $X2=1.46 $Y2=1.055
r133 7 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.095 $Y=1.725
+ $X2=1.095 $Y2=1.65
r134 7 9 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.095 $Y=1.725 $X2=1.095
+ $Y2=2.665
r135 2 52 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=2.455 $X2=3.445 $Y2=2.665
r136 1 42 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.675 $X2=3.115 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LP__HA_0%B 3 7 10 13 15 17 18 19 22 24 25 26 27 39
c71 22 0 1.58215e-19 $X=3.36 $Y=1.28
c72 15 0 1.04272e-19 $X=3.36 $Y=1.205
c73 3 0 7.08146e-21 $X=1.89 $Y=0.445
r74 36 39 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.04 $Y=2 $X2=3.23
+ $Y2=2
r75 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.76
+ $Y=2.13 $X2=1.76 $Y2=2.13
r76 27 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04 $Y=2
+ $X2=3.04 $Y2=2
r77 26 27 12.131 $w=3.78e-07 $l=4e-07 $layer=LI1_cond $X=2.64 $Y=2.105 $X2=3.04
+ $Y2=2.105
r78 25 26 14.5572 $w=3.78e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.105
+ $X2=2.64 $Y2=2.105
r79 25 34 12.131 $w=3.78e-07 $l=4e-07 $layer=LI1_cond $X=2.16 $Y=2.105 $X2=1.76
+ $Y2=2.105
r80 24 34 2.4262 $w=3.78e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=2.105 $X2=1.76
+ $Y2=2.105
r81 20 22 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=3.23 $Y=1.28
+ $X2=3.36 $Y2=1.28
r82 18 33 8.03333 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.815 $Y=2.13
+ $X2=1.76 $Y2=2.13
r83 18 19 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.815 $Y=2.13
+ $X2=1.89 $Y2=2.13
r84 15 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.36 $Y=1.205
+ $X2=3.36 $Y2=1.28
r85 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.36 $Y=1.205
+ $X2=3.36 $Y2=0.885
r86 11 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=2.165
+ $X2=3.23 $Y2=2
r87 11 13 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.23 $Y=2.165 $X2=3.23
+ $Y2=2.665
r88 10 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.835
+ $X2=3.23 $Y2=2
r89 9 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.23 $Y=1.355
+ $X2=3.23 $Y2=1.28
r90 9 10 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.23 $Y=1.355
+ $X2=3.23 $Y2=1.835
r91 5 19 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=2.295
+ $X2=1.89 $Y2=2.13
r92 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.89 $Y=2.295 $X2=1.89
+ $Y2=2.665
r93 1 19 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.965
+ $X2=1.89 $Y2=2.13
r94 1 3 779.404 $w=1.5e-07 $l=1.52e-06 $layer=POLY_cond $X=1.89 $Y=1.965
+ $X2=1.89 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__HA_0%A 3 7 10 11 12 15 20 22 23 25 26 27
c69 27 0 2.62487e-19 $X=2.64 $Y=1.295
r70 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.22 $X2=2.48 $Y2=1.22
r71 27 32 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.64 $Y=1.22 $X2=2.48
+ $Y2=1.22
r72 26 32 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.16 $Y=1.22
+ $X2=2.48 $Y2=1.22
r73 24 25 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=3.69 $Y=1.565
+ $X2=3.69 $Y2=1.715
r74 23 31 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=2.735 $Y=1.22
+ $X2=2.48 $Y2=1.22
r75 21 31 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=2.395 $Y=1.22
+ $X2=2.48 $Y2=1.22
r76 21 22 5.03009 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.395 $Y=1.22
+ $X2=2.3 $Y2=1.22
r77 20 24 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.72 $Y=0.885
+ $X2=3.72 $Y2=1.565
r78 17 20 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.72 $Y=0.335
+ $X2=3.72 $Y2=0.885
r79 15 25 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.66 $Y=2.665
+ $X2=3.66 $Y2=1.715
r80 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.645 $Y=0.26
+ $X2=3.72 $Y2=0.335
r81 11 12 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.645 $Y=0.26
+ $X2=2.885 $Y2=0.26
r82 10 23 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.81 $Y=1.055
+ $X2=2.735 $Y2=1.22
r83 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.81 $Y=0.335
+ $X2=2.885 $Y2=0.26
r84 9 10 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.81 $Y=0.335
+ $X2=2.81 $Y2=1.055
r85 5 22 37.0704 $w=1.5e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.32 $Y=1.055
+ $X2=2.3 $Y2=1.22
r86 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.32 $Y=1.055 $X2=2.32
+ $Y2=0.445
r87 1 22 37.0704 $w=1.5e-07 $l=1.74714e-07 $layer=POLY_cond $X=2.28 $Y=1.385
+ $X2=2.3 $Y2=1.22
r88 1 3 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=2.28 $Y=1.385 $X2=2.28
+ $Y2=2.665
.ends

.subckt PM_SKY130_FD_SC_LP__HA_0%SUM 1 2 7 8 9 10 11 12 13 39 43
r21 43 44 5.12173 $w=4.03e-07 $l=1.05e-07 $layer=LI1_cond $X=0.297 $Y=2.6
+ $X2=0.297 $Y2=2.495
r22 22 39 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.26 $Y=1.26
+ $X2=0.26 $Y2=1.295
r23 13 43 4.97969 $w=4.03e-07 $l=1.75e-07 $layer=LI1_cond $X=0.297 $Y=2.775
+ $X2=0.297 $Y2=2.6
r24 12 44 4.50956 $w=2.28e-07 $l=9e-08 $layer=LI1_cond $X=0.21 $Y=2.405 $X2=0.21
+ $Y2=2.495
r25 11 12 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=2.035
+ $X2=0.21 $Y2=2.405
r26 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=2.035
r27 10 41 12.0255 $w=2.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=1.425
r28 9 41 4.73726 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.26 $Y=1.32
+ $X2=0.26 $Y2=1.425
r29 9 39 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.26 $Y=1.32
+ $X2=0.26 $Y2=1.295
r30 9 22 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.26 $Y=1.235
+ $X2=0.26 $Y2=1.26
r31 8 9 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.26 $Y=0.925 $X2=0.26
+ $Y2=1.235
r32 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.555 $X2=0.26
+ $Y2=0.925
r33 2 43 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.21
+ $Y=2.455 $X2=0.335 $Y2=2.6
r34 1 7 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.43 $X2=0.26 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_LP__HA_0%VPWR 1 2 3 14 18 21 22 23 38 39 42 47 50
r55 49 50 12.3619 $w=9.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=2.957
+ $X2=3.18 $Y2=2.957
r56 45 49 5 $w=9.13e-07 $l=3.75e-07 $layer=LI1_cond $X=2.64 $Y=2.957 $X2=3.015
+ $Y2=2.957
r57 45 47 14.2952 $w=9.13e-07 $l=3.1e-07 $layer=LI1_cond $X=2.64 $Y=2.957
+ $X2=2.33 $Y2=2.957
r58 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r62 36 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 35 50 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=3.18
+ $Y2=3.33
r64 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r65 31 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.33 $Y2=3.33
r66 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r67 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r68 29 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 28 31 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r70 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r71 26 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=0.835
+ $Y2=3.33
r72 26 28 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=1.2
+ $Y2=3.33
r73 23 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r74 23 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 21 35 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.78 $Y=3.33 $X2=3.6
+ $Y2=3.33
r76 21 22 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.78 $Y=3.33
+ $X2=3.932 $Y2=3.33
r77 20 38 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.085 $Y=3.33
+ $X2=4.56 $Y2=3.33
r78 20 22 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.085 $Y=3.33
+ $X2=3.932 $Y2=3.33
r79 16 22 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.932 $Y=3.245
+ $X2=3.932 $Y2=3.33
r80 16 18 24.3713 $w=3.03e-07 $l=6.45e-07 $layer=LI1_cond $X=3.932 $Y=3.245
+ $X2=3.932 $Y2=2.6
r81 12 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=3.245
+ $X2=0.835 $Y2=3.33
r82 12 14 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=0.835 $Y=3.245
+ $X2=0.835 $Y2=2.6
r83 3 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.735
+ $Y=2.455 $X2=3.875 $Y2=2.6
r84 2 49 300 $w=1.7e-07 $l=7.5776e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=2.455 $X2=3.015 $Y2=2.665
r85 1 14 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=0.645
+ $Y=2.455 $X2=0.88 $Y2=2.6
.ends

.subckt PM_SKY130_FD_SC_LP__HA_0%COUT 1 2 9 12 13 14 15 16 38
r21 23 38 1.60062 $w=3.58e-07 $l=5e-08 $layer=LI1_cond $X=4.535 $Y=1.245
+ $X2=4.535 $Y2=1.295
r22 15 16 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.575 $Y=1.665
+ $X2=4.575 $Y2=2.035
r23 15 40 9.87808 $w=2.78e-07 $l=2.4e-07 $layer=LI1_cond $X=4.575 $Y=1.665
+ $X2=4.575 $Y2=1.425
r24 14 40 4.21726 $w=3.58e-07 $l=1.13e-07 $layer=LI1_cond $X=4.535 $Y=1.312
+ $X2=4.535 $Y2=1.425
r25 14 38 0.544209 $w=3.58e-07 $l=1.7e-08 $layer=LI1_cond $X=4.535 $Y=1.312
+ $X2=4.535 $Y2=1.295
r26 14 23 0.576222 $w=3.58e-07 $l=1.8e-08 $layer=LI1_cond $X=4.535 $Y=1.227
+ $X2=4.535 $Y2=1.245
r27 13 14 9.66772 $w=3.58e-07 $l=3.02e-07 $layer=LI1_cond $X=4.535 $Y=0.925
+ $X2=4.535 $Y2=1.227
r28 13 28 3.36129 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=4.535 $Y=0.925
+ $X2=4.535 $Y2=0.82
r29 12 28 8.48326 $w=3.58e-07 $l=2.65e-07 $layer=LI1_cond $X=4.535 $Y=0.555
+ $X2=4.535 $Y2=0.82
r30 10 16 16.4635 $w=2.78e-07 $l=4e-07 $layer=LI1_cond $X=4.575 $Y=2.435
+ $X2=4.575 $Y2=2.035
r31 9 10 6.10861 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=2.6
+ $X2=4.485 $Y2=2.435
r32 2 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.28
+ $Y=2.455 $X2=4.42 $Y2=2.6
r33 1 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.4
+ $Y=0.675 $X2=4.54 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__HA_0%VGND 1 2 3 12 16 20 22 24 29 34 44 45 48 51 54
r58 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r59 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r60 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r62 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r63 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.02
+ $Y2=0
r64 42 44 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.56
+ $Y2=0
r65 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r66 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r67 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r68 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r69 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r70 35 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.105
+ $Y2=0
r71 35 37 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.64
+ $Y2=0
r72 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=4.02
+ $Y2=0
r73 34 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=3.6
+ $Y2=0
r74 33 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r75 33 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r76 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r77 30 48 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.7
+ $Y2=0
r78 30 32 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=0.805 $Y=0 $X2=1.68
+ $Y2=0
r79 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.105
+ $Y2=0
r80 29 32 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.68
+ $Y2=0
r81 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r82 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r83 24 48 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.7
+ $Y2=0
r84 24 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.24
+ $Y2=0
r85 22 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r86 22 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r87 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r88 18 20 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=4.02 $Y=0.085 $X2=4.02
+ $Y2=0.885
r89 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r90 14 16 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.445
r91 10 48 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r92 10 12 29.3117 $w=2.08e-07 $l=5.55e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.64
r93 3 20 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=3.795
+ $Y=0.675 $X2=4.02 $Y2=0.885
r94 2 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.235 $X2=2.105 $Y2=0.445
r95 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.43 $X2=0.69 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_LP__HA_0%A_307_47# 1 2 9 11 12 15
c29 12 0 1.08071e-19 $X=1.77 $Y=0.8
r30 13 15 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=2.57 $Y=0.715
+ $X2=2.57 $Y2=0.445
r31 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.44 $Y=0.8
+ $X2=2.57 $Y2=0.715
r32 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.44 $Y=0.8 $X2=1.77
+ $Y2=0.8
r33 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.665 $Y=0.715
+ $X2=1.77 $Y2=0.8
r34 7 9 14.2597 $w=2.08e-07 $l=2.7e-07 $layer=LI1_cond $X=1.665 $Y=0.715
+ $X2=1.665 $Y2=0.445
r35 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.235 $X2=2.535 $Y2=0.445
r36 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.675 $Y2=0.445
.ends

