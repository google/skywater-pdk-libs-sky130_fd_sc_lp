* File: sky130_fd_sc_lp__o31ai_2.pex.spice
* Created: Fri Aug 28 11:16:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31AI_2%A1 3 5 7 10 12 14 15 16 17 31
r50 30 31 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.99 $Y=1.44 $X2=1.06
+ $Y2=1.44
r51 28 30 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.97 $Y=1.44 $X2=0.99
+ $Y2=1.44
r52 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.44 $X2=0.97 $Y2=1.44
r53 26 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.63 $Y=1.44
+ $X2=0.97 $Y2=1.44
r54 25 26 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.56 $Y=1.44 $X2=0.63
+ $Y2=1.44
r55 22 25 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.54 $Y=1.44 $X2=0.56
+ $Y2=1.44
r56 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.44 $X2=0.54 $Y2=1.44
r57 17 29 8.41466 $w=3.13e-07 $l=2.3e-07 $layer=LI1_cond $X=1.2 $Y=1.367
+ $X2=0.97 $Y2=1.367
r58 16 29 9.14637 $w=3.13e-07 $l=2.5e-07 $layer=LI1_cond $X=0.72 $Y=1.367
+ $X2=0.97 $Y2=1.367
r59 16 23 6.58539 $w=3.13e-07 $l=1.8e-07 $layer=LI1_cond $X=0.72 $Y=1.367
+ $X2=0.54 $Y2=1.367
r60 15 23 10.9756 $w=3.13e-07 $l=3e-07 $layer=LI1_cond $X=0.24 $Y=1.367 $X2=0.54
+ $Y2=1.367
r61 12 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.275
+ $X2=1.06 $Y2=1.44
r62 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.06 $Y=1.275
+ $X2=1.06 $Y2=0.745
r63 8 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.605
+ $X2=0.99 $Y2=1.44
r64 8 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.99 $Y=1.605
+ $X2=0.99 $Y2=2.465
r65 5 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.275
+ $X2=0.63 $Y2=1.44
r66 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.63 $Y=1.275 $X2=0.63
+ $Y2=0.745
r67 1 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=1.605
+ $X2=0.56 $Y2=1.44
r68 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.56 $Y=1.605 $X2=0.56
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_2%A2 3 5 7 10 12 14 15 20 21 22
c56 22 0 2.83291e-20 $X=2.16 $Y=1.295
r57 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.11
+ $Y=1.44 $X2=2.11 $Y2=1.44
r58 22 27 1.82927 $w=3.13e-07 $l=5e-08 $layer=LI1_cond $X=2.16 $Y=1.367 $X2=2.11
+ $Y2=1.367
r59 21 27 15.7318 $w=3.13e-07 $l=4.3e-07 $layer=LI1_cond $X=1.68 $Y=1.367
+ $X2=2.11 $Y2=1.367
r60 20 26 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.265 $Y=1.44
+ $X2=2.11 $Y2=1.44
r61 18 19 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.49 $Y=1.44
+ $X2=1.85 $Y2=1.44
r62 16 18 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.42 $Y=1.44 $X2=1.49
+ $Y2=1.44
r63 15 26 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.925 $Y=1.44
+ $X2=2.11 $Y2=1.44
r64 15 19 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=1.44
+ $X2=1.85 $Y2=1.44
r65 12 20 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.34 $Y=1.275
+ $X2=2.265 $Y2=1.44
r66 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.34 $Y=1.275
+ $X2=2.34 $Y2=0.745
r67 8 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.605
+ $X2=1.85 $Y2=1.44
r68 8 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.85 $Y=1.605
+ $X2=1.85 $Y2=2.465
r69 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.275
+ $X2=1.49 $Y2=1.44
r70 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.49 $Y=1.275 $X2=1.49
+ $Y2=0.745
r71 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.605
+ $X2=1.42 $Y2=1.44
r72 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.42 $Y=1.605 $X2=1.42
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_2%A3 3 7 11 15 17 23 24
c56 23 0 2.83291e-20 $X=3.25 $Y=1.51
c57 15 0 1.17964e-19 $X=3.31 $Y=2.465
r58 23 25 8.98137 $w=3.22e-07 $l=6e-08 $layer=POLY_cond $X=3.25 $Y=1.51 $X2=3.31
+ $Y2=1.51
r59 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.51 $X2=3.25 $Y2=1.51
r60 21 23 7.48447 $w=3.22e-07 $l=5e-08 $layer=POLY_cond $X=3.2 $Y=1.51 $X2=3.25
+ $Y2=1.51
r61 20 21 59.8758 $w=3.22e-07 $l=4e-07 $layer=POLY_cond $X=2.8 $Y=1.51 $X2=3.2
+ $Y2=1.51
r62 19 20 4.49068 $w=3.22e-07 $l=3e-08 $layer=POLY_cond $X=2.77 $Y=1.51 $X2=2.8
+ $Y2=1.51
r63 17 24 4.70075 $w=3.78e-07 $l=1.55e-07 $layer=LI1_cond $X=3.225 $Y=1.665
+ $X2=3.225 $Y2=1.51
r64 13 25 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.675
+ $X2=3.31 $Y2=1.51
r65 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.31 $Y=1.675
+ $X2=3.31 $Y2=2.465
r66 9 21 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.2 $Y=1.345 $X2=3.2
+ $Y2=1.51
r67 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.2 $Y=1.345 $X2=3.2
+ $Y2=0.745
r68 5 20 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=1.675 $X2=2.8
+ $Y2=1.51
r69 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.8 $Y=1.675 $X2=2.8
+ $Y2=2.465
r70 1 19 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.345
+ $X2=2.77 $Y2=1.51
r71 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.77 $Y=1.345 $X2=2.77
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_2%B1 1 3 6 8 10 13 20 26 31
r44 29 31 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=1.397
+ $X2=4.26 $Y2=1.397
r45 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.425
+ $Y=1.44 $X2=4.425 $Y2=1.44
r46 26 28 12.7513 $w=3.78e-07 $l=1e-07 $layer=POLY_cond $X=4.325 $Y=1.47
+ $X2=4.425 $Y2=1.47
r47 25 26 24.8651 $w=3.78e-07 $l=1.95e-07 $layer=POLY_cond $X=4.13 $Y=1.47
+ $X2=4.325 $Y2=1.47
r48 24 25 29.9656 $w=3.78e-07 $l=2.35e-07 $layer=POLY_cond $X=3.895 $Y=1.47
+ $X2=4.13 $Y2=1.47
r49 20 29 4.14879 $w=3.73e-07 $l=1.35e-07 $layer=LI1_cond $X=4.56 $Y=1.397
+ $X2=4.425 $Y2=1.397
r50 18 24 10.8386 $w=3.78e-07 $l=8.5e-08 $layer=POLY_cond $X=3.81 $Y=1.47
+ $X2=3.895 $Y2=1.47
r51 18 22 14.0265 $w=3.78e-07 $l=1.1e-07 $layer=POLY_cond $X=3.81 $Y=1.47
+ $X2=3.7 $Y2=1.47
r52 17 31 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.81 $Y=1.5 $X2=4.26
+ $Y2=1.5
r53 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.81
+ $Y=1.5 $X2=3.81 $Y2=1.5
r54 11 26 24.4846 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.325 $Y=1.665
+ $X2=4.325 $Y2=1.47
r55 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.325 $Y=1.665
+ $X2=4.325 $Y2=2.465
r56 8 25 24.4846 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.13 $Y=1.275
+ $X2=4.13 $Y2=1.47
r57 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.13 $Y=1.275
+ $X2=4.13 $Y2=0.745
r58 4 24 24.4846 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.895 $Y=1.665
+ $X2=3.895 $Y2=1.47
r59 4 6 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.895 $Y=1.665 $X2=3.895
+ $Y2=2.465
r60 1 22 24.4846 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.7 $Y=1.275 $X2=3.7
+ $Y2=1.47
r61 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.7 $Y=1.275 $X2=3.7
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_2%A_44_367# 1 2 3 12 16 17 20 24 28 30
r51 26 28 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.065 $Y=1.865
+ $X2=2.065 $Y2=1.98
r52 25 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=1.78
+ $X2=1.205 $Y2=1.78
r53 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.9 $Y=1.78
+ $X2=2.065 $Y2=1.865
r54 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.9 $Y=1.78 $X2=1.37
+ $Y2=1.78
r55 20 22 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=1.205 $Y=1.98
+ $X2=1.205 $Y2=2.91
r56 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=1.865
+ $X2=1.205 $Y2=1.78
r57 18 20 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.205 $Y=1.865
+ $X2=1.205 $Y2=1.98
r58 16 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=1.78
+ $X2=1.205 $Y2=1.78
r59 16 17 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.04 $Y=1.78
+ $X2=0.51 $Y2=1.78
r60 12 14 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=0.345 $Y=1.98
+ $X2=0.345 $Y2=2.91
r61 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.345 $Y=1.865
+ $X2=0.51 $Y2=1.78
r62 10 12 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.345 $Y=1.865
+ $X2=0.345 $Y2=1.98
r63 3 28 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.925
+ $Y=1.835 $X2=2.065 $Y2=1.98
r64 2 22 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.835 $X2=1.205 $Y2=2.91
r65 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.835 $X2=1.205 $Y2=1.98
r66 1 14 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.835 $X2=0.345 $Y2=2.91
r67 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.835 $X2=0.345 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_2%VPWR 1 2 11 17 21 23 33 34 37 40
r53 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 34 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 31 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.11 $Y2=3.33
r58 31 33 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r61 27 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 26 29 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r63 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r64 24 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.87 $Y=3.33
+ $X2=0.775 $Y2=3.33
r65 24 26 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.87 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 23 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=4.11 $Y2=3.33
r67 23 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=3.6 $Y2=3.33
r68 21 30 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r69 21 27 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r70 17 20 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=4.11 $Y=2.18
+ $X2=4.11 $Y2=2.95
r71 15 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=3.33
r72 15 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=2.95
r73 11 14 43.7799 $w=1.88e-07 $l=7.5e-07 $layer=LI1_cond $X=0.775 $Y=2.2
+ $X2=0.775 $Y2=2.95
r74 9 37 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=3.245
+ $X2=0.775 $Y2=3.33
r75 9 14 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.775 $Y=3.245
+ $X2=0.775 $Y2=2.95
r76 2 20 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.97
+ $Y=1.835 $X2=4.11 $Y2=2.95
r77 2 17 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=3.97
+ $Y=1.835 $X2=4.11 $Y2=2.18
r78 1 14 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.835 $X2=0.775 $Y2=2.95
r79 1 11 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.835 $X2=0.775 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_2%A_299_367# 1 2 7 9 11 15
r17 13 15 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=3.05 $Y=2.905
+ $X2=3.05 $Y2=2.455
r18 12 18 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.73 $Y=2.99
+ $X2=1.635 $Y2=2.99
r19 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.92 $Y=2.99
+ $X2=3.05 $Y2=2.905
r20 11 12 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.92 $Y=2.99
+ $X2=1.73 $Y2=2.99
r21 7 18 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.635 $Y=2.905
+ $X2=1.635 $Y2=2.99
r22 7 9 41.1531 $w=1.88e-07 $l=7.05e-07 $layer=LI1_cond $X=1.635 $Y=2.905
+ $X2=1.635 $Y2=2.2
r23 2 15 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=2.875
+ $Y=1.835 $X2=3.015 $Y2=2.455
r24 1 18 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.835 $X2=1.635 $Y2=2.91
r25 1 9 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.835 $X2=1.635 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_2%Y 1 2 3 4 15 16 19 21 25 29 30 31 37 48 52
+ 53
c73 52 0 1.17964e-19 $X=2.585 $Y=1.98
r74 60 61 0.530435 $w=2.76e-07 $l=1.2e-08 $layer=LI1_cond $X=3.595 $Y=2.01
+ $X2=3.595 $Y2=2.022
r75 58 60 7.51449 $w=2.76e-07 $l=1.7e-07 $layer=LI1_cond $X=3.595 $Y=1.84
+ $X2=3.595 $Y2=2.01
r76 52 54 1.1127 $w=4.33e-07 $l=4.2e-08 $layer=LI1_cond $X=2.637 $Y=1.98
+ $X2=2.637 $Y2=2.022
r77 52 53 8.80985 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=2.637 $Y=1.98
+ $X2=2.637 $Y2=1.815
r78 38 54 5.46954 $w=1.95e-07 $l=2.18e-07 $layer=LI1_cond $X=2.855 $Y=2.022
+ $X2=2.637 $Y2=2.022
r79 37 61 2.79433 $w=1.95e-07 $l=1.8e-07 $layer=LI1_cond $X=3.415 $Y=2.022
+ $X2=3.595 $Y2=2.022
r80 31 61 0.574638 $w=2.76e-07 $l=1.3e-08 $layer=LI1_cond $X=3.595 $Y=2.035
+ $X2=3.595 $Y2=2.022
r81 31 48 8.9106 $w=5.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.595 $Y=2.12
+ $X2=3.595 $Y2=2.46
r82 30 37 16.7786 $w=1.93e-07 $l=2.95e-07 $layer=LI1_cond $X=3.12 $Y=2.022
+ $X2=3.415 $Y2=2.022
r83 30 38 15.0723 $w=1.93e-07 $l=2.65e-07 $layer=LI1_cond $X=3.12 $Y=2.022
+ $X2=2.855 $Y2=2.022
r84 29 42 2.95094 $w=4.33e-07 $l=8.5e-08 $layer=LI1_cond $X=2.637 $Y=2.035
+ $X2=2.637 $Y2=2.12
r85 29 54 0.344408 $w=4.33e-07 $l=1.3e-08 $layer=LI1_cond $X=2.637 $Y=2.035
+ $X2=2.637 $Y2=2.022
r86 29 42 1.06966 $w=6.13e-07 $l=5.5e-08 $layer=LI1_cond $X=2.64 $Y=2.427
+ $X2=2.585 $Y2=2.427
r87 25 27 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=4.575 $Y=1.98
+ $X2=4.575 $Y2=2.91
r88 23 25 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=4.575 $Y=1.925
+ $X2=4.575 $Y2=1.98
r89 22 58 3.57235 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.775 $Y=1.84
+ $X2=3.595 $Y2=1.84
r90 21 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.445 $Y=1.84
+ $X2=4.575 $Y2=1.925
r91 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.445 $Y=1.84
+ $X2=3.775 $Y2=1.84
r92 17 19 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.915 $Y=1.075
+ $X2=3.915 $Y2=0.68
r93 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.75 $Y=1.16
+ $X2=3.915 $Y2=1.075
r94 15 16 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.75 $Y=1.16
+ $X2=2.855 $Y2=1.16
r95 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=1.245
+ $X2=2.855 $Y2=1.16
r96 13 53 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.77 $Y=1.245
+ $X2=2.77 $Y2=1.815
r97 4 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.835 $X2=4.54 $Y2=2.91
r98 4 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.835 $X2=4.54 $Y2=1.98
r99 3 60 600 $w=1.7e-07 $l=2.68608e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.835 $X2=3.58 $Y2=2.01
r100 3 48 300 $w=1.7e-07 $l=7.15891e-07 $layer=licon1_PDIFF $count=2 $X=3.385
+ $Y=1.835 $X2=3.58 $Y2=2.46
r101 2 52 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.46
+ $Y=1.835 $X2=2.585 $Y2=1.98
r102 1 19 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=3.775
+ $Y=0.325 $X2=3.915 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_2%A_58_65# 1 2 3 4 5 16 18 20 24 26 30 32 35
+ 38 39 42 47 49
r67 49 50 6.72245 $w=2.45e-07 $l=1.35e-07 $layer=LI1_cond $X=2.497 $Y=0.82
+ $X2=2.497 $Y2=0.955
r68 40 42 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=4.38 $Y=0.425
+ $X2=4.38 $Y2=0.47
r69 38 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.25 $Y=0.34
+ $X2=4.38 $Y2=0.425
r70 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.25 $Y=0.34
+ $X2=3.58 $Y2=0.34
r71 35 52 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=0.735
+ $X2=3.45 $Y2=0.82
r72 35 37 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=3.45 $Y=0.735
+ $X2=3.45 $Y2=0.45
r73 34 39 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.45 $Y=0.425
+ $X2=3.58 $Y2=0.34
r74 34 37 1.10812 $w=2.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.45 $Y=0.425
+ $X2=3.45 $Y2=0.45
r75 33 49 2.87745 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=2.65 $Y=0.82
+ $X2=2.497 $Y2=0.82
r76 32 52 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.32 $Y=0.82 $X2=3.45
+ $Y2=0.82
r77 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.32 $Y=0.82
+ $X2=2.65 $Y2=0.82
r78 28 49 3.90749 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.497 $Y=0.735
+ $X2=2.497 $Y2=0.82
r79 28 30 10.7687 $w=3.03e-07 $l=2.85e-07 $layer=LI1_cond $X=2.497 $Y=0.735
+ $X2=2.497 $Y2=0.45
r80 27 47 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.41 $Y=0.955
+ $X2=1.295 $Y2=0.955
r81 26 50 2.87745 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=2.345 $Y=0.955
+ $X2=2.497 $Y2=0.955
r82 26 27 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.345 $Y=0.955 $X2=1.41
+ $Y2=0.955
r83 22 47 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.87
+ $X2=1.295 $Y2=0.955
r84 22 24 19.5414 $w=2.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.295 $Y=0.87
+ $X2=1.295 $Y2=0.48
r85 21 45 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.51 $Y=0.955
+ $X2=0.38 $Y2=0.955
r86 20 47 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.18 $Y=0.955
+ $X2=1.295 $Y2=0.955
r87 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.18 $Y=0.955
+ $X2=0.51 $Y2=0.955
r88 16 45 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.38 $Y=0.87 $X2=0.38
+ $Y2=0.955
r89 16 18 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=0.38 $Y=0.87
+ $X2=0.38 $Y2=0.48
r90 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.205
+ $Y=0.325 $X2=4.345 $Y2=0.47
r91 4 52 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=3.275
+ $Y=0.325 $X2=3.415 $Y2=0.82
r92 4 37 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.275
+ $Y=0.325 $X2=3.415 $Y2=0.45
r93 3 49 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.325 $X2=2.555 $Y2=0.82
r94 3 30 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.325 $X2=2.555 $Y2=0.45
r95 2 47 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=1.135
+ $Y=0.325 $X2=1.275 $Y2=0.955
r96 2 24 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.135
+ $Y=0.325 $X2=1.275 $Y2=0.48
r97 1 45 182 $w=1.7e-07 $l=6.89674e-07 $layer=licon1_NDIFF $count=1 $X=0.29
+ $Y=0.325 $X2=0.415 $Y2=0.955
r98 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.29
+ $Y=0.325 $X2=0.415 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_2%VGND 1 2 3 14 18 22 24 26 31 38 39 42 45 48
r61 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r62 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r63 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r64 39 49 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.12
+ $Y2=0
r65 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r66 36 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=0 $X2=2.985
+ $Y2=0
r67 36 38 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=3.15 $Y=0 $X2=4.56
+ $Y2=0
r68 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r69 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r70 32 45 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=1.877
+ $Y2=0
r71 32 34 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.64
+ $Y2=0
r72 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=2.985
+ $Y2=0
r73 31 34 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=2.64
+ $Y2=0
r74 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r75 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r76 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r77 27 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.845
+ $Y2=0
r78 27 29 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.2
+ $Y2=0
r79 26 45 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=1.877
+ $Y2=0
r80 26 29 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=1.2
+ $Y2=0
r81 24 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r82 24 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r83 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=0.085
+ $X2=2.985 $Y2=0
r84 20 22 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.985 $Y=0.085
+ $X2=2.985 $Y2=0.45
r85 16 45 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.877 $Y=0.085
+ $X2=1.877 $Y2=0
r86 16 18 9.04597 $w=5.93e-07 $l=4.5e-07 $layer=LI1_cond $X=1.877 $Y=0.085
+ $X2=1.877 $Y2=0.535
r87 12 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=0.085
+ $X2=0.845 $Y2=0
r88 12 14 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.845 $Y=0.085
+ $X2=0.845 $Y2=0.575
r89 3 22 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.845
+ $Y=0.325 $X2=2.985 $Y2=0.45
r90 2 18 91 $w=1.7e-07 $l=6.21188e-07 $layer=licon1_NDIFF $count=2 $X=1.565
+ $Y=0.325 $X2=2.09 $Y2=0.535
r91 1 14 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.705
+ $Y=0.325 $X2=0.845 $Y2=0.575
.ends

