* File: sky130_fd_sc_lp__a211oi_lp.spice
* Created: Wed Sep  2 09:18:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a211oi_lp.pex.spice"
.subckt sky130_fd_sc_lp__a211oi_lp  VNB VPB C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1008 A_137_57# N_C1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_C1_M1005_g A_137_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1000 A_295_57# N_B1_M1000_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75001.4 A=0.063
+ P=1.14 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g A_295_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1003 A_453_57# N_A1_M1003_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=24.276 NRS=0 M=1 R=2.8 SA=75001.8 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g A_453_57# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=24.276 M=1 R=2.8 SA=75002.2 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 A_181_409# N_C1_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.49 PD=1.24 PS=2.98 NRD=12.7853 NRS=40.3653 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1002 N_A_279_409#_M1002_d N_B1_M1002_g A_181_409# VPB PHIGHVT L=0.25 W=1
+ AD=0.16 AS=0.12 PD=1.32 PS=1.24 NRD=7.8603 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_279_409#_M1002_d VPB PHIGHVT L=0.25 W=1
+ AD=0.29 AS=0.16 PD=1.58 PS=1.32 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_A_279_409#_M1006_d N_A2_M1006_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.29 PD=2.57 PS=1.58 NRD=0 NRS=59.0803 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a211oi_lp.pxi.spice"
*
.ends
*
*
