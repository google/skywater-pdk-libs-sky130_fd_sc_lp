* File: sky130_fd_sc_lp__bufkapwr_2.pex.spice
* Created: Fri Aug 28 10:11:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_2%A 3 6 8 11 13
r32 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.94
+ $X2=0.51 $Y2=1.105
r33 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.94
+ $X2=0.51 $Y2=0.775
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=0.94 $X2=0.51 $Y2=0.94
r35 8 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=0.94 $X2=0.51
+ $Y2=0.94
r36 6 14 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.105
r37 3 13 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_2%A_27_47# 1 2 9 13 17 21 24 27 33 39 41 45
r68 45 46 0.710914 $w=3.39e-07 $l=5e-09 $layer=POLY_cond $X=1.385 $Y=1.375
+ $X2=1.39 $Y2=1.375
r69 42 43 0.710914 $w=3.39e-07 $l=5e-09 $layer=POLY_cond $X=0.955 $Y=1.375
+ $X2=0.96 $Y2=1.375
r70 36 39 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.435 $X2=0.26
+ $Y2=0.435
r71 34 45 47.6313 $w=3.39e-07 $l=3.35e-07 $layer=POLY_cond $X=1.05 $Y=1.375
+ $X2=1.385 $Y2=1.375
r72 34 43 12.7965 $w=3.39e-07 $l=9e-08 $layer=POLY_cond $X=1.05 $Y=1.375
+ $X2=0.96 $Y2=1.375
r73 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.38 $X2=1.05 $Y2=1.38
r74 31 41 1.05597 $w=2.6e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=1.405
+ $X2=0.24 $Y2=1.405
r75 31 33 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=0.395 $Y=1.405
+ $X2=1.05 $Y2=1.405
r76 27 29 31.2275 $w=3.08e-07 $l=8.4e-07 $layer=LI1_cond $X=0.24 $Y=2.04
+ $X2=0.24 $Y2=2.88
r77 25 41 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=0.24 $Y=1.535
+ $X2=0.24 $Y2=1.405
r78 25 27 18.7737 $w=3.08e-07 $l=5.05e-07 $layer=LI1_cond $X=0.24 $Y=1.535
+ $X2=0.24 $Y2=2.04
r79 24 41 5.51899 $w=2.4e-07 $l=1.61245e-07 $layer=LI1_cond $X=0.17 $Y=1.275
+ $X2=0.24 $Y2=1.405
r80 23 36 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.17 $Y=0.605
+ $X2=0.17 $Y2=0.435
r81 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=0.605
+ $X2=0.17 $Y2=1.275
r82 19 46 21.8644 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.39 $Y=1.205
+ $X2=1.39 $Y2=1.375
r83 19 21 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.39 $Y=1.205
+ $X2=1.39 $Y2=0.445
r84 15 45 21.8644 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.385 $Y=1.545
+ $X2=1.385 $Y2=1.375
r85 15 17 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=1.385 $Y=1.545
+ $X2=1.385 $Y2=2.465
r86 11 43 21.8644 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.96 $Y=1.205
+ $X2=0.96 $Y2=1.375
r87 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.96 $Y=1.205
+ $X2=0.96 $Y2=0.445
r88 7 42 21.8644 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.955 $Y=1.545
+ $X2=0.955 $Y2=1.375
r89 7 9 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=0.955 $Y=1.545
+ $X2=0.955 $Y2=2.465
r90 2 29 400 $w=1.7e-07 $l=1.10574e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.88
r91 2 27 400 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.04
r92 1 39 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_2%KAPWR 1 2 7 10 18 22
r24 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.595 $Y=2.81
+ $X2=1.595 $Y2=2.81
r25 18 21 26.2124 $w=2.53e-07 $l=5.8e-07 $layer=LI1_cond $X=1.602 $Y=2.23
+ $X2=1.602 $Y2=2.81
r26 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.71 $Y=2.81
+ $X2=0.71 $Y2=2.81
r27 10 13 28.6252 $w=3.08e-07 $l=7.7e-07 $layer=LI1_cond $X=0.72 $Y=2.04
+ $X2=0.72 $Y2=2.81
r28 7 22 0.367476 $w=2.55e-07 $l=6.35e-07 $layer=MET1_cond $X=0.96 $Y=2.817
+ $X2=1.595 $Y2=2.817
r29 7 14 0.144675 $w=2.55e-07 $l=2.5e-07 $layer=MET1_cond $X=0.96 $Y=2.817
+ $X2=0.71 $Y2=2.817
r30 2 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.91
r31 2 18 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.23
r32 1 13 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.88
r33 1 10 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_2%X 1 2 9 13 14 15 16 17 26 36
r39 31 36 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=1.6 $Y=1.725 $X2=1.6
+ $Y2=1.665
r40 17 31 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=1.81 $X2=1.6
+ $Y2=1.81
r41 17 36 0.348413 $w=4.28e-07 $l=1.3e-08 $layer=LI1_cond $X=1.6 $Y=1.652
+ $X2=1.6 $Y2=1.665
r42 16 17 9.56796 $w=4.28e-07 $l=3.57e-07 $layer=LI1_cond $X=1.6 $Y=1.295
+ $X2=1.6 $Y2=1.652
r43 16 30 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.6 $Y=1.295 $X2=1.6
+ $Y2=1.105
r44 15 30 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=0.942 $X2=1.6
+ $Y2=0.942
r45 14 30 14.1839 $w=3.23e-07 $l=4e-07 $layer=LI1_cond $X=1.2 $Y=0.942 $X2=1.6
+ $Y2=0.942
r46 14 24 0.886495 $w=3.23e-07 $l=2.5e-08 $layer=LI1_cond $X=1.2 $Y=0.942
+ $X2=1.175 $Y2=0.942
r47 13 24 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=1.175 $Y=0.555
+ $X2=1.175 $Y2=0.78
r48 13 26 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=1.175 $Y=0.555
+ $X2=1.175 $Y2=0.44
r49 9 11 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=1.175 $Y=2.04
+ $X2=1.175 $Y2=2.88
r50 7 31 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.175 $Y=1.81
+ $X2=1.6 $Y2=1.81
r51 7 9 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.175 $Y=1.895
+ $X2=1.175 $Y2=2.04
r52 2 11 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.88
r53 2 9 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.04
r54 1 26 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.175 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_2%VGND 1 2 9 11 13 15 17 22 28 32
r29 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r30 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r31 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r32 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 23 28 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.692
+ $Y2=0
r34 23 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.2
+ $Y2=0
r35 22 31 3.96354 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.697
+ $Y2=0
r36 22 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.2
+ $Y2=0
r37 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r38 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 17 28 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.692
+ $Y2=0
r40 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.24
+ $Y2=0
r41 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r42 15 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r43 11 31 3.21368 $w=2.55e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.697 $Y2=0
r44 11 13 16.2698 $w=2.53e-07 $l=3.6e-07 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.602 $Y2=0.445
r45 7 28 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0
r46 7 9 14.877 $w=2.73e-07 $l=3.55e-07 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0.44
r47 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.235 $X2=1.605 $Y2=0.445
r48 1 9 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__BUFKAPWR_2%VPWR 1 8 14
r23 5 14 0.0081048 $w=1.92e-06 $l=1.22e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.96 $Y2=3.208
r24 5 8 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33 $X2=1.68
+ $Y2=3.33
r25 4 8 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.68
+ $Y2=3.33
r26 4 5 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33 $X2=0.24
+ $Y2=3.33
r27 1 14 6.64328e-05 $w=1.92e-06 $l=1e-09 $layer=MET1_cond $X=0.96 $Y=3.207
+ $X2=0.96 $Y2=3.208
.ends

