* File: sky130_fd_sc_lp__and4_lp2.pxi.spice
* Created: Wed Sep  2 09:33:05 2020
* 
x_PM_SKY130_FD_SC_LP__AND4_LP2%A_84_21# N_A_84_21#_M1000_d N_A_84_21#_M1009_d
+ N_A_84_21#_M1007_d N_A_84_21#_c_74_n N_A_84_21#_M1005_g N_A_84_21#_M1010_g
+ N_A_84_21#_M1008_g N_A_84_21#_c_76_n N_A_84_21#_c_77_n N_A_84_21#_c_78_n
+ N_A_84_21#_c_79_n N_A_84_21#_c_80_n N_A_84_21#_c_81_n N_A_84_21#_c_87_n
+ N_A_84_21#_c_147_p N_A_84_21#_c_88_n N_A_84_21#_c_89_n N_A_84_21#_c_90_n
+ N_A_84_21#_c_82_n N_A_84_21#_c_83_n N_A_84_21#_c_84_n N_A_84_21#_c_91_n
+ PM_SKY130_FD_SC_LP__AND4_LP2%A_84_21#
x_PM_SKY130_FD_SC_LP__AND4_LP2%D N_D_M1009_g N_D_c_183_n N_D_M1004_g N_D_c_184_n
+ N_D_c_185_n N_D_c_186_n N_D_c_187_n D D N_D_c_189_n
+ PM_SKY130_FD_SC_LP__AND4_LP2%D
x_PM_SKY130_FD_SC_LP__AND4_LP2%C N_C_M1006_g N_C_M1002_g N_C_c_238_n N_C_c_239_n
+ C C N_C_c_241_n PM_SKY130_FD_SC_LP__AND4_LP2%C
x_PM_SKY130_FD_SC_LP__AND4_LP2%B N_B_M1003_g N_B_c_278_n N_B_M1007_g N_B_c_279_n
+ B B N_B_c_280_n N_B_c_281_n PM_SKY130_FD_SC_LP__AND4_LP2%B
x_PM_SKY130_FD_SC_LP__AND4_LP2%A N_A_c_317_n N_A_M1000_g N_A_M1001_g N_A_c_318_n
+ N_A_c_319_n N_A_c_320_n N_A_c_321_n A A N_A_c_322_n N_A_c_323_n
+ PM_SKY130_FD_SC_LP__AND4_LP2%A
x_PM_SKY130_FD_SC_LP__AND4_LP2%X N_X_M1005_s N_X_M1010_s N_X_c_353_n X X X
+ N_X_c_354_n X PM_SKY130_FD_SC_LP__AND4_LP2%X
x_PM_SKY130_FD_SC_LP__AND4_LP2%VPWR N_VPWR_M1010_d N_VPWR_M1006_d N_VPWR_M1001_d
+ N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n
+ N_VPWR_c_381_n VPWR N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_375_n
+ PM_SKY130_FD_SC_LP__AND4_LP2%VPWR
x_PM_SKY130_FD_SC_LP__AND4_LP2%VGND N_VGND_M1008_d N_VGND_c_423_n VGND
+ N_VGND_c_424_n N_VGND_c_425_n N_VGND_c_426_n N_VGND_c_427_n
+ PM_SKY130_FD_SC_LP__AND4_LP2%VGND
cc_1 VNB N_A_84_21#_c_74_n 0.0325119f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_2 VNB N_A_84_21#_M1010_g 0.00282885f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.545
cc_3 VNB N_A_84_21#_c_76_n 0.0200515f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.88
cc_4 VNB N_A_84_21#_c_77_n 0.0149226f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.61
cc_5 VNB N_A_84_21#_c_78_n 0.00222358f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.12
cc_6 VNB N_A_84_21#_c_79_n 0.00191586f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.43
cc_7 VNB N_A_84_21#_c_80_n 2.70146e-19 $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.97
cc_8 VNB N_A_84_21#_c_81_n 0.0536063f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.855
cc_9 VNB N_A_84_21#_c_82_n 0.0191244f $X=-0.19 $Y=-0.245 $X2=2.78 $Y2=0.47
cc_10 VNB N_A_84_21#_c_83_n 0.0411451f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.105
cc_11 VNB N_A_84_21#_c_84_n 0.00111966f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.61
cc_12 VNB N_D_c_183_n 0.0152548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D_c_184_n 0.0140408f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_14 VNB N_D_c_185_n 0.0231052f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_15 VNB N_D_c_186_n 0.00215656f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.61
cc_16 VNB N_D_c_187_n 0.0178014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB D 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_18 VNB N_D_c_189_n 0.0163625f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.438
cc_19 VNB N_C_M1002_g 0.0333697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_c_238_n 0.0234675f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_21 VNB N_C_c_239_n 0.00208291f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_22 VNB C 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.61
cc_23 VNB N_C_c_241_n 0.0165645f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_24 VNB N_B_M1003_g 0.0335716f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=2.045
cc_25 VNB N_B_c_278_n 0.00193406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_c_279_n 0.0217904f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_27 VNB N_B_c_280_n 0.015746f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_28 VNB N_B_c_281_n 0.00559843f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_29 VNB N_A_c_317_n 0.0177151f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.235
cc_30 VNB N_A_c_318_n 0.0217667f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_31 VNB N_A_c_319_n 0.0192868f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.545
cc_32 VNB N_A_c_320_n 0.027533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_c_321_n 0.00244376f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_34 VNB N_A_c_322_n 0.0185781f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.438
cc_35 VNB N_A_c_323_n 0.035306f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.61
cc_36 VNB N_X_c_353_n 0.0219529f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_37 VNB N_X_c_354_n 0.0460252f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.055
cc_38 VNB N_VPWR_c_375_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.9
cc_39 VNB N_VGND_c_423_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_424_n 0.026731f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_41 VNB N_VGND_c_425_n 0.066739f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_42 VNB N_VGND_c_426_n 0.201826f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_43 VNB N_VGND_c_427_n 0.00510817f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.73
cc_44 VPB N_A_84_21#_M1010_g 0.0453264f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_45 VPB N_A_84_21#_c_80_n 0.00257114f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.97
cc_46 VPB N_A_84_21#_c_87_n 0.00623881f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=2.055
cc_47 VPB N_A_84_21#_c_88_n 0.00207453f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=2.19
cc_48 VPB N_A_84_21#_c_89_n 0.0177179f $X=-0.19 $Y=1.655 $X2=2.365 $Y2=2.055
cc_49 VPB N_A_84_21#_c_90_n 0.00207453f $X=-0.19 $Y=1.655 $X2=2.53 $Y2=2.19
cc_50 VPB N_A_84_21#_c_91_n 0.00902579f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=2.055
cc_51 VPB N_D_M1009_g 0.0319341f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.045
cc_52 VPB N_D_c_186_n 0.0119306f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.61
cc_53 VPB D 7.4543e-19 $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_54 VPB N_C_M1006_g 0.0321773f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.045
cc_55 VPB N_C_c_239_n 0.0116277f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_56 VPB C 7.56276e-19 $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.61
cc_57 VPB N_B_c_278_n 0.010958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_B_M1007_g 0.0326253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_B_c_281_n 0.00212235f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_60 VPB N_A_M1001_g 0.0407138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_c_321_n 0.0132804f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.73
cc_62 VPB N_A_c_323_n 0.00925731f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.61
cc_63 VPB X 0.054923f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.61
cc_64 VPB N_X_c_354_n 0.0126158f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=2.055
cc_65 VPB N_VPWR_c_376_n 0.0041643f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_66 VPB N_VPWR_c_377_n 0.00417575f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_67 VPB N_VPWR_c_378_n 0.0119948f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=0.88
cc_68 VPB N_VPWR_c_379_n 0.0470736f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.88
cc_69 VPB N_VPWR_c_380_n 0.0205366f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.61
cc_70 VPB N_VPWR_c_381_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.97
cc_71 VPB N_VPWR_c_382_n 0.0219685f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=2.19
cc_72 VPB N_VPWR_c_383_n 0.0246129f $X=-0.19 $Y=1.655 $X2=1.555 $Y2=2.055
cc_73 VPB N_VPWR_c_375_n 0.0546651f $X=-0.19 $Y=1.655 $X2=2.53 $Y2=2.9
cc_74 N_A_84_21#_M1010_g N_D_M1009_g 0.0251349f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_75 N_A_84_21#_c_80_n N_D_M1009_g 0.003755f $X=0.725 $Y=1.97 $X2=0 $Y2=0
cc_76 N_A_84_21#_c_87_n N_D_M1009_g 0.0187754f $X=1.225 $Y=2.055 $X2=0 $Y2=0
cc_77 N_A_84_21#_c_88_n N_D_M1009_g 0.0145863f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_78 N_A_84_21#_c_91_n N_D_M1009_g 0.00163378f $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_79 N_A_84_21#_c_74_n N_D_c_183_n 0.0131268f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_80 N_A_84_21#_c_78_n N_D_c_184_n 0.00360238f $X=0.63 $Y=1.12 $X2=0 $Y2=0
cc_81 N_A_84_21#_c_81_n N_D_c_184_n 0.00465822f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_82 N_A_84_21#_c_83_n N_D_c_184_n 0.0065402f $X=0.615 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A_84_21#_M1010_g N_D_c_185_n 0.00687047f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_84 N_A_84_21#_c_77_n N_D_c_185_n 0.0153097f $X=0.607 $Y=1.61 $X2=0 $Y2=0
cc_85 N_A_84_21#_c_84_n N_D_c_185_n 0.00131808f $X=0.63 $Y=1.61 $X2=0 $Y2=0
cc_86 N_A_84_21#_c_80_n N_D_c_186_n 0.00131808f $X=0.725 $Y=1.97 $X2=0 $Y2=0
cc_87 N_A_84_21#_c_91_n N_D_c_186_n 5.35752e-19 $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_88 N_A_84_21#_c_76_n N_D_c_187_n 0.00877648f $X=0.675 $Y=0.88 $X2=0 $Y2=0
cc_89 N_A_84_21#_c_81_n N_D_c_187_n 0.0129296f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_90 N_A_84_21#_c_79_n D 0.0501772f $X=0.63 $Y=1.43 $X2=0 $Y2=0
cc_91 N_A_84_21#_c_81_n D 0.0245051f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_92 N_A_84_21#_c_87_n D 0.017002f $X=1.225 $Y=2.055 $X2=0 $Y2=0
cc_93 N_A_84_21#_c_83_n D 5.82133e-19 $X=0.615 $Y=1.105 $X2=0 $Y2=0
cc_94 N_A_84_21#_c_91_n D 0.00790183f $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_95 N_A_84_21#_c_79_n N_D_c_189_n 0.00131808f $X=0.63 $Y=1.43 $X2=0 $Y2=0
cc_96 N_A_84_21#_c_81_n N_D_c_189_n 0.00123003f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_97 N_A_84_21#_c_83_n N_D_c_189_n 0.0153097f $X=0.615 $Y=1.105 $X2=0 $Y2=0
cc_98 N_A_84_21#_c_88_n N_C_M1006_g 0.0168806f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_99 N_A_84_21#_c_89_n N_C_M1006_g 0.0182829f $X=2.365 $Y=2.055 $X2=0 $Y2=0
cc_100 N_A_84_21#_c_90_n N_C_M1006_g 9.22258e-19 $X=2.53 $Y=2.19 $X2=0 $Y2=0
cc_101 N_A_84_21#_c_91_n N_C_M1006_g 0.00161889f $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_102 N_A_84_21#_c_81_n N_C_M1002_g 0.0114638f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_103 N_A_84_21#_c_89_n N_C_c_239_n 5.42828e-19 $X=2.365 $Y=2.055 $X2=0 $Y2=0
cc_104 N_A_84_21#_c_81_n C 0.0245051f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_105 N_A_84_21#_c_89_n C 0.0223517f $X=2.365 $Y=2.055 $X2=0 $Y2=0
cc_106 N_A_84_21#_c_91_n C 0.00193735f $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_107 N_A_84_21#_c_81_n N_C_c_241_n 0.00122995f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_108 N_A_84_21#_c_81_n N_B_M1003_g 0.0115229f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_109 N_A_84_21#_c_82_n N_B_M1003_g 0.00249736f $X=2.78 $Y=0.47 $X2=0 $Y2=0
cc_110 N_A_84_21#_c_89_n N_B_c_278_n 5.77992e-19 $X=2.365 $Y=2.055 $X2=0 $Y2=0
cc_111 N_A_84_21#_c_88_n N_B_M1007_g 9.15887e-19 $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_112 N_A_84_21#_c_89_n N_B_M1007_g 0.0206408f $X=2.365 $Y=2.055 $X2=0 $Y2=0
cc_113 N_A_84_21#_c_90_n N_B_M1007_g 0.0155619f $X=2.53 $Y=2.19 $X2=0 $Y2=0
cc_114 N_A_84_21#_c_81_n N_B_c_280_n 0.00123028f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_115 N_A_84_21#_c_81_n N_B_c_281_n 0.0289521f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_116 N_A_84_21#_c_89_n N_B_c_281_n 0.0290891f $X=2.365 $Y=2.055 $X2=0 $Y2=0
cc_117 N_A_84_21#_c_82_n N_A_c_317_n 0.0101133f $X=2.78 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_84_21#_c_89_n N_A_M1001_g 0.00597021f $X=2.365 $Y=2.055 $X2=0 $Y2=0
cc_119 N_A_84_21#_c_90_n N_A_M1001_g 0.016587f $X=2.53 $Y=2.19 $X2=0 $Y2=0
cc_120 N_A_84_21#_c_81_n N_A_c_318_n 0.0118201f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_121 N_A_84_21#_c_82_n N_A_c_318_n 0.00600519f $X=2.78 $Y=0.47 $X2=0 $Y2=0
cc_122 N_A_84_21#_c_81_n N_A_c_319_n 0.00497558f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_123 N_A_84_21#_c_81_n N_A_c_322_n 9.65096e-19 $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_124 N_A_84_21#_c_81_n N_A_c_323_n 0.0226737f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_125 N_A_84_21#_c_89_n N_A_c_323_n 0.00193735f $X=2.365 $Y=2.055 $X2=0 $Y2=0
cc_126 N_A_84_21#_c_74_n N_X_c_353_n 0.00986136f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_127 N_A_84_21#_M1010_g X 0.0240034f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_128 N_A_84_21#_c_80_n X 0.00340231f $X=0.725 $Y=1.97 $X2=0 $Y2=0
cc_129 N_A_84_21#_c_147_p X 0.0130043f $X=0.81 $Y=2.055 $X2=0 $Y2=0
cc_130 N_A_84_21#_c_84_n X 4.16515e-19 $X=0.63 $Y=1.61 $X2=0 $Y2=0
cc_131 N_A_84_21#_c_74_n N_X_c_354_n 0.0047922f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_132 N_A_84_21#_c_78_n N_X_c_354_n 0.0206395f $X=0.63 $Y=1.12 $X2=0 $Y2=0
cc_133 N_A_84_21#_c_79_n N_X_c_354_n 0.0354f $X=0.63 $Y=1.43 $X2=0 $Y2=0
cc_134 N_A_84_21#_c_80_n N_X_c_354_n 0.010399f $X=0.725 $Y=1.97 $X2=0 $Y2=0
cc_135 N_A_84_21#_c_83_n N_X_c_354_n 0.0228828f $X=0.615 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A_84_21#_c_87_n N_VPWR_M1010_d 0.00143726f $X=1.225 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_84_21#_c_147_p N_VPWR_M1010_d 7.70949e-19 $X=0.81 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_84_21#_c_89_n N_VPWR_M1006_d 0.00267852f $X=2.365 $Y=2.055 $X2=0
+ $Y2=0
cc_139 N_A_84_21#_M1010_g N_VPWR_c_376_n 0.0185453f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_140 N_A_84_21#_c_87_n N_VPWR_c_376_n 0.0103329f $X=1.225 $Y=2.055 $X2=0 $Y2=0
cc_141 N_A_84_21#_c_147_p N_VPWR_c_376_n 0.00777198f $X=0.81 $Y=2.055 $X2=0
+ $Y2=0
cc_142 N_A_84_21#_c_88_n N_VPWR_c_376_n 0.0222114f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_143 N_A_84_21#_c_88_n N_VPWR_c_377_n 0.0490886f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_144 N_A_84_21#_c_89_n N_VPWR_c_377_n 0.0208822f $X=2.365 $Y=2.055 $X2=0 $Y2=0
cc_145 N_A_84_21#_c_90_n N_VPWR_c_377_n 0.0193194f $X=2.53 $Y=2.19 $X2=0 $Y2=0
cc_146 N_A_84_21#_c_89_n N_VPWR_c_379_n 0.00805415f $X=2.365 $Y=2.055 $X2=0
+ $Y2=0
cc_147 N_A_84_21#_c_90_n N_VPWR_c_379_n 0.0609159f $X=2.53 $Y=2.19 $X2=0 $Y2=0
cc_148 N_A_84_21#_c_88_n N_VPWR_c_380_n 0.021949f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_149 N_A_84_21#_c_90_n N_VPWR_c_382_n 0.021949f $X=2.53 $Y=2.19 $X2=0 $Y2=0
cc_150 N_A_84_21#_M1010_g N_VPWR_c_383_n 0.00769046f $X=0.56 $Y=2.545 $X2=0
+ $Y2=0
cc_151 N_A_84_21#_M1010_g N_VPWR_c_375_n 0.0140941f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_152 N_A_84_21#_c_88_n N_VPWR_c_375_n 0.0124703f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_153 N_A_84_21#_c_90_n N_VPWR_c_375_n 0.0124703f $X=2.53 $Y=2.19 $X2=0 $Y2=0
cc_154 N_A_84_21#_c_74_n N_VGND_c_423_n 0.0131302f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_155 N_A_84_21#_c_81_n N_VGND_c_423_n 0.0222521f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_156 N_A_84_21#_c_74_n N_VGND_c_424_n 0.0103533f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_157 N_A_84_21#_c_76_n N_VGND_c_424_n 6.21075e-19 $X=0.675 $Y=0.88 $X2=0 $Y2=0
cc_158 N_A_84_21#_c_82_n N_VGND_c_425_n 0.0197788f $X=2.78 $Y=0.47 $X2=0 $Y2=0
cc_159 N_A_84_21#_M1000_d N_VGND_c_426_n 0.00232985f $X=2.64 $Y=0.235 $X2=0
+ $Y2=0
cc_160 N_A_84_21#_c_74_n N_VGND_c_426_n 0.015166f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_161 N_A_84_21#_c_76_n N_VGND_c_426_n 8.18184e-19 $X=0.675 $Y=0.88 $X2=0 $Y2=0
cc_162 N_A_84_21#_c_78_n N_VGND_c_426_n 0.00634285f $X=0.63 $Y=1.12 $X2=0 $Y2=0
cc_163 N_A_84_21#_c_81_n N_VGND_c_426_n 0.0502596f $X=2.615 $Y=0.855 $X2=0 $Y2=0
cc_164 N_A_84_21#_c_82_n N_VGND_c_426_n 0.0125782f $X=2.78 $Y=0.47 $X2=0 $Y2=0
cc_165 N_D_M1009_g N_C_M1006_g 0.0196434f $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_166 N_D_c_183_n N_C_M1002_g 0.0437936f $X=1.395 $Y=0.73 $X2=0 $Y2=0
cc_167 N_D_c_184_n N_C_M1002_g 0.00845519f $X=1.155 $Y=1.12 $X2=0 $Y2=0
cc_168 N_D_c_185_n N_C_c_238_n 0.0135694f $X=1.155 $Y=1.625 $X2=0 $Y2=0
cc_169 N_D_c_186_n N_C_c_239_n 0.0135694f $X=1.155 $Y=1.79 $X2=0 $Y2=0
cc_170 D C 0.0423335f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_171 N_D_c_189_n C 0.00232658f $X=1.155 $Y=1.285 $X2=0 $Y2=0
cc_172 D N_C_c_241_n 0.00232658f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_173 N_D_c_189_n N_C_c_241_n 0.0135694f $X=1.155 $Y=1.285 $X2=0 $Y2=0
cc_174 N_D_M1009_g X 8.80684e-19 $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_175 N_D_M1009_g N_VPWR_c_376_n 0.00314852f $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_176 N_D_M1009_g N_VPWR_c_377_n 8.63241e-19 $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_177 N_D_M1009_g N_VPWR_c_380_n 0.0086001f $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_178 N_D_M1009_g N_VPWR_c_375_n 0.0156118f $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_179 N_D_c_183_n N_VGND_c_423_n 0.0124929f $X=1.395 $Y=0.73 $X2=0 $Y2=0
cc_180 N_D_c_187_n N_VGND_c_423_n 0.00181468f $X=1.395 $Y=0.805 $X2=0 $Y2=0
cc_181 N_D_c_183_n N_VGND_c_425_n 0.00585385f $X=1.395 $Y=0.73 $X2=0 $Y2=0
cc_182 N_D_c_187_n N_VGND_c_425_n 0.0017538f $X=1.395 $Y=0.805 $X2=0 $Y2=0
cc_183 N_D_c_183_n N_VGND_c_426_n 0.00652711f $X=1.395 $Y=0.73 $X2=0 $Y2=0
cc_184 N_D_c_187_n N_VGND_c_426_n 0.00234546f $X=1.395 $Y=0.805 $X2=0 $Y2=0
cc_185 N_C_M1002_g N_B_M1003_g 0.0235099f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_186 N_C_c_239_n N_B_c_278_n 0.0235099f $X=1.695 $Y=1.79 $X2=0 $Y2=0
cc_187 N_C_M1006_g N_B_M1007_g 0.0332064f $X=1.655 $Y=2.545 $X2=0 $Y2=0
cc_188 N_C_c_238_n N_B_c_279_n 0.0235099f $X=1.695 $Y=1.625 $X2=0 $Y2=0
cc_189 C N_B_c_280_n 7.64905e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_190 N_C_c_241_n N_B_c_280_n 0.0235099f $X=1.695 $Y=1.285 $X2=0 $Y2=0
cc_191 C N_B_c_281_n 0.0503126f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_192 N_C_c_241_n N_B_c_281_n 0.00411812f $X=1.695 $Y=1.285 $X2=0 $Y2=0
cc_193 N_C_M1006_g N_VPWR_c_377_n 0.0176406f $X=1.655 $Y=2.545 $X2=0 $Y2=0
cc_194 N_C_M1006_g N_VPWR_c_380_n 0.00769046f $X=1.655 $Y=2.545 $X2=0 $Y2=0
cc_195 N_C_M1006_g N_VPWR_c_375_n 0.0134474f $X=1.655 $Y=2.545 $X2=0 $Y2=0
cc_196 N_C_M1002_g N_VGND_c_425_n 0.00585385f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_197 N_C_M1002_g N_VGND_c_426_n 0.00619611f $X=1.785 $Y=0.445 $X2=0 $Y2=0
cc_198 N_B_M1003_g N_A_c_317_n 0.0426524f $X=2.175 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_199 N_B_M1007_g N_A_M1001_g 0.0196512f $X=2.265 $Y=2.545 $X2=0 $Y2=0
cc_200 N_B_M1003_g N_A_c_319_n 0.00782887f $X=2.175 $Y=0.445 $X2=0 $Y2=0
cc_201 N_B_c_279_n N_A_c_320_n 0.0115267f $X=2.265 $Y=1.625 $X2=0 $Y2=0
cc_202 N_B_c_278_n N_A_c_321_n 0.0115267f $X=2.265 $Y=1.79 $X2=0 $Y2=0
cc_203 N_B_c_280_n N_A_c_322_n 0.0115267f $X=2.265 $Y=1.285 $X2=0 $Y2=0
cc_204 N_B_c_281_n N_A_c_322_n 0.00245756f $X=2.265 $Y=1.285 $X2=0 $Y2=0
cc_205 N_B_c_280_n N_A_c_323_n 0.00245345f $X=2.265 $Y=1.285 $X2=0 $Y2=0
cc_206 N_B_c_281_n N_A_c_323_n 0.0401411f $X=2.265 $Y=1.285 $X2=0 $Y2=0
cc_207 N_B_M1007_g N_VPWR_c_377_n 0.00711482f $X=2.265 $Y=2.545 $X2=0 $Y2=0
cc_208 N_B_M1007_g N_VPWR_c_379_n 9.45246e-19 $X=2.265 $Y=2.545 $X2=0 $Y2=0
cc_209 N_B_M1007_g N_VPWR_c_382_n 0.0086001f $X=2.265 $Y=2.545 $X2=0 $Y2=0
cc_210 N_B_M1007_g N_VPWR_c_375_n 0.0158034f $X=2.265 $Y=2.545 $X2=0 $Y2=0
cc_211 N_B_M1003_g N_VGND_c_425_n 0.00585385f $X=2.175 $Y=0.445 $X2=0 $Y2=0
cc_212 N_B_M1003_g N_VGND_c_426_n 0.00619611f $X=2.175 $Y=0.445 $X2=0 $Y2=0
cc_213 N_A_M1001_g N_VPWR_c_379_n 0.0237533f $X=2.795 $Y=2.545 $X2=0 $Y2=0
cc_214 N_A_c_321_n N_VPWR_c_379_n 6.02959e-19 $X=2.835 $Y=1.79 $X2=0 $Y2=0
cc_215 N_A_c_323_n N_VPWR_c_379_n 0.0238273f $X=2.835 $Y=1.285 $X2=0 $Y2=0
cc_216 N_A_M1001_g N_VPWR_c_382_n 0.00769046f $X=2.795 $Y=2.545 $X2=0 $Y2=0
cc_217 N_A_M1001_g N_VPWR_c_375_n 0.0134474f $X=2.795 $Y=2.545 $X2=0 $Y2=0
cc_218 N_A_c_317_n N_VGND_c_425_n 0.00549284f $X=2.565 $Y=0.73 $X2=0 $Y2=0
cc_219 N_A_c_318_n N_VGND_c_425_n 4.17622e-19 $X=2.745 $Y=0.805 $X2=0 $Y2=0
cc_220 N_A_c_317_n N_VGND_c_426_n 0.00751205f $X=2.565 $Y=0.73 $X2=0 $Y2=0
cc_221 X N_VPWR_c_376_n 0.0494176f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_222 X N_VPWR_c_383_n 0.0240548f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_223 X N_VPWR_c_375_n 0.0137416f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_224 N_X_c_353_n N_VGND_c_423_n 0.0109108f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_225 N_X_c_353_n N_VGND_c_424_n 0.0205268f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_226 N_X_M1005_s N_VGND_c_426_n 0.00232985f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_227 N_X_c_353_n N_VGND_c_426_n 0.0130725f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_228 A_114_47# N_VGND_c_426_n 0.00490351f $X=0.57 $Y=0.235 $X2=3.12 $Y2=0
cc_229 N_VGND_c_426_n A_294_47# 0.00327011f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_230 N_VGND_c_426_n A_372_47# 0.00327011f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_231 N_VGND_c_426_n A_450_47# 0.00327011f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
