* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__lsbufiso1p_lp A DESTPWR DESTVPB SLEEP VGND VPB VPWR X
M1000 a_278_718# A a_206_718# VGND nshort w=840000u l=150000u
+  ad=4.578e+11p pd=4.45e+06u as=1.764e+11p ps=2.1e+06u
M1001 a_364_718# a_278_47# a_278_718# VGND nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1002 a_717_1085# SLEEP DESTPWR DESTVPB phighvt w=1e+06u l=150000u
+  ad=2.1e+11p pd=2.42e+06u as=5.6e+11p ps=5.12e+06u
M1003 a_517_420# SLEEP a_717_1085# DESTVPB phighvt w=1e+06u l=150000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1004 a_278_47# A a_206_47# VPB phighvt w=1e+06u l=150000u
+  ad=2.65e+11p pd=2.53e+06u as=2.1e+11p ps=2.42e+06u
M1005 DESTPWR a_517_420# a_1033_1085# DESTVPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.1e+11p ps=2.42e+06u
M1006 a_206_718# A a_123_718# VGND nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1007 a_364_1085# a_123_718# a_278_1085# DESTVPB phighvt w=1e+06u l=150000u
+  ad=2.1e+11p pd=2.42e+06u as=5.5e+11p ps=5.1e+06u
M1008 a_176_987# a_123_718# a_364_1085# DESTVPB phighvt w=1e+06u l=150000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1009 X a_123_718# a_1191_718# VGND nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=1.764e+11p ps=2.1e+06u
M1010 a_278_47# A a_206_446# VGND nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1011 a_206_47# A VPWR VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1012 a_1191_718# a_517_420# VGND VGND nshort w=840000u l=150000u
+  ad=0p pd=0u as=7.014e+11p ps=7.24e+06u
M1013 a_517_420# SLEEP a_631_802# VGND nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1014 a_206_446# A VGND VGND nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 DESTPWR SLEEP a_278_1085# DESTVPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_123_718# a_1191_1085# DESTVPB phighvt w=1e+06u l=150000u
+  ad=5.5e+11p pd=5.1e+06u as=2.1e+11p ps=2.42e+06u
M1017 a_1191_1085# a_123_718# DESTPWR DESTVPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_631_802# SLEEP VGND VGND nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_278_1085# a_176_987# a_206_1085# DESTVPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.1e+11p ps=2.42e+06u
M1020 a_206_1085# a_176_987# a_123_718# DESTVPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1021 a_1033_1085# a_517_420# X DESTVPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_176_987# a_278_47# a_364_718# VGND nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1023 VGND a_517_420# a_278_718# VGND nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
