* File: sky130_fd_sc_lp__lsbufiso1p_lp.spice
* Created: Fri Aug 28 10:42:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__lsbufiso1p_lp.pex.spice"
.subckt sky130_fd_sc_lp__lsbufiso1p_lp  VGND VPB DESTVPB A SLEEP VPWR DESTPWR X
* 
* X	X
* DESTPWR	DESTPWR
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* DESTVPB	DESTVPB
* VPB	VPB
* VGND	VGND
MM1014 A_206_446# N_A_M1014_g N_VGND_M1014_s N_VGND_M1014_b NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 A_206_718# N_A_M1006_g N_A_123_718#_M1006_s N_VGND_M1014_b NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1010 N_A_278_47#_M1010_d N_A_M1010_g A_206_446# N_VGND_M1014_b NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_278_718#_M1000_d N_A_M1000_g A_206_718# N_VGND_M1014_b NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.0882 PD=1.12 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1001 A_364_718# N_A_278_47#_M1001_g N_A_278_718#_M1000_d N_VGND_M1014_b NSHORT
+ L=0.15 W=0.84 AD=0.0882 AS=0.1176 PD=1.05 PS=1.12 NRD=7.14 NRS=0 M=1 R=5.6
+ SA=75001 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1022 N_A_176_987#_M1022_d N_A_278_47#_M1022_g A_364_718# N_VGND_M1014_b NSHORT
+ L=0.15 W=0.84 AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6
+ SA=75001.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1023 N_VGND_M1023_d N_A_517_420#_M1023_g N_A_278_718#_M1023_s N_VGND_M1014_b
+ NSHORT L=0.15 W=0.84 AD=0.2394 AS=0.2226 PD=2.25 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1018 A_631_802# N_SLEEP_M1018_g N_VGND_M1018_s N_VGND_M1014_b NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_517_420#_M1013_d N_SLEEP_M1013_g A_631_802# N_VGND_M1014_b NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 A_1191_718# N_A_517_420#_M1012_g N_VGND_M1012_s N_VGND_M1014_b NSHORT
+ L=0.15 W=0.84 AD=0.0882 AS=0.2394 PD=1.05 PS=2.25 NRD=7.14 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_X_M1009_d N_A_123_718#_M1009_g A_1191_718# N_VGND_M1014_b NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 A_206_47# N_A_M1011_g N_VPWR_M1011_s N_VPB_M1011_b PHIGHVT L=0.15 W=1
+ AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=9.8303 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75000.5 A=0.15 P=2.3 MULT=1
MM1020 A_206_1085# N_A_176_987#_M1020_g N_A_123_718#_M1020_s N_DESTVPB_M1020_b
+ PHIGHVT L=0.15 W=1 AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=9.8303 NRS=0 M=1
+ R=6.66667 SA=75000.2 SB=75001.4 A=0.15 P=2.3 MULT=1
MM1004 N_A_278_47#_M1004_d N_A_M1004_g A_206_47# N_VPB_M1011_b PHIGHVT L=0.15
+ W=1 AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667
+ SA=75000.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1019 N_A_278_1085#_M1019_d N_A_176_987#_M1019_g A_206_1085# N_DESTVPB_M1020_b
+ PHIGHVT L=0.15 W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=9.8303 M=1
+ R=6.66667 SA=75000.5 SB=75001 A=0.15 P=2.3 MULT=1
MM1007 A_364_1085# N_A_123_718#_M1007_g N_A_278_1085#_M1019_d N_DESTVPB_M1020_b
+ PHIGHVT L=0.15 W=1 AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=9.8303 NRS=0 M=1
+ R=6.66667 SA=75001 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1008 N_A_176_987#_M1008_d N_A_123_718#_M1008_g A_364_1085# N_DESTVPB_M1020_b
+ PHIGHVT L=0.15 W=1 AD=0.285 AS=0.105 PD=2.57 PS=1.21 NRD=0 NRS=9.8303 M=1
+ R=6.66667 SA=75001.3 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1015 N_DESTPWR_M1015_d N_SLEEP_M1015_g N_A_278_1085#_M1015_s N_DESTVPB_M1020_b
+ PHIGHVT L=0.15 W=1 AD=0.14 AS=0.27 PD=1.28 PS=2.54 NRD=0 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001 A=0.15 P=2.3 MULT=1
MM1002 A_717_1085# N_SLEEP_M1002_g N_DESTPWR_M1015_d N_DESTVPB_M1020_b PHIGHVT
+ L=0.15 W=1 AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=9.8303 NRS=0 M=1 R=6.66667
+ SA=75000.6 SB=75000.6 A=0.15 P=2.3 MULT=1
MM1003 N_A_517_420#_M1003_d N_SLEEP_M1003_g A_717_1085# N_DESTVPB_M1020_b
+ PHIGHVT L=0.15 W=1 AD=0.285 AS=0.105 PD=2.57 PS=1.21 NRD=0 NRS=9.8303 M=1
+ R=6.66667 SA=75001 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1021 A_1033_1085# N_A_517_420#_M1021_g N_X_M1021_s N_DESTVPB_M1020_b PHIGHVT
+ L=0.15 W=1 AD=0.105 AS=0.285 PD=1.21 PS=2.57 NRD=9.8303 NRS=0 M=1 R=6.66667
+ SA=75000.2 SB=75001.3 A=0.15 P=2.3 MULT=1
MM1005 N_DESTPWR_M1005_d N_A_517_420#_M1005_g A_1033_1085# N_DESTVPB_M1020_b
+ PHIGHVT L=0.15 W=1 AD=0.14 AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=9.8303 M=1
+ R=6.66667 SA=75000.6 SB=75001 A=0.15 P=2.3 MULT=1
MM1017 A_1191_1085# N_A_123_718#_M1017_g N_DESTPWR_M1005_d N_DESTVPB_M1020_b
+ PHIGHVT L=0.15 W=1 AD=0.105 AS=0.14 PD=1.21 PS=1.28 NRD=9.8303 NRS=0 M=1
+ R=6.66667 SA=75001 SB=75000.5 A=0.15 P=2.3 MULT=1
MM1016 N_X_M1016_d N_A_123_718#_M1016_g A_1191_1085# N_DESTVPB_M1020_b PHIGHVT
+ L=0.15 W=1 AD=0.265 AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=9.8303 M=1 R=6.66667
+ SA=75001.4 SB=75000.2 A=0.15 P=2.3 MULT=1
DX24_noxref N_VGND_M1014_b N_VPB_M1011_b NWDIODE A=13.5212 P=18.23
DX25_noxref N_VGND_M1014_b N_DESTVPB_M1020_b NWDIODE A=13.5212 P=18.23
*
.include "sky130_fd_sc_lp__lsbufiso1p_lp.pxi.spice"
*
.ends
*
*
