* File: sky130_fd_sc_lp__a41o_0.pxi.spice
* Created: Fri Aug 28 10:02:23 2020
* 
x_PM_SKY130_FD_SC_LP__A41O_0%A_80_309# N_A_80_309#_M1006_d N_A_80_309#_M1008_s
+ N_A_80_309#_c_100_n N_A_80_309#_M1001_g N_A_80_309#_M1002_g
+ N_A_80_309#_c_102_n N_A_80_309#_c_103_n N_A_80_309#_c_94_n N_A_80_309#_c_95_n
+ N_A_80_309#_c_104_n N_A_80_309#_c_105_n N_A_80_309#_c_106_n N_A_80_309#_c_96_n
+ N_A_80_309#_c_97_n N_A_80_309#_c_98_n N_A_80_309#_c_99_n N_A_80_309#_c_133_p
+ PM_SKY130_FD_SC_LP__A41O_0%A_80_309#
x_PM_SKY130_FD_SC_LP__A41O_0%B1 N_B1_M1006_g N_B1_c_176_n N_B1_M1008_g
+ N_B1_c_172_n N_B1_c_173_n N_B1_c_179_n B1 B1 N_B1_c_175_n
+ PM_SKY130_FD_SC_LP__A41O_0%B1
x_PM_SKY130_FD_SC_LP__A41O_0%A1 N_A1_M1011_g N_A1_M1005_g N_A1_c_227_n
+ N_A1_c_232_n A1 A1 A1 N_A1_c_229_n PM_SKY130_FD_SC_LP__A41O_0%A1
x_PM_SKY130_FD_SC_LP__A41O_0%A2 N_A2_M1007_g N_A2_M1000_g N_A2_c_278_n
+ N_A2_c_279_n N_A2_c_280_n A2 A2 A2 A2 N_A2_c_282_n
+ PM_SKY130_FD_SC_LP__A41O_0%A2
x_PM_SKY130_FD_SC_LP__A41O_0%A3 N_A3_M1003_g N_A3_c_325_n N_A3_M1009_g
+ N_A3_c_326_n A3 A3 A3 N_A3_c_328_n PM_SKY130_FD_SC_LP__A41O_0%A3
x_PM_SKY130_FD_SC_LP__A41O_0%A4 N_A4_c_366_n N_A4_M1004_g N_A4_M1010_g
+ N_A4_c_367_n N_A4_c_368_n N_A4_c_374_n N_A4_c_369_n A4 A4 A4 N_A4_c_371_n
+ PM_SKY130_FD_SC_LP__A41O_0%A4
x_PM_SKY130_FD_SC_LP__A41O_0%X N_X_M1002_s N_X_M1001_s X X X X X X X N_X_c_408_n
+ N_X_c_406_n X PM_SKY130_FD_SC_LP__A41O_0%X
x_PM_SKY130_FD_SC_LP__A41O_0%VPWR N_VPWR_M1001_d N_VPWR_M1005_d N_VPWR_M1009_d
+ N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n
+ VPWR N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_423_n
+ N_VPWR_c_433_n N_VPWR_c_434_n PM_SKY130_FD_SC_LP__A41O_0%VPWR
x_PM_SKY130_FD_SC_LP__A41O_0%A_321_473# N_A_321_473#_M1008_d
+ N_A_321_473#_M1000_d N_A_321_473#_M1010_d N_A_321_473#_c_473_n
+ N_A_321_473#_c_474_n N_A_321_473#_c_475_n N_A_321_473#_c_476_n
+ N_A_321_473#_c_477_n N_A_321_473#_c_478_n N_A_321_473#_c_479_n
+ PM_SKY130_FD_SC_LP__A41O_0%A_321_473#
x_PM_SKY130_FD_SC_LP__A41O_0%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_c_518_n
+ N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n
+ VGND N_VGND_c_524_n N_VGND_c_525_n PM_SKY130_FD_SC_LP__A41O_0%VGND
cc_1 VNB N_A_80_309#_M1002_g 0.063893f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.445
cc_2 VNB N_A_80_309#_c_94_n 0.00960329f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=0.825
cc_3 VNB N_A_80_309#_c_95_n 0.00219325f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.825
cc_4 VNB N_A_80_309#_c_96_n 0.0019275f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=0.74
cc_5 VNB N_A_80_309#_c_97_n 0.00345798f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.71
cc_6 VNB N_A_80_309#_c_98_n 0.0166659f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.71
cc_7 VNB N_A_80_309#_c_99_n 0.0114255f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.545
cc_8 VNB N_B1_M1006_g 0.0370093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_172_n 0.0221031f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.545
cc_10 VNB N_B1_c_173_n 0.00450606f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.445
cc_11 VNB B1 0.00591895f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.045
cc_12 VNB N_B1_c_175_n 0.0164755f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.13
cc_13 VNB N_A1_M1011_g 0.0403657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_227_n 0.024595f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.725
cc_15 VNB A1 0.00524554f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.545
cc_16 VNB N_A1_c_229_n 0.0192441f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.91
cc_17 VNB N_A2_M1000_g 0.0108404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_278_n 0.0163723f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.215
cc_19 VNB N_A2_c_279_n 0.0209075f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.725
cc_20 VNB N_A2_c_280_n 0.0153438f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.725
cc_21 VNB A2 0.00629845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_c_282_n 0.0160353f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.545
cc_23 VNB N_A3_M1003_g 0.03492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A3_c_325_n 0.0208835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A3_c_326_n 6.78035e-19 $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.725
cc_26 VNB A3 0.00840684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A3_c_328_n 0.0181985f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.045
cc_28 VNB N_A4_c_366_n 0.0206184f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.235
cc_29 VNB N_A4_c_367_n 0.00907722f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.215
cc_30 VNB N_A4_c_368_n 0.0373297f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.545
cc_31 VNB N_A4_c_369_n 0.0187513f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.91
cc_32 VNB A4 0.035726f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.545
cc_33 VNB N_A4_c_371_n 0.0368995f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=2.51
cc_34 VNB X 0.0559629f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.722
cc_35 VNB N_X_c_406_n 0.017882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_423_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_518_n 0.00519343f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.215
cc_38 VNB N_VGND_c_519_n 0.0182436f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.545
cc_39 VNB N_VGND_c_520_n 0.0213005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_521_n 0.004878f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=2.215
cc_41 VNB N_VGND_c_522_n 0.0579646f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.045
cc_42 VNB N_VGND_c_523_n 0.00621103f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.91
cc_43 VNB N_VGND_c_524_n 0.0120081f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.71
cc_44 VNB N_VGND_c_525_n 0.211918f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.545
cc_45 VPB N_A_80_309#_c_100_n 0.0246489f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=2.038
cc_46 VPB N_A_80_309#_M1001_g 0.0280249f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.725
cc_47 VPB N_A_80_309#_c_102_n 0.0198331f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=2.215
cc_48 VPB N_A_80_309#_c_103_n 0.00305146f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.045
cc_49 VPB N_A_80_309#_c_104_n 0.0178059f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=2.13
cc_50 VPB N_A_80_309#_c_105_n 0.00482188f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=2.13
cc_51 VPB N_A_80_309#_c_106_n 0.0128017f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=2.51
cc_52 VPB N_A_80_309#_c_97_n 5.04473e-19 $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.71
cc_53 VPB N_A_80_309#_c_98_n 0.00486145f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.71
cc_54 VPB N_B1_c_176_n 0.0192409f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B1_M1008_g 0.0216357f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_56 VPB N_B1_c_173_n 0.0112454f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=0.445
cc_57 VPB N_B1_c_179_n 0.0313831f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=2.215
cc_58 VPB B1 0.00309378f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.045
cc_59 VPB N_A1_M1005_g 0.0406786f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_60 VPB N_A1_c_227_n 0.00150301f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.725
cc_61 VPB N_A1_c_232_n 0.0261805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB A1 0.00276112f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.545
cc_63 VPB N_A2_M1000_g 0.0465733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB A2 0.00274746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A3_M1009_g 0.0402437f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_66 VPB N_A3_c_326_n 0.0173646f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.725
cc_67 VPB A3 0.00401886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A4_M1010_g 0.0229278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A4_c_367_n 0.0298367f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_70 VPB N_A4_c_374_n 0.0169855f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=2.215
cc_71 VPB A4 0.0133476f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1.545
cc_72 VPB X 0.037593f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.722
cc_73 VPB N_X_c_408_n 0.0229413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB X 0.00835826f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_424_n 0.0165813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_425_n 0.00981896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_426_n 0.0100229f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.91
cc_78 VPB N_VPWR_c_427_n 0.0166607f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=0.825
cc_79 VPB N_VPWR_c_428_n 0.00555219f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=2.13
cc_80 VPB N_VPWR_c_429_n 0.0171682f $X=-0.19 $Y=1.655 $X2=1.297 $Y2=2.51
cc_81 VPB N_VPWR_c_430_n 0.032936f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.71
cc_82 VPB N_VPWR_c_431_n 0.0203278f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.545
cc_83 VPB N_VPWR_c_423_n 0.0751285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_433_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_434_n 0.00507132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_321_473#_c_473_n 0.00561114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_321_473#_c_474_n 0.00647708f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=0.445
cc_88 VPB N_A_321_473#_c_475_n 0.003515f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=0.445
cc_89 VPB N_A_321_473#_c_476_n 0.0055099f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.74
cc_90 VPB N_A_321_473#_c_477_n 0.0180476f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.91
cc_91 VPB N_A_321_473#_c_478_n 0.0360849f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=2.13
cc_92 VPB N_A_321_473#_c_479_n 0.0087752f $X=-0.19 $Y=1.655 $X2=1.297 $Y2=2.215
cc_93 N_A_80_309#_M1002_g N_B1_M1006_g 0.0261432f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_80_309#_c_94_n N_B1_M1006_g 0.0146897f $X=1.165 $Y=0.825 $X2=0 $Y2=0
cc_95 N_A_80_309#_c_96_n N_B1_M1006_g 0.00275763f $X=1.29 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A_80_309#_c_99_n N_B1_M1006_g 0.0037634f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_97 N_A_80_309#_c_100_n N_B1_c_176_n 0.00574679f $X=0.577 $Y=2.038 $X2=0 $Y2=0
cc_98 N_A_80_309#_c_103_n N_B1_c_176_n 0.0050709f $X=0.7 $Y=2.045 $X2=0 $Y2=0
cc_99 N_A_80_309#_c_104_n N_B1_c_176_n 0.00324623f $X=1.15 $Y=2.13 $X2=0 $Y2=0
cc_100 N_A_80_309#_c_106_n N_B1_M1008_g 0.00398238f $X=1.315 $Y=2.51 $X2=0 $Y2=0
cc_101 N_A_80_309#_c_97_n N_B1_c_172_n 0.00155952f $X=0.59 $Y=1.71 $X2=0 $Y2=0
cc_102 N_A_80_309#_c_98_n N_B1_c_172_n 0.00532237f $X=0.59 $Y=1.71 $X2=0 $Y2=0
cc_103 N_A_80_309#_c_100_n N_B1_c_173_n 0.00532237f $X=0.577 $Y=2.038 $X2=0
+ $Y2=0
cc_104 N_A_80_309#_c_103_n N_B1_c_173_n 0.00155952f $X=0.7 $Y=2.045 $X2=0 $Y2=0
cc_105 N_A_80_309#_c_104_n N_B1_c_173_n 0.00319316f $X=1.15 $Y=2.13 $X2=0 $Y2=0
cc_106 N_A_80_309#_c_102_n N_B1_c_179_n 0.00574679f $X=0.577 $Y=2.215 $X2=0
+ $Y2=0
cc_107 N_A_80_309#_c_104_n N_B1_c_179_n 0.015899f $X=1.15 $Y=2.13 $X2=0 $Y2=0
cc_108 N_A_80_309#_c_100_n B1 2.19503e-19 $X=0.577 $Y=2.038 $X2=0 $Y2=0
cc_109 N_A_80_309#_c_94_n B1 0.0244269f $X=1.165 $Y=0.825 $X2=0 $Y2=0
cc_110 N_A_80_309#_c_104_n B1 0.0215596f $X=1.15 $Y=2.13 $X2=0 $Y2=0
cc_111 N_A_80_309#_c_99_n B1 0.0575644f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_112 N_A_80_309#_M1002_g N_B1_c_175_n 0.0182165f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_80_309#_c_94_n N_B1_c_175_n 0.00164565f $X=1.165 $Y=0.825 $X2=0 $Y2=0
cc_114 N_A_80_309#_c_99_n N_B1_c_175_n 0.00155952f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_115 N_A_80_309#_c_94_n N_A1_M1011_g 7.85718e-19 $X=1.165 $Y=0.825 $X2=0 $Y2=0
cc_116 N_A_80_309#_c_96_n N_A1_M1011_g 0.00116945f $X=1.29 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A_80_309#_c_133_p N_A1_M1011_g 0.00504314f $X=1.635 $Y=0.445 $X2=0
+ $Y2=0
cc_118 N_A_80_309#_c_94_n A1 0.0116577f $X=1.165 $Y=0.825 $X2=0 $Y2=0
cc_119 N_A_80_309#_c_133_p A1 0.0145962f $X=1.635 $Y=0.445 $X2=0 $Y2=0
cc_120 N_A_80_309#_c_133_p N_A1_c_229_n 0.00142678f $X=1.635 $Y=0.445 $X2=0
+ $Y2=0
cc_121 N_A_80_309#_c_133_p N_A2_c_278_n 6.627e-19 $X=1.635 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_80_309#_c_94_n A2 0.00110837f $X=1.165 $Y=0.825 $X2=0 $Y2=0
cc_123 N_A_80_309#_c_96_n A2 0.00458747f $X=1.29 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A_80_309#_c_133_p A2 0.0150333f $X=1.635 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_80_309#_M1002_g X 0.019999f $X=0.65 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_80_309#_c_95_n X 0.00748974f $X=0.895 $Y=0.825 $X2=0 $Y2=0
cc_127 N_A_80_309#_c_105_n X 0.0139714f $X=0.895 $Y=2.13 $X2=0 $Y2=0
cc_128 N_A_80_309#_c_97_n X 0.0390399f $X=0.59 $Y=1.71 $X2=0 $Y2=0
cc_129 N_A_80_309#_c_98_n X 0.024186f $X=0.59 $Y=1.71 $X2=0 $Y2=0
cc_130 N_A_80_309#_c_99_n X 0.0275989f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_131 N_A_80_309#_M1001_g X 9.38286e-19 $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_132 N_A_80_309#_M1001_g N_VPWR_c_424_n 0.00515749f $X=0.475 $Y=2.725 $X2=0
+ $Y2=0
cc_133 N_A_80_309#_c_102_n N_VPWR_c_424_n 0.00151751f $X=0.577 $Y=2.215 $X2=0
+ $Y2=0
cc_134 N_A_80_309#_c_105_n N_VPWR_c_424_n 0.0265564f $X=0.895 $Y=2.13 $X2=0
+ $Y2=0
cc_135 N_A_80_309#_c_106_n N_VPWR_c_424_n 0.0357486f $X=1.315 $Y=2.51 $X2=0
+ $Y2=0
cc_136 N_A_80_309#_M1001_g N_VPWR_c_429_n 0.0053602f $X=0.475 $Y=2.725 $X2=0
+ $Y2=0
cc_137 N_A_80_309#_c_106_n N_VPWR_c_430_n 0.0159397f $X=1.315 $Y=2.51 $X2=0
+ $Y2=0
cc_138 N_A_80_309#_M1001_g N_VPWR_c_423_n 0.01173f $X=0.475 $Y=2.725 $X2=0 $Y2=0
cc_139 N_A_80_309#_c_106_n N_VPWR_c_423_n 0.0111051f $X=1.315 $Y=2.51 $X2=0
+ $Y2=0
cc_140 N_A_80_309#_c_104_n N_A_321_473#_c_473_n 0.00325194f $X=1.15 $Y=2.13
+ $X2=0 $Y2=0
cc_141 N_A_80_309#_c_106_n N_A_321_473#_c_473_n 0.0135529f $X=1.315 $Y=2.51
+ $X2=0 $Y2=0
cc_142 N_A_80_309#_c_104_n N_A_321_473#_c_475_n 0.0116792f $X=1.15 $Y=2.13 $X2=0
+ $Y2=0
cc_143 N_A_80_309#_M1002_g N_VGND_c_518_n 0.0030614f $X=0.65 $Y=0.445 $X2=0
+ $Y2=0
cc_144 N_A_80_309#_c_94_n N_VGND_c_518_n 0.00580777f $X=1.165 $Y=0.825 $X2=0
+ $Y2=0
cc_145 N_A_80_309#_c_95_n N_VGND_c_518_n 0.0117747f $X=0.895 $Y=0.825 $X2=0
+ $Y2=0
cc_146 N_A_80_309#_M1002_g N_VGND_c_520_n 0.00585385f $X=0.65 $Y=0.445 $X2=0
+ $Y2=0
cc_147 N_A_80_309#_c_95_n N_VGND_c_520_n 2.40268e-19 $X=0.895 $Y=0.825 $X2=0
+ $Y2=0
cc_148 N_A_80_309#_c_94_n N_VGND_c_522_n 0.00222198f $X=1.165 $Y=0.825 $X2=0
+ $Y2=0
cc_149 N_A_80_309#_c_133_p N_VGND_c_522_n 0.03344f $X=1.635 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_80_309#_M1006_d N_VGND_c_525_n 0.00513926f $X=1.155 $Y=0.235 $X2=0
+ $Y2=0
cc_151 N_A_80_309#_M1002_g N_VGND_c_525_n 0.0118122f $X=0.65 $Y=0.445 $X2=0
+ $Y2=0
cc_152 N_A_80_309#_c_94_n N_VGND_c_525_n 0.00405009f $X=1.165 $Y=0.825 $X2=0
+ $Y2=0
cc_153 N_A_80_309#_c_95_n N_VGND_c_525_n 0.00105576f $X=0.895 $Y=0.825 $X2=0
+ $Y2=0
cc_154 N_A_80_309#_c_133_p N_VGND_c_525_n 0.023753f $X=1.635 $Y=0.445 $X2=0
+ $Y2=0
cc_155 N_B1_M1006_g N_A1_M1011_g 0.00809117f $X=1.08 $Y=0.445 $X2=0 $Y2=0
cc_156 B1 N_A1_M1011_g 2.08568e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_157 N_B1_c_175_n N_A1_M1011_g 0.0017201f $X=1.16 $Y=1.245 $X2=0 $Y2=0
cc_158 N_B1_c_176_n N_A1_M1005_g 0.00559378f $X=1.25 $Y=2.065 $X2=0 $Y2=0
cc_159 N_B1_c_179_n N_A1_M1005_g 0.0174007f $X=1.53 $Y=2.14 $X2=0 $Y2=0
cc_160 N_B1_c_172_n N_A1_c_227_n 0.0119085f $X=1.16 $Y=1.585 $X2=0 $Y2=0
cc_161 N_B1_c_173_n N_A1_c_232_n 0.0119085f $X=1.16 $Y=1.75 $X2=0 $Y2=0
cc_162 N_B1_c_179_n N_A1_c_232_n 0.00279326f $X=1.53 $Y=2.14 $X2=0 $Y2=0
cc_163 N_B1_M1006_g A1 0.00343054f $X=1.08 $Y=0.445 $X2=0 $Y2=0
cc_164 N_B1_c_179_n A1 2.37496e-19 $X=1.53 $Y=2.14 $X2=0 $Y2=0
cc_165 B1 A1 0.0462872f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_166 N_B1_c_175_n A1 0.00103107f $X=1.16 $Y=1.245 $X2=0 $Y2=0
cc_167 B1 N_A1_c_229_n 0.00434954f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_168 N_B1_c_175_n N_A1_c_229_n 0.0119085f $X=1.16 $Y=1.245 $X2=0 $Y2=0
cc_169 N_B1_M1008_g N_VPWR_c_424_n 0.00328525f $X=1.53 $Y=2.685 $X2=0 $Y2=0
cc_170 N_B1_M1008_g N_VPWR_c_430_n 0.00499542f $X=1.53 $Y=2.685 $X2=0 $Y2=0
cc_171 N_B1_M1008_g N_VPWR_c_423_n 0.0104152f $X=1.53 $Y=2.685 $X2=0 $Y2=0
cc_172 N_B1_c_179_n N_A_321_473#_c_473_n 0.00171168f $X=1.53 $Y=2.14 $X2=0 $Y2=0
cc_173 N_B1_c_176_n N_A_321_473#_c_475_n 0.0011152f $X=1.25 $Y=2.065 $X2=0 $Y2=0
cc_174 N_B1_c_179_n N_A_321_473#_c_475_n 0.00111345f $X=1.53 $Y=2.14 $X2=0 $Y2=0
cc_175 N_B1_M1006_g N_VGND_c_518_n 0.00309118f $X=1.08 $Y=0.445 $X2=0 $Y2=0
cc_176 N_B1_M1006_g N_VGND_c_522_n 0.00439878f $X=1.08 $Y=0.445 $X2=0 $Y2=0
cc_177 N_B1_M1006_g N_VGND_c_525_n 0.00668005f $X=1.08 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A1_c_227_n N_A2_M1000_g 0.00636276f $X=1.8 $Y=1.675 $X2=0 $Y2=0
cc_179 N_A1_c_232_n N_A2_M1000_g 0.0365108f $X=1.8 $Y=1.825 $X2=0 $Y2=0
cc_180 A1 N_A2_M1000_g 2.71485e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_181 N_A1_M1011_g N_A2_c_278_n 0.0254853f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_182 N_A1_c_229_n N_A2_c_279_n 0.013384f $X=1.73 $Y=1.32 $X2=0 $Y2=0
cc_183 N_A1_c_227_n N_A2_c_280_n 0.013384f $X=1.8 $Y=1.675 $X2=0 $Y2=0
cc_184 N_A1_M1011_g A2 0.0106286f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A1_M1005_g A2 4.94343e-19 $X=1.96 $Y=2.685 $X2=0 $Y2=0
cc_186 N_A1_c_232_n A2 0.00479929f $X=1.8 $Y=1.825 $X2=0 $Y2=0
cc_187 A1 A2 0.0825842f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_188 N_A1_M1011_g N_A2_c_282_n 0.013384f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_189 A1 N_A2_c_282_n 5.71963e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_190 N_A1_M1005_g N_VPWR_c_425_n 0.00315007f $X=1.96 $Y=2.685 $X2=0 $Y2=0
cc_191 N_A1_M1005_g N_VPWR_c_430_n 0.00499542f $X=1.96 $Y=2.685 $X2=0 $Y2=0
cc_192 N_A1_M1005_g N_VPWR_c_423_n 0.00971452f $X=1.96 $Y=2.685 $X2=0 $Y2=0
cc_193 N_A1_M1005_g N_A_321_473#_c_473_n 0.00272746f $X=1.96 $Y=2.685 $X2=0
+ $Y2=0
cc_194 N_A1_M1005_g N_A_321_473#_c_474_n 0.0184889f $X=1.96 $Y=2.685 $X2=0 $Y2=0
cc_195 N_A1_c_232_n N_A_321_473#_c_474_n 5.98754e-19 $X=1.8 $Y=1.825 $X2=0 $Y2=0
cc_196 N_A1_c_232_n N_A_321_473#_c_475_n 0.00318797f $X=1.8 $Y=1.825 $X2=0 $Y2=0
cc_197 A1 N_A_321_473#_c_475_n 0.0209841f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_198 N_A1_M1011_g N_VGND_c_522_n 0.0054833f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_199 N_A1_M1011_g N_VGND_c_525_n 0.0096471f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_200 A1 N_VGND_c_525_n 0.00174213f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_201 N_A2_c_278_n N_A3_M1003_g 0.0299133f $X=2.3 $Y=0.765 $X2=0 $Y2=0
cc_202 A2 N_A3_M1003_g 0.00573087f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_203 N_A2_c_282_n N_A3_M1003_g 0.0160567f $X=2.3 $Y=0.93 $X2=0 $Y2=0
cc_204 N_A2_c_280_n N_A3_c_325_n 0.0160567f $X=2.3 $Y=1.435 $X2=0 $Y2=0
cc_205 N_A2_M1000_g N_A3_M1009_g 0.0290211f $X=2.39 $Y=2.685 $X2=0 $Y2=0
cc_206 N_A2_M1000_g N_A3_c_326_n 0.0160567f $X=2.39 $Y=2.685 $X2=0 $Y2=0
cc_207 A2 A3 0.0408233f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_208 N_A2_c_282_n A3 0.00310096f $X=2.3 $Y=0.93 $X2=0 $Y2=0
cc_209 N_A2_c_279_n N_A3_c_328_n 0.0160567f $X=2.3 $Y=1.27 $X2=0 $Y2=0
cc_210 N_A2_M1000_g N_VPWR_c_425_n 0.00179007f $X=2.39 $Y=2.685 $X2=0 $Y2=0
cc_211 N_A2_M1000_g N_VPWR_c_427_n 0.00499542f $X=2.39 $Y=2.685 $X2=0 $Y2=0
cc_212 N_A2_M1000_g N_VPWR_c_423_n 0.00972572f $X=2.39 $Y=2.685 $X2=0 $Y2=0
cc_213 N_A2_M1000_g N_A_321_473#_c_474_n 0.0174517f $X=2.39 $Y=2.685 $X2=0 $Y2=0
cc_214 N_A2_c_280_n N_A_321_473#_c_474_n 5.47318e-19 $X=2.3 $Y=1.435 $X2=0 $Y2=0
cc_215 A2 N_A_321_473#_c_474_n 0.0307332f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_216 N_A2_M1000_g N_A_321_473#_c_476_n 0.00275529f $X=2.39 $Y=2.685 $X2=0
+ $Y2=0
cc_217 N_A2_c_278_n N_VGND_c_522_n 0.00384725f $X=2.3 $Y=0.765 $X2=0 $Y2=0
cc_218 A2 N_VGND_c_522_n 0.0128989f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_219 N_A2_c_282_n N_VGND_c_522_n 0.00183649f $X=2.3 $Y=0.93 $X2=0 $Y2=0
cc_220 N_A2_c_278_n N_VGND_c_525_n 0.00566682f $X=2.3 $Y=0.765 $X2=0 $Y2=0
cc_221 A2 N_VGND_c_525_n 0.0127525f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_222 N_A2_c_282_n N_VGND_c_525_n 0.00213786f $X=2.3 $Y=0.93 $X2=0 $Y2=0
cc_223 A2 A_385_47# 0.00531707f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_224 N_A3_M1003_g N_A4_c_366_n 0.0511956f $X=2.75 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_225 N_A3_M1009_g N_A4_c_367_n 0.00800061f $X=2.82 $Y=2.685 $X2=0 $Y2=0
cc_226 N_A3_c_326_n N_A4_c_367_n 0.00969829f $X=2.855 $Y=1.825 $X2=0 $Y2=0
cc_227 A3 N_A4_c_368_n 0.013731f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_228 N_A3_M1009_g N_A4_c_374_n 0.0161932f $X=2.82 $Y=2.685 $X2=0 $Y2=0
cc_229 N_A3_c_325_n N_A4_c_369_n 0.00969829f $X=2.855 $Y=1.645 $X2=0 $Y2=0
cc_230 N_A3_M1003_g A4 2.27792e-19 $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_231 A3 A4 0.0852459f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_232 N_A3_c_328_n A4 5.54225e-19 $X=2.87 $Y=1.32 $X2=0 $Y2=0
cc_233 N_A3_M1003_g N_A4_c_371_n 0.00455089f $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_234 A3 N_A4_c_371_n 0.00747825f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_235 N_A3_c_328_n N_A4_c_371_n 0.00969829f $X=2.87 $Y=1.32 $X2=0 $Y2=0
cc_236 N_A3_M1009_g N_VPWR_c_426_n 0.00188236f $X=2.82 $Y=2.685 $X2=0 $Y2=0
cc_237 N_A3_M1009_g N_VPWR_c_427_n 0.00499542f $X=2.82 $Y=2.685 $X2=0 $Y2=0
cc_238 N_A3_M1009_g N_VPWR_c_423_n 0.00973735f $X=2.82 $Y=2.685 $X2=0 $Y2=0
cc_239 N_A3_M1009_g N_A_321_473#_c_476_n 0.0027772f $X=2.82 $Y=2.685 $X2=0 $Y2=0
cc_240 N_A3_M1009_g N_A_321_473#_c_477_n 0.0165955f $X=2.82 $Y=2.685 $X2=0 $Y2=0
cc_241 N_A3_c_326_n N_A_321_473#_c_477_n 0.00156189f $X=2.855 $Y=1.825 $X2=0
+ $Y2=0
cc_242 A3 N_A_321_473#_c_477_n 0.0331587f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_243 N_A3_c_326_n N_A_321_473#_c_479_n 0.00263262f $X=2.855 $Y=1.825 $X2=0
+ $Y2=0
cc_244 N_A3_M1003_g N_VGND_c_519_n 0.00312909f $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_245 A3 N_VGND_c_519_n 0.00512795f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_246 N_A3_M1003_g N_VGND_c_522_n 0.00585385f $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_247 N_A3_M1003_g N_VGND_c_525_n 0.00966365f $X=2.75 $Y=0.445 $X2=0 $Y2=0
cc_248 A3 N_VGND_c_525_n 0.0138772f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_249 N_A4_M1010_g N_VPWR_c_426_n 0.00321847f $X=3.275 $Y=2.685 $X2=0 $Y2=0
cc_250 N_A4_M1010_g N_VPWR_c_431_n 0.00499542f $X=3.275 $Y=2.685 $X2=0 $Y2=0
cc_251 N_A4_M1010_g N_VPWR_c_423_n 0.0101262f $X=3.275 $Y=2.685 $X2=0 $Y2=0
cc_252 N_A4_c_367_n N_A_321_473#_c_477_n 0.00754492f $X=3.38 $Y=2.065 $X2=0
+ $Y2=0
cc_253 N_A4_c_374_n N_A_321_473#_c_477_n 0.0145833f $X=3.38 $Y=2.14 $X2=0 $Y2=0
cc_254 N_A4_c_369_n N_A_321_473#_c_477_n 7.05524e-19 $X=3.47 $Y=1.51 $X2=0 $Y2=0
cc_255 A4 N_A_321_473#_c_477_n 0.0245803f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_256 N_A4_M1010_g N_A_321_473#_c_478_n 0.00489157f $X=3.275 $Y=2.685 $X2=0
+ $Y2=0
cc_257 N_A4_c_374_n N_A_321_473#_c_478_n 0.00412141f $X=3.38 $Y=2.14 $X2=0 $Y2=0
cc_258 N_A4_c_366_n N_VGND_c_519_n 0.0145968f $X=3.11 $Y=0.765 $X2=0 $Y2=0
cc_259 N_A4_c_368_n N_VGND_c_519_n 0.0113852f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_260 A4 N_VGND_c_519_n 0.0122642f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_261 N_A4_c_366_n N_VGND_c_522_n 0.00388479f $X=3.11 $Y=0.765 $X2=0 $Y2=0
cc_262 N_A4_c_368_n N_VGND_c_524_n 0.00207886f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_263 N_A4_c_366_n N_VGND_c_525_n 0.00352586f $X=3.11 $Y=0.765 $X2=0 $Y2=0
cc_264 N_A4_c_368_n N_VGND_c_525_n 0.00283267f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_265 A4 N_VGND_c_525_n 0.00954475f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_266 X N_VPWR_c_424_n 0.00311658f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_267 N_X_c_408_n N_VPWR_c_429_n 0.0204296f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_268 N_X_c_408_n N_VPWR_c_423_n 0.011724f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_269 N_X_c_406_n N_VGND_c_520_n 0.0266288f $X=0.435 $Y=0.445 $X2=0 $Y2=0
cc_270 N_X_M1002_s N_VGND_c_525_n 0.00234325f $X=0.31 $Y=0.235 $X2=0 $Y2=0
cc_271 N_X_c_406_n N_VGND_c_525_n 0.018252f $X=0.435 $Y=0.445 $X2=0 $Y2=0
cc_272 N_VPWR_c_425_n N_A_321_473#_c_473_n 0.00304975f $X=2.175 $Y=2.51 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_430_n N_A_321_473#_c_473_n 0.0137636f $X=2.04 $Y=3.33 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_423_n N_A_321_473#_c_473_n 0.00958901f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_425_n N_A_321_473#_c_474_n 0.0222131f $X=2.175 $Y=2.51 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_425_n N_A_321_473#_c_476_n 0.00304975f $X=2.175 $Y=2.51 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_426_n N_A_321_473#_c_476_n 0.00307077f $X=3.035 $Y=2.51 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_427_n N_A_321_473#_c_476_n 0.0137636f $X=2.9 $Y=3.33 $X2=0 $Y2=0
cc_279 N_VPWR_c_423_n N_A_321_473#_c_476_n 0.00958901f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_426_n N_A_321_473#_c_477_n 0.0243245f $X=3.035 $Y=2.51 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_426_n N_A_321_473#_c_478_n 0.0031047f $X=3.035 $Y=2.51 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_431_n N_A_321_473#_c_478_n 0.0159397f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_283 N_VPWR_c_423_n N_A_321_473#_c_478_n 0.0111051f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_284 N_VGND_c_525_n A_385_47# 0.0056148f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_285 N_VGND_c_525_n A_477_47# 0.0105766f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_286 N_VGND_c_525_n A_565_47# 0.0028582f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
