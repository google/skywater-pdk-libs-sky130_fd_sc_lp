* File: sky130_fd_sc_lp__a21bo_2.pex.spice
* Created: Wed Sep  2 09:18:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BO_2%A_22_259# 1 2 7 9 12 14 16 18 21 23 26 29 30
+ 31 34 37 41 42 45 47 48 52
c91 47 0 9.79989e-20 $X=2.222 $Y=1.815
r92 51 52 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.49 $Y=1.46
+ $X2=0.565 $Y2=1.46
r93 43 45 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=2.715 $Y=0.86
+ $X2=2.715 $Y2=0.42
r94 41 43 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.585 $Y=0.945
+ $X2=2.715 $Y2=0.86
r95 41 42 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.585 $Y=0.945
+ $X2=2.36 $Y2=0.945
r96 39 42 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=2.272 $Y=1.03
+ $X2=2.36 $Y2=0.945
r97 39 47 49.7506 $w=1.73e-07 $l=7.85e-07 $layer=LI1_cond $X=2.272 $Y=1.03
+ $X2=2.272 $Y2=1.815
r98 35 48 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.222 $Y=2.495
+ $X2=2.222 $Y2=2.41
r99 35 37 17.3914 $w=2.73e-07 $l=4.15e-07 $layer=LI1_cond $X=2.222 $Y=2.495
+ $X2=2.222 $Y2=2.91
r100 32 48 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.222 $Y=2.325
+ $X2=2.222 $Y2=2.41
r101 32 34 14.4579 $w=2.73e-07 $l=3.45e-07 $layer=LI1_cond $X=2.222 $Y=2.325
+ $X2=2.222 $Y2=1.98
r102 31 47 7.25931 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.222 $Y=1.952
+ $X2=2.222 $Y2=1.815
r103 31 34 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=2.222 $Y=1.952
+ $X2=2.222 $Y2=1.98
r104 29 48 3.11956 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=2.085 $Y=2.41
+ $X2=2.222 $Y2=2.41
r105 29 30 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=2.085 $Y=2.41
+ $X2=0.44 $Y2=2.41
r106 27 51 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.275 $Y=1.46
+ $X2=0.49 $Y2=1.46
r107 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.46 $X2=0.275 $Y2=1.46
r108 24 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.275 $Y=2.325
+ $X2=0.44 $Y2=2.41
r109 24 26 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.275 $Y=2.325
+ $X2=0.275 $Y2=1.46
r110 19 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.92 $Y=1.445
+ $X2=0.92 $Y2=1.37
r111 19 21 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=0.92 $Y=1.445
+ $X2=0.92 $Y2=2.465
r112 16 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.92 $Y=1.295
+ $X2=0.92 $Y2=1.37
r113 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.92 $Y=1.295
+ $X2=0.92 $Y2=0.765
r114 14 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=1.37
+ $X2=0.92 $Y2=1.37
r115 14 52 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.845 $Y=1.37
+ $X2=0.565 $Y2=1.37
r116 10 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.625
+ $X2=0.49 $Y2=1.46
r117 10 12 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.49 $Y=1.625
+ $X2=0.49 $Y2=2.465
r118 7 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.295
+ $X2=0.49 $Y2=1.46
r119 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.49 $Y=1.295
+ $X2=0.49 $Y2=0.765
r120 2 37 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=1.835 $X2=2.25 $Y2=2.91
r121 2 34 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.125
+ $Y=1.835 $X2=2.25 $Y2=1.98
r122 1 45 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.54
+ $Y=0.235 $X2=2.68 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_2%B1_N 3 6 8 9 10 15 17
c28 15 0 1.16806e-19 $X=1.37 $Y=1.46
r29 15 18 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.372 $Y=1.46
+ $X2=1.372 $Y2=1.625
r30 15 17 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.372 $Y=1.46
+ $X2=1.372 $Y2=1.295
r31 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.46 $X2=1.37 $Y2=1.46
r32 9 10 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.257 $Y=1.665
+ $X2=1.257 $Y2=2.035
r33 9 16 5.98103 $w=3.93e-07 $l=2.05e-07 $layer=LI1_cond $X=1.257 $Y=1.665
+ $X2=1.257 $Y2=1.46
r34 8 16 4.814 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.257 $Y=1.295
+ $X2=1.257 $Y2=1.46
r35 6 18 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.465 $Y=2.045
+ $X2=1.465 $Y2=1.625
r36 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.445 $Y=0.975
+ $X2=1.445 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_2%A_304_153# 1 2 7 11 15 17 18 20 27
r44 26 27 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.915 $Y=1.46
+ $X2=1.915 $Y2=1.37
r45 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.46 $X2=1.915 $Y2=1.46
r46 23 25 16.4408 $w=3.97e-07 $l=5.35e-07 $layer=LI1_cond $X=1.755 $Y=0.925
+ $X2=1.755 $Y2=1.46
r47 18 25 6.52282 $w=3.97e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=1.625
+ $X2=1.755 $Y2=1.46
r48 18 20 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=1.755 $Y=1.625
+ $X2=1.755 $Y2=1.99
r49 13 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.465 $Y=1.445
+ $X2=2.465 $Y2=1.37
r50 13 15 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.465 $Y=1.445
+ $X2=2.465 $Y2=2.465
r51 9 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.465 $Y=1.295
+ $X2=2.465 $Y2=1.37
r52 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.465 $Y=1.295
+ $X2=2.465 $Y2=0.655
r53 8 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.08 $Y=1.37
+ $X2=1.915 $Y2=1.37
r54 7 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.39 $Y=1.37
+ $X2=2.465 $Y2=1.37
r55 7 8 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=2.39 $Y=1.37 $X2=2.08
+ $Y2=1.37
r56 2 20 600 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.835 $X2=1.72 $Y2=1.99
r57 1 23 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.765 $X2=1.66 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_2%A1 3 6 8 9 13 15
c34 13 0 9.79989e-20 $X=2.915 $Y=1.35
r35 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=1.515
r36 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=1.185
r37 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.35 $X2=2.915 $Y2=1.35
r38 9 14 7.50003 $w=3.13e-07 $l=2.05e-07 $layer=LI1_cond $X=3.12 $Y=1.357
+ $X2=2.915 $Y2=1.357
r39 8 14 10.061 $w=3.13e-07 $l=2.75e-07 $layer=LI1_cond $X=2.64 $Y=1.357
+ $X2=2.915 $Y2=1.357
r40 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.895 $Y=2.465
+ $X2=2.895 $Y2=1.515
r41 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.895 $Y=0.655
+ $X2=2.895 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_2%A2 3 6 8 11 13
r24 11 14 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.462 $Y=1.35
+ $X2=3.462 $Y2=1.515
r25 11 13 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.462 $Y=1.35
+ $X2=3.462 $Y2=1.185
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.47
+ $Y=1.35 $X2=3.47 $Y2=1.35
r27 8 12 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.6 $Y=1.35 $X2=3.47
+ $Y2=1.35
r28 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.365 $Y=2.465
+ $X2=3.365 $Y2=1.515
r29 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.365 $Y=0.655
+ $X2=3.365 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_2%VPWR 1 2 3 10 12 16 20 24 26 31 41 42 48 51
r48 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.13 $Y2=3.33
r54 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.6 $Y2=3.33
r55 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r59 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.135 $Y2=3.33
r61 32 34 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=1.68
+ $Y2=3.33
r62 31 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.13 $Y2=3.33
r63 31 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 30 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 27 45 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r68 27 29 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 26 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.135 $Y2=3.33
r70 26 29 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 24 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r72 24 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 20 23 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=3.13 $Y=2.11
+ $X2=3.13 $Y2=2.95
r74 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=3.33
r75 18 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=2.95
r76 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=3.33
r77 14 16 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=2.785
r78 10 45 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r79 10 12 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.785
r80 3 23 400 $w=1.7e-07 $l=1.19232e-06 $layer=licon1_PDIFF $count=1 $X=2.97
+ $Y=1.835 $X2=3.13 $Y2=2.95
r81 3 20 400 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.97
+ $Y=1.835 $X2=3.13 $Y2=2.11
r82 2 16 600 $w=1.7e-07 $l=1.0176e-06 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.785
r83 1 12 600 $w=1.7e-07 $l=1.01057e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_2%X 1 2 7 8 9 10 11
c16 7 0 1.16806e-19 $X=0.72 $Y=0.555
r17 10 11 16.8846 $w=2.13e-07 $l=3.15e-07 $layer=LI1_cond $X=0.717 $Y=1.665
+ $X2=0.717 $Y2=1.98
r18 9 10 19.8327 $w=2.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.717 $Y=1.295
+ $X2=0.717 $Y2=1.665
r19 8 9 19.8327 $w=2.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.717 $Y=0.925
+ $X2=0.717 $Y2=1.295
r20 7 8 23.3169 $w=2.13e-07 $l=4.35e-07 $layer=LI1_cond $X=0.717 $Y=0.49
+ $X2=0.717 $Y2=0.925
r21 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=1.98
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.345 $X2=0.705 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_2%A_508_367# 1 2 9 13 14 17
r23 17 19 38.2776 $w=2.78e-07 $l=9.3e-07 $layer=LI1_cond $X=3.605 $Y=1.98
+ $X2=3.605 $Y2=2.91
r24 15 17 5.14483 $w=2.78e-07 $l=1.25e-07 $layer=LI1_cond $X=3.605 $Y=1.855
+ $X2=3.605 $Y2=1.98
r25 13 15 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.465 $Y=1.77
+ $X2=3.605 $Y2=1.855
r26 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.465 $Y=1.77
+ $X2=2.795 $Y2=1.77
r27 9 11 40.4442 $w=2.63e-07 $l=9.3e-07 $layer=LI1_cond $X=2.662 $Y=1.98
+ $X2=2.662 $Y2=2.91
r28 7 14 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=2.662 $Y=1.855
+ $X2=2.795 $Y2=1.77
r29 7 9 5.43605 $w=2.63e-07 $l=1.25e-07 $layer=LI1_cond $X=2.662 $Y=1.855
+ $X2=2.662 $Y2=1.98
r30 2 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.835 $X2=3.58 $Y2=2.91
r31 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.835 $X2=3.58 $Y2=1.98
r32 1 11 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=1.835 $X2=2.68 $Y2=2.91
r33 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=1.835 $X2=2.68 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_2%VGND 1 2 3 4 13 15 19 23 27 29 31 33 35 40
+ 49 52 56
r59 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r60 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r61 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r62 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 44 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r64 44 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r65 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r66 41 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.25
+ $Y2=0
r67 41 43 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=3.12
+ $Y2=0
r68 40 55 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.627
+ $Y2=0
r69 40 43 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.12
+ $Y2=0
r70 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r71 39 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r72 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r73 36 46 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r74 36 38 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.72
+ $Y2=0
r75 35 49 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.147
+ $Y2=0
r76 35 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.72
+ $Y2=0
r77 33 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r78 33 50 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r79 29 55 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.627 $Y2=0
r80 29 31 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.58 $Y2=0.38
r81 25 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=0.085
+ $X2=2.25 $Y2=0
r82 25 27 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2.25 $Y=0.085
+ $X2=2.25 $Y2=0.54
r83 24 49 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.147
+ $Y2=0
r84 23 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.25
+ $Y2=0
r85 23 24 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=1.3
+ $Y2=0
r86 19 21 14.5472 $w=3.03e-07 $l=3.85e-07 $layer=LI1_cond $X=1.147 $Y=0.49
+ $X2=1.147 $Y2=0.875
r87 17 49 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.147 $Y=0.085
+ $X2=1.147 $Y2=0
r88 17 19 15.3029 $w=3.03e-07 $l=4.05e-07 $layer=LI1_cond $X=1.147 $Y=0.085
+ $X2=1.147 $Y2=0.49
r89 13 46 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r90 13 15 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.49
r91 4 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.44
+ $Y=0.235 $X2=3.58 $Y2=0.38
r92 3 27 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=2.125
+ $Y=0.235 $X2=2.25 $Y2=0.54
r93 2 21 182 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.345 $X2=1.135 $Y2=0.875
r94 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.345 $X2=1.135 $Y2=0.49
r95 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.345 $X2=0.275 $Y2=0.49
.ends

