* File: sky130_fd_sc_lp__and4bb_lp.spice
* Created: Wed Sep  2 09:34:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4bb_lp.pex.spice"
.subckt sky130_fd_sc_lp__and4bb_lp  VNB VPB A_N B_N C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1009 A_114_51# N_A_N_M1009_g N_A_27_51#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_N_M1002_g A_114_51# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1010 A_272_51# N_B_N_M1010_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1011 N_A_291_409#_M1011_d N_B_N_M1011_g A_272_51# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 A_548_47# N_A_27_51#_M1014_g N_A_461_47#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1006 A_626_47# N_A_291_409#_M1006_g A_548_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1007 A_704_47# N_C_M1007_g A_626_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_D_M1008_g A_704_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1016 A_896_47# N_A_461_47#_M1016_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0882 PD=0.63 PS=0.84 NRD=14.28 NRS=39.996 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_461_47#_M1000_g A_896_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_A_N_M1012_g N_A_27_51#_M1012_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_B_N_M1003_g N_A_291_409#_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1013 N_A_461_47#_M1013_d N_A_27_51#_M1013_g N_VPWR_M1003_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_A_291_409#_M1005_g N_A_461_47#_M1013_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.18 AS=0.14 PD=1.36 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1004 N_A_461_47#_M1004_d N_C_M1004_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.18 PD=1.28 PS=1.36 NRD=0 NRS=15.7403 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_D_M1001_g N_A_461_47#_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.1925 AS=0.14 PD=1.385 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1015 N_X_M1015_d N_A_461_47#_M1015_g N_VPWR_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.1925 PD=2.57 PS=1.385 NRD=0 NRS=20.685 M=1 R=4 SA=125003
+ SB=125000 A=0.25 P=2.5 MULT=1
DX17_noxref VNB VPB NWDIODE A=10.5559 P=15.05
c_67 VNB 0 1.66554e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__and4bb_lp.pxi.spice"
*
.ends
*
*
