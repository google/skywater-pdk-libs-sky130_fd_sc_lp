* File: sky130_fd_sc_lp__and4b_lp.pxi.spice
* Created: Wed Sep  2 09:33:47 2020
* 
x_PM_SKY130_FD_SC_LP__AND4B_LP%A_84_21# N_A_84_21#_M1010_d N_A_84_21#_M1013_d
+ N_A_84_21#_M1011_d N_A_84_21#_c_95_n N_A_84_21#_M1006_g N_A_84_21#_M1004_g
+ N_A_84_21#_c_96_n N_A_84_21#_c_97_n N_A_84_21#_M1012_g N_A_84_21#_c_98_n
+ N_A_84_21#_c_99_n N_A_84_21#_c_100_n N_A_84_21#_c_107_n N_A_84_21#_c_101_n
+ N_A_84_21#_c_102_n N_A_84_21#_c_109_n N_A_84_21#_c_110_n N_A_84_21#_c_111_n
+ N_A_84_21#_c_112_n N_A_84_21#_c_113_n N_A_84_21#_c_103_n N_A_84_21#_c_115_n
+ N_A_84_21#_c_116_n N_A_84_21#_c_104_n PM_SKY130_FD_SC_LP__AND4B_LP%A_84_21#
x_PM_SKY130_FD_SC_LP__AND4B_LP%D N_D_c_210_n N_D_M1013_g N_D_c_211_n N_D_M1000_g
+ N_D_c_212_n N_D_c_213_n N_D_c_214_n D D N_D_c_216_n
+ PM_SKY130_FD_SC_LP__AND4B_LP%D
x_PM_SKY130_FD_SC_LP__AND4B_LP%C N_C_M1009_g N_C_M1001_g N_C_c_264_n N_C_c_265_n
+ C C C C N_C_c_267_n PM_SKY130_FD_SC_LP__AND4B_LP%C
x_PM_SKY130_FD_SC_LP__AND4B_LP%B N_B_M1002_g N_B_c_314_n N_B_M1011_g N_B_c_315_n
+ N_B_c_316_n N_B_c_317_n N_B_c_318_n B B B B N_B_c_320_n
+ PM_SKY130_FD_SC_LP__AND4B_LP%B
x_PM_SKY130_FD_SC_LP__AND4B_LP%A_480_21# N_A_480_21#_M1003_d N_A_480_21#_M1005_d
+ N_A_480_21#_c_365_n N_A_480_21#_M1010_g N_A_480_21#_c_366_n
+ N_A_480_21#_c_367_n N_A_480_21#_c_368_n N_A_480_21#_M1007_g
+ N_A_480_21#_c_369_n N_A_480_21#_c_370_n N_A_480_21#_c_371_n
+ N_A_480_21#_c_378_n N_A_480_21#_c_372_n N_A_480_21#_c_373_n
+ PM_SKY130_FD_SC_LP__AND4B_LP%A_480_21#
x_PM_SKY130_FD_SC_LP__AND4B_LP%A_N N_A_N_M1008_g N_A_N_M1005_g N_A_N_M1003_g
+ N_A_N_c_438_n A_N N_A_N_c_439_n N_A_N_c_440_n PM_SKY130_FD_SC_LP__AND4B_LP%A_N
x_PM_SKY130_FD_SC_LP__AND4B_LP%X N_X_M1006_s N_X_M1004_s N_X_c_479_n N_X_c_477_n
+ X PM_SKY130_FD_SC_LP__AND4B_LP%X
x_PM_SKY130_FD_SC_LP__AND4B_LP%VPWR N_VPWR_M1004_d N_VPWR_M1009_d N_VPWR_M1007_d
+ N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n
+ VPWR N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_497_n N_VPWR_c_506_n
+ N_VPWR_c_507_n PM_SKY130_FD_SC_LP__AND4B_LP%VPWR
x_PM_SKY130_FD_SC_LP__AND4B_LP%VGND N_VGND_M1012_d N_VGND_M1008_s N_VGND_c_552_n
+ N_VGND_c_553_n N_VGND_c_554_n VGND N_VGND_c_555_n N_VGND_c_556_n
+ N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n PM_SKY130_FD_SC_LP__AND4B_LP%VGND
cc_1 VNB N_A_84_21#_c_95_n 0.0168575f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_2 VNB N_A_84_21#_c_96_n 0.0221815f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_3 VNB N_A_84_21#_c_97_n 0.0137388f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_4 VNB N_A_84_21#_c_98_n 0.0061567f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_5 VNB N_A_84_21#_c_99_n 0.0185761f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.165
cc_6 VNB N_A_84_21#_c_100_n 0.0245124f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.67
cc_7 VNB N_A_84_21#_c_101_n 0.00223075f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.33
cc_8 VNB N_A_84_21#_c_102_n 0.0148989f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.33
cc_9 VNB N_A_84_21#_c_103_n 0.0142817f $X=-0.19 $Y=-0.245 $X2=2.61 $Y2=1.97
cc_10 VNB N_A_84_21#_c_104_n 0.00350484f $X=-0.19 $Y=-0.245 $X2=2.69 $Y2=0.445
cc_11 VNB N_D_c_210_n 0.00185394f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=0.235
cc_12 VNB N_D_c_211_n 0.0142181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D_c_212_n 0.0154759f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_14 VNB N_D_c_213_n 0.0208877f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_15 VNB N_D_c_214_n 0.0154999f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.835
cc_16 VNB D 0.00616653f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.545
cc_17 VNB N_D_c_216_n 0.0156218f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_18 VNB N_C_M1001_g 0.0296622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_C_c_264_n 0.0230546f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_20 VNB N_C_c_265_n 0.00204627f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_21 VNB C 0.00783771f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_22 VNB N_C_c_267_n 0.0163348f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_23 VNB N_B_c_314_n 0.00219226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_c_315_n 0.0136386f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_25 VNB N_B_c_316_n 0.00953377f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_26 VNB N_B_c_317_n 0.013129f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_27 VNB N_B_c_318_n 0.0246995f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.165
cc_28 VNB B 0.00297804f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.835
cc_29 VNB N_B_c_320_n 0.017879f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_30 VNB N_A_480_21#_c_365_n 0.0176959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_480_21#_c_366_n 0.0357181f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_32 VNB N_A_480_21#_c_367_n 0.0125706f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_33 VNB N_A_480_21#_c_368_n 0.0161908f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_34 VNB N_A_480_21#_c_369_n 0.0499792f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.545
cc_35 VNB N_A_480_21#_c_370_n 0.00217589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_480_21#_c_371_n 0.0304066f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_37 VNB N_A_480_21#_c_372_n 0.0329251f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.33
cc_38 VNB N_A_480_21#_c_373_n 0.0209565f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.055
cc_39 VNB N_A_N_M1008_g 0.0224905f $X=-0.19 $Y=-0.245 $X2=2.33 $Y2=2.045
cc_40 VNB N_A_N_M1005_g 0.0332631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_N_M1003_g 0.0246614f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_42 VNB N_A_N_c_438_n 0.00295838f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.835
cc_43 VNB N_A_N_c_439_n 0.0374988f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_44 VNB N_A_N_c_440_n 0.00144844f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.97
cc_45 VNB N_X_c_477_n 0.0477299f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.88
cc_46 VNB X 0.0230781f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.165
cc_47 VNB N_VPWR_c_497_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.305 $Y2=2.055
cc_48 VNB N_VGND_c_552_n 0.00432289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_553_n 0.0506035f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_50 VNB N_VGND_c_554_n 0.00662781f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.835
cc_51 VNB N_VGND_c_555_n 0.0266231f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_52 VNB N_VGND_c_556_n 0.0268694f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.165
cc_53 VNB N_VGND_c_557_n 0.233029f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.67
cc_54 VNB N_VGND_c_558_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.33
cc_55 VNB N_VGND_c_559_n 0.00511011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VPB N_A_84_21#_M1004_g 0.032289f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.545
cc_57 VPB N_A_84_21#_c_100_n 0.00105918f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.67
cc_58 VPB N_A_84_21#_c_107_n 0.014908f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.835
cc_59 VPB N_A_84_21#_c_101_n 0.00274054f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.33
cc_60 VPB N_A_84_21#_c_109_n 0.00745329f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=2.055
cc_61 VPB N_A_84_21#_c_110_n 7.08592e-19 $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.055
cc_62 VPB N_A_84_21#_c_111_n 0.00207453f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=2.19
cc_63 VPB N_A_84_21#_c_112_n 0.00782233f $X=-0.19 $Y=1.655 $X2=2.305 $Y2=2.055
cc_64 VPB N_A_84_21#_c_113_n 0.00207453f $X=-0.19 $Y=1.655 $X2=2.47 $Y2=2.19
cc_65 VPB N_A_84_21#_c_103_n 0.00279657f $X=-0.19 $Y=1.655 $X2=2.61 $Y2=1.97
cc_66 VPB N_A_84_21#_c_115_n 0.0082777f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=2.055
cc_67 VPB N_A_84_21#_c_116_n 0.00669815f $X=-0.19 $Y=1.655 $X2=2.5 $Y2=2.055
cc_68 VPB N_D_c_210_n 0.0105975f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=0.235
cc_69 VPB N_D_M1013_g 0.0309416f $X=-0.19 $Y=1.655 $X2=2.33 $Y2=2.045
cc_70 VPB D 0.00183349f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.545
cc_71 VPB N_C_M1009_g 0.0313463f $X=-0.19 $Y=1.655 $X2=2.33 $Y2=2.045
cc_72 VPB N_C_c_265_n 0.0114346f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_73 VPB C 7.46359e-19 $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.88
cc_74 VPB N_B_c_314_n 0.0116871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_B_M1011_g 0.0313001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB B 5.07246e-19 $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.835
cc_77 VPB N_A_480_21#_c_368_n 0.0247463f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_78 VPB N_A_480_21#_M1007_g 0.0322058f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.165
cc_79 VPB N_A_480_21#_c_370_n 0.00833911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_480_21#_c_371_n 0.00181403f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_81 VPB N_A_480_21#_c_378_n 0.0556681f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.33
cc_82 VPB N_A_N_M1005_g 0.0515394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_X_c_479_n 0.0339041f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_84 VPB N_X_c_477_n 0.0285895f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.88
cc_85 VPB N_VPWR_c_498_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.165
cc_86 VPB N_VPWR_c_499_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_500_n 0.0105883f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_88 VPB N_VPWR_c_501_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.67
cc_89 VPB N_VPWR_c_502_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.835
cc_90 VPB N_VPWR_c_503_n 0.0207786f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.055
cc_91 VPB N_VPWR_c_504_n 0.034586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_497_n 0.0726148f $X=-0.19 $Y=1.655 $X2=2.305 $Y2=2.055
cc_93 VPB N_VPWR_c_506_n 0.024803f $X=-0.19 $Y=1.655 $X2=2.5 $Y2=2.19
cc_94 VPB N_VPWR_c_507_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.47 $Y2=2.9
cc_95 N_A_84_21#_c_107_n N_D_c_210_n 0.0126553f $X=0.585 $Y=1.835 $X2=-0.19
+ $Y2=-0.245
cc_96 N_A_84_21#_c_109_n N_D_c_210_n 2.68303e-19 $X=1.225 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_84_21#_c_115_n N_D_c_210_n 3.10581e-19 $X=1.39 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_84_21#_M1004_g N_D_M1013_g 0.0280273f $X=0.595 $Y=2.545 $X2=0 $Y2=0
cc_99 N_A_84_21#_c_107_n N_D_M1013_g 0.00246552f $X=0.585 $Y=1.835 $X2=0 $Y2=0
cc_100 N_A_84_21#_c_101_n N_D_M1013_g 0.00318388f $X=0.585 $Y=1.33 $X2=0 $Y2=0
cc_101 N_A_84_21#_c_109_n N_D_M1013_g 0.0178513f $X=1.225 $Y=2.055 $X2=0 $Y2=0
cc_102 N_A_84_21#_c_111_n N_D_M1013_g 0.0165176f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_103 N_A_84_21#_c_115_n N_D_M1013_g 0.00163378f $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_104 N_A_84_21#_c_97_n N_D_c_211_n 0.00978158f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_105 N_A_84_21#_c_99_n N_D_c_212_n 0.0063149f $X=0.585 $Y=1.165 $X2=0 $Y2=0
cc_106 N_A_84_21#_c_100_n N_D_c_213_n 0.0126553f $X=0.585 $Y=1.67 $X2=0 $Y2=0
cc_107 N_A_84_21#_c_96_n N_D_c_214_n 0.0108032f $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_108 N_A_84_21#_c_99_n D 2.57027e-19 $X=0.585 $Y=1.165 $X2=0 $Y2=0
cc_109 N_A_84_21#_c_101_n D 0.0395155f $X=0.585 $Y=1.33 $X2=0 $Y2=0
cc_110 N_A_84_21#_c_102_n D 0.00216912f $X=0.585 $Y=1.33 $X2=0 $Y2=0
cc_111 N_A_84_21#_c_109_n D 0.0192947f $X=1.225 $Y=2.055 $X2=0 $Y2=0
cc_112 N_A_84_21#_c_115_n D 0.0075854f $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_113 N_A_84_21#_c_99_n N_D_c_216_n 0.00151221f $X=0.585 $Y=1.165 $X2=0 $Y2=0
cc_114 N_A_84_21#_c_101_n N_D_c_216_n 0.00217048f $X=0.585 $Y=1.33 $X2=0 $Y2=0
cc_115 N_A_84_21#_c_102_n N_D_c_216_n 0.0126553f $X=0.585 $Y=1.33 $X2=0 $Y2=0
cc_116 N_A_84_21#_c_111_n N_C_M1009_g 0.0166112f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_117 N_A_84_21#_c_112_n N_C_M1009_g 0.0179678f $X=2.305 $Y=2.055 $X2=0 $Y2=0
cc_118 N_A_84_21#_c_113_n N_C_M1009_g 9.17538e-19 $X=2.47 $Y=2.19 $X2=0 $Y2=0
cc_119 N_A_84_21#_c_115_n N_C_M1009_g 0.00163378f $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_120 N_A_84_21#_c_112_n N_C_c_265_n 3.37098e-19 $X=2.305 $Y=2.055 $X2=0 $Y2=0
cc_121 N_A_84_21#_c_115_n N_C_c_265_n 2.25414e-19 $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_122 N_A_84_21#_c_112_n C 0.0200838f $X=2.305 $Y=2.055 $X2=0 $Y2=0
cc_123 N_A_84_21#_c_115_n C 0.00449587f $X=1.39 $Y=2.055 $X2=0 $Y2=0
cc_124 N_A_84_21#_c_112_n N_B_c_314_n 2.67978e-19 $X=2.305 $Y=2.055 $X2=0 $Y2=0
cc_125 N_A_84_21#_c_116_n N_B_c_314_n 0.0013432f $X=2.5 $Y=2.055 $X2=0 $Y2=0
cc_126 N_A_84_21#_c_111_n N_B_M1011_g 9.03227e-19 $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_127 N_A_84_21#_c_112_n N_B_M1011_g 0.018515f $X=2.305 $Y=2.055 $X2=0 $Y2=0
cc_128 N_A_84_21#_c_113_n N_B_M1011_g 0.0173065f $X=2.47 $Y=2.19 $X2=0 $Y2=0
cc_129 N_A_84_21#_c_103_n N_B_M1011_g 0.0036611f $X=2.61 $Y=1.97 $X2=0 $Y2=0
cc_130 N_A_84_21#_c_116_n N_B_M1011_g 0.00163378f $X=2.5 $Y=2.055 $X2=0 $Y2=0
cc_131 N_A_84_21#_c_104_n N_B_c_315_n 0.0010912f $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A_84_21#_c_103_n N_B_c_317_n 6.30807e-19 $X=2.61 $Y=1.97 $X2=0 $Y2=0
cc_133 N_A_84_21#_c_112_n B 0.0193186f $X=2.305 $Y=2.055 $X2=0 $Y2=0
cc_134 N_A_84_21#_c_116_n B 0.00321542f $X=2.5 $Y=2.055 $X2=0 $Y2=0
cc_135 N_A_84_21#_c_104_n B 0.089716f $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_136 N_A_84_21#_c_103_n N_B_c_320_n 0.00473665f $X=2.61 $Y=1.97 $X2=0 $Y2=0
cc_137 N_A_84_21#_c_103_n N_A_480_21#_c_365_n 0.00254758f $X=2.61 $Y=1.97 $X2=0
+ $Y2=0
cc_138 N_A_84_21#_c_104_n N_A_480_21#_c_365_n 0.00525439f $X=2.69 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A_84_21#_c_103_n N_A_480_21#_c_366_n 0.0115778f $X=2.61 $Y=1.97 $X2=0
+ $Y2=0
cc_140 N_A_84_21#_c_104_n N_A_480_21#_c_366_n 0.00756954f $X=2.69 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_84_21#_c_103_n N_A_480_21#_c_367_n 0.00214739f $X=2.61 $Y=1.97 $X2=0
+ $Y2=0
cc_142 N_A_84_21#_c_103_n N_A_480_21#_c_368_n 0.0085358f $X=2.61 $Y=1.97 $X2=0
+ $Y2=0
cc_143 N_A_84_21#_c_113_n N_A_480_21#_M1007_g 0.0170862f $X=2.47 $Y=2.19 $X2=0
+ $Y2=0
cc_144 N_A_84_21#_c_103_n N_A_480_21#_M1007_g 0.00771553f $X=2.61 $Y=1.97 $X2=0
+ $Y2=0
cc_145 N_A_84_21#_c_116_n N_A_480_21#_M1007_g 0.00582846f $X=2.5 $Y=2.055 $X2=0
+ $Y2=0
cc_146 N_A_84_21#_c_103_n N_A_480_21#_c_369_n 0.0127695f $X=2.61 $Y=1.97 $X2=0
+ $Y2=0
cc_147 N_A_84_21#_c_103_n N_A_480_21#_c_370_n 0.0250523f $X=2.61 $Y=1.97 $X2=0
+ $Y2=0
cc_148 N_A_84_21#_c_103_n N_A_N_M1008_g 0.00221821f $X=2.61 $Y=1.97 $X2=0 $Y2=0
cc_149 N_A_84_21#_c_104_n N_A_N_M1008_g 6.66399e-19 $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_84_21#_c_103_n N_A_N_c_440_n 0.0184874f $X=2.61 $Y=1.97 $X2=0 $Y2=0
cc_151 N_A_84_21#_M1004_g N_X_c_479_n 0.0140251f $X=0.595 $Y=2.545 $X2=0 $Y2=0
cc_152 N_A_84_21#_c_110_n N_X_c_479_n 0.00189912f $X=0.75 $Y=2.055 $X2=0 $Y2=0
cc_153 N_A_84_21#_c_95_n N_X_c_477_n 0.0329711f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_154 N_A_84_21#_M1004_g N_X_c_477_n 0.00767711f $X=0.595 $Y=2.545 $X2=0 $Y2=0
cc_155 N_A_84_21#_c_101_n N_X_c_477_n 0.0581196f $X=0.585 $Y=1.33 $X2=0 $Y2=0
cc_156 N_A_84_21#_c_110_n N_X_c_477_n 0.00935721f $X=0.75 $Y=2.055 $X2=0 $Y2=0
cc_157 N_A_84_21#_c_95_n X 0.00852454f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_158 N_A_84_21#_c_97_n X 0.00111159f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_159 N_A_84_21#_c_109_n N_VPWR_M1004_d 0.00180746f $X=1.225 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_84_21#_c_112_n N_VPWR_M1009_d 0.00202522f $X=2.305 $Y=2.055 $X2=0
+ $Y2=0
cc_161 N_A_84_21#_M1004_g N_VPWR_c_498_n 0.0186219f $X=0.595 $Y=2.545 $X2=0
+ $Y2=0
cc_162 N_A_84_21#_c_109_n N_VPWR_c_498_n 0.0146459f $X=1.225 $Y=2.055 $X2=0
+ $Y2=0
cc_163 N_A_84_21#_c_110_n N_VPWR_c_498_n 0.00189912f $X=0.75 $Y=2.055 $X2=0
+ $Y2=0
cc_164 N_A_84_21#_c_111_n N_VPWR_c_498_n 0.0490886f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_165 N_A_84_21#_c_111_n N_VPWR_c_499_n 0.0490886f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_166 N_A_84_21#_c_112_n N_VPWR_c_499_n 0.0164557f $X=2.305 $Y=2.055 $X2=0
+ $Y2=0
cc_167 N_A_84_21#_c_113_n N_VPWR_c_499_n 0.0460829f $X=2.47 $Y=2.19 $X2=0 $Y2=0
cc_168 N_A_84_21#_c_113_n N_VPWR_c_500_n 0.0347341f $X=2.47 $Y=2.19 $X2=0 $Y2=0
cc_169 N_A_84_21#_c_116_n N_VPWR_c_500_n 0.00538816f $X=2.5 $Y=2.055 $X2=0 $Y2=0
cc_170 N_A_84_21#_c_111_n N_VPWR_c_501_n 0.021949f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_171 N_A_84_21#_c_113_n N_VPWR_c_503_n 0.0257867f $X=2.47 $Y=2.19 $X2=0 $Y2=0
cc_172 N_A_84_21#_M1004_g N_VPWR_c_497_n 0.0141137f $X=0.595 $Y=2.545 $X2=0
+ $Y2=0
cc_173 N_A_84_21#_c_111_n N_VPWR_c_497_n 0.0124703f $X=1.39 $Y=2.19 $X2=0 $Y2=0
cc_174 N_A_84_21#_c_113_n N_VPWR_c_497_n 0.0145155f $X=2.47 $Y=2.19 $X2=0 $Y2=0
cc_175 N_A_84_21#_M1004_g N_VPWR_c_506_n 0.00769046f $X=0.595 $Y=2.545 $X2=0
+ $Y2=0
cc_176 N_A_84_21#_c_95_n N_VGND_c_552_n 0.00240189f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_177 N_A_84_21#_c_97_n N_VGND_c_552_n 0.0136342f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_178 N_A_84_21#_c_104_n N_VGND_c_553_n 0.0192986f $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_179 N_A_84_21#_c_104_n N_VGND_c_554_n 0.0246077f $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_180 N_A_84_21#_c_95_n N_VGND_c_555_n 0.00547815f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_181 N_A_84_21#_c_96_n N_VGND_c_555_n 4.87571e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_182 N_A_84_21#_c_97_n N_VGND_c_555_n 0.00486043f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_183 N_A_84_21#_M1010_d N_VGND_c_557_n 0.00232985f $X=2.55 $Y=0.235 $X2=0
+ $Y2=0
cc_184 N_A_84_21#_c_95_n N_VGND_c_557_n 0.010868f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_185 N_A_84_21#_c_96_n N_VGND_c_557_n 6.51792e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_186 N_A_84_21#_c_97_n N_VGND_c_557_n 0.00814425f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_187 N_A_84_21#_c_104_n N_VGND_c_557_n 0.0124718f $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_188 N_D_M1013_g N_C_M1009_g 0.0196369f $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_189 N_D_c_211_n N_C_M1001_g 0.0407119f $X=1.305 $Y=0.73 $X2=0 $Y2=0
cc_190 N_D_c_212_n N_C_M1001_g 0.0078056f $X=1.125 $Y=1.12 $X2=0 $Y2=0
cc_191 N_D_c_213_n N_C_c_264_n 0.0139518f $X=1.125 $Y=1.625 $X2=0 $Y2=0
cc_192 N_D_c_210_n N_C_c_265_n 0.0139518f $X=1.125 $Y=1.79 $X2=0 $Y2=0
cc_193 N_D_c_211_n C 0.00682848f $X=1.305 $Y=0.73 $X2=0 $Y2=0
cc_194 N_D_c_212_n C 0.00549467f $X=1.125 $Y=1.12 $X2=0 $Y2=0
cc_195 D C 0.0499848f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_196 N_D_c_216_n C 7.98982e-19 $X=1.125 $Y=1.285 $X2=0 $Y2=0
cc_197 D N_C_c_267_n 0.00382414f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_198 N_D_c_216_n N_C_c_267_n 0.0139518f $X=1.125 $Y=1.285 $X2=0 $Y2=0
cc_199 N_D_M1013_g N_X_c_479_n 2.04297e-19 $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_200 N_D_M1013_g N_VPWR_c_498_n 0.0175722f $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_201 N_D_M1013_g N_VPWR_c_499_n 8.63241e-19 $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_202 N_D_M1013_g N_VPWR_c_501_n 0.00769046f $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_203 N_D_M1013_g N_VPWR_c_497_n 0.0134474f $X=1.125 $Y=2.545 $X2=0 $Y2=0
cc_204 N_D_c_211_n N_VGND_c_552_n 0.0107229f $X=1.305 $Y=0.73 $X2=0 $Y2=0
cc_205 N_D_c_214_n N_VGND_c_552_n 0.00327338f $X=1.305 $Y=0.805 $X2=0 $Y2=0
cc_206 D N_VGND_c_552_n 0.0117644f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_207 N_D_c_216_n N_VGND_c_552_n 0.00122441f $X=1.125 $Y=1.285 $X2=0 $Y2=0
cc_208 N_D_c_211_n N_VGND_c_553_n 0.00564095f $X=1.305 $Y=0.73 $X2=0 $Y2=0
cc_209 N_D_c_211_n N_VGND_c_557_n 0.00950947f $X=1.305 $Y=0.73 $X2=0 $Y2=0
cc_210 N_C_c_265_n N_B_c_314_n 0.0135694f $X=1.665 $Y=1.79 $X2=0 $Y2=0
cc_211 N_C_M1009_g N_B_M1011_g 0.0290426f $X=1.655 $Y=2.545 $X2=0 $Y2=0
cc_212 N_C_M1001_g N_B_c_315_n 0.0416847f $X=1.695 $Y=0.445 $X2=0 $Y2=0
cc_213 C N_B_c_315_n 0.00260749f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_214 N_C_M1001_g N_B_c_317_n 0.0102342f $X=1.695 $Y=0.445 $X2=0 $Y2=0
cc_215 C N_B_c_317_n 0.00140033f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_216 N_C_c_264_n N_B_c_318_n 0.0135694f $X=1.665 $Y=1.625 $X2=0 $Y2=0
cc_217 N_C_M1001_g B 7.6356e-19 $X=1.695 $Y=0.445 $X2=0 $Y2=0
cc_218 C B 0.0873337f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_219 N_C_c_267_n B 0.00232743f $X=1.665 $Y=1.285 $X2=0 $Y2=0
cc_220 C N_B_c_320_n 0.00232658f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_221 N_C_c_267_n N_B_c_320_n 0.0135694f $X=1.665 $Y=1.285 $X2=0 $Y2=0
cc_222 N_C_M1009_g N_VPWR_c_498_n 8.63241e-19 $X=1.655 $Y=2.545 $X2=0 $Y2=0
cc_223 N_C_M1009_g N_VPWR_c_499_n 0.017679f $X=1.655 $Y=2.545 $X2=0 $Y2=0
cc_224 N_C_M1009_g N_VPWR_c_501_n 0.00769046f $X=1.655 $Y=2.545 $X2=0 $Y2=0
cc_225 N_C_M1009_g N_VPWR_c_497_n 0.0134474f $X=1.655 $Y=2.545 $X2=0 $Y2=0
cc_226 N_C_M1001_g N_VGND_c_552_n 0.00222745f $X=1.695 $Y=0.445 $X2=0 $Y2=0
cc_227 C N_VGND_c_552_n 0.0130116f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_228 N_C_M1001_g N_VGND_c_553_n 0.00393362f $X=1.695 $Y=0.445 $X2=0 $Y2=0
cc_229 C N_VGND_c_553_n 0.00843335f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_230 N_C_M1001_g N_VGND_c_557_n 0.00544199f $X=1.695 $Y=0.445 $X2=0 $Y2=0
cc_231 C N_VGND_c_557_n 0.0106746f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_232 C A_276_47# 0.00302196f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_233 C A_354_47# 0.00200068f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_234 N_B_c_315_n N_A_480_21#_c_365_n 0.0330224f $X=2.1 $Y=0.73 $X2=0 $Y2=0
cc_235 B N_A_480_21#_c_365_n 0.00250837f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_236 N_B_c_316_n N_A_480_21#_c_367_n 0.00978005f $X=2.1 $Y=0.88 $X2=0 $Y2=0
cc_237 N_B_c_314_n N_A_480_21#_c_368_n 0.00498561f $X=2.205 $Y=1.79 $X2=0 $Y2=0
cc_238 N_B_M1011_g N_A_480_21#_c_368_n 0.0174109f $X=2.205 $Y=2.545 $X2=0 $Y2=0
cc_239 N_B_c_318_n N_A_480_21#_c_368_n 0.00884207f $X=2.205 $Y=1.625 $X2=0 $Y2=0
cc_240 N_B_c_317_n N_A_480_21#_c_369_n 0.00403073f $X=2.205 $Y=1.12 $X2=0 $Y2=0
cc_241 N_B_c_320_n N_A_480_21#_c_369_n 0.00884207f $X=2.205 $Y=1.285 $X2=0 $Y2=0
cc_242 N_B_M1011_g N_VPWR_c_499_n 0.0158808f $X=2.205 $Y=2.545 $X2=0 $Y2=0
cc_243 N_B_M1011_g N_VPWR_c_503_n 0.00840515f $X=2.205 $Y=2.545 $X2=0 $Y2=0
cc_244 N_B_M1011_g N_VPWR_c_497_n 0.0146909f $X=2.205 $Y=2.545 $X2=0 $Y2=0
cc_245 N_B_c_315_n N_VGND_c_553_n 0.00433047f $X=2.1 $Y=0.73 $X2=0 $Y2=0
cc_246 B N_VGND_c_553_n 0.00854282f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_247 N_B_c_315_n N_VGND_c_557_n 0.00655311f $X=2.1 $Y=0.73 $X2=0 $Y2=0
cc_248 B N_VGND_c_557_n 0.00996452f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_249 B A_432_47# 0.00176828f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_250 N_A_480_21#_c_366_n N_A_N_M1008_g 0.0149926f $X=2.71 $Y=0.805 $X2=0 $Y2=0
cc_251 N_A_480_21#_c_373_n N_A_N_M1008_g 0.00121917f $X=4.04 $Y=0.47 $X2=0 $Y2=0
cc_252 N_A_480_21#_c_368_n N_A_N_M1005_g 0.0192612f $X=2.735 $Y=1.82 $X2=0 $Y2=0
cc_253 N_A_480_21#_c_369_n N_A_N_M1005_g 0.0300488f $X=2.945 $Y=1.46 $X2=0 $Y2=0
cc_254 N_A_480_21#_c_370_n N_A_N_M1005_g 0.0242314f $X=3.645 $Y=1.53 $X2=0 $Y2=0
cc_255 N_A_480_21#_c_371_n N_A_N_M1005_g 0.00826078f $X=3.81 $Y=1.695 $X2=0
+ $Y2=0
cc_256 N_A_480_21#_c_378_n N_A_N_M1005_g 0.0427348f $X=3.81 $Y=2.19 $X2=0 $Y2=0
cc_257 N_A_480_21#_c_372_n N_A_N_M1005_g 0.0038234f $X=4.12 $Y=1.365 $X2=0 $Y2=0
cc_258 N_A_480_21#_c_372_n N_A_N_M1003_g 0.0131282f $X=4.12 $Y=1.365 $X2=0 $Y2=0
cc_259 N_A_480_21#_c_373_n N_A_N_M1003_g 0.00850185f $X=4.04 $Y=0.47 $X2=0 $Y2=0
cc_260 N_A_480_21#_c_371_n N_A_N_c_438_n 0.0164462f $X=3.81 $Y=1.695 $X2=0 $Y2=0
cc_261 N_A_480_21#_c_372_n N_A_N_c_438_n 0.0245788f $X=4.12 $Y=1.365 $X2=0 $Y2=0
cc_262 N_A_480_21#_c_369_n N_A_N_c_439_n 0.0149926f $X=2.945 $Y=1.46 $X2=0 $Y2=0
cc_263 N_A_480_21#_c_370_n N_A_N_c_439_n 7.9644e-19 $X=3.645 $Y=1.53 $X2=0 $Y2=0
cc_264 N_A_480_21#_c_371_n N_A_N_c_439_n 0.00726817f $X=3.81 $Y=1.695 $X2=0
+ $Y2=0
cc_265 N_A_480_21#_c_366_n N_A_N_c_440_n 0.0053175f $X=2.71 $Y=0.805 $X2=0 $Y2=0
cc_266 N_A_480_21#_c_369_n N_A_N_c_440_n 0.0149968f $X=2.945 $Y=1.46 $X2=0 $Y2=0
cc_267 N_A_480_21#_c_370_n N_A_N_c_440_n 0.0478347f $X=3.645 $Y=1.53 $X2=0 $Y2=0
cc_268 N_A_480_21#_M1007_g N_VPWR_c_499_n 8.46437e-19 $X=2.735 $Y=2.545 $X2=0
+ $Y2=0
cc_269 N_A_480_21#_c_368_n N_VPWR_c_500_n 0.00745268f $X=2.735 $Y=1.82 $X2=0
+ $Y2=0
cc_270 N_A_480_21#_M1007_g N_VPWR_c_500_n 0.003604f $X=2.735 $Y=2.545 $X2=0
+ $Y2=0
cc_271 N_A_480_21#_c_370_n N_VPWR_c_500_n 0.0169963f $X=3.645 $Y=1.53 $X2=0
+ $Y2=0
cc_272 N_A_480_21#_c_378_n N_VPWR_c_500_n 0.0387929f $X=3.81 $Y=2.19 $X2=0 $Y2=0
cc_273 N_A_480_21#_M1007_g N_VPWR_c_503_n 0.0077662f $X=2.735 $Y=2.545 $X2=0
+ $Y2=0
cc_274 N_A_480_21#_c_378_n N_VPWR_c_504_n 0.0220321f $X=3.81 $Y=2.19 $X2=0 $Y2=0
cc_275 N_A_480_21#_M1007_g N_VPWR_c_497_n 0.0137168f $X=2.735 $Y=2.545 $X2=0
+ $Y2=0
cc_276 N_A_480_21#_c_378_n N_VPWR_c_497_n 0.0125808f $X=3.81 $Y=2.19 $X2=0 $Y2=0
cc_277 N_A_480_21#_c_365_n N_VGND_c_553_n 0.00549284f $X=2.475 $Y=0.73 $X2=0
+ $Y2=0
cc_278 N_A_480_21#_c_366_n N_VGND_c_553_n 0.00521502f $X=2.71 $Y=0.805 $X2=0
+ $Y2=0
cc_279 N_A_480_21#_c_365_n N_VGND_c_554_n 0.002414f $X=2.475 $Y=0.73 $X2=0 $Y2=0
cc_280 N_A_480_21#_c_366_n N_VGND_c_554_n 0.0028014f $X=2.71 $Y=0.805 $X2=0
+ $Y2=0
cc_281 N_A_480_21#_c_373_n N_VGND_c_554_n 0.0122119f $X=4.04 $Y=0.47 $X2=0 $Y2=0
cc_282 N_A_480_21#_c_373_n N_VGND_c_556_n 0.0195507f $X=4.04 $Y=0.47 $X2=0 $Y2=0
cc_283 N_A_480_21#_M1003_d N_VGND_c_557_n 0.00232985f $X=3.9 $Y=0.235 $X2=0
+ $Y2=0
cc_284 N_A_480_21#_c_365_n N_VGND_c_557_n 0.0114101f $X=2.475 $Y=0.73 $X2=0
+ $Y2=0
cc_285 N_A_480_21#_c_366_n N_VGND_c_557_n 0.00633619f $X=2.71 $Y=0.805 $X2=0
+ $Y2=0
cc_286 N_A_480_21#_c_373_n N_VGND_c_557_n 0.0124998f $X=4.04 $Y=0.47 $X2=0 $Y2=0
cc_287 N_A_N_M1005_g N_VPWR_c_500_n 0.0142936f $X=3.545 $Y=2.545 $X2=0 $Y2=0
cc_288 N_A_N_M1005_g N_VPWR_c_504_n 0.0086001f $X=3.545 $Y=2.545 $X2=0 $Y2=0
cc_289 N_A_N_M1005_g N_VPWR_c_497_n 0.0169093f $X=3.545 $Y=2.545 $X2=0 $Y2=0
cc_290 N_A_N_M1008_g N_VGND_c_554_n 0.0129216f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_291 N_A_N_M1003_g N_VGND_c_554_n 0.00227546f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_292 N_A_N_c_438_n N_VGND_c_554_n 0.00983511f $X=3.685 $Y=1.02 $X2=0 $Y2=0
cc_293 N_A_N_c_440_n N_VGND_c_554_n 0.0118246f $X=3.235 $Y=0.997 $X2=0 $Y2=0
cc_294 N_A_N_M1008_g N_VGND_c_556_n 0.00486043f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_295 N_A_N_M1003_g N_VGND_c_556_n 0.00549284f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_296 N_A_N_M1008_g N_VGND_c_557_n 0.00443987f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_297 N_A_N_M1003_g N_VGND_c_557_n 0.00796501f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_298 N_A_N_c_438_n N_VGND_c_557_n 0.0140331f $X=3.685 $Y=1.02 $X2=0 $Y2=0
cc_299 N_A_N_c_439_n N_VGND_c_557_n 7.60946e-19 $X=3.825 $Y=1.02 $X2=0 $Y2=0
cc_300 N_A_N_c_440_n N_VGND_c_557_n 0.00330605f $X=3.235 $Y=0.997 $X2=0 $Y2=0
cc_301 N_X_c_479_n N_VPWR_c_498_n 0.0498359f $X=0.33 $Y=2.485 $X2=0 $Y2=0
cc_302 N_X_c_479_n N_VPWR_c_497_n 0.0154828f $X=0.33 $Y=2.485 $X2=0 $Y2=0
cc_303 N_X_c_479_n N_VPWR_c_506_n 0.0270889f $X=0.33 $Y=2.485 $X2=0 $Y2=0
cc_304 X N_VGND_c_552_n 0.0137589f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_305 X N_VGND_c_555_n 0.0207696f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_306 N_X_M1006_s N_VGND_c_557_n 0.00233022f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_307 X N_VGND_c_557_n 0.0134309f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_308 A_114_47# N_VGND_c_557_n 0.00829524f $X=0.57 $Y=0.235 $X2=4.08 $Y2=0
cc_309 N_VGND_c_557_n A_276_47# 0.00626835f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_310 N_VGND_c_557_n A_354_47# 0.00829053f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_311 N_VGND_c_557_n A_432_47# 0.00407766f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_312 N_VGND_c_557_n A_708_47# 0.00312872f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
