* File: sky130_fd_sc_lp__einvn_lp.spice
* Created: Fri Aug 28 10:33:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvn_lp.pex.spice"
.subckt sky130_fd_sc_lp__einvn_lp  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1003 A_115_148# N_TE_B_M1003_g N_A_28_148#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_TE_B_M1001_g A_115_148# VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.0441 PD=0.755 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1000 A_284_148# N_A_28_148#_M1000_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.07035 PD=0.745 PS=0.755 NRD=30.708 NRS=15.708 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_Z_M1005_d N_A_M1005_g A_284_148# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.06825 PD=1.41 PS=0.745 NRD=0 NRS=30.708 M=1 R=2.8 SA=75001.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_TE_B_M1004_g N_A_28_148#_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1002 A_252_414# N_TE_B_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.14 PD=1.24 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_Z_M1006_d N_A_M1006_g A_252_414# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.12 PD=2.57 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125000 A=0.25
+ P=2.5 MULT=1
DX7_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__einvn_lp.pxi.spice"
*
.ends
*
*
