* NGSPICE file created from sky130_fd_sc_lp__o221a_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o221a_0 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 a_127_106# B2 a_213_106# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.352e+11p ps=2.8e+06u
M1001 a_213_106# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1002 a_32_484# B2 a_269_484# VPB phighvt w=640000u l=150000u
+  ad=4.192e+11p pd=3.87e+06u as=1.344e+11p ps=1.7e+06u
M1003 a_269_484# B1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=7.936e+11p ps=5.04e+06u
M1004 VPWR A1 a_449_484# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1005 VPWR C1 a_32_484# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_32_484# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1007 a_213_106# B1 a_127_106# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_127_106# C1 a_32_484# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 VGND A1 a_213_106# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_32_484# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 a_449_484# A2 a_32_484# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

