* File: sky130_fd_sc_lp__inv_0.spice
* Created: Fri Aug 28 10:37:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__inv_0.pex.spice"
.subckt sky130_fd_sc_lp__inv_0  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.2 A=0.063
+ P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX2_noxref VNB VPB NWDIODE A=2.4991 P=6.41
*
.include "sky130_fd_sc_lp__inv_0.pxi.spice"
*
.ends
*
*
