* File: sky130_fd_sc_lp__a22oi_2.pex.spice
* Created: Fri Aug 28 09:54:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22OI_2%A1 3 7 11 15 17 18 19 20 32 33 37 38 40
c87 15 0 1.73976e-19 $X=2.54 $Y=2.465
r88 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.29
+ $Y=1.51 $X2=2.29 $Y2=1.51
r89 35 37 3.51825 $w=2.74e-07 $l=2e-08 $layer=POLY_cond $X=2.27 $Y=1.51 $X2=2.29
+ $Y2=1.51
r90 31 33 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=0.72 $Y=1.51 $X2=0.82
+ $Y2=1.51
r91 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.51 $X2=0.72 $Y2=1.51
r92 28 31 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.585 $Y=1.51
+ $X2=0.72 $Y2=1.51
r93 20 40 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.25 $Y=2.035
+ $X2=2.125 $Y2=2.035
r94 20 38 14.9227 $w=3.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.25 $Y=1.95
+ $X2=2.25 $Y2=1.51
r95 20 40 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.1 $Y=2.035
+ $X2=2.125 $Y2=2.035
r96 19 20 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=2.1 $Y2=2.035
r97 18 19 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=1.68 $Y2=2.035
r98 18 41 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=0.885 $Y2=2.035
r99 17 41 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.755 $Y=2.035
+ $X2=0.885 $Y2=2.035
r100 17 32 13.5803 $w=4.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.755 $Y=1.95
+ $X2=0.755 $Y2=1.51
r101 13 37 43.9781 $w=2.74e-07 $l=3.22102e-07 $layer=POLY_cond $X=2.54 $Y=1.675
+ $X2=2.29 $Y2=1.51
r102 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.54 $Y=1.675
+ $X2=2.54 $Y2=2.465
r103 9 35 16.847 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.345
+ $X2=2.27 $Y2=1.51
r104 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.27 $Y=1.345
+ $X2=2.27 $Y2=0.655
r105 5 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.82 $Y=1.345
+ $X2=0.82 $Y2=1.51
r106 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.82 $Y=1.345
+ $X2=0.82 $Y2=0.655
r107 1 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.675
+ $X2=0.585 $Y2=1.51
r108 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.585 $Y=1.675
+ $X2=0.585 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_2%A2 3 7 9 13 17 19 20 21 24 28
r61 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.51
+ $X2=1.75 $Y2=1.675
r62 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.51 $X2=1.75 $Y2=1.51
r63 24 27 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.75 $Y=1.42 $X2=1.75
+ $Y2=1.51
r64 24 25 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=1.42 $X2=1.75
+ $Y2=1.345
r65 21 28 1.85451 $w=4.33e-07 $l=7e-08 $layer=LI1_cond $X=1.68 $Y=1.562 $X2=1.75
+ $Y2=1.562
r66 20 21 12.7166 $w=4.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.562
+ $X2=1.68 $Y2=1.562
r67 17 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.84 $Y=0.655
+ $X2=1.84 $Y2=1.345
r68 13 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.66 $Y=2.465
+ $X2=1.66 $Y2=1.675
r69 10 19 5.30422 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.325 $Y=1.42
+ $X2=1.24 $Y2=1.42
r70 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.42
+ $X2=1.75 $Y2=1.42
r71 9 10 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.585 $Y=1.42
+ $X2=1.325 $Y2=1.42
r72 5 19 20.4101 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=1.25 $Y=1.345
+ $X2=1.24 $Y2=1.42
r73 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.25 $Y=1.345 $X2=1.25
+ $Y2=0.655
r74 1 19 20.4101 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=1.23 $Y=1.495
+ $X2=1.24 $Y2=1.42
r75 1 3 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=1.23 $Y=1.495 $X2=1.23
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_2%B1 3 7 11 15 19 20 22 23 24 25 32 33
c75 23 0 1.73976e-19 $X=3.155 $Y=2.01
c76 22 0 2.25787e-20 $X=3.985 $Y=2.01
c77 7 0 8.0434e-20 $X=2.97 $Y=2.465
r78 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.39 $Y=1.51
+ $X2=4.39 $Y2=1.675
r79 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.39 $Y=1.51
+ $X2=4.39 $Y2=1.345
r80 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.39
+ $Y=1.51 $X2=4.39 $Y2=1.51
r81 25 33 8.82117 $w=4.03e-07 $l=3.1e-07 $layer=LI1_cond $X=4.08 $Y=1.547
+ $X2=4.39 $Y2=1.547
r82 25 38 0.142277 $w=4.03e-07 $l=5e-09 $layer=LI1_cond $X=4.08 $Y=1.547
+ $X2=4.075 $Y2=1.547
r83 25 38 5.50734 $w=1.8e-07 $l=2.03e-07 $layer=LI1_cond $X=4.075 $Y=1.75
+ $X2=4.075 $Y2=1.547
r84 24 25 7.15827 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=4.075 $Y=1.925
+ $X2=4.075 $Y2=1.75
r85 22 24 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.985 $Y=2.01
+ $X2=4.075 $Y2=1.925
r86 22 23 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.985 $Y=2.01
+ $X2=3.155 $Y2=2.01
r87 20 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.51
+ $X2=2.99 $Y2=1.675
r88 20 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.99 $Y=1.51
+ $X2=2.99 $Y2=1.345
r89 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.51 $X2=2.99 $Y2=1.51
r90 17 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.03 $Y=1.925
+ $X2=3.155 $Y2=2.01
r91 17 19 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=3.03 $Y=1.925
+ $X2=3.03 $Y2=1.51
r92 15 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.3 $Y=2.465 $X2=4.3
+ $Y2=1.675
r93 11 34 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.3 $Y=0.655 $X2=4.3
+ $Y2=1.345
r94 7 30 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.97 $Y=2.465
+ $X2=2.97 $Y2=1.675
r95 3 29 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.9 $Y=0.655 $X2=2.9
+ $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_2%B2 3 7 11 15 17 23 24
c50 23 0 8.0434e-20 $X=3.73 $Y=1.51
r51 22 24 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.73 $Y=1.51
+ $X2=3.87 $Y2=1.51
r52 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.51 $X2=3.73 $Y2=1.51
r53 19 22 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=3.44 $Y=1.51
+ $X2=3.73 $Y2=1.51
r54 17 23 4.11983 $w=4.48e-07 $l=1.55e-07 $layer=LI1_cond $X=3.59 $Y=1.665
+ $X2=3.59 $Y2=1.51
r55 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.87 $Y=1.675
+ $X2=3.87 $Y2=1.51
r56 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.87 $Y=1.675
+ $X2=3.87 $Y2=2.465
r57 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.87 $Y=1.345
+ $X2=3.87 $Y2=1.51
r58 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.87 $Y=1.345
+ $X2=3.87 $Y2=0.655
r59 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=1.675
+ $X2=3.44 $Y2=1.51
r60 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.44 $Y=1.675 $X2=3.44
+ $Y2=2.465
r61 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=1.345
+ $X2=3.44 $Y2=1.51
r62 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.44 $Y=1.345 $X2=3.44
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_2%A_49_367# 1 2 3 4 5 18 22 26 28 31 33 34 35
+ 36 38 40 43 45 48 51
c73 36 0 2.25787e-20 $X=4.41 $Y=2.92
r74 50 51 3.16842 $w=4.68e-07 $l=7e-08 $layer=LI1_cond $X=3.655 $Y=2.84
+ $X2=3.725 $Y2=2.84
r75 47 48 9.33757 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=2.84
+ $X2=2.59 $Y2=2.84
r76 38 53 3.66588 $w=2.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.545 $Y=2.765
+ $X2=4.545 $Y2=2.92
r77 38 40 26.0367 $w=2.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.545 $Y=2.765
+ $X2=4.545 $Y2=2.155
r78 36 53 3.19286 $w=3.1e-07 $l=1.35e-07 $layer=LI1_cond $X=4.41 $Y=2.92
+ $X2=4.545 $Y2=2.92
r79 36 51 25.4653 $w=3.08e-07 $l=6.85e-07 $layer=LI1_cond $X=4.41 $Y=2.92
+ $X2=3.725 $Y2=2.92
r80 35 47 7.76179 $w=4.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.06 $Y=2.84
+ $X2=2.755 $Y2=2.84
r81 34 50 4.199 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.49 $Y=2.84
+ $X2=3.655 $Y2=2.84
r82 34 35 10.9428 $w=4.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.49 $Y=2.84
+ $X2=3.06 $Y2=2.84
r83 33 48 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.38 $Y=2.69
+ $X2=2.59 $Y2=2.69
r84 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=2.605
+ $X2=2.38 $Y2=2.69
r85 30 31 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.295 $Y=2.46
+ $X2=2.295 $Y2=2.605
r86 29 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.54 $Y=2.375
+ $X2=1.41 $Y2=2.375
r87 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.21 $Y=2.375
+ $X2=2.295 $Y2=2.46
r88 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.21 $Y=2.375
+ $X2=1.54 $Y2=2.375
r89 24 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=2.46
+ $X2=1.41 $Y2=2.375
r90 24 26 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=1.41 $Y=2.46
+ $X2=1.41 $Y2=2.91
r91 23 43 3.3199 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=2.375
+ $X2=0.37 $Y2=2.375
r92 22 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.28 $Y=2.375
+ $X2=1.41 $Y2=2.375
r93 22 23 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.28 $Y=2.375
+ $X2=0.535 $Y2=2.375
r94 16 43 3.24686 $w=2.9e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.33 $Y=2.29
+ $X2=0.37 $Y2=2.375
r95 16 18 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=0.33 $Y=2.29
+ $X2=0.33 $Y2=2.02
r96 5 53 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.375
+ $Y=1.835 $X2=4.515 $Y2=2.91
r97 5 40 300 $w=1.7e-07 $l=3.83667e-07 $layer=licon1_PDIFF $count=2 $X=4.375
+ $Y=1.835 $X2=4.515 $Y2=2.155
r98 4 50 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.835 $X2=3.655 $Y2=2.895
r99 3 47 600 $w=1.7e-07 $l=1.00256e-06 $layer=licon1_PDIFF $count=1 $X=2.615
+ $Y=1.835 $X2=2.755 $Y2=2.77
r100 2 45 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=1.305
+ $Y=1.835 $X2=1.445 $Y2=2.375
r101 2 26 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.305
+ $Y=1.835 $X2=1.445 $Y2=2.91
r102 1 43 300 $w=1.7e-07 $l=6.79632e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.455
r103 1 18 600 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_2%VPWR 1 2 9 12 13 14 20 29 30 37
r65 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 35 37 5.86751 $w=5.51e-07 $l=2.65e-07 $layer=LI1_cond $X=2.06 $Y=3.065
+ $X2=2.06 $Y2=3.33
r67 33 35 6.86388 $w=5.51e-07 $l=3.91727e-07 $layer=LI1_cond $X=1.875 $Y=2.755
+ $X2=2.06 $Y2=3.065
r68 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r69 27 30 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r70 26 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r71 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r72 24 37 7.77084 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=2.41 $Y=3.33 $X2=2.06
+ $Y2=3.33
r73 24 26 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.64 $Y2=3.33
r74 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 20 37 7.77084 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=1.71 $Y=3.33 $X2=2.06
+ $Y2=3.33
r77 20 22 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.71 $Y=3.33 $X2=1.68
+ $Y2=3.33
r78 18 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 14 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 14 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 12 17 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.75 $Y=3.33 $X2=0.72
+ $Y2=3.33
r83 12 13 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=3.33
+ $X2=0.915 $Y2=3.33
r84 11 22 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.08 $Y=3.33 $X2=1.68
+ $Y2=3.33
r85 11 13 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=3.33
+ $X2=0.915 $Y2=3.33
r86 7 13 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.915 $Y=3.245
+ $X2=0.915 $Y2=3.33
r87 7 9 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.915 $Y=3.245
+ $X2=0.915 $Y2=2.755
r88 2 35 600 $w=1.7e-07 $l=1.46294e-06 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=1.835 $X2=2.245 $Y2=3.065
r89 2 33 600 $w=1.7e-07 $l=9.87522e-07 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=1.835 $X2=1.875 $Y2=2.755
r90 1 9 600 $w=1.7e-07 $l=1.03971e-06 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.915 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_2%Y 1 2 3 4 5 18 20 21 24 26 27 30 34 37 39 44
+ 45
r97 44 45 22.1818 $w=1.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.642 $Y=1.665
+ $X2=2.642 $Y2=2.035
r98 39 42 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=4.08 $Y=2.35 $X2=4.08
+ $Y2=2.43
r99 38 45 13.7887 $w=1.83e-07 $l=2.3e-07 $layer=LI1_cond $X=2.642 $Y=2.265
+ $X2=2.642 $Y2=2.035
r100 36 44 29.3759 $w=1.83e-07 $l=4.9e-07 $layer=LI1_cond $X=2.642 $Y=1.175
+ $X2=2.642 $Y2=1.665
r101 36 37 1.88775 $w=1.85e-07 $l=3.09167e-07 $layer=LI1_cond $X=2.642 $Y=1.175
+ $X2=2.41 $Y2=0.995
r102 32 34 24.0778 $w=2.78e-07 $l=5.85e-07 $layer=LI1_cond $X=4.54 $Y=1.005
+ $X2=4.54 $Y2=0.42
r103 31 37 4.40132 $w=1.7e-07 $l=3.745e-07 $layer=LI1_cond $X=2.74 $Y=1.09
+ $X2=2.41 $Y2=0.995
r104 30 32 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.4 $Y=1.09
+ $X2=4.54 $Y2=1.005
r105 30 31 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=4.4 $Y=1.09
+ $X2=2.74 $Y2=1.09
r106 27 38 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=2.735 $Y=2.35
+ $X2=2.642 $Y2=2.265
r107 27 29 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.735 $Y=2.35
+ $X2=3.225 $Y2=2.35
r108 26 39 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.92 $Y=2.35
+ $X2=4.08 $Y2=2.35
r109 26 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.92 $Y=2.35
+ $X2=3.225 $Y2=2.35
r110 22 37 1.88775 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0.995
+ $X2=2.41 $Y2=0.995
r111 22 24 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=2.575 $Y=0.995
+ $X2=2.575 $Y2=0.41
r112 20 37 4.40132 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=1.08
+ $X2=2.41 $Y2=0.995
r113 20 21 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=2.41 $Y=1.08
+ $X2=0.69 $Y2=1.08
r114 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.565 $Y=0.995
+ $X2=0.69 $Y2=1.08
r115 16 18 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=0.565 $Y=0.995
+ $X2=0.565 $Y2=0.42
r116 5 42 600 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.835 $X2=4.085 $Y2=2.43
r117 4 29 600 $w=1.7e-07 $l=5.98268e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=1.835 $X2=3.225 $Y2=2.35
r118 3 34 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.375
+ $Y=0.235 $X2=4.515 $Y2=0.42
r119 2 24 91 $w=1.7e-07 $l=3.05205e-07 $layer=licon1_NDIFF $count=2 $X=2.345
+ $Y=0.235 $X2=2.575 $Y2=0.41
r120 1 18 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.48
+ $Y=0.235 $X2=0.605 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_2%A_179_47# 1 2 9 11 12 15
r28 13 15 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.055 $Y=0.655
+ $X2=2.055 $Y2=0.37
r29 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.89 $Y=0.74
+ $X2=2.055 $Y2=0.655
r30 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.89 $Y=0.74 $X2=1.2
+ $Y2=0.74
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.035 $Y=0.655
+ $X2=1.2 $Y2=0.74
r32 7 9 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.035 $Y=0.655
+ $X2=1.035 $Y2=0.37
r33 2 15 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.915
+ $Y=0.235 $X2=2.055 $Y2=0.37
r34 1 9 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=0.895
+ $Y=0.235 $X2=1.035 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_2%VGND 1 2 9 13 15 17 25 32 33 36 39
r63 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r64 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r65 33 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r66 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r67 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.82 $Y=0 $X2=3.655
+ $Y2=0
r68 30 32 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.82 $Y=0 $X2=4.56
+ $Y2=0
r69 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r70 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r71 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.545
+ $Y2=0
r72 26 28 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=1.71 $Y=0 $X2=3.12
+ $Y2=0
r73 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.49 $Y=0 $X2=3.655
+ $Y2=0
r74 25 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.49 $Y=0 $X2=3.12
+ $Y2=0
r75 24 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r76 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r77 20 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r78 19 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r79 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r80 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=0 $X2=1.545
+ $Y2=0
r81 17 23 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.38 $Y=0 $X2=1.2
+ $Y2=0
r82 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r83 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r84 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0.085
+ $X2=3.655 $Y2=0
r85 11 13 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.655 $Y=0.085
+ $X2=3.655 $Y2=0.395
r86 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=0.085
+ $X2=1.545 $Y2=0
r87 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.545 $Y=0.085
+ $X2=1.545 $Y2=0.36
r88 2 13 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.655 $Y2=0.395
r89 1 9 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=1.325
+ $Y=0.235 $X2=1.545 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_2%A_595_47# 1 2 9 11 12 14
r19 14 16 3.84148 $w=2.38e-07 $l=8e-08 $layer=LI1_cond $X=4.11 $Y=0.67 $X2=4.11
+ $Y2=0.75
r20 11 16 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.99 $Y=0.75 $X2=4.11
+ $Y2=0.75
r21 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.99 $Y=0.75
+ $X2=3.32 $Y2=0.75
r22 7 12 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.15 $Y=0.665
+ $X2=3.32 $Y2=0.75
r23 7 9 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=3.15 $Y=0.665
+ $X2=3.15 $Y2=0.37
r24 2 14 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=3.945
+ $Y=0.235 $X2=4.085 $Y2=0.67
r25 1 9 91 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=2 $X=2.975
+ $Y=0.235 $X2=3.145 $Y2=0.37
.ends

