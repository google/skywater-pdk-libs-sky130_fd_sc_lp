* File: sky130_fd_sc_lp__o41ai_4.pex.spice
* Created: Fri Aug 28 11:20:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41AI_4%B1 3 7 11 15 19 23 27 31 33 34 35 36 37 38
+ 45 65 66
r90 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.65
+ $Y=1.46 $X2=2.65 $Y2=1.46
r91 63 65 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.59 $Y=1.46 $X2=2.65
+ $Y2=1.46
r92 62 63 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.16 $Y=1.46
+ $X2=2.59 $Y2=1.46
r93 60 62 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.97 $Y=1.46
+ $X2=2.16 $Y2=1.46
r94 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.46 $X2=1.97 $Y2=1.46
r95 58 60 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.73 $Y=1.46
+ $X2=1.97 $Y2=1.46
r96 56 58 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.63 $Y=1.46 $X2=1.73
+ $Y2=1.46
r97 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.46 $X2=1.63 $Y2=1.46
r98 54 56 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.3 $Y=1.46 $X2=1.63
+ $Y2=1.46
r99 53 57 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=1.29 $Y=1.567
+ $X2=1.63 $Y2=1.567
r100 52 54 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.29 $Y=1.46 $X2=1.3
+ $Y2=1.46
r101 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.29
+ $Y=1.46 $X2=1.29 $Y2=1.46
r102 50 52 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.87 $Y=1.46
+ $X2=1.29 $Y2=1.46
r103 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.46 $X2=0.61 $Y2=1.46
r104 45 50 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.795 $Y=1.46
+ $X2=0.87 $Y2=1.46
r105 45 47 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.795 $Y=1.46
+ $X2=0.61 $Y2=1.46
r106 38 66 0.299336 $w=3.83e-07 $l=1e-08 $layer=LI1_cond $X=2.64 $Y=1.567
+ $X2=2.65 $Y2=1.567
r107 37 38 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.567
+ $X2=2.64 $Y2=1.567
r108 37 61 5.68738 $w=3.83e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=1.567
+ $X2=1.97 $Y2=1.567
r109 36 61 8.68074 $w=3.83e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=1.567
+ $X2=1.97 $Y2=1.567
r110 36 57 1.49668 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=1.68 $Y=1.567
+ $X2=1.63 $Y2=1.567
r111 35 53 2.69402 $w=3.83e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.567 $X2=1.29
+ $Y2=1.567
r112 34 35 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.567
+ $X2=1.2 $Y2=1.567
r113 34 48 3.29269 $w=3.83e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.567
+ $X2=0.61 $Y2=1.567
r114 33 48 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.567
+ $X2=0.61 $Y2=1.567
r115 29 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.295
+ $X2=2.59 $Y2=1.46
r116 29 31 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.59 $Y=1.295
+ $X2=2.59 $Y2=0.655
r117 25 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.625
+ $X2=2.16 $Y2=1.46
r118 25 27 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.16 $Y=1.625
+ $X2=2.16 $Y2=2.465
r119 21 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.46
r120 21 23 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=0.655
r121 17 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.625
+ $X2=1.73 $Y2=1.46
r122 17 19 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.73 $Y=1.625
+ $X2=1.73 $Y2=2.465
r123 13 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.46
r124 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=0.655
r125 9 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.3 $Y=1.625
+ $X2=1.3 $Y2=1.46
r126 9 11 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.3 $Y=1.625 $X2=1.3
+ $Y2=2.465
r127 5 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.3 $Y=1.295
+ $X2=1.3 $Y2=1.46
r128 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.3 $Y=1.295 $X2=1.3
+ $Y2=0.655
r129 1 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.87 $Y=1.625
+ $X2=0.87 $Y2=1.46
r130 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.87 $Y=1.625
+ $X2=0.87 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%A4 1 3 6 10 12 14 17 19 21 24 26 28 31 34 35
+ 48 50 57
c97 24 0 5.30626e-20 $X=4.4 $Y=2.435
r98 45 46 8.58524 $w=3.93e-07 $l=7e-08 $layer=POLY_cond $X=3.97 $Y=1.395
+ $X2=4.04 $Y2=1.395
r99 44 45 44.1527 $w=3.93e-07 $l=3.6e-07 $layer=POLY_cond $X=3.61 $Y=1.395
+ $X2=3.97 $Y2=1.395
r100 43 44 8.58524 $w=3.93e-07 $l=7e-08 $layer=POLY_cond $X=3.54 $Y=1.395
+ $X2=3.61 $Y2=1.395
r101 42 50 8.05287 $w=4.03e-07 $l=2.83e-07 $layer=LI1_cond $X=3.2 $Y=1.557
+ $X2=3.483 $Y2=1.557
r102 41 43 41.6997 $w=3.93e-07 $l=3.4e-07 $layer=POLY_cond $X=3.2 $Y=1.395
+ $X2=3.54 $Y2=1.395
r103 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.44 $X2=3.2 $Y2=1.44
r104 39 41 11.0382 $w=3.93e-07 $l=9e-08 $layer=POLY_cond $X=3.11 $Y=1.395
+ $X2=3.2 $Y2=1.395
r105 38 39 1.22646 $w=3.93e-07 $l=1e-08 $layer=POLY_cond $X=3.1 $Y=1.395
+ $X2=3.11 $Y2=1.395
r106 35 57 6.39237 $w=4.03e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=1.557
+ $X2=3.685 $Y2=1.557
r107 35 50 3.32928 $w=4.03e-07 $l=1.17e-07 $layer=LI1_cond $X=3.6 $Y=1.557
+ $X2=3.483 $Y2=1.557
r108 34 42 2.27643 $w=4.03e-07 $l=8e-08 $layer=LI1_cond $X=3.12 $Y=1.557 $X2=3.2
+ $Y2=1.557
r109 32 48 38.0204 $w=3.93e-07 $l=3.1e-07 $layer=POLY_cond $X=4.09 $Y=1.395
+ $X2=4.4 $Y2=1.395
r110 32 46 6.13232 $w=3.93e-07 $l=5e-08 $layer=POLY_cond $X=4.09 $Y=1.395
+ $X2=4.04 $Y2=1.395
r111 31 57 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.09 $Y=1.44
+ $X2=3.685 $Y2=1.44
r112 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.09
+ $Y=1.44 $X2=4.09 $Y2=1.44
r113 26 48 19.6234 $w=3.93e-07 $l=2.78747e-07 $layer=POLY_cond $X=4.56 $Y=1.185
+ $X2=4.4 $Y2=1.395
r114 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.56 $Y=1.185
+ $X2=4.56 $Y2=0.655
r115 22 48 25.4309 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.4 $Y=1.605
+ $X2=4.4 $Y2=1.395
r116 22 24 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.4 $Y=1.605
+ $X2=4.4 $Y2=2.435
r117 19 46 25.4309 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.04 $Y=1.185
+ $X2=4.04 $Y2=1.395
r118 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.04 $Y=1.185
+ $X2=4.04 $Y2=0.655
r119 15 45 25.4309 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.97 $Y=1.605
+ $X2=3.97 $Y2=1.395
r120 15 17 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.97 $Y=1.605
+ $X2=3.97 $Y2=2.435
r121 12 44 25.4309 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.61 $Y=1.185
+ $X2=3.61 $Y2=1.395
r122 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.61 $Y=1.185
+ $X2=3.61 $Y2=0.655
r123 8 43 25.4309 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.54 $Y=1.605
+ $X2=3.54 $Y2=1.395
r124 8 10 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.54 $Y=1.605
+ $X2=3.54 $Y2=2.435
r125 4 39 25.4309 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=1.395
r126 4 6 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=2.435
r127 1 38 25.4309 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.1 $Y=1.185 $X2=3.1
+ $Y2=1.395
r128 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.1 $Y=1.185 $X2=3.1
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%A3 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 48
c100 48 0 1.2076e-19 $X=6.37 $Y=1.48
c101 22 0 1.91349e-19 $X=6.12 $Y=1.695
c102 1 0 7.8353e-20 $X=4.83 $Y=1.695
r103 48 50 7.8587 $w=3.68e-07 $l=6e-08 $layer=POLY_cond $X=6.37 $Y=1.505
+ $X2=6.43 $Y2=1.505
r104 48 49 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.37
+ $Y=1.48 $X2=6.37 $Y2=1.48
r105 46 48 32.7446 $w=3.68e-07 $l=2.5e-07 $layer=POLY_cond $X=6.12 $Y=1.505
+ $X2=6.37 $Y2=1.505
r106 45 46 15.7174 $w=3.68e-07 $l=1.2e-07 $layer=POLY_cond $X=6 $Y=1.505
+ $X2=6.12 $Y2=1.505
r107 44 45 40.6033 $w=3.68e-07 $l=3.1e-07 $layer=POLY_cond $X=5.69 $Y=1.505
+ $X2=6 $Y2=1.505
r108 43 44 15.7174 $w=3.68e-07 $l=1.2e-07 $layer=POLY_cond $X=5.57 $Y=1.505
+ $X2=5.69 $Y2=1.505
r109 42 43 40.6033 $w=3.68e-07 $l=3.1e-07 $layer=POLY_cond $X=5.26 $Y=1.505
+ $X2=5.57 $Y2=1.505
r110 41 42 26.1957 $w=3.68e-07 $l=2e-07 $layer=POLY_cond $X=5.06 $Y=1.505
+ $X2=5.26 $Y2=1.505
r111 39 41 6.54891 $w=3.68e-07 $l=5e-08 $layer=POLY_cond $X=5.01 $Y=1.505
+ $X2=5.06 $Y2=1.505
r112 39 40 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.01
+ $Y=1.48 $X2=5.01 $Y2=1.48
r113 32 49 3.13009 $w=4.03e-07 $l=1.1e-07 $layer=LI1_cond $X=6.48 $Y=1.547
+ $X2=6.37 $Y2=1.547
r114 31 49 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=6 $Y=1.547 $X2=6.37
+ $Y2=1.547
r115 30 31 13.6586 $w=4.03e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.547 $X2=6
+ $Y2=1.547
r116 29 30 13.6586 $w=4.03e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.547
+ $X2=5.52 $Y2=1.547
r117 29 40 0.853661 $w=4.03e-07 $l=3e-08 $layer=LI1_cond $X=5.04 $Y=1.547
+ $X2=5.01 $Y2=1.547
r118 25 50 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.43 $Y=1.315
+ $X2=6.43 $Y2=1.505
r119 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.43 $Y=1.315
+ $X2=6.43 $Y2=0.655
r120 22 46 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.12 $Y=1.695
+ $X2=6.12 $Y2=1.505
r121 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.12 $Y=1.695
+ $X2=6.12 $Y2=2.435
r122 18 45 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6 $Y=1.315 $X2=6
+ $Y2=1.505
r123 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6 $Y=1.315 $X2=6
+ $Y2=0.655
r124 15 44 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.69 $Y=1.695
+ $X2=5.69 $Y2=1.505
r125 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.69 $Y=1.695
+ $X2=5.69 $Y2=2.435
r126 11 43 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.57 $Y=1.315
+ $X2=5.57 $Y2=1.505
r127 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.57 $Y=1.315
+ $X2=5.57 $Y2=0.655
r128 8 42 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.26 $Y=1.695
+ $X2=5.26 $Y2=1.505
r129 8 10 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.26 $Y=1.695
+ $X2=5.26 $Y2=2.435
r130 4 41 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.06 $Y=1.315
+ $X2=5.06 $Y2=1.505
r131 4 6 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.06 $Y=1.315
+ $X2=5.06 $Y2=0.655
r132 1 39 23.5761 $w=3.68e-07 $l=2.65141e-07 $layer=POLY_cond $X=4.83 $Y=1.695
+ $X2=5.01 $Y2=1.505
r133 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.83 $Y=1.695
+ $X2=4.83 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%A2 3 7 11 15 19 23 27 31 38 41 56 62
c101 62 0 1.91349e-19 $X=7.335 $Y=1.547
c102 38 0 2.82898e-20 $X=8.27 $Y=1.44
r103 55 56 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.285 $Y=1.44
+ $X2=8.36 $Y2=1.44
r104 52 53 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.72 $Y=1.44
+ $X2=7.93 $Y2=1.44
r105 49 50 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.29 $Y=1.44
+ $X2=7.5 $Y2=1.44
r106 48 62 6.02733 $w=4.03e-07 $l=8.5e-08 $layer=LI1_cond $X=7.25 $Y=1.547
+ $X2=7.335 $Y2=1.547
r107 47 49 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=7.25 $Y=1.44 $X2=7.29
+ $Y2=1.44
r108 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.25
+ $Y=1.44 $X2=7.25 $Y2=1.44
r109 45 47 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.07 $Y=1.44
+ $X2=7.25 $Y2=1.44
r110 43 45 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=6.86 $Y=1.44
+ $X2=7.07 $Y2=1.44
r111 41 48 8.25206 $w=4.03e-07 $l=2.9e-07 $layer=LI1_cond $X=6.96 $Y=1.547
+ $X2=7.25 $Y2=1.547
r112 39 55 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.27 $Y=1.44
+ $X2=8.285 $Y2=1.44
r113 39 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.27 $Y=1.44
+ $X2=7.93 $Y2=1.44
r114 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.27
+ $Y=1.44 $X2=8.27 $Y2=1.44
r115 36 52 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=7.59 $Y=1.44
+ $X2=7.72 $Y2=1.44
r116 36 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.59 $Y=1.44 $X2=7.5
+ $Y2=1.44
r117 35 38 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=7.59 $Y=1.435
+ $X2=8.27 $Y2=1.435
r118 35 62 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=7.59 $Y=1.435
+ $X2=7.335 $Y2=1.435
r119 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.59
+ $Y=1.44 $X2=7.59 $Y2=1.44
r120 29 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.36 $Y=1.605
+ $X2=8.36 $Y2=1.44
r121 29 31 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.36 $Y=1.605
+ $X2=8.36 $Y2=2.465
r122 25 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.285 $Y=1.275
+ $X2=8.285 $Y2=1.44
r123 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.285 $Y=1.275
+ $X2=8.285 $Y2=0.655
r124 21 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.93 $Y=1.605
+ $X2=7.93 $Y2=1.44
r125 21 23 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.93 $Y=1.605
+ $X2=7.93 $Y2=2.465
r126 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.72 $Y=1.275
+ $X2=7.72 $Y2=1.44
r127 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.72 $Y=1.275
+ $X2=7.72 $Y2=0.655
r128 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.5 $Y=1.605
+ $X2=7.5 $Y2=1.44
r129 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.5 $Y=1.605
+ $X2=7.5 $Y2=2.465
r130 9 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.29 $Y=1.275
+ $X2=7.29 $Y2=1.44
r131 9 11 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.29 $Y=1.275
+ $X2=7.29 $Y2=0.655
r132 5 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.07 $Y=1.605
+ $X2=7.07 $Y2=1.44
r133 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.07 $Y=1.605
+ $X2=7.07 $Y2=2.465
r134 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.86 $Y=1.275
+ $X2=6.86 $Y2=1.44
r135 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.86 $Y=1.275
+ $X2=6.86 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 46
c69 6 0 2.82898e-20 $X=8.79 $Y=2.465
r70 44 46 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=10.08 $Y=1.35
+ $X2=10.29 $Y2=1.35
r71 43 44 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=10.01 $Y=1.35
+ $X2=10.08 $Y2=1.35
r72 42 43 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=9.65 $Y=1.35
+ $X2=10.01 $Y2=1.35
r73 41 42 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=9.58 $Y=1.35 $X2=9.65
+ $Y2=1.35
r74 40 41 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=9.22 $Y=1.35
+ $X2=9.58 $Y2=1.35
r75 39 40 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=9.15 $Y=1.35 $X2=9.22
+ $Y2=1.35
r76 37 39 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=8.93 $Y=1.35
+ $X2=9.15 $Y2=1.35
r77 37 38 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.93
+ $Y=1.35 $X2=8.93 $Y2=1.35
r78 35 37 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=8.79 $Y=1.35
+ $X2=8.93 $Y2=1.35
r79 33 35 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.72 $Y=1.35 $X2=8.79
+ $Y2=1.35
r80 30 46 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=10.29
+ $Y=1.35 $X2=10.29 $Y2=1.35
r81 29 30 16.4635 $w=3.13e-07 $l=4.5e-07 $layer=LI1_cond $X=9.84 $Y=1.367
+ $X2=10.29 $Y2=1.367
r82 29 38 33.2928 $w=3.13e-07 $l=9.1e-07 $layer=LI1_cond $X=9.84 $Y=1.367
+ $X2=8.93 $Y2=1.367
r83 25 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.08 $Y=1.515
+ $X2=10.08 $Y2=1.35
r84 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=10.08 $Y=1.515
+ $X2=10.08 $Y2=2.465
r85 22 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.01 $Y=1.185
+ $X2=10.01 $Y2=1.35
r86 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.01 $Y=1.185
+ $X2=10.01 $Y2=0.655
r87 18 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.65 $Y=1.515
+ $X2=9.65 $Y2=1.35
r88 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.65 $Y=1.515
+ $X2=9.65 $Y2=2.465
r89 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.58 $Y=1.185
+ $X2=9.58 $Y2=1.35
r90 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.58 $Y=1.185
+ $X2=9.58 $Y2=0.655
r91 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.22 $Y=1.515
+ $X2=9.22 $Y2=1.35
r92 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.22 $Y=1.515
+ $X2=9.22 $Y2=2.465
r93 8 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.15 $Y=1.185
+ $X2=9.15 $Y2=1.35
r94 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.15 $Y=1.185
+ $X2=9.15 $Y2=0.655
r95 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.79 $Y=1.515
+ $X2=8.79 $Y2=1.35
r96 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.79 $Y=1.515 $X2=8.79
+ $Y2=2.465
r97 1 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.72 $Y=1.185
+ $X2=8.72 $Y2=1.35
r98 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.72 $Y=1.185 $X2=8.72
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%VPWR 1 2 3 4 5 18 24 28 32 38 43 44 46 47 48
+ 50 62 66 73 74 77 80 83
r129 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r130 80 81 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r131 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r132 74 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r133 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r134 71 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.03 $Y=3.33
+ $X2=9.865 $Y2=3.33
r135 71 73 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.03 $Y=3.33
+ $X2=10.32 $Y2=3.33
r136 70 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r137 70 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r138 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r139 67 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.17 $Y=3.33
+ $X2=9.005 $Y2=3.33
r140 67 69 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.17 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 66 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.7 $Y=3.33
+ $X2=9.865 $Y2=3.33
r142 66 69 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.7 $Y=3.33
+ $X2=9.36 $Y2=3.33
r143 64 65 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r144 62 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.84 $Y=3.33
+ $X2=9.005 $Y2=3.33
r145 62 64 404.492 $w=1.68e-07 $l=6.2e-06 $layer=LI1_cond $X=8.84 $Y=3.33
+ $X2=2.64 $Y2=3.33
r146 61 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r147 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r148 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r149 58 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r150 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r151 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.655 $Y2=3.33
r152 55 57 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=1.2 $Y2=3.33
r153 53 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r155 50 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.49 $Y=3.33
+ $X2=0.655 $Y2=3.33
r156 50 52 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.49 $Y=3.33
+ $X2=0.24 $Y2=3.33
r157 48 81 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=8.88 $Y2=3.33
r158 48 65 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=2.64 $Y2=3.33
r159 46 60 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.21 $Y=3.33 $X2=2.16
+ $Y2=3.33
r160 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=3.33
+ $X2=2.375 $Y2=3.33
r161 45 64 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.54 $Y=3.33 $X2=2.64
+ $Y2=3.33
r162 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=3.33
+ $X2=2.375 $Y2=3.33
r163 43 57 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.35 $Y=3.33 $X2=1.2
+ $Y2=3.33
r164 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.515 $Y2=3.33
r165 42 60 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r166 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=1.515 $Y2=3.33
r167 38 41 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=9.865 $Y=2.13
+ $X2=9.865 $Y2=2.95
r168 36 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.865 $Y=3.245
+ $X2=9.865 $Y2=3.33
r169 36 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.865 $Y=3.245
+ $X2=9.865 $Y2=2.95
r170 32 35 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=9.005 $Y=2.13
+ $X2=9.005 $Y2=2.95
r171 30 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.005 $Y=3.245
+ $X2=9.005 $Y2=3.33
r172 30 35 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.005 $Y=3.245
+ $X2=9.005 $Y2=2.95
r173 26 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=3.245
+ $X2=2.375 $Y2=3.33
r174 26 28 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=2.375 $Y=3.245
+ $X2=2.375 $Y2=2.395
r175 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.515 $Y=3.245
+ $X2=1.515 $Y2=3.33
r176 22 24 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=1.515 $Y=3.245
+ $X2=1.515 $Y2=2.395
r177 18 21 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=0.655 $Y=2.015
+ $X2=0.655 $Y2=2.95
r178 16 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.655 $Y=3.245
+ $X2=0.655 $Y2=3.33
r179 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.655 $Y=3.245
+ $X2=0.655 $Y2=2.95
r180 5 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.725
+ $Y=1.835 $X2=9.865 $Y2=2.95
r181 5 38 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=9.725
+ $Y=1.835 $X2=9.865 $Y2=2.13
r182 4 35 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.865
+ $Y=1.835 $X2=9.005 $Y2=2.95
r183 4 32 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=8.865
+ $Y=1.835 $X2=9.005 $Y2=2.13
r184 3 28 300 $w=1.7e-07 $l=6.26099e-07 $layer=licon1_PDIFF $count=2 $X=2.235
+ $Y=1.835 $X2=2.375 $Y2=2.395
r185 2 24 300 $w=1.7e-07 $l=6.26099e-07 $layer=licon1_PDIFF $count=2 $X=1.375
+ $Y=1.835 $X2=1.515 $Y2=2.395
r186 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.53
+ $Y=1.835 $X2=0.655 $Y2=2.95
r187 1 18 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.53
+ $Y=1.835 $X2=0.655 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%Y 1 2 3 4 5 6 19 21 23 27 29 30 33 35 39 41
+ 45 49 54 55 57 59 60 64 69
r109 64 71 15.735 $w=2.83e-07 $l=4.52913e-07 $layer=LI1_cond $X=4.55 $Y=1.705
+ $X2=4.185 $Y2=1.902
r110 64 69 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=4.55 $Y=1.705
+ $X2=4.55 $Y2=1.665
r111 60 64 0.431095 $w=2.83e-07 $l=2.6533e-08 $layer=LI1_cond $X=4.56 $Y=1.727
+ $X2=4.55 $Y2=1.705
r112 60 69 1.06025 $w=2.48e-07 $l=2.3e-08 $layer=LI1_cond $X=4.55 $Y=1.642
+ $X2=4.55 $Y2=1.665
r113 59 60 15.9959 $w=2.48e-07 $l=3.47e-07 $layer=LI1_cond $X=4.55 $Y=1.295
+ $X2=4.55 $Y2=1.642
r114 58 59 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=4.55 $Y=1.185
+ $X2=4.55 $Y2=1.295
r115 49 71 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=4.185 $Y=2.64
+ $X2=4.185 $Y2=2.1
r116 46 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.49 $Y=2.015
+ $X2=3.325 $Y2=2.015
r117 45 71 9.04317 $w=2.83e-07 $l=2.14173e-07 $layer=LI1_cond $X=4.02 $Y=2.015
+ $X2=4.185 $Y2=1.902
r118 45 46 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.02 $Y=2.015
+ $X2=3.49 $Y2=2.015
r119 42 55 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.47 $Y=1.1
+ $X2=2.375 $Y2=1.1
r120 41 58 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.425 $Y=1.1
+ $X2=4.55 $Y2=1.185
r121 41 42 127.545 $w=1.68e-07 $l=1.955e-06 $layer=LI1_cond $X=4.425 $Y=1.1
+ $X2=2.47 $Y2=1.1
r122 37 55 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=1.015
+ $X2=2.375 $Y2=1.1
r123 37 39 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=2.375 $Y=1.015
+ $X2=2.375 $Y2=0.76
r124 36 54 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.04 $Y=2.015 $X2=1.95
+ $Y2=2.015
r125 35 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=2.015
+ $X2=3.325 $Y2=2.015
r126 35 36 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=3.16 $Y=2.015
+ $X2=2.04 $Y2=2.015
r127 31 54 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=2.1 $X2=1.95
+ $Y2=2.015
r128 31 33 24.6465 $w=1.78e-07 $l=4e-07 $layer=LI1_cond $X=1.95 $Y=2.1 $X2=1.95
+ $Y2=2.5
r129 29 55 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.28 $Y=1.1
+ $X2=2.375 $Y2=1.1
r130 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.28 $Y=1.1
+ $X2=1.61 $Y2=1.1
r131 25 30 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.497 $Y=1.015
+ $X2=1.61 $Y2=1.1
r132 25 27 13.061 $w=2.23e-07 $l=2.55e-07 $layer=LI1_cond $X=1.497 $Y=1.015
+ $X2=1.497 $Y2=0.76
r133 24 52 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.18 $Y=2.015
+ $X2=1.085 $Y2=2.015
r134 23 54 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.86 $Y=2.015 $X2=1.95
+ $Y2=2.015
r135 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.86 $Y=2.015
+ $X2=1.18 $Y2=2.015
r136 19 52 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=2.1
+ $X2=1.085 $Y2=2.015
r137 19 21 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=1.085 $Y=2.1
+ $X2=1.085 $Y2=2.91
r138 6 71 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.805 $X2=4.185 $Y2=1.93
r139 6 49 400 $w=1.7e-07 $l=9.02289e-07 $layer=licon1_PDIFF $count=1 $X=4.045
+ $Y=1.805 $X2=4.185 $Y2=2.64
r140 5 57 300 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=2 $X=3.185
+ $Y=1.805 $X2=3.325 $Y2=2.045
r141 4 54 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=1.805
+ $Y=1.835 $X2=1.945 $Y2=2.015
r142 4 33 300 $w=1.7e-07 $l=7.31659e-07 $layer=licon1_PDIFF $count=2 $X=1.805
+ $Y=1.835 $X2=1.945 $Y2=2.5
r143 3 52 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=0.945
+ $Y=1.835 $X2=1.085 $Y2=2.095
r144 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.945
+ $Y=1.835 $X2=1.085 $Y2=2.91
r145 2 39 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.235 $X2=2.375 $Y2=0.76
r146 1 27 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=1.375
+ $Y=0.235 $X2=1.515 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%A_554_361# 1 2 3 4 5 18 20 21 24 26 29 30 31
+ 34 36 38 40 42 48
c66 29 0 7.8353e-20 $X=4.615 $Y=2.895
r67 38 50 3.71573 $w=2.6e-07 $l=1.53e-07 $layer=LI1_cond $X=6.37 $Y=2.225
+ $X2=6.37 $Y2=2.072
r68 38 40 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.37 $Y=2.225
+ $X2=6.37 $Y2=2.52
r69 37 48 3.42911 $w=3.05e-07 $l=9.5e-08 $layer=LI1_cond $X=5.57 $Y=2.072
+ $X2=5.475 $Y2=2.072
r70 36 50 3.15716 $w=3.05e-07 $l=1.3e-07 $layer=LI1_cond $X=6.24 $Y=2.072
+ $X2=6.37 $Y2=2.072
r71 36 37 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=6.24 $Y=2.072
+ $X2=5.57 $Y2=2.072
r72 32 48 3.09063 $w=1.9e-07 $l=1.53e-07 $layer=LI1_cond $X=5.475 $Y=2.225
+ $X2=5.475 $Y2=2.072
r73 32 34 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=5.475 $Y=2.225
+ $X2=5.475 $Y2=2.52
r74 31 44 16.2691 $w=3.05e-07 $l=3.82e-07 $layer=LI1_cond $X=4.997 $Y=2.072
+ $X2=4.615 $Y2=2.072
r75 30 48 3.42911 $w=3.05e-07 $l=9.5e-08 $layer=LI1_cond $X=5.38 $Y=2.072
+ $X2=5.475 $Y2=2.072
r76 30 31 14.4717 $w=3.03e-07 $l=3.83e-07 $layer=LI1_cond $X=5.38 $Y=2.072
+ $X2=4.997 $Y2=2.072
r77 29 46 3.31928 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=4.615 $Y=2.895
+ $X2=4.615 $Y2=2.985
r78 28 44 1.56892 $w=1.9e-07 $l=1.53e-07 $layer=LI1_cond $X=4.615 $Y=2.225
+ $X2=4.615 $Y2=2.072
r79 28 29 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=4.615 $Y=2.225
+ $X2=4.615 $Y2=2.895
r80 27 42 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.85 $Y=2.985
+ $X2=3.755 $Y2=2.985
r81 26 46 3.50369 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.52 $Y=2.985
+ $X2=4.615 $Y2=2.985
r82 26 27 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.52 $Y=2.985
+ $X2=3.85 $Y2=2.985
r83 22 42 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=3.755 $Y=2.895
+ $X2=3.755 $Y2=2.985
r84 22 24 26.8517 $w=1.88e-07 $l=4.6e-07 $layer=LI1_cond $X=3.755 $Y=2.895
+ $X2=3.755 $Y2=2.435
r85 20 42 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.66 $Y=2.985
+ $X2=3.755 $Y2=2.985
r86 20 21 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.66 $Y=2.985
+ $X2=2.99 $Y2=2.985
r87 16 21 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=2.86 $Y=2.895
+ $X2=2.99 $Y2=2.985
r88 16 18 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=2.86 $Y=2.895
+ $X2=2.86 $Y2=2.435
r89 5 50 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=6.195
+ $Y=1.805 $X2=6.335 $Y2=2.005
r90 5 40 600 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_PDIFF $count=1 $X=6.195
+ $Y=1.805 $X2=6.335 $Y2=2.52
r91 4 48 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.805 $X2=5.475 $Y2=2.085
r92 4 34 600 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.805 $X2=5.475 $Y2=2.52
r93 3 46 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.805 $X2=4.615 $Y2=2.91
r94 3 44 400 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.805 $X2=4.615 $Y2=2.21
r95 2 24 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=3.615
+ $Y=1.805 $X2=3.755 $Y2=2.435
r96 1 18 300 $w=1.7e-07 $l=6.89674e-07 $layer=licon1_PDIFF $count=2 $X=2.77
+ $Y=1.805 $X2=2.895 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%A_981_361# 1 2 3 4 15 17 18 21 23 27 29 31
+ 33 35 36
c66 18 0 5.30626e-20 $X=5.21 $Y=2.965
c67 15 0 1.2076e-19 $X=5.045 $Y=2.48
r68 31 38 3.95267 $w=2.6e-07 $l=1.7e-07 $layer=LI1_cond $X=8.18 $Y=2.735
+ $X2=8.18 $Y2=2.905
r69 31 33 23.2705 $w=2.58e-07 $l=5.25e-07 $layer=LI1_cond $X=8.18 $Y=2.735
+ $X2=8.18 $Y2=2.21
r70 30 36 5.90962 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=2.905
+ $X2=7.285 $Y2=2.905
r71 29 38 3.02263 $w=3.4e-07 $l=1.3e-07 $layer=LI1_cond $X=8.05 $Y=2.905
+ $X2=8.18 $Y2=2.905
r72 29 30 20.3372 $w=3.38e-07 $l=6e-07 $layer=LI1_cond $X=8.05 $Y=2.905 $X2=7.45
+ $Y2=2.905
r73 25 36 0.758147 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=7.285 $Y=2.735
+ $X2=7.285 $Y2=2.905
r74 25 27 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=7.285 $Y=2.735
+ $X2=7.285 $Y2=2.355
r75 24 35 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.07 $Y=2.965
+ $X2=5.905 $Y2=2.965
r76 23 36 5.90962 $w=2.8e-07 $l=1.92678e-07 $layer=LI1_cond $X=7.12 $Y=2.965
+ $X2=7.285 $Y2=2.905
r77 23 24 55.003 $w=2.18e-07 $l=1.05e-06 $layer=LI1_cond $X=7.12 $Y=2.965
+ $X2=6.07 $Y2=2.965
r78 19 35 0.067832 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=5.905 $Y=2.855
+ $X2=5.905 $Y2=2.965
r79 19 21 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.905 $Y=2.855
+ $X2=5.905 $Y2=2.48
r80 17 35 7.13466 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.74 $Y=2.965
+ $X2=5.905 $Y2=2.965
r81 17 18 27.7634 $w=2.18e-07 $l=5.3e-07 $layer=LI1_cond $X=5.74 $Y=2.965
+ $X2=5.21 $Y2=2.965
r82 13 18 7.17723 $w=2.2e-07 $l=2.13014e-07 $layer=LI1_cond $X=5.045 $Y=2.855
+ $X2=5.21 $Y2=2.965
r83 13 15 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.045 $Y=2.855
+ $X2=5.045 $Y2=2.48
r84 4 38 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.005
+ $Y=1.835 $X2=8.145 $Y2=2.91
r85 4 33 300 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=2 $X=8.005
+ $Y=1.835 $X2=8.145 $Y2=2.21
r86 3 27 300 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=2 $X=7.145
+ $Y=1.835 $X2=7.285 $Y2=2.355
r87 2 21 300 $w=1.7e-07 $l=7.41704e-07 $layer=licon1_PDIFF $count=2 $X=5.765
+ $Y=1.805 $X2=5.905 $Y2=2.48
r88 1 15 300 $w=1.7e-07 $l=7.41704e-07 $layer=licon1_PDIFF $count=2 $X=4.905
+ $Y=1.805 $X2=5.045 $Y2=2.48
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%A_1346_367# 1 2 3 4 5 16 18 20 24 26 30 34
+ 38 42 46 52 57 58
r70 55 56 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=7.75 $Y=1.98 $X2=7.75
+ $Y2=2.01
r71 52 55 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=7.75 $Y=1.785
+ $X2=7.75 $Y2=1.98
r72 46 48 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=10.33 $Y=1.98
+ $X2=10.33 $Y2=2.91
r73 44 46 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=10.33 $Y=1.875
+ $X2=10.33 $Y2=1.98
r74 43 58 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=9.53 $Y=1.785
+ $X2=9.435 $Y2=1.785
r75 42 44 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=10.2 $Y=1.785
+ $X2=10.33 $Y2=1.875
r76 42 43 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=10.2 $Y=1.785
+ $X2=9.53 $Y2=1.785
r77 38 40 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=9.435 $Y=1.98
+ $X2=9.435 $Y2=2.91
r78 36 58 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=9.435 $Y=1.875
+ $X2=9.435 $Y2=1.785
r79 36 38 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=9.435 $Y=1.875
+ $X2=9.435 $Y2=1.98
r80 35 57 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=8.67 $Y=1.785
+ $X2=8.575 $Y2=1.785
r81 34 58 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=9.34 $Y=1.785
+ $X2=9.435 $Y2=1.785
r82 34 35 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=9.34 $Y=1.785
+ $X2=8.67 $Y2=1.785
r83 30 32 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=8.575 $Y=1.98
+ $X2=8.575 $Y2=2.91
r84 28 57 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=8.575 $Y=1.875
+ $X2=8.575 $Y2=1.785
r85 28 30 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=8.575 $Y=1.875
+ $X2=8.575 $Y2=1.98
r86 27 52 2.89065 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=7.88 $Y=1.785
+ $X2=7.75 $Y2=1.785
r87 26 57 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=8.48 $Y=1.785
+ $X2=8.575 $Y2=1.785
r88 26 27 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=8.48 $Y=1.785 $X2=7.88
+ $Y2=1.785
r89 22 56 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=7.75 $Y=2.1 $X2=7.75
+ $Y2=2.01
r90 22 24 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=7.75 $Y=2.1
+ $X2=7.75 $Y2=2.325
r91 21 51 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=6.95 $Y=2.01 $X2=6.82
+ $Y2=2.01
r92 20 56 2.89065 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=7.62 $Y=2.01 $X2=7.75
+ $Y2=2.01
r93 20 21 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.62 $Y=2.01
+ $X2=6.95 $Y2=2.01
r94 16 51 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=6.82 $Y=2.1 $X2=6.82
+ $Y2=2.01
r95 16 18 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=6.82 $Y=2.1 $X2=6.82
+ $Y2=2.52
r96 5 48 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.835 $X2=10.295 $Y2=2.91
r97 5 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.835 $X2=10.295 $Y2=1.98
r98 4 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.295
+ $Y=1.835 $X2=9.435 $Y2=2.91
r99 4 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.295
+ $Y=1.835 $X2=9.435 $Y2=1.98
r100 3 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.435
+ $Y=1.835 $X2=8.575 $Y2=2.91
r101 3 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.435
+ $Y=1.835 $X2=8.575 $Y2=1.98
r102 2 55 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.575
+ $Y=1.835 $X2=7.715 $Y2=1.98
r103 2 24 600 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=1 $X=7.575
+ $Y=1.835 $X2=7.715 $Y2=2.325
r104 1 51 600 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.835 $X2=6.855 $Y2=2.005
r105 1 18 600 $w=1.7e-07 $l=7.44883e-07 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.835 $X2=6.855 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%A_192_47# 1 2 3 4 5 6 7 8 9 10 11 36 38 39
+ 42 44 45 46 47 50 52 56 59 60 61 64 66 70 72 76 78 82 84 88 90 94 97 100 101
+ 102 103 104 105 107
r169 105 106 6.16854 $w=2.67e-07 $l=1.35e-07 $layer=LI1_cond $X=8.482 $Y=0.955
+ $X2=8.482 $Y2=1.09
r170 92 94 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=10.25 $Y=0.87
+ $X2=10.25 $Y2=0.42
r171 91 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.49 $Y=0.955
+ $X2=9.365 $Y2=0.955
r172 90 92 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=10.11 $Y=0.955
+ $X2=10.25 $Y2=0.87
r173 90 91 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=10.11 $Y=0.955
+ $X2=9.49 $Y2=0.955
r174 86 107 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.365 $Y=0.87
+ $X2=9.365 $Y2=0.955
r175 86 88 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=9.365 $Y=0.87
+ $X2=9.365 $Y2=0.42
r176 85 105 3.37873 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=8.625 $Y=0.955
+ $X2=8.482 $Y2=0.955
r177 84 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.24 $Y=0.955
+ $X2=9.365 $Y2=0.955
r178 84 85 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=9.24 $Y=0.955
+ $X2=8.625 $Y2=0.955
r179 80 105 3.70346 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=8.482 $Y=0.87
+ $X2=8.482 $Y2=0.955
r180 80 82 18.1965 $w=2.83e-07 $l=4.5e-07 $layer=LI1_cond $X=8.482 $Y=0.87
+ $X2=8.482 $Y2=0.42
r181 79 104 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.67 $Y=1.09
+ $X2=7.54 $Y2=1.09
r182 78 106 3.37873 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=8.34 $Y=1.09
+ $X2=8.482 $Y2=1.09
r183 78 79 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.34 $Y=1.09
+ $X2=7.67 $Y2=1.09
r184 74 104 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.54 $Y=1.005
+ $X2=7.54 $Y2=1.09
r185 74 76 25.93 $w=2.58e-07 $l=5.85e-07 $layer=LI1_cond $X=7.54 $Y=1.005
+ $X2=7.54 $Y2=0.42
r186 73 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.74 $Y=1.09
+ $X2=6.645 $Y2=1.09
r187 72 104 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.41 $Y=1.09
+ $X2=7.54 $Y2=1.09
r188 72 73 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.41 $Y=1.09
+ $X2=6.74 $Y2=1.09
r189 68 103 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=1.005
+ $X2=6.645 $Y2=1.09
r190 68 70 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=6.645 $Y=1.005
+ $X2=6.645 $Y2=0.42
r191 67 102 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.88 $Y=1.09
+ $X2=5.785 $Y2=1.09
r192 66 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.55 $Y=1.09
+ $X2=6.645 $Y2=1.09
r193 66 67 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.55 $Y=1.09
+ $X2=5.88 $Y2=1.09
r194 62 102 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=1.005
+ $X2=5.785 $Y2=1.09
r195 62 64 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=5.785 $Y=1.005
+ $X2=5.785 $Y2=0.42
r196 60 102 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.69 $Y=1.09
+ $X2=5.785 $Y2=1.09
r197 60 61 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.69 $Y=1.09
+ $X2=5.015 $Y2=1.09
r198 59 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.93 $Y=1.005
+ $X2=5.015 $Y2=1.09
r199 58 101 3.67481 $w=2.52e-07 $l=1.19499e-07 $layer=LI1_cond $X=4.93 $Y=0.845
+ $X2=4.847 $Y2=0.76
r200 58 59 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.93 $Y=0.845
+ $X2=4.93 $Y2=1.005
r201 54 101 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=4.847 $Y=0.675
+ $X2=4.847 $Y2=0.76
r202 54 56 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=4.847 $Y=0.675
+ $X2=4.847 $Y2=0.38
r203 53 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=0.76
+ $X2=3.825 $Y2=0.76
r204 52 101 2.79892 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=4.68 $Y=0.76
+ $X2=4.847 $Y2=0.76
r205 52 53 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.68 $Y=0.76
+ $X2=3.99 $Y2=0.76
r206 48 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=0.675
+ $X2=3.825 $Y2=0.76
r207 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.825 $Y=0.675
+ $X2=3.825 $Y2=0.38
r208 46 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.66 $Y=0.76
+ $X2=3.825 $Y2=0.76
r209 46 47 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.66 $Y=0.76
+ $X2=2.97 $Y2=0.76
r210 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.805 $Y=0.675
+ $X2=2.97 $Y2=0.76
r211 44 99 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=0.425
+ $X2=2.805 $Y2=0.34
r212 44 45 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.805 $Y=0.425
+ $X2=2.805 $Y2=0.675
r213 43 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=0.34
+ $X2=1.945 $Y2=0.34
r214 42 99 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=0.34
+ $X2=2.805 $Y2=0.34
r215 42 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.64 $Y=0.34
+ $X2=2.11 $Y2=0.34
r216 38 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0.34
+ $X2=1.945 $Y2=0.34
r217 38 39 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.78 $Y=0.34
+ $X2=1.215 $Y2=0.34
r218 34 39 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.067 $Y=0.425
+ $X2=1.215 $Y2=0.34
r219 34 36 0.585988 $w=2.93e-07 $l=1.5e-08 $layer=LI1_cond $X=1.067 $Y=0.425
+ $X2=1.067 $Y2=0.44
r220 11 94 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=10.085
+ $Y=0.235 $X2=10.225 $Y2=0.42
r221 10 88 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.225
+ $Y=0.235 $X2=9.365 $Y2=0.42
r222 9 82 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.36
+ $Y=0.235 $X2=8.5 $Y2=0.42
r223 8 76 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.365
+ $Y=0.235 $X2=7.505 $Y2=0.42
r224 7 70 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.505
+ $Y=0.235 $X2=6.645 $Y2=0.42
r225 6 64 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.645
+ $Y=0.235 $X2=5.785 $Y2=0.42
r226 5 56 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=4.635
+ $Y=0.235 $X2=4.845 $Y2=0.38
r227 4 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.685
+ $Y=0.235 $X2=3.825 $Y2=0.38
r228 3 99 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.665
+ $Y=0.235 $X2=2.805 $Y2=0.38
r229 2 97 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.805
+ $Y=0.235 $X2=1.945 $Y2=0.38
r230 1 36 91 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=2 $X=0.96
+ $Y=0.235 $X2=1.085 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 41 45 47 51
+ 55 59 62 63 65 66 68 69 70 71 72 90 95 102 103 106 109 112 115
r152 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r153 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r154 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r155 107 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.92 $Y2=0
r156 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r157 103 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r158 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r159 100 115 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=9.94 $Y=0 $X2=9.8
+ $Y2=0
r160 100 102 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.94 $Y=0
+ $X2=10.32 $Y2=0
r161 99 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r162 99 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r163 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r164 96 112 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=9.07 $Y=0
+ $X2=8.932 $Y2=0
r165 96 98 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.07 $Y=0 $X2=9.36
+ $Y2=0
r166 95 115 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=9.66 $Y=0 $X2=9.8
+ $Y2=0
r167 95 98 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=9.66 $Y=0 $X2=9.36
+ $Y2=0
r168 94 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r169 94 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r170 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r171 91 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.17 $Y=0
+ $X2=8.005 $Y2=0
r172 91 93 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.17 $Y=0 $X2=8.4
+ $Y2=0
r173 90 112 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=8.795 $Y=0
+ $X2=8.932 $Y2=0
r174 90 93 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.4
+ $Y2=0
r175 89 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r176 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r177 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r178 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r179 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r180 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r181 79 80 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r182 76 80 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=3.12 $Y2=0
r183 75 79 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.12
+ $Y2=0
r184 75 76 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r185 72 89 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=6
+ $Y2=0
r186 72 86 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.04 $Y2=0
r187 70 88 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.05 $Y=0 $X2=6 $Y2=0
r188 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.05 $Y=0 $X2=6.215
+ $Y2=0
r189 68 85 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.185 $Y=0
+ $X2=5.04 $Y2=0
r190 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.185 $Y=0 $X2=5.35
+ $Y2=0
r191 67 88 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.515 $Y=0 $X2=6
+ $Y2=0
r192 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.515 $Y=0 $X2=5.35
+ $Y2=0
r193 65 82 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.17 $Y=0 $X2=4.08
+ $Y2=0
r194 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.17 $Y=0 $X2=4.335
+ $Y2=0
r195 64 85 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=5.04
+ $Y2=0
r196 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=4.335
+ $Y2=0
r197 62 79 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.15 $Y=0 $X2=3.12
+ $Y2=0
r198 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=0 $X2=3.315
+ $Y2=0
r199 61 82 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.48 $Y=0 $X2=4.08
+ $Y2=0
r200 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.48 $Y=0 $X2=3.315
+ $Y2=0
r201 57 115 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.8 $Y=0.085
+ $X2=9.8 $Y2=0
r202 57 59 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=9.8 $Y=0.085
+ $X2=9.8 $Y2=0.535
r203 53 112 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=8.932 $Y=0.085
+ $X2=8.932 $Y2=0
r204 53 55 18.8582 $w=2.73e-07 $l=4.5e-07 $layer=LI1_cond $X=8.932 $Y=0.085
+ $X2=8.932 $Y2=0.535
r205 49 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.005 $Y=0.085
+ $X2=8.005 $Y2=0
r206 49 51 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.005 $Y=0.085
+ $X2=8.005 $Y2=0.38
r207 48 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.24 $Y=0
+ $X2=7.075 $Y2=0
r208 47 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.84 $Y=0
+ $X2=8.005 $Y2=0
r209 47 48 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.84 $Y=0 $X2=7.24
+ $Y2=0
r210 43 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=0.085
+ $X2=7.075 $Y2=0
r211 43 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.075 $Y=0.085
+ $X2=7.075 $Y2=0.38
r212 42 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.38 $Y=0 $X2=6.215
+ $Y2=0
r213 41 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.91 $Y=0
+ $X2=7.075 $Y2=0
r214 41 42 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.91 $Y=0 $X2=6.38
+ $Y2=0
r215 37 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.215 $Y=0.085
+ $X2=6.215 $Y2=0
r216 37 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.215 $Y=0.085
+ $X2=6.215 $Y2=0.38
r217 33 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.35 $Y=0.085
+ $X2=5.35 $Y2=0
r218 33 35 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.35 $Y=0.085
+ $X2=5.35 $Y2=0.38
r219 29 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.335 $Y=0.085
+ $X2=4.335 $Y2=0
r220 29 31 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.335 $Y=0.085
+ $X2=4.335 $Y2=0.38
r221 25 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0
r222 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0.38
r223 8 59 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=9.655
+ $Y=0.235 $X2=9.795 $Y2=0.535
r224 7 55 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=8.795
+ $Y=0.235 $X2=8.935 $Y2=0.535
r225 6 51 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.795
+ $Y=0.235 $X2=8.005 $Y2=0.38
r226 5 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.935
+ $Y=0.235 $X2=7.075 $Y2=0.38
r227 4 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.075
+ $Y=0.235 $X2=6.215 $Y2=0.38
r228 3 35 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=5.135
+ $Y=0.235 $X2=5.35 $Y2=0.38
r229 2 31 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=4.115
+ $Y=0.235 $X2=4.335 $Y2=0.38
r230 1 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.235 $X2=3.315 $Y2=0.38
.ends

