* File: sky130_fd_sc_lp__nand4b_lp.pxi.spice
* Created: Wed Sep  2 10:06:24 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4B_LP%A_87_231# N_A_87_231#_M1010_d
+ N_A_87_231#_M1001_d N_A_87_231#_c_74_n N_A_87_231#_M1008_g N_A_87_231#_M1000_g
+ N_A_87_231#_c_77_n N_A_87_231#_c_83_n N_A_87_231#_c_78_n N_A_87_231#_c_79_n
+ N_A_87_231#_c_84_n N_A_87_231#_c_80_n N_A_87_231#_c_81_n
+ PM_SKY130_FD_SC_LP__NAND4B_LP%A_87_231#
x_PM_SKY130_FD_SC_LP__NAND4B_LP%B N_B_M1003_g N_B_M1009_g B N_B_c_148_n
+ N_B_c_149_n PM_SKY130_FD_SC_LP__NAND4B_LP%B
x_PM_SKY130_FD_SC_LP__NAND4B_LP%C N_C_M1005_g N_C_M1007_g N_C_c_192_n
+ N_C_c_197_n C C N_C_c_194_n PM_SKY130_FD_SC_LP__NAND4B_LP%C
x_PM_SKY130_FD_SC_LP__NAND4B_LP%D N_D_c_236_n N_D_M1006_g N_D_M1004_g
+ N_D_c_237_n N_D_c_238_n N_D_c_239_n N_D_c_244_n D D N_D_c_241_n
+ PM_SKY130_FD_SC_LP__NAND4B_LP%D
x_PM_SKY130_FD_SC_LP__NAND4B_LP%A_N N_A_N_c_283_n N_A_N_M1002_g N_A_N_M1001_g
+ N_A_N_c_284_n N_A_N_M1010_g N_A_N_c_285_n N_A_N_c_286_n N_A_N_c_287_n
+ N_A_N_c_292_n A_N A_N N_A_N_c_289_n PM_SKY130_FD_SC_LP__NAND4B_LP%A_N
x_PM_SKY130_FD_SC_LP__NAND4B_LP%VPWR N_VPWR_M1008_s N_VPWR_M1003_d
+ N_VPWR_M1004_d N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n N_VPWR_c_337_n
+ N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n VPWR N_VPWR_c_341_n
+ N_VPWR_c_333_n N_VPWR_c_343_n PM_SKY130_FD_SC_LP__NAND4B_LP%VPWR
x_PM_SKY130_FD_SC_LP__NAND4B_LP%Y N_Y_M1000_s N_Y_M1008_d N_Y_M1007_d
+ N_Y_c_386_n N_Y_c_387_n N_Y_c_388_n N_Y_c_389_n N_Y_c_390_n N_Y_c_391_n
+ N_Y_c_384_n N_Y_c_392_n Y Y PM_SKY130_FD_SC_LP__NAND4B_LP%Y
x_PM_SKY130_FD_SC_LP__NAND4B_LP%VGND N_VGND_M1006_d N_VGND_c_447_n VGND
+ N_VGND_c_448_n N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_451_n
+ PM_SKY130_FD_SC_LP__NAND4B_LP%VGND
cc_1 VNB N_A_87_231#_c_74_n 0.0471712f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.28
cc_2 VNB N_A_87_231#_M1008_g 0.0248587f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.545
cc_3 VNB N_A_87_231#_M1000_g 0.0231154f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.445
cc_4 VNB N_A_87_231#_c_77_n 0.0421495f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=0.91
cc_5 VNB N_A_87_231#_c_78_n 0.0220231f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=0.47
cc_6 VNB N_A_87_231#_c_79_n 0.0036521f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.91
cc_7 VNB N_A_87_231#_c_80_n 0.0314582f $X=-0.19 $Y=-0.245 $X2=3.027 $Y2=2.025
cc_8 VNB N_A_87_231#_c_81_n 0.0164212f $X=-0.19 $Y=-0.245 $X2=3.067 $Y2=0.91
cc_9 VNB N_B_M1009_g 0.0504199f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.28
cc_10 VNB N_B_c_148_n 0.0172997f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.445
cc_11 VNB N_B_c_149_n 0.0036033f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.445
cc_12 VNB N_C_M1005_g 0.0361987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C_c_192_n 0.0214367f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.825
cc_14 VNB C 0.00170402f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.445
cc_15 VNB N_C_c_194_n 0.016359f $X=-0.19 $Y=-0.245 $X2=3.027 $Y2=2.9
cc_16 VNB N_D_c_236_n 0.014806f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=0.235
cc_17 VNB N_D_c_237_n 0.0154323f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.445
cc_18 VNB N_D_c_238_n 0.016868f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=0.91
cc_19 VNB N_D_c_239_n 0.0218023f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.91
cc_20 VNB D 0.00171359f $X=-0.19 $Y=-0.245 $X2=3.027 $Y2=2.9
cc_21 VNB N_D_c_241_n 0.0165654f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=0.47
cc_22 VNB N_A_N_c_283_n 0.0145676f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=0.235
cc_23 VNB N_A_N_c_284_n 0.0172366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_N_c_285_n 0.0234538f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.91
cc_25 VNB N_A_N_c_286_n 0.0199726f $X=-0.19 $Y=-0.245 $X2=2.965 $Y2=2.9
cc_26 VNB N_A_N_c_287_n 0.0222717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A_N 0.00457311f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=0.47
cc_28 VNB N_A_N_c_289_n 0.0141921f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.91
cc_29 VNB N_VPWR_c_333_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.99
cc_30 VNB N_Y_c_384_n 0.0225304f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=0.47
cc_31 VNB Y 0.0527694f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.99
cc_32 VNB N_VGND_c_447_n 0.002833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_448_n 0.0602728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_449_n 0.0315757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_450_n 0.193212f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=0.825
cc_36 VNB N_VGND_c_451_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A_87_231#_M1008_g 0.0429968f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_38 VPB N_A_87_231#_c_83_n 0.0390561f $X=-0.19 $Y=1.655 $X2=2.965 $Y2=2.9
cc_39 VPB N_A_87_231#_c_84_n 0.0179524f $X=-0.19 $Y=1.655 $X2=2.965 $Y2=2.19
cc_40 VPB N_A_87_231#_c_80_n 0.0177864f $X=-0.19 $Y=1.655 $X2=3.027 $Y2=2.025
cc_41 VPB N_B_M1003_g 0.0318863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_B_c_148_n 0.00914787f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.445
cc_43 VPB N_B_c_149_n 0.00309836f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.445
cc_44 VPB N_C_M1007_g 0.0280974f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.28
cc_45 VPB N_C_c_192_n 0.00163736f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.825
cc_46 VPB N_C_c_197_n 0.0135841f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.445
cc_47 VPB C 7.45799e-19 $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.445
cc_48 VPB N_D_M1004_g 0.0283904f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_49 VPB N_D_c_239_n 0.00166642f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.91
cc_50 VPB N_D_c_244_n 0.0136829f $X=-0.19 $Y=1.655 $X2=3.027 $Y2=2.252
cc_51 VPB D 7.45264e-19 $X=-0.19 $Y=1.655 $X2=3.027 $Y2=2.9
cc_52 VPB N_A_N_M1001_g 0.0335899f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_53 VPB N_A_N_c_287_n 0.00170229f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_N_c_292_n 0.0139582f $X=-0.19 $Y=1.655 $X2=3.045 $Y2=0.825
cc_55 VPB A_N 0.00243168f $X=-0.19 $Y=1.655 $X2=3.045 $Y2=0.47
cc_56 VPB N_VPWR_c_334_n 0.0117329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_335_n 0.0334288f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.445
cc_58 VPB N_VPWR_c_336_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_337_n 0.00177638f $X=-0.19 $Y=1.655 $X2=3.027 $Y2=2.9
cc_60 VPB N_VPWR_c_338_n 0.010434f $X=-0.19 $Y=1.655 $X2=3.045 $Y2=0.47
cc_61 VPB N_VPWR_c_339_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.91
cc_62 VPB N_VPWR_c_340_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_341_n 0.0220676f $X=-0.19 $Y=1.655 $X2=3.067 $Y2=0.91
cc_64 VPB N_VPWR_c_333_n 0.0527973f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=0.99
cc_65 VPB N_VPWR_c_343_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_Y_c_386_n 0.00271393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_Y_c_387_n 0.00779619f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.825
cc_68 VPB N_Y_c_388_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_Y_c_389_n 0.00770712f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.91
cc_70 VPB N_Y_c_390_n 0.00906025f $X=-0.19 $Y=1.655 $X2=3.027 $Y2=2.9
cc_71 VPB N_Y_c_391_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_Y_c_392_n 0.00254917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB Y 0.0152712f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.99
cc_74 N_A_87_231#_M1008_g N_B_M1003_g 0.0194569f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_75 N_A_87_231#_c_74_n N_B_M1009_g 0.0107575f $X=0.56 $Y=1.28 $X2=0 $Y2=0
cc_76 N_A_87_231#_M1000_g N_B_M1009_g 0.0585636f $X=0.79 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A_87_231#_c_77_n N_B_M1009_g 0.0128841f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_78 N_A_87_231#_c_79_n N_B_M1009_g 0.00115306f $X=0.7 $Y=0.91 $X2=0 $Y2=0
cc_79 N_A_87_231#_M1008_g N_B_c_148_n 0.0181444f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_80 N_A_87_231#_c_77_n N_B_c_148_n 0.00367189f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_81 N_A_87_231#_c_74_n N_B_c_149_n 0.00119725f $X=0.56 $Y=1.28 $X2=0 $Y2=0
cc_82 N_A_87_231#_M1008_g N_B_c_149_n 0.0123212f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_83 N_A_87_231#_c_77_n N_B_c_149_n 0.0137011f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_84 N_A_87_231#_c_79_n N_B_c_149_n 0.0133077f $X=0.7 $Y=0.91 $X2=0 $Y2=0
cc_85 N_A_87_231#_c_77_n N_C_M1005_g 0.0119252f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_86 N_A_87_231#_c_77_n C 0.0245014f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_87 N_A_87_231#_c_77_n N_C_c_194_n 0.00122373f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_88 N_A_87_231#_c_84_n N_D_M1004_g 2.87643e-19 $X=2.965 $Y=2.19 $X2=0 $Y2=0
cc_89 N_A_87_231#_c_77_n N_D_c_237_n 0.00874789f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_90 N_A_87_231#_c_77_n N_D_c_238_n 0.0070824f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_91 N_A_87_231#_c_77_n D 0.0245051f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_92 N_A_87_231#_c_77_n N_D_c_241_n 0.00123044f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_93 N_A_87_231#_c_78_n N_A_N_c_283_n 0.00150158f $X=3.045 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_87_231#_c_83_n N_A_N_M1001_g 0.0150161f $X=2.965 $Y=2.9 $X2=0 $Y2=0
cc_95 N_A_87_231#_c_84_n N_A_N_M1001_g 0.00480265f $X=2.965 $Y=2.19 $X2=0 $Y2=0
cc_96 N_A_87_231#_c_80_n N_A_N_M1001_g 0.00427061f $X=3.027 $Y=2.025 $X2=0 $Y2=0
cc_97 N_A_87_231#_c_78_n N_A_N_c_284_n 0.00990318f $X=3.045 $Y=0.47 $X2=0 $Y2=0
cc_98 N_A_87_231#_c_77_n N_A_N_c_285_n 0.0184498f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_99 N_A_87_231#_c_78_n N_A_N_c_285_n 0.0063278f $X=3.045 $Y=0.47 $X2=0 $Y2=0
cc_100 N_A_87_231#_c_81_n N_A_N_c_285_n 0.00144114f $X=3.067 $Y=0.91 $X2=0 $Y2=0
cc_101 N_A_87_231#_c_77_n N_A_N_c_286_n 0.00806361f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_102 N_A_87_231#_c_80_n N_A_N_c_286_n 0.00362326f $X=3.027 $Y=2.025 $X2=0
+ $Y2=0
cc_103 N_A_87_231#_c_84_n N_A_N_c_292_n 6.14058e-19 $X=2.965 $Y=2.19 $X2=0 $Y2=0
cc_104 N_A_87_231#_c_77_n A_N 0.0266762f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_105 N_A_87_231#_c_84_n A_N 0.00867382f $X=2.965 $Y=2.19 $X2=0 $Y2=0
cc_106 N_A_87_231#_c_80_n A_N 0.0486831f $X=3.027 $Y=2.025 $X2=0 $Y2=0
cc_107 N_A_87_231#_c_81_n A_N 0.00204652f $X=3.067 $Y=0.91 $X2=0 $Y2=0
cc_108 N_A_87_231#_c_77_n N_A_N_c_289_n 4.94304e-19 $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_109 N_A_87_231#_c_80_n N_A_N_c_289_n 0.0148853f $X=3.027 $Y=2.025 $X2=0 $Y2=0
cc_110 N_A_87_231#_M1008_g N_VPWR_c_335_n 0.0192403f $X=0.56 $Y=2.545 $X2=0
+ $Y2=0
cc_111 N_A_87_231#_M1008_g N_VPWR_c_336_n 0.00769046f $X=0.56 $Y=2.545 $X2=0
+ $Y2=0
cc_112 N_A_87_231#_M1008_g N_VPWR_c_337_n 8.49223e-19 $X=0.56 $Y=2.545 $X2=0
+ $Y2=0
cc_113 N_A_87_231#_c_84_n N_VPWR_c_338_n 0.0650754f $X=2.965 $Y=2.19 $X2=0 $Y2=0
cc_114 N_A_87_231#_c_83_n N_VPWR_c_341_n 0.0304602f $X=2.965 $Y=2.9 $X2=0 $Y2=0
cc_115 N_A_87_231#_M1008_g N_VPWR_c_333_n 0.0134474f $X=0.56 $Y=2.545 $X2=0
+ $Y2=0
cc_116 N_A_87_231#_c_83_n N_VPWR_c_333_n 0.0174175f $X=2.965 $Y=2.9 $X2=0 $Y2=0
cc_117 N_A_87_231#_M1008_g N_Y_c_386_n 0.024414f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_118 N_A_87_231#_M1008_g N_Y_c_388_n 0.0187085f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_119 N_A_87_231#_c_74_n N_Y_c_384_n 0.0043208f $X=0.56 $Y=1.28 $X2=0 $Y2=0
cc_120 N_A_87_231#_M1000_g N_Y_c_384_n 0.00752285f $X=0.79 $Y=0.445 $X2=0 $Y2=0
cc_121 N_A_87_231#_c_79_n N_Y_c_384_n 0.0126596f $X=0.7 $Y=0.91 $X2=0 $Y2=0
cc_122 N_A_87_231#_M1008_g N_Y_c_392_n 0.00489696f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_123 N_A_87_231#_c_74_n Y 0.0353093f $X=0.56 $Y=1.28 $X2=0 $Y2=0
cc_124 N_A_87_231#_M1000_g Y 0.00512192f $X=0.79 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_87_231#_c_79_n Y 0.0243167f $X=0.7 $Y=0.91 $X2=0 $Y2=0
cc_126 N_A_87_231#_c_77_n N_VGND_c_447_n 0.0222143f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_127 N_A_87_231#_M1000_g N_VGND_c_448_n 0.0054778f $X=0.79 $Y=0.445 $X2=0
+ $Y2=0
cc_128 N_A_87_231#_c_78_n N_VGND_c_449_n 0.0197885f $X=3.045 $Y=0.47 $X2=0 $Y2=0
cc_129 N_A_87_231#_M1010_d N_VGND_c_450_n 0.00232985f $X=2.905 $Y=0.235 $X2=0
+ $Y2=0
cc_130 N_A_87_231#_M1000_g N_VGND_c_450_n 0.00742906f $X=0.79 $Y=0.445 $X2=0
+ $Y2=0
cc_131 N_A_87_231#_c_77_n N_VGND_c_450_n 0.0543174f $X=2.88 $Y=0.91 $X2=0 $Y2=0
cc_132 N_A_87_231#_c_78_n N_VGND_c_450_n 0.0125808f $X=3.045 $Y=0.47 $X2=0 $Y2=0
cc_133 N_A_87_231#_c_79_n N_VGND_c_450_n 0.00397468f $X=0.7 $Y=0.91 $X2=0 $Y2=0
cc_134 N_A_87_231#_c_81_n N_VGND_c_450_n 0.00179786f $X=3.067 $Y=0.91 $X2=0
+ $Y2=0
cc_135 N_B_M1009_g N_C_M1005_g 0.0615638f $X=1.18 $Y=0.445 $X2=0 $Y2=0
cc_136 N_B_M1003_g N_C_M1007_g 0.0299962f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_137 N_B_c_148_n N_C_c_192_n 0.0191671f $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_138 N_B_c_149_n N_C_c_192_n 0.0011377f $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_139 N_B_M1003_g N_C_c_197_n 0.0035718f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_140 N_B_M1003_g C 4.35377e-19 $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_141 N_B_M1009_g C 0.00183384f $X=1.18 $Y=0.445 $X2=0 $Y2=0
cc_142 N_B_c_148_n C 4.1366e-19 $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_143 N_B_c_149_n C 0.0219784f $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_144 N_B_M1009_g N_C_c_194_n 0.0191671f $X=1.18 $Y=0.445 $X2=0 $Y2=0
cc_145 N_B_M1003_g N_VPWR_c_335_n 8.6579e-19 $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_146 N_B_M1003_g N_VPWR_c_336_n 0.00769046f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_147 N_B_M1003_g N_VPWR_c_337_n 0.0163548f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_148 N_B_M1003_g N_VPWR_c_333_n 0.0134474f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_149 N_B_c_149_n N_Y_c_386_n 0.00371935f $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_150 N_B_M1003_g N_Y_c_388_n 0.0155966f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_151 N_B_M1003_g N_Y_c_389_n 0.0184281f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_152 N_B_c_148_n N_Y_c_389_n 9.97824e-19 $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_153 N_B_c_149_n N_Y_c_389_n 0.0142612f $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_154 N_B_M1003_g N_Y_c_391_n 8.93705e-19 $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_155 N_B_M1009_g N_Y_c_384_n 0.00187941f $X=1.18 $Y=0.445 $X2=0 $Y2=0
cc_156 N_B_M1003_g N_Y_c_392_n 0.00317911f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_157 N_B_c_148_n N_Y_c_392_n 9.27233e-19 $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_158 N_B_c_149_n N_Y_c_392_n 0.02743f $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_159 N_B_c_149_n Y 0.0199626f $X=1.09 $Y=1.615 $X2=0 $Y2=0
cc_160 N_B_M1009_g N_VGND_c_448_n 0.00585385f $X=1.18 $Y=0.445 $X2=0 $Y2=0
cc_161 N_B_M1009_g N_VGND_c_450_n 0.00633367f $X=1.18 $Y=0.445 $X2=0 $Y2=0
cc_162 N_C_M1005_g N_D_c_236_n 0.0434803f $X=1.57 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_163 N_C_M1007_g N_D_M1004_g 0.0171479f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_164 N_C_M1005_g N_D_c_238_n 0.0109452f $X=1.57 $Y=0.445 $X2=0 $Y2=0
cc_165 N_C_c_192_n N_D_c_239_n 0.0135694f $X=1.63 $Y=1.68 $X2=0 $Y2=0
cc_166 N_C_c_197_n N_D_c_244_n 0.0135694f $X=1.63 $Y=1.845 $X2=0 $Y2=0
cc_167 C D 0.0423335f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_168 N_C_c_194_n D 0.00232658f $X=1.63 $Y=1.34 $X2=0 $Y2=0
cc_169 C N_D_c_241_n 0.00232658f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_170 N_C_c_194_n N_D_c_241_n 0.0135694f $X=1.63 $Y=1.34 $X2=0 $Y2=0
cc_171 N_C_M1007_g N_VPWR_c_337_n 0.0163548f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_172 N_C_M1007_g N_VPWR_c_338_n 9.45181e-19 $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_173 N_C_M1007_g N_VPWR_c_339_n 0.00769046f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_174 N_C_M1007_g N_VPWR_c_333_n 0.0134474f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_175 N_C_M1007_g N_Y_c_388_n 8.93705e-19 $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_176 N_C_M1007_g N_Y_c_389_n 0.0178513f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_177 C N_Y_c_389_n 0.0185305f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_178 N_C_M1007_g N_Y_c_390_n 9.81754e-19 $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_179 N_C_c_197_n N_Y_c_390_n 3.80871e-19 $X=1.63 $Y=1.845 $X2=0 $Y2=0
cc_180 C N_Y_c_390_n 0.00619639f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_181 N_C_M1007_g N_Y_c_391_n 0.0155966f $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_182 N_C_M1007_g N_Y_c_392_n 2.77272e-19 $X=1.62 $Y=2.545 $X2=0 $Y2=0
cc_183 N_C_M1005_g N_VGND_c_447_n 0.00312012f $X=1.57 $Y=0.445 $X2=0 $Y2=0
cc_184 N_C_M1005_g N_VGND_c_448_n 0.00585385f $X=1.57 $Y=0.445 $X2=0 $Y2=0
cc_185 N_C_M1005_g N_VGND_c_450_n 0.00633367f $X=1.57 $Y=0.445 $X2=0 $Y2=0
cc_186 N_D_c_236_n N_A_N_c_283_n 0.0132973f $X=1.96 $Y=0.73 $X2=-0.19 $Y2=-0.245
cc_187 N_D_M1004_g N_A_N_M1001_g 0.015445f $X=2.15 $Y=2.545 $X2=0 $Y2=0
cc_188 N_D_c_237_n N_A_N_c_285_n 0.00941174f $X=2.08 $Y=0.805 $X2=0 $Y2=0
cc_189 N_D_c_238_n N_A_N_c_286_n 0.00923257f $X=2.17 $Y=1.175 $X2=0 $Y2=0
cc_190 N_D_c_239_n N_A_N_c_287_n 0.0117733f $X=2.17 $Y=1.68 $X2=0 $Y2=0
cc_191 N_D_c_244_n N_A_N_c_292_n 0.0117733f $X=2.17 $Y=1.845 $X2=0 $Y2=0
cc_192 D A_N 0.0492677f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_193 N_D_c_241_n A_N 0.00411803f $X=2.17 $Y=1.34 $X2=0 $Y2=0
cc_194 D N_A_N_c_289_n 7.73334e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_195 N_D_c_241_n N_A_N_c_289_n 0.0117733f $X=2.17 $Y=1.34 $X2=0 $Y2=0
cc_196 N_D_M1004_g N_VPWR_c_337_n 8.49223e-19 $X=2.15 $Y=2.545 $X2=0 $Y2=0
cc_197 N_D_M1004_g N_VPWR_c_338_n 0.0225513f $X=2.15 $Y=2.545 $X2=0 $Y2=0
cc_198 N_D_c_244_n N_VPWR_c_338_n 4.586e-19 $X=2.17 $Y=1.845 $X2=0 $Y2=0
cc_199 D N_VPWR_c_338_n 0.00696838f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_200 N_D_M1004_g N_VPWR_c_339_n 0.00769046f $X=2.15 $Y=2.545 $X2=0 $Y2=0
cc_201 N_D_M1004_g N_VPWR_c_333_n 0.0134474f $X=2.15 $Y=2.545 $X2=0 $Y2=0
cc_202 N_D_M1004_g N_Y_c_390_n 0.00354188f $X=2.15 $Y=2.545 $X2=0 $Y2=0
cc_203 D N_Y_c_390_n 0.00363823f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_204 N_D_M1004_g N_Y_c_391_n 0.0150096f $X=2.15 $Y=2.545 $X2=0 $Y2=0
cc_205 N_D_c_236_n N_VGND_c_447_n 0.0127111f $X=1.96 $Y=0.73 $X2=0 $Y2=0
cc_206 N_D_c_237_n N_VGND_c_447_n 0.00342512f $X=2.08 $Y=0.805 $X2=0 $Y2=0
cc_207 N_D_c_236_n N_VGND_c_448_n 0.00486043f $X=1.96 $Y=0.73 $X2=0 $Y2=0
cc_208 N_D_c_236_n N_VGND_c_450_n 0.00450668f $X=1.96 $Y=0.73 $X2=0 $Y2=0
cc_209 N_A_N_M1001_g N_VPWR_c_338_n 0.0217145f $X=2.7 $Y=2.545 $X2=0 $Y2=0
cc_210 A_N N_VPWR_c_338_n 0.00472567f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_211 N_A_N_M1001_g N_VPWR_c_341_n 0.00840515f $X=2.7 $Y=2.545 $X2=0 $Y2=0
cc_212 N_A_N_M1001_g N_VPWR_c_333_n 0.0153885f $X=2.7 $Y=2.545 $X2=0 $Y2=0
cc_213 N_A_N_M1001_g N_Y_c_391_n 2.18111e-19 $X=2.7 $Y=2.545 $X2=0 $Y2=0
cc_214 N_A_N_c_283_n N_VGND_c_447_n 0.00516266f $X=2.47 $Y=0.73 $X2=0 $Y2=0
cc_215 N_A_N_c_283_n N_VGND_c_449_n 0.00585385f $X=2.47 $Y=0.73 $X2=0 $Y2=0
cc_216 N_A_N_c_284_n N_VGND_c_449_n 0.00549284f $X=2.83 $Y=0.73 $X2=0 $Y2=0
cc_217 N_A_N_c_285_n N_VGND_c_449_n 6.21075e-19 $X=2.83 $Y=0.805 $X2=0 $Y2=0
cc_218 N_A_N_c_283_n N_VGND_c_450_n 0.00638707f $X=2.47 $Y=0.73 $X2=0 $Y2=0
cc_219 N_A_N_c_284_n N_VGND_c_450_n 0.00715351f $X=2.83 $Y=0.73 $X2=0 $Y2=0
cc_220 N_A_N_c_285_n N_VGND_c_450_n 8.18184e-19 $X=2.83 $Y=0.805 $X2=0 $Y2=0
cc_221 N_VPWR_M1008_s N_Y_c_386_n 2.39543e-19 $X=0.15 $Y=2.045 $X2=0 $Y2=0
cc_222 N_VPWR_c_335_n N_Y_c_386_n 0.00346358f $X=0.295 $Y=2.475 $X2=0 $Y2=0
cc_223 N_VPWR_M1008_s N_Y_c_387_n 0.00281819f $X=0.15 $Y=2.045 $X2=0 $Y2=0
cc_224 N_VPWR_c_335_n N_Y_c_387_n 0.019414f $X=0.295 $Y=2.475 $X2=0 $Y2=0
cc_225 N_VPWR_c_335_n N_Y_c_388_n 0.0497475f $X=0.295 $Y=2.475 $X2=0 $Y2=0
cc_226 N_VPWR_c_336_n N_Y_c_388_n 0.021949f $X=1.19 $Y=3.33 $X2=0 $Y2=0
cc_227 N_VPWR_c_337_n N_Y_c_388_n 0.0454646f $X=1.355 $Y=2.54 $X2=0 $Y2=0
cc_228 N_VPWR_c_333_n N_Y_c_388_n 0.0124703f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_229 N_VPWR_M1003_d N_Y_c_389_n 0.00180746f $X=1.215 $Y=2.045 $X2=0 $Y2=0
cc_230 N_VPWR_c_337_n N_Y_c_389_n 0.0163515f $X=1.355 $Y=2.54 $X2=0 $Y2=0
cc_231 N_VPWR_c_338_n N_Y_c_390_n 0.0119061f $X=2.415 $Y=2.19 $X2=0 $Y2=0
cc_232 N_VPWR_c_337_n N_Y_c_391_n 0.0454646f $X=1.355 $Y=2.54 $X2=0 $Y2=0
cc_233 N_VPWR_c_338_n N_Y_c_391_n 0.0572919f $X=2.415 $Y=2.19 $X2=0 $Y2=0
cc_234 N_VPWR_c_339_n N_Y_c_391_n 0.021949f $X=2.25 $Y=3.33 $X2=0 $Y2=0
cc_235 N_VPWR_c_333_n N_Y_c_391_n 0.0124703f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_236 N_Y_c_384_n N_VGND_c_448_n 0.027436f $X=0.24 $Y=0.645 $X2=0 $Y2=0
cc_237 N_Y_M1000_s N_VGND_c_450_n 0.0023218f $X=0.43 $Y=0.235 $X2=0 $Y2=0
cc_238 N_Y_c_384_n N_VGND_c_450_n 0.022061f $X=0.24 $Y=0.645 $X2=0 $Y2=0
cc_239 A_173_47# N_VGND_c_450_n 0.00346804f $X=0.865 $Y=0.235 $X2=3.12 $Y2=0
cc_240 A_251_47# N_VGND_c_450_n 0.00346804f $X=1.255 $Y=0.235 $X2=3.12 $Y2=0
cc_241 A_329_47# N_VGND_c_450_n 0.00346804f $X=1.645 $Y=0.235 $X2=3.12 $Y2=0
cc_242 N_VGND_c_450_n A_509_47# 0.00303453f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
