* File: sky130_fd_sc_lp__lsbuf_lp.pxi.spice
* Created: Wed Sep  2 09:58:57 2020
* 
x_PM_SKY130_FD_SC_LP__LSBUF_LP%VGND N_VGND_M1011_s N_VGND_M1005_d N_VGND_M1000_s
+ N_VGND_M1011_b N_VGND_c_17_p N_VGND_c_21_p N_VGND_c_7_p N_VGND_c_18_p VGND
+ N_VGND_c_71_p N_VGND_c_12_p N_VGND_c_13_p PM_SKY130_FD_SC_LP__LSBUF_LP%VGND
x_PM_SKY130_FD_SC_LP__LSBUF_LP%VPB N_VPB_M1009_b VPB VPB VPB VPB VPB VPB
+ PM_SKY130_FD_SC_LP__LSBUF_LP%VPB
x_PM_SKY130_FD_SC_LP__LSBUF_LP%DESTVPB N_DESTVPB_M1014_b DESTVPB DESTVPB DESTVPB
+ DESTVPB DESTVPB DESTVPB PM_SKY130_FD_SC_LP__LSBUF_LP%DESTVPB
x_PM_SKY130_FD_SC_LP__LSBUF_LP%A_246_987# N_A_246_987#_M1002_d
+ N_A_246_987#_M1012_d N_A_246_987#_M1014_g N_A_246_987#_M1015_g
+ N_A_246_987#_c_171_n N_A_246_987#_c_172_n N_A_246_987#_c_173_n
+ N_A_246_987#_c_159_n N_A_246_987#_c_162_n N_A_246_987#_c_163_n
+ N_A_246_987#_c_175_n N_A_246_987#_c_164_n N_A_246_987#_c_168_n
+ PM_SKY130_FD_SC_LP__LSBUF_LP%A_246_987#
x_PM_SKY130_FD_SC_LP__LSBUF_LP%A N_A_M1009_g N_A_c_243_n N_A_M1011_g N_A_M1010_g
+ N_A_M1001_g N_A_M1008_g N_A_M1005_g N_A_c_258_n N_A_c_260_n N_A_c_264_n A
+ N_A_c_267_n N_A_c_269_n N_A_c_273_n PM_SKY130_FD_SC_LP__LSBUF_LP%A
x_PM_SKY130_FD_SC_LP__LSBUF_LP%A_278_47# N_A_278_47#_M1008_d N_A_278_47#_M1001_d
+ N_A_278_47#_c_306_n N_A_278_47#_M1007_g N_A_278_47#_c_309_n
+ N_A_278_47#_c_310_n N_A_278_47#_c_311_n N_A_278_47#_M1002_g
+ N_A_278_47#_c_325_n N_A_278_47#_c_315_n N_A_278_47#_c_316_n
+ N_A_278_47#_c_319_n N_A_278_47#_c_327_n N_A_278_47#_c_324_n
+ PM_SKY130_FD_SC_LP__LSBUF_LP%A_278_47#
x_PM_SKY130_FD_SC_LP__LSBUF_LP%A_193_718# N_A_193_718#_M1010_s
+ N_A_193_718#_M1014_s N_A_193_718#_c_396_n N_A_193_718#_M1006_g
+ N_A_193_718#_c_397_n N_A_193_718#_M1012_g N_A_193_718#_c_398_n
+ N_A_193_718#_c_373_n N_A_193_718#_c_374_n N_A_193_718#_M1000_g
+ N_A_193_718#_M1004_g N_A_193_718#_c_379_n N_A_193_718#_M1013_g
+ N_A_193_718#_M1003_g N_A_193_718#_c_384_n N_A_193_718#_c_385_n
+ N_A_193_718#_c_386_n N_A_193_718#_c_387_n N_A_193_718#_c_408_n
+ N_A_193_718#_c_391_n N_A_193_718#_c_393_n N_A_193_718#_c_394_n
+ N_A_193_718#_c_410_n N_A_193_718#_c_395_n N_A_193_718#_c_413_n
+ PM_SKY130_FD_SC_LP__LSBUF_LP%A_193_718#
x_PM_SKY130_FD_SC_LP__LSBUF_LP%VPWR N_VPWR_M1009_s N_VPWR_c_490_n VPWR
+ N_VPWR_c_492_n N_VPWR_c_494_n N_VPWR_c_489_n N_VPWR_c_499_n
+ PM_SKY130_FD_SC_LP__LSBUF_LP%VPWR
x_PM_SKY130_FD_SC_LP__LSBUF_LP%DESTPWR N_DESTPWR_M1015_d N_DESTPWR_M1004_s
+ N_DESTPWR_c_517_n N_DESTPWR_c_518_n N_DESTPWR_c_519_n N_DESTPWR_c_521_n
+ DESTPWR N_DESTPWR_c_522_n N_DESTPWR_c_523_n N_DESTPWR_c_516_n
+ N_DESTPWR_c_528_n PM_SKY130_FD_SC_LP__LSBUF_LP%DESTPWR
x_PM_SKY130_FD_SC_LP__LSBUF_LP%X N_X_M1013_d N_X_M1003_d X X X X X X N_X_c_572_n
+ PM_SKY130_FD_SC_LP__LSBUF_LP%X
cc_1 N_VGND_M1011_b VPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_2 N_VGND_M1011_b VPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=4.475 $Y2=0.47
cc_3 N_VGND_M1011_b DESTVPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_4 N_VGND_M1011_b DESTVPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=4.475 $Y2=0.47
cc_5 N_VGND_M1000_s N_A_246_987#_c_159_n 8.76384e-19 $X=3.125 $Y=3.59 $X2=0
+ $Y2=0
cc_6 N_VGND_M1011_b N_A_246_987#_c_159_n 0.0156489f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_7 N_VGND_c_7_p N_A_246_987#_c_159_n 0.00493592f $X=3.27 $Y=3.715 $X2=0 $Y2=0
cc_8 N_VGND_M1011_b N_A_246_987#_c_162_n 0.00411745f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_9 N_VGND_M1011_b N_A_246_987#_c_163_n 0.00736044f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_10 N_VGND_M1011_b N_A_246_987#_c_164_n 0.00939378f $X=-0.025 $Y=-0.245
+ $X2=4.56 $Y2=0.925
cc_11 N_VGND_c_7_p N_A_246_987#_c_164_n 0.0546974f $X=3.27 $Y=3.715 $X2=4.56
+ $Y2=0.925
cc_12 N_VGND_c_12_p N_A_246_987#_c_164_n 0.0305519f $X=3.12 $Y=3.33 $X2=4.56
+ $Y2=0.925
cc_13 N_VGND_c_13_p N_A_246_987#_c_164_n 0.0165209f $X=4.56 $Y=3.33 $X2=4.56
+ $Y2=0.925
cc_14 N_VGND_M1011_b N_A_246_987#_c_168_n 0.0169579f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_15 N_VGND_M1011_b N_A_M1009_g 0.00622578f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_16 N_VGND_M1011_b N_A_c_243_n 0.0227707f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_17 N_VGND_c_17_p N_A_c_243_n 0.00857607f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_18 N_VGND_c_18_p N_A_c_243_n 0.00322089f $X=1.715 $Y=3.33 $X2=0 $Y2=0
cc_19 N_VGND_c_13_p N_A_c_243_n 0.00381775f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_20 N_VGND_M1011_b N_A_M1010_g 0.0392728f $X=-0.025 $Y=-0.245 $X2=0.155
+ $Y2=0.84
cc_21 N_VGND_c_21_p N_A_M1010_g 0.00388479f $X=1.88 $Y=3.715 $X2=0.155 $Y2=0.84
cc_22 N_VGND_c_18_p N_A_M1010_g 0.012665f $X=1.715 $Y=3.33 $X2=0.155 $Y2=0.84
cc_23 N_VGND_c_13_p N_A_M1010_g 0.0142323f $X=4.56 $Y=3.33 $X2=0.155 $Y2=0.84
cc_24 N_VGND_M1011_b N_A_M1001_g 0.00537455f $X=-0.025 $Y=-0.245 $X2=4.475
+ $Y2=1.21
cc_25 N_VGND_M1011_b N_A_M1008_g 0.0125692f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_26 N_VGND_c_17_p N_A_M1008_g 3.66739e-19 $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_27 N_VGND_M1011_b N_A_M1005_g 0.0357211f $X=-0.025 $Y=-0.245 $X2=0.24
+ $Y2=0.525
cc_28 N_VGND_c_21_p N_A_M1005_g 0.0232744f $X=1.88 $Y=3.715 $X2=0.24 $Y2=0.525
cc_29 N_VGND_c_18_p N_A_M1005_g 0.011296f $X=1.715 $Y=3.33 $X2=0.24 $Y2=0.525
cc_30 N_VGND_c_13_p N_A_M1005_g 0.0101853f $X=4.56 $Y=3.33 $X2=0.24 $Y2=0.525
cc_31 N_VGND_M1011_b N_A_c_258_n 0.00200096f $X=-0.025 $Y=-0.245 $X2=0.24
+ $Y2=0.925
cc_32 N_VGND_c_17_p N_A_c_258_n 0.0222632f $X=0.74 $Y=2.44 $X2=0.24 $Y2=0.925
cc_33 N_VGND_M1011_b N_A_c_260_n 0.00392808f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_34 N_VGND_c_17_p N_A_c_260_n 0.0265164f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_35 N_VGND_c_18_p N_A_c_260_n 0.012059f $X=1.715 $Y=3.33 $X2=0 $Y2=0
cc_36 N_VGND_c_13_p N_A_c_260_n 0.00653588f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_37 N_VGND_M1011_b N_A_c_264_n 0.00325622f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_38 N_VGND_c_18_p N_A_c_264_n 0.0419863f $X=1.715 $Y=3.33 $X2=0 $Y2=0
cc_39 N_VGND_c_13_p N_A_c_264_n 0.0222748f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_40 N_VGND_M1011_b N_A_c_267_n 0.0674831f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_41 N_VGND_c_17_p N_A_c_267_n 0.00213349f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_42 N_VGND_M1011_b N_A_c_269_n 0.062954f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_43 N_VGND_c_17_p N_A_c_269_n 0.00526872f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_44 N_VGND_c_18_p N_A_c_269_n 0.00346729f $X=1.715 $Y=3.33 $X2=0 $Y2=0
cc_45 N_VGND_c_13_p N_A_c_269_n 0.00867339f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_46 N_VGND_M1011_b N_A_c_273_n 0.0344679f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_47 N_VGND_c_17_p N_A_c_273_n 0.0262117f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_48 N_VGND_M1011_b N_A_278_47#_c_306_n 0.0153045f $X=-0.025 $Y=-0.245
+ $X2=-0.025 $Y2=-0.19
cc_49 N_VGND_c_21_p N_A_278_47#_c_306_n 0.00216224f $X=1.88 $Y=3.715 $X2=-0.025
+ $Y2=-0.19
cc_50 N_VGND_c_13_p N_A_278_47#_c_306_n 0.00937715f $X=4.56 $Y=3.33 $X2=-0.025
+ $Y2=-0.19
cc_51 N_VGND_M1011_b N_A_278_47#_c_309_n 0.00847207f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=0.84
cc_52 N_VGND_M1011_b N_A_278_47#_c_310_n 0.0114697f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=1.21
cc_53 N_VGND_M1011_b N_A_278_47#_c_311_n 0.0180803f $X=-0.025 $Y=-0.245
+ $X2=4.475 $Y2=0.47
cc_54 N_VGND_c_7_p N_A_278_47#_c_311_n 0.00287368f $X=3.27 $Y=3.715 $X2=4.475
+ $Y2=0.47
cc_55 N_VGND_c_12_p N_A_278_47#_c_311_n 5.83419e-19 $X=3.12 $Y=3.33 $X2=4.475
+ $Y2=0.47
cc_56 N_VGND_c_13_p N_A_278_47#_c_311_n 0.010645f $X=4.56 $Y=3.33 $X2=4.475
+ $Y2=0.47
cc_57 N_VGND_M1011_b N_A_278_47#_c_315_n 0.0382462f $X=-0.025 $Y=-0.245 $X2=0.24
+ $Y2=0.525
cc_58 N_VGND_M1011_b N_A_278_47#_c_316_n 0.0378754f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_59 N_VGND_c_18_p N_A_278_47#_c_316_n 0.001325f $X=1.715 $Y=3.33 $X2=0 $Y2=0
cc_60 N_VGND_c_13_p N_A_278_47#_c_316_n 0.00908544f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_61 N_VGND_M1011_b N_A_278_47#_c_319_n 0.0443455f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_62 N_VGND_c_21_p N_A_278_47#_c_319_n 0.0444661f $X=1.88 $Y=3.715 $X2=0 $Y2=0
cc_63 N_VGND_c_18_p N_A_278_47#_c_319_n 0.0123326f $X=1.715 $Y=3.33 $X2=0 $Y2=0
cc_64 N_VGND_c_12_p N_A_278_47#_c_319_n 0.0121875f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_65 N_VGND_c_13_p N_A_278_47#_c_319_n 0.0503784f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_66 N_VGND_M1011_b N_A_278_47#_c_324_n 0.0436885f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_67 N_VGND_M1011_b N_A_193_718#_c_373_n 0.00977309f $X=-0.025 $Y=-0.245
+ $X2=4.475 $Y2=1.21
cc_68 N_VGND_M1011_b N_A_193_718#_c_374_n 0.0134026f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_69 N_VGND_M1011_b N_A_193_718#_M1000_g 0.0402979f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_70 N_VGND_c_7_p N_A_193_718#_M1000_g 0.0178969f $X=3.27 $Y=3.715 $X2=0 $Y2=0
cc_71 N_VGND_c_71_p N_A_193_718#_M1000_g 0.00465098f $X=4.41 $Y=3.33 $X2=0 $Y2=0
cc_72 N_VGND_c_13_p N_A_193_718#_M1000_g 0.00805442f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_73 N_VGND_M1011_b N_A_193_718#_c_379_n 0.00251633f $X=-0.025 $Y=-0.245
+ $X2=0.24 $Y2=0.925
cc_74 N_VGND_M1011_b N_A_193_718#_M1013_g 0.0475006f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_75 N_VGND_c_7_p N_A_193_718#_M1013_g 0.0027764f $X=3.27 $Y=3.715 $X2=0 $Y2=0
cc_76 N_VGND_c_71_p N_A_193_718#_M1013_g 0.00525141f $X=4.41 $Y=3.33 $X2=0 $Y2=0
cc_77 N_VGND_c_13_p N_A_193_718#_M1013_g 0.0107926f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_78 N_VGND_M1011_b N_A_193_718#_c_384_n 0.00608676f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_79 N_VGND_M1011_b N_A_193_718#_c_385_n 7.95968e-19 $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_80 N_VGND_M1011_b N_A_193_718#_c_386_n 0.00222291f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_81 N_VGND_M1011_b N_A_193_718#_c_387_n 0.0653551f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_82 N_VGND_c_21_p N_A_193_718#_c_387_n 0.0143416f $X=1.88 $Y=3.715 $X2=0 $Y2=0
cc_83 N_VGND_c_18_p N_A_193_718#_c_387_n 0.0199289f $X=1.715 $Y=3.33 $X2=0 $Y2=0
cc_84 N_VGND_c_13_p N_A_193_718#_c_387_n 0.010808f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_85 N_VGND_M1011_b N_A_193_718#_c_391_n 0.0242504f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_86 N_VGND_c_21_p N_A_193_718#_c_391_n 0.0239528f $X=1.88 $Y=3.715 $X2=0 $Y2=0
cc_87 N_VGND_M1011_b N_A_193_718#_c_393_n 0.00542866f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_88 N_VGND_M1011_b N_A_193_718#_c_394_n 0.0107473f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_89 N_VGND_M1011_b N_A_193_718#_c_395_n 0.0119951f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_90 N_VGND_M1011_b N_VPWR_c_489_n 0.203486f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_91 N_VGND_M1011_b N_DESTPWR_c_516_n 0.203486f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_92 N_VGND_M1011_b N_X_c_572_n 0.117645f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_93 N_VGND_c_7_p N_X_c_572_n 0.02158f $X=3.27 $Y=3.715 $X2=0 $Y2=0
cc_94 N_VGND_c_71_p N_X_c_572_n 0.0234289f $X=4.41 $Y=3.33 $X2=0 $Y2=0
cc_95 N_VGND_c_13_p N_X_c_572_n 0.0126421f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_96 N_VPB_M1009_b N_A_M1009_g 0.0389027f $X=-0.025 $Y=-0.19 $X2=3.125 $Y2=3.59
cc_97 VPB N_A_M1009_g 0.00621856f $X=0.155 $Y=0.47 $X2=3.125 $Y2=3.59
cc_98 N_VPB_M1009_b N_A_M1001_g 0.0358449f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_99 N_VPB_M1009_b N_A_c_273_n 0.0183257f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_100 N_VPB_M1009_b N_A_278_47#_c_325_n 0.0369401f $X=-0.025 $Y=-0.19 $X2=0
+ $Y2=0
cc_101 N_VPB_M1009_b N_A_278_47#_c_315_n 0.0164461f $X=-0.025 $Y=-0.19 $X2=0
+ $Y2=0
cc_102 N_VPB_M1009_b N_A_278_47#_c_327_n 0.00836222f $X=-0.025 $Y=-0.19 $X2=0
+ $Y2=0
cc_103 N_VPB_M1009_b N_VPWR_c_490_n 0.0144492f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_490_n 0.0708842f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_105 N_VPB_M1009_b N_VPWR_c_492_n 0.0176917f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_492_n 0.0200925f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_107 N_VPB_M1009_b N_VPWR_c_494_n 0.119083f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_494_n 0.0200925f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_109 N_VPB_M1009_b N_VPWR_c_489_n 0.169196f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_489_n 0.0115306f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_489_n 0.0115306f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_112 N_VPB_M1009_b N_VPWR_c_499_n 0.00513431f $X=-0.025 $Y=-0.19 $X2=-0.025
+ $Y2=-0.245
cc_113 N_DESTVPB_M1014_b N_A_246_987#_M1014_g 0.0210833f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_114 N_DESTVPB_M1014_b N_A_246_987#_M1015_g 0.0168025f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_115 N_DESTVPB_M1014_b N_A_246_987#_c_171_n 0.00503307f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_116 N_DESTVPB_M1014_b N_A_246_987#_c_172_n 0.00748677f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_117 N_DESTVPB_M1014_b N_A_246_987#_c_173_n 0.00839347f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_118 N_DESTVPB_M1014_b N_A_246_987#_c_163_n 0.00415241f $X=-0.025 $Y=4.985
+ $X2=0.24 $Y2=3.245
cc_119 N_DESTVPB_M1014_b N_A_246_987#_c_175_n 0.00229064f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_120 N_DESTVPB_M1014_b N_A_246_987#_c_168_n 0.0274464f $X=-0.025 $Y=4.985
+ $X2=1.855 $Y2=3.415
cc_121 N_DESTVPB_M1014_b N_A_278_47#_c_319_n 0.00275879f $X=-0.025 $Y=4.985
+ $X2=-0.025 $Y2=-0.245
cc_122 N_DESTVPB_M1014_b N_A_278_47#_c_324_n 0.00363258f $X=-0.025 $Y=4.985
+ $X2=0.24 $Y2=3.415
cc_123 N_DESTVPB_M1014_b N_A_193_718#_c_396_n 0.0128194f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_124 N_DESTVPB_M1014_b N_A_193_718#_c_397_n 0.0167244f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_125 N_DESTVPB_M1014_b N_A_193_718#_c_398_n 0.0326863f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_126 N_DESTVPB_M1014_b N_A_193_718#_c_373_n 0.0340845f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_127 N_DESTVPB_M1014_b N_A_193_718#_c_374_n 0.00374597f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_128 N_DESTVPB_M1014_b N_A_193_718#_M1004_g 0.0285516f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_129 N_DESTVPB_M1014_b N_A_193_718#_c_379_n 0.00362008f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_130 N_DESTVPB_M1014_b N_A_193_718#_M1003_g 0.0328677f $X=-0.025 $Y=4.985
+ $X2=0.24 $Y2=3.415
cc_131 DESTVPB N_A_193_718#_M1003_g 0.00224388f $X=4.475 $Y=5.28 $X2=0.24
+ $Y2=3.415
cc_132 N_DESTVPB_M1014_b N_A_193_718#_c_384_n 0.0216804f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_133 N_DESTVPB_M1014_b N_A_193_718#_c_385_n 0.00159194f $X=-0.025 $Y=4.985
+ $X2=0.39 $Y2=3.33
cc_134 N_DESTVPB_M1014_b N_A_193_718#_c_386_n 0.00444583f $X=-0.025 $Y=4.985
+ $X2=0.74 $Y2=3.245
cc_135 N_DESTVPB_M1014_b N_A_193_718#_c_408_n 0.0137457f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_136 N_DESTVPB_M1014_b N_A_193_718#_c_393_n 3.94425e-19 $X=-0.025 $Y=4.985
+ $X2=4.56 $Y2=3.245
cc_137 N_DESTVPB_M1014_b N_A_193_718#_c_410_n 0.00291786f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_138 N_DESTVPB_M1014_b N_A_193_718#_c_395_n 0.0177627f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_139 DESTVPB N_A_193_718#_c_395_n 0.0438681f $X=0.155 $Y=5.28 $X2=0 $Y2=0
cc_140 N_DESTVPB_M1014_b N_A_193_718#_c_413_n 0.00803899f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_141 N_DESTVPB_M1014_b N_DESTPWR_c_517_n 4.89148e-19 $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_142 N_DESTVPB_M1014_b N_DESTPWR_c_518_n 0.0119037f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_143 N_DESTVPB_M1014_b N_DESTPWR_c_519_n 0.049514f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_144 DESTVPB N_DESTPWR_c_519_n 0.0200925f $X=0.155 $Y=5.28 $X2=0 $Y2=0
cc_145 N_DESTVPB_M1014_b N_DESTPWR_c_521_n 0.00436868f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_146 N_DESTVPB_M1014_b N_DESTPWR_c_522_n 0.0295949f $X=-0.025 $Y=4.985
+ $X2=0.24 $Y2=2.39
cc_147 N_DESTVPB_M1014_b N_DESTPWR_c_523_n 0.0385711f $X=-0.025 $Y=4.985
+ $X2=0.575 $Y2=3.33
cc_148 DESTVPB N_DESTPWR_c_523_n 0.0200925f $X=4.475 $Y=5.28 $X2=0.575 $Y2=3.33
cc_149 N_DESTVPB_M1014_b N_DESTPWR_c_516_n 0.091183f $X=-0.025 $Y=4.985 $X2=0.39
+ $Y2=3.33
cc_150 DESTVPB N_DESTPWR_c_516_n 0.0115306f $X=0.155 $Y=5.28 $X2=0.39 $Y2=3.33
cc_151 DESTVPB N_DESTPWR_c_516_n 0.0115306f $X=4.475 $Y=5.28 $X2=0.39 $Y2=3.33
cc_152 N_DESTVPB_M1014_b N_DESTPWR_c_528_n 0.00510842f $X=-0.025 $Y=4.985
+ $X2=0.74 $Y2=2.44
cc_153 N_DESTVPB_M1014_b N_X_c_572_n 0.0240847f $X=-0.025 $Y=4.985 $X2=0 $Y2=0
cc_154 DESTVPB N_X_c_572_n 0.0915263f $X=4.475 $Y=5.28 $X2=0 $Y2=0
cc_155 N_A_246_987#_c_168_n N_A_M1010_g 0.00436304f $X=1.665 $Y=5.1 $X2=0 $Y2=0
cc_156 N_A_246_987#_c_168_n N_A_M1005_g 0.00436304f $X=1.665 $Y=5.1 $X2=0 $Y2=0
cc_157 N_A_246_987#_c_164_n N_A_278_47#_c_306_n 4.25494e-19 $X=2.67 $Y=3.715
+ $X2=0 $Y2=0
cc_158 N_A_246_987#_c_171_n N_A_278_47#_c_309_n 4.27514e-19 $X=2.505 $Y=5.44
+ $X2=0 $Y2=0
cc_159 N_A_246_987#_c_159_n N_A_278_47#_c_311_n 0.00228462f $X=2.742 $Y=4.4
+ $X2=0 $Y2=0
cc_160 N_A_246_987#_c_164_n N_A_278_47#_c_311_n 0.0099858f $X=2.67 $Y=3.715
+ $X2=0 $Y2=0
cc_161 N_A_246_987#_c_171_n N_A_278_47#_c_319_n 0.00842185f $X=2.505 $Y=5.44
+ $X2=-0.025 $Y2=-0.245
cc_162 N_A_246_987#_c_172_n N_A_278_47#_c_319_n 0.0204053f $X=2.67 $Y=5.525
+ $X2=-0.025 $Y2=-0.245
cc_163 N_A_246_987#_c_159_n N_A_278_47#_c_319_n 0.0249802f $X=2.742 $Y=4.4
+ $X2=-0.025 $Y2=-0.245
cc_164 N_A_246_987#_c_163_n N_A_278_47#_c_319_n 0.0242161f $X=3.075 $Y=5.16
+ $X2=-0.025 $Y2=-0.245
cc_165 N_A_246_987#_c_164_n N_A_278_47#_c_319_n 0.0229888f $X=2.67 $Y=3.715
+ $X2=-0.025 $Y2=-0.245
cc_166 N_A_246_987#_c_172_n N_A_278_47#_c_324_n 6.09952e-19 $X=2.67 $Y=5.525
+ $X2=0.24 $Y2=3.415
cc_167 N_A_246_987#_c_159_n N_A_278_47#_c_324_n 0.00783532f $X=2.742 $Y=4.4
+ $X2=0.24 $Y2=3.415
cc_168 N_A_246_987#_c_163_n N_A_278_47#_c_324_n 0.00285919f $X=3.075 $Y=5.16
+ $X2=0.24 $Y2=3.415
cc_169 N_A_246_987#_c_171_n N_A_193_718#_c_396_n 0.013726f $X=2.505 $Y=5.44
+ $X2=0 $Y2=0
cc_170 N_A_246_987#_c_173_n N_A_193_718#_c_396_n 0.0027548f $X=2.67 $Y=5.55
+ $X2=0 $Y2=0
cc_171 N_A_246_987#_c_171_n N_A_193_718#_c_397_n 0.0108698f $X=2.505 $Y=5.44
+ $X2=0 $Y2=0
cc_172 N_A_246_987#_c_172_n N_A_193_718#_c_397_n 0.00226275f $X=2.67 $Y=5.525
+ $X2=0 $Y2=0
cc_173 N_A_246_987#_c_173_n N_A_193_718#_c_397_n 0.0146785f $X=2.67 $Y=5.55
+ $X2=0 $Y2=0
cc_174 N_A_246_987#_c_172_n N_A_193_718#_c_398_n 0.0298679f $X=2.67 $Y=5.525
+ $X2=0 $Y2=0
cc_175 N_A_246_987#_c_159_n N_A_193_718#_c_398_n 7.1387e-19 $X=2.742 $Y=4.4
+ $X2=0 $Y2=0
cc_176 N_A_246_987#_M1015_g N_A_193_718#_c_373_n 0.0268657f $X=1.665 $Y=5.925
+ $X2=0 $Y2=0
cc_177 N_A_246_987#_c_171_n N_A_193_718#_c_373_n 0.00266703f $X=2.505 $Y=5.44
+ $X2=0 $Y2=0
cc_178 N_A_246_987#_c_172_n N_A_193_718#_c_373_n 7.0281e-19 $X=2.67 $Y=5.525
+ $X2=0 $Y2=0
cc_179 N_A_246_987#_c_175_n N_A_193_718#_c_373_n 0.00130944f $X=1.515 $Y=5.1
+ $X2=0 $Y2=0
cc_180 N_A_246_987#_c_168_n N_A_193_718#_c_373_n 0.0219836f $X=1.665 $Y=5.1
+ $X2=0 $Y2=0
cc_181 N_A_246_987#_c_159_n N_A_193_718#_M1000_g 0.00601097f $X=2.742 $Y=4.4
+ $X2=0 $Y2=0
cc_182 N_A_246_987#_c_162_n N_A_193_718#_M1000_g 0.00330223f $X=2.67 $Y=4.275
+ $X2=0 $Y2=0
cc_183 N_A_246_987#_c_163_n N_A_193_718#_M1000_g 0.00898098f $X=3.075 $Y=5.16
+ $X2=0 $Y2=0
cc_184 N_A_246_987#_c_164_n N_A_193_718#_M1000_g 0.00109863f $X=2.67 $Y=3.715
+ $X2=0 $Y2=0
cc_185 N_A_246_987#_c_172_n N_A_193_718#_M1004_g 0.00431398f $X=2.67 $Y=5.525
+ $X2=0 $Y2=0
cc_186 N_A_246_987#_c_163_n N_A_193_718#_M1004_g 4.59228e-19 $X=3.075 $Y=5.16
+ $X2=0 $Y2=0
cc_187 N_A_246_987#_c_172_n N_A_193_718#_c_384_n 0.00891125f $X=2.67 $Y=5.525
+ $X2=0 $Y2=0
cc_188 N_A_246_987#_c_163_n N_A_193_718#_c_384_n 0.0164207f $X=3.075 $Y=5.16
+ $X2=0 $Y2=0
cc_189 N_A_246_987#_M1014_g N_A_193_718#_c_408_n 0.0139697f $X=1.305 $Y=5.925
+ $X2=0 $Y2=0
cc_190 N_A_246_987#_c_171_n N_A_193_718#_c_391_n 0.00619807f $X=2.505 $Y=5.44
+ $X2=3.27 $Y2=3.715
cc_191 N_A_246_987#_c_175_n N_A_193_718#_c_391_n 0.0252464f $X=1.515 $Y=5.1
+ $X2=3.27 $Y2=3.715
cc_192 N_A_246_987#_c_168_n N_A_193_718#_c_391_n 0.0102483f $X=1.665 $Y=5.1
+ $X2=3.27 $Y2=3.715
cc_193 N_A_246_987#_c_175_n N_A_193_718#_c_393_n 0.00138846f $X=1.515 $Y=5.1
+ $X2=4.56 $Y2=3.245
cc_194 N_A_246_987#_c_168_n N_A_193_718#_c_393_n 0.00132465f $X=1.665 $Y=5.1
+ $X2=4.56 $Y2=3.245
cc_195 N_A_246_987#_M1014_g N_A_193_718#_c_410_n 0.00381798f $X=1.305 $Y=5.925
+ $X2=0 $Y2=0
cc_196 N_A_246_987#_M1015_g N_A_193_718#_c_410_n 0.0029638f $X=1.665 $Y=5.925
+ $X2=0 $Y2=0
cc_197 N_A_246_987#_c_175_n N_A_193_718#_c_410_n 0.00581585f $X=1.515 $Y=5.1
+ $X2=0 $Y2=0
cc_198 N_A_246_987#_c_175_n N_A_193_718#_c_395_n 0.0299155f $X=1.515 $Y=5.1
+ $X2=0 $Y2=0
cc_199 N_A_246_987#_c_168_n N_A_193_718#_c_395_n 0.0143834f $X=1.665 $Y=5.1
+ $X2=0 $Y2=0
cc_200 N_A_246_987#_c_171_n N_A_193_718#_c_413_n 0.0290917f $X=2.505 $Y=5.44
+ $X2=0 $Y2=0
cc_201 N_A_246_987#_c_172_n N_A_193_718#_c_413_n 0.00109068f $X=2.67 $Y=5.525
+ $X2=0 $Y2=0
cc_202 N_A_246_987#_c_175_n N_A_193_718#_c_413_n 0.0129286f $X=1.515 $Y=5.1
+ $X2=0 $Y2=0
cc_203 N_A_246_987#_c_168_n N_A_193_718#_c_413_n 0.00119275f $X=1.665 $Y=5.1
+ $X2=0 $Y2=0
cc_204 N_A_246_987#_c_175_n A_276_1085# 0.00200208f $X=1.515 $Y=5.1 $X2=0.615
+ $Y2=2.23
cc_205 N_A_246_987#_c_171_n N_DESTPWR_M1015_d 0.00176461f $X=2.505 $Y=5.44
+ $X2=0.615 $Y2=2.23
cc_206 N_A_246_987#_M1014_g N_DESTPWR_c_517_n 0.00314212f $X=1.305 $Y=5.925
+ $X2=0 $Y2=0
cc_207 N_A_246_987#_M1015_g N_DESTPWR_c_517_n 0.0180441f $X=1.665 $Y=5.925 $X2=0
+ $Y2=0
cc_208 N_A_246_987#_c_171_n N_DESTPWR_c_517_n 0.0170777f $X=2.505 $Y=5.44 $X2=0
+ $Y2=0
cc_209 N_A_246_987#_c_173_n N_DESTPWR_c_517_n 0.0234201f $X=2.67 $Y=5.55 $X2=0
+ $Y2=0
cc_210 N_A_246_987#_c_172_n N_DESTPWR_c_518_n 0.00631144f $X=2.67 $Y=5.525 $X2=0
+ $Y2=0
cc_211 N_A_246_987#_c_173_n N_DESTPWR_c_518_n 0.0524911f $X=2.67 $Y=5.55 $X2=0
+ $Y2=0
cc_212 N_A_246_987#_M1014_g N_DESTPWR_c_519_n 0.00518588f $X=1.305 $Y=5.925
+ $X2=0 $Y2=0
cc_213 N_A_246_987#_M1015_g N_DESTPWR_c_519_n 0.00486043f $X=1.665 $Y=5.925
+ $X2=0 $Y2=0
cc_214 N_A_246_987#_c_173_n N_DESTPWR_c_522_n 0.019758f $X=2.67 $Y=5.55 $X2=0.24
+ $Y2=2.39
cc_215 N_A_246_987#_M1012_d N_DESTPWR_c_516_n 0.0023218f $X=2.53 $Y=5.425
+ $X2=0.39 $Y2=3.33
cc_216 N_A_246_987#_M1014_g N_DESTPWR_c_516_n 0.0103683f $X=1.305 $Y=5.925
+ $X2=0.39 $Y2=3.33
cc_217 N_A_246_987#_M1015_g N_DESTPWR_c_516_n 0.00814425f $X=1.665 $Y=5.925
+ $X2=0.39 $Y2=3.33
cc_218 N_A_246_987#_c_173_n N_DESTPWR_c_516_n 0.012508f $X=2.67 $Y=5.55 $X2=0.39
+ $Y2=3.33
cc_219 N_A_246_987#_c_171_n A_434_1085# 0.00366293f $X=2.505 $Y=5.44 $X2=0.615
+ $Y2=2.23
cc_220 N_A_M1005_g N_A_278_47#_c_306_n 0.0198552f $X=1.665 $Y=4.01 $X2=0 $Y2=0
cc_221 N_A_M1009_g N_A_278_47#_c_325_n 0.00339963f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_222 N_A_M1001_g N_A_278_47#_c_325_n 0.0148505f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_223 N_A_M1001_g N_A_278_47#_c_315_n 0.0266813f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_224 N_A_c_258_n N_A_278_47#_c_315_n 0.0140219f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_225 N_A_c_264_n N_A_278_47#_c_315_n 0.0223669f $X=1.745 $Y=2.925 $X2=0 $Y2=0
cc_226 N_A_c_269_n N_A_278_47#_c_315_n 0.00809784f $X=1.665 $Y=2.925 $X2=0 $Y2=0
cc_227 N_A_c_273_n N_A_278_47#_c_315_n 0.0500336f $X=1.16 $Y=1.832 $X2=0 $Y2=0
cc_228 N_A_c_264_n N_A_278_47#_c_316_n 0.0139563f $X=1.745 $Y=2.925 $X2=0 $Y2=0
cc_229 N_A_c_269_n N_A_278_47#_c_316_n 0.00454742f $X=1.665 $Y=2.925 $X2=0 $Y2=0
cc_230 N_A_M1005_g N_A_278_47#_c_319_n 0.00401063f $X=1.665 $Y=4.01 $X2=-0.025
+ $Y2=-0.245
cc_231 N_A_c_264_n N_A_278_47#_c_319_n 0.0175426f $X=1.745 $Y=2.925 $X2=-0.025
+ $Y2=-0.245
cc_232 N_A_c_269_n N_A_278_47#_c_319_n 0.00305169f $X=1.665 $Y=2.925 $X2=-0.025
+ $Y2=-0.245
cc_233 N_A_M1001_g N_A_278_47#_c_327_n 0.00684213f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_234 N_A_M1010_g N_A_193_718#_c_387_n 0.00781956f $X=1.305 $Y=4.01 $X2=0 $Y2=0
cc_235 N_A_M1010_g N_A_193_718#_c_391_n 0.00392017f $X=1.305 $Y=4.01 $X2=3.27
+ $Y2=3.715
cc_236 N_A_M1005_g N_A_193_718#_c_391_n 0.00352781f $X=1.665 $Y=4.01 $X2=3.27
+ $Y2=3.715
cc_237 N_A_M1009_g N_VPWR_c_490_n 0.0213886f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_238 N_A_M1001_g N_VPWR_c_490_n 0.00375886f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_239 N_A_c_267_n N_VPWR_c_490_n 0.00119966f $X=1.315 $Y=1.96 $X2=0 $Y2=0
cc_240 N_A_c_273_n N_VPWR_c_490_n 0.0154497f $X=1.16 $Y=1.832 $X2=0 $Y2=0
cc_241 N_A_M1009_g N_VPWR_c_494_n 0.00486043f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_242 N_A_M1001_g N_VPWR_c_494_n 0.00549284f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_243 N_A_M1009_g N_VPWR_c_489_n 0.00814425f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_244 N_A_M1001_g N_VPWR_c_489_n 0.0111098f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_245 N_A_278_47#_c_309_n N_A_193_718#_c_373_n 0.00233791f $X=2.38 $Y=4.615
+ $X2=0 $Y2=0
cc_246 N_A_278_47#_c_310_n N_A_193_718#_c_373_n 0.0157124f $X=2.17 $Y=4.615
+ $X2=0 $Y2=0
cc_247 N_A_278_47#_c_319_n N_A_193_718#_c_373_n 0.003329f $X=2.25 $Y=4.31 $X2=0
+ $Y2=0
cc_248 N_A_278_47#_c_324_n N_A_193_718#_c_373_n 0.0241477f $X=2.6 $Y=4.615 $X2=0
+ $Y2=0
cc_249 N_A_278_47#_c_324_n N_A_193_718#_M1000_g 0.00356709f $X=2.6 $Y=4.615
+ $X2=0 $Y2=0
cc_250 N_A_278_47#_c_324_n N_A_193_718#_c_384_n 0.00358313f $X=2.6 $Y=4.615
+ $X2=0 $Y2=0
cc_251 N_A_278_47#_c_310_n N_A_193_718#_c_391_n 0.00278759f $X=2.17 $Y=4.615
+ $X2=3.27 $Y2=3.715
cc_252 N_A_278_47#_c_319_n N_A_193_718#_c_391_n 0.0151734f $X=2.25 $Y=4.31
+ $X2=3.27 $Y2=3.715
cc_253 N_A_278_47#_c_324_n N_A_193_718#_c_391_n 5.58194e-19 $X=2.6 $Y=4.615
+ $X2=3.27 $Y2=3.715
cc_254 N_A_278_47#_c_319_n N_A_193_718#_c_393_n 0.00796579f $X=2.25 $Y=4.31
+ $X2=4.56 $Y2=3.245
cc_255 N_A_278_47#_c_324_n N_A_193_718#_c_393_n 6.34113e-19 $X=2.6 $Y=4.615
+ $X2=4.56 $Y2=3.245
cc_256 N_A_278_47#_c_310_n N_A_193_718#_c_413_n 0.00100861f $X=2.17 $Y=4.615
+ $X2=0 $Y2=0
cc_257 N_A_278_47#_c_319_n N_A_193_718#_c_413_n 0.0071736f $X=2.25 $Y=4.31 $X2=0
+ $Y2=0
cc_258 N_A_278_47#_c_325_n N_VPWR_c_490_n 0.0305839f $X=1.53 $Y=0.38 $X2=0 $Y2=0
cc_259 N_A_278_47#_c_325_n N_VPWR_c_494_n 0.0211337f $X=1.53 $Y=0.38 $X2=0 $Y2=0
cc_260 N_A_278_47#_M1001_d N_VPWR_c_489_n 0.00215406f $X=1.39 $Y=0.235 $X2=0
+ $Y2=0
cc_261 N_A_278_47#_c_325_n N_VPWR_c_489_n 0.0132819f $X=1.53 $Y=0.38 $X2=0 $Y2=0
cc_262 N_A_193_718#_c_396_n N_DESTPWR_c_517_n 0.0183086f $X=2.095 $Y=5.35 $X2=0
+ $Y2=0
cc_263 N_A_193_718#_c_397_n N_DESTPWR_c_517_n 0.00318727f $X=2.455 $Y=5.35 $X2=0
+ $Y2=0
cc_264 N_A_193_718#_c_408_n N_DESTPWR_c_517_n 0.0247854f $X=1.09 $Y=6.28 $X2=0
+ $Y2=0
cc_265 N_A_193_718#_c_397_n N_DESTPWR_c_518_n 0.00386407f $X=2.455 $Y=5.35 $X2=0
+ $Y2=0
cc_266 N_A_193_718#_c_374_n N_DESTPWR_c_518_n 0.00158632f $X=3.41 $Y=5.01 $X2=0
+ $Y2=0
cc_267 N_A_193_718#_M1004_g N_DESTPWR_c_518_n 0.0218301f $X=3.485 $Y=5.925 $X2=0
+ $Y2=0
cc_268 N_A_193_718#_M1003_g N_DESTPWR_c_518_n 0.00369509f $X=3.845 $Y=5.925
+ $X2=0 $Y2=0
cc_269 N_A_193_718#_c_384_n N_DESTPWR_c_518_n 0.00227815f $X=3.105 $Y=5.01 $X2=0
+ $Y2=0
cc_270 N_A_193_718#_c_408_n N_DESTPWR_c_519_n 0.0224101f $X=1.09 $Y=6.28 $X2=0
+ $Y2=0
cc_271 N_A_193_718#_c_396_n N_DESTPWR_c_522_n 0.00486043f $X=2.095 $Y=5.35
+ $X2=0.24 $Y2=2.39
cc_272 N_A_193_718#_c_397_n N_DESTPWR_c_522_n 0.00549284f $X=2.455 $Y=5.35
+ $X2=0.24 $Y2=2.39
cc_273 N_A_193_718#_M1004_g N_DESTPWR_c_523_n 0.00486043f $X=3.485 $Y=5.925
+ $X2=0.575 $Y2=3.33
cc_274 N_A_193_718#_M1003_g N_DESTPWR_c_523_n 0.0054895f $X=3.845 $Y=5.925
+ $X2=0.575 $Y2=3.33
cc_275 N_A_193_718#_M1014_s N_DESTPWR_c_516_n 0.00215158f $X=0.965 $Y=5.425
+ $X2=0.39 $Y2=3.33
cc_276 N_A_193_718#_c_396_n N_DESTPWR_c_516_n 0.00814425f $X=2.095 $Y=5.35
+ $X2=0.39 $Y2=3.33
cc_277 N_A_193_718#_c_397_n N_DESTPWR_c_516_n 0.0111098f $X=2.455 $Y=5.35
+ $X2=0.39 $Y2=3.33
cc_278 N_A_193_718#_M1004_g N_DESTPWR_c_516_n 0.00814425f $X=3.485 $Y=5.925
+ $X2=0.39 $Y2=3.33
cc_279 N_A_193_718#_M1003_g N_DESTPWR_c_516_n 0.0111095f $X=3.845 $Y=5.925
+ $X2=0.39 $Y2=3.33
cc_280 N_A_193_718#_c_408_n N_DESTPWR_c_516_n 0.0132444f $X=1.09 $Y=6.28
+ $X2=0.39 $Y2=3.33
cc_281 N_A_193_718#_M1000_g N_X_c_572_n 0.00528658f $X=3.485 $Y=4.01 $X2=0 $Y2=0
cc_282 N_A_193_718#_M1004_g N_X_c_572_n 0.00453972f $X=3.485 $Y=5.925 $X2=0
+ $Y2=0
cc_283 N_A_193_718#_M1013_g N_X_c_572_n 0.036079f $X=3.845 $Y=4.01 $X2=0 $Y2=0
cc_284 N_A_193_718#_M1003_g N_X_c_572_n 0.0286173f $X=3.845 $Y=5.925 $X2=0 $Y2=0
cc_285 N_A_193_718#_c_386_n N_X_c_572_n 0.0105303f $X=3.845 $Y=5.01 $X2=0 $Y2=0
cc_286 N_VPWR_c_489_n A_206_47# 0.00899413f $X=4.56 $Y=0 $X2=0.615 $Y2=2.23
cc_287 A_276_1085# N_DESTPWR_c_516_n 0.00899413f $X=1.38 $Y=5.425 $X2=2.742
+ $Y2=4.4
cc_288 N_DESTPWR_c_516_n A_434_1085# 0.00899413f $X=4.56 $Y=6.66 $X2=0.615
+ $Y2=2.23
cc_289 N_DESTPWR_c_516_n A_712_1085# 0.00899413f $X=4.56 $Y=6.66 $X2=0.615
+ $Y2=2.23
cc_290 N_DESTPWR_c_516_n N_X_M1003_d 0.00215158f $X=4.56 $Y=6.66 $X2=1.74
+ $Y2=3.59
cc_291 N_DESTPWR_c_518_n N_X_c_572_n 0.0302789f $X=3.27 $Y=5.585 $X2=0 $Y2=0
cc_292 N_DESTPWR_c_523_n N_X_c_572_n 0.0210467f $X=4.56 $Y=6.66 $X2=0 $Y2=0
cc_293 N_DESTPWR_c_516_n N_X_c_572_n 0.0125689f $X=4.56 $Y=6.66 $X2=0 $Y2=0
