* File: sky130_fd_sc_lp__mux2i_lp2.spice
* Created: Fri Aug 28 10:45:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2i_lp2.pex.spice"
.subckt sky130_fd_sc_lp__mux2i_lp2  VNB VPB S A0 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1005 A_256_47# N_S_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.3192 PD=0.66 PS=2.36 NRD=18.564 NRS=135.708 M=1 R=2.8 SA=75000.7
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A1_M1004_g A_256_47# VNB NSHORT L=0.15 W=0.42 AD=0.0609
+ AS=0.0504 PD=0.71 PS=0.66 NRD=1.428 NRS=18.564 M=1 R=2.8 SA=75001.1 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1010 A_422_47# N_A0_M1010_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.0714
+ AS=0.0609 PD=0.76 PS=0.71 NRD=32.856 NRS=1.428 M=1 R=2.8 SA=75001.5 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_490_21#_M1002_g A_422_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.0714 PD=0.715 PS=0.76 NRD=1.428 NRS=32.856 M=1 R=2.8 SA=75002
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1000 A_609_47# N_S_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.06195 PD=0.63 PS=0.715 NRD=14.28 NRS=2.856 M=1 R=2.8 SA=75002.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_490_21#_M1009_d N_S_M1009_g A_609_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_148_419# N_S_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.295 PD=1.24 PS=2.59 NRD=12.7853 NRS=1.9503 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1007 N_Y_M1007_d N_A0_M1007_g A_148_419# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.12 PD=1.57 PS=1.24 NRD=57.13 NRS=12.7853 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1008 A_410_419# N_A1_M1008_g N_Y_M1007_d VPB PHIGHVT L=0.25 W=1 AD=0.215
+ AS=0.285 PD=1.43 PS=1.57 NRD=31.5003 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A_490_21#_M1001_g A_410_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.16 AS=0.215 PD=1.32 PS=1.43 NRD=0 NRS=31.5003 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1003 N_A_490_21#_M1003_d N_S_M1003_g N_VPWR_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=7.8603 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX11_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__mux2i_lp2.pxi.spice"
*
.ends
*
*
