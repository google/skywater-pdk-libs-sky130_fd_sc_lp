* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2111o_m A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 X a_85_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_503_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A2 a_411_369# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND B1 a_85_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_85_21# A1 a_503_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_411_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_339_369# B1 a_411_369# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND D1 a_85_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_85_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_85_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_85_21# D1 a_267_369# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_267_369# C1 a_339_369# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
