* File: sky130_fd_sc_lp__sdlclkp_2.pex.spice
* Created: Wed Sep  2 10:37:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%SCE 2 5 8 10 11 12 13 14 20 22
r27 20 22 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.352 $Y=1.045
+ $X2=0.352 $Y2=0.88
r28 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.32
+ $Y=1.045 $X2=0.32 $Y2=1.045
r29 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.665
+ $X2=0.25 $Y2=2.035
r30 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.665
r31 12 21 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.045
r32 11 21 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.25 $Y=0.925
+ $X2=0.25 $Y2=1.045
r33 8 10 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.475 $Y=2.66
+ $X2=0.475 $Y2=1.55
r34 5 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.56
+ $X2=0.475 $Y2=0.88
r35 2 10 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.352 $Y=1.353
+ $X2=0.352 $Y2=1.55
r36 1 20 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.352 $Y=1.077
+ $X2=0.352 $Y2=1.045
r37 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.352 $Y=1.077
+ $X2=0.352 $Y2=1.353
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%GATE 3 7 11 12 13 16
c45 3 0 1.90777e-19 $X=0.835 $Y=2.66
r46 16 18 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.007 $Y=1.47
+ $X2=1.007 $Y2=1.305
r47 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.02
+ $Y=1.47 $X2=1.02 $Y2=1.47
r48 13 17 3.21335 $w=6.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.2 $Y=1.64 $X2=1.02
+ $Y2=1.64
r49 11 12 44.0658 $w=3.55e-07 $l=1.5e-07 $layer=POLY_cond $X=0.972 $Y=1.825
+ $X2=0.972 $Y2=1.975
r50 9 16 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=1.007 $Y=1.482
+ $X2=1.007 $Y2=1.47
r51 9 11 55.7537 $w=3.55e-07 $l=3.43e-07 $layer=POLY_cond $X=1.007 $Y=1.482
+ $X2=1.007 $Y2=1.825
r52 7 18 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.905 $Y=0.56
+ $X2=0.905 $Y2=1.305
r53 3 12 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.835 $Y=2.66
+ $X2=0.835 $Y2=1.975
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%A_282_70# 1 2 7 9 13 17 19 22 27 30 31 32
+ 33 35 37
c77 7 0 1.68021e-19 $X=3.35 $Y=1.66
r78 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.43
+ $Y=1.75 $X2=2.43 $Y2=1.75
r79 33 39 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=1.915
+ $X2=2.415 $Y2=1.75
r80 33 35 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=2.415 $Y=1.915
+ $X2=2.415 $Y2=2.21
r81 31 39 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.305 $Y=1.75
+ $X2=2.415 $Y2=1.75
r82 31 32 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.305 $Y=1.75
+ $X2=1.715 $Y2=1.75
r83 30 32 7.10306 $w=3.3e-07 $l=2.14942e-07 $layer=LI1_cond $X=1.6 $Y=1.585
+ $X2=1.715 $Y2=1.75
r84 30 37 23.0489 $w=2.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.6 $Y=1.585 $X2=1.6
+ $Y2=1.125
r85 25 37 6.3332 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=1.567 $Y=0.978
+ $X2=1.567 $Y2=1.125
r86 25 27 16.3295 $w=2.93e-07 $l=4.18e-07 $layer=LI1_cond $X=1.567 $Y=0.978
+ $X2=1.567 $Y2=0.56
r87 22 40 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.62 $Y=1.75
+ $X2=2.43 $Y2=1.75
r88 22 23 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.695 $Y=1.75 $X2=2.695
+ $Y2=2.05
r89 19 22 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.695 $Y=1.66
+ $X2=2.695 $Y2=1.75
r90 15 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.425 $Y=1.585
+ $X2=3.425 $Y2=0.875
r91 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.225 $Y=2.125
+ $X2=3.225 $Y2=2.495
r92 10 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.77 $Y=2.05
+ $X2=2.695 $Y2=2.05
r93 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.15 $Y=2.05
+ $X2=3.225 $Y2=2.125
r94 9 10 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=3.15 $Y=2.05 $X2=2.77
+ $Y2=2.05
r95 8 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.77 $Y=1.66
+ $X2=2.695 $Y2=1.66
r96 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.35 $Y=1.66
+ $X2=3.425 $Y2=1.585
r97 7 8 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.35 $Y=1.66 $X2=2.77
+ $Y2=1.66
r98 2 35 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=2.055
+ $Y=2.085 $X2=2.39 $Y2=2.21
r99 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.35 $X2=1.55 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%A_250_443# 1 2 8 9 11 12 13 15 18 20 21 22
+ 24 27 31 38 41 43 44 49 56
c130 31 0 1.75311e-19 $X=1.505 $Y=2.29
c131 27 0 1.0624e-19 $X=3.655 $Y=2.495
r132 53 56 6.36149 $w=2.48e-07 $l=1.38e-07 $layer=LI1_cond $X=5.157 $Y=2.24
+ $X2=5.295 $Y2=2.24
r133 51 52 5.00426 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=0.61
+ $X2=5.115 $Y2=0.695
r134 49 51 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=5.115 $Y=0.53
+ $X2=5.115 $Y2=0.61
r135 43 46 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.07 $Y=0.35
+ $X2=2.07 $Y2=0.61
r136 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.07
+ $Y=0.35 $X2=2.07 $Y2=0.35
r137 41 53 2.85067 $w=1.75e-07 $l=1.25e-07 $layer=LI1_cond $X=5.157 $Y=2.115
+ $X2=5.157 $Y2=2.24
r138 41 52 89.9948 $w=1.73e-07 $l=1.42e-06 $layer=LI1_cond $X=5.157 $Y=2.115
+ $X2=5.157 $Y2=0.695
r139 39 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=0.61
+ $X2=2.07 $Y2=0.61
r140 38 51 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.985 $Y=0.61
+ $X2=5.115 $Y2=0.61
r141 38 39 179.412 $w=1.68e-07 $l=2.75e-06 $layer=LI1_cond $X=4.985 $Y=0.61
+ $X2=2.235 $Y2=0.61
r142 37 44 92.6765 $w=3.3e-07 $l=5.3e-07 $layer=POLY_cond $X=2.07 $Y=0.88
+ $X2=2.07 $Y2=0.35
r143 36 37 7.94458 $w=3.3e-07 $l=2.32e-07 $layer=POLY_cond $X=2.07 $Y=1.112
+ $X2=2.07 $Y2=0.88
r144 35 36 10.5805 $w=4.1e-07 $l=9e-08 $layer=POLY_cond $X=1.98 $Y=1.112
+ $X2=2.07 $Y2=1.112
r145 34 35 55.8415 $w=4.1e-07 $l=4.75e-07 $layer=POLY_cond $X=1.505 $Y=1.112
+ $X2=1.98 $Y2=1.112
r146 29 31 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.325 $Y=2.29
+ $X2=1.505 $Y2=2.29
r147 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.655 $Y=3.075
+ $X2=3.655 $Y2=2.495
r148 22 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.995 $Y=1.195
+ $X2=2.995 $Y2=0.875
r149 21 36 39.7867 $w=4.1e-07 $l=2.30857e-07 $layer=POLY_cond $X=2.235 $Y=1.27
+ $X2=2.07 $Y2=1.112
r150 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.92 $Y=1.27
+ $X2=2.995 $Y2=1.195
r151 20 21 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.92 $Y=1.27
+ $X2=2.235 $Y2=1.27
r152 16 35 26.4667 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.98 $Y=1.345
+ $X2=1.98 $Y2=1.112
r153 16 18 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=1.98 $Y=1.345
+ $X2=1.98 $Y2=2.405
r154 15 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.505 $Y=2.215
+ $X2=1.505 $Y2=2.29
r155 14 34 26.4667 $w=1.5e-07 $l=2.33e-07 $layer=POLY_cond $X=1.505 $Y=1.345
+ $X2=1.505 $Y2=1.112
r156 14 15 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.505 $Y=1.345
+ $X2=1.505 $Y2=2.215
r157 12 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.58 $Y=3.15
+ $X2=3.655 $Y2=3.075
r158 12 13 1117.83 $w=1.5e-07 $l=2.18e-06 $layer=POLY_cond $X=3.58 $Y=3.15
+ $X2=1.4 $Y2=3.15
r159 9 34 19.9854 $w=4.1e-07 $l=3.05392e-07 $layer=POLY_cond $X=1.335 $Y=0.88
+ $X2=1.505 $Y2=1.112
r160 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.335 $Y=0.88
+ $X2=1.335 $Y2=0.56
r161 8 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.325 $Y=3.075
+ $X2=1.4 $Y2=3.15
r162 7 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.325 $Y=2.365
+ $X2=1.325 $Y2=2.29
r163 7 8 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.325 $Y=2.365
+ $X2=1.325 $Y2=3.075
r164 2 56 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.15
+ $Y=2.145 $X2=5.295 $Y2=2.28
r165 1 49 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=5.025
+ $Y=0.37 $X2=5.15 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%A_742_107# 1 2 9 13 17 19 20 23 27 28 30
+ 37 40 43 44 47 48 49 52 53 56 61 62 67
c139 56 0 2.74261e-19 $X=3.875 $Y=1.75
r140 57 67 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.875 $Y=1.75
+ $X2=4.015 $Y2=1.75
r141 57 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.875 $Y=1.75
+ $X2=3.785 $Y2=1.75
r142 56 59 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=3.877 $Y=1.75
+ $X2=3.877 $Y2=1.83
r143 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.875
+ $Y=1.75 $X2=3.875 $Y2=1.75
r144 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.55
+ $Y=1.48 $X2=6.55 $Y2=1.48
r145 50 52 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.55 $Y=1.735
+ $X2=6.55 $Y2=1.48
r146 48 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.385 $Y=1.82
+ $X2=6.55 $Y2=1.735
r147 48 49 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.385 $Y=1.82
+ $X2=5.955 $Y2=1.82
r148 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.87 $Y=1.905
+ $X2=5.955 $Y2=1.82
r149 46 47 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.87 $Y=1.905
+ $X2=5.87 $Y2=2.535
r150 45 62 2.76166 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.92 $Y=2.62
+ $X2=4.79 $Y2=2.62
r151 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.785 $Y=2.62
+ $X2=5.87 $Y2=2.535
r152 44 45 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=5.785 $Y=2.62
+ $X2=4.92 $Y2=2.62
r153 43 61 4.40882 $w=2.05e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.815 $Y=1.745
+ $X2=4.78 $Y2=1.83
r154 42 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.815 $Y=1.055
+ $X2=4.815 $Y2=1.745
r155 38 62 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.79 $Y=2.705
+ $X2=4.79 $Y2=2.62
r156 38 40 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=4.79 $Y=2.705
+ $X2=4.79 $Y2=2.91
r157 35 62 3.70735 $w=2.5e-07 $l=8.9861e-08 $layer=LI1_cond $X=4.78 $Y=2.535
+ $X2=4.79 $Y2=2.62
r158 35 37 27.1304 $w=2.38e-07 $l=5.65e-07 $layer=LI1_cond $X=4.78 $Y=2.535
+ $X2=4.78 $Y2=1.97
r159 34 61 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=1.915
+ $X2=4.78 $Y2=1.83
r160 34 37 2.64102 $w=2.38e-07 $l=5.5e-08 $layer=LI1_cond $X=4.78 $Y=1.915
+ $X2=4.78 $Y2=1.97
r161 30 42 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.73 $Y=0.96
+ $X2=4.815 $Y2=1.055
r162 30 32 8.17225 $w=1.88e-07 $l=1.4e-07 $layer=LI1_cond $X=4.73 $Y=0.96
+ $X2=4.59 $Y2=0.96
r163 29 59 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=4.04 $Y=1.83
+ $X2=3.877 $Y2=1.83
r164 28 61 2.0246 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.66 $Y=1.83 $X2=4.78
+ $Y2=1.83
r165 28 29 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.66 $Y=1.83
+ $X2=4.04 $Y2=1.83
r166 26 53 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.55 $Y=1.82
+ $X2=6.55 $Y2=1.48
r167 26 27 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=1.82
+ $X2=6.55 $Y2=1.985
r168 25 53 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.55 $Y=1.465
+ $X2=6.55 $Y2=1.48
r169 23 27 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.53 $Y=2.465
+ $X2=6.53 $Y2=1.985
r170 19 25 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.385 $Y=1.39
+ $X2=6.55 $Y2=1.465
r171 19 20 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=6.385 $Y=1.39
+ $X2=6.23 $Y2=1.39
r172 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.155 $Y=1.315
+ $X2=6.23 $Y2=1.39
r173 15 17 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=6.155 $Y=1.315
+ $X2=6.155 $Y2=0.58
r174 11 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.915
+ $X2=4.015 $Y2=1.75
r175 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.015 $Y=1.915
+ $X2=4.015 $Y2=2.495
r176 7 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.585
+ $X2=3.785 $Y2=1.75
r177 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.785 $Y=1.585
+ $X2=3.785 $Y2=0.875
r178 2 40 400 $w=1.7e-07 $l=1.15288e-06 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=1.825 $X2=4.755 $Y2=2.91
r179 2 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=1.825 $X2=4.755 $Y2=1.97
r180 1 32 182 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_NDIFF $count=1 $X=4.45
+ $Y=0.245 $X2=4.59 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%A_614_133# 1 2 9 13 17 19 22 26 30
c63 13 0 1.40694e-19 $X=4.54 $Y=2.455
r64 30 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.465 $Y=1.39
+ $X2=4.465 $Y2=1.555
r65 30 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.465 $Y=1.39
+ $X2=4.465 $Y2=1.225
r66 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.465
+ $Y=1.39 $X2=4.465 $Y2=1.39
r67 26 29 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=4.43 $Y=1.31 $X2=4.43
+ $Y2=1.39
r68 24 25 5.27994 $w=4.98e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=1.31
+ $X2=3.295 $Y2=1.395
r69 22 24 8.61176 $w=4.98e-07 $l=3.6e-07 $layer=LI1_cond $X=3.295 $Y=0.95
+ $X2=3.295 $Y2=1.31
r70 20 24 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=3.545 $Y=1.31
+ $X2=3.295 $Y2=1.31
r71 19 26 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.3 $Y=1.31 $X2=4.43
+ $Y2=1.31
r72 19 20 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.3 $Y=1.31
+ $X2=3.545 $Y2=1.31
r73 17 25 52.5802 $w=2.38e-07 $l=1.095e-06 $layer=LI1_cond $X=3.425 $Y=2.49
+ $X2=3.425 $Y2=1.395
r74 13 34 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=4.54 $Y=2.455 $X2=4.54
+ $Y2=1.555
r75 9 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.375 $Y=0.665
+ $X2=4.375 $Y2=1.225
r76 2 17 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=2.285 $X2=3.44 $Y2=2.49
r77 1 22 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.665 $X2=3.21 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%CLK 1 3 4 6 8 10 11 15 17 18 19 35
c66 4 0 1.40694e-19 $X=5.51 $Y=1.855
r67 28 35 2.55074 $w=3.73e-07 $l=8.3e-08 $layer=LI1_cond $X=5.602 $Y=1.378
+ $X2=5.602 $Y2=1.295
r68 25 27 64.2966 $w=5.36e-07 $l=7.15e-07 $layer=POLY_cond $X=5.58 $Y=1.065
+ $X2=5.58 $Y2=1.78
r69 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.52
+ $Y=1.065 $X2=5.52 $Y2=1.065
r70 18 19 12.8279 $w=2.72e-07 $l=2.86e-07 $layer=LI1_cond $X=5.602 $Y=1.379
+ $X2=5.602 $Y2=1.665
r71 18 28 0.974138 $w=3.75e-07 $l=1e-09 $layer=LI1_cond $X=5.602 $Y=1.379
+ $X2=5.602 $Y2=1.378
r72 18 35 0.0307318 $w=3.73e-07 $l=1e-09 $layer=LI1_cond $X=5.602 $Y=1.294
+ $X2=5.602 $Y2=1.295
r73 18 26 7.03759 $w=3.73e-07 $l=2.29e-07 $layer=LI1_cond $X=5.602 $Y=1.294
+ $X2=5.602 $Y2=1.065
r74 17 26 4.30245 $w=3.73e-07 $l=1.4e-07 $layer=LI1_cond $X=5.602 $Y=0.925
+ $X2=5.602 $Y2=1.065
r75 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.1 $Y=1.855 $X2=6.1
+ $Y2=2.465
r76 12 27 33.1734 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.87 $Y=1.78
+ $X2=5.58 $Y2=1.78
r77 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.025 $Y=1.78
+ $X2=6.1 $Y2=1.855
r78 11 12 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=6.025 $Y=1.78
+ $X2=5.87 $Y2=1.78
r79 8 25 31.7333 $w=2.68e-07 $l=2.85832e-07 $layer=POLY_cond $X=5.795 $Y=0.9
+ $X2=5.58 $Y2=1.065
r80 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.795 $Y=0.9
+ $X2=5.795 $Y2=0.58
r81 4 27 34.7758 $w=5.36e-07 $l=1.04283e-07 $layer=POLY_cond $X=5.51 $Y=1.855
+ $X2=5.58 $Y2=1.78
r82 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.51 $Y=1.855 $X2=5.51
+ $Y2=2.465
r83 1 25 31.7333 $w=2.68e-07 $l=2.85832e-07 $layer=POLY_cond $X=5.365 $Y=0.9
+ $X2=5.58 $Y2=1.065
r84 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.365 $Y=0.9 $X2=5.365
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%A_1235_429# 1 2 9 13 19 23 25 30 32 34 35
+ 37 38 42 43 46 47 49
r98 48 49 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.665 $Y=1.46
+ $X2=7.59 $Y2=1.46
r99 43 48 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.88 $Y=1.46
+ $X2=7.665 $Y2=1.46
r100 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.88
+ $Y=1.46 $X2=7.88 $Y2=1.46
r101 40 42 33.4652 $w=2.58e-07 $l=7.55e-07 $layer=LI1_cond $X=7.915 $Y=2.215
+ $X2=7.915 $Y2=1.46
r102 39 47 4.80229 $w=2.4e-07 $l=1.40712e-07 $layer=LI1_cond $X=7.115 $Y=2.3
+ $X2=7.005 $Y2=2.23
r103 38 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.785 $Y=2.3
+ $X2=7.915 $Y2=2.215
r104 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.785 $Y=2.3
+ $X2=7.115 $Y2=2.3
r105 37 47 1.65768 $w=2.2e-07 $l=1.55e-07 $layer=LI1_cond $X=7.005 $Y=2.075
+ $X2=7.005 $Y2=2.23
r106 36 37 45.05 $w=2.18e-07 $l=8.6e-07 $layer=LI1_cond $X=7.005 $Y=1.215
+ $X2=7.005 $Y2=2.075
r107 34 36 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.895 $Y=1.13
+ $X2=7.005 $Y2=1.215
r108 34 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.895 $Y=1.13
+ $X2=6.535 $Y2=1.13
r109 33 46 3.1405 $w=3.1e-07 $l=1.3e-07 $layer=LI1_cond $X=6.41 $Y=2.23 $X2=6.28
+ $Y2=2.23
r110 32 47 4.80229 $w=2.4e-07 $l=1.1e-07 $layer=LI1_cond $X=6.895 $Y=2.23
+ $X2=7.005 $Y2=2.23
r111 32 33 18.0302 $w=3.08e-07 $l=4.85e-07 $layer=LI1_cond $X=6.895 $Y=2.23
+ $X2=6.41 $Y2=2.23
r112 28 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.37 $Y=1.045
+ $X2=6.535 $Y2=1.13
r113 28 30 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.37 $Y=1.045
+ $X2=6.37 $Y2=0.555
r114 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.665 $Y=1.625
+ $X2=7.665 $Y2=1.46
r115 21 23 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=7.665 $Y=1.625
+ $X2=7.665 $Y2=2.465
r116 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.665 $Y=1.295
+ $X2=7.665 $Y2=1.46
r117 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.665 $Y=1.295
+ $X2=7.665 $Y2=0.695
r118 16 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.31 $Y=1.37
+ $X2=7.235 $Y2=1.37
r119 16 49 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.31 $Y=1.37
+ $X2=7.59 $Y2=1.37
r120 11 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.235 $Y=1.445
+ $X2=7.235 $Y2=1.37
r121 11 13 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=7.235 $Y=1.445
+ $X2=7.235 $Y2=2.465
r122 7 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.235 $Y=1.295
+ $X2=7.235 $Y2=1.37
r123 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.235 $Y=1.295 $X2=7.235
+ $Y2=0.695
r124 2 46 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=6.175
+ $Y=2.145 $X2=6.315 $Y2=2.32
r125 1 30 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.23
+ $Y=0.37 $X2=6.37 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%VPWR 1 2 3 4 5 6 19 21 25 29 35 39 43 45
+ 48 49 50 52 57 69 73 82 85 88 92
c100 25 0 1.90777e-19 $X=1.63 $Y=2.6
r101 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r102 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r103 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 77 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 77 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r107 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r108 74 88 12.6176 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=7.185 $Y=3.33
+ $X2=6.882 $Y2=3.33
r109 74 76 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.185 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 73 91 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.937 $Y2=3.33
r111 73 76 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 72 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r113 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 69 88 12.6176 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=6.58 $Y=3.33
+ $X2=6.882 $Y2=3.33
r115 69 71 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.58 $Y=3.33 $X2=6.48
+ $Y2=3.33
r116 68 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r117 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r118 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r120 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r121 62 85 10.508 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=4.267 $Y2=3.33
r122 62 64 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.49 $Y=3.33 $X2=4.56
+ $Y2=3.33
r123 61 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r124 60 61 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r125 58 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.63 $Y2=3.33
r126 58 60 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=2.16 $Y2=3.33
r127 57 85 10.508 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.267 $Y2=3.33
r128 57 60 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 56 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r130 56 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r131 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 53 79 4.68586 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.207 $Y2=3.33
r133 53 55 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=1.2 $Y2=3.33
r134 52 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.63 $Y2=3.33
r135 52 55 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 50 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r137 50 61 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 50 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r139 48 67 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=5.64 $Y=3.33
+ $X2=5.52 $Y2=3.33
r140 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.64 $Y=3.33
+ $X2=5.805 $Y2=3.33
r141 47 71 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.97 $Y=3.33
+ $X2=6.48 $Y2=3.33
r142 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.97 $Y=3.33
+ $X2=5.805 $Y2=3.33
r143 43 91 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.937 $Y2=3.33
r144 43 45 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.88 $Y2=2.72
r145 39 42 6.12867 $w=6.03e-07 $l=3.1e-07 $layer=LI1_cond $X=6.882 $Y=2.64
+ $X2=6.882 $Y2=2.95
r146 37 88 2.53987 $w=6.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.882 $Y=3.245
+ $X2=6.882 $Y2=3.33
r147 37 42 5.83212 $w=6.03e-07 $l=2.95e-07 $layer=LI1_cond $X=6.882 $Y=3.245
+ $X2=6.882 $Y2=2.95
r148 33 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.805 $Y=3.245
+ $X2=5.805 $Y2=3.33
r149 33 35 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.805 $Y=3.245
+ $X2=5.805 $Y2=2.96
r150 29 32 19.9411 $w=4.43e-07 $l=7.7e-07 $layer=LI1_cond $X=4.267 $Y=2.17
+ $X2=4.267 $Y2=2.94
r151 27 85 1.76584 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.267 $Y=3.245
+ $X2=4.267 $Y2=3.33
r152 27 32 7.89877 $w=4.43e-07 $l=3.05e-07 $layer=LI1_cond $X=4.267 $Y=3.245
+ $X2=4.267 $Y2=2.94
r153 23 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r154 23 25 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.6
r155 19 79 2.99625 $w=3.2e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.207 $Y2=3.33
r156 19 21 27.0104 $w=3.18e-07 $l=7.5e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.495
r157 6 45 600 $w=1.7e-07 $l=9.52431e-07 $layer=licon1_PDIFF $count=1 $X=7.74
+ $Y=1.835 $X2=7.88 $Y2=2.72
r158 5 42 600 $w=1.7e-07 $l=9.9101e-07 $layer=licon1_PDIFF $count=1 $X=6.605
+ $Y=2.145 $X2=7.02 $Y2=2.95
r159 5 39 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=6.605
+ $Y=2.145 $X2=6.745 $Y2=2.64
r160 4 35 600 $w=1.7e-07 $l=9.18436e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=2.145 $X2=5.805 $Y2=2.96
r161 3 32 600 $w=1.7e-07 $l=7.63512e-07 $layer=licon1_PDIFF $count=1 $X=4.09
+ $Y=2.285 $X2=4.325 $Y2=2.94
r162 3 29 300 $w=1.7e-07 $l=2.86793e-07 $layer=licon1_PDIFF $count=2 $X=4.09
+ $Y=2.285 $X2=4.325 $Y2=2.17
r163 2 25 600 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_PDIFF $count=1 $X=1.475
+ $Y=2.44 $X2=1.63 $Y2=2.6
r164 1 21 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.34 $X2=0.26 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%A_110_70# 1 2 3 4 14 17 21 23 26 27 28 32
+ 34 35 37 41 42
c82 26 0 1.75311e-19 $X=2.05 $Y=2.895
r83 41 42 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=2.49
+ $X2=2.915 $Y2=2.325
r84 39 42 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=2.78 $Y=1.125
+ $X2=2.78 $Y2=2.325
r85 37 39 8.8114 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.7 $Y=0.95 $X2=2.7
+ $Y2=1.125
r86 33 34 10.4473 $w=2.23e-07 $l=1.9e-07 $layer=LI1_cond $X=0.702 $Y=0.74
+ $X2=0.702 $Y2=0.93
r87 31 41 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=2.915 $Y=2.545
+ $X2=2.915 $Y2=2.49
r88 31 32 9.16716 $w=4.38e-07 $l=3.5e-07 $layer=LI1_cond $X=2.915 $Y=2.545
+ $X2=2.915 $Y2=2.895
r89 27 32 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=2.695 $Y=2.98
+ $X2=2.915 $Y2=2.895
r90 27 28 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.695 $Y=2.98
+ $X2=2.135 $Y2=2.98
r91 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.05 $Y=2.895
+ $X2=2.135 $Y2=2.98
r92 25 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.05 $Y=2.335
+ $X2=2.05 $Y2=2.895
r93 24 35 4.54334 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=1.215 $Y=2.25
+ $X2=0.9 $Y2=2.25
r94 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.965 $Y=2.25
+ $X2=2.05 $Y2=2.335
r95 23 24 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.965 $Y=2.25
+ $X2=1.215 $Y2=2.25
r96 21 33 9.21954 $w=2.23e-07 $l=1.8e-07 $layer=LI1_cond $X=0.707 $Y=0.56
+ $X2=0.707 $Y2=0.74
r97 15 35 2.41844 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=2.335 $X2=0.9
+ $Y2=2.25
r98 15 17 2.84781 $w=6.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.9 $Y=2.335 $X2=0.9
+ $Y2=2.485
r99 14 35 2.41844 $w=4e-07 $l=2.69165e-07 $layer=LI1_cond $X=0.67 $Y=2.165
+ $X2=0.9 $Y2=2.25
r100 14 34 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=0.67 $Y=2.165
+ $X2=0.67 $Y2=0.93
r101 4 41 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=2.885
+ $Y=2.285 $X2=3.01 $Y2=2.49
r102 3 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=2.34 $X2=1.05 $Y2=2.485
r103 2 37 182 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.665 $X2=2.7 $Y2=0.95
r104 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.35 $X2=0.69 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%GCLK 1 2 9 12 13 14 15 21
r20 14 15 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.48 $Y=1.295
+ $X2=7.48 $Y2=1.665
r21 13 14 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.48 $Y=0.925
+ $X2=7.48 $Y2=1.295
r22 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.48 $Y=0.555
+ $X2=7.48 $Y2=0.925
r23 12 21 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.48 $Y=0.555
+ $X2=7.48 $Y2=0.42
r24 10 15 8.10978 $w=2.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.48 $Y=1.855
+ $X2=7.48 $Y2=1.665
r25 9 10 4.08188 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.45 $Y=1.96
+ $X2=7.45 $Y2=1.855
r26 2 9 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.31
+ $Y=1.835 $X2=7.45 $Y2=1.96
r27 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.31
+ $Y=0.275 $X2=7.45 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_2%VGND 1 2 3 4 5 6 19 21 25 29 33 35 37 39
+ 41 46 51 56 61 70 74 80 83 87
r91 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r92 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r93 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r94 74 77 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=4.08
+ $Y2=0.27
r95 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r96 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r97 65 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r98 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r99 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r100 62 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=0 $X2=7.01
+ $Y2=0
r101 62 64 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.175 $Y=0
+ $X2=7.44 $Y2=0
r102 61 86 4.09935 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=7.785 $Y=0
+ $X2=7.972 $Y2=0
r103 61 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.785 $Y=0 $X2=7.44
+ $Y2=0
r104 60 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r105 60 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=5.52
+ $Y2=0
r106 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r107 57 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.745 $Y=0 $X2=5.58
+ $Y2=0
r108 57 59 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=5.745 $Y=0
+ $X2=6.48 $Y2=0
r109 56 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=0 $X2=7.01
+ $Y2=0
r110 56 59 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.845 $Y=0
+ $X2=6.48 $Y2=0
r111 55 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r112 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r113 52 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.245 $Y=0 $X2=4.08
+ $Y2=0
r114 52 54 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.245 $Y=0
+ $X2=5.04 $Y2=0
r115 51 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.415 $Y=0 $X2=5.58
+ $Y2=0
r116 51 54 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.415 $Y=0
+ $X2=5.04 $Y2=0
r117 50 71 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=1.2
+ $Y2=0
r118 49 50 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r119 47 70 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.12
+ $Y2=0
r120 47 49 153.316 $w=1.68e-07 $l=2.35e-06 $layer=LI1_cond $X=1.25 $Y=0 $X2=3.6
+ $Y2=0
r121 46 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=4.08
+ $Y2=0
r122 46 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=3.6
+ $Y2=0
r123 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r124 45 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r125 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r126 42 67 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r127 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r128 41 70 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.12
+ $Y2=0
r129 41 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r130 39 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r131 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r132 39 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r133 35 86 3.11287 $w=2.6e-07 $l=1.09864e-07 $layer=LI1_cond $X=7.915 $Y=0.085
+ $X2=7.972 $Y2=0
r134 35 37 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=7.915 $Y=0.085
+ $X2=7.915 $Y2=0.42
r135 31 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.01 $Y=0.085
+ $X2=7.01 $Y2=0
r136 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.01 $Y=0.085
+ $X2=7.01 $Y2=0.42
r137 27 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=0.085
+ $X2=5.58 $Y2=0
r138 27 29 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=5.58 $Y=0.085
+ $X2=5.58 $Y2=0.545
r139 23 70 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r140 23 25 21.0542 $w=2.58e-07 $l=4.75e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.56
r141 19 67 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r142 19 21 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.545
r143 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.275 $X2=7.88 $Y2=0.42
r144 5 33 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.885
+ $Y=0.275 $X2=7.01 $Y2=0.42
r145 4 29 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=5.44
+ $Y=0.37 $X2=5.58 $Y2=0.545
r146 3 77 182 $w=1.7e-07 $l=4.92874e-07 $layer=licon1_NDIFF $count=1 $X=3.86
+ $Y=0.665 $X2=4.08 $Y2=0.27
r147 2 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.35 $X2=1.12 $Y2=0.56
r148 1 21 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.35 $X2=0.26 $Y2=0.545
.ends

