* File: sky130_fd_sc_lp__a2bb2oi_4.pxi.spice
* Created: Wed Sep  2 09:24:36 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%B1 N_B1_M1002_g N_B1_M1003_g N_B1_M1005_g
+ N_B1_M1013_g N_B1_M1014_g N_B1_M1025_g N_B1_M1035_g N_B1_c_164_n N_B1_M1018_g
+ N_B1_c_166_n N_B1_c_175_n B1 B1 N_B1_c_168_n N_B1_c_169_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_4%B1
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%B2 N_B2_M1000_g N_B2_M1004_g N_B2_M1012_g
+ N_B2_M1010_g N_B2_M1021_g N_B2_M1020_g N_B2_M1034_g N_B2_M1023_g B2 B2 B2
+ N_B2_c_286_n N_B2_c_287_n N_B2_c_288_n B2 PM_SKY130_FD_SC_LP__A2BB2OI_4%B2
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%A_832_21# N_A_832_21#_M1006_d
+ N_A_832_21#_M1022_d N_A_832_21#_M1007_d N_A_832_21#_M1027_d
+ N_A_832_21#_M1009_d N_A_832_21#_M1032_d N_A_832_21#_M1017_g
+ N_A_832_21#_M1001_g N_A_832_21#_M1030_g N_A_832_21#_M1016_g
+ N_A_832_21#_M1031_g N_A_832_21#_M1028_g N_A_832_21#_M1037_g
+ N_A_832_21#_M1036_g N_A_832_21#_c_363_n N_A_832_21#_c_364_n
+ N_A_832_21#_c_526_p N_A_832_21#_c_365_n N_A_832_21#_c_366_n
+ N_A_832_21#_c_534_p N_A_832_21#_c_367_n N_A_832_21#_c_420_p
+ N_A_832_21#_c_535_p N_A_832_21#_c_506_p N_A_832_21#_c_423_p
+ N_A_832_21#_c_379_n N_A_832_21#_c_380_n N_A_832_21#_c_536_p
+ N_A_832_21#_c_509_p N_A_832_21#_c_368_n N_A_832_21#_c_381_n
+ N_A_832_21#_c_369_n N_A_832_21#_c_383_n N_A_832_21#_c_384_n
+ N_A_832_21#_c_370_n N_A_832_21#_c_371_n N_A_832_21#_c_443_p
+ N_A_832_21#_c_372_n N_A_832_21#_c_385_n N_A_832_21#_c_373_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_4%A_832_21#
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%A1_N N_A1_N_M1006_g N_A1_N_M1011_g
+ N_A1_N_M1008_g N_A1_N_M1022_g N_A1_N_M1019_g N_A1_N_M1026_g N_A1_N_M1029_g
+ N_A1_N_M1038_g A1_N A1_N A1_N A1_N N_A1_N_c_557_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_4%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%A2_N N_A2_N_M1007_g N_A2_N_M1009_g
+ N_A2_N_M1024_g N_A2_N_M1015_g N_A2_N_M1027_g N_A2_N_M1032_g N_A2_N_M1039_g
+ N_A2_N_M1033_g A2_N A2_N N_A2_N_c_672_n N_A2_N_c_654_n N_A2_N_c_655_n A2_N
+ PM_SKY130_FD_SC_LP__A2BB2OI_4%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%A_73_367# N_A_73_367#_M1002_d
+ N_A_73_367#_M1005_d N_A_73_367#_M1000_d N_A_73_367#_M1021_d
+ N_A_73_367#_M1018_d N_A_73_367#_M1016_s N_A_73_367#_M1036_s
+ N_A_73_367#_c_728_n N_A_73_367#_c_729_n N_A_73_367#_c_730_n
+ N_A_73_367#_c_776_p N_A_73_367#_c_741_n N_A_73_367#_c_787_p
+ N_A_73_367#_c_744_n N_A_73_367#_c_788_p N_A_73_367#_c_745_n
+ N_A_73_367#_c_747_n N_A_73_367#_c_750_n N_A_73_367#_c_763_n
+ N_A_73_367#_c_751_n N_A_73_367#_c_811_p N_A_73_367#_c_765_n
+ N_A_73_367#_c_731_n N_A_73_367#_c_732_n N_A_73_367#_c_733_n
+ N_A_73_367#_c_756_n N_A_73_367#_c_757_n N_A_73_367#_c_786_p
+ PM_SKY130_FD_SC_LP__A2BB2OI_4%A_73_367#
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%VPWR N_VPWR_M1002_s N_VPWR_M1014_s
+ N_VPWR_M1012_s N_VPWR_M1034_s N_VPWR_M1008_s N_VPWR_M1029_s N_VPWR_c_819_n
+ N_VPWR_c_820_n N_VPWR_c_821_n N_VPWR_c_822_n N_VPWR_c_823_n N_VPWR_c_824_n
+ N_VPWR_c_825_n N_VPWR_c_826_n N_VPWR_c_827_n N_VPWR_c_828_n N_VPWR_c_829_n
+ N_VPWR_c_830_n N_VPWR_c_831_n VPWR N_VPWR_c_832_n N_VPWR_c_833_n
+ N_VPWR_c_834_n N_VPWR_c_818_n N_VPWR_c_836_n N_VPWR_c_837_n N_VPWR_c_838_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%Y N_Y_M1004_d N_Y_M1020_d N_Y_M1017_s
+ N_Y_M1031_s N_Y_M1001_d N_Y_M1028_d N_Y_c_968_n N_Y_c_963_n N_Y_c_1043_p
+ N_Y_c_976_n N_Y_c_964_n N_Y_c_965_n N_Y_c_1000_n N_Y_c_1045_p N_Y_c_1005_n
+ N_Y_c_1009_n Y PM_SKY130_FD_SC_LP__A2BB2OI_4%Y
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%A_1241_367# N_A_1241_367#_M1008_d
+ N_A_1241_367#_M1019_d N_A_1241_367#_M1038_d N_A_1241_367#_M1015_s
+ N_A_1241_367#_M1033_s N_A_1241_367#_c_1059_n N_A_1241_367#_c_1060_n
+ N_A_1241_367#_c_1073_n N_A_1241_367#_c_1101_n N_A_1241_367#_c_1077_n
+ N_A_1241_367#_c_1081_n N_A_1241_367#_c_1105_n N_A_1241_367#_c_1065_n
+ N_A_1241_367#_c_1067_n N_A_1241_367#_c_1068_n N_A_1241_367#_c_1061_n
+ N_A_1241_367#_c_1062_n N_A_1241_367#_c_1082_n N_A_1241_367#_c_1113_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_4%A_1241_367#
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%VGND N_VGND_M1003_d N_VGND_M1013_d
+ N_VGND_M1035_d N_VGND_M1030_d N_VGND_M1037_d N_VGND_M1011_s N_VGND_M1026_s
+ N_VGND_M1024_s N_VGND_M1039_s N_VGND_c_1115_n N_VGND_c_1116_n N_VGND_c_1117_n
+ N_VGND_c_1118_n N_VGND_c_1119_n N_VGND_c_1120_n N_VGND_c_1121_n
+ N_VGND_c_1122_n N_VGND_c_1123_n N_VGND_c_1124_n N_VGND_c_1125_n
+ N_VGND_c_1126_n N_VGND_c_1127_n N_VGND_c_1128_n N_VGND_c_1129_n
+ N_VGND_c_1130_n N_VGND_c_1131_n N_VGND_c_1132_n N_VGND_c_1133_n VGND
+ N_VGND_c_1134_n N_VGND_c_1135_n N_VGND_c_1136_n N_VGND_c_1137_n
+ N_VGND_c_1138_n N_VGND_c_1139_n N_VGND_c_1140_n N_VGND_c_1141_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_4%VGND
x_PM_SKY130_FD_SC_LP__A2BB2OI_4%A_157_47# N_A_157_47#_M1003_s
+ N_A_157_47#_M1025_s N_A_157_47#_M1010_s N_A_157_47#_M1023_s
+ N_A_157_47#_c_1299_n N_A_157_47#_c_1274_n N_A_157_47#_c_1275_n
+ N_A_157_47#_c_1304_n N_A_157_47#_c_1285_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_4%A_157_47#
cc_1 VNB N_B1_M1002_g 0.00233375f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.465
cc_2 VNB N_B1_M1003_g 0.0303807f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.655
cc_3 VNB N_B1_M1005_g 0.00147296f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=2.465
cc_4 VNB N_B1_M1013_g 0.0206884f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.655
cc_5 VNB N_B1_M1014_g 0.00135569f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=2.465
cc_6 VNB N_B1_M1025_g 0.0209252f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=0.655
cc_7 VNB N_B1_M1035_g 0.0186883f $X=-0.19 $Y=-0.245 $X2=3.72 $Y2=0.655
cc_8 VNB N_B1_c_164_n 0.034187f $X=-0.19 $Y=-0.245 $X2=3.875 $Y2=1.54
cc_9 VNB N_B1_M1018_g 0.00579185f $X=-0.19 $Y=-0.245 $X2=3.875 $Y2=2.465
cc_10 VNB N_B1_c_166_n 0.0121355f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.452
cc_11 VNB B1 0.00508327f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.21
cc_12 VNB N_B1_c_168_n 0.042574f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.46
cc_13 VNB N_B1_c_169_n 0.0500674f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=1.46
cc_14 VNB N_B2_M1000_g 0.00463918f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.465
cc_15 VNB N_B2_M1004_g 0.0188931f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.655
cc_16 VNB N_B2_M1012_g 0.00452371f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=2.465
cc_17 VNB N_B2_M1010_g 0.0184678f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.655
cc_18 VNB N_B2_M1021_g 0.00452421f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=2.465
cc_19 VNB N_B2_M1020_g 0.0184723f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=0.655
cc_20 VNB N_B2_M1034_g 0.00510447f $X=-0.19 $Y=-0.245 $X2=3.72 $Y2=0.655
cc_21 VNB N_B2_M1023_g 0.0188574f $X=-0.19 $Y=-0.245 $X2=3.875 $Y2=2.465
cc_22 VNB N_B2_c_286_n 0.00678485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B2_c_287_n 0.0787107f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.46
cc_24 VNB N_B2_c_288_n 9.89949e-19 $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=1.46
cc_25 VNB N_A_832_21#_M1017_g 0.0230011f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=1.295
cc_26 VNB N_A_832_21#_M1030_g 0.0218419f $X=-0.19 $Y=-0.245 $X2=3.875 $Y2=1.54
cc_27 VNB N_A_832_21#_M1031_g 0.0218789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_832_21#_M1037_g 0.0210156f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.75
cc_29 VNB N_A_832_21#_c_363_n 0.00329067f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.46
cc_30 VNB N_A_832_21#_c_364_n 0.00118656f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.46
cc_31 VNB N_A_832_21#_c_365_n 0.00304888f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=1.375
cc_32 VNB N_A_832_21#_c_366_n 0.00487646f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=1.375
cc_33 VNB N_A_832_21#_c_367_n 0.0060272f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=1.375
cc_34 VNB N_A_832_21#_c_368_n 0.0133826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_832_21#_c_369_n 0.0238383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_832_21#_c_370_n 0.00144499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_832_21#_c_371_n 0.00359511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_832_21#_c_372_n 0.00261354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_832_21#_c_373_n 0.0703377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A1_N_M1006_g 0.0224266f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.465
cc_41 VNB N_A1_N_M1011_g 0.0227357f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.655
cc_42 VNB N_A1_N_M1022_g 0.0227528f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.655
cc_43 VNB N_A1_N_M1026_g 0.0304638f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=0.655
cc_44 VNB A1_N 0.003338f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.46
cc_45 VNB N_A1_N_c_557_n 0.0972745f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.46
cc_46 VNB N_A2_N_M1007_g 0.0241499f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.465
cc_47 VNB N_A2_N_M1009_g 0.00256139f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.655
cc_48 VNB N_A2_N_M1024_g 0.020016f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=2.465
cc_49 VNB N_A2_N_M1015_g 0.00249089f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=0.655
cc_50 VNB N_A2_N_M1027_g 0.0205117f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=2.465
cc_51 VNB N_A2_N_M1032_g 0.00249043f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=0.655
cc_52 VNB N_A2_N_M1039_g 0.0236548f $X=-0.19 $Y=-0.245 $X2=3.72 $Y2=0.655
cc_53 VNB N_A2_N_M1033_g 0.00269253f $X=-0.19 $Y=-0.245 $X2=3.875 $Y2=2.465
cc_54 VNB A2_N 0.00214223f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.452
cc_55 VNB N_A2_N_c_654_n 0.0893876f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.46
cc_56 VNB N_A2_N_c_655_n 0.00358962f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.46
cc_57 VNB N_VPWR_c_818_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Y_c_963_n 0.00386207f $X=-0.19 $Y=-0.245 $X2=3.72 $Y2=0.655
cc_59 VNB N_Y_c_964_n 0.00313013f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.46
cc_60 VNB N_Y_c_965_n 0.00212745f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.46
cc_61 VNB Y 0.00460961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1115_n 0.0396521f $X=-0.19 $Y=-0.245 $X2=3.875 $Y2=2.465
cc_63 VNB N_VGND_c_1116_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1117_n 4.06069e-19 $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.46
cc_65 VNB N_VGND_c_1118_n 0.00497428f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.46
cc_66 VNB N_VGND_c_1119_n 3.16879e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1120_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.58
cc_68 VNB N_VGND_c_1121_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1122_n 3.08929e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1123_n 3.1072e-19 $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.46
cc_71 VNB N_VGND_c_1124_n 0.0141935f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.46
cc_72 VNB N_VGND_c_1125_n 0.0261041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1126_n 0.0126445f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=1.375
cc_74 VNB N_VGND_c_1127_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=3.74 $Y2=1.375
cc_75 VNB N_VGND_c_1128_n 0.0523266f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=1.295
cc_76 VNB N_VGND_c_1129_n 0.00632108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1130_n 0.0143903f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=1.375
cc_78 VNB N_VGND_c_1131_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=1.622
cc_79 VNB N_VGND_c_1132_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1133_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1134_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1135_n 0.0131581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1136_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1137_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1138_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1139_n 0.0165581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1140_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1141_n 0.481574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_157_47#_c_1274_n 0.00626045f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.625
cc_90 VNB N_A_157_47#_c_1275_n 0.00317756f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=2.465
cc_91 VPB N_B1_M1002_g 0.0250717f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.465
cc_92 VPB N_B1_M1005_g 0.0186586f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.465
cc_93 VPB N_B1_M1014_g 0.0188208f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=2.465
cc_94 VPB N_B1_M1018_g 0.0210863f $X=-0.19 $Y=1.655 $X2=3.875 $Y2=2.465
cc_95 VPB N_B1_c_166_n 4.21112e-19 $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.452
cc_96 VPB N_B1_c_175_n 0.0224175f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=1.75
cc_97 VPB B1 3.40277e-19 $X=-0.19 $Y=1.655 $X2=3.515 $Y2=1.58
cc_98 VPB N_B2_M1000_g 0.0182009f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.465
cc_99 VPB N_B2_M1012_g 0.0181771f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.465
cc_100 VPB N_B2_M1021_g 0.0181597f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=2.465
cc_101 VPB N_B2_M1034_g 0.020104f $X=-0.19 $Y=1.655 $X2=3.72 $Y2=0.655
cc_102 VPB N_A_832_21#_M1001_g 0.019819f $X=-0.19 $Y=1.655 $X2=3.72 $Y2=1.21
cc_103 VPB N_A_832_21#_M1016_g 0.0192755f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.452
cc_104 VPB N_A_832_21#_M1028_g 0.0192386f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=1.75
cc_105 VPB N_A_832_21#_M1036_g 0.0253127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_832_21#_c_363_n 0.00975558f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.46
cc_107 VPB N_A_832_21#_c_379_n 0.00236792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_832_21#_c_380_n 0.00272206f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_832_21#_c_381_n 0.00968219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_832_21#_c_369_n 0.00191807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_832_21#_c_383_n 0.00381232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_832_21#_c_384_n 0.00139422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_832_21#_c_385_n 0.00209282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_832_21#_c_373_n 0.0103314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A1_N_M1008_g 0.024141f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.465
cc_116 VPB N_A1_N_M1019_g 0.0178969f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=2.465
cc_117 VPB N_A1_N_M1029_g 0.0178969f $X=-0.19 $Y=1.655 $X2=3.72 $Y2=0.655
cc_118 VPB N_A1_N_M1038_g 0.0180878f $X=-0.19 $Y=1.655 $X2=3.875 $Y2=2.465
cc_119 VPB A1_N 0.0131966f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.46
cc_120 VPB N_A1_N_c_557_n 0.0329f $X=-0.19 $Y=1.655 $X2=1.48 $Y2=1.46
cc_121 VPB N_A2_N_M1009_g 0.0195486f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.655
cc_122 VPB N_A2_N_M1015_g 0.0186105f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=0.655
cc_123 VPB N_A2_N_M1032_g 0.0185927f $X=-0.19 $Y=1.655 $X2=1.57 $Y2=0.655
cc_124 VPB N_A2_N_M1033_g 0.0235239f $X=-0.19 $Y=1.655 $X2=3.875 $Y2=2.465
cc_125 VPB N_A_73_367#_c_728_n 0.0446588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_73_367#_c_729_n 0.0031252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_73_367#_c_730_n 0.00903419f $X=-0.19 $Y=1.655 $X2=3.875 $Y2=1.54
cc_128 VPB N_A_73_367#_c_731_n 0.001829f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.46
cc_129 VPB N_A_73_367#_c_732_n 0.00949083f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.46
cc_130 VPB N_A_73_367#_c_733_n 0.00268916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_819_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.57 $Y2=1.295
cc_132 VPB N_VPWR_c_820_n 0.0129398f $X=-0.19 $Y=1.655 $X2=3.72 $Y2=1.21
cc_133 VPB N_VPWR_c_821_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=3.875 $Y2=1.54
cc_134 VPB N_VPWR_c_822_n 3.22457e-19 $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.452
cc_135 VPB N_VPWR_c_823_n 0.0045419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_824_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=3.505 $Y2=1.75
cc_137 VPB N_VPWR_c_825_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.72 $Y2=1.75
cc_138 VPB N_VPWR_c_826_n 0.0226949f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=1.21
cc_139 VPB N_VPWR_c_827_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=1.58
cc_140 VPB N_VPWR_c_828_n 0.0671635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_829_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_830_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.46
cc_143 VPB N_VPWR_c_831_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_832_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.57 $Y2=1.46
cc_145 VPB N_VPWR_c_833_n 0.0164383f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_834_n 0.0549843f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_818_n 0.0661226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_836_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_837_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_838_n 0.00631788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_Y_c_963_n 0.00247048f $X=-0.19 $Y=1.655 $X2=3.72 $Y2=0.655
cc_152 VPB N_A_1241_367#_c_1059_n 0.00202346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_1241_367#_c_1060_n 0.00893455f $X=-0.19 $Y=1.655 $X2=1.565
+ $Y2=2.465
cc_154 VPB N_A_1241_367#_c_1061_n 0.00745909f $X=-0.19 $Y=1.655 $X2=1.48
+ $Y2=1.452
cc_155 VPB N_A_1241_367#_c_1062_n 0.0331155f $X=-0.19 $Y=1.655 $X2=1.48 $Y2=1.46
cc_156 N_B1_M1014_g N_B2_M1000_g 0.0389471f $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_157 N_B1_c_166_n N_B2_M1000_g 2.17836e-19 $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_158 N_B1_c_175_n N_B2_M1000_g 0.0116372f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_159 N_B1_c_169_n N_B2_M1000_g 0.009427f $X=1.57 $Y=1.46 $X2=0 $Y2=0
cc_160 N_B1_M1025_g N_B2_M1004_g 0.0182161f $X=1.57 $Y=0.655 $X2=0 $Y2=0
cc_161 N_B1_c_175_n N_B2_M1012_g 0.0105687f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_162 N_B1_c_175_n N_B2_M1021_g 0.0106152f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_163 N_B1_c_175_n N_B2_M1034_g 0.0116939f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_164 N_B1_M1035_g N_B2_M1023_g 0.0345081f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_165 N_B1_c_164_n N_B2_M1023_g 0.0113432f $X=3.875 $Y=1.54 $X2=0 $Y2=0
cc_166 B1 N_B2_M1023_g 0.00120083f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_167 N_B1_c_164_n N_B2_c_286_n 2.81496e-19 $X=3.875 $Y=1.54 $X2=0 $Y2=0
cc_168 N_B1_c_175_n N_B2_c_286_n 0.0804507f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_169 B1 N_B2_c_286_n 0.0236501f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_170 N_B1_M1025_g N_B2_c_287_n 0.009427f $X=1.57 $Y=0.655 $X2=0 $Y2=0
cc_171 N_B1_c_164_n N_B2_c_287_n 0.00993704f $X=3.875 $Y=1.54 $X2=0 $Y2=0
cc_172 N_B1_M1018_g N_B2_c_287_n 0.0378985f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_173 N_B1_c_166_n N_B2_c_287_n 0.00517446f $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_174 N_B1_c_175_n N_B2_c_287_n 0.007546f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_175 B1 N_B2_c_287_n 0.00528302f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_176 N_B1_M1025_g N_B2_c_288_n 5.77136e-19 $X=1.57 $Y=0.655 $X2=0 $Y2=0
cc_177 N_B1_c_166_n N_B2_c_288_n 0.0103286f $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_178 N_B1_c_175_n N_B2_c_288_n 0.0136253f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_179 N_B1_c_169_n N_B2_c_288_n 3.43472e-19 $X=1.57 $Y=1.46 $X2=0 $Y2=0
cc_180 N_B1_M1035_g N_A_832_21#_M1017_g 0.0229521f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_181 N_B1_c_164_n N_A_832_21#_M1017_g 0.00862923f $X=3.875 $Y=1.54 $X2=0 $Y2=0
cc_182 B1 N_A_832_21#_M1017_g 3.76346e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_183 N_B1_M1018_g N_A_832_21#_M1001_g 0.0323692f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_184 N_B1_c_164_n N_A_832_21#_c_373_n 0.0161016f $X=3.875 $Y=1.54 $X2=0 $Y2=0
cc_185 N_B1_M1002_g N_A_73_367#_c_729_n 0.0144188f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B1_M1005_g N_A_73_367#_c_729_n 0.0127594f $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_187 N_B1_c_166_n N_A_73_367#_c_729_n 0.0473917f $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_188 N_B1_c_168_n N_A_73_367#_c_729_n 0.00107159f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_189 N_B1_c_169_n N_A_73_367#_c_729_n 0.00245668f $X=1.57 $Y=1.46 $X2=0 $Y2=0
cc_190 N_B1_c_166_n N_A_73_367#_c_730_n 0.0212343f $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_191 N_B1_c_168_n N_A_73_367#_c_730_n 0.0065941f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_192 N_B1_M1014_g N_A_73_367#_c_741_n 0.013604f $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_193 N_B1_c_166_n N_A_73_367#_c_741_n 0.0155513f $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_194 N_B1_c_175_n N_A_73_367#_c_741_n 0.0174841f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_195 N_B1_c_175_n N_A_73_367#_c_744_n 0.0385167f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_196 N_B1_c_175_n N_A_73_367#_c_745_n 0.0203099f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_197 B1 N_A_73_367#_c_745_n 7.83599e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_198 N_B1_c_164_n N_A_73_367#_c_747_n 5.53111e-19 $X=3.875 $Y=1.54 $X2=0 $Y2=0
cc_199 N_B1_M1018_g N_A_73_367#_c_747_n 0.0204538f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_200 B1 N_A_73_367#_c_747_n 0.0199509f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_201 N_B1_M1018_g N_A_73_367#_c_750_n 0.00778311f $X=3.875 $Y=2.465 $X2=0
+ $Y2=0
cc_202 N_B1_M1018_g N_A_73_367#_c_751_n 0.00217191f $X=3.875 $Y=2.465 $X2=0
+ $Y2=0
cc_203 N_B1_M1005_g N_A_73_367#_c_733_n 2.39613e-19 $X=1.135 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_B1_M1014_g N_A_73_367#_c_733_n 8.31919e-19 $X=1.565 $Y=2.465 $X2=0
+ $Y2=0
cc_205 N_B1_c_166_n N_A_73_367#_c_733_n 0.0249025f $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_206 N_B1_c_169_n N_A_73_367#_c_733_n 0.00255747f $X=1.57 $Y=1.46 $X2=0 $Y2=0
cc_207 N_B1_c_175_n N_A_73_367#_c_756_n 0.0140367f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_208 N_B1_c_175_n N_A_73_367#_c_757_n 0.0143997f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_209 N_B1_c_166_n N_VPWR_M1014_s 0.00184459f $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_210 B1 N_VPWR_M1034_s 0.00380464f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_211 N_B1_M1002_g N_VPWR_c_819_n 0.0168197f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_212 N_B1_M1005_g N_VPWR_c_819_n 0.014823f $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_213 N_B1_M1014_g N_VPWR_c_819_n 7.04153e-19 $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_214 N_B1_M1005_g N_VPWR_c_820_n 0.00486043f $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_215 N_B1_M1014_g N_VPWR_c_820_n 0.00486043f $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_216 N_B1_M1005_g N_VPWR_c_821_n 6.53615e-19 $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_217 N_B1_M1014_g N_VPWR_c_821_n 0.0129237f $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B1_M1018_g N_VPWR_c_823_n 0.00627696f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_219 N_B1_M1002_g N_VPWR_c_826_n 0.00486043f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_220 N_B1_M1018_g N_VPWR_c_828_n 0.00532251f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_221 N_B1_M1002_g N_VPWR_c_818_n 0.0093368f $X=0.705 $Y=2.465 $X2=0 $Y2=0
cc_222 N_B1_M1005_g N_VPWR_c_818_n 0.00824727f $X=1.135 $Y=2.465 $X2=0 $Y2=0
cc_223 N_B1_M1014_g N_VPWR_c_818_n 0.00824727f $X=1.565 $Y=2.465 $X2=0 $Y2=0
cc_224 N_B1_M1018_g N_VPWR_c_818_n 0.00990847f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_225 N_B1_M1035_g N_Y_c_968_n 0.0169614f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_226 N_B1_c_164_n N_Y_c_968_n 0.00491361f $X=3.875 $Y=1.54 $X2=0 $Y2=0
cc_227 N_B1_c_175_n N_Y_c_968_n 0.00401809f $X=3.505 $Y=1.75 $X2=0 $Y2=0
cc_228 B1 N_Y_c_968_n 0.0227242f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_229 N_B1_M1035_g N_Y_c_963_n 0.00354456f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_230 N_B1_c_164_n N_Y_c_963_n 0.00447991f $X=3.875 $Y=1.54 $X2=0 $Y2=0
cc_231 B1 N_Y_c_963_n 0.0348277f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_232 B1 N_Y_c_963_n 0.0135461f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B1_M1018_g N_Y_c_976_n 6.36367e-19 $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_234 N_B1_M1003_g N_VGND_c_1115_n 0.00702716f $X=0.71 $Y=0.655 $X2=0 $Y2=0
cc_235 N_B1_c_166_n N_VGND_c_1115_n 0.0173953f $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_236 N_B1_c_168_n N_VGND_c_1115_n 0.00684551f $X=0.63 $Y=1.46 $X2=0 $Y2=0
cc_237 N_B1_M1003_g N_VGND_c_1116_n 0.00585385f $X=0.71 $Y=0.655 $X2=0 $Y2=0
cc_238 N_B1_M1013_g N_VGND_c_1116_n 0.00486043f $X=1.14 $Y=0.655 $X2=0 $Y2=0
cc_239 N_B1_M1003_g N_VGND_c_1117_n 6.31647e-19 $X=0.71 $Y=0.655 $X2=0 $Y2=0
cc_240 N_B1_M1013_g N_VGND_c_1117_n 0.0103796f $X=1.14 $Y=0.655 $X2=0 $Y2=0
cc_241 N_B1_M1025_g N_VGND_c_1117_n 0.011457f $X=1.57 $Y=0.655 $X2=0 $Y2=0
cc_242 N_B1_M1035_g N_VGND_c_1118_n 0.00347238f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_243 N_B1_M1025_g N_VGND_c_1128_n 0.00486043f $X=1.57 $Y=0.655 $X2=0 $Y2=0
cc_244 N_B1_M1035_g N_VGND_c_1128_n 0.00441875f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_245 N_B1_M1003_g N_VGND_c_1141_n 0.0116279f $X=0.71 $Y=0.655 $X2=0 $Y2=0
cc_246 N_B1_M1013_g N_VGND_c_1141_n 0.00824727f $X=1.14 $Y=0.655 $X2=0 $Y2=0
cc_247 N_B1_M1025_g N_VGND_c_1141_n 0.0082726f $X=1.57 $Y=0.655 $X2=0 $Y2=0
cc_248 N_B1_M1035_g N_VGND_c_1141_n 0.00627331f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_249 N_B1_M1013_g N_A_157_47#_c_1274_n 0.0132652f $X=1.14 $Y=0.655 $X2=0 $Y2=0
cc_250 N_B1_M1025_g N_A_157_47#_c_1274_n 0.0131569f $X=1.57 $Y=0.655 $X2=0 $Y2=0
cc_251 N_B1_c_166_n N_A_157_47#_c_1274_n 0.0582186f $X=1.635 $Y=1.452 $X2=0
+ $Y2=0
cc_252 N_B1_c_175_n N_A_157_47#_c_1274_n 0.00265181f $X=3.505 $Y=1.75 $X2=0
+ $Y2=0
cc_253 N_B1_c_169_n N_A_157_47#_c_1274_n 0.0024132f $X=1.57 $Y=1.46 $X2=0 $Y2=0
cc_254 N_B1_M1003_g N_A_157_47#_c_1275_n 0.00303715f $X=0.71 $Y=0.655 $X2=0
+ $Y2=0
cc_255 N_B1_c_166_n N_A_157_47#_c_1275_n 0.018788f $X=1.635 $Y=1.452 $X2=0 $Y2=0
cc_256 N_B1_c_169_n N_A_157_47#_c_1275_n 0.00251095f $X=1.57 $Y=1.46 $X2=0 $Y2=0
cc_257 N_B2_M1000_g N_A_73_367#_c_741_n 0.0122738f $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_258 N_B2_M1012_g N_A_73_367#_c_744_n 0.0123204f $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_259 N_B2_M1021_g N_A_73_367#_c_744_n 0.0123204f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_260 N_B2_M1034_g N_A_73_367#_c_745_n 0.021091f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_261 N_B2_M1034_g N_A_73_367#_c_750_n 7.96233e-19 $X=3.285 $Y=2.465 $X2=0
+ $Y2=0
cc_262 N_B2_M1000_g N_VPWR_c_821_n 0.0129672f $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_263 N_B2_M1012_g N_VPWR_c_821_n 6.53615e-19 $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_264 N_B2_M1000_g N_VPWR_c_822_n 6.53615e-19 $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_265 N_B2_M1012_g N_VPWR_c_822_n 0.0130363f $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_266 N_B2_M1021_g N_VPWR_c_822_n 0.0132068f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_267 N_B2_M1034_g N_VPWR_c_822_n 6.68961e-19 $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_268 N_B2_M1034_g N_VPWR_c_823_n 0.00485824f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_269 N_B2_M1000_g N_VPWR_c_832_n 0.00486043f $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_270 N_B2_M1012_g N_VPWR_c_832_n 0.00486043f $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_271 N_B2_M1021_g N_VPWR_c_833_n 0.00486043f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_272 N_B2_M1034_g N_VPWR_c_833_n 0.00585385f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_273 N_B2_M1000_g N_VPWR_c_818_n 0.00824727f $X=1.995 $Y=2.465 $X2=0 $Y2=0
cc_274 N_B2_M1012_g N_VPWR_c_818_n 0.00824727f $X=2.425 $Y=2.465 $X2=0 $Y2=0
cc_275 N_B2_M1021_g N_VPWR_c_818_n 0.00824727f $X=2.855 $Y=2.465 $X2=0 $Y2=0
cc_276 N_B2_M1034_g N_VPWR_c_818_n 0.0111432f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_277 N_B2_M1004_g N_Y_c_968_n 0.00349339f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_278 N_B2_M1010_g N_Y_c_968_n 0.0112456f $X=2.43 $Y=0.655 $X2=0 $Y2=0
cc_279 N_B2_M1020_g N_Y_c_968_n 0.0112456f $X=2.86 $Y=0.655 $X2=0 $Y2=0
cc_280 N_B2_M1023_g N_Y_c_968_n 0.0115875f $X=3.29 $Y=0.655 $X2=0 $Y2=0
cc_281 N_B2_c_286_n N_Y_c_968_n 0.0779176f $X=3.17 $Y=1.4 $X2=0 $Y2=0
cc_282 N_B2_c_287_n N_Y_c_968_n 0.00200533f $X=3.285 $Y=1.4 $X2=0 $Y2=0
cc_283 N_B2_c_288_n N_Y_c_968_n 0.00814247f $X=2.182 $Y=1.342 $X2=0 $Y2=0
cc_284 N_B2_M1004_g N_VGND_c_1117_n 0.00109252f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_285 N_B2_M1004_g N_VGND_c_1128_n 0.00357877f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_286 N_B2_M1010_g N_VGND_c_1128_n 0.00357877f $X=2.43 $Y=0.655 $X2=0 $Y2=0
cc_287 N_B2_M1020_g N_VGND_c_1128_n 0.00357877f $X=2.86 $Y=0.655 $X2=0 $Y2=0
cc_288 N_B2_M1023_g N_VGND_c_1128_n 0.00357877f $X=3.29 $Y=0.655 $X2=0 $Y2=0
cc_289 N_B2_M1004_g N_VGND_c_1141_n 0.00537654f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_290 N_B2_M1010_g N_VGND_c_1141_n 0.0053512f $X=2.43 $Y=0.655 $X2=0 $Y2=0
cc_291 N_B2_M1020_g N_VGND_c_1141_n 0.0053512f $X=2.86 $Y=0.655 $X2=0 $Y2=0
cc_292 N_B2_M1023_g N_VGND_c_1141_n 0.00537654f $X=3.29 $Y=0.655 $X2=0 $Y2=0
cc_293 N_B2_M1004_g N_A_157_47#_c_1274_n 0.00329514f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_294 N_B2_M1004_g N_A_157_47#_c_1285_n 0.0158838f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_295 N_B2_M1010_g N_A_157_47#_c_1285_n 0.0118112f $X=2.43 $Y=0.655 $X2=0 $Y2=0
cc_296 N_B2_M1020_g N_A_157_47#_c_1285_n 0.0118112f $X=2.86 $Y=0.655 $X2=0 $Y2=0
cc_297 N_B2_M1023_g N_A_157_47#_c_1285_n 0.0119021f $X=3.29 $Y=0.655 $X2=0 $Y2=0
cc_298 N_B2_c_288_n N_A_157_47#_c_1285_n 2.56135e-19 $X=2.182 $Y=1.342 $X2=0
+ $Y2=0
cc_299 N_A_832_21#_M1037_g N_A1_N_M1006_g 0.0222502f $X=5.525 $Y=0.655 $X2=0
+ $Y2=0
cc_300 N_A_832_21#_c_364_n N_A1_N_M1006_g 0.00287337f $X=5.965 $Y=1.55 $X2=0
+ $Y2=0
cc_301 N_A_832_21#_c_366_n N_A1_N_M1006_g 0.010615f $X=6.265 $Y=1.15 $X2=0 $Y2=0
cc_302 N_A_832_21#_c_373_n N_A1_N_M1006_g 0.0121012f $X=5.595 $Y=1.49 $X2=0
+ $Y2=0
cc_303 N_A_832_21#_c_364_n N_A1_N_M1011_g 0.00203834f $X=5.965 $Y=1.55 $X2=0
+ $Y2=0
cc_304 N_A_832_21#_c_365_n N_A1_N_M1011_g 0.0141753f $X=6.935 $Y=1.15 $X2=0
+ $Y2=0
cc_305 N_A_832_21#_c_363_n N_A1_N_M1008_g 2.0382e-19 $X=5.88 $Y=1.635 $X2=0
+ $Y2=0
cc_306 N_A_832_21#_c_365_n N_A1_N_M1022_g 0.0141753f $X=6.935 $Y=1.15 $X2=0
+ $Y2=0
cc_307 N_A_832_21#_c_367_n N_A1_N_M1026_g 0.017016f $X=7.87 $Y=1.137 $X2=0 $Y2=0
cc_308 N_A_832_21#_c_371_n N_A1_N_M1026_g 0.00310109f $X=7.955 $Y=0.955 $X2=0
+ $Y2=0
cc_309 N_A_832_21#_c_380_n N_A1_N_M1038_g 5.07515e-19 $X=8.615 $Y=1.785 $X2=0
+ $Y2=0
cc_310 N_A_832_21#_M1036_g A1_N 0.00111363f $X=5.595 $Y=2.465 $X2=0 $Y2=0
cc_311 N_A_832_21#_c_363_n A1_N 0.0147976f $X=5.88 $Y=1.635 $X2=0 $Y2=0
cc_312 N_A_832_21#_c_364_n A1_N 0.0109352f $X=5.965 $Y=1.55 $X2=0 $Y2=0
cc_313 N_A_832_21#_c_366_n A1_N 0.0527857f $X=6.265 $Y=1.15 $X2=0 $Y2=0
cc_314 N_A_832_21#_c_367_n A1_N 0.0562224f $X=7.87 $Y=1.137 $X2=0 $Y2=0
cc_315 N_A_832_21#_c_380_n A1_N 0.00343266f $X=8.615 $Y=1.785 $X2=0 $Y2=0
cc_316 N_A_832_21#_c_370_n A1_N 0.0160892f $X=7.03 $Y=1.137 $X2=0 $Y2=0
cc_317 N_A_832_21#_c_371_n A1_N 0.0140619f $X=7.955 $Y=0.955 $X2=0 $Y2=0
cc_318 N_A_832_21#_M1036_g N_A1_N_c_557_n 0.0121012f $X=5.595 $Y=2.465 $X2=0
+ $Y2=0
cc_319 N_A_832_21#_c_363_n N_A1_N_c_557_n 0.00748794f $X=5.88 $Y=1.635 $X2=0
+ $Y2=0
cc_320 N_A_832_21#_c_364_n N_A1_N_c_557_n 0.0100696f $X=5.965 $Y=1.55 $X2=0
+ $Y2=0
cc_321 N_A_832_21#_c_365_n N_A1_N_c_557_n 0.00282707f $X=6.935 $Y=1.15 $X2=0
+ $Y2=0
cc_322 N_A_832_21#_c_366_n N_A1_N_c_557_n 0.00400953f $X=6.265 $Y=1.15 $X2=0
+ $Y2=0
cc_323 N_A_832_21#_c_367_n N_A1_N_c_557_n 0.0151722f $X=7.87 $Y=1.137 $X2=0
+ $Y2=0
cc_324 N_A_832_21#_c_384_n N_A1_N_c_557_n 5.07268e-19 $X=5.185 $Y=1.552 $X2=0
+ $Y2=0
cc_325 N_A_832_21#_c_370_n N_A1_N_c_557_n 0.00292626f $X=7.03 $Y=1.137 $X2=0
+ $Y2=0
cc_326 N_A_832_21#_c_371_n N_A1_N_c_557_n 0.00112198f $X=7.955 $Y=0.955 $X2=0
+ $Y2=0
cc_327 N_A_832_21#_c_420_p N_A2_N_M1007_g 0.0157862f $X=8.305 $Y=0.955 $X2=0
+ $Y2=0
cc_328 N_A_832_21#_c_371_n N_A2_N_M1007_g 0.00825827f $X=7.955 $Y=0.955 $X2=0
+ $Y2=0
cc_329 N_A_832_21#_c_380_n N_A2_N_M1009_g 0.00344778f $X=8.615 $Y=1.785 $X2=0
+ $Y2=0
cc_330 N_A_832_21#_c_423_p N_A2_N_M1024_g 0.0122129f $X=9.165 $Y=0.955 $X2=0
+ $Y2=0
cc_331 N_A_832_21#_c_379_n N_A2_N_M1015_g 0.0149389f $X=9.215 $Y=1.785 $X2=0
+ $Y2=0
cc_332 N_A_832_21#_c_423_p N_A2_N_M1027_g 0.0130197f $X=9.165 $Y=0.955 $X2=0
+ $Y2=0
cc_333 N_A_832_21#_c_372_n N_A2_N_M1027_g 0.00250412f $X=9.265 $Y=0.955 $X2=0
+ $Y2=0
cc_334 N_A_832_21#_c_379_n N_A2_N_M1032_g 0.0149141f $X=9.215 $Y=1.785 $X2=0
+ $Y2=0
cc_335 N_A_832_21#_c_368_n N_A2_N_M1039_g 0.0142666f $X=9.73 $Y=1.09 $X2=0 $Y2=0
cc_336 N_A_832_21#_c_369_n N_A2_N_M1039_g 0.00346516f $X=9.832 $Y=1.695 $X2=0
+ $Y2=0
cc_337 N_A_832_21#_c_372_n N_A2_N_M1039_g 2.17608e-19 $X=9.265 $Y=0.955 $X2=0
+ $Y2=0
cc_338 N_A_832_21#_c_381_n N_A2_N_M1033_g 0.0170416f $X=9.73 $Y=1.785 $X2=0
+ $Y2=0
cc_339 N_A_832_21#_c_423_p N_A2_N_c_672_n 0.00742672f $X=9.165 $Y=0.955 $X2=0
+ $Y2=0
cc_340 N_A_832_21#_c_368_n N_A2_N_c_672_n 0.0134448f $X=9.73 $Y=1.09 $X2=0 $Y2=0
cc_341 N_A_832_21#_c_381_n N_A2_N_c_672_n 0.00579321f $X=9.73 $Y=1.785 $X2=0
+ $Y2=0
cc_342 N_A_832_21#_c_369_n N_A2_N_c_672_n 0.0144179f $X=9.832 $Y=1.695 $X2=0
+ $Y2=0
cc_343 N_A_832_21#_c_372_n N_A2_N_c_672_n 0.0159884f $X=9.265 $Y=0.955 $X2=0
+ $Y2=0
cc_344 N_A_832_21#_c_385_n N_A2_N_c_672_n 0.0210583f $X=9.345 $Y=1.785 $X2=0
+ $Y2=0
cc_345 N_A_832_21#_c_423_p N_A2_N_c_654_n 6.05796e-19 $X=9.165 $Y=0.955 $X2=0
+ $Y2=0
cc_346 N_A_832_21#_c_379_n N_A2_N_c_654_n 0.00276902f $X=9.215 $Y=1.785 $X2=0
+ $Y2=0
cc_347 N_A_832_21#_c_380_n N_A2_N_c_654_n 0.00286879f $X=8.615 $Y=1.785 $X2=0
+ $Y2=0
cc_348 N_A_832_21#_c_368_n N_A2_N_c_654_n 0.00229216f $X=9.73 $Y=1.09 $X2=0
+ $Y2=0
cc_349 N_A_832_21#_c_369_n N_A2_N_c_654_n 0.0154035f $X=9.832 $Y=1.695 $X2=0
+ $Y2=0
cc_350 N_A_832_21#_c_443_p N_A2_N_c_654_n 6.63344e-19 $X=8.405 $Y=0.955 $X2=0
+ $Y2=0
cc_351 N_A_832_21#_c_372_n N_A2_N_c_654_n 0.00283411f $X=9.265 $Y=0.955 $X2=0
+ $Y2=0
cc_352 N_A_832_21#_c_385_n N_A2_N_c_654_n 0.00286879f $X=9.345 $Y=1.785 $X2=0
+ $Y2=0
cc_353 N_A_832_21#_c_420_p N_A2_N_c_655_n 0.00568189f $X=8.305 $Y=0.955 $X2=0
+ $Y2=0
cc_354 N_A_832_21#_c_423_p N_A2_N_c_655_n 0.0294415f $X=9.165 $Y=0.955 $X2=0
+ $Y2=0
cc_355 N_A_832_21#_c_379_n N_A2_N_c_655_n 0.0430879f $X=9.215 $Y=1.785 $X2=0
+ $Y2=0
cc_356 N_A_832_21#_c_380_n N_A2_N_c_655_n 0.0231206f $X=8.615 $Y=1.785 $X2=0
+ $Y2=0
cc_357 N_A_832_21#_c_371_n N_A2_N_c_655_n 0.00191778f $X=7.955 $Y=0.955 $X2=0
+ $Y2=0
cc_358 N_A_832_21#_c_443_p N_A2_N_c_655_n 0.0157534f $X=8.405 $Y=0.955 $X2=0
+ $Y2=0
cc_359 N_A_832_21#_M1001_g N_A_73_367#_c_763_n 0.0115031f $X=4.305 $Y=2.465
+ $X2=0 $Y2=0
cc_360 N_A_832_21#_M1016_g N_A_73_367#_c_763_n 0.0115031f $X=4.735 $Y=2.465
+ $X2=0 $Y2=0
cc_361 N_A_832_21#_M1028_g N_A_73_367#_c_765_n 0.0115031f $X=5.165 $Y=2.465
+ $X2=0 $Y2=0
cc_362 N_A_832_21#_M1036_g N_A_73_367#_c_765_n 0.0115031f $X=5.595 $Y=2.465
+ $X2=0 $Y2=0
cc_363 N_A_832_21#_c_363_n N_A_73_367#_c_732_n 0.0215235f $X=5.88 $Y=1.635 $X2=0
+ $Y2=0
cc_364 N_A_832_21#_M1001_g N_VPWR_c_828_n 0.00357877f $X=4.305 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_A_832_21#_M1016_g N_VPWR_c_828_n 0.00357877f $X=4.735 $Y=2.465 $X2=0
+ $Y2=0
cc_366 N_A_832_21#_M1028_g N_VPWR_c_828_n 0.00357877f $X=5.165 $Y=2.465 $X2=0
+ $Y2=0
cc_367 N_A_832_21#_M1036_g N_VPWR_c_828_n 0.00357877f $X=5.595 $Y=2.465 $X2=0
+ $Y2=0
cc_368 N_A_832_21#_M1009_d N_VPWR_c_818_n 0.00224381f $X=8.34 $Y=1.835 $X2=0
+ $Y2=0
cc_369 N_A_832_21#_M1032_d N_VPWR_c_818_n 0.00225186f $X=9.2 $Y=1.835 $X2=0
+ $Y2=0
cc_370 N_A_832_21#_M1001_g N_VPWR_c_818_n 0.00537654f $X=4.305 $Y=2.465 $X2=0
+ $Y2=0
cc_371 N_A_832_21#_M1016_g N_VPWR_c_818_n 0.0053512f $X=4.735 $Y=2.465 $X2=0
+ $Y2=0
cc_372 N_A_832_21#_M1028_g N_VPWR_c_818_n 0.0053512f $X=5.165 $Y=2.465 $X2=0
+ $Y2=0
cc_373 N_A_832_21#_M1036_g N_VPWR_c_818_n 0.00665089f $X=5.595 $Y=2.465 $X2=0
+ $Y2=0
cc_374 N_A_832_21#_M1017_g N_Y_c_963_n 0.00588823f $X=4.235 $Y=0.655 $X2=0 $Y2=0
cc_375 N_A_832_21#_M1001_g N_Y_c_963_n 0.00442826f $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_376 N_A_832_21#_M1030_g N_Y_c_963_n 6.27328e-19 $X=4.665 $Y=0.655 $X2=0 $Y2=0
cc_377 N_A_832_21#_c_383_n N_Y_c_963_n 0.0251635f $X=4.94 $Y=1.552 $X2=0 $Y2=0
cc_378 N_A_832_21#_c_373_n N_Y_c_963_n 0.00854596f $X=5.595 $Y=1.49 $X2=0 $Y2=0
cc_379 N_A_832_21#_M1001_g N_Y_c_976_n 0.00846541f $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A_832_21#_M1016_g N_Y_c_976_n 0.00821665f $X=4.735 $Y=2.465 $X2=0 $Y2=0
cc_381 N_A_832_21#_M1028_g N_Y_c_976_n 5.71429e-19 $X=5.165 $Y=2.465 $X2=0 $Y2=0
cc_382 N_A_832_21#_M1030_g N_Y_c_964_n 0.0135632f $X=4.665 $Y=0.655 $X2=0 $Y2=0
cc_383 N_A_832_21#_M1031_g N_Y_c_964_n 0.0138595f $X=5.095 $Y=0.655 $X2=0 $Y2=0
cc_384 N_A_832_21#_c_363_n N_Y_c_964_n 0.0012536f $X=5.88 $Y=1.635 $X2=0 $Y2=0
cc_385 N_A_832_21#_c_383_n N_Y_c_964_n 0.0469263f $X=4.94 $Y=1.552 $X2=0 $Y2=0
cc_386 N_A_832_21#_c_373_n N_Y_c_964_n 0.00270092f $X=5.595 $Y=1.49 $X2=0 $Y2=0
cc_387 N_A_832_21#_M1017_g N_Y_c_965_n 0.0166544f $X=4.235 $Y=0.655 $X2=0 $Y2=0
cc_388 N_A_832_21#_c_383_n N_Y_c_965_n 0.0168679f $X=4.94 $Y=1.552 $X2=0 $Y2=0
cc_389 N_A_832_21#_c_373_n N_Y_c_965_n 0.00279997f $X=5.595 $Y=1.49 $X2=0 $Y2=0
cc_390 N_A_832_21#_M1016_g N_Y_c_1000_n 0.00531166f $X=4.735 $Y=2.465 $X2=0
+ $Y2=0
cc_391 N_A_832_21#_M1028_g N_Y_c_1000_n 0.0118386f $X=5.165 $Y=2.465 $X2=0 $Y2=0
cc_392 N_A_832_21#_c_383_n N_Y_c_1000_n 0.0106959f $X=4.94 $Y=1.552 $X2=0 $Y2=0
cc_393 N_A_832_21#_c_384_n N_Y_c_1000_n 0.0185548f $X=5.185 $Y=1.552 $X2=0 $Y2=0
cc_394 N_A_832_21#_c_373_n N_Y_c_1000_n 6.14176e-19 $X=5.595 $Y=1.49 $X2=0 $Y2=0
cc_395 N_A_832_21#_M1001_g N_Y_c_1005_n 0.0157034f $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_396 N_A_832_21#_M1016_g N_Y_c_1005_n 0.00748343f $X=4.735 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_A_832_21#_c_383_n N_Y_c_1005_n 0.0289674f $X=4.94 $Y=1.552 $X2=0 $Y2=0
cc_398 N_A_832_21#_c_373_n N_Y_c_1005_n 0.00224921f $X=5.595 $Y=1.49 $X2=0 $Y2=0
cc_399 N_A_832_21#_M1016_g N_Y_c_1009_n 5.70646e-19 $X=4.735 $Y=2.465 $X2=0
+ $Y2=0
cc_400 N_A_832_21#_M1028_g N_Y_c_1009_n 0.0113838f $X=5.165 $Y=2.465 $X2=0 $Y2=0
cc_401 N_A_832_21#_M1036_g N_Y_c_1009_n 0.0121432f $X=5.595 $Y=2.465 $X2=0 $Y2=0
cc_402 N_A_832_21#_c_363_n N_Y_c_1009_n 0.021761f $X=5.88 $Y=1.635 $X2=0 $Y2=0
cc_403 N_A_832_21#_c_373_n N_Y_c_1009_n 6.63344e-19 $X=5.595 $Y=1.49 $X2=0 $Y2=0
cc_404 N_A_832_21#_M1031_g Y 0.00256815f $X=5.095 $Y=0.655 $X2=0 $Y2=0
cc_405 N_A_832_21#_M1037_g Y 0.0142577f $X=5.525 $Y=0.655 $X2=0 $Y2=0
cc_406 N_A_832_21#_c_363_n Y 0.032077f $X=5.88 $Y=1.635 $X2=0 $Y2=0
cc_407 N_A_832_21#_c_364_n Y 0.0105456f $X=5.965 $Y=1.55 $X2=0 $Y2=0
cc_408 N_A_832_21#_c_366_n Y 0.0142421f $X=6.265 $Y=1.15 $X2=0 $Y2=0
cc_409 N_A_832_21#_c_373_n Y 0.0133003f $X=5.595 $Y=1.49 $X2=0 $Y2=0
cc_410 N_A_832_21#_c_379_n N_A_1241_367#_M1015_s 0.00176773f $X=9.215 $Y=1.785
+ $X2=0 $Y2=0
cc_411 N_A_832_21#_c_381_n N_A_1241_367#_M1033_s 0.00246138f $X=9.73 $Y=1.785
+ $X2=0 $Y2=0
cc_412 N_A_832_21#_M1009_d N_A_1241_367#_c_1065_n 0.00332344f $X=8.34 $Y=1.835
+ $X2=0 $Y2=0
cc_413 N_A_832_21#_c_506_p N_A_1241_367#_c_1065_n 0.0126348f $X=8.48 $Y=1.98
+ $X2=0 $Y2=0
cc_414 N_A_832_21#_c_379_n N_A_1241_367#_c_1067_n 0.0135577f $X=9.215 $Y=1.785
+ $X2=0 $Y2=0
cc_415 N_A_832_21#_M1032_d N_A_1241_367#_c_1068_n 0.00332344f $X=9.2 $Y=1.835
+ $X2=0 $Y2=0
cc_416 N_A_832_21#_c_509_p N_A_1241_367#_c_1068_n 0.0126348f $X=9.34 $Y=1.98
+ $X2=0 $Y2=0
cc_417 N_A_832_21#_c_381_n N_A_1241_367#_c_1062_n 0.022006f $X=9.73 $Y=1.785
+ $X2=0 $Y2=0
cc_418 N_A_832_21#_c_365_n N_VGND_M1011_s 0.00176461f $X=6.935 $Y=1.15 $X2=0
+ $Y2=0
cc_419 N_A_832_21#_c_367_n N_VGND_M1026_s 0.00705089f $X=7.87 $Y=1.137 $X2=0
+ $Y2=0
cc_420 N_A_832_21#_c_420_p N_VGND_M1026_s 0.00161883f $X=8.305 $Y=0.955 $X2=0
+ $Y2=0
cc_421 N_A_832_21#_c_371_n N_VGND_M1026_s 0.00624606f $X=7.955 $Y=0.955 $X2=0
+ $Y2=0
cc_422 N_A_832_21#_c_423_p N_VGND_M1024_s 0.003325f $X=9.165 $Y=0.955 $X2=0
+ $Y2=0
cc_423 N_A_832_21#_c_368_n N_VGND_M1039_s 0.00257121f $X=9.73 $Y=1.09 $X2=0
+ $Y2=0
cc_424 N_A_832_21#_M1017_g N_VGND_c_1118_n 0.00191339f $X=4.235 $Y=0.655 $X2=0
+ $Y2=0
cc_425 N_A_832_21#_M1017_g N_VGND_c_1119_n 6.09599e-19 $X=4.235 $Y=0.655 $X2=0
+ $Y2=0
cc_426 N_A_832_21#_M1030_g N_VGND_c_1119_n 0.0109519f $X=4.665 $Y=0.655 $X2=0
+ $Y2=0
cc_427 N_A_832_21#_M1031_g N_VGND_c_1119_n 0.0108513f $X=5.095 $Y=0.655 $X2=0
+ $Y2=0
cc_428 N_A_832_21#_M1037_g N_VGND_c_1119_n 6.22495e-19 $X=5.525 $Y=0.655 $X2=0
+ $Y2=0
cc_429 N_A_832_21#_M1031_g N_VGND_c_1120_n 6.25324e-19 $X=5.095 $Y=0.655 $X2=0
+ $Y2=0
cc_430 N_A_832_21#_M1037_g N_VGND_c_1120_n 0.0110149f $X=5.525 $Y=0.655 $X2=0
+ $Y2=0
cc_431 N_A_832_21#_c_363_n N_VGND_c_1120_n 0.00452069f $X=5.88 $Y=1.635 $X2=0
+ $Y2=0
cc_432 N_A_832_21#_c_366_n N_VGND_c_1120_n 0.00163297f $X=6.265 $Y=1.15 $X2=0
+ $Y2=0
cc_433 N_A_832_21#_c_526_p N_VGND_c_1121_n 0.0124525f $X=6.17 $Y=0.59 $X2=0
+ $Y2=0
cc_434 N_A_832_21#_c_365_n N_VGND_c_1122_n 0.0170777f $X=6.935 $Y=1.15 $X2=0
+ $Y2=0
cc_435 N_A_832_21#_c_423_p N_VGND_c_1123_n 0.0170777f $X=9.165 $Y=0.955 $X2=0
+ $Y2=0
cc_436 N_A_832_21#_c_368_n N_VGND_c_1125_n 0.0231627f $X=9.73 $Y=1.09 $X2=0
+ $Y2=0
cc_437 N_A_832_21#_M1017_g N_VGND_c_1130_n 0.00441743f $X=4.235 $Y=0.655 $X2=0
+ $Y2=0
cc_438 N_A_832_21#_M1030_g N_VGND_c_1130_n 0.00486043f $X=4.665 $Y=0.655 $X2=0
+ $Y2=0
cc_439 N_A_832_21#_M1031_g N_VGND_c_1132_n 0.00486043f $X=5.095 $Y=0.655 $X2=0
+ $Y2=0
cc_440 N_A_832_21#_M1037_g N_VGND_c_1132_n 0.00486043f $X=5.525 $Y=0.655 $X2=0
+ $Y2=0
cc_441 N_A_832_21#_c_534_p N_VGND_c_1134_n 0.0124525f $X=7.03 $Y=0.42 $X2=0
+ $Y2=0
cc_442 N_A_832_21#_c_535_p N_VGND_c_1135_n 0.0128073f $X=8.41 $Y=0.42 $X2=0
+ $Y2=0
cc_443 N_A_832_21#_c_536_p N_VGND_c_1136_n 0.0124525f $X=9.27 $Y=0.42 $X2=0
+ $Y2=0
cc_444 N_A_832_21#_c_367_n N_VGND_c_1139_n 0.0343065f $X=7.87 $Y=1.137 $X2=0
+ $Y2=0
cc_445 N_A_832_21#_c_420_p N_VGND_c_1139_n 0.00297175f $X=8.305 $Y=0.955 $X2=0
+ $Y2=0
cc_446 N_A_832_21#_c_371_n N_VGND_c_1139_n 0.0144796f $X=7.955 $Y=0.955 $X2=0
+ $Y2=0
cc_447 N_A_832_21#_M1006_d N_VGND_c_1141_n 0.00545212f $X=6.03 $Y=0.235 $X2=0
+ $Y2=0
cc_448 N_A_832_21#_M1022_d N_VGND_c_1141_n 0.00536646f $X=6.89 $Y=0.235 $X2=0
+ $Y2=0
cc_449 N_A_832_21#_M1007_d N_VGND_c_1141_n 0.00501859f $X=8.27 $Y=0.235 $X2=0
+ $Y2=0
cc_450 N_A_832_21#_M1027_d N_VGND_c_1141_n 0.00536646f $X=9.13 $Y=0.235 $X2=0
+ $Y2=0
cc_451 N_A_832_21#_M1017_g N_VGND_c_1141_n 0.00625916f $X=4.235 $Y=0.655 $X2=0
+ $Y2=0
cc_452 N_A_832_21#_M1030_g N_VGND_c_1141_n 0.00824727f $X=4.665 $Y=0.655 $X2=0
+ $Y2=0
cc_453 N_A_832_21#_M1031_g N_VGND_c_1141_n 0.00824727f $X=5.095 $Y=0.655 $X2=0
+ $Y2=0
cc_454 N_A_832_21#_M1037_g N_VGND_c_1141_n 0.00824727f $X=5.525 $Y=0.655 $X2=0
+ $Y2=0
cc_455 N_A_832_21#_c_526_p N_VGND_c_1141_n 0.00730901f $X=6.17 $Y=0.59 $X2=0
+ $Y2=0
cc_456 N_A_832_21#_c_534_p N_VGND_c_1141_n 0.00730901f $X=7.03 $Y=0.42 $X2=0
+ $Y2=0
cc_457 N_A_832_21#_c_535_p N_VGND_c_1141_n 0.00769778f $X=8.41 $Y=0.42 $X2=0
+ $Y2=0
cc_458 N_A_832_21#_c_536_p N_VGND_c_1141_n 0.00730901f $X=9.27 $Y=0.42 $X2=0
+ $Y2=0
cc_459 A1_N N_A2_N_M1009_g 0.00305234f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_460 N_A1_N_c_557_n N_A2_N_M1009_g 0.0204653f $X=7.835 $Y=1.51 $X2=0 $Y2=0
cc_461 A1_N N_A2_N_c_654_n 0.00347148f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_462 N_A1_N_c_557_n N_A2_N_c_654_n 0.0178008f $X=7.835 $Y=1.51 $X2=0 $Y2=0
cc_463 A1_N N_A2_N_c_655_n 0.010519f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_464 N_A1_N_c_557_n N_A2_N_c_655_n 4.76398e-19 $X=7.835 $Y=1.51 $X2=0 $Y2=0
cc_465 N_A1_N_M1008_g N_A_73_367#_c_732_n 6.65533e-19 $X=6.545 $Y=2.465 $X2=0
+ $Y2=0
cc_466 N_A1_N_c_557_n N_A_73_367#_c_732_n 6.51314e-19 $X=7.835 $Y=1.51 $X2=0
+ $Y2=0
cc_467 N_A1_N_M1008_g N_VPWR_c_824_n 0.0168028f $X=6.545 $Y=2.465 $X2=0 $Y2=0
cc_468 N_A1_N_M1019_g N_VPWR_c_824_n 0.0149184f $X=6.975 $Y=2.465 $X2=0 $Y2=0
cc_469 N_A1_N_M1029_g N_VPWR_c_824_n 6.77662e-19 $X=7.405 $Y=2.465 $X2=0 $Y2=0
cc_470 N_A1_N_M1019_g N_VPWR_c_825_n 6.77662e-19 $X=6.975 $Y=2.465 $X2=0 $Y2=0
cc_471 N_A1_N_M1029_g N_VPWR_c_825_n 0.0146776f $X=7.405 $Y=2.465 $X2=0 $Y2=0
cc_472 N_A1_N_M1038_g N_VPWR_c_825_n 0.0158505f $X=7.835 $Y=2.465 $X2=0 $Y2=0
cc_473 N_A1_N_M1008_g N_VPWR_c_828_n 0.00486043f $X=6.545 $Y=2.465 $X2=0 $Y2=0
cc_474 N_A1_N_M1019_g N_VPWR_c_830_n 0.00486043f $X=6.975 $Y=2.465 $X2=0 $Y2=0
cc_475 N_A1_N_M1029_g N_VPWR_c_830_n 0.00486043f $X=7.405 $Y=2.465 $X2=0 $Y2=0
cc_476 N_A1_N_M1038_g N_VPWR_c_834_n 0.00486043f $X=7.835 $Y=2.465 $X2=0 $Y2=0
cc_477 N_A1_N_M1008_g N_VPWR_c_818_n 0.00954696f $X=6.545 $Y=2.465 $X2=0 $Y2=0
cc_478 N_A1_N_M1019_g N_VPWR_c_818_n 0.00824727f $X=6.975 $Y=2.465 $X2=0 $Y2=0
cc_479 N_A1_N_M1029_g N_VPWR_c_818_n 0.00824727f $X=7.405 $Y=2.465 $X2=0 $Y2=0
cc_480 N_A1_N_M1038_g N_VPWR_c_818_n 0.0082726f $X=7.835 $Y=2.465 $X2=0 $Y2=0
cc_481 N_A1_N_M1006_g Y 0.00176992f $X=5.955 $Y=0.655 $X2=0 $Y2=0
cc_482 A1_N N_A_1241_367#_c_1059_n 0.0169473f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_483 N_A1_N_c_557_n N_A_1241_367#_c_1059_n 0.00350654f $X=7.835 $Y=1.51 $X2=0
+ $Y2=0
cc_484 N_A1_N_M1008_g N_A_1241_367#_c_1073_n 0.01229f $X=6.545 $Y=2.465 $X2=0
+ $Y2=0
cc_485 N_A1_N_M1019_g N_A_1241_367#_c_1073_n 0.01229f $X=6.975 $Y=2.465 $X2=0
+ $Y2=0
cc_486 A1_N N_A_1241_367#_c_1073_n 0.0420923f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_487 N_A1_N_c_557_n N_A_1241_367#_c_1073_n 5.62401e-19 $X=7.835 $Y=1.51 $X2=0
+ $Y2=0
cc_488 N_A1_N_M1029_g N_A_1241_367#_c_1077_n 0.0122435f $X=7.405 $Y=2.465 $X2=0
+ $Y2=0
cc_489 N_A1_N_M1038_g N_A_1241_367#_c_1077_n 0.01229f $X=7.835 $Y=2.465 $X2=0
+ $Y2=0
cc_490 A1_N N_A_1241_367#_c_1077_n 0.0420923f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_491 N_A1_N_c_557_n N_A_1241_367#_c_1077_n 5.69728e-19 $X=7.835 $Y=1.51 $X2=0
+ $Y2=0
cc_492 A1_N N_A_1241_367#_c_1081_n 0.00671851f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_493 A1_N N_A_1241_367#_c_1082_n 0.0151418f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_494 N_A1_N_c_557_n N_A_1241_367#_c_1082_n 6.37626e-19 $X=7.835 $Y=1.51 $X2=0
+ $Y2=0
cc_495 N_A1_N_M1006_g N_VGND_c_1120_n 0.0110358f $X=5.955 $Y=0.655 $X2=0 $Y2=0
cc_496 N_A1_N_M1011_g N_VGND_c_1120_n 6.61513e-19 $X=6.385 $Y=0.655 $X2=0 $Y2=0
cc_497 N_A1_N_M1006_g N_VGND_c_1121_n 0.00486043f $X=5.955 $Y=0.655 $X2=0 $Y2=0
cc_498 N_A1_N_M1011_g N_VGND_c_1121_n 0.00486043f $X=6.385 $Y=0.655 $X2=0 $Y2=0
cc_499 N_A1_N_M1006_g N_VGND_c_1122_n 6.67171e-19 $X=5.955 $Y=0.655 $X2=0 $Y2=0
cc_500 N_A1_N_M1011_g N_VGND_c_1122_n 0.0107833f $X=6.385 $Y=0.655 $X2=0 $Y2=0
cc_501 N_A1_N_M1022_g N_VGND_c_1122_n 0.0107809f $X=6.815 $Y=0.655 $X2=0 $Y2=0
cc_502 N_A1_N_M1026_g N_VGND_c_1122_n 6.30572e-19 $X=7.245 $Y=0.655 $X2=0 $Y2=0
cc_503 N_A1_N_M1022_g N_VGND_c_1134_n 0.00486043f $X=6.815 $Y=0.655 $X2=0 $Y2=0
cc_504 N_A1_N_M1026_g N_VGND_c_1134_n 0.00486043f $X=7.245 $Y=0.655 $X2=0 $Y2=0
cc_505 N_A1_N_M1022_g N_VGND_c_1139_n 6.40525e-19 $X=6.815 $Y=0.655 $X2=0 $Y2=0
cc_506 N_A1_N_M1026_g N_VGND_c_1139_n 0.0130128f $X=7.245 $Y=0.655 $X2=0 $Y2=0
cc_507 N_A1_N_c_557_n N_VGND_c_1139_n 6.87646e-19 $X=7.835 $Y=1.51 $X2=0 $Y2=0
cc_508 N_A1_N_M1006_g N_VGND_c_1141_n 0.00835506f $X=5.955 $Y=0.655 $X2=0 $Y2=0
cc_509 N_A1_N_M1011_g N_VGND_c_1141_n 0.00835506f $X=6.385 $Y=0.655 $X2=0 $Y2=0
cc_510 N_A1_N_M1022_g N_VGND_c_1141_n 0.00824727f $X=6.815 $Y=0.655 $X2=0 $Y2=0
cc_511 N_A1_N_M1026_g N_VGND_c_1141_n 0.00819843f $X=7.245 $Y=0.655 $X2=0 $Y2=0
cc_512 N_A2_N_M1009_g N_VPWR_c_825_n 0.00109252f $X=8.265 $Y=2.465 $X2=0 $Y2=0
cc_513 N_A2_N_M1009_g N_VPWR_c_834_n 0.00357877f $X=8.265 $Y=2.465 $X2=0 $Y2=0
cc_514 N_A2_N_M1015_g N_VPWR_c_834_n 0.00357877f $X=8.695 $Y=2.465 $X2=0 $Y2=0
cc_515 N_A2_N_M1032_g N_VPWR_c_834_n 0.00357877f $X=9.125 $Y=2.465 $X2=0 $Y2=0
cc_516 N_A2_N_M1033_g N_VPWR_c_834_n 0.00357877f $X=9.555 $Y=2.465 $X2=0 $Y2=0
cc_517 N_A2_N_M1009_g N_VPWR_c_818_n 0.00537654f $X=8.265 $Y=2.465 $X2=0 $Y2=0
cc_518 N_A2_N_M1015_g N_VPWR_c_818_n 0.0053512f $X=8.695 $Y=2.465 $X2=0 $Y2=0
cc_519 N_A2_N_M1032_g N_VPWR_c_818_n 0.0053512f $X=9.125 $Y=2.465 $X2=0 $Y2=0
cc_520 N_A2_N_M1033_g N_VPWR_c_818_n 0.00632779f $X=9.555 $Y=2.465 $X2=0 $Y2=0
cc_521 N_A2_N_c_654_n N_A_1241_367#_c_1081_n 0.00129197f $X=9.555 $Y=1.44 $X2=0
+ $Y2=0
cc_522 N_A2_N_M1009_g N_A_1241_367#_c_1065_n 0.012237f $X=8.265 $Y=2.465 $X2=0
+ $Y2=0
cc_523 N_A2_N_M1015_g N_A_1241_367#_c_1065_n 0.0121905f $X=8.695 $Y=2.465 $X2=0
+ $Y2=0
cc_524 N_A2_N_M1032_g N_A_1241_367#_c_1068_n 0.012237f $X=9.125 $Y=2.465 $X2=0
+ $Y2=0
cc_525 N_A2_N_M1033_g N_A_1241_367#_c_1068_n 0.012237f $X=9.555 $Y=2.465 $X2=0
+ $Y2=0
cc_526 N_A2_N_M1007_g N_VGND_c_1123_n 5.79502e-19 $X=8.195 $Y=0.655 $X2=0 $Y2=0
cc_527 N_A2_N_M1024_g N_VGND_c_1123_n 0.0101098f $X=8.625 $Y=0.655 $X2=0 $Y2=0
cc_528 N_A2_N_M1027_g N_VGND_c_1123_n 0.0100888f $X=9.055 $Y=0.655 $X2=0 $Y2=0
cc_529 N_A2_N_M1039_g N_VGND_c_1123_n 5.75816e-19 $X=9.485 $Y=0.655 $X2=0 $Y2=0
cc_530 N_A2_N_M1027_g N_VGND_c_1125_n 6.14008e-19 $X=9.055 $Y=0.655 $X2=0 $Y2=0
cc_531 N_A2_N_M1039_g N_VGND_c_1125_n 0.0112405f $X=9.485 $Y=0.655 $X2=0 $Y2=0
cc_532 N_A2_N_M1007_g N_VGND_c_1135_n 0.00525069f $X=8.195 $Y=0.655 $X2=0 $Y2=0
cc_533 N_A2_N_M1024_g N_VGND_c_1135_n 0.00486043f $X=8.625 $Y=0.655 $X2=0 $Y2=0
cc_534 N_A2_N_M1027_g N_VGND_c_1136_n 0.00486043f $X=9.055 $Y=0.655 $X2=0 $Y2=0
cc_535 N_A2_N_M1039_g N_VGND_c_1136_n 0.00486043f $X=9.485 $Y=0.655 $X2=0 $Y2=0
cc_536 N_A2_N_M1007_g N_VGND_c_1139_n 0.0164209f $X=8.195 $Y=0.655 $X2=0 $Y2=0
cc_537 N_A2_N_M1024_g N_VGND_c_1139_n 5.8213e-19 $X=8.625 $Y=0.655 $X2=0 $Y2=0
cc_538 N_A2_N_M1007_g N_VGND_c_1141_n 0.00881625f $X=8.195 $Y=0.655 $X2=0 $Y2=0
cc_539 N_A2_N_M1024_g N_VGND_c_1141_n 0.00824727f $X=8.625 $Y=0.655 $X2=0 $Y2=0
cc_540 N_A2_N_M1027_g N_VGND_c_1141_n 0.00824727f $X=9.055 $Y=0.655 $X2=0 $Y2=0
cc_541 N_A2_N_M1039_g N_VGND_c_1141_n 0.00824727f $X=9.485 $Y=0.655 $X2=0 $Y2=0
cc_542 N_A_73_367#_c_729_n N_VPWR_M1002_s 0.00176461f $X=1.255 $Y=1.81 $X2=-0.19
+ $Y2=1.655
cc_543 N_A_73_367#_c_741_n N_VPWR_M1014_s 0.00356267f $X=2.115 $Y=2.1 $X2=0
+ $Y2=0
cc_544 N_A_73_367#_c_744_n N_VPWR_M1012_s 0.00343737f $X=2.975 $Y=2.1 $X2=0
+ $Y2=0
cc_545 N_A_73_367#_c_745_n N_VPWR_M1034_s 0.00214538f $X=3.515 $Y=2.215 $X2=0
+ $Y2=0
cc_546 N_A_73_367#_c_747_n N_VPWR_M1034_s 0.0100957f $X=4.05 $Y=2.425 $X2=0
+ $Y2=0
cc_547 N_A_73_367#_c_729_n N_VPWR_c_819_n 0.0170777f $X=1.255 $Y=1.81 $X2=0
+ $Y2=0
cc_548 N_A_73_367#_c_776_p N_VPWR_c_820_n 0.0124525f $X=1.35 $Y=2.44 $X2=0 $Y2=0
cc_549 N_A_73_367#_c_741_n N_VPWR_c_821_n 0.0170777f $X=2.115 $Y=2.1 $X2=0 $Y2=0
cc_550 N_A_73_367#_c_744_n N_VPWR_c_822_n 0.0170777f $X=2.975 $Y=2.1 $X2=0 $Y2=0
cc_551 N_A_73_367#_c_745_n N_VPWR_c_823_n 0.0084195f $X=3.515 $Y=2.215 $X2=0
+ $Y2=0
cc_552 N_A_73_367#_c_747_n N_VPWR_c_823_n 0.0196399f $X=4.05 $Y=2.425 $X2=0
+ $Y2=0
cc_553 N_A_73_367#_c_728_n N_VPWR_c_826_n 0.0178111f $X=0.49 $Y=1.98 $X2=0 $Y2=0
cc_554 N_A_73_367#_c_763_n N_VPWR_c_828_n 0.0361172f $X=4.855 $Y=2.99 $X2=0
+ $Y2=0
cc_555 N_A_73_367#_c_751_n N_VPWR_c_828_n 0.0164734f $X=4.185 $Y=2.99 $X2=0
+ $Y2=0
cc_556 N_A_73_367#_c_765_n N_VPWR_c_828_n 0.0361172f $X=5.715 $Y=2.99 $X2=0
+ $Y2=0
cc_557 N_A_73_367#_c_731_n N_VPWR_c_828_n 0.0179183f $X=5.845 $Y=2.905 $X2=0
+ $Y2=0
cc_558 N_A_73_367#_c_786_p N_VPWR_c_828_n 0.0125234f $X=4.95 $Y=2.99 $X2=0 $Y2=0
cc_559 N_A_73_367#_c_787_p N_VPWR_c_832_n 0.0124525f $X=2.21 $Y=2.91 $X2=0 $Y2=0
cc_560 N_A_73_367#_c_788_p N_VPWR_c_833_n 0.0128073f $X=3.07 $Y=2.545 $X2=0
+ $Y2=0
cc_561 N_A_73_367#_M1002_d N_VPWR_c_818_n 0.00371702f $X=0.365 $Y=1.835 $X2=0
+ $Y2=0
cc_562 N_A_73_367#_M1005_d N_VPWR_c_818_n 0.00536646f $X=1.21 $Y=1.835 $X2=0
+ $Y2=0
cc_563 N_A_73_367#_M1000_d N_VPWR_c_818_n 0.00536646f $X=2.07 $Y=1.835 $X2=0
+ $Y2=0
cc_564 N_A_73_367#_M1021_d N_VPWR_c_818_n 0.00501859f $X=2.93 $Y=1.835 $X2=0
+ $Y2=0
cc_565 N_A_73_367#_M1018_d N_VPWR_c_818_n 0.00223562f $X=3.95 $Y=1.835 $X2=0
+ $Y2=0
cc_566 N_A_73_367#_M1016_s N_VPWR_c_818_n 0.00223565f $X=4.81 $Y=1.835 $X2=0
+ $Y2=0
cc_567 N_A_73_367#_M1036_s N_VPWR_c_818_n 0.00215161f $X=5.67 $Y=1.835 $X2=0
+ $Y2=0
cc_568 N_A_73_367#_c_728_n N_VPWR_c_818_n 0.0100304f $X=0.49 $Y=1.98 $X2=0 $Y2=0
cc_569 N_A_73_367#_c_776_p N_VPWR_c_818_n 0.00730901f $X=1.35 $Y=2.44 $X2=0
+ $Y2=0
cc_570 N_A_73_367#_c_787_p N_VPWR_c_818_n 0.00730901f $X=2.21 $Y=2.91 $X2=0
+ $Y2=0
cc_571 N_A_73_367#_c_788_p N_VPWR_c_818_n 0.00769778f $X=3.07 $Y=2.545 $X2=0
+ $Y2=0
cc_572 N_A_73_367#_c_763_n N_VPWR_c_818_n 0.023676f $X=4.855 $Y=2.99 $X2=0 $Y2=0
cc_573 N_A_73_367#_c_751_n N_VPWR_c_818_n 0.0102636f $X=4.185 $Y=2.99 $X2=0
+ $Y2=0
cc_574 N_A_73_367#_c_765_n N_VPWR_c_818_n 0.023676f $X=5.715 $Y=2.99 $X2=0 $Y2=0
cc_575 N_A_73_367#_c_731_n N_VPWR_c_818_n 0.0101082f $X=5.845 $Y=2.905 $X2=0
+ $Y2=0
cc_576 N_A_73_367#_c_786_p N_VPWR_c_818_n 0.00738676f $X=4.95 $Y=2.99 $X2=0
+ $Y2=0
cc_577 N_A_73_367#_c_763_n N_Y_M1001_d 0.00332344f $X=4.855 $Y=2.99 $X2=0 $Y2=0
cc_578 N_A_73_367#_c_765_n N_Y_M1028_d 0.00332344f $X=5.715 $Y=2.99 $X2=0 $Y2=0
cc_579 N_A_73_367#_M1018_d N_Y_c_963_n 0.00113401f $X=3.95 $Y=1.835 $X2=0 $Y2=0
cc_580 N_A_73_367#_c_747_n N_Y_c_976_n 0.00497351f $X=4.05 $Y=2.425 $X2=0 $Y2=0
cc_581 N_A_73_367#_c_763_n N_Y_c_976_n 0.0159249f $X=4.855 $Y=2.99 $X2=0 $Y2=0
cc_582 N_A_73_367#_M1016_s N_Y_c_1000_n 0.00334718f $X=4.81 $Y=1.835 $X2=0 $Y2=0
cc_583 N_A_73_367#_c_811_p N_Y_c_1000_n 0.0136314f $X=4.95 $Y=2.42 $X2=0 $Y2=0
cc_584 N_A_73_367#_M1018_d N_Y_c_1005_n 0.002775f $X=3.95 $Y=1.835 $X2=0 $Y2=0
cc_585 N_A_73_367#_c_747_n N_Y_c_1005_n 0.0136549f $X=4.05 $Y=2.425 $X2=0 $Y2=0
cc_586 N_A_73_367#_c_765_n N_Y_c_1009_n 0.0159805f $X=5.715 $Y=2.99 $X2=0 $Y2=0
cc_587 N_A_73_367#_c_732_n N_A_1241_367#_c_1059_n 0.0136671f $X=5.81 $Y=2.055
+ $X2=0 $Y2=0
cc_588 N_A_73_367#_c_731_n N_A_1241_367#_c_1060_n 0.0136671f $X=5.845 $Y=2.905
+ $X2=0 $Y2=0
cc_589 N_A_73_367#_c_732_n N_A_1241_367#_c_1060_n 0.0597152f $X=5.81 $Y=2.055
+ $X2=0 $Y2=0
cc_590 N_VPWR_c_818_n N_Y_M1001_d 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_591 N_VPWR_c_818_n N_Y_M1028_d 0.00225186f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_592 N_VPWR_c_818_n N_A_1241_367#_M1008_d 0.00371702f $X=9.84 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_593 N_VPWR_c_818_n N_A_1241_367#_M1019_d 0.00536646f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_818_n N_A_1241_367#_M1038_d 0.00376625f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_818_n N_A_1241_367#_M1015_s 0.00220343f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_818_n N_A_1241_367#_M1033_s 0.00215159f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_828_n N_A_1241_367#_c_1060_n 0.0178111f $X=6.595 $Y=3.33 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_818_n N_A_1241_367#_c_1060_n 0.0100304f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_599 N_VPWR_M1008_s N_A_1241_367#_c_1073_n 0.00334983f $X=6.62 $Y=1.835 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_824_n N_A_1241_367#_c_1073_n 0.0170777f $X=6.76 $Y=2.375 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_830_n N_A_1241_367#_c_1101_n 0.0124525f $X=7.455 $Y=3.33 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_818_n N_A_1241_367#_c_1101_n 0.00730901f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_603 N_VPWR_M1029_s N_A_1241_367#_c_1077_n 0.00334983f $X=7.48 $Y=1.835 $X2=0
+ $Y2=0
cc_604 N_VPWR_c_825_n N_A_1241_367#_c_1077_n 0.0170777f $X=7.62 $Y=2.375 $X2=0
+ $Y2=0
cc_605 N_VPWR_c_834_n N_A_1241_367#_c_1105_n 0.0134105f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_606 N_VPWR_c_818_n N_A_1241_367#_c_1105_n 0.0083587f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_607 N_VPWR_c_834_n N_A_1241_367#_c_1065_n 0.0341772f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_608 N_VPWR_c_818_n N_A_1241_367#_c_1065_n 0.0216081f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_609 N_VPWR_c_834_n N_A_1241_367#_c_1068_n 0.0336481f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_610 N_VPWR_c_818_n N_A_1241_367#_c_1068_n 0.0210442f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_611 N_VPWR_c_834_n N_A_1241_367#_c_1061_n 0.0189465f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_612 N_VPWR_c_818_n N_A_1241_367#_c_1061_n 0.0112692f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_613 N_VPWR_c_834_n N_A_1241_367#_c_1113_n 0.0150071f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_614 N_VPWR_c_818_n N_A_1241_367#_c_1113_n 0.0101082f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_615 N_Y_c_968_n N_VGND_M1035_d 0.00465758f $X=3.995 $Y=0.892 $X2=0 $Y2=0
cc_616 N_Y_c_963_n N_VGND_M1035_d 5.21174e-19 $X=4.08 $Y=1.885 $X2=0 $Y2=0
cc_617 N_Y_c_965_n N_VGND_M1035_d 0.0011696f $X=4.545 $Y=1.13 $X2=0 $Y2=0
cc_618 N_Y_c_964_n N_VGND_M1030_d 0.00180746f $X=5.215 $Y=1.13 $X2=0 $Y2=0
cc_619 Y N_VGND_M1037_d 7.8956e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_620 N_Y_c_968_n N_VGND_c_1118_n 0.0115964f $X=3.995 $Y=0.892 $X2=0 $Y2=0
cc_621 N_Y_c_965_n N_VGND_c_1118_n 0.0094036f $X=4.545 $Y=1.13 $X2=0 $Y2=0
cc_622 N_Y_c_964_n N_VGND_c_1119_n 0.0163515f $X=5.215 $Y=1.13 $X2=0 $Y2=0
cc_623 Y N_VGND_c_1120_n 0.00556928f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_624 N_Y_c_968_n N_VGND_c_1128_n 0.00207897f $X=3.995 $Y=0.892 $X2=0 $Y2=0
cc_625 N_Y_c_1043_p N_VGND_c_1130_n 0.0140491f $X=4.45 $Y=0.42 $X2=0 $Y2=0
cc_626 N_Y_c_965_n N_VGND_c_1130_n 0.00213656f $X=4.545 $Y=1.13 $X2=0 $Y2=0
cc_627 N_Y_c_1045_p N_VGND_c_1132_n 0.0124525f $X=5.31 $Y=0.42 $X2=0 $Y2=0
cc_628 N_Y_M1004_d N_VGND_c_1141_n 0.00225186f $X=2.075 $Y=0.235 $X2=0 $Y2=0
cc_629 N_Y_M1020_d N_VGND_c_1141_n 0.00225186f $X=2.935 $Y=0.235 $X2=0 $Y2=0
cc_630 N_Y_M1017_s N_VGND_c_1141_n 0.00380103f $X=4.31 $Y=0.235 $X2=0 $Y2=0
cc_631 N_Y_M1031_s N_VGND_c_1141_n 0.00536646f $X=5.17 $Y=0.235 $X2=0 $Y2=0
cc_632 N_Y_c_968_n N_VGND_c_1141_n 0.00705887f $X=3.995 $Y=0.892 $X2=0 $Y2=0
cc_633 N_Y_c_1043_p N_VGND_c_1141_n 0.0090585f $X=4.45 $Y=0.42 $X2=0 $Y2=0
cc_634 N_Y_c_965_n N_VGND_c_1141_n 0.00443737f $X=4.545 $Y=1.13 $X2=0 $Y2=0
cc_635 N_Y_c_1045_p N_VGND_c_1141_n 0.00730901f $X=5.31 $Y=0.42 $X2=0 $Y2=0
cc_636 N_Y_c_968_n N_A_157_47#_M1010_s 0.0033307f $X=3.995 $Y=0.892 $X2=0 $Y2=0
cc_637 N_Y_c_968_n N_A_157_47#_M1023_s 0.00434417f $X=3.995 $Y=0.892 $X2=0 $Y2=0
cc_638 N_Y_M1004_d N_A_157_47#_c_1285_n 0.0033152f $X=2.075 $Y=0.235 $X2=0 $Y2=0
cc_639 N_Y_M1020_d N_A_157_47#_c_1285_n 0.0033152f $X=2.935 $Y=0.235 $X2=0 $Y2=0
cc_640 N_Y_c_968_n N_A_157_47#_c_1285_n 0.0844995f $X=3.995 $Y=0.892 $X2=0 $Y2=0
cc_641 N_VGND_c_1141_n N_A_157_47#_M1003_s 0.00397496f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_642 N_VGND_c_1141_n N_A_157_47#_M1025_s 0.00376627f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_643 N_VGND_c_1141_n N_A_157_47#_M1010_s 0.00223577f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_644 N_VGND_c_1141_n N_A_157_47#_M1023_s 0.0022036f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_645 N_VGND_c_1116_n N_A_157_47#_c_1299_n 0.0138717f $X=1.19 $Y=0 $X2=0 $Y2=0
cc_646 N_VGND_c_1141_n N_A_157_47#_c_1299_n 0.00886411f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_647 N_VGND_M1013_d N_A_157_47#_c_1274_n 0.00176461f $X=1.215 $Y=0.235 $X2=0
+ $Y2=0
cc_648 N_VGND_c_1117_n N_A_157_47#_c_1274_n 0.0170777f $X=1.355 $Y=0.36 $X2=0
+ $Y2=0
cc_649 N_VGND_c_1115_n N_A_157_47#_c_1275_n 0.00166417f $X=0.495 $Y=0.38 $X2=0
+ $Y2=0
cc_650 N_VGND_c_1128_n N_A_157_47#_c_1304_n 0.0121686f $X=3.81 $Y=0 $X2=0 $Y2=0
cc_651 N_VGND_c_1141_n N_A_157_47#_c_1304_n 0.00698742f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_652 N_VGND_c_1128_n N_A_157_47#_c_1285_n 0.100358f $X=3.81 $Y=0 $X2=0 $Y2=0
cc_653 N_VGND_c_1141_n N_A_157_47#_c_1285_n 0.0645089f $X=9.84 $Y=0 $X2=0 $Y2=0
