* File: sky130_fd_sc_lp__a221o_4.pxi.spice
* Created: Fri Aug 28 09:52:41 2020
* 
x_PM_SKY130_FD_SC_LP__A221O_4%A_83_21# N_A_83_21#_M1013_s N_A_83_21#_M1020_s
+ N_A_83_21#_M1011_s N_A_83_21#_M1024_d N_A_83_21#_M1016_s N_A_83_21#_M1003_g
+ N_A_83_21#_M1007_g N_A_83_21#_M1012_g N_A_83_21#_M1008_g N_A_83_21#_M1014_g
+ N_A_83_21#_M1018_g N_A_83_21#_M1021_g N_A_83_21#_M1023_g N_A_83_21#_c_191_p
+ N_A_83_21#_c_133_n N_A_83_21#_c_154_p N_A_83_21#_c_261_p N_A_83_21#_c_124_n
+ N_A_83_21#_c_135_n N_A_83_21#_c_163_p N_A_83_21#_c_165_p N_A_83_21#_c_263_p
+ N_A_83_21#_c_125_n N_A_83_21#_c_126_n N_A_83_21#_c_127_n N_A_83_21#_c_137_n
+ N_A_83_21#_c_128_n PM_SKY130_FD_SC_LP__A221O_4%A_83_21#
x_PM_SKY130_FD_SC_LP__A221O_4%A2 N_A2_c_289_n N_A2_M1000_g N_A2_M1002_g
+ N_A2_c_291_n N_A2_M1009_g N_A2_M1017_g A2 A2 N_A2_c_294_n
+ PM_SKY130_FD_SC_LP__A221O_4%A2
x_PM_SKY130_FD_SC_LP__A221O_4%A1 N_A1_M1015_g N_A1_M1025_g N_A1_c_338_n
+ N_A1_M1013_g N_A1_c_339_n N_A1_M1020_g A1 N_A1_c_351_n N_A1_c_340_n
+ PM_SKY130_FD_SC_LP__A221O_4%A1
x_PM_SKY130_FD_SC_LP__A221O_4%C1 N_C1_c_382_n N_C1_M1001_g N_C1_M1016_g
+ N_C1_c_384_n N_C1_M1011_g N_C1_M1026_g C1 C1 N_C1_c_387_n
+ PM_SKY130_FD_SC_LP__A221O_4%C1
x_PM_SKY130_FD_SC_LP__A221O_4%B1 N_B1_c_430_n N_B1_M1005_g N_B1_M1004_g
+ N_B1_c_432_n N_B1_M1024_g N_B1_M1019_g B1 B1 N_B1_c_435_n
+ PM_SKY130_FD_SC_LP__A221O_4%B1
x_PM_SKY130_FD_SC_LP__A221O_4%B2 N_B2_M1010_g N_B2_M1027_g N_B2_M1006_g
+ N_B2_M1022_g B2 B2 N_B2_c_483_n N_B2_c_488_n B2 PM_SKY130_FD_SC_LP__A221O_4%B2
x_PM_SKY130_FD_SC_LP__A221O_4%VPWR N_VPWR_M1007_d N_VPWR_M1008_d N_VPWR_M1023_d
+ N_VPWR_M1017_s N_VPWR_M1025_d N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n
+ N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n
+ N_VPWR_c_535_n N_VPWR_c_536_n N_VPWR_c_537_n VPWR N_VPWR_c_538_n
+ N_VPWR_c_539_n N_VPWR_c_526_n N_VPWR_c_541_n N_VPWR_c_542_n
+ PM_SKY130_FD_SC_LP__A221O_4%VPWR
x_PM_SKY130_FD_SC_LP__A221O_4%X N_X_M1003_d N_X_M1014_d N_X_M1007_s N_X_M1018_s
+ N_X_c_635_n N_X_c_640_n N_X_c_641_n N_X_c_686_p N_X_c_673_n N_X_c_642_n
+ N_X_c_636_n N_X_c_685_p N_X_c_677_n N_X_c_637_n N_X_c_643_n X X N_X_c_638_n X
+ PM_SKY130_FD_SC_LP__A221O_4%X
x_PM_SKY130_FD_SC_LP__A221O_4%A_457_367# N_A_457_367#_M1002_d
+ N_A_457_367#_M1015_s N_A_457_367#_M1004_d N_A_457_367#_M1010_d
+ N_A_457_367#_c_698_n N_A_457_367#_c_737_n N_A_457_367#_c_699_n
+ N_A_457_367#_c_741_n N_A_457_367#_c_691_n N_A_457_367#_c_692_n
+ N_A_457_367#_c_705_n N_A_457_367#_c_693_n N_A_457_367#_c_708_n
+ N_A_457_367#_c_694_n N_A_457_367#_c_695_n N_A_457_367#_c_757_p
+ N_A_457_367#_c_710_n PM_SKY130_FD_SC_LP__A221O_4%A_457_367#
x_PM_SKY130_FD_SC_LP__A221O_4%A_822_367# N_A_822_367#_M1016_d
+ N_A_822_367#_M1026_d N_A_822_367#_M1019_s N_A_822_367#_M1027_s
+ N_A_822_367#_c_759_n N_A_822_367#_c_769_n N_A_822_367#_c_774_n
+ N_A_822_367#_c_760_n N_A_822_367#_c_761_n N_A_822_367#_c_771_n
+ PM_SKY130_FD_SC_LP__A221O_4%A_822_367#
x_PM_SKY130_FD_SC_LP__A221O_4%VGND N_VGND_M1003_s N_VGND_M1012_s N_VGND_M1021_s
+ N_VGND_M1009_s N_VGND_M1001_d N_VGND_M1006_d N_VGND_c_807_n N_VGND_c_808_n
+ N_VGND_c_809_n N_VGND_c_810_n N_VGND_c_811_n N_VGND_c_812_n N_VGND_c_813_n
+ N_VGND_c_814_n N_VGND_c_815_n N_VGND_c_816_n N_VGND_c_817_n VGND
+ N_VGND_c_818_n N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n
+ N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n PM_SKY130_FD_SC_LP__A221O_4%VGND
x_PM_SKY130_FD_SC_LP__A221O_4%A_457_47# N_A_457_47#_M1000_d N_A_457_47#_M1013_d
+ N_A_457_47#_c_942_n N_A_457_47#_c_922_n N_A_457_47#_c_932_n
+ N_A_457_47#_c_928_n PM_SKY130_FD_SC_LP__A221O_4%A_457_47#
x_PM_SKY130_FD_SC_LP__A221O_4%A_1077_47# N_A_1077_47#_M1005_s
+ N_A_1077_47#_M1006_s N_A_1077_47#_M1022_s N_A_1077_47#_c_947_n
+ N_A_1077_47#_c_948_n N_A_1077_47#_c_949_n N_A_1077_47#_c_950_n
+ N_A_1077_47#_c_951_n PM_SKY130_FD_SC_LP__A221O_4%A_1077_47#
cc_1 VNB N_A_83_21#_M1003_g 0.0264787f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_2 VNB N_A_83_21#_M1012_g 0.0217751f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.655
cc_3 VNB N_A_83_21#_M1014_g 0.021796f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_4 VNB N_A_83_21#_M1021_g 0.0233423f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_5 VNB N_A_83_21#_c_124_n 0.0113078f $X=-0.19 $Y=-0.245 $X2=4.21 $Y2=1.69
cc_6 VNB N_A_83_21#_c_125_n 0.00299093f $X=-0.19 $Y=-0.245 $X2=5.955 $Y2=0.4
cc_7 VNB N_A_83_21#_c_126_n 0.00409881f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.492
cc_8 VNB N_A_83_21#_c_127_n 0.0043152f $X=-0.19 $Y=-0.245 $X2=3.37 $Y2=0.34
cc_9 VNB N_A_83_21#_c_128_n 0.0704017f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.49
cc_10 VNB N_A2_c_289_n 0.0161955f $X=-0.19 $Y=-0.245 $X2=3.25 $Y2=0.235
cc_11 VNB N_A2_M1002_g 0.00718672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_291_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_M1017_g 0.00703883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A2 0.00392191f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.325
cc_15 VNB N_A2_c_294_n 0.0429085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_M1015_g 0.0072287f $X=-0.19 $Y=-0.245 $X2=4.955 $Y2=0.235
cc_17 VNB N_A1_M1025_g 0.00863263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_338_n 0.0220758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_339_n 0.0164051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_340_n 0.0800248f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.325
cc_21 VNB N_C1_c_382_n 0.0169108f $X=-0.19 $Y=-0.245 $X2=3.25 $Y2=0.235
cc_22 VNB N_C1_M1016_g 0.00706954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C1_c_384_n 0.0169651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C1_M1026_g 0.00677515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB C1 0.00986389f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.325
cc_26 VNB N_C1_c_387_n 0.0357404f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.325
cc_27 VNB N_B1_c_430_n 0.0169694f $X=-0.19 $Y=-0.245 $X2=3.25 $Y2=0.235
cc_28 VNB N_B1_M1004_g 0.00677981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B1_c_432_n 0.0207694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B1_M1019_g 0.00677981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB B1 0.00630591f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.325
cc_32 VNB N_B1_c_435_n 0.0455013f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.325
cc_33 VNB N_B2_M1006_g 0.0271803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B2_M1022_g 0.0289145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB B2 0.0133486f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_36 VNB N_B2_c_483_n 0.076578f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.655
cc_37 VNB N_VPWR_c_526_n 0.322901f $X=-0.19 $Y=-0.245 $X2=4.665 $Y2=2.14
cc_38 VNB N_X_c_635_n 0.00143138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_636_n 0.00631347f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_40 VNB N_X_c_637_n 0.00144228f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_41 VNB N_X_c_638_n 0.00802798f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.492
cc_42 VNB X 0.0209285f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.49
cc_43 VNB N_VGND_c_807_n 0.0108441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_808_n 0.0282332f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_45 VNB N_VGND_c_809_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.655
cc_46 VNB N_VGND_c_810_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.465
cc_47 VNB N_VGND_c_811_n 0.00711269f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.655
cc_48 VNB N_VGND_c_812_n 0.00522139f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.465
cc_49 VNB N_VGND_c_813_n 7.46595e-19 $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=0.655
cc_50 VNB N_VGND_c_814_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.655
cc_51 VNB N_VGND_c_815_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.465
cc_52 VNB N_VGND_c_816_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_817_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.492
cc_54 VNB N_VGND_c_818_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.49
cc_55 VNB N_VGND_c_819_n 0.0370061f $X=-0.19 $Y=-0.245 $X2=4.21 $Y2=1.69
cc_56 VNB N_VGND_c_820_n 0.0465179f $X=-0.19 $Y=-0.245 $X2=4.365 $Y2=0.94
cc_57 VNB N_VGND_c_821_n 0.0181466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_822_n 0.378113f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.492
cc_59 VNB N_VGND_c_823_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.37 $Y2=0.51
cc_60 VNB N_VGND_c_824_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.245 $Y2=0.34
cc_61 VNB N_VGND_c_825_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=4.21 $Y2=1.782
cc_62 VNB N_A_457_47#_c_922_n 0.00744826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1077_47#_c_947_n 0.00821659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1077_47#_c_948_n 0.00511077f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.325
cc_65 VNB N_A_1077_47#_c_949_n 0.012746f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_66 VNB N_A_1077_47#_c_950_n 0.0307328f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_67 VNB N_A_1077_47#_c_951_n 0.00540181f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.325
cc_68 VPB N_A_83_21#_M1007_g 0.0224142f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_69 VPB N_A_83_21#_M1008_g 0.0188421f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_70 VPB N_A_83_21#_M1018_g 0.0188567f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_71 VPB N_A_83_21#_M1023_g 0.0188007f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_72 VPB N_A_83_21#_c_133_n 0.0193682f $X=-0.19 $Y=1.655 $X2=4.125 $Y2=1.782
cc_73 VPB N_A_83_21#_c_124_n 8.42598e-19 $X=-0.19 $Y=1.655 $X2=4.21 $Y2=1.69
cc_74 VPB N_A_83_21#_c_135_n 0.00505798f $X=-0.19 $Y=1.655 $X2=4.5 $Y2=1.79
cc_75 VPB N_A_83_21#_c_126_n 6.07831e-19 $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.492
cc_76 VPB N_A_83_21#_c_137_n 5.36628e-19 $X=-0.19 $Y=1.655 $X2=4.21 $Y2=1.782
cc_77 VPB N_A_83_21#_c_128_n 0.00700947f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=1.49
cc_78 VPB N_A2_M1002_g 0.0184403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A2_M1017_g 0.0184505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A1_M1015_g 0.0184515f $X=-0.19 $Y=1.655 $X2=4.955 $Y2=0.235
cc_81 VPB N_A1_M1025_g 0.02294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_C1_M1016_g 0.0234833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_C1_M1026_g 0.0196034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_B1_M1004_g 0.0196052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_B1_M1019_g 0.0188441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_B2_M1010_g 0.017738f $X=-0.19 $Y=1.655 $X2=4.955 $Y2=0.235
cc_87 VPB N_B2_M1027_g 0.0246989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB B2 0.0241822f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.655
cc_89 VPB N_B2_c_483_n 0.0236431f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.655
cc_90 VPB N_B2_c_488_n 0.00304121f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_91 VPB N_VPWR_c_527_n 0.0108182f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.325
cc_92 VPB N_VPWR_c_528_n 0.0415885f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.655
cc_93 VPB N_VPWR_c_529_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.325
cc_94 VPB N_VPWR_c_530_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.465
cc_95 VPB N_VPWR_c_531_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.655
cc_96 VPB N_VPWR_c_532_n 0.012974f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.465
cc_97 VPB N_VPWR_c_533_n 0.0107183f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=0.655
cc_98 VPB N_VPWR_c_534_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_99 VPB N_VPWR_c_535_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.78 $Y2=2.465
cc_100 VPB N_VPWR_c_536_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_537_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.85 $Y2=1.492
cc_102 VPB N_VPWR_c_538_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.49
cc_103 VPB N_VPWR_c_539_n 0.0962607f $X=-0.19 $Y=1.655 $X2=4.665 $Y2=1.875
cc_104 VPB N_VPWR_c_526_n 0.0787088f $X=-0.19 $Y=1.655 $X2=4.665 $Y2=2.14
cc_105 VPB N_VPWR_c_541_n 0.00436868f $X=-0.19 $Y=1.655 $X2=5.955 $Y2=0.385
cc_106 VPB N_VPWR_c_542_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.492
cc_107 VPB N_X_c_640_n 0.00143138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_X_c_641_n 0.00779219f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.325
cc_109 VPB N_X_c_642_n 0.00520893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_X_c_643_n 0.00134924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB X 0.00491218f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.49
cc_112 VPB N_A_457_367#_c_691_n 0.0105496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_457_367#_c_692_n 0.0030259f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.655
cc_114 VPB N_A_457_367#_c_693_n 0.00188293f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.655
cc_115 VPB N_A_457_367#_c_694_n 0.00888893f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=0.655
cc_116 VPB N_A_457_367#_c_695_n 0.00192029f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=0.655
cc_117 VPB N_A_822_367#_c_759_n 0.00317703f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_822_367#_c_760_n 0.00747154f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.655
cc_119 VPB N_A_822_367#_c_761_n 0.0379527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 N_A_83_21#_M1021_g N_A2_c_289_n 0.0172225f $X=1.78 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_83_21#_c_133_n N_A2_M1002_g 0.0153271f $X=4.125 $Y=1.782 $X2=0 $Y2=0
cc_122 N_A_83_21#_c_126_n N_A2_M1002_g 0.00412851f $X=1.935 $Y=1.492 $X2=0 $Y2=0
cc_123 N_A_83_21#_c_128_n N_A2_M1002_g 0.025802f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_124 N_A_83_21#_c_127_n N_A2_c_291_n 7.89306e-19 $X=3.37 $Y=0.34 $X2=0 $Y2=0
cc_125 N_A_83_21#_c_133_n N_A2_M1017_g 0.0110074f $X=4.125 $Y=1.782 $X2=0 $Y2=0
cc_126 N_A_83_21#_M1021_g A2 0.00111729f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_127 N_A_83_21#_c_133_n A2 0.0744914f $X=4.125 $Y=1.782 $X2=0 $Y2=0
cc_128 N_A_83_21#_c_126_n A2 0.00910954f $X=1.935 $Y=1.492 $X2=0 $Y2=0
cc_129 N_A_83_21#_M1021_g N_A2_c_294_n 0.0182491f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_130 N_A_83_21#_c_133_n N_A2_c_294_n 0.00450442f $X=4.125 $Y=1.782 $X2=0 $Y2=0
cc_131 N_A_83_21#_c_126_n N_A2_c_294_n 8.95767e-19 $X=1.935 $Y=1.492 $X2=0 $Y2=0
cc_132 N_A_83_21#_c_133_n N_A1_M1015_g 0.0110581f $X=4.125 $Y=1.782 $X2=0 $Y2=0
cc_133 N_A_83_21#_c_133_n N_A1_M1025_g 0.0133316f $X=4.125 $Y=1.782 $X2=0 $Y2=0
cc_134 N_A_83_21#_c_124_n N_A1_M1025_g 0.00400735f $X=4.21 $Y=1.69 $X2=0 $Y2=0
cc_135 N_A_83_21#_c_154_p N_A1_c_338_n 0.00882437f $X=4.125 $Y=0.34 $X2=0 $Y2=0
cc_136 N_A_83_21#_c_127_n N_A1_c_338_n 0.00601598f $X=3.37 $Y=0.34 $X2=0 $Y2=0
cc_137 N_A_83_21#_c_154_p N_A1_c_339_n 0.0119618f $X=4.125 $Y=0.34 $X2=0 $Y2=0
cc_138 N_A_83_21#_c_124_n N_A1_c_339_n 0.00586364f $X=4.21 $Y=1.69 $X2=0 $Y2=0
cc_139 N_A_83_21#_c_127_n N_A1_c_339_n 5.19462e-19 $X=3.37 $Y=0.34 $X2=0 $Y2=0
cc_140 N_A_83_21#_c_133_n N_A1_c_351_n 0.0423552f $X=4.125 $Y=1.782 $X2=0 $Y2=0
cc_141 N_A_83_21#_c_124_n N_A1_c_351_n 0.0258783f $X=4.21 $Y=1.69 $X2=0 $Y2=0
cc_142 N_A_83_21#_c_133_n N_A1_c_340_n 0.0181687f $X=4.125 $Y=1.782 $X2=0 $Y2=0
cc_143 N_A_83_21#_c_124_n N_C1_c_382_n 0.0128739f $X=4.21 $Y=1.69 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A_83_21#_c_163_p N_C1_c_382_n 0.0127044f $X=4.965 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_83_21#_c_135_n N_C1_M1016_g 0.0165495f $X=4.5 $Y=1.79 $X2=0 $Y2=0
cc_146 N_A_83_21#_c_165_p N_C1_M1016_g 0.011021f $X=4.665 $Y=2.14 $X2=0 $Y2=0
cc_147 N_A_83_21#_c_137_n N_C1_M1016_g 6.80097e-19 $X=4.21 $Y=1.782 $X2=0 $Y2=0
cc_148 N_A_83_21#_c_163_p N_C1_c_384_n 0.00998618f $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_149 N_A_83_21#_c_135_n N_C1_M1026_g 0.00537419f $X=4.5 $Y=1.79 $X2=0 $Y2=0
cc_150 N_A_83_21#_c_165_p N_C1_M1026_g 0.00812327f $X=4.665 $Y=2.14 $X2=0 $Y2=0
cc_151 N_A_83_21#_c_124_n C1 0.026147f $X=4.21 $Y=1.69 $X2=0 $Y2=0
cc_152 N_A_83_21#_c_135_n C1 0.0284092f $X=4.5 $Y=1.79 $X2=0 $Y2=0
cc_153 N_A_83_21#_c_163_p C1 0.0436749f $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_154 N_A_83_21#_c_135_n N_C1_c_387_n 0.00230174f $X=4.5 $Y=1.79 $X2=0 $Y2=0
cc_155 N_A_83_21#_c_163_p N_C1_c_387_n 0.00224206f $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_156 N_A_83_21#_c_125_n N_B1_c_430_n 0.0149068f $X=5.955 $Y=0.4 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A_83_21#_c_135_n N_B1_M1004_g 4.98432e-19 $X=4.5 $Y=1.79 $X2=0 $Y2=0
cc_158 N_A_83_21#_c_165_p N_B1_M1004_g 0.00117675f $X=4.665 $Y=2.14 $X2=0 $Y2=0
cc_159 N_A_83_21#_c_125_n N_B1_c_432_n 0.0099907f $X=5.955 $Y=0.4 $X2=0 $Y2=0
cc_160 N_A_83_21#_c_133_n N_VPWR_M1023_d 7.12265e-19 $X=4.125 $Y=1.782 $X2=0
+ $Y2=0
cc_161 N_A_83_21#_c_126_n N_VPWR_M1023_d 0.00126408f $X=1.935 $Y=1.492 $X2=0
+ $Y2=0
cc_162 N_A_83_21#_c_133_n N_VPWR_M1017_s 0.00177354f $X=4.125 $Y=1.782 $X2=0
+ $Y2=0
cc_163 N_A_83_21#_c_133_n N_VPWR_M1025_d 0.00240575f $X=4.125 $Y=1.782 $X2=0
+ $Y2=0
cc_164 N_A_83_21#_M1007_g N_VPWR_c_528_n 0.0153838f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_83_21#_M1008_g N_VPWR_c_528_n 7.27171e-19 $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_83_21#_M1007_g N_VPWR_c_529_n 7.42371e-19 $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_83_21#_M1008_g N_VPWR_c_529_n 0.0144441f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A_83_21#_M1018_g N_VPWR_c_529_n 0.0142189f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_83_21#_M1023_g N_VPWR_c_529_n 7.27171e-19 $X=1.78 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_83_21#_M1018_g N_VPWR_c_530_n 7.41316e-19 $X=1.35 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_83_21#_M1023_g N_VPWR_c_530_n 0.0153036f $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A_83_21#_c_191_p N_VPWR_c_530_n 6.474e-19 $X=1.85 $Y=1.492 $X2=0 $Y2=0
cc_173 N_A_83_21#_c_133_n N_VPWR_c_530_n 0.00654259f $X=4.125 $Y=1.782 $X2=0
+ $Y2=0
cc_174 N_A_83_21#_c_126_n N_VPWR_c_530_n 0.00968462f $X=1.935 $Y=1.492 $X2=0
+ $Y2=0
cc_175 N_A_83_21#_M1018_g N_VPWR_c_534_n 0.00486043f $X=1.35 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_83_21#_M1023_g N_VPWR_c_534_n 0.00486043f $X=1.78 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_83_21#_M1007_g N_VPWR_c_538_n 0.00486043f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_83_21#_M1008_g N_VPWR_c_538_n 0.00486043f $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A_83_21#_M1016_s N_VPWR_c_526_n 0.00225465f $X=4.525 $Y=1.835 $X2=0
+ $Y2=0
cc_180 N_A_83_21#_M1007_g N_VPWR_c_526_n 0.00824727f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_83_21#_M1008_g N_VPWR_c_526_n 0.00824727f $X=0.92 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_83_21#_M1018_g N_VPWR_c_526_n 0.00824727f $X=1.35 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_83_21#_M1023_g N_VPWR_c_526_n 0.00824727f $X=1.78 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_83_21#_M1003_g N_X_c_635_n 0.0164915f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_185 N_A_83_21#_c_191_p N_X_c_635_n 0.00729511f $X=1.85 $Y=1.492 $X2=0 $Y2=0
cc_186 N_A_83_21#_M1007_g N_X_c_640_n 0.0155886f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A_83_21#_c_191_p N_X_c_640_n 0.00729511f $X=1.85 $Y=1.492 $X2=0 $Y2=0
cc_188 N_A_83_21#_M1008_g N_X_c_642_n 0.0131657f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_83_21#_M1018_g N_X_c_642_n 0.0130035f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A_83_21#_M1023_g N_X_c_642_n 6.8937e-19 $X=1.78 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_83_21#_c_191_p N_X_c_642_n 0.0631595f $X=1.85 $Y=1.492 $X2=0 $Y2=0
cc_192 N_A_83_21#_c_126_n N_X_c_642_n 0.0071394f $X=1.935 $Y=1.492 $X2=0 $Y2=0
cc_193 N_A_83_21#_c_128_n N_X_c_642_n 0.00497162f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_194 N_A_83_21#_M1012_g N_X_c_636_n 0.0145172f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A_83_21#_M1014_g N_X_c_636_n 0.0141546f $X=1.35 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A_83_21#_M1021_g N_X_c_636_n 0.00417933f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_197 N_A_83_21#_c_191_p N_X_c_636_n 0.062752f $X=1.85 $Y=1.492 $X2=0 $Y2=0
cc_198 N_A_83_21#_c_128_n N_X_c_636_n 0.00500688f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_199 N_A_83_21#_c_191_p N_X_c_637_n 0.0154156f $X=1.85 $Y=1.492 $X2=0 $Y2=0
cc_200 N_A_83_21#_c_128_n N_X_c_637_n 0.00255183f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_201 N_A_83_21#_c_191_p N_X_c_643_n 0.0146041f $X=1.85 $Y=1.492 $X2=0 $Y2=0
cc_202 N_A_83_21#_c_128_n N_X_c_643_n 0.00253619f $X=1.78 $Y=1.49 $X2=0 $Y2=0
cc_203 N_A_83_21#_M1003_g X 0.0198406f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_204 N_A_83_21#_c_191_p X 0.0149238f $X=1.85 $Y=1.492 $X2=0 $Y2=0
cc_205 N_A_83_21#_c_133_n N_A_457_367#_M1002_d 0.00176922f $X=4.125 $Y=1.782
+ $X2=-0.19 $Y2=-0.245
cc_206 N_A_83_21#_c_133_n N_A_457_367#_M1015_s 0.00176922f $X=4.125 $Y=1.782
+ $X2=0 $Y2=0
cc_207 N_A_83_21#_c_133_n N_A_457_367#_c_698_n 0.0135828f $X=4.125 $Y=1.782
+ $X2=0 $Y2=0
cc_208 N_A_83_21#_c_133_n N_A_457_367#_c_699_n 0.0326748f $X=4.125 $Y=1.782
+ $X2=0 $Y2=0
cc_209 N_A_83_21#_c_133_n N_A_457_367#_c_691_n 0.0473196f $X=4.125 $Y=1.782
+ $X2=0 $Y2=0
cc_210 N_A_83_21#_c_135_n N_A_457_367#_c_691_n 0.00156751f $X=4.5 $Y=1.79 $X2=0
+ $Y2=0
cc_211 N_A_83_21#_c_165_p N_A_457_367#_c_691_n 0.0131487f $X=4.665 $Y=2.14 $X2=0
+ $Y2=0
cc_212 N_A_83_21#_c_137_n N_A_457_367#_c_691_n 0.0151295f $X=4.21 $Y=1.782 $X2=0
+ $Y2=0
cc_213 N_A_83_21#_c_165_p N_A_457_367#_c_692_n 0.00422906f $X=4.665 $Y=2.14
+ $X2=0 $Y2=0
cc_214 N_A_83_21#_M1016_s N_A_457_367#_c_705_n 0.00348701f $X=4.525 $Y=1.835
+ $X2=0 $Y2=0
cc_215 N_A_83_21#_c_135_n N_A_457_367#_c_705_n 0.00316052f $X=4.5 $Y=1.79 $X2=0
+ $Y2=0
cc_216 N_A_83_21#_c_165_p N_A_457_367#_c_705_n 0.0168339f $X=4.665 $Y=2.14 $X2=0
+ $Y2=0
cc_217 N_A_83_21#_c_165_p N_A_457_367#_c_708_n 0.0115866f $X=4.665 $Y=2.14 $X2=0
+ $Y2=0
cc_218 N_A_83_21#_c_135_n N_A_457_367#_c_695_n 0.00563554f $X=4.5 $Y=1.79 $X2=0
+ $Y2=0
cc_219 N_A_83_21#_c_133_n N_A_457_367#_c_710_n 0.0135828f $X=4.125 $Y=1.782
+ $X2=0 $Y2=0
cc_220 N_A_83_21#_c_135_n N_A_822_367#_M1016_d 2.01974e-19 $X=4.5 $Y=1.79
+ $X2=-0.19 $Y2=-0.245
cc_221 N_A_83_21#_c_137_n N_A_822_367#_M1016_d 0.00203624f $X=4.21 $Y=1.782
+ $X2=-0.19 $Y2=-0.245
cc_222 N_A_83_21#_M1016_s N_A_822_367#_c_759_n 0.00341454f $X=4.525 $Y=1.835
+ $X2=0 $Y2=0
cc_223 N_A_83_21#_c_163_p N_VGND_M1001_d 0.00328279f $X=4.965 $Y=0.94 $X2=0
+ $Y2=0
cc_224 N_A_83_21#_M1003_g N_VGND_c_808_n 0.0125061f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_225 N_A_83_21#_M1012_g N_VGND_c_808_n 6.29568e-19 $X=0.92 $Y=0.655 $X2=0
+ $Y2=0
cc_226 N_A_83_21#_M1003_g N_VGND_c_809_n 6.25324e-19 $X=0.49 $Y=0.655 $X2=0
+ $Y2=0
cc_227 N_A_83_21#_M1012_g N_VGND_c_809_n 0.0110627f $X=0.92 $Y=0.655 $X2=0 $Y2=0
cc_228 N_A_83_21#_M1014_g N_VGND_c_809_n 0.0110627f $X=1.35 $Y=0.655 $X2=0 $Y2=0
cc_229 N_A_83_21#_M1021_g N_VGND_c_809_n 6.25324e-19 $X=1.78 $Y=0.655 $X2=0
+ $Y2=0
cc_230 N_A_83_21#_M1014_g N_VGND_c_810_n 6.64931e-19 $X=1.35 $Y=0.655 $X2=0
+ $Y2=0
cc_231 N_A_83_21#_M1021_g N_VGND_c_810_n 0.0137058f $X=1.78 $Y=0.655 $X2=0 $Y2=0
cc_232 N_A_83_21#_c_191_p N_VGND_c_810_n 7.52263e-19 $X=1.85 $Y=1.492 $X2=0
+ $Y2=0
cc_233 N_A_83_21#_c_133_n N_VGND_c_810_n 0.00315204f $X=4.125 $Y=1.782 $X2=0
+ $Y2=0
cc_234 N_A_83_21#_c_126_n N_VGND_c_810_n 0.00689755f $X=1.935 $Y=1.492 $X2=0
+ $Y2=0
cc_235 N_A_83_21#_c_127_n N_VGND_c_811_n 0.0322659f $X=3.37 $Y=0.34 $X2=0 $Y2=0
cc_236 N_A_83_21#_c_163_p N_VGND_c_812_n 0.0132261f $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_237 N_A_83_21#_M1014_g N_VGND_c_814_n 0.00486043f $X=1.35 $Y=0.655 $X2=0
+ $Y2=0
cc_238 N_A_83_21#_M1021_g N_VGND_c_814_n 0.00486043f $X=1.78 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_A_83_21#_M1003_g N_VGND_c_818_n 0.00486043f $X=0.49 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_83_21#_M1012_g N_VGND_c_818_n 0.00486043f $X=0.92 $Y=0.655 $X2=0
+ $Y2=0
cc_241 N_A_83_21#_c_154_p N_VGND_c_819_n 0.0331045f $X=4.125 $Y=0.34 $X2=0 $Y2=0
cc_242 N_A_83_21#_c_261_p N_VGND_c_819_n 0.0142975f $X=4.245 $Y=0.425 $X2=0
+ $Y2=0
cc_243 N_A_83_21#_c_127_n N_VGND_c_819_n 0.0197669f $X=3.37 $Y=0.34 $X2=0 $Y2=0
cc_244 N_A_83_21#_c_263_p N_VGND_c_820_n 0.0153619f $X=5.1 $Y=0.515 $X2=0 $Y2=0
cc_245 N_A_83_21#_c_125_n N_VGND_c_820_n 0.05201f $X=5.955 $Y=0.4 $X2=0 $Y2=0
cc_246 N_A_83_21#_M1013_s N_VGND_c_822_n 0.00215962f $X=3.25 $Y=0.235 $X2=0
+ $Y2=0
cc_247 N_A_83_21#_M1020_s N_VGND_c_822_n 0.00229732f $X=4.095 $Y=0.235 $X2=0
+ $Y2=0
cc_248 N_A_83_21#_M1011_s N_VGND_c_822_n 0.0022973f $X=4.955 $Y=0.235 $X2=0
+ $Y2=0
cc_249 N_A_83_21#_M1024_d N_VGND_c_822_n 0.00215176f $X=5.815 $Y=0.235 $X2=0
+ $Y2=0
cc_250 N_A_83_21#_M1003_g N_VGND_c_822_n 0.00824727f $X=0.49 $Y=0.655 $X2=0
+ $Y2=0
cc_251 N_A_83_21#_M1012_g N_VGND_c_822_n 0.00824727f $X=0.92 $Y=0.655 $X2=0
+ $Y2=0
cc_252 N_A_83_21#_M1014_g N_VGND_c_822_n 0.00824727f $X=1.35 $Y=0.655 $X2=0
+ $Y2=0
cc_253 N_A_83_21#_M1021_g N_VGND_c_822_n 0.00824727f $X=1.78 $Y=0.655 $X2=0
+ $Y2=0
cc_254 N_A_83_21#_c_154_p N_VGND_c_822_n 0.0209991f $X=4.125 $Y=0.34 $X2=0 $Y2=0
cc_255 N_A_83_21#_c_261_p N_VGND_c_822_n 0.00933065f $X=4.245 $Y=0.425 $X2=0
+ $Y2=0
cc_256 N_A_83_21#_c_163_p N_VGND_c_822_n 0.0101042f $X=4.965 $Y=0.94 $X2=0 $Y2=0
cc_257 N_A_83_21#_c_263_p N_VGND_c_822_n 0.0104581f $X=5.1 $Y=0.515 $X2=0 $Y2=0
cc_258 N_A_83_21#_c_125_n N_VGND_c_822_n 0.0321116f $X=5.955 $Y=0.4 $X2=0 $Y2=0
cc_259 N_A_83_21#_c_127_n N_VGND_c_822_n 0.0121489f $X=3.37 $Y=0.34 $X2=0 $Y2=0
cc_260 N_A_83_21#_c_154_p N_A_457_47#_M1013_d 0.00332344f $X=4.125 $Y=0.34 $X2=0
+ $Y2=0
cc_261 N_A_83_21#_M1013_s N_A_457_47#_c_922_n 0.00548084f $X=3.25 $Y=0.235 $X2=0
+ $Y2=0
cc_262 N_A_83_21#_c_133_n N_A_457_47#_c_922_n 0.00467503f $X=4.125 $Y=1.782
+ $X2=0 $Y2=0
cc_263 N_A_83_21#_c_154_p N_A_457_47#_c_922_n 0.00375322f $X=4.125 $Y=0.34 $X2=0
+ $Y2=0
cc_264 N_A_83_21#_c_127_n N_A_457_47#_c_922_n 0.0199738f $X=3.37 $Y=0.34 $X2=0
+ $Y2=0
cc_265 N_A_83_21#_c_154_p N_A_457_47#_c_928_n 0.012764f $X=4.125 $Y=0.34 $X2=0
+ $Y2=0
cc_266 N_A_83_21#_c_125_n N_A_1077_47#_M1005_s 0.00329748f $X=5.955 $Y=0.4
+ $X2=-0.19 $Y2=-0.245
cc_267 N_A_83_21#_M1024_d N_A_1077_47#_c_947_n 0.00602235f $X=5.815 $Y=0.235
+ $X2=0 $Y2=0
cc_268 N_A_83_21#_c_125_n N_A_1077_47#_c_947_n 0.0417784f $X=5.955 $Y=0.4 $X2=0
+ $Y2=0
cc_269 N_A_83_21#_c_125_n N_A_1077_47#_c_948_n 0.0207418f $X=5.955 $Y=0.4 $X2=0
+ $Y2=0
cc_270 N_A2_M1017_g N_A1_M1015_g 0.0456599f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_271 A2 N_A1_c_351_n 0.0274335f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_272 A2 N_A1_c_340_n 0.0182412f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_273 N_A2_c_294_n N_A1_c_340_n 0.0219201f $X=2.64 $Y=1.352 $X2=0 $Y2=0
cc_274 N_A2_M1002_g N_VPWR_c_530_n 0.0151389f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A2_M1017_g N_VPWR_c_530_n 6.90674e-19 $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A2_M1002_g N_VPWR_c_531_n 6.42299e-19 $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A2_M1017_g N_VPWR_c_531_n 0.0120926f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_278 N_A2_M1002_g N_VPWR_c_536_n 0.00486043f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_279 N_A2_M1017_g N_VPWR_c_536_n 0.00486043f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_280 N_A2_M1002_g N_VPWR_c_526_n 0.00824727f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_281 N_A2_M1017_g N_VPWR_c_526_n 0.00824727f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_282 A2 N_X_c_636_n 0.0016503f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_283 N_A2_M1017_g N_A_457_367#_c_699_n 0.0125125f $X=2.64 $Y=2.465 $X2=0 $Y2=0
cc_284 N_A2_c_289_n N_VGND_c_810_n 0.0139645f $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_285 N_A2_c_291_n N_VGND_c_810_n 6.17119e-19 $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_286 N_A2_c_289_n N_VGND_c_811_n 5.68743e-19 $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_287 N_A2_c_291_n N_VGND_c_811_n 0.0112665f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_288 N_A2_c_289_n N_VGND_c_816_n 0.00486043f $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_289 N_A2_c_291_n N_VGND_c_816_n 0.00486043f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_290 N_A2_c_289_n N_VGND_c_822_n 0.00824727f $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_291 N_A2_c_291_n N_VGND_c_822_n 0.00455156f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_292 N_A2_c_291_n N_A_457_47#_c_922_n 0.0117904f $X=2.64 $Y=1.185 $X2=0 $Y2=0
cc_293 A2 N_A_457_47#_c_922_n 0.0476379f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_294 N_A2_c_294_n N_A_457_47#_c_922_n 0.00144925f $X=2.64 $Y=1.352 $X2=0 $Y2=0
cc_295 A2 N_A_457_47#_c_932_n 0.0146133f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_296 N_A2_c_294_n N_A_457_47#_c_932_n 0.00232957f $X=2.64 $Y=1.352 $X2=0 $Y2=0
cc_297 N_A1_c_339_n N_C1_c_382_n 0.0135768f $X=4.02 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_298 N_A1_c_340_n N_C1_c_387_n 0.0135768f $X=4.02 $Y=1.35 $X2=0 $Y2=0
cc_299 N_A1_M1015_g N_VPWR_c_531_n 0.012166f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A1_M1025_g N_VPWR_c_531_n 6.47302e-19 $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A1_M1015_g N_VPWR_c_532_n 0.00486043f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A1_M1025_g N_VPWR_c_532_n 0.00486043f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A1_M1015_g N_VPWR_c_533_n 6.50131e-19 $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A1_M1025_g N_VPWR_c_533_n 0.0142509f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A1_M1015_g N_VPWR_c_526_n 0.00824727f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_306 N_A1_M1025_g N_VPWR_c_526_n 0.00824727f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_307 N_A1_M1015_g N_A_457_367#_c_699_n 0.0125125f $X=3.07 $Y=2.465 $X2=0 $Y2=0
cc_308 N_A1_M1025_g N_A_457_367#_c_691_n 0.0143f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_309 N_A1_M1025_g N_A_457_367#_c_692_n 0.00298777f $X=3.5 $Y=2.465 $X2=0 $Y2=0
cc_310 N_A1_c_338_n N_VGND_c_811_n 0.00329003f $X=3.59 $Y=1.185 $X2=0 $Y2=0
cc_311 N_A1_c_338_n N_VGND_c_819_n 0.00359375f $X=3.59 $Y=1.185 $X2=0 $Y2=0
cc_312 N_A1_c_339_n N_VGND_c_819_n 0.00357877f $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_313 N_A1_c_338_n N_VGND_c_822_n 0.0068125f $X=3.59 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A1_c_339_n N_VGND_c_822_n 0.00537654f $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_315 N_A1_c_338_n N_A_457_47#_c_922_n 0.0118781f $X=3.59 $Y=1.185 $X2=0 $Y2=0
cc_316 N_A1_c_351_n N_A_457_47#_c_922_n 0.0202925f $X=3.835 $Y=1.35 $X2=0 $Y2=0
cc_317 N_A1_c_340_n N_A_457_47#_c_922_n 0.0140324f $X=4.02 $Y=1.35 $X2=0 $Y2=0
cc_318 N_A1_c_339_n N_A_457_47#_c_928_n 0.00460003f $X=4.02 $Y=1.185 $X2=0 $Y2=0
cc_319 N_A1_c_351_n N_A_457_47#_c_928_n 0.0168269f $X=3.835 $Y=1.35 $X2=0 $Y2=0
cc_320 N_A1_c_340_n N_A_457_47#_c_928_n 0.00229431f $X=4.02 $Y=1.35 $X2=0 $Y2=0
cc_321 N_C1_c_384_n N_B1_c_430_n 0.0153433f $X=4.88 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_322 N_C1_M1026_g N_B1_M1004_g 0.058668f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_323 C1 B1 0.0291708f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_324 N_C1_c_387_n B1 2.70249e-19 $X=4.88 $Y=1.36 $X2=0 $Y2=0
cc_325 C1 N_B1_c_435_n 0.0028427f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_326 N_C1_c_387_n N_B1_c_435_n 0.0163878f $X=4.88 $Y=1.36 $X2=0 $Y2=0
cc_327 N_C1_M1016_g N_VPWR_c_533_n 0.00676995f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_328 N_C1_M1016_g N_VPWR_c_539_n 0.00359964f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_329 N_C1_M1026_g N_VPWR_c_539_n 0.00359964f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_330 N_C1_M1016_g N_VPWR_c_526_n 0.00665257f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_331 N_C1_M1026_g N_VPWR_c_526_n 0.00537821f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_332 N_C1_M1016_g N_A_457_367#_c_691_n 0.00394375f $X=4.45 $Y=2.465 $X2=0
+ $Y2=0
cc_333 N_C1_M1016_g N_A_457_367#_c_692_n 0.00816609f $X=4.45 $Y=2.465 $X2=0
+ $Y2=0
cc_334 N_C1_M1016_g N_A_457_367#_c_705_n 0.0134612f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_335 N_C1_M1026_g N_A_457_367#_c_705_n 0.014279f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_336 N_C1_M1026_g N_A_457_367#_c_708_n 0.00200765f $X=4.88 $Y=2.465 $X2=0
+ $Y2=0
cc_337 N_C1_M1026_g N_A_457_367#_c_695_n 4.98432e-19 $X=4.88 $Y=2.465 $X2=0
+ $Y2=0
cc_338 N_C1_M1016_g N_A_822_367#_c_759_n 0.0106561f $X=4.45 $Y=2.465 $X2=0 $Y2=0
cc_339 N_C1_M1026_g N_A_822_367#_c_759_n 0.0106561f $X=4.88 $Y=2.465 $X2=0 $Y2=0
cc_340 N_C1_c_382_n N_VGND_c_812_n 0.00350831f $X=4.45 $Y=1.195 $X2=0 $Y2=0
cc_341 N_C1_c_384_n N_VGND_c_812_n 0.00350831f $X=4.88 $Y=1.195 $X2=0 $Y2=0
cc_342 N_C1_c_382_n N_VGND_c_819_n 0.00585385f $X=4.45 $Y=1.195 $X2=0 $Y2=0
cc_343 N_C1_c_384_n N_VGND_c_820_n 0.00585385f $X=4.88 $Y=1.195 $X2=0 $Y2=0
cc_344 N_C1_c_382_n N_VGND_c_822_n 0.00627451f $X=4.45 $Y=1.195 $X2=0 $Y2=0
cc_345 N_C1_c_384_n N_VGND_c_822_n 0.00627451f $X=4.88 $Y=1.195 $X2=0 $Y2=0
cc_346 B1 N_B2_M1006_g 0.00354769f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_347 N_B1_M1019_g N_B2_c_483_n 0.02745f $X=5.74 $Y=2.465 $X2=0 $Y2=0
cc_348 B1 N_B2_c_483_n 0.00982175f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_349 N_B1_c_435_n N_B2_c_483_n 0.0117871f $X=5.74 $Y=1.36 $X2=0 $Y2=0
cc_350 B1 N_B2_c_488_n 0.00419158f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_351 N_B1_M1004_g N_VPWR_c_539_n 0.00359964f $X=5.31 $Y=2.465 $X2=0 $Y2=0
cc_352 N_B1_M1019_g N_VPWR_c_539_n 0.0035993f $X=5.74 $Y=2.465 $X2=0 $Y2=0
cc_353 N_B1_M1004_g N_VPWR_c_526_n 0.00537821f $X=5.31 $Y=2.465 $X2=0 $Y2=0
cc_354 N_B1_M1019_g N_VPWR_c_526_n 0.00537818f $X=5.74 $Y=2.465 $X2=0 $Y2=0
cc_355 N_B1_M1004_g N_A_457_367#_c_705_n 0.0118214f $X=5.31 $Y=2.465 $X2=0 $Y2=0
cc_356 N_B1_M1004_g N_A_457_367#_c_708_n 0.0107219f $X=5.31 $Y=2.465 $X2=0 $Y2=0
cc_357 N_B1_M1019_g N_A_457_367#_c_694_n 0.0138387f $X=5.74 $Y=2.465 $X2=0 $Y2=0
cc_358 B1 N_A_457_367#_c_694_n 0.0371963f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_359 N_B1_c_435_n N_A_457_367#_c_694_n 0.00155936f $X=5.74 $Y=1.36 $X2=0 $Y2=0
cc_360 N_B1_M1004_g N_A_457_367#_c_695_n 0.00489838f $X=5.31 $Y=2.465 $X2=0
+ $Y2=0
cc_361 B1 N_A_457_367#_c_695_n 0.0208919f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_362 N_B1_c_435_n N_A_457_367#_c_695_n 0.00231808f $X=5.74 $Y=1.36 $X2=0 $Y2=0
cc_363 N_B1_M1004_g N_A_822_367#_c_759_n 0.0106551f $X=5.31 $Y=2.465 $X2=0 $Y2=0
cc_364 N_B1_M1019_g N_A_822_367#_c_759_n 0.013501f $X=5.74 $Y=2.465 $X2=0 $Y2=0
cc_365 N_B1_M1004_g N_A_822_367#_c_769_n 9.55923e-19 $X=5.31 $Y=2.465 $X2=0
+ $Y2=0
cc_366 N_B1_M1019_g N_A_822_367#_c_769_n 0.0090699f $X=5.74 $Y=2.465 $X2=0 $Y2=0
cc_367 N_B1_M1019_g N_A_822_367#_c_771_n 8.49285e-19 $X=5.74 $Y=2.465 $X2=0
+ $Y2=0
cc_368 N_B1_c_430_n N_VGND_c_820_n 0.00357877f $X=5.31 $Y=1.195 $X2=0 $Y2=0
cc_369 N_B1_c_432_n N_VGND_c_820_n 0.00357877f $X=5.74 $Y=1.195 $X2=0 $Y2=0
cc_370 N_B1_c_430_n N_VGND_c_822_n 0.00537654f $X=5.31 $Y=1.195 $X2=0 $Y2=0
cc_371 N_B1_c_432_n N_VGND_c_822_n 0.00665089f $X=5.74 $Y=1.195 $X2=0 $Y2=0
cc_372 N_B1_c_432_n N_A_1077_47#_c_947_n 0.0167471f $X=5.74 $Y=1.195 $X2=0 $Y2=0
cc_373 B1 N_A_1077_47#_c_947_n 0.0491164f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_374 N_B1_c_435_n N_A_1077_47#_c_947_n 0.00370003f $X=5.74 $Y=1.36 $X2=0 $Y2=0
cc_375 N_B1_c_432_n N_A_1077_47#_c_948_n 0.00339302f $X=5.74 $Y=1.195 $X2=0
+ $Y2=0
cc_376 N_B1_c_432_n N_A_1077_47#_c_951_n 0.00473581f $X=5.74 $Y=1.195 $X2=0
+ $Y2=0
cc_377 B1 N_A_1077_47#_c_951_n 0.00290769f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_378 N_B2_M1010_g N_VPWR_c_539_n 0.0035993f $X=6.17 $Y=2.465 $X2=0 $Y2=0
cc_379 N_B2_M1027_g N_VPWR_c_539_n 0.0035993f $X=6.6 $Y=2.465 $X2=0 $Y2=0
cc_380 N_B2_M1010_g N_VPWR_c_526_n 0.00537818f $X=6.17 $Y=2.465 $X2=0 $Y2=0
cc_381 N_B2_M1027_g N_VPWR_c_526_n 0.00665253f $X=6.6 $Y=2.465 $X2=0 $Y2=0
cc_382 N_B2_M1010_g N_A_457_367#_c_694_n 0.0163884f $X=6.17 $Y=2.465 $X2=0 $Y2=0
cc_383 N_B2_M1027_g N_A_457_367#_c_694_n 0.00302481f $X=6.6 $Y=2.465 $X2=0 $Y2=0
cc_384 N_B2_c_483_n N_A_457_367#_c_694_n 0.00398532f $X=7.12 $Y=1.5 $X2=0 $Y2=0
cc_385 N_B2_c_488_n N_A_457_367#_c_694_n 0.0040114f $X=6.985 $Y=1.577 $X2=0
+ $Y2=0
cc_386 N_B2_M1010_g N_A_822_367#_c_769_n 0.00814308f $X=6.17 $Y=2.465 $X2=0
+ $Y2=0
cc_387 N_B2_M1027_g N_A_822_367#_c_769_n 3.00577e-19 $X=6.6 $Y=2.465 $X2=0 $Y2=0
cc_388 N_B2_M1010_g N_A_822_367#_c_774_n 0.0105769f $X=6.17 $Y=2.465 $X2=0 $Y2=0
cc_389 N_B2_M1027_g N_A_822_367#_c_774_n 0.0105769f $X=6.6 $Y=2.465 $X2=0 $Y2=0
cc_390 N_B2_M1027_g N_A_822_367#_c_760_n 6.00691e-19 $X=6.6 $Y=2.465 $X2=0 $Y2=0
cc_391 N_B2_M1010_g N_A_822_367#_c_761_n 6.74942e-19 $X=6.17 $Y=2.465 $X2=0
+ $Y2=0
cc_392 N_B2_M1027_g N_A_822_367#_c_761_n 0.0139311f $X=6.6 $Y=2.465 $X2=0 $Y2=0
cc_393 N_B2_c_483_n N_A_822_367#_c_761_n 0.0018156f $X=7.12 $Y=1.5 $X2=0 $Y2=0
cc_394 N_B2_c_488_n N_A_822_367#_c_761_n 0.0259536f $X=6.985 $Y=1.577 $X2=0
+ $Y2=0
cc_395 N_B2_M1010_g N_A_822_367#_c_771_n 0.0025256f $X=6.17 $Y=2.465 $X2=0 $Y2=0
cc_396 N_B2_M1027_g N_A_822_367#_c_771_n 3.22649e-19 $X=6.6 $Y=2.465 $X2=0 $Y2=0
cc_397 N_B2_M1006_g N_VGND_c_813_n 0.0127147f $X=6.69 $Y=0.665 $X2=0 $Y2=0
cc_398 N_B2_M1022_g N_VGND_c_813_n 0.0127286f $X=7.12 $Y=0.665 $X2=0 $Y2=0
cc_399 N_B2_M1006_g N_VGND_c_820_n 0.00477554f $X=6.69 $Y=0.665 $X2=0 $Y2=0
cc_400 N_B2_M1022_g N_VGND_c_821_n 0.00477554f $X=7.12 $Y=0.665 $X2=0 $Y2=0
cc_401 N_B2_M1006_g N_VGND_c_822_n 0.00955784f $X=6.69 $Y=0.665 $X2=0 $Y2=0
cc_402 N_B2_M1022_g N_VGND_c_822_n 0.0092618f $X=7.12 $Y=0.665 $X2=0 $Y2=0
cc_403 N_B2_c_483_n N_A_1077_47#_c_947_n 0.00673362f $X=7.12 $Y=1.5 $X2=0 $Y2=0
cc_404 N_B2_M1006_g N_A_1077_47#_c_949_n 0.0155838f $X=6.69 $Y=0.665 $X2=0 $Y2=0
cc_405 N_B2_M1022_g N_A_1077_47#_c_949_n 0.0152307f $X=7.12 $Y=0.665 $X2=0 $Y2=0
cc_406 B2 N_A_1077_47#_c_949_n 0.0414175f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_407 N_B2_c_483_n N_A_1077_47#_c_949_n 0.00714658f $X=7.12 $Y=1.5 $X2=0 $Y2=0
cc_408 N_B2_c_488_n N_A_1077_47#_c_949_n 0.0263729f $X=6.985 $Y=1.577 $X2=0
+ $Y2=0
cc_409 N_B2_c_483_n N_A_1077_47#_c_951_n 0.0106437f $X=7.12 $Y=1.5 $X2=0 $Y2=0
cc_410 N_VPWR_c_526_n N_X_M1007_s 0.00571434f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_411 N_VPWR_c_526_n N_X_M1018_s 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_412 N_VPWR_M1007_d N_X_c_640_n 2.33864e-19 $X=0.15 $Y=1.835 $X2=0 $Y2=0
cc_413 N_VPWR_c_528_n N_X_c_640_n 0.00362085f $X=0.275 $Y=2.18 $X2=0 $Y2=0
cc_414 N_VPWR_M1007_d N_X_c_641_n 0.00247068f $X=0.15 $Y=1.835 $X2=0 $Y2=0
cc_415 N_VPWR_c_528_n N_X_c_641_n 0.0203341f $X=0.275 $Y=2.18 $X2=0 $Y2=0
cc_416 N_VPWR_c_538_n N_X_c_673_n 0.0120977f $X=0.97 $Y=3.33 $X2=0 $Y2=0
cc_417 N_VPWR_c_526_n N_X_c_673_n 0.00691495f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_418 N_VPWR_M1008_d N_X_c_642_n 0.00176461f $X=0.995 $Y=1.835 $X2=0 $Y2=0
cc_419 N_VPWR_c_529_n N_X_c_642_n 0.0170777f $X=1.135 $Y=2.18 $X2=0 $Y2=0
cc_420 N_VPWR_c_534_n N_X_c_677_n 0.0124525f $X=1.83 $Y=3.33 $X2=0 $Y2=0
cc_421 N_VPWR_c_526_n N_X_c_677_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_422 N_VPWR_c_526_n N_A_457_367#_M1002_d 0.00536646f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_423 N_VPWR_c_526_n N_A_457_367#_M1015_s 0.00536823f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_526_n N_A_457_367#_M1004_d 0.00225465f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_526_n N_A_457_367#_M1010_d 0.00225465f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_536_n N_A_457_367#_c_737_n 0.0124525f $X=2.69 $Y=3.33 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_526_n N_A_457_367#_c_737_n 0.00730901f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_428 N_VPWR_M1017_s N_A_457_367#_c_699_n 0.00352528f $X=2.715 $Y=1.835 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_531_n N_A_457_367#_c_699_n 0.0171443f $X=2.855 $Y=2.48 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_532_n N_A_457_367#_c_741_n 0.0117038f $X=3.55 $Y=3.33 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_526_n N_A_457_367#_c_741_n 0.00727431f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_432 N_VPWR_M1025_d N_A_457_367#_c_691_n 0.00498953f $X=3.575 $Y=1.835 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_533_n N_A_457_367#_c_691_n 0.0220026f $X=3.715 $Y=2.47 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_533_n N_A_457_367#_c_692_n 0.00448147f $X=3.715 $Y=2.47 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_533_n N_A_457_367#_c_693_n 0.0139f $X=3.715 $Y=2.47 $X2=0 $Y2=0
cc_436 N_VPWR_c_526_n N_A_822_367#_M1016_d 0.00215439f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_437 N_VPWR_c_526_n N_A_822_367#_M1026_d 0.00223855f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_526_n N_A_822_367#_M1019_s 0.00223819f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_526_n N_A_822_367#_M1027_s 0.00215406f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_533_n N_A_822_367#_c_759_n 0.0227306f $X=3.715 $Y=2.47 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_539_n N_A_822_367#_c_759_n 0.0935607f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_526_n N_A_822_367#_c_759_n 0.062161f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_443 N_VPWR_c_539_n N_A_822_367#_c_774_n 0.0280869f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_526_n N_A_822_367#_c_774_n 0.0186561f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_539_n N_A_822_367#_c_760_n 0.0199166f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_446 N_VPWR_c_526_n N_A_822_367#_c_760_n 0.0125808f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_447 N_VPWR_c_539_n N_A_822_367#_c_771_n 0.0179231f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_448 N_VPWR_c_526_n N_A_822_367#_c_771_n 0.0123929f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_449 N_X_c_635_n N_VGND_M1003_s 2.33864e-19 $X=0.61 $Y=1.145 $X2=-0.19
+ $Y2=-0.245
cc_450 N_X_c_638_n N_VGND_M1003_s 0.00211783f $X=0.222 $Y=1.23 $X2=-0.19
+ $Y2=-0.245
cc_451 N_X_c_636_n N_VGND_M1012_s 0.00176922f $X=1.47 $Y=1.137 $X2=0 $Y2=0
cc_452 N_X_c_635_n N_VGND_c_808_n 0.00362085f $X=0.61 $Y=1.145 $X2=0 $Y2=0
cc_453 N_X_c_638_n N_VGND_c_808_n 0.0203341f $X=0.222 $Y=1.23 $X2=0 $Y2=0
cc_454 N_X_c_636_n N_VGND_c_809_n 0.0171764f $X=1.47 $Y=1.137 $X2=0 $Y2=0
cc_455 N_X_c_685_p N_VGND_c_814_n 0.0124525f $X=1.565 $Y=0.42 $X2=0 $Y2=0
cc_456 N_X_c_686_p N_VGND_c_818_n 0.0124525f $X=0.705 $Y=0.42 $X2=0 $Y2=0
cc_457 N_X_M1003_d N_VGND_c_822_n 0.00536646f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_458 N_X_M1014_d N_VGND_c_822_n 0.00536646f $X=1.425 $Y=0.235 $X2=0 $Y2=0
cc_459 N_X_c_686_p N_VGND_c_822_n 0.00730901f $X=0.705 $Y=0.42 $X2=0 $Y2=0
cc_460 N_X_c_685_p N_VGND_c_822_n 0.00730901f $X=1.565 $Y=0.42 $X2=0 $Y2=0
cc_461 N_A_457_367#_c_691_n N_A_822_367#_M1016_d 0.00561479f $X=4.07 $Y=2.13
+ $X2=-0.19 $Y2=1.655
cc_462 N_A_457_367#_c_692_n N_A_822_367#_M1016_d 0.00384659f $X=4.192 $Y=2.445
+ $X2=-0.19 $Y2=1.655
cc_463 N_A_457_367#_c_693_n N_A_822_367#_M1016_d 0.00300215f $X=4.315 $Y=2.53
+ $X2=-0.19 $Y2=1.655
cc_464 N_A_457_367#_c_705_n N_A_822_367#_M1026_d 0.00805622f $X=5.36 $Y=2.53
+ $X2=0 $Y2=0
cc_465 N_A_457_367#_c_694_n N_A_822_367#_M1019_s 0.00180746f $X=6.29 $Y=1.79
+ $X2=0 $Y2=0
cc_466 N_A_457_367#_M1004_d N_A_822_367#_c_759_n 0.00341017f $X=5.385 $Y=1.835
+ $X2=0 $Y2=0
cc_467 N_A_457_367#_c_705_n N_A_822_367#_c_759_n 0.0681402f $X=5.36 $Y=2.53
+ $X2=0 $Y2=0
cc_468 N_A_457_367#_c_693_n N_A_822_367#_c_759_n 0.0196292f $X=4.315 $Y=2.53
+ $X2=0 $Y2=0
cc_469 N_A_457_367#_c_694_n N_A_822_367#_c_769_n 0.0163515f $X=6.29 $Y=1.79
+ $X2=0 $Y2=0
cc_470 N_A_457_367#_M1010_d N_A_822_367#_c_774_n 0.00335807f $X=6.245 $Y=1.835
+ $X2=0 $Y2=0
cc_471 N_A_457_367#_c_757_p N_A_822_367#_c_774_n 0.012662f $X=6.385 $Y=1.98
+ $X2=0 $Y2=0
cc_472 N_A_457_367#_c_694_n N_A_1077_47#_c_951_n 0.00458286f $X=6.29 $Y=1.79
+ $X2=0 $Y2=0
cc_473 N_VGND_c_822_n N_A_457_47#_M1000_d 0.00408812f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_474 N_VGND_c_822_n N_A_457_47#_M1013_d 0.00224381f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_475 N_VGND_c_816_n N_A_457_47#_c_942_n 0.0124525f $X=2.69 $Y=0 $X2=0 $Y2=0
cc_476 N_VGND_c_822_n N_A_457_47#_c_942_n 0.00730901f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_477 N_VGND_M1009_s N_A_457_47#_c_922_n 0.00512142f $X=2.715 $Y=0.235 $X2=0
+ $Y2=0
cc_478 N_VGND_c_811_n N_A_457_47#_c_922_n 0.021529f $X=2.855 $Y=0.51 $X2=0 $Y2=0
cc_479 N_VGND_c_822_n N_A_457_47#_c_922_n 0.0134553f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_480 N_VGND_c_822_n N_A_1077_47#_M1005_s 0.00225186f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_481 N_VGND_c_822_n N_A_1077_47#_M1006_s 0.00368844f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_482 N_VGND_c_822_n N_A_1077_47#_M1022_s 0.00368844f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_483 N_VGND_c_820_n N_A_1077_47#_c_947_n 0.00327408f $X=6.74 $Y=0 $X2=0 $Y2=0
cc_484 N_VGND_c_822_n N_A_1077_47#_c_947_n 0.00677337f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_485 N_VGND_c_820_n N_A_1077_47#_c_948_n 0.0178111f $X=6.74 $Y=0 $X2=0 $Y2=0
cc_486 N_VGND_c_822_n N_A_1077_47#_c_948_n 0.0100304f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_M1006_d N_A_1077_47#_c_949_n 0.00176461f $X=6.765 $Y=0.245 $X2=0
+ $Y2=0
cc_488 N_VGND_c_813_n N_A_1077_47#_c_949_n 0.0170777f $X=6.905 $Y=0.39 $X2=0
+ $Y2=0
cc_489 N_VGND_c_821_n N_A_1077_47#_c_950_n 0.0178111f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_490 N_VGND_c_822_n N_A_1077_47#_c_950_n 0.0100304f $X=7.44 $Y=0 $X2=0 $Y2=0
