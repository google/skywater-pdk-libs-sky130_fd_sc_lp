* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fa_lp A B CIN VGND VNB VPB VPWR COUT SUM
X0 a_1049_419# CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_84_209# CIN a_458_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_1720_419# B a_1818_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VPWR A a_458_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_1005_141# CIN VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1574_141# CIN a_1686_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_1574_141# a_1956_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1574_141# CIN a_1720_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VPWR a_1574_141# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_1956_66# a_1574_141# SUM VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_458_409# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 VGND A a_1005_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1049_419# a_84_209# a_1574_141# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_1686_141# B a_1764_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND A a_577_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 COUT a_84_209# a_134_85# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_245_409# B a_84_209# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_134_85# a_84_209# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 COUT a_84_209# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X19 a_245_409# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 VPWR A a_1049_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 a_1764_141# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1005_141# a_84_209# a_1574_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_577_141# B a_84_209# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VGND B a_1005_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_355_141# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_355_141# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_1818_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X28 a_84_209# CIN a_355_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR B a_1049_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
