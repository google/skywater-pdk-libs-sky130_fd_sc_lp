* File: sky130_fd_sc_lp__and4_lp2.spice
* Created: Wed Sep  2 09:33:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4_lp2.pex.spice"
.subckt sky130_fd_sc_lp__and4_lp2  VNB VPB D C B A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1005 A_114_47# N_A_84_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_84_21#_M1008_g A_114_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1004 A_294_47# N_D_M1004_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=31.428 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 A_372_47# N_C_M1002_g A_294_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.5 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1003 A_450_47# N_B_M1003_g A_372_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_84_21#_M1000_d N_A_M1000_g A_450_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_84_21#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.25 W=1
+ AD=0.1575 AS=0.285 PD=1.315 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1009 N_A_84_21#_M1009_d N_D_M1009_g N_VPWR_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.1575 PD=1.28 PS=1.315 NRD=0 NRS=6.8753 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_A_84_21#_M1009_d VPB PHIGHVT L=0.25 W=1
+ AD=0.18 AS=0.14 PD=1.36 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1007 N_A_84_21#_M1007_d N_B_M1007_g N_VPWR_M1006_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.18 PD=1.28 PS=1.36 NRD=0 NRS=15.7403 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_84_21#_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX11_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__and4_lp2.pxi.spice"
*
.ends
*
*
