* File: sky130_fd_sc_lp__o221ai_m.spice
* Created: Wed Sep  2 10:19:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221ai_m.pex.spice"
.subckt sky130_fd_sc_lp__o221ai_m  VNB VPB C1 B1 A2 A1 B2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* B2	B2
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1000 N_A_148_47#_M1000_d N_C1_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_234_47#_M1005_d N_B1_M1005_g N_A_148_47#_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.06195 AS=0.0588 PD=0.715 PS=0.7 NRD=4.284 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_234_47#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.06195 PD=0.84 PS=0.715 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_234_47#_M1003_d N_A1_M1003_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0882 PD=0.7 PS=0.84 NRD=0 NRS=34.284 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_148_47#_M1004_d N_B2_M1004_g N_A_234_47#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_C1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0915 AS=0.1113 PD=0.88 PS=1.37 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1009 A_245_480# N_B1_M1009_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0915 PD=0.63 PS=0.88 NRD=23.443 NRS=30.4759 M=1 R=2.8
+ SA=75000.7 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g A_245_480# VPB PHIGHVT L=0.15 W=0.42 AD=0.109325
+ AS=0.0441 PD=0.975 PS=0.63 NRD=46.886 NRS=23.443 M=1 R=2.8 SA=75001.1 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1007 A_441_463# N_A2_M1007_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.109325 PD=0.63 PS=0.975 NRD=23.443 NRS=44.5417 M=1 R=2.8 SA=75001.4
+ SB=75000.5 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_441_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o221ai_m.pxi.spice"
*
.ends
*
*
