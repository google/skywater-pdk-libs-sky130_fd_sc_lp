* File: sky130_fd_sc_lp__dfrtp_1.pxi.spice
* Created: Wed Sep  2 09:43:41 2020
* 
x_PM_SKY130_FD_SC_LP__DFRTP_1%CLK N_CLK_M1013_g N_CLK_M1020_g N_CLK_c_236_n
+ N_CLK_c_241_n CLK CLK N_CLK_c_237_n N_CLK_c_238_n
+ PM_SKY130_FD_SC_LP__DFRTP_1%CLK
x_PM_SKY130_FD_SC_LP__DFRTP_1%A_27_114# N_A_27_114#_M1013_s N_A_27_114#_M1020_s
+ N_A_27_114#_c_272_n N_A_27_114#_M1006_g N_A_27_114#_M1026_g
+ N_A_27_114#_M1004_g N_A_27_114#_M1009_g N_A_27_114#_M1011_g
+ N_A_27_114#_c_274_n N_A_27_114#_M1030_g N_A_27_114#_c_275_n
+ N_A_27_114#_c_276_n N_A_27_114#_c_310_n N_A_27_114#_c_277_n
+ N_A_27_114#_c_278_n N_A_27_114#_c_279_n N_A_27_114#_c_311_n
+ N_A_27_114#_c_280_n N_A_27_114#_c_281_n N_A_27_114#_c_282_n
+ N_A_27_114#_c_283_n N_A_27_114#_c_284_n N_A_27_114#_c_285_n
+ N_A_27_114#_c_286_n N_A_27_114#_c_287_n N_A_27_114#_c_288_n
+ N_A_27_114#_c_289_n N_A_27_114#_c_290_n N_A_27_114#_c_291_n
+ N_A_27_114#_c_292_n N_A_27_114#_c_293_n N_A_27_114#_c_294_n
+ N_A_27_114#_c_312_n N_A_27_114#_c_295_n N_A_27_114#_c_296_n
+ N_A_27_114#_c_297_n N_A_27_114#_c_298_n N_A_27_114#_c_299_n
+ N_A_27_114#_c_300_n N_A_27_114#_c_301_n N_A_27_114#_c_314_n
+ N_A_27_114#_c_315_n N_A_27_114#_c_302_n N_A_27_114#_c_303_n
+ N_A_27_114#_c_304_n N_A_27_114#_c_305_n PM_SKY130_FD_SC_LP__DFRTP_1%A_27_114#
x_PM_SKY130_FD_SC_LP__DFRTP_1%D N_D_M1021_g N_D_M1002_g D N_D_c_542_n
+ N_D_c_543_n PM_SKY130_FD_SC_LP__DFRTP_1%D
x_PM_SKY130_FD_SC_LP__DFRTP_1%A_196_462# N_A_196_462#_M1026_d
+ N_A_196_462#_M1006_d N_A_196_462#_M1015_g N_A_196_462#_M1027_g
+ N_A_196_462#_M1031_g N_A_196_462#_c_585_n N_A_196_462#_c_586_n
+ N_A_196_462#_M1005_g N_A_196_462#_c_594_n N_A_196_462#_c_595_n
+ N_A_196_462#_c_587_n N_A_196_462#_c_597_n N_A_196_462#_c_598_n
+ N_A_196_462#_c_599_n N_A_196_462#_c_588_n N_A_196_462#_c_589_n
+ N_A_196_462#_c_601_n N_A_196_462#_c_602_n N_A_196_462#_c_603_n
+ N_A_196_462#_c_604_n N_A_196_462#_c_707_p N_A_196_462#_c_605_n
+ N_A_196_462#_c_590_n N_A_196_462#_c_607_n
+ PM_SKY130_FD_SC_LP__DFRTP_1%A_196_462#
x_PM_SKY130_FD_SC_LP__DFRTP_1%A_695_375# N_A_695_375#_M1028_d
+ N_A_695_375#_M1012_d N_A_695_375#_M1029_g N_A_695_375#_c_790_n
+ N_A_695_375#_c_791_n N_A_695_375#_M1018_g N_A_695_375#_c_782_n
+ N_A_695_375#_c_783_n N_A_695_375#_c_784_n N_A_695_375#_c_794_n
+ N_A_695_375#_c_785_n N_A_695_375#_c_786_n N_A_695_375#_c_787_n
+ N_A_695_375#_c_788_n N_A_695_375#_c_809_n
+ PM_SKY130_FD_SC_LP__DFRTP_1%A_695_375#
x_PM_SKY130_FD_SC_LP__DFRTP_1%RESET_B N_RESET_B_M1007_g N_RESET_B_c_889_n
+ N_RESET_B_c_890_n N_RESET_B_M1010_g N_RESET_B_c_892_n N_RESET_B_c_900_n
+ N_RESET_B_M1022_g N_RESET_B_c_901_n N_RESET_B_c_902_n N_RESET_B_M1014_g
+ N_RESET_B_M1001_g N_RESET_B_M1003_g N_RESET_B_c_895_n N_RESET_B_c_905_n
+ N_RESET_B_c_906_n N_RESET_B_c_907_n N_RESET_B_c_896_n N_RESET_B_c_909_n
+ N_RESET_B_c_976_p N_RESET_B_c_910_n N_RESET_B_c_933_n RESET_B
+ N_RESET_B_c_897_n N_RESET_B_c_898_n RESET_B
+ PM_SKY130_FD_SC_LP__DFRTP_1%RESET_B
x_PM_SKY130_FD_SC_LP__DFRTP_1%A_559_533# N_A_559_533#_M1004_d
+ N_A_559_533#_M1015_d N_A_559_533#_M1022_d N_A_559_533#_c_1075_n
+ N_A_559_533#_M1028_g N_A_559_533#_c_1080_n N_A_559_533#_M1012_g
+ N_A_559_533#_c_1099_n N_A_559_533#_c_1082_n N_A_559_533#_c_1101_n
+ N_A_559_533#_c_1083_n N_A_559_533#_c_1084_n N_A_559_533#_c_1076_n
+ N_A_559_533#_c_1085_n N_A_559_533#_c_1086_n N_A_559_533#_c_1087_n
+ N_A_559_533#_c_1088_n N_A_559_533#_c_1125_n N_A_559_533#_c_1089_n
+ N_A_559_533#_c_1077_n N_A_559_533#_c_1090_n N_A_559_533#_c_1091_n
+ N_A_559_533#_c_1078_n N_A_559_533#_c_1079_n
+ PM_SKY130_FD_SC_LP__DFRTP_1%A_559_533#
x_PM_SKY130_FD_SC_LP__DFRTP_1%A_1467_419# N_A_1467_419#_M1025_d
+ N_A_1467_419#_M1003_d N_A_1467_419#_M1016_g N_A_1467_419#_M1000_g
+ N_A_1467_419#_c_1231_n N_A_1467_419#_c_1232_n N_A_1467_419#_c_1233_n
+ N_A_1467_419#_c_1227_n N_A_1467_419#_c_1234_n N_A_1467_419#_c_1228_n
+ N_A_1467_419#_c_1236_n PM_SKY130_FD_SC_LP__DFRTP_1%A_1467_419#
x_PM_SKY130_FD_SC_LP__DFRTP_1%A_1247_89# N_A_1247_89#_M1031_d
+ N_A_1247_89#_M1011_d N_A_1247_89#_c_1304_n N_A_1247_89#_M1025_g
+ N_A_1247_89#_M1008_g N_A_1247_89#_c_1305_n N_A_1247_89#_c_1306_n
+ N_A_1247_89#_M1023_g N_A_1247_89#_M1017_g N_A_1247_89#_c_1309_n
+ N_A_1247_89#_c_1318_n N_A_1247_89#_c_1310_n N_A_1247_89#_c_1311_n
+ N_A_1247_89#_c_1319_n N_A_1247_89#_c_1312_n N_A_1247_89#_c_1313_n
+ N_A_1247_89#_c_1314_n N_A_1247_89#_c_1315_n
+ PM_SKY130_FD_SC_LP__DFRTP_1%A_1247_89#
x_PM_SKY130_FD_SC_LP__DFRTP_1%A_1832_367# N_A_1832_367#_M1017_s
+ N_A_1832_367#_M1023_s N_A_1832_367#_M1024_g N_A_1832_367#_M1019_g
+ N_A_1832_367#_c_1419_n N_A_1832_367#_c_1425_n N_A_1832_367#_c_1420_n
+ N_A_1832_367#_c_1421_n N_A_1832_367#_c_1422_n N_A_1832_367#_c_1423_n
+ PM_SKY130_FD_SC_LP__DFRTP_1%A_1832_367#
x_PM_SKY130_FD_SC_LP__DFRTP_1%VPWR N_VPWR_M1020_d N_VPWR_M1007_d N_VPWR_M1029_d
+ N_VPWR_M1012_s N_VPWR_M1016_d N_VPWR_M1008_d N_VPWR_M1023_d N_VPWR_c_1467_n
+ N_VPWR_c_1468_n N_VPWR_c_1469_n N_VPWR_c_1470_n N_VPWR_c_1471_n
+ N_VPWR_c_1472_n N_VPWR_c_1473_n N_VPWR_c_1474_n N_VPWR_c_1475_n
+ N_VPWR_c_1476_n N_VPWR_c_1477_n N_VPWR_c_1478_n VPWR N_VPWR_c_1479_n
+ N_VPWR_c_1480_n N_VPWR_c_1481_n N_VPWR_c_1482_n N_VPWR_c_1483_n
+ N_VPWR_c_1466_n N_VPWR_c_1485_n N_VPWR_c_1486_n N_VPWR_c_1487_n
+ N_VPWR_c_1488_n PM_SKY130_FD_SC_LP__DFRTP_1%VPWR
x_PM_SKY130_FD_SC_LP__DFRTP_1%A_304_533# N_A_304_533#_M1002_d
+ N_A_304_533#_M1007_s N_A_304_533#_M1021_d N_A_304_533#_c_1606_n
+ N_A_304_533#_c_1607_n N_A_304_533#_c_1608_n N_A_304_533#_c_1674_n
+ N_A_304_533#_c_1609_n N_A_304_533#_c_1605_n N_A_304_533#_c_1611_n
+ N_A_304_533#_c_1612_n N_A_304_533#_c_1613_n
+ PM_SKY130_FD_SC_LP__DFRTP_1%A_304_533#
x_PM_SKY130_FD_SC_LP__DFRTP_1%Q N_Q_M1019_d N_Q_M1024_d N_Q_c_1684_n
+ N_Q_c_1685_n Q Q Q Q PM_SKY130_FD_SC_LP__DFRTP_1%Q
x_PM_SKY130_FD_SC_LP__DFRTP_1%VGND N_VGND_M1013_d N_VGND_M1010_s N_VGND_M1014_d
+ N_VGND_M1000_d N_VGND_M1017_d N_VGND_c_1697_n N_VGND_c_1698_n N_VGND_c_1699_n
+ N_VGND_c_1700_n N_VGND_c_1701_n N_VGND_c_1702_n VGND N_VGND_c_1703_n
+ N_VGND_c_1704_n N_VGND_c_1705_n N_VGND_c_1706_n N_VGND_c_1707_n
+ N_VGND_c_1708_n N_VGND_c_1709_n N_VGND_c_1710_n N_VGND_c_1711_n
+ N_VGND_c_1712_n PM_SKY130_FD_SC_LP__DFRTP_1%VGND
cc_1 VNB N_CLK_M1013_g 0.0481971f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.78
cc_2 VNB N_CLK_c_236_n 0.00323314f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.955
cc_3 VNB N_CLK_c_237_n 0.0188165f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_4 VNB N_CLK_c_238_n 0.0106096f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_5 VNB N_A_27_114#_c_272_n 0.0210472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_114#_M1009_g 0.0029533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_114#_c_274_n 0.0178453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_114#_c_275_n 0.00806754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_114#_c_276_n 0.0193914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_114#_c_277_n 0.00615948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_114#_c_278_n 0.0103811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_114#_c_279_n 0.00232923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_114#_c_280_n 0.0018044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_114#_c_281_n 0.0151462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_114#_c_282_n 0.00286516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_114#_c_283_n 0.00531767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_114#_c_284_n 0.0133101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_114#_c_285_n 0.00389653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_114#_c_286_n 6.79085e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_114#_c_287_n 0.00795713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_114#_c_288_n 0.00224585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_114#_c_289_n 0.00474729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_114#_c_290_n 0.0388787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_114#_c_291_n 0.00353494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_114#_c_292_n 0.0011223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_114#_c_293_n 0.0101746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_114#_c_294_n 0.0465667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_114#_c_295_n 0.00807085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_114#_c_296_n 0.0255263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_114#_c_297_n 7.17315e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_114#_c_298_n 0.00107849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_114#_c_299_n 0.018078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_114#_c_300_n 0.00334703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_114#_c_301_n 0.0011466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_114#_c_302_n 0.00466019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_114#_c_303_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_114#_c_304_n 0.0193678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_114#_c_305_n 0.0152115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_D_M1002_g 0.0294199f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.63
cc_40 VNB N_D_c_542_n 0.0244567f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_41 VNB N_D_c_543_n 0.00378305f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_42 VNB N_A_196_462#_M1027_g 0.0177192f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_43 VNB N_A_196_462#_M1031_g 0.030803f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_44 VNB N_A_196_462#_c_585_n 0.061204f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_45 VNB N_A_196_462#_c_586_n 0.00859381f $X=-0.19 $Y=-0.245 $X2=0.282
+ $Y2=1.615
cc_46 VNB N_A_196_462#_c_587_n 0.013695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_196_462#_c_588_n 3.60697e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_196_462#_c_589_n 0.0309113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_196_462#_c_590_n 0.00146971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_695_375#_M1018_g 0.0190438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_695_375#_c_782_n 0.00844421f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.615
cc_52 VNB N_A_695_375#_c_783_n 0.0115515f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.615
cc_53 VNB N_A_695_375#_c_784_n 0.0102589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_695_375#_c_785_n 0.00182429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_695_375#_c_786_n 0.0162307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_695_375#_c_787_n 7.37641e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_695_375#_c_788_n 0.00293346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_M1007_g 0.0798099f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.78
cc_59 VNB N_RESET_B_c_889_n 0.0225367f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.12
cc_60 VNB N_RESET_B_c_890_n 0.0128168f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.63
cc_61 VNB N_RESET_B_M1010_g 0.0288417f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_62 VNB N_RESET_B_c_892_n 0.169186f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.955
cc_63 VNB N_RESET_B_M1014_g 0.0432348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_RESET_B_M1001_g 0.034336f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=2.035
cc_65 VNB N_RESET_B_c_895_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_RESET_B_c_896_n 0.00215951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_RESET_B_c_897_n 0.00270331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_RESET_B_c_898_n 0.0125006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_559_533#_c_1075_n 0.0216785f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=2.12
cc_70 VNB N_A_559_533#_c_1076_n 0.0049201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_559_533#_c_1077_n 2.20412e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_559_533#_c_1078_n 0.0425957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_559_533#_c_1079_n 0.0148049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1467_419#_M1000_g 0.0430821f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_75 VNB N_A_1467_419#_c_1227_n 0.015014f $X=-0.19 $Y=-0.245 $X2=0.282
+ $Y2=2.035
cc_76 VNB N_A_1467_419#_c_1228_n 0.00805764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1247_89#_c_1304_n 0.0217027f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.63
cc_78 VNB N_A_1247_89#_c_1305_n 0.0496641f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_79 VNB N_A_1247_89#_c_1306_n 0.028256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1247_89#_M1023_g 0.0154203f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_81 VNB N_A_1247_89#_M1017_g 0.0240627f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.665
cc_82 VNB N_A_1247_89#_c_1309_n 0.0250027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1247_89#_c_1310_n 0.00268567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1247_89#_c_1311_n 0.0387684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1247_89#_c_1312_n 0.00128739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1247_89#_c_1313_n 0.00138645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1247_89#_c_1314_n 0.00224376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1247_89#_c_1315_n 0.0264435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1832_367#_c_1419_n 0.0168763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1832_367#_c_1420_n 0.00336326f $X=-0.19 $Y=-0.245 $X2=0.282
+ $Y2=2.035
cc_91 VNB N_A_1832_367#_c_1421_n 0.0290259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1832_367#_c_1422_n 0.00258614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1832_367#_c_1423_n 0.0204406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VPWR_c_1466_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_304_533#_c_1605_n 0.0097213f $X=-0.19 $Y=-0.245 $X2=0.282
+ $Y2=2.035
cc_96 VNB Q 0.0581212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1697_n 0.0189118f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_98 VNB N_VGND_c_1698_n 0.0089408f $X=-0.19 $Y=-0.245 $X2=0.282 $Y2=1.665
cc_99 VNB N_VGND_c_1699_n 0.0206764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1700_n 0.0106566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1701_n 0.05223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1702_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1703_n 0.019573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1704_n 0.0307173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1705_n 0.0694445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1706_n 0.0538347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1707_n 0.0167577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1708_n 0.573213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1709_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1710_n 0.00585925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1711_n 0.0129533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1712_n 0.006464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VPB N_CLK_M1020_g 0.0283555f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.63
cc_114 VPB N_CLK_c_236_n 0.0247874f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_115 VPB N_CLK_c_241_n 0.0188165f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_116 VPB N_CLK_c_238_n 0.0208317f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_117 VPB N_A_27_114#_M1006_g 0.0399341f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_118 VPB N_A_27_114#_M1009_g 0.0632124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_27_114#_M1011_g 0.0225691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_27_114#_c_275_n 0.0171453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_27_114#_c_310_n 0.0041814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_27_114#_c_311_n 0.00377063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_27_114#_c_312_n 0.0304915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_27_114#_c_297_n 0.00334346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_27_114#_c_314_n 0.00135413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_27_114#_c_315_n 0.0371187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_27_114#_c_302_n 0.00167956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_D_M1021_g 0.0522229f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.78
cc_129 VPB N_D_c_542_n 0.0245939f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_130 VPB N_D_c_543_n 0.0074657f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_131 VPB N_A_196_462#_M1015_g 0.0234837f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_132 VPB N_A_196_462#_c_585_n 0.00944119f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.615
cc_133 VPB N_A_196_462#_M1005_g 0.0348803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_196_462#_c_594_n 0.0219798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_196_462#_c_595_n 0.00912064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_196_462#_c_587_n 0.0072546f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_196_462#_c_597_n 0.0160583f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_196_462#_c_598_n 0.0312687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_196_462#_c_599_n 0.00842961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_196_462#_c_588_n 0.00381616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_196_462#_c_601_n 0.031982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_196_462#_c_602_n 0.00420229f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_196_462#_c_603_n 0.0238404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_196_462#_c_604_n 6.84794e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_196_462#_c_605_n 0.0264966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_196_462#_c_590_n 0.006464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_196_462#_c_607_n 0.0217007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_695_375#_M1029_g 0.0450758f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_149 VPB N_A_695_375#_c_790_n 0.0536938f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_150 VPB N_A_695_375#_c_791_n 0.012181f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_151 VPB N_A_695_375#_c_782_n 0.0166986f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_152 VPB N_A_695_375#_c_783_n 0.00679601f $X=-0.19 $Y=1.655 $X2=0.282
+ $Y2=1.615
cc_153 VPB N_A_695_375#_c_794_n 0.0075829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_695_375#_c_788_n 6.41825e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_RESET_B_M1007_g 0.0739316f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.78
cc_156 VPB N_RESET_B_c_900_n 0.0201938f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_157 VPB N_RESET_B_c_901_n 0.0225517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_RESET_B_c_902_n 0.00881958f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_159 VPB N_RESET_B_M1014_g 0.0441931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_M1003_g 0.0475849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_RESET_B_c_905_n 0.0180666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_RESET_B_c_906_n 0.00872221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_RESET_B_c_907_n 0.00413066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_RESET_B_c_896_n 0.00137539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_RESET_B_c_909_n 0.00531886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_RESET_B_c_910_n 0.059003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_RESET_B_c_897_n 0.00197619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_RESET_B_c_898_n 0.0216318f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_559_533#_c_1080_n 0.0222427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_559_533#_M1012_g 0.0230242f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_171 VPB N_A_559_533#_c_1082_n 2.91352e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_559_533#_c_1083_n 0.00699968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_559_533#_c_1084_n 0.00183865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_559_533#_c_1085_n 2.96747e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_559_533#_c_1086_n 0.00468957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_559_533#_c_1087_n 0.0116051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_559_533#_c_1088_n 0.00389911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_559_533#_c_1089_n 4.29785e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_559_533#_c_1090_n 0.00338439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_559_533#_c_1091_n 0.0347696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_559_533#_c_1079_n 0.00657257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_1467_419#_M1016_g 0.0228055f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.615
cc_183 VPB N_A_1467_419#_M1000_g 0.0210653f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_184 VPB N_A_1467_419#_c_1231_n 0.0070546f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1467_419#_c_1232_n 0.044898f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.615
cc_186 VPB N_A_1467_419#_c_1233_n 0.00204491f $X=-0.19 $Y=1.655 $X2=0.282
+ $Y2=1.665
cc_187 VPB N_A_1467_419#_c_1234_n 0.014134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_1467_419#_c_1228_n 0.00913838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_1467_419#_c_1236_n 0.0090738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_1247_89#_M1008_g 0.0571308f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_191 VPB N_A_1247_89#_M1023_g 0.0278503f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_192 VPB N_A_1247_89#_c_1318_n 0.018263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_1247_89#_c_1319_n 0.00346963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_1247_89#_c_1312_n 0.00930182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_1247_89#_c_1314_n 0.00113069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1247_89#_c_1315_n 0.0035373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_1832_367#_M1024_g 0.0251752f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.615
cc_198 VPB N_A_1832_367#_c_1425_n 0.00821505f $X=-0.19 $Y=1.655 $X2=0.282
+ $Y2=1.615
cc_199 VPB N_A_1832_367#_c_1420_n 0.0022917f $X=-0.19 $Y=1.655 $X2=0.282
+ $Y2=2.035
cc_200 VPB N_A_1832_367#_c_1421_n 0.00767213f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1832_367#_c_1422_n 0.00152607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1467_n 0.00446608f $X=-0.19 $Y=1.655 $X2=0.282 $Y2=2.035
cc_203 VPB N_VPWR_c_1468_n 7.46595e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1469_n 0.00525747f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1470_n 0.00832364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1471_n 0.0147008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1472_n 0.0131738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1473_n 0.03553f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1474_n 0.00419999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1475_n 0.0460827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1476_n 0.00651023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1477_n 0.0208776f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1478_n 0.00545601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1479_n 0.0167813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1480_n 0.0275062f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1481_n 0.0331879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1482_n 0.021098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1483_n 0.0169629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1466_n 0.110047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1485_n 0.00613849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1486_n 0.0044848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1487_n 0.0131092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1488_n 0.00597398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_304_533#_c_1606_n 0.00382819f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=2.12
cc_225 VPB N_A_304_533#_c_1607_n 0.00298515f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_226 VPB N_A_304_533#_c_1608_n 0.00419285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_304_533#_c_1609_n 0.00249815f $X=-0.19 $Y=1.655 $X2=0.282
+ $Y2=1.615
cc_228 VPB N_A_304_533#_c_1605_n 0.00307129f $X=-0.19 $Y=1.655 $X2=0.282
+ $Y2=2.035
cc_229 VPB N_A_304_533#_c_1611_n 0.00543994f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_304_533#_c_1612_n 0.00154182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_304_533#_c_1613_n 0.00672637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_Q_c_1684_n 0.0453583f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_233 VPB N_Q_c_1685_n 0.00723403f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_234 VPB Q 0.0103667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 N_CLK_c_237_n N_A_27_114#_c_272_n 0.0170356f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_236 N_CLK_c_238_n N_A_27_114#_c_272_n 5.92621e-19 $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_237 N_CLK_c_241_n N_A_27_114#_M1006_g 0.0170356f $X=0.385 $Y=2.12 $X2=0 $Y2=0
cc_238 N_CLK_c_236_n N_A_27_114#_c_275_n 0.0170356f $X=0.385 $Y=1.955 $X2=0
+ $Y2=0
cc_239 N_CLK_M1013_g N_A_27_114#_c_276_n 0.00919221f $X=0.475 $Y=0.78 $X2=0
+ $Y2=0
cc_240 N_CLK_M1020_g N_A_27_114#_c_310_n 0.0122586f $X=0.475 $Y=2.63 $X2=0 $Y2=0
cc_241 N_CLK_c_241_n N_A_27_114#_c_310_n 3.02199e-19 $X=0.385 $Y=2.12 $X2=0
+ $Y2=0
cc_242 N_CLK_c_238_n N_A_27_114#_c_310_n 0.00901834f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_243 N_CLK_M1013_g N_A_27_114#_c_277_n 0.0136942f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_244 N_CLK_c_238_n N_A_27_114#_c_277_n 0.0033306f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_245 N_CLK_M1013_g N_A_27_114#_c_278_n 0.00440676f $X=0.475 $Y=0.78 $X2=0
+ $Y2=0
cc_246 N_CLK_c_237_n N_A_27_114#_c_278_n 0.00139848f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_247 N_CLK_c_238_n N_A_27_114#_c_278_n 0.0297142f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_248 N_CLK_M1013_g N_A_27_114#_c_279_n 0.00446922f $X=0.475 $Y=0.78 $X2=0
+ $Y2=0
cc_249 N_CLK_c_238_n N_A_27_114#_c_279_n 0.0476093f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_250 N_CLK_c_241_n N_A_27_114#_c_311_n 0.00446922f $X=0.385 $Y=2.12 $X2=0
+ $Y2=0
cc_251 N_CLK_M1013_g N_A_27_114#_c_280_n 0.00188094f $X=0.475 $Y=0.78 $X2=0
+ $Y2=0
cc_252 N_CLK_M1020_g N_A_27_114#_c_312_n 4.46816e-19 $X=0.475 $Y=2.63 $X2=0
+ $Y2=0
cc_253 N_CLK_c_241_n N_A_27_114#_c_312_n 0.00102088f $X=0.385 $Y=2.12 $X2=0
+ $Y2=0
cc_254 N_CLK_c_238_n N_A_27_114#_c_312_n 0.0242383f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_255 N_CLK_M1013_g N_A_27_114#_c_296_n 0.0170356f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_256 N_CLK_c_237_n N_A_27_114#_c_297_n 0.00446922f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_257 N_CLK_M1013_g N_A_27_114#_c_304_n 0.007168f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_258 N_CLK_M1020_g N_VPWR_c_1467_n 0.010629f $X=0.475 $Y=2.63 $X2=0 $Y2=0
cc_259 N_CLK_M1020_g N_VPWR_c_1479_n 0.0047441f $X=0.475 $Y=2.63 $X2=0 $Y2=0
cc_260 N_CLK_M1020_g N_VPWR_c_1466_n 0.00455844f $X=0.475 $Y=2.63 $X2=0 $Y2=0
cc_261 N_CLK_M1013_g N_VGND_c_1697_n 0.00360998f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_262 N_CLK_M1013_g N_VGND_c_1703_n 0.00428973f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_263 N_CLK_M1013_g N_VGND_c_1708_n 0.00484898f $X=0.475 $Y=0.78 $X2=0 $Y2=0
cc_264 N_A_27_114#_c_284_n N_D_M1002_g 0.00429574f $X=2.515 $Y=1.26 $X2=0 $Y2=0
cc_265 N_A_27_114#_c_286_n N_D_M1002_g 0.00940627f $X=2.6 $Y=1.175 $X2=0 $Y2=0
cc_266 N_A_27_114#_c_287_n N_D_M1002_g 0.00735348f $X=3.225 $Y=0.555 $X2=0 $Y2=0
cc_267 N_A_27_114#_c_288_n N_D_M1002_g 2.7459e-19 $X=2.685 $Y=0.555 $X2=0 $Y2=0
cc_268 N_A_27_114#_c_289_n N_D_M1002_g 6.67626e-19 $X=3.31 $Y=1.44 $X2=0 $Y2=0
cc_269 N_A_27_114#_c_305_n N_D_M1002_g 0.0116914f $X=3.287 $Y=1.275 $X2=0 $Y2=0
cc_270 N_A_27_114#_M1009_g N_D_c_542_n 0.00428431f $X=3.19 $Y=2.875 $X2=0 $Y2=0
cc_271 N_A_27_114#_c_284_n N_D_c_542_n 0.0105211f $X=2.515 $Y=1.26 $X2=0 $Y2=0
cc_272 N_A_27_114#_c_290_n N_D_c_542_n 0.0116914f $X=3.31 $Y=1.44 $X2=0 $Y2=0
cc_273 N_A_27_114#_c_284_n N_D_c_543_n 0.0443491f $X=2.515 $Y=1.26 $X2=0 $Y2=0
cc_274 N_A_27_114#_M1009_g N_A_196_462#_M1015_g 0.018437f $X=3.19 $Y=2.875 $X2=0
+ $Y2=0
cc_275 N_A_27_114#_c_289_n N_A_196_462#_M1027_g 0.00498063f $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_276 N_A_27_114#_c_290_n N_A_196_462#_M1027_g 0.00103472f $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_277 N_A_27_114#_c_299_n N_A_196_462#_M1027_g 0.00400712f $X=4.47 $Y=0.587
+ $X2=0 $Y2=0
cc_278 N_A_27_114#_c_305_n N_A_196_462#_M1027_g 0.00608067f $X=3.287 $Y=1.275
+ $X2=0 $Y2=0
cc_279 N_A_27_114#_c_274_n N_A_196_462#_M1031_g 0.00620831f $X=7.01 $Y=0.555
+ $X2=0 $Y2=0
cc_280 N_A_27_114#_c_291_n N_A_196_462#_M1031_g 0.015933f $X=6.175 $Y=0.48 $X2=0
+ $Y2=0
cc_281 N_A_27_114#_c_294_n N_A_196_462#_M1031_g 0.00319828f $X=7.01 $Y=0.39
+ $X2=0 $Y2=0
cc_282 N_A_27_114#_c_302_n N_A_196_462#_M1031_g 0.0197973f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_283 N_A_27_114#_c_303_n N_A_196_462#_M1031_g 0.00952336f $X=6.26 $Y=0.48
+ $X2=0 $Y2=0
cc_284 N_A_27_114#_c_274_n N_A_196_462#_c_585_n 0.00552376f $X=7.01 $Y=0.555
+ $X2=0 $Y2=0
cc_285 N_A_27_114#_c_302_n N_A_196_462#_c_585_n 0.00835447f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_286 N_A_27_114#_c_314_n N_A_196_462#_c_586_n 5.2361e-19 $X=6.2 $Y=1.92 $X2=0
+ $Y2=0
cc_287 N_A_27_114#_c_315_n N_A_196_462#_c_586_n 0.0159935f $X=6.2 $Y=1.92 $X2=0
+ $Y2=0
cc_288 N_A_27_114#_c_302_n N_A_196_462#_c_586_n 0.00284443f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_289 N_A_27_114#_M1011_g N_A_196_462#_c_594_n 0.0148928f $X=6.295 $Y=2.665
+ $X2=0 $Y2=0
cc_290 N_A_27_114#_M1006_g N_A_196_462#_c_595_n 2.21843e-19 $X=0.905 $Y=2.63
+ $X2=0 $Y2=0
cc_291 N_A_27_114#_M1006_g N_A_196_462#_c_587_n 0.00312784f $X=0.905 $Y=2.63
+ $X2=0 $Y2=0
cc_292 N_A_27_114#_c_279_n N_A_196_462#_c_587_n 0.0379362f $X=0.895 $Y=1.54
+ $X2=0 $Y2=0
cc_293 N_A_27_114#_c_311_n N_A_196_462#_c_587_n 0.00552727f $X=0.75 $Y=2.3 $X2=0
+ $Y2=0
cc_294 N_A_27_114#_c_280_n N_A_196_462#_c_587_n 0.0204043f $X=1.04 $Y=1.1 $X2=0
+ $Y2=0
cc_295 N_A_27_114#_c_281_n N_A_196_462#_c_587_n 0.0141951f $X=1.655 $Y=0.365
+ $X2=0 $Y2=0
cc_296 N_A_27_114#_c_283_n N_A_196_462#_c_587_n 0.0416034f $X=1.74 $Y=1.175
+ $X2=0 $Y2=0
cc_297 N_A_27_114#_c_285_n N_A_196_462#_c_587_n 0.0144665f $X=1.825 $Y=1.26
+ $X2=0 $Y2=0
cc_298 N_A_27_114#_c_295_n N_A_196_462#_c_587_n 0.0144989f $X=0.995 $Y=1.265
+ $X2=0 $Y2=0
cc_299 N_A_27_114#_c_304_n N_A_196_462#_c_587_n 0.009374f $X=1.04 $Y=1.1 $X2=0
+ $Y2=0
cc_300 N_A_27_114#_M1009_g N_A_196_462#_c_597_n 2.29197e-19 $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_301 N_A_27_114#_M1009_g N_A_196_462#_c_598_n 0.0211744f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_302 N_A_27_114#_M1009_g N_A_196_462#_c_599_n 0.00146304f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_303 N_A_27_114#_c_290_n N_A_196_462#_c_599_n 7.19867e-19 $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_304 N_A_27_114#_M1009_g N_A_196_462#_c_588_n 0.00434504f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_305 N_A_27_114#_c_289_n N_A_196_462#_c_588_n 0.0137454f $X=3.31 $Y=1.44 $X2=0
+ $Y2=0
cc_306 N_A_27_114#_c_290_n N_A_196_462#_c_588_n 0.00111562f $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_307 N_A_27_114#_M1009_g N_A_196_462#_c_589_n 7.79521e-19 $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_308 N_A_27_114#_c_289_n N_A_196_462#_c_589_n 9.44736e-19 $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_309 N_A_27_114#_c_290_n N_A_196_462#_c_589_n 0.0187638f $X=3.31 $Y=1.44 $X2=0
+ $Y2=0
cc_310 N_A_27_114#_M1009_g N_A_196_462#_c_601_n 0.0017875f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_311 N_A_27_114#_c_284_n N_A_196_462#_c_601_n 0.00483077f $X=2.515 $Y=1.26
+ $X2=0 $Y2=0
cc_312 N_A_27_114#_c_285_n N_A_196_462#_c_601_n 0.00558496f $X=1.825 $Y=1.26
+ $X2=0 $Y2=0
cc_313 N_A_27_114#_c_289_n N_A_196_462#_c_601_n 0.00586127f $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_314 N_A_27_114#_c_290_n N_A_196_462#_c_601_n 0.00130725f $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_315 N_A_27_114#_M1006_g N_A_196_462#_c_602_n 5.29328e-19 $X=0.905 $Y=2.63
+ $X2=0 $Y2=0
cc_316 N_A_27_114#_c_275_n N_A_196_462#_c_602_n 0.00377308f $X=1.04 $Y=1.77
+ $X2=0 $Y2=0
cc_317 N_A_27_114#_c_311_n N_A_196_462#_c_602_n 0.00193898f $X=0.75 $Y=2.3 $X2=0
+ $Y2=0
cc_318 N_A_27_114#_c_297_n N_A_196_462#_c_602_n 0.00196952f $X=0.895 $Y=1.77
+ $X2=0 $Y2=0
cc_319 N_A_27_114#_M1011_g N_A_196_462#_c_603_n 0.00647094f $X=6.295 $Y=2.665
+ $X2=0 $Y2=0
cc_320 N_A_27_114#_c_314_n N_A_196_462#_c_603_n 0.0139799f $X=6.2 $Y=1.92 $X2=0
+ $Y2=0
cc_321 N_A_27_114#_c_315_n N_A_196_462#_c_603_n 0.0056652f $X=6.2 $Y=1.92 $X2=0
+ $Y2=0
cc_322 N_A_27_114#_c_315_n N_A_196_462#_c_605_n 0.0195126f $X=6.2 $Y=1.92 $X2=0
+ $Y2=0
cc_323 N_A_27_114#_M1006_g N_A_196_462#_c_607_n 0.00867852f $X=0.905 $Y=2.63
+ $X2=0 $Y2=0
cc_324 N_A_27_114#_c_275_n N_A_196_462#_c_607_n 0.00563771f $X=1.04 $Y=1.77
+ $X2=0 $Y2=0
cc_325 N_A_27_114#_c_310_n N_A_196_462#_c_607_n 0.00170421f $X=0.665 $Y=2.385
+ $X2=0 $Y2=0
cc_326 N_A_27_114#_c_311_n N_A_196_462#_c_607_n 0.0248176f $X=0.75 $Y=2.3 $X2=0
+ $Y2=0
cc_327 N_A_27_114#_c_297_n N_A_196_462#_c_607_n 0.00740586f $X=0.895 $Y=1.77
+ $X2=0 $Y2=0
cc_328 N_A_27_114#_c_291_n N_A_695_375#_M1028_d 0.00756935f $X=6.175 $Y=0.48
+ $X2=-0.19 $Y2=-0.245
cc_329 N_A_27_114#_c_292_n N_A_695_375#_M1028_d 0.00215999f $X=5.73 $Y=0.48
+ $X2=-0.19 $Y2=-0.245
cc_330 N_A_27_114#_M1009_g N_A_695_375#_c_791_n 0.0830148f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_331 N_A_27_114#_c_299_n N_A_695_375#_M1018_g 0.0045995f $X=4.47 $Y=0.587
+ $X2=0 $Y2=0
cc_332 N_A_27_114#_c_300_n N_A_695_375#_M1018_g 0.00201117f $X=4.835 $Y=0.587
+ $X2=0 $Y2=0
cc_333 N_A_27_114#_c_302_n N_A_695_375#_c_784_n 0.0245837f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_334 N_A_27_114#_M1011_g N_A_695_375#_c_794_n 0.00146327f $X=6.295 $Y=2.665
+ $X2=0 $Y2=0
cc_335 N_A_27_114#_c_314_n N_A_695_375#_c_794_n 0.0235435f $X=6.2 $Y=1.92 $X2=0
+ $Y2=0
cc_336 N_A_27_114#_c_315_n N_A_695_375#_c_794_n 0.00285789f $X=6.2 $Y=1.92 $X2=0
+ $Y2=0
cc_337 N_A_27_114#_c_302_n N_A_695_375#_c_794_n 0.005269f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_338 N_A_27_114#_c_292_n N_A_695_375#_c_787_n 0.0280606f $X=5.73 $Y=0.48 $X2=0
+ $Y2=0
cc_339 N_A_27_114#_c_302_n N_A_695_375#_c_787_n 0.013453f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_340 N_A_27_114#_c_302_n N_A_695_375#_c_788_n 0.0111958f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_341 N_A_27_114#_c_314_n N_A_695_375#_c_809_n 0.00451428f $X=6.2 $Y=1.92 $X2=0
+ $Y2=0
cc_342 N_A_27_114#_c_315_n N_A_695_375#_c_809_n 0.00287452f $X=6.2 $Y=1.92 $X2=0
+ $Y2=0
cc_343 N_A_27_114#_c_280_n N_RESET_B_M1007_g 2.26442e-19 $X=1.04 $Y=1.1 $X2=0
+ $Y2=0
cc_344 N_A_27_114#_c_281_n N_RESET_B_M1007_g 0.00258609f $X=1.655 $Y=0.365 $X2=0
+ $Y2=0
cc_345 N_A_27_114#_c_283_n N_RESET_B_M1007_g 0.0180822f $X=1.74 $Y=1.175 $X2=0
+ $Y2=0
cc_346 N_A_27_114#_c_284_n N_RESET_B_M1007_g 0.0143341f $X=2.515 $Y=1.26 $X2=0
+ $Y2=0
cc_347 N_A_27_114#_c_285_n N_RESET_B_M1007_g 0.00375834f $X=1.825 $Y=1.26 $X2=0
+ $Y2=0
cc_348 N_A_27_114#_c_304_n N_RESET_B_M1007_g 0.0177651f $X=1.04 $Y=1.1 $X2=0
+ $Y2=0
cc_349 N_A_27_114#_c_281_n N_RESET_B_c_890_n 0.00443325f $X=1.655 $Y=0.365 $X2=0
+ $Y2=0
cc_350 N_A_27_114#_c_283_n N_RESET_B_M1010_g 8.52563e-19 $X=1.74 $Y=1.175 $X2=0
+ $Y2=0
cc_351 N_A_27_114#_c_284_n N_RESET_B_M1010_g 0.0108072f $X=2.515 $Y=1.26 $X2=0
+ $Y2=0
cc_352 N_A_27_114#_c_286_n N_RESET_B_M1010_g 0.00219874f $X=2.6 $Y=1.175 $X2=0
+ $Y2=0
cc_353 N_A_27_114#_c_288_n N_RESET_B_M1010_g 0.00355358f $X=2.685 $Y=0.555 $X2=0
+ $Y2=0
cc_354 N_A_27_114#_c_287_n N_RESET_B_c_892_n 0.00884495f $X=3.225 $Y=0.555 $X2=0
+ $Y2=0
cc_355 N_A_27_114#_c_288_n N_RESET_B_c_892_n 0.00324383f $X=2.685 $Y=0.555 $X2=0
+ $Y2=0
cc_356 N_A_27_114#_c_292_n N_RESET_B_c_892_n 8.57535e-19 $X=5.73 $Y=0.48 $X2=0
+ $Y2=0
cc_357 N_A_27_114#_c_298_n N_RESET_B_c_892_n 0.00399336f $X=3.31 $Y=0.555 $X2=0
+ $Y2=0
cc_358 N_A_27_114#_c_299_n N_RESET_B_c_892_n 0.0257939f $X=4.47 $Y=0.587 $X2=0
+ $Y2=0
cc_359 N_A_27_114#_c_305_n N_RESET_B_c_892_n 0.0074428f $X=3.287 $Y=1.275 $X2=0
+ $Y2=0
cc_360 N_A_27_114#_c_300_n N_RESET_B_M1014_g 0.00934553f $X=4.835 $Y=0.587 $X2=0
+ $Y2=0
cc_361 N_A_27_114#_c_301_n N_RESET_B_M1014_g 0.00714923f $X=5.505 $Y=0.48 $X2=0
+ $Y2=0
cc_362 N_A_27_114#_M1011_g N_RESET_B_c_907_n 0.014834f $X=6.295 $Y=2.665 $X2=0
+ $Y2=0
cc_363 N_A_27_114#_M1011_g N_RESET_B_c_933_n 0.00416455f $X=6.295 $Y=2.665 $X2=0
+ $Y2=0
cc_364 N_A_27_114#_c_289_n N_A_559_533#_M1004_d 0.0044492f $X=3.31 $Y=1.44
+ $X2=-0.19 $Y2=-0.245
cc_365 N_A_27_114#_c_292_n N_A_559_533#_c_1075_n 0.0191618f $X=5.73 $Y=0.48
+ $X2=0 $Y2=0
cc_366 N_A_27_114#_c_301_n N_A_559_533#_c_1075_n 0.00776506f $X=5.505 $Y=0.48
+ $X2=0 $Y2=0
cc_367 N_A_27_114#_c_302_n N_A_559_533#_c_1075_n 9.00297e-19 $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_368 N_A_27_114#_M1011_g N_A_559_533#_c_1080_n 0.0272237f $X=6.295 $Y=2.665
+ $X2=0 $Y2=0
cc_369 N_A_27_114#_c_315_n N_A_559_533#_c_1080_n 0.00942378f $X=6.2 $Y=1.92
+ $X2=0 $Y2=0
cc_370 N_A_27_114#_M1009_g N_A_559_533#_c_1099_n 0.00919f $X=3.19 $Y=2.875 $X2=0
+ $Y2=0
cc_371 N_A_27_114#_M1009_g N_A_559_533#_c_1082_n 0.00374419f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_372 N_A_27_114#_c_289_n N_A_559_533#_c_1101_n 0.0265609f $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_373 N_A_27_114#_c_299_n N_A_559_533#_c_1101_n 0.0384846f $X=4.47 $Y=0.587
+ $X2=0 $Y2=0
cc_374 N_A_27_114#_c_305_n N_A_559_533#_c_1101_n 0.00112264f $X=3.287 $Y=1.275
+ $X2=0 $Y2=0
cc_375 N_A_27_114#_M1009_g N_A_559_533#_c_1084_n 9.93271e-19 $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_376 N_A_27_114#_c_299_n N_A_559_533#_c_1076_n 0.0127847f $X=4.47 $Y=0.587
+ $X2=0 $Y2=0
cc_377 N_A_27_114#_c_300_n N_A_559_533#_c_1076_n 0.0340728f $X=4.835 $Y=0.587
+ $X2=0 $Y2=0
cc_378 N_A_27_114#_c_301_n N_A_559_533#_c_1077_n 0.0168728f $X=5.505 $Y=0.48
+ $X2=0 $Y2=0
cc_379 N_A_27_114#_c_315_n N_A_559_533#_c_1091_n 0.00266077f $X=6.2 $Y=1.92
+ $X2=0 $Y2=0
cc_380 N_A_27_114#_c_301_n N_A_559_533#_c_1078_n 0.001215f $X=5.505 $Y=0.48
+ $X2=0 $Y2=0
cc_381 N_A_27_114#_c_274_n N_A_1467_419#_M1000_g 0.0270687f $X=7.01 $Y=0.555
+ $X2=0 $Y2=0
cc_382 N_A_27_114#_c_294_n N_A_1467_419#_M1000_g 0.00129738f $X=7.01 $Y=0.39
+ $X2=0 $Y2=0
cc_383 N_A_27_114#_c_293_n N_A_1247_89#_M1031_d 0.0103142f $X=7.01 $Y=0.39
+ $X2=-0.19 $Y2=-0.245
cc_384 N_A_27_114#_c_302_n N_A_1247_89#_M1031_d 0.00368341f $X=6.225 $Y=1.755
+ $X2=-0.19 $Y2=-0.245
cc_385 N_A_27_114#_c_303_n N_A_1247_89#_M1031_d 0.00339727f $X=6.26 $Y=0.48
+ $X2=-0.19 $Y2=-0.245
cc_386 N_A_27_114#_c_274_n N_A_1247_89#_c_1310_n 0.0132881f $X=7.01 $Y=0.555
+ $X2=0 $Y2=0
cc_387 N_A_27_114#_c_293_n N_A_1247_89#_c_1310_n 0.020747f $X=7.01 $Y=0.39 $X2=0
+ $Y2=0
cc_388 N_A_27_114#_c_302_n N_A_1247_89#_c_1310_n 0.0369888f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_389 N_A_27_114#_c_303_n N_A_1247_89#_c_1310_n 8.37543e-19 $X=6.26 $Y=0.48
+ $X2=0 $Y2=0
cc_390 N_A_27_114#_c_274_n N_A_1247_89#_c_1311_n 0.00646191f $X=7.01 $Y=0.555
+ $X2=0 $Y2=0
cc_391 N_A_27_114#_c_293_n N_A_1247_89#_c_1311_n 0.0101095f $X=7.01 $Y=0.39
+ $X2=0 $Y2=0
cc_392 N_A_27_114#_c_294_n N_A_1247_89#_c_1311_n 0.0028231f $X=7.01 $Y=0.39
+ $X2=0 $Y2=0
cc_393 N_A_27_114#_c_315_n N_A_1247_89#_c_1312_n 0.00431327f $X=6.2 $Y=1.92
+ $X2=0 $Y2=0
cc_394 N_A_27_114#_c_302_n N_A_1247_89#_c_1312_n 0.0517836f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_395 N_A_27_114#_c_302_n N_A_1247_89#_c_1313_n 0.0143568f $X=6.225 $Y=1.755
+ $X2=0 $Y2=0
cc_396 N_A_27_114#_c_310_n N_VPWR_M1020_d 0.00177916f $X=0.665 $Y=2.385
+ $X2=-0.19 $Y2=-0.245
cc_397 N_A_27_114#_M1006_g N_VPWR_c_1467_n 0.00996799f $X=0.905 $Y=2.63 $X2=0
+ $Y2=0
cc_398 N_A_27_114#_c_310_n N_VPWR_c_1467_n 0.0162291f $X=0.665 $Y=2.385 $X2=0
+ $Y2=0
cc_399 N_A_27_114#_c_312_n N_VPWR_c_1467_n 0.0131449f $X=0.26 $Y=2.465 $X2=0
+ $Y2=0
cc_400 N_A_27_114#_M1009_g N_VPWR_c_1473_n 0.00351226f $X=3.19 $Y=2.875 $X2=0
+ $Y2=0
cc_401 N_A_27_114#_M1011_g N_VPWR_c_1475_n 0.00351226f $X=6.295 $Y=2.665 $X2=0
+ $Y2=0
cc_402 N_A_27_114#_c_312_n N_VPWR_c_1479_n 0.0110559f $X=0.26 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A_27_114#_M1006_g N_VPWR_c_1480_n 0.0047441f $X=0.905 $Y=2.63 $X2=0
+ $Y2=0
cc_404 N_A_27_114#_M1006_g N_VPWR_c_1466_n 0.00455844f $X=0.905 $Y=2.63 $X2=0
+ $Y2=0
cc_405 N_A_27_114#_M1009_g N_VPWR_c_1466_n 0.00526607f $X=3.19 $Y=2.875 $X2=0
+ $Y2=0
cc_406 N_A_27_114#_M1011_g N_VPWR_c_1466_n 0.00648053f $X=6.295 $Y=2.665 $X2=0
+ $Y2=0
cc_407 N_A_27_114#_c_310_n N_VPWR_c_1466_n 0.00636496f $X=0.665 $Y=2.385 $X2=0
+ $Y2=0
cc_408 N_A_27_114#_c_312_n N_VPWR_c_1466_n 0.00946638f $X=0.26 $Y=2.465 $X2=0
+ $Y2=0
cc_409 N_A_27_114#_M1006_g N_A_304_533#_c_1606_n 0.00163718f $X=0.905 $Y=2.63
+ $X2=0 $Y2=0
cc_410 N_A_27_114#_M1009_g N_A_304_533#_c_1609_n 0.00696411f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_411 N_A_27_114#_M1009_g N_A_304_533#_c_1605_n 0.00275155f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_412 N_A_27_114#_c_284_n N_A_304_533#_c_1605_n 0.0137445f $X=2.515 $Y=1.26
+ $X2=0 $Y2=0
cc_413 N_A_27_114#_c_286_n N_A_304_533#_c_1605_n 0.0126831f $X=2.6 $Y=1.175
+ $X2=0 $Y2=0
cc_414 N_A_27_114#_c_287_n N_A_304_533#_c_1605_n 0.0145268f $X=3.225 $Y=0.555
+ $X2=0 $Y2=0
cc_415 N_A_27_114#_c_289_n N_A_304_533#_c_1605_n 0.0438387f $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_416 N_A_27_114#_c_305_n N_A_304_533#_c_1605_n 0.00350959f $X=3.287 $Y=1.275
+ $X2=0 $Y2=0
cc_417 N_A_27_114#_M1009_g N_A_304_533#_c_1611_n 0.0144474f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_418 N_A_27_114#_M1009_g N_A_304_533#_c_1613_n 0.012202f $X=3.19 $Y=2.875
+ $X2=0 $Y2=0
cc_419 N_A_27_114#_c_289_n N_A_304_533#_c_1613_n 0.00128451f $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_420 N_A_27_114#_c_290_n N_A_304_533#_c_1613_n 6.15908e-19 $X=3.31 $Y=1.44
+ $X2=0 $Y2=0
cc_421 N_A_27_114#_c_280_n N_VGND_M1013_d 0.00413533f $X=1.04 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_422 N_A_27_114#_c_301_n N_VGND_M1014_d 0.00940607f $X=5.505 $Y=0.48 $X2=0
+ $Y2=0
cc_423 N_A_27_114#_c_277_n N_VGND_c_1697_n 0.00519653f $X=0.665 $Y=1.19 $X2=0
+ $Y2=0
cc_424 N_A_27_114#_c_280_n N_VGND_c_1697_n 0.0354425f $X=1.04 $Y=1.1 $X2=0 $Y2=0
cc_425 N_A_27_114#_c_282_n N_VGND_c_1697_n 0.0144678f $X=1.125 $Y=0.365 $X2=0
+ $Y2=0
cc_426 N_A_27_114#_c_295_n N_VGND_c_1697_n 0.0109396f $X=0.995 $Y=1.265 $X2=0
+ $Y2=0
cc_427 N_A_27_114#_c_304_n N_VGND_c_1697_n 0.00135451f $X=1.04 $Y=1.1 $X2=0
+ $Y2=0
cc_428 N_A_27_114#_c_281_n N_VGND_c_1698_n 0.0132272f $X=1.655 $Y=0.365 $X2=0
+ $Y2=0
cc_429 N_A_27_114#_c_283_n N_VGND_c_1698_n 0.040112f $X=1.74 $Y=1.175 $X2=0
+ $Y2=0
cc_430 N_A_27_114#_c_284_n N_VGND_c_1698_n 0.0244345f $X=2.515 $Y=1.26 $X2=0
+ $Y2=0
cc_431 N_A_27_114#_c_286_n N_VGND_c_1698_n 0.016804f $X=2.6 $Y=1.175 $X2=0 $Y2=0
cc_432 N_A_27_114#_c_288_n N_VGND_c_1698_n 0.0137302f $X=2.685 $Y=0.555 $X2=0
+ $Y2=0
cc_433 N_A_27_114#_c_274_n N_VGND_c_1699_n 0.00227001f $X=7.01 $Y=0.555 $X2=0
+ $Y2=0
cc_434 N_A_27_114#_c_293_n N_VGND_c_1699_n 0.0135276f $X=7.01 $Y=0.39 $X2=0
+ $Y2=0
cc_435 N_A_27_114#_c_294_n N_VGND_c_1699_n 0.00306163f $X=7.01 $Y=0.39 $X2=0
+ $Y2=0
cc_436 N_A_27_114#_c_292_n N_VGND_c_1701_n 0.0459634f $X=5.73 $Y=0.48 $X2=0
+ $Y2=0
cc_437 N_A_27_114#_c_293_n N_VGND_c_1701_n 0.0541731f $X=7.01 $Y=0.39 $X2=0
+ $Y2=0
cc_438 N_A_27_114#_c_294_n N_VGND_c_1701_n 0.00601136f $X=7.01 $Y=0.39 $X2=0
+ $Y2=0
cc_439 N_A_27_114#_c_301_n N_VGND_c_1701_n 0.00321687f $X=5.505 $Y=0.48 $X2=0
+ $Y2=0
cc_440 N_A_27_114#_c_303_n N_VGND_c_1701_n 0.0121867f $X=6.26 $Y=0.48 $X2=0
+ $Y2=0
cc_441 N_A_27_114#_c_276_n N_VGND_c_1703_n 0.00596511f $X=0.26 $Y=0.785 $X2=0
+ $Y2=0
cc_442 N_A_27_114#_c_281_n N_VGND_c_1704_n 0.0398657f $X=1.655 $Y=0.365 $X2=0
+ $Y2=0
cc_443 N_A_27_114#_c_282_n N_VGND_c_1704_n 0.0105206f $X=1.125 $Y=0.365 $X2=0
+ $Y2=0
cc_444 N_A_27_114#_c_304_n N_VGND_c_1704_n 6.40413e-19 $X=1.04 $Y=1.1 $X2=0
+ $Y2=0
cc_445 N_A_27_114#_c_287_n N_VGND_c_1705_n 0.0146104f $X=3.225 $Y=0.555 $X2=0
+ $Y2=0
cc_446 N_A_27_114#_c_288_n N_VGND_c_1705_n 0.00508759f $X=2.685 $Y=0.555 $X2=0
+ $Y2=0
cc_447 N_A_27_114#_c_298_n N_VGND_c_1705_n 0.00508515f $X=3.31 $Y=0.555 $X2=0
+ $Y2=0
cc_448 N_A_27_114#_c_299_n N_VGND_c_1705_n 0.0390696f $X=4.47 $Y=0.587 $X2=0
+ $Y2=0
cc_449 N_A_27_114#_c_301_n N_VGND_c_1705_n 0.00383594f $X=5.505 $Y=0.48 $X2=0
+ $Y2=0
cc_450 N_A_27_114#_c_276_n N_VGND_c_1708_n 0.0100079f $X=0.26 $Y=0.785 $X2=0
+ $Y2=0
cc_451 N_A_27_114#_c_281_n N_VGND_c_1708_n 0.0259601f $X=1.655 $Y=0.365 $X2=0
+ $Y2=0
cc_452 N_A_27_114#_c_282_n N_VGND_c_1708_n 0.00652894f $X=1.125 $Y=0.365 $X2=0
+ $Y2=0
cc_453 N_A_27_114#_c_287_n N_VGND_c_1708_n 0.0153373f $X=3.225 $Y=0.555 $X2=0
+ $Y2=0
cc_454 N_A_27_114#_c_288_n N_VGND_c_1708_n 0.00512732f $X=2.685 $Y=0.555 $X2=0
+ $Y2=0
cc_455 N_A_27_114#_c_292_n N_VGND_c_1708_n 0.0254292f $X=5.73 $Y=0.48 $X2=0
+ $Y2=0
cc_456 N_A_27_114#_c_293_n N_VGND_c_1708_n 0.0300145f $X=7.01 $Y=0.39 $X2=0
+ $Y2=0
cc_457 N_A_27_114#_c_294_n N_VGND_c_1708_n 0.00828645f $X=7.01 $Y=0.39 $X2=0
+ $Y2=0
cc_458 N_A_27_114#_c_298_n N_VGND_c_1708_n 0.00512732f $X=3.31 $Y=0.555 $X2=0
+ $Y2=0
cc_459 N_A_27_114#_c_299_n N_VGND_c_1708_n 0.0409596f $X=4.47 $Y=0.587 $X2=0
+ $Y2=0
cc_460 N_A_27_114#_c_301_n N_VGND_c_1708_n 0.0117232f $X=5.505 $Y=0.48 $X2=0
+ $Y2=0
cc_461 N_A_27_114#_c_303_n N_VGND_c_1708_n 0.00660921f $X=6.26 $Y=0.48 $X2=0
+ $Y2=0
cc_462 N_A_27_114#_c_292_n N_VGND_c_1711_n 0.00824664f $X=5.73 $Y=0.48 $X2=0
+ $Y2=0
cc_463 N_A_27_114#_c_301_n N_VGND_c_1711_n 0.0241876f $X=5.505 $Y=0.48 $X2=0
+ $Y2=0
cc_464 N_A_27_114#_c_300_n A_875_149# 0.0025911f $X=4.835 $Y=0.587 $X2=-0.19
+ $Y2=-0.245
cc_465 N_D_M1021_g N_A_196_462#_M1015_g 0.0201301f $X=2.29 $Y=2.875 $X2=0 $Y2=0
cc_466 N_D_c_543_n N_A_196_462#_c_587_n 0.0130063f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_467 N_D_M1021_g N_A_196_462#_c_597_n 0.0115205f $X=2.29 $Y=2.875 $X2=0 $Y2=0
cc_468 N_D_c_542_n N_A_196_462#_c_597_n 0.00332609f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_469 N_D_c_543_n N_A_196_462#_c_597_n 0.0178266f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_470 N_D_M1021_g N_A_196_462#_c_598_n 0.0220509f $X=2.29 $Y=2.875 $X2=0 $Y2=0
cc_471 N_D_c_542_n N_A_196_462#_c_598_n 0.00745362f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_472 N_D_M1021_g N_A_196_462#_c_601_n 0.00612539f $X=2.29 $Y=2.875 $X2=0 $Y2=0
cc_473 N_D_c_542_n N_A_196_462#_c_601_n 0.0037916f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_474 N_D_c_543_n N_A_196_462#_c_601_n 0.016162f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_475 N_D_c_542_n N_RESET_B_M1007_g 0.0634747f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_476 N_D_c_543_n N_RESET_B_M1007_g 0.00448711f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_477 N_D_M1002_g N_RESET_B_M1010_g 0.0402981f $X=2.745 $Y=0.955 $X2=0 $Y2=0
cc_478 N_D_c_542_n N_RESET_B_M1010_g 0.00960888f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_479 N_D_M1002_g N_RESET_B_c_892_n 0.00744285f $X=2.745 $Y=0.955 $X2=0 $Y2=0
cc_480 N_D_M1021_g N_VPWR_c_1468_n 0.00789591f $X=2.29 $Y=2.875 $X2=0 $Y2=0
cc_481 N_D_M1021_g N_VPWR_c_1473_n 0.00348975f $X=2.29 $Y=2.875 $X2=0 $Y2=0
cc_482 N_D_M1021_g N_VPWR_c_1466_n 0.00420719f $X=2.29 $Y=2.875 $X2=0 $Y2=0
cc_483 N_D_M1021_g N_A_304_533#_c_1607_n 0.0115676f $X=2.29 $Y=2.875 $X2=0 $Y2=0
cc_484 N_D_M1002_g N_A_304_533#_c_1605_n 0.00722174f $X=2.745 $Y=0.955 $X2=0
+ $Y2=0
cc_485 N_D_c_542_n N_A_304_533#_c_1605_n 5.30613e-19 $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_486 N_D_c_543_n N_A_304_533#_c_1605_n 0.0136643f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_487 N_D_M1021_g N_A_304_533#_c_1613_n 0.00311905f $X=2.29 $Y=2.875 $X2=0
+ $Y2=0
cc_488 N_D_c_542_n N_A_304_533#_c_1613_n 2.24569e-19 $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_489 N_D_c_543_n N_A_304_533#_c_1613_n 0.0028641f $X=2.38 $Y=1.67 $X2=0 $Y2=0
cc_490 N_D_M1002_g N_VGND_c_1698_n 3.08645e-19 $X=2.745 $Y=0.955 $X2=0 $Y2=0
cc_491 N_A_196_462#_c_599_n N_A_695_375#_M1029_g 0.00837493f $X=3.85 $Y=1.875
+ $X2=0 $Y2=0
cc_492 N_A_196_462#_c_599_n N_A_695_375#_c_790_n 0.0195026f $X=3.85 $Y=1.875
+ $X2=0 $Y2=0
cc_493 N_A_196_462#_c_588_n N_A_695_375#_c_790_n 0.00136392f $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_494 N_A_196_462#_c_589_n N_A_695_375#_c_790_n 0.0181259f $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_495 N_A_196_462#_c_603_n N_A_695_375#_c_790_n 0.0126894f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_496 N_A_196_462#_c_599_n N_A_695_375#_c_791_n 0.00822711f $X=3.85 $Y=1.875
+ $X2=0 $Y2=0
cc_497 N_A_196_462#_M1027_g N_A_695_375#_M1018_g 0.0321064f $X=3.94 $Y=0.955
+ $X2=0 $Y2=0
cc_498 N_A_196_462#_c_588_n N_A_695_375#_M1018_g 0.00127f $X=3.85 $Y=1.47 $X2=0
+ $Y2=0
cc_499 N_A_196_462#_c_588_n N_A_695_375#_c_782_n 0.00531873f $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_500 N_A_196_462#_c_603_n N_A_695_375#_c_783_n 0.0228092f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_501 N_A_196_462#_M1031_g N_A_695_375#_c_784_n 0.00586816f $X=6.16 $Y=0.765
+ $X2=0 $Y2=0
cc_502 N_A_196_462#_c_603_n N_A_695_375#_c_794_n 0.0171347f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_503 N_A_196_462#_c_599_n N_A_695_375#_c_785_n 0.00510245f $X=3.85 $Y=1.875
+ $X2=0 $Y2=0
cc_504 N_A_196_462#_c_588_n N_A_695_375#_c_785_n 0.0338985f $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_505 N_A_196_462#_c_589_n N_A_695_375#_c_785_n 9.74578e-19 $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_506 N_A_196_462#_c_603_n N_A_695_375#_c_785_n 0.00888897f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_507 N_A_196_462#_c_589_n N_A_695_375#_c_786_n 0.0321064f $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_508 N_A_196_462#_M1031_g N_A_695_375#_c_787_n 0.00183779f $X=6.16 $Y=0.765
+ $X2=0 $Y2=0
cc_509 N_A_196_462#_c_586_n N_A_695_375#_c_788_n 5.68329e-19 $X=6.235 $Y=1.44
+ $X2=0 $Y2=0
cc_510 N_A_196_462#_c_603_n N_A_695_375#_c_788_n 0.00425903f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_511 N_A_196_462#_c_603_n N_A_695_375#_c_809_n 0.0112806f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_512 N_A_196_462#_c_595_n N_RESET_B_M1007_g 0.00542593f $X=1.12 $Y=2.455 $X2=0
+ $Y2=0
cc_513 N_A_196_462#_c_587_n N_RESET_B_M1007_g 0.0121503f $X=1.39 $Y=0.785 $X2=0
+ $Y2=0
cc_514 N_A_196_462#_c_597_n N_RESET_B_M1007_g 0.0141308f $X=2.74 $Y=2.24 $X2=0
+ $Y2=0
cc_515 N_A_196_462#_c_601_n N_RESET_B_M1007_g 0.0104207f $X=3.455 $Y=2.035 $X2=0
+ $Y2=0
cc_516 N_A_196_462#_c_607_n N_RESET_B_M1007_g 0.00504473f $X=1.485 $Y=2.137
+ $X2=0 $Y2=0
cc_517 N_A_196_462#_M1027_g N_RESET_B_c_892_n 0.00743797f $X=3.94 $Y=0.955 $X2=0
+ $Y2=0
cc_518 N_A_196_462#_c_603_n N_RESET_B_c_902_n 0.00242864f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_519 N_A_196_462#_c_603_n N_RESET_B_M1014_g 0.0061786f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_520 N_A_196_462#_c_603_n N_RESET_B_c_906_n 0.0108664f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_521 N_A_196_462#_M1005_g N_RESET_B_c_907_n 0.01515f $X=6.82 $Y=2.795 $X2=0
+ $Y2=0
cc_522 N_A_196_462#_c_594_n N_RESET_B_c_907_n 0.00300807f $X=6.935 $Y=2.215
+ $X2=0 $Y2=0
cc_523 N_A_196_462#_c_585_n N_RESET_B_c_896_n 0.00267841f $X=6.575 $Y=1.44 $X2=0
+ $Y2=0
cc_524 N_A_196_462#_c_590_n N_RESET_B_c_896_n 0.0267823f $X=6.96 $Y=1.71 $X2=0
+ $Y2=0
cc_525 N_A_196_462#_M1005_g N_RESET_B_c_909_n 0.00731848f $X=6.82 $Y=2.795 $X2=0
+ $Y2=0
cc_526 N_A_196_462#_c_707_p N_RESET_B_c_909_n 0.00669343f $X=6.96 $Y=2.035 $X2=0
+ $Y2=0
cc_527 N_A_196_462#_c_605_n N_RESET_B_c_909_n 0.00219977f $X=6.96 $Y=1.71 $X2=0
+ $Y2=0
cc_528 N_A_196_462#_c_590_n N_RESET_B_c_909_n 0.0215141f $X=6.96 $Y=1.71 $X2=0
+ $Y2=0
cc_529 N_A_196_462#_M1031_g N_A_559_533#_c_1075_n 0.0095923f $X=6.16 $Y=0.765
+ $X2=0 $Y2=0
cc_530 N_A_196_462#_c_603_n N_A_559_533#_c_1080_n 0.0044583f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_531 N_A_196_462#_c_603_n N_A_559_533#_M1012_g 0.00138046f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_532 N_A_196_462#_M1027_g N_A_559_533#_c_1101_n 0.00657099f $X=3.94 $Y=0.955
+ $X2=0 $Y2=0
cc_533 N_A_196_462#_c_588_n N_A_559_533#_c_1101_n 0.0238888f $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_534 N_A_196_462#_c_589_n N_A_559_533#_c_1101_n 0.00399404f $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_535 N_A_196_462#_c_599_n N_A_559_533#_c_1083_n 0.0213733f $X=3.85 $Y=1.875
+ $X2=0 $Y2=0
cc_536 N_A_196_462#_c_603_n N_A_559_533#_c_1083_n 0.00619918f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_537 N_A_196_462#_c_604_n N_A_559_533#_c_1083_n 0.00105234f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_538 N_A_196_462#_c_599_n N_A_559_533#_c_1084_n 0.00627087f $X=3.85 $Y=1.875
+ $X2=0 $Y2=0
cc_539 N_A_196_462#_c_601_n N_A_559_533#_c_1084_n 0.00174943f $X=3.455 $Y=2.035
+ $X2=0 $Y2=0
cc_540 N_A_196_462#_c_604_n N_A_559_533#_c_1084_n 9.34656e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_541 N_A_196_462#_c_603_n N_A_559_533#_c_1087_n 0.0246756f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_542 N_A_196_462#_c_599_n N_A_559_533#_c_1088_n 0.00468108f $X=3.85 $Y=1.875
+ $X2=0 $Y2=0
cc_543 N_A_196_462#_c_603_n N_A_559_533#_c_1088_n 0.00780264f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_544 N_A_196_462#_M1027_g N_A_559_533#_c_1125_n 0.00450683f $X=3.94 $Y=0.955
+ $X2=0 $Y2=0
cc_545 N_A_196_462#_c_603_n N_A_559_533#_c_1089_n 0.00197326f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_546 N_A_196_462#_c_603_n N_A_559_533#_c_1090_n 0.0208625f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_547 N_A_196_462#_c_603_n N_A_559_533#_c_1091_n 7.31737e-19 $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_548 N_A_196_462#_c_586_n N_A_559_533#_c_1078_n 0.0095923f $X=6.235 $Y=1.44
+ $X2=0 $Y2=0
cc_549 N_A_196_462#_c_585_n N_A_1467_419#_M1000_g 0.0299111f $X=6.575 $Y=1.44
+ $X2=0 $Y2=0
cc_550 N_A_196_462#_c_590_n N_A_1467_419#_M1000_g 6.00385e-19 $X=6.96 $Y=1.71
+ $X2=0 $Y2=0
cc_551 N_A_196_462#_M1005_g N_A_1467_419#_c_1232_n 0.0211083f $X=6.82 $Y=2.795
+ $X2=0 $Y2=0
cc_552 N_A_196_462#_c_594_n N_A_1467_419#_c_1232_n 0.00752726f $X=6.935 $Y=2.215
+ $X2=0 $Y2=0
cc_553 N_A_196_462#_M1031_g N_A_1247_89#_c_1310_n 0.00169042f $X=6.16 $Y=0.765
+ $X2=0 $Y2=0
cc_554 N_A_196_462#_c_585_n N_A_1247_89#_c_1311_n 0.00691077f $X=6.575 $Y=1.44
+ $X2=0 $Y2=0
cc_555 N_A_196_462#_c_603_n N_A_1247_89#_c_1311_n 0.00105285f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_556 N_A_196_462#_c_707_p N_A_1247_89#_c_1311_n 0.0036902f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_557 N_A_196_462#_c_590_n N_A_1247_89#_c_1311_n 0.0139133f $X=6.96 $Y=1.71
+ $X2=0 $Y2=0
cc_558 N_A_196_462#_c_594_n N_A_1247_89#_c_1319_n 0.00585487f $X=6.935 $Y=2.215
+ $X2=0 $Y2=0
cc_559 N_A_196_462#_c_603_n N_A_1247_89#_c_1319_n 0.00735778f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_560 N_A_196_462#_c_585_n N_A_1247_89#_c_1312_n 0.0189138f $X=6.575 $Y=1.44
+ $X2=0 $Y2=0
cc_561 N_A_196_462#_c_603_n N_A_1247_89#_c_1312_n 0.0202337f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_562 N_A_196_462#_c_707_p N_A_1247_89#_c_1312_n 0.00237532f $X=6.96 $Y=2.035
+ $X2=0 $Y2=0
cc_563 N_A_196_462#_c_605_n N_A_1247_89#_c_1312_n 0.00585487f $X=6.96 $Y=1.71
+ $X2=0 $Y2=0
cc_564 N_A_196_462#_c_590_n N_A_1247_89#_c_1312_n 0.0463998f $X=6.96 $Y=1.71
+ $X2=0 $Y2=0
cc_565 N_A_196_462#_M1031_g N_A_1247_89#_c_1313_n 9.88984e-19 $X=6.16 $Y=0.765
+ $X2=0 $Y2=0
cc_566 N_A_196_462#_c_585_n N_A_1247_89#_c_1313_n 0.00792363f $X=6.575 $Y=1.44
+ $X2=0 $Y2=0
cc_567 N_A_196_462#_c_603_n N_A_1247_89#_c_1313_n 0.00259098f $X=6.815 $Y=2.035
+ $X2=0 $Y2=0
cc_568 N_A_196_462#_c_595_n N_VPWR_c_1467_n 0.0123683f $X=1.12 $Y=2.455 $X2=0
+ $Y2=0
cc_569 N_A_196_462#_M1015_g N_VPWR_c_1468_n 0.00116179f $X=2.72 $Y=2.875 $X2=0
+ $Y2=0
cc_570 N_A_196_462#_M1015_g N_VPWR_c_1473_n 0.00419621f $X=2.72 $Y=2.875 $X2=0
+ $Y2=0
cc_571 N_A_196_462#_M1005_g N_VPWR_c_1475_n 0.00302501f $X=6.82 $Y=2.795 $X2=0
+ $Y2=0
cc_572 N_A_196_462#_c_595_n N_VPWR_c_1480_n 0.0105907f $X=1.12 $Y=2.455 $X2=0
+ $Y2=0
cc_573 N_A_196_462#_M1015_g N_VPWR_c_1466_n 0.00609424f $X=2.72 $Y=2.875 $X2=0
+ $Y2=0
cc_574 N_A_196_462#_M1005_g N_VPWR_c_1466_n 0.00457741f $X=6.82 $Y=2.795 $X2=0
+ $Y2=0
cc_575 N_A_196_462#_c_595_n N_VPWR_c_1466_n 0.00938517f $X=1.12 $Y=2.455 $X2=0
+ $Y2=0
cc_576 N_A_196_462#_c_595_n N_A_304_533#_c_1606_n 0.02075f $X=1.12 $Y=2.455
+ $X2=0 $Y2=0
cc_577 N_A_196_462#_c_597_n N_A_304_533#_c_1607_n 0.0463162f $X=2.74 $Y=2.24
+ $X2=0 $Y2=0
cc_578 N_A_196_462#_c_595_n N_A_304_533#_c_1608_n 0.0134196f $X=1.12 $Y=2.455
+ $X2=0 $Y2=0
cc_579 N_A_196_462#_c_607_n N_A_304_533#_c_1608_n 0.0205416f $X=1.485 $Y=2.137
+ $X2=0 $Y2=0
cc_580 N_A_196_462#_M1015_g N_A_304_533#_c_1609_n 0.0120525f $X=2.72 $Y=2.875
+ $X2=0 $Y2=0
cc_581 N_A_196_462#_c_597_n N_A_304_533#_c_1609_n 0.0176411f $X=2.74 $Y=2.24
+ $X2=0 $Y2=0
cc_582 N_A_196_462#_c_598_n N_A_304_533#_c_1609_n 0.00279821f $X=2.74 $Y=2.24
+ $X2=0 $Y2=0
cc_583 N_A_196_462#_c_601_n N_A_304_533#_c_1609_n 0.00441803f $X=3.455 $Y=2.035
+ $X2=0 $Y2=0
cc_584 N_A_196_462#_c_588_n N_A_304_533#_c_1605_n 0.00561466f $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_585 N_A_196_462#_M1015_g N_A_304_533#_c_1611_n 0.00182823f $X=2.72 $Y=2.875
+ $X2=0 $Y2=0
cc_586 N_A_196_462#_c_597_n N_A_304_533#_c_1611_n 0.015789f $X=2.74 $Y=2.24
+ $X2=0 $Y2=0
cc_587 N_A_196_462#_c_598_n N_A_304_533#_c_1611_n 0.00313854f $X=2.74 $Y=2.24
+ $X2=0 $Y2=0
cc_588 N_A_196_462#_c_599_n N_A_304_533#_c_1611_n 0.0126042f $X=3.85 $Y=1.875
+ $X2=0 $Y2=0
cc_589 N_A_196_462#_c_601_n N_A_304_533#_c_1611_n 0.0195435f $X=3.455 $Y=2.035
+ $X2=0 $Y2=0
cc_590 N_A_196_462#_c_604_n N_A_304_533#_c_1611_n 3.73542e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_591 N_A_196_462#_c_597_n N_A_304_533#_c_1612_n 0.0179742f $X=2.74 $Y=2.24
+ $X2=0 $Y2=0
cc_592 N_A_196_462#_c_598_n N_A_304_533#_c_1612_n 0.00163335f $X=2.74 $Y=2.24
+ $X2=0 $Y2=0
cc_593 N_A_196_462#_c_597_n N_A_304_533#_c_1613_n 0.00259173f $X=2.74 $Y=2.24
+ $X2=0 $Y2=0
cc_594 N_A_196_462#_c_598_n N_A_304_533#_c_1613_n 9.34852e-19 $X=2.74 $Y=2.24
+ $X2=0 $Y2=0
cc_595 N_A_196_462#_c_599_n N_A_304_533#_c_1613_n 0.0050339f $X=3.85 $Y=1.875
+ $X2=0 $Y2=0
cc_596 N_A_196_462#_c_588_n N_A_304_533#_c_1613_n 0.00351315f $X=3.85 $Y=1.47
+ $X2=0 $Y2=0
cc_597 N_A_196_462#_c_601_n N_A_304_533#_c_1613_n 0.0122951f $X=3.455 $Y=2.035
+ $X2=0 $Y2=0
cc_598 N_A_196_462#_c_604_n N_A_304_533#_c_1613_n 2.49749e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_599 N_A_196_462#_M1031_g N_VGND_c_1701_n 8.34806e-19 $X=6.16 $Y=0.765 $X2=0
+ $Y2=0
cc_600 N_A_695_375#_M1018_g N_RESET_B_c_892_n 0.00743797f $X=4.3 $Y=0.955 $X2=0
+ $Y2=0
cc_601 N_A_695_375#_M1029_g N_RESET_B_c_902_n 0.0192094f $X=3.55 $Y=2.875 $X2=0
+ $Y2=0
cc_602 N_A_695_375#_c_790_n N_RESET_B_c_902_n 0.0193903f $X=4.225 $Y=1.95 $X2=0
+ $Y2=0
cc_603 N_A_695_375#_M1018_g N_RESET_B_M1014_g 0.0244377f $X=4.3 $Y=0.955 $X2=0
+ $Y2=0
cc_604 N_A_695_375#_c_783_n N_RESET_B_M1014_g 0.012019f $X=5.665 $Y=1.58 $X2=0
+ $Y2=0
cc_605 N_A_695_375#_c_785_n N_RESET_B_M1014_g 0.00268792f $X=4.39 $Y=1.52 $X2=0
+ $Y2=0
cc_606 N_A_695_375#_c_786_n N_RESET_B_M1014_g 0.0435538f $X=4.39 $Y=1.52 $X2=0
+ $Y2=0
cc_607 N_A_695_375#_M1012_d N_RESET_B_c_907_n 0.00671307f $X=5.825 $Y=2.255
+ $X2=0 $Y2=0
cc_608 N_A_695_375#_c_809_n N_RESET_B_c_907_n 0.0083139f $X=6.035 $Y=2.38 $X2=0
+ $Y2=0
cc_609 N_A_695_375#_M1012_d N_RESET_B_c_933_n 0.0049542f $X=5.825 $Y=2.255 $X2=0
+ $Y2=0
cc_610 N_A_695_375#_c_809_n N_RESET_B_c_933_n 0.0082346f $X=6.035 $Y=2.38 $X2=0
+ $Y2=0
cc_611 N_A_695_375#_c_787_n N_A_559_533#_c_1075_n 0.0040101f $X=5.83 $Y=0.96
+ $X2=0 $Y2=0
cc_612 N_A_695_375#_c_783_n N_A_559_533#_c_1080_n 0.00454312f $X=5.665 $Y=1.58
+ $X2=0 $Y2=0
cc_613 N_A_695_375#_c_794_n N_A_559_533#_c_1080_n 0.00496769f $X=5.85 $Y=2.265
+ $X2=0 $Y2=0
cc_614 N_A_695_375#_c_788_n N_A_559_533#_c_1080_n 0.00422132f $X=5.8 $Y=1.58
+ $X2=0 $Y2=0
cc_615 N_A_695_375#_c_794_n N_A_559_533#_M1012_g 0.00431972f $X=5.85 $Y=2.265
+ $X2=0 $Y2=0
cc_616 N_A_695_375#_c_809_n N_A_559_533#_M1012_g 0.0122613f $X=6.035 $Y=2.38
+ $X2=0 $Y2=0
cc_617 N_A_695_375#_M1029_g N_A_559_533#_c_1099_n 0.00664262f $X=3.55 $Y=2.875
+ $X2=0 $Y2=0
cc_618 N_A_695_375#_M1029_g N_A_559_533#_c_1082_n 0.00581307f $X=3.55 $Y=2.875
+ $X2=0 $Y2=0
cc_619 N_A_695_375#_M1029_g N_A_559_533#_c_1083_n 0.00475318f $X=3.55 $Y=2.875
+ $X2=0 $Y2=0
cc_620 N_A_695_375#_c_790_n N_A_559_533#_c_1083_n 0.0024148f $X=4.225 $Y=1.95
+ $X2=0 $Y2=0
cc_621 N_A_695_375#_M1029_g N_A_559_533#_c_1084_n 0.00425424f $X=3.55 $Y=2.875
+ $X2=0 $Y2=0
cc_622 N_A_695_375#_M1018_g N_A_559_533#_c_1076_n 0.0128779f $X=4.3 $Y=0.955
+ $X2=0 $Y2=0
cc_623 N_A_695_375#_c_783_n N_A_559_533#_c_1076_n 0.0263151f $X=5.665 $Y=1.58
+ $X2=0 $Y2=0
cc_624 N_A_695_375#_c_785_n N_A_559_533#_c_1076_n 0.01942f $X=4.39 $Y=1.52 $X2=0
+ $Y2=0
cc_625 N_A_695_375#_c_786_n N_A_559_533#_c_1076_n 0.00106084f $X=4.39 $Y=1.52
+ $X2=0 $Y2=0
cc_626 N_A_695_375#_M1029_g N_A_559_533#_c_1085_n 5.87988e-19 $X=3.55 $Y=2.875
+ $X2=0 $Y2=0
cc_627 N_A_695_375#_M1029_g N_A_559_533#_c_1086_n 0.00252449f $X=3.55 $Y=2.875
+ $X2=0 $Y2=0
cc_628 N_A_695_375#_c_790_n N_A_559_533#_c_1087_n 0.00105302f $X=4.225 $Y=1.95
+ $X2=0 $Y2=0
cc_629 N_A_695_375#_c_783_n N_A_559_533#_c_1087_n 0.0102259f $X=5.665 $Y=1.58
+ $X2=0 $Y2=0
cc_630 N_A_695_375#_c_785_n N_A_559_533#_c_1087_n 0.00850757f $X=4.39 $Y=1.52
+ $X2=0 $Y2=0
cc_631 N_A_695_375#_M1029_g N_A_559_533#_c_1088_n 0.00333898f $X=3.55 $Y=2.875
+ $X2=0 $Y2=0
cc_632 N_A_695_375#_c_790_n N_A_559_533#_c_1088_n 0.00252998f $X=4.225 $Y=1.95
+ $X2=0 $Y2=0
cc_633 N_A_695_375#_c_785_n N_A_559_533#_c_1088_n 0.0129951f $X=4.39 $Y=1.52
+ $X2=0 $Y2=0
cc_634 N_A_695_375#_M1018_g N_A_559_533#_c_1125_n 0.00339057f $X=4.3 $Y=0.955
+ $X2=0 $Y2=0
cc_635 N_A_695_375#_c_790_n N_A_559_533#_c_1089_n 2.18144e-19 $X=4.225 $Y=1.95
+ $X2=0 $Y2=0
cc_636 N_A_695_375#_c_783_n N_A_559_533#_c_1077_n 0.0234393f $X=5.665 $Y=1.58
+ $X2=0 $Y2=0
cc_637 N_A_695_375#_c_787_n N_A_559_533#_c_1077_n 0.0287726f $X=5.83 $Y=0.96
+ $X2=0 $Y2=0
cc_638 N_A_695_375#_c_783_n N_A_559_533#_c_1090_n 0.0220123f $X=5.665 $Y=1.58
+ $X2=0 $Y2=0
cc_639 N_A_695_375#_c_794_n N_A_559_533#_c_1090_n 0.0196657f $X=5.85 $Y=2.265
+ $X2=0 $Y2=0
cc_640 N_A_695_375#_c_785_n N_A_559_533#_c_1090_n 0.00288732f $X=4.39 $Y=1.52
+ $X2=0 $Y2=0
cc_641 N_A_695_375#_c_809_n N_A_559_533#_c_1090_n 0.00157212f $X=6.035 $Y=2.38
+ $X2=0 $Y2=0
cc_642 N_A_695_375#_c_783_n N_A_559_533#_c_1091_n 0.00154727f $X=5.665 $Y=1.58
+ $X2=0 $Y2=0
cc_643 N_A_695_375#_c_794_n N_A_559_533#_c_1091_n 0.00255927f $X=5.85 $Y=2.265
+ $X2=0 $Y2=0
cc_644 N_A_695_375#_c_783_n N_A_559_533#_c_1078_n 0.00417135f $X=5.665 $Y=1.58
+ $X2=0 $Y2=0
cc_645 N_A_695_375#_c_784_n N_A_559_533#_c_1078_n 0.0040101f $X=5.8 $Y=1.495
+ $X2=0 $Y2=0
cc_646 N_A_695_375#_c_783_n N_A_559_533#_c_1079_n 0.0121666f $X=5.665 $Y=1.58
+ $X2=0 $Y2=0
cc_647 N_A_695_375#_c_784_n N_A_559_533#_c_1079_n 0.00292747f $X=5.8 $Y=1.495
+ $X2=0 $Y2=0
cc_648 N_A_695_375#_c_794_n N_A_559_533#_c_1079_n 0.00249776f $X=5.85 $Y=2.265
+ $X2=0 $Y2=0
cc_649 N_A_695_375#_c_794_n N_A_1247_89#_c_1312_n 0.00541588f $X=5.85 $Y=2.265
+ $X2=0 $Y2=0
cc_650 N_A_695_375#_M1029_g N_VPWR_c_1469_n 0.00475138f $X=3.55 $Y=2.875 $X2=0
+ $Y2=0
cc_651 N_A_695_375#_M1029_g N_VPWR_c_1473_n 0.00371521f $X=3.55 $Y=2.875 $X2=0
+ $Y2=0
cc_652 N_A_695_375#_M1012_d N_VPWR_c_1466_n 0.00318038f $X=5.825 $Y=2.255 $X2=0
+ $Y2=0
cc_653 N_A_695_375#_M1029_g N_VPWR_c_1466_n 0.00562668f $X=3.55 $Y=2.875 $X2=0
+ $Y2=0
cc_654 N_A_695_375#_M1029_g N_A_304_533#_c_1611_n 0.0017691f $X=3.55 $Y=2.875
+ $X2=0 $Y2=0
cc_655 N_A_695_375#_c_791_n N_A_304_533#_c_1611_n 3.48151e-19 $X=3.625 $Y=1.95
+ $X2=0 $Y2=0
cc_656 N_RESET_B_c_892_n N_A_559_533#_c_1075_n 0.0188764f $X=4.765 $Y=0.3 $X2=0
+ $Y2=0
cc_657 N_RESET_B_c_906_n N_A_559_533#_M1012_g 0.009771f $X=5.765 $Y=2.72 $X2=0
+ $Y2=0
cc_658 N_RESET_B_c_907_n N_A_559_533#_M1012_g 3.03723e-19 $X=7.225 $Y=2.99 $X2=0
+ $Y2=0
cc_659 N_RESET_B_c_933_n N_A_559_533#_M1012_g 0.0153755f $X=5.85 $Y=2.72 $X2=0
+ $Y2=0
cc_660 N_RESET_B_c_900_n N_A_559_533#_c_1082_n 5.71856e-19 $X=4.085 $Y=2.545
+ $X2=0 $Y2=0
cc_661 N_RESET_B_c_900_n N_A_559_533#_c_1083_n 0.00522226f $X=4.085 $Y=2.545
+ $X2=0 $Y2=0
cc_662 N_RESET_B_c_902_n N_A_559_533#_c_1083_n 0.00356673f $X=4.16 $Y=2.47 $X2=0
+ $Y2=0
cc_663 N_RESET_B_M1014_g N_A_559_533#_c_1076_n 0.0141489f $X=4.84 $Y=0.745 $X2=0
+ $Y2=0
cc_664 N_RESET_B_c_900_n N_A_559_533#_c_1085_n 0.00635942f $X=4.085 $Y=2.545
+ $X2=0 $Y2=0
cc_665 N_RESET_B_c_976_p N_A_559_533#_c_1085_n 0.0283158f $X=4.75 $Y=2.56 $X2=0
+ $Y2=0
cc_666 N_RESET_B_c_910_n N_A_559_533#_c_1085_n 0.00427871f $X=4.75 $Y=2.56 $X2=0
+ $Y2=0
cc_667 N_RESET_B_c_901_n N_A_559_533#_c_1086_n 0.00656475f $X=4.585 $Y=2.47
+ $X2=0 $Y2=0
cc_668 N_RESET_B_M1014_g N_A_559_533#_c_1086_n 2.76286e-19 $X=4.84 $Y=0.745
+ $X2=0 $Y2=0
cc_669 N_RESET_B_c_901_n N_A_559_533#_c_1087_n 0.00983999f $X=4.585 $Y=2.47
+ $X2=0 $Y2=0
cc_670 N_RESET_B_M1014_g N_A_559_533#_c_1087_n 0.0147143f $X=4.84 $Y=0.745 $X2=0
+ $Y2=0
cc_671 N_RESET_B_c_906_n N_A_559_533#_c_1087_n 0.00979089f $X=5.765 $Y=2.72
+ $X2=0 $Y2=0
cc_672 N_RESET_B_c_976_p N_A_559_533#_c_1087_n 0.0224038f $X=4.75 $Y=2.56 $X2=0
+ $Y2=0
cc_673 N_RESET_B_c_900_n N_A_559_533#_c_1089_n 9.64993e-19 $X=4.085 $Y=2.545
+ $X2=0 $Y2=0
cc_674 N_RESET_B_c_901_n N_A_559_533#_c_1089_n 0.00879464f $X=4.585 $Y=2.47
+ $X2=0 $Y2=0
cc_675 N_RESET_B_c_902_n N_A_559_533#_c_1089_n 2.42145e-19 $X=4.16 $Y=2.47 $X2=0
+ $Y2=0
cc_676 N_RESET_B_c_976_p N_A_559_533#_c_1089_n 0.0114534f $X=4.75 $Y=2.56 $X2=0
+ $Y2=0
cc_677 N_RESET_B_c_910_n N_A_559_533#_c_1089_n 6.10593e-19 $X=4.75 $Y=2.56 $X2=0
+ $Y2=0
cc_678 N_RESET_B_M1014_g N_A_559_533#_c_1077_n 0.00135923f $X=4.84 $Y=0.745
+ $X2=0 $Y2=0
cc_679 N_RESET_B_M1014_g N_A_559_533#_c_1090_n 0.00350706f $X=4.84 $Y=0.745
+ $X2=0 $Y2=0
cc_680 N_RESET_B_c_906_n N_A_559_533#_c_1090_n 0.0140334f $X=5.765 $Y=2.72 $X2=0
+ $Y2=0
cc_681 N_RESET_B_c_906_n N_A_559_533#_c_1091_n 0.00429327f $X=5.765 $Y=2.72
+ $X2=0 $Y2=0
cc_682 N_RESET_B_M1014_g N_A_559_533#_c_1078_n 0.0584323f $X=4.84 $Y=0.745 $X2=0
+ $Y2=0
cc_683 N_RESET_B_M1003_g N_A_1467_419#_M1016_g 0.0104552f $X=8.11 $Y=2.795 $X2=0
+ $Y2=0
cc_684 N_RESET_B_c_907_n N_A_1467_419#_M1016_g 0.00533768f $X=7.225 $Y=2.99
+ $X2=0 $Y2=0
cc_685 N_RESET_B_c_909_n N_A_1467_419#_M1016_g 0.0128907f $X=7.31 $Y=2.905 $X2=0
+ $Y2=0
cc_686 N_RESET_B_M1001_g N_A_1467_419#_M1000_g 0.0452f $X=7.89 $Y=0.875 $X2=0
+ $Y2=0
cc_687 N_RESET_B_M1003_g N_A_1467_419#_M1000_g 0.00527981f $X=8.11 $Y=2.795
+ $X2=0 $Y2=0
cc_688 N_RESET_B_c_896_n N_A_1467_419#_M1000_g 0.00283556f $X=7.31 $Y=1.885
+ $X2=0 $Y2=0
cc_689 N_RESET_B_c_909_n N_A_1467_419#_M1000_g 0.00546195f $X=7.31 $Y=2.905
+ $X2=0 $Y2=0
cc_690 N_RESET_B_c_897_n N_A_1467_419#_M1000_g 0.0167089f $X=7.98 $Y=1.72 $X2=0
+ $Y2=0
cc_691 N_RESET_B_M1003_g N_A_1467_419#_c_1231_n 0.0150551f $X=8.11 $Y=2.795
+ $X2=0 $Y2=0
cc_692 N_RESET_B_c_909_n N_A_1467_419#_c_1231_n 0.0248018f $X=7.31 $Y=2.905
+ $X2=0 $Y2=0
cc_693 N_RESET_B_c_897_n N_A_1467_419#_c_1231_n 0.038688f $X=7.98 $Y=1.72 $X2=0
+ $Y2=0
cc_694 N_RESET_B_c_898_n N_A_1467_419#_c_1231_n 0.00523955f $X=8.11 $Y=1.72
+ $X2=0 $Y2=0
cc_695 N_RESET_B_M1003_g N_A_1467_419#_c_1232_n 0.0213808f $X=8.11 $Y=2.795
+ $X2=0 $Y2=0
cc_696 N_RESET_B_c_909_n N_A_1467_419#_c_1232_n 0.00988262f $X=7.31 $Y=2.905
+ $X2=0 $Y2=0
cc_697 N_RESET_B_c_897_n N_A_1467_419#_c_1232_n 0.00675699f $X=7.98 $Y=1.72
+ $X2=0 $Y2=0
cc_698 N_RESET_B_c_898_n N_A_1467_419#_c_1232_n 6.47558e-19 $X=8.11 $Y=1.72
+ $X2=0 $Y2=0
cc_699 N_RESET_B_M1003_g N_A_1467_419#_c_1233_n 0.0106908f $X=8.11 $Y=2.795
+ $X2=0 $Y2=0
cc_700 N_RESET_B_M1001_g N_A_1467_419#_c_1227_n 8.89028e-19 $X=7.89 $Y=0.875
+ $X2=0 $Y2=0
cc_701 N_RESET_B_M1003_g N_A_1467_419#_c_1236_n 0.00585482f $X=8.11 $Y=2.795
+ $X2=0 $Y2=0
cc_702 N_RESET_B_c_907_n N_A_1247_89#_M1011_d 0.00486719f $X=7.225 $Y=2.99 $X2=0
+ $Y2=0
cc_703 N_RESET_B_M1001_g N_A_1247_89#_c_1304_n 0.0494163f $X=7.89 $Y=0.875 $X2=0
+ $Y2=0
cc_704 N_RESET_B_c_898_n N_A_1247_89#_M1008_g 0.0392301f $X=8.11 $Y=1.72 $X2=0
+ $Y2=0
cc_705 N_RESET_B_c_898_n N_A_1247_89#_c_1309_n 6.67584e-19 $X=8.11 $Y=1.72 $X2=0
+ $Y2=0
cc_706 N_RESET_B_M1001_g N_A_1247_89#_c_1311_n 0.0138719f $X=7.89 $Y=0.875 $X2=0
+ $Y2=0
cc_707 N_RESET_B_c_896_n N_A_1247_89#_c_1311_n 0.0131874f $X=7.31 $Y=1.885 $X2=0
+ $Y2=0
cc_708 N_RESET_B_c_897_n N_A_1247_89#_c_1311_n 0.0518816f $X=7.98 $Y=1.72 $X2=0
+ $Y2=0
cc_709 N_RESET_B_c_898_n N_A_1247_89#_c_1311_n 0.00583141f $X=8.11 $Y=1.72 $X2=0
+ $Y2=0
cc_710 N_RESET_B_c_907_n N_A_1247_89#_c_1319_n 0.0196796f $X=7.225 $Y=2.99 $X2=0
+ $Y2=0
cc_711 N_RESET_B_c_933_n N_A_1247_89#_c_1319_n 0.00396914f $X=5.85 $Y=2.72 $X2=0
+ $Y2=0
cc_712 N_RESET_B_c_909_n N_A_1247_89#_c_1312_n 0.0154424f $X=7.31 $Y=2.905 $X2=0
+ $Y2=0
cc_713 N_RESET_B_M1001_g N_A_1247_89#_c_1314_n 0.0010658f $X=7.89 $Y=0.875 $X2=0
+ $Y2=0
cc_714 N_RESET_B_c_897_n N_A_1247_89#_c_1314_n 0.0177637f $X=7.98 $Y=1.72 $X2=0
+ $Y2=0
cc_715 N_RESET_B_c_898_n N_A_1247_89#_c_1314_n 0.00114018f $X=8.11 $Y=1.72 $X2=0
+ $Y2=0
cc_716 N_RESET_B_M1001_g N_A_1247_89#_c_1315_n 0.00630584f $X=7.89 $Y=0.875
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_897_n N_A_1247_89#_c_1315_n 0.0010088f $X=7.98 $Y=1.72 $X2=0
+ $Y2=0
cc_718 N_RESET_B_c_898_n N_A_1247_89#_c_1315_n 0.0191641f $X=8.11 $Y=1.72 $X2=0
+ $Y2=0
cc_719 N_RESET_B_c_906_n N_VPWR_M1012_s 0.00930157f $X=5.765 $Y=2.72 $X2=0 $Y2=0
cc_720 N_RESET_B_M1007_g N_VPWR_c_1468_n 0.00926909f $X=1.86 $Y=2.875 $X2=0
+ $Y2=0
cc_721 N_RESET_B_c_900_n N_VPWR_c_1469_n 0.00296786f $X=4.085 $Y=2.545 $X2=0
+ $Y2=0
cc_722 N_RESET_B_M1003_g N_VPWR_c_1470_n 0.00795407f $X=8.11 $Y=2.795 $X2=0
+ $Y2=0
cc_723 N_RESET_B_c_907_n N_VPWR_c_1470_n 0.014145f $X=7.225 $Y=2.99 $X2=0 $Y2=0
cc_724 N_RESET_B_c_909_n N_VPWR_c_1470_n 0.0203633f $X=7.31 $Y=2.905 $X2=0 $Y2=0
cc_725 N_RESET_B_c_906_n N_VPWR_c_1475_n 0.0034313f $X=5.765 $Y=2.72 $X2=0 $Y2=0
cc_726 N_RESET_B_c_907_n N_VPWR_c_1475_n 0.0903674f $X=7.225 $Y=2.99 $X2=0 $Y2=0
cc_727 N_RESET_B_c_933_n N_VPWR_c_1475_n 0.00946397f $X=5.85 $Y=2.72 $X2=0 $Y2=0
cc_728 N_RESET_B_M1003_g N_VPWR_c_1477_n 0.0047088f $X=8.11 $Y=2.795 $X2=0 $Y2=0
cc_729 N_RESET_B_M1007_g N_VPWR_c_1480_n 0.00348975f $X=1.86 $Y=2.875 $X2=0
+ $Y2=0
cc_730 N_RESET_B_c_900_n N_VPWR_c_1481_n 0.00422451f $X=4.085 $Y=2.545 $X2=0
+ $Y2=0
cc_731 N_RESET_B_c_906_n N_VPWR_c_1481_n 0.00798338f $X=5.765 $Y=2.72 $X2=0
+ $Y2=0
cc_732 N_RESET_B_c_976_p N_VPWR_c_1481_n 0.0136773f $X=4.75 $Y=2.56 $X2=0 $Y2=0
cc_733 N_RESET_B_c_910_n N_VPWR_c_1481_n 0.00865497f $X=4.75 $Y=2.56 $X2=0 $Y2=0
cc_734 N_RESET_B_M1007_g N_VPWR_c_1466_n 0.00548155f $X=1.86 $Y=2.875 $X2=0
+ $Y2=0
cc_735 N_RESET_B_c_900_n N_VPWR_c_1466_n 0.00739128f $X=4.085 $Y=2.545 $X2=0
+ $Y2=0
cc_736 N_RESET_B_c_901_n N_VPWR_c_1466_n 0.00169585f $X=4.585 $Y=2.47 $X2=0
+ $Y2=0
cc_737 N_RESET_B_M1003_g N_VPWR_c_1466_n 0.00924756f $X=8.11 $Y=2.795 $X2=0
+ $Y2=0
cc_738 N_RESET_B_c_906_n N_VPWR_c_1466_n 0.0176487f $X=5.765 $Y=2.72 $X2=0 $Y2=0
cc_739 N_RESET_B_c_907_n N_VPWR_c_1466_n 0.053462f $X=7.225 $Y=2.99 $X2=0 $Y2=0
cc_740 N_RESET_B_c_976_p N_VPWR_c_1466_n 0.0117745f $X=4.75 $Y=2.56 $X2=0 $Y2=0
cc_741 N_RESET_B_c_910_n N_VPWR_c_1466_n 0.0117576f $X=4.75 $Y=2.56 $X2=0 $Y2=0
cc_742 N_RESET_B_c_933_n N_VPWR_c_1466_n 0.00618975f $X=5.85 $Y=2.72 $X2=0 $Y2=0
cc_743 N_RESET_B_c_906_n N_VPWR_c_1487_n 0.0240991f $X=5.765 $Y=2.72 $X2=0 $Y2=0
cc_744 N_RESET_B_c_976_p N_VPWR_c_1487_n 4.72826e-19 $X=4.75 $Y=2.56 $X2=0 $Y2=0
cc_745 N_RESET_B_c_910_n N_VPWR_c_1487_n 0.00290215f $X=4.75 $Y=2.56 $X2=0 $Y2=0
cc_746 N_RESET_B_c_933_n N_VPWR_c_1487_n 0.00708052f $X=5.85 $Y=2.72 $X2=0 $Y2=0
cc_747 N_RESET_B_M1007_g N_A_304_533#_c_1607_n 0.0130017f $X=1.86 $Y=2.875 $X2=0
+ $Y2=0
cc_748 N_RESET_B_c_907_n A_1379_517# 0.00732703f $X=7.225 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_749 N_RESET_B_c_909_n A_1379_517# 0.00440575f $X=7.31 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_750 N_RESET_B_M1007_g N_VGND_c_1698_n 0.00538482f $X=1.86 $Y=2.875 $X2=0
+ $Y2=0
cc_751 N_RESET_B_c_889_n N_VGND_c_1698_n 0.018267f $X=2.31 $Y=0.3 $X2=0 $Y2=0
cc_752 N_RESET_B_M1010_g N_VGND_c_1698_n 0.0145814f $X=2.385 $Y=0.955 $X2=0
+ $Y2=0
cc_753 N_RESET_B_c_895_n N_VGND_c_1698_n 0.00751259f $X=2.385 $Y=0.3 $X2=0 $Y2=0
cc_754 N_RESET_B_M1001_g N_VGND_c_1699_n 0.0104136f $X=7.89 $Y=0.875 $X2=0 $Y2=0
cc_755 N_RESET_B_c_890_n N_VGND_c_1704_n 0.0064269f $X=1.935 $Y=0.3 $X2=0 $Y2=0
cc_756 N_RESET_B_c_895_n N_VGND_c_1705_n 0.0498401f $X=2.385 $Y=0.3 $X2=0 $Y2=0
cc_757 N_RESET_B_M1001_g N_VGND_c_1706_n 0.0032821f $X=7.89 $Y=0.875 $X2=0 $Y2=0
cc_758 N_RESET_B_c_889_n N_VGND_c_1708_n 0.00417944f $X=2.31 $Y=0.3 $X2=0 $Y2=0
cc_759 N_RESET_B_c_890_n N_VGND_c_1708_n 0.00794683f $X=1.935 $Y=0.3 $X2=0 $Y2=0
cc_760 N_RESET_B_c_892_n N_VGND_c_1708_n 0.0610514f $X=4.765 $Y=0.3 $X2=0 $Y2=0
cc_761 N_RESET_B_M1001_g N_VGND_c_1708_n 0.00385154f $X=7.89 $Y=0.875 $X2=0
+ $Y2=0
cc_762 N_RESET_B_c_895_n N_VGND_c_1708_n 0.00755729f $X=2.385 $Y=0.3 $X2=0 $Y2=0
cc_763 N_RESET_B_c_892_n N_VGND_c_1711_n 0.00392069f $X=4.765 $Y=0.3 $X2=0 $Y2=0
cc_764 N_A_559_533#_c_1090_n N_VPWR_M1012_s 0.00381762f $X=5.32 $Y=1.93 $X2=0
+ $Y2=0
cc_765 N_A_559_533#_c_1099_n N_VPWR_c_1469_n 0.0184082f $X=3.415 $Y=2.96 $X2=0
+ $Y2=0
cc_766 N_A_559_533#_c_1082_n N_VPWR_c_1469_n 0.00354788f $X=3.5 $Y=2.845 $X2=0
+ $Y2=0
cc_767 N_A_559_533#_c_1083_n N_VPWR_c_1469_n 0.0155633f $X=4.145 $Y=2.53 $X2=0
+ $Y2=0
cc_768 N_A_559_533#_c_1099_n N_VPWR_c_1473_n 0.0437869f $X=3.415 $Y=2.96 $X2=0
+ $Y2=0
cc_769 N_A_559_533#_c_1083_n N_VPWR_c_1473_n 0.00254765f $X=4.145 $Y=2.53 $X2=0
+ $Y2=0
cc_770 N_A_559_533#_M1012_g N_VPWR_c_1475_n 0.00389381f $X=5.75 $Y=2.675 $X2=0
+ $Y2=0
cc_771 N_A_559_533#_c_1083_n N_VPWR_c_1481_n 0.002372f $X=4.145 $Y=2.53 $X2=0
+ $Y2=0
cc_772 N_A_559_533#_c_1085_n N_VPWR_c_1481_n 0.0133686f $X=4.3 $Y=2.87 $X2=0
+ $Y2=0
cc_773 N_A_559_533#_M1015_d N_VPWR_c_1466_n 0.00261173f $X=2.795 $Y=2.665 $X2=0
+ $Y2=0
cc_774 N_A_559_533#_M1022_d N_VPWR_c_1466_n 0.00228073f $X=4.16 $Y=2.665 $X2=0
+ $Y2=0
cc_775 N_A_559_533#_M1012_g N_VPWR_c_1466_n 0.00737537f $X=5.75 $Y=2.675 $X2=0
+ $Y2=0
cc_776 N_A_559_533#_c_1099_n N_VPWR_c_1466_n 0.028214f $X=3.415 $Y=2.96 $X2=0
+ $Y2=0
cc_777 N_A_559_533#_c_1083_n N_VPWR_c_1466_n 0.00911237f $X=4.145 $Y=2.53 $X2=0
+ $Y2=0
cc_778 N_A_559_533#_c_1085_n N_VPWR_c_1466_n 0.0101282f $X=4.3 $Y=2.87 $X2=0
+ $Y2=0
cc_779 N_A_559_533#_M1012_g N_VPWR_c_1487_n 0.00712182f $X=5.75 $Y=2.675 $X2=0
+ $Y2=0
cc_780 N_A_559_533#_M1015_d N_A_304_533#_c_1609_n 0.00211743f $X=2.795 $Y=2.665
+ $X2=0 $Y2=0
cc_781 N_A_559_533#_c_1099_n N_A_304_533#_c_1609_n 0.0241781f $X=3.415 $Y=2.96
+ $X2=0 $Y2=0
cc_782 N_A_559_533#_c_1082_n N_A_304_533#_c_1609_n 0.00474389f $X=3.5 $Y=2.845
+ $X2=0 $Y2=0
cc_783 N_A_559_533#_c_1084_n N_A_304_533#_c_1609_n 0.00980672f $X=3.585 $Y=2.53
+ $X2=0 $Y2=0
cc_784 N_A_559_533#_c_1084_n N_A_304_533#_c_1611_n 0.00480683f $X=3.585 $Y=2.53
+ $X2=0 $Y2=0
cc_785 N_A_559_533#_c_1099_n A_653_533# 0.00451309f $X=3.415 $Y=2.96 $X2=-0.19
+ $Y2=-0.245
cc_786 N_A_559_533#_c_1082_n A_653_533# 0.00201007f $X=3.5 $Y=2.845 $X2=-0.19
+ $Y2=-0.245
cc_787 N_A_559_533#_c_1076_n N_VGND_M1014_d 0.00227919f $X=5.155 $Y=1.035 $X2=0
+ $Y2=0
cc_788 N_A_559_533#_c_1077_n N_VGND_M1014_d 0.00267456f $X=5.32 $Y=1.035 $X2=0
+ $Y2=0
cc_789 N_A_559_533#_c_1075_n N_VGND_c_1701_n 0.00329948f $X=5.5 $Y=1.065 $X2=0
+ $Y2=0
cc_790 N_A_559_533#_c_1075_n N_VGND_c_1708_n 0.00576296f $X=5.5 $Y=1.065 $X2=0
+ $Y2=0
cc_791 N_A_559_533#_c_1075_n N_VGND_c_1711_n 0.00300633f $X=5.5 $Y=1.065 $X2=0
+ $Y2=0
cc_792 N_A_559_533#_c_1076_n A_803_149# 0.00112882f $X=5.155 $Y=1.035 $X2=-0.19
+ $Y2=-0.245
cc_793 N_A_559_533#_c_1125_n A_803_149# 0.00522443f $X=4.145 $Y=0.975 $X2=-0.19
+ $Y2=-0.245
cc_794 N_A_559_533#_c_1076_n A_875_149# 0.00564184f $X=5.155 $Y=1.035 $X2=-0.19
+ $Y2=-0.245
cc_795 N_A_1467_419#_c_1227_n N_A_1247_89#_c_1304_n 0.00603276f $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_796 N_A_1467_419#_c_1228_n N_A_1247_89#_c_1304_n 0.00373494f $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_797 N_A_1467_419#_c_1233_n N_A_1247_89#_M1008_g 0.00460242f $X=8.325 $Y=2.795
+ $X2=0 $Y2=0
cc_798 N_A_1467_419#_c_1234_n N_A_1247_89#_M1008_g 0.0149048f $X=8.825 $Y=2.18
+ $X2=0 $Y2=0
cc_799 N_A_1467_419#_c_1228_n N_A_1247_89#_M1008_g 0.00750966f $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_800 N_A_1467_419#_c_1236_n N_A_1247_89#_M1008_g 0.0110747f $X=8.312 $Y=2.26
+ $X2=0 $Y2=0
cc_801 N_A_1467_419#_c_1228_n N_A_1247_89#_c_1305_n 0.0142898f $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_802 N_A_1467_419#_c_1227_n N_A_1247_89#_c_1306_n 3.57913e-19 $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_803 N_A_1467_419#_c_1228_n N_A_1247_89#_c_1306_n 6.74571e-19 $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_804 N_A_1467_419#_c_1228_n N_A_1247_89#_M1023_g 7.27987e-19 $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_805 N_A_1467_419#_c_1227_n N_A_1247_89#_M1017_g 7.62659e-19 $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_806 N_A_1467_419#_c_1227_n N_A_1247_89#_c_1309_n 0.00915388f $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_807 N_A_1467_419#_c_1234_n N_A_1247_89#_c_1318_n 0.00299181f $X=8.825 $Y=2.18
+ $X2=0 $Y2=0
cc_808 N_A_1467_419#_c_1236_n N_A_1247_89#_c_1318_n 5.21175e-19 $X=8.312 $Y=2.26
+ $X2=0 $Y2=0
cc_809 N_A_1467_419#_M1000_g N_A_1247_89#_c_1311_n 0.0160561f $X=7.46 $Y=0.875
+ $X2=0 $Y2=0
cc_810 N_A_1467_419#_c_1227_n N_A_1247_89#_c_1311_n 0.00460758f $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_811 N_A_1467_419#_M1000_g N_A_1247_89#_c_1312_n 8.25022e-19 $X=7.46 $Y=0.875
+ $X2=0 $Y2=0
cc_812 N_A_1467_419#_c_1227_n N_A_1247_89#_c_1314_n 0.0214989f $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_813 N_A_1467_419#_c_1234_n N_A_1247_89#_c_1314_n 0.0114023f $X=8.825 $Y=2.18
+ $X2=0 $Y2=0
cc_814 N_A_1467_419#_c_1228_n N_A_1247_89#_c_1314_n 0.0498119f $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_815 N_A_1467_419#_c_1236_n N_A_1247_89#_c_1314_n 0.00489233f $X=8.312 $Y=2.26
+ $X2=0 $Y2=0
cc_816 N_A_1467_419#_c_1228_n N_A_1247_89#_c_1315_n 0.0063593f $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_817 N_A_1467_419#_c_1227_n N_A_1832_367#_c_1419_n 0.029425f $X=8.825 $Y=0.86
+ $X2=0 $Y2=0
cc_818 N_A_1467_419#_c_1228_n N_A_1832_367#_c_1419_n 0.0235646f $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_819 N_A_1467_419#_c_1234_n N_A_1832_367#_c_1425_n 0.0143977f $X=8.825 $Y=2.18
+ $X2=0 $Y2=0
cc_820 N_A_1467_419#_c_1228_n N_A_1832_367#_c_1425_n 0.0326383f $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_821 N_A_1467_419#_c_1228_n N_A_1832_367#_c_1422_n 0.0277882f $X=8.91 $Y=2.095
+ $X2=0 $Y2=0
cc_822 N_A_1467_419#_M1016_g N_VPWR_c_1470_n 0.00596873f $X=7.41 $Y=2.795 $X2=0
+ $Y2=0
cc_823 N_A_1467_419#_c_1231_n N_VPWR_c_1470_n 0.0244885f $X=8.16 $Y=2.26 $X2=0
+ $Y2=0
cc_824 N_A_1467_419#_c_1232_n N_VPWR_c_1470_n 0.00592599f $X=7.66 $Y=2.26 $X2=0
+ $Y2=0
cc_825 N_A_1467_419#_c_1233_n N_VPWR_c_1470_n 0.0187069f $X=8.325 $Y=2.795 $X2=0
+ $Y2=0
cc_826 N_A_1467_419#_c_1234_n N_VPWR_c_1471_n 0.0131255f $X=8.825 $Y=2.18 $X2=0
+ $Y2=0
cc_827 N_A_1467_419#_M1016_g N_VPWR_c_1475_n 0.0042066f $X=7.41 $Y=2.795 $X2=0
+ $Y2=0
cc_828 N_A_1467_419#_c_1233_n N_VPWR_c_1477_n 0.00997522f $X=8.325 $Y=2.795
+ $X2=0 $Y2=0
cc_829 N_A_1467_419#_M1016_g N_VPWR_c_1466_n 0.00798794f $X=7.41 $Y=2.795 $X2=0
+ $Y2=0
cc_830 N_A_1467_419#_c_1233_n N_VPWR_c_1466_n 0.0109258f $X=8.325 $Y=2.795 $X2=0
+ $Y2=0
cc_831 N_A_1467_419#_M1000_g N_VGND_c_1699_n 0.0114811f $X=7.46 $Y=0.875 $X2=0
+ $Y2=0
cc_832 N_A_1467_419#_c_1227_n N_VGND_c_1699_n 0.01166f $X=8.825 $Y=0.86 $X2=0
+ $Y2=0
cc_833 N_A_1467_419#_M1000_g N_VGND_c_1701_n 0.0032821f $X=7.46 $Y=0.875 $X2=0
+ $Y2=0
cc_834 N_A_1467_419#_c_1227_n N_VGND_c_1706_n 0.0112173f $X=8.825 $Y=0.86 $X2=0
+ $Y2=0
cc_835 N_A_1467_419#_M1000_g N_VGND_c_1708_n 0.00385154f $X=7.46 $Y=0.875 $X2=0
+ $Y2=0
cc_836 N_A_1467_419#_c_1227_n N_VGND_c_1708_n 0.0196111f $X=8.825 $Y=0.86 $X2=0
+ $Y2=0
cc_837 N_A_1247_89#_M1023_g N_A_1832_367#_M1024_g 0.0116128f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_838 N_A_1247_89#_c_1305_n N_A_1832_367#_c_1419_n 0.00941398f $X=9.425 $Y=1.27
+ $X2=0 $Y2=0
cc_839 N_A_1247_89#_c_1306_n N_A_1832_367#_c_1419_n 0.014703f $X=9.5 $Y=1.345
+ $X2=0 $Y2=0
cc_840 N_A_1247_89#_M1017_g N_A_1832_367#_c_1419_n 0.00875644f $X=9.575 $Y=0.595
+ $X2=0 $Y2=0
cc_841 N_A_1247_89#_M1008_g N_A_1832_367#_c_1425_n 0.00620472f $X=8.54 $Y=2.795
+ $X2=0 $Y2=0
cc_842 N_A_1247_89#_M1023_g N_A_1832_367#_c_1425_n 0.00550743f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_843 N_A_1247_89#_c_1306_n N_A_1832_367#_c_1420_n 0.00555047f $X=9.5 $Y=1.345
+ $X2=0 $Y2=0
cc_844 N_A_1247_89#_M1023_g N_A_1832_367#_c_1420_n 0.00665567f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_845 N_A_1247_89#_c_1306_n N_A_1832_367#_c_1421_n 0.021329f $X=9.5 $Y=1.345
+ $X2=0 $Y2=0
cc_846 N_A_1247_89#_c_1305_n N_A_1832_367#_c_1422_n 0.00448416f $X=9.425 $Y=1.27
+ $X2=0 $Y2=0
cc_847 N_A_1247_89#_M1023_g N_A_1832_367#_c_1422_n 0.0133801f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_848 N_A_1247_89#_c_1306_n N_A_1832_367#_c_1423_n 0.00448381f $X=9.5 $Y=1.345
+ $X2=0 $Y2=0
cc_849 N_A_1247_89#_M1017_g N_A_1832_367#_c_1423_n 0.0148089f $X=9.575 $Y=0.595
+ $X2=0 $Y2=0
cc_850 N_A_1247_89#_M1008_g N_VPWR_c_1471_n 0.00553306f $X=8.54 $Y=2.795 $X2=0
+ $Y2=0
cc_851 N_A_1247_89#_M1023_g N_VPWR_c_1472_n 0.00520367f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_852 N_A_1247_89#_M1008_g N_VPWR_c_1477_n 0.00499542f $X=8.54 $Y=2.795 $X2=0
+ $Y2=0
cc_853 N_A_1247_89#_M1023_g N_VPWR_c_1482_n 0.00312414f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_854 N_A_1247_89#_M1011_d N_VPWR_c_1466_n 0.00212318f $X=6.37 $Y=2.245 $X2=0
+ $Y2=0
cc_855 N_A_1247_89#_M1008_g N_VPWR_c_1466_n 0.0102383f $X=8.54 $Y=2.795 $X2=0
+ $Y2=0
cc_856 N_A_1247_89#_M1023_g N_VPWR_c_1466_n 0.00410284f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_857 N_A_1247_89#_c_1304_n N_VGND_c_1699_n 0.00170478f $X=8.25 $Y=1.195 $X2=0
+ $Y2=0
cc_858 N_A_1247_89#_c_1311_n N_VGND_c_1699_n 0.0216087f $X=8.395 $Y=1.28 $X2=0
+ $Y2=0
cc_859 N_A_1247_89#_c_1306_n N_VGND_c_1700_n 5.76509e-19 $X=9.5 $Y=1.345 $X2=0
+ $Y2=0
cc_860 N_A_1247_89#_M1017_g N_VGND_c_1700_n 0.0085264f $X=9.575 $Y=0.595 $X2=0
+ $Y2=0
cc_861 N_A_1247_89#_c_1304_n N_VGND_c_1706_n 0.00380579f $X=8.25 $Y=1.195 $X2=0
+ $Y2=0
cc_862 N_A_1247_89#_M1017_g N_VGND_c_1706_n 0.00542223f $X=9.575 $Y=0.595 $X2=0
+ $Y2=0
cc_863 N_A_1247_89#_c_1304_n N_VGND_c_1708_n 0.00458517f $X=8.25 $Y=1.195 $X2=0
+ $Y2=0
cc_864 N_A_1247_89#_M1017_g N_VGND_c_1708_n 0.0054106f $X=9.575 $Y=0.595 $X2=0
+ $Y2=0
cc_865 N_A_1832_367#_M1024_g N_VPWR_c_1472_n 0.0230777f $X=10.01 $Y=2.465 $X2=0
+ $Y2=0
cc_866 N_A_1832_367#_c_1425_n N_VPWR_c_1472_n 0.0010381f $X=9.285 $Y=1.985 $X2=0
+ $Y2=0
cc_867 N_A_1832_367#_c_1420_n N_VPWR_c_1472_n 0.0257576f $X=9.95 $Y=1.5 $X2=0
+ $Y2=0
cc_868 N_A_1832_367#_c_1421_n N_VPWR_c_1472_n 0.00329759f $X=9.95 $Y=1.5 $X2=0
+ $Y2=0
cc_869 N_A_1832_367#_M1024_g N_VPWR_c_1483_n 0.00486043f $X=10.01 $Y=2.465 $X2=0
+ $Y2=0
cc_870 N_A_1832_367#_M1024_g N_VPWR_c_1466_n 0.00924348f $X=10.01 $Y=2.465 $X2=0
+ $Y2=0
cc_871 N_A_1832_367#_c_1425_n N_VPWR_c_1466_n 0.0087929f $X=9.285 $Y=1.985 $X2=0
+ $Y2=0
cc_872 N_A_1832_367#_c_1421_n N_Q_c_1685_n 0.00112485f $X=9.95 $Y=1.5 $X2=0
+ $Y2=0
cc_873 N_A_1832_367#_M1024_g Q 0.00665999f $X=10.01 $Y=2.465 $X2=0 $Y2=0
cc_874 N_A_1832_367#_c_1420_n Q 0.0271104f $X=9.95 $Y=1.5 $X2=0 $Y2=0
cc_875 N_A_1832_367#_c_1423_n Q 0.0170182f $X=9.972 $Y=1.335 $X2=0 $Y2=0
cc_876 N_A_1832_367#_c_1419_n N_VGND_c_1700_n 0.042915f $X=9.36 $Y=0.595 $X2=0
+ $Y2=0
cc_877 N_A_1832_367#_c_1420_n N_VGND_c_1700_n 0.0256984f $X=9.95 $Y=1.5 $X2=0
+ $Y2=0
cc_878 N_A_1832_367#_c_1421_n N_VGND_c_1700_n 0.00536365f $X=9.95 $Y=1.5 $X2=0
+ $Y2=0
cc_879 N_A_1832_367#_c_1423_n N_VGND_c_1700_n 0.0176733f $X=9.972 $Y=1.335 $X2=0
+ $Y2=0
cc_880 N_A_1832_367#_c_1419_n N_VGND_c_1706_n 0.0108386f $X=9.36 $Y=0.595 $X2=0
+ $Y2=0
cc_881 N_A_1832_367#_c_1423_n N_VGND_c_1707_n 0.00471276f $X=9.972 $Y=1.335
+ $X2=0 $Y2=0
cc_882 N_A_1832_367#_c_1419_n N_VGND_c_1708_n 0.0125299f $X=9.36 $Y=0.595 $X2=0
+ $Y2=0
cc_883 N_A_1832_367#_c_1423_n N_VGND_c_1708_n 0.0045449f $X=9.972 $Y=1.335 $X2=0
+ $Y2=0
cc_884 N_VPWR_c_1466_n N_A_304_533#_M1007_s 0.00231379f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_885 N_VPWR_c_1466_n N_A_304_533#_M1021_d 0.00244643f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_886 N_VPWR_c_1467_n N_A_304_533#_c_1606_n 0.00216868f $X=0.69 $Y=2.76 $X2=0
+ $Y2=0
cc_887 N_VPWR_c_1480_n N_A_304_533#_c_1606_n 0.0139215f $X=1.91 $Y=3.33 $X2=0
+ $Y2=0
cc_888 N_VPWR_c_1466_n N_A_304_533#_c_1606_n 0.00975953f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_889 N_VPWR_M1007_d N_A_304_533#_c_1607_n 0.0017023f $X=1.935 $Y=2.665 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_1468_n N_A_304_533#_c_1607_n 0.016098f $X=2.075 $Y=2.96 $X2=0
+ $Y2=0
cc_891 N_VPWR_c_1473_n N_A_304_533#_c_1607_n 0.00235807f $X=3.755 $Y=3.33 $X2=0
+ $Y2=0
cc_892 N_VPWR_c_1480_n N_A_304_533#_c_1607_n 0.00235807f $X=1.91 $Y=3.33 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_1466_n N_A_304_533#_c_1607_n 0.00976846f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_894 N_VPWR_c_1473_n N_A_304_533#_c_1674_n 0.0108952f $X=3.755 $Y=3.33 $X2=0
+ $Y2=0
cc_895 N_VPWR_c_1466_n N_A_304_533#_c_1674_n 0.0086247f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_896 N_VPWR_c_1473_n N_A_304_533#_c_1609_n 0.00252511f $X=3.755 $Y=3.33 $X2=0
+ $Y2=0
cc_897 N_VPWR_c_1466_n N_A_304_533#_c_1609_n 0.00448663f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_898 N_VPWR_c_1466_n A_653_533# 0.00168885f $X=10.32 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_899 N_VPWR_c_1466_n N_Q_M1024_d 0.00371702f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_900 N_VPWR_c_1483_n N_Q_c_1684_n 0.0239045f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_901 N_VPWR_c_1466_n N_Q_c_1684_n 0.013335f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_902 Q N_VGND_c_1700_n 0.0309222f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_903 Q N_VGND_c_1707_n 0.0112788f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_904 Q N_VGND_c_1708_n 0.00980826f $X=10.235 $Y=0.47 $X2=0 $Y2=0
