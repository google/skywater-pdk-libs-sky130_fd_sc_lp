* File: sky130_fd_sc_lp__sdfstp_1.pxi.spice
* Created: Wed Sep  2 10:35:37 2020
* 
x_PM_SKY130_FD_SC_LP__SDFSTP_1%SCD N_SCD_M1013_g N_SCD_M1014_g N_SCD_c_268_n
+ N_SCD_c_269_n N_SCD_c_274_n SCD SCD N_SCD_c_271_n
+ PM_SKY130_FD_SC_LP__SDFSTP_1%SCD
x_PM_SKY130_FD_SC_LP__SDFSTP_1%D N_D_M1036_g N_D_M1003_g D D D N_D_c_300_n
+ PM_SKY130_FD_SC_LP__SDFSTP_1%D
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_324_102# N_A_324_102#_M1038_d
+ N_A_324_102#_M1026_d N_A_324_102#_c_335_n N_A_324_102#_M1034_g
+ N_A_324_102#_c_336_n N_A_324_102#_M1009_g N_A_324_102#_c_338_n
+ N_A_324_102#_c_339_n N_A_324_102#_c_340_n N_A_324_102#_c_341_n
+ N_A_324_102#_c_342_n N_A_324_102#_c_346_n N_A_324_102#_c_347_n
+ PM_SKY130_FD_SC_LP__SDFSTP_1%A_324_102#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%SCE N_SCE_M1000_g N_SCE_M1033_g N_SCE_c_417_n
+ N_SCE_c_418_n N_SCE_M1038_g N_SCE_c_420_n N_SCE_c_421_n N_SCE_c_422_n
+ N_SCE_c_423_n N_SCE_M1026_g N_SCE_c_424_n N_SCE_c_425_n N_SCE_c_431_n SCE SCE
+ N_SCE_c_427_n PM_SKY130_FD_SC_LP__SDFSTP_1%SCE
x_PM_SKY130_FD_SC_LP__SDFSTP_1%CLK N_CLK_M1025_g N_CLK_M1027_g CLK CLK CLK
+ N_CLK_c_507_n PM_SKY130_FD_SC_LP__SDFSTP_1%CLK
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_871_47# N_A_871_47#_M1037_d N_A_871_47#_M1016_d
+ N_A_871_47#_M1023_g N_A_871_47#_M1019_g N_A_871_47#_M1001_g
+ N_A_871_47#_M1002_g N_A_871_47#_c_548_n N_A_871_47#_c_555_n
+ N_A_871_47#_c_549_n N_A_871_47#_c_557_n N_A_871_47#_c_550_n
+ N_A_871_47#_c_559_n N_A_871_47#_c_560_n N_A_871_47#_c_561_n
+ N_A_871_47#_c_562_n N_A_871_47#_c_563_n N_A_871_47#_c_564_n
+ N_A_871_47#_c_592_p N_A_871_47#_c_551_n N_A_871_47#_c_565_n
+ N_A_871_47#_c_566_n N_A_871_47#_c_567_n N_A_871_47#_c_568_n
+ N_A_871_47#_c_569_n PM_SKY130_FD_SC_LP__SDFSTP_1%A_871_47#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_1263_31# N_A_1263_31#_M1039_s
+ N_A_1263_31#_M1004_d N_A_1263_31#_c_719_n N_A_1263_31#_M1022_g
+ N_A_1263_31#_c_726_n N_A_1263_31#_M1032_g N_A_1263_31#_c_727_n
+ N_A_1263_31#_c_728_n N_A_1263_31#_c_729_n N_A_1263_31#_c_720_n
+ N_A_1263_31#_c_721_n N_A_1263_31#_c_722_n N_A_1263_31#_c_732_n
+ N_A_1263_31#_c_723_n N_A_1263_31#_c_724_n N_A_1263_31#_c_725_n
+ PM_SKY130_FD_SC_LP__SDFSTP_1%A_1263_31#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_1135_57# N_A_1135_57#_M1018_d
+ N_A_1135_57#_M1023_d N_A_1135_57#_c_809_n N_A_1135_57#_M1004_g
+ N_A_1135_57#_c_797_n N_A_1135_57#_c_798_n N_A_1135_57#_M1039_g
+ N_A_1135_57#_M1029_g N_A_1135_57#_c_799_n N_A_1135_57#_c_800_n
+ N_A_1135_57#_M1007_g N_A_1135_57#_c_812_n N_A_1135_57#_c_908_p
+ N_A_1135_57#_c_801_n N_A_1135_57#_c_802_n N_A_1135_57#_c_803_n
+ N_A_1135_57#_c_804_n N_A_1135_57#_c_805_n N_A_1135_57#_c_806_n
+ N_A_1135_57#_c_807_n N_A_1135_57#_c_808_n
+ PM_SKY130_FD_SC_LP__SDFSTP_1%A_1135_57#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%SET_B N_SET_B_M1020_g N_SET_B_M1021_g
+ N_SET_B_M1012_g N_SET_B_c_913_n N_SET_B_M1035_g N_SET_B_c_914_n
+ N_SET_B_c_915_n N_SET_B_c_916_n N_SET_B_c_925_n N_SET_B_c_917_n
+ N_SET_B_c_918_n N_SET_B_c_919_n SET_B SET_B SET_B SET_B SET_B SET_B
+ N_SET_B_c_920_n N_SET_B_c_921_n PM_SKY130_FD_SC_LP__SDFSTP_1%SET_B
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_702_47# N_A_702_47#_M1025_s N_A_702_47#_M1027_s
+ N_A_702_47#_c_1013_n N_A_702_47#_M1037_g N_A_702_47#_c_1014_n
+ N_A_702_47#_M1016_g N_A_702_47#_c_1015_n N_A_702_47#_c_1027_n
+ N_A_702_47#_c_1028_n N_A_702_47#_c_1029_n N_A_702_47#_c_1030_n
+ N_A_702_47#_M1018_g N_A_702_47#_M1028_g N_A_702_47#_c_1032_n
+ N_A_702_47#_c_1033_n N_A_702_47#_M1017_g N_A_702_47#_c_1017_n
+ N_A_702_47#_c_1018_n N_A_702_47#_M1006_g N_A_702_47#_c_1020_n
+ N_A_702_47#_c_1037_n N_A_702_47#_c_1021_n N_A_702_47#_c_1022_n
+ N_A_702_47#_c_1038_n N_A_702_47#_c_1039_n N_A_702_47#_c_1023_n
+ N_A_702_47#_c_1041_n N_A_702_47#_c_1024_n N_A_702_47#_c_1025_n
+ N_A_702_47#_c_1043_n PM_SKY130_FD_SC_LP__SDFSTP_1%A_702_47#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_2158_231# N_A_2158_231#_M1031_d
+ N_A_2158_231#_M1011_d N_A_2158_231#_M1010_g N_A_2158_231#_M1024_g
+ N_A_2158_231#_c_1194_n N_A_2158_231#_c_1195_n N_A_2158_231#_c_1196_n
+ N_A_2158_231#_c_1197_n N_A_2158_231#_c_1198_n N_A_2158_231#_c_1199_n
+ N_A_2158_231#_c_1200_n PM_SKY130_FD_SC_LP__SDFSTP_1%A_2158_231#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_1912_463# N_A_1912_463#_M1002_d
+ N_A_1912_463#_M1001_d N_A_1912_463#_M1035_d N_A_1912_463#_M1031_g
+ N_A_1912_463#_M1011_g N_A_1912_463#_c_1262_n N_A_1912_463#_M1005_g
+ N_A_1912_463#_c_1269_n N_A_1912_463#_M1008_g N_A_1912_463#_c_1264_n
+ N_A_1912_463#_c_1271_n N_A_1912_463#_c_1265_n N_A_1912_463#_c_1273_n
+ N_A_1912_463#_c_1266_n N_A_1912_463#_c_1275_n N_A_1912_463#_c_1276_n
+ N_A_1912_463#_c_1277_n N_A_1912_463#_c_1298_n N_A_1912_463#_c_1278_n
+ N_A_1912_463#_c_1279_n PM_SKY130_FD_SC_LP__SDFSTP_1%A_1912_463#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_2598_153# N_A_2598_153#_M1005_s
+ N_A_2598_153#_M1008_s N_A_2598_153#_M1015_g N_A_2598_153#_M1030_g
+ N_A_2598_153#_c_1372_n N_A_2598_153#_c_1378_n N_A_2598_153#_c_1373_n
+ N_A_2598_153#_c_1374_n N_A_2598_153#_c_1375_n N_A_2598_153#_c_1376_n
+ PM_SKY130_FD_SC_LP__SDFSTP_1%A_2598_153#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_27_408# N_A_27_408#_M1013_s N_A_27_408#_M1009_d
+ N_A_27_408#_c_1413_n N_A_27_408#_c_1414_n N_A_27_408#_c_1415_n
+ N_A_27_408#_c_1416_n PM_SKY130_FD_SC_LP__SDFSTP_1%A_27_408#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%VPWR N_VPWR_M1013_d N_VPWR_M1026_s N_VPWR_M1027_d
+ N_VPWR_M1032_d N_VPWR_M1020_d N_VPWR_M1010_d N_VPWR_M1011_s N_VPWR_M1008_d
+ N_VPWR_c_1446_n N_VPWR_c_1447_n N_VPWR_c_1448_n N_VPWR_c_1449_n
+ N_VPWR_c_1450_n N_VPWR_c_1451_n N_VPWR_c_1452_n N_VPWR_c_1453_n
+ N_VPWR_c_1454_n N_VPWR_c_1455_n N_VPWR_c_1456_n N_VPWR_c_1457_n
+ N_VPWR_c_1458_n VPWR N_VPWR_c_1459_n N_VPWR_c_1460_n N_VPWR_c_1461_n
+ N_VPWR_c_1462_n N_VPWR_c_1463_n N_VPWR_c_1464_n N_VPWR_c_1445_n
+ N_VPWR_c_1466_n N_VPWR_c_1467_n N_VPWR_c_1468_n N_VPWR_c_1469_n
+ N_VPWR_c_1470_n N_VPWR_c_1471_n PM_SKY130_FD_SC_LP__SDFSTP_1%VPWR
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_196_128# N_A_196_128#_M1000_d
+ N_A_196_128#_M1018_s N_A_196_128#_M1036_d N_A_196_128#_M1023_s
+ N_A_196_128#_c_1622_n N_A_196_128#_c_1609_n N_A_196_128#_c_1610_n
+ N_A_196_128#_c_1614_n N_A_196_128#_c_1611_n N_A_196_128#_c_1649_n
+ N_A_196_128#_c_1663_n N_A_196_128#_c_1616_n N_A_196_128#_c_1617_n
+ N_A_196_128#_c_1654_n N_A_196_128#_c_1667_n N_A_196_128#_c_1655_n
+ N_A_196_128#_c_1618_n N_A_196_128#_c_1612_n N_A_196_128#_c_1720_n
+ N_A_196_128#_c_1746_n N_A_196_128#_c_1620_n N_A_196_128#_c_1613_n
+ N_A_196_128#_c_1621_n PM_SKY130_FD_SC_LP__SDFSTP_1%A_196_128#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_1703_379# N_A_1703_379#_M1029_d
+ N_A_1703_379#_M1017_d N_A_1703_379#_c_1758_n N_A_1703_379#_c_1759_n
+ N_A_1703_379#_c_1760_n PM_SKY130_FD_SC_LP__SDFSTP_1%A_1703_379#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%A_1810_463# N_A_1810_463#_M1001_s
+ N_A_1810_463#_M1010_s N_A_1810_463#_c_1791_n N_A_1810_463#_c_1792_n
+ N_A_1810_463#_c_1793_n PM_SKY130_FD_SC_LP__SDFSTP_1%A_1810_463#
x_PM_SKY130_FD_SC_LP__SDFSTP_1%Q N_Q_M1015_d N_Q_M1030_d Q Q Q Q Q Q Q
+ N_Q_c_1817_n Q Q PM_SKY130_FD_SC_LP__SDFSTP_1%Q
x_PM_SKY130_FD_SC_LP__SDFSTP_1%VGND N_VGND_M1014_s N_VGND_M1034_d N_VGND_M1025_d
+ N_VGND_M1022_d N_VGND_M1021_d N_VGND_M1012_d N_VGND_M1005_d N_VGND_c_1833_n
+ N_VGND_c_1834_n N_VGND_c_1835_n N_VGND_c_1836_n N_VGND_c_1837_n
+ N_VGND_c_1838_n N_VGND_c_1911_n N_VGND_c_1913_n N_VGND_c_1839_n
+ N_VGND_c_1840_n N_VGND_c_1841_n N_VGND_c_1842_n N_VGND_c_1843_n
+ N_VGND_c_1844_n N_VGND_c_1845_n N_VGND_c_1846_n VGND N_VGND_c_1847_n
+ N_VGND_c_1848_n N_VGND_c_1849_n N_VGND_c_1850_n N_VGND_c_1851_n
+ N_VGND_c_1852_n N_VGND_c_1853_n N_VGND_c_1854_n
+ PM_SKY130_FD_SC_LP__SDFSTP_1%VGND
cc_1 VNB N_SCD_c_268_n 0.0211419f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.17
cc_2 VNB N_SCD_c_269_n 0.0256058f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.675
cc_3 VNB SCD 0.0221048f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_SCD_c_271_n 0.0183831f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_5 VNB N_D_M1003_g 0.0316516f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.85
cc_6 VNB D 0.00474758f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.84
cc_7 VNB N_D_c_300_n 0.0113905f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_8 VNB N_A_324_102#_c_335_n 0.0144542f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.85
cc_9 VNB N_A_324_102#_c_336_n 0.0278018f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.675
cc_10 VNB N_A_324_102#_M1009_g 0.00405205f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A_324_102#_c_338_n 0.0487022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_324_102#_c_339_n 0.00929145f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.335
cc_13 VNB N_A_324_102#_c_340_n 0.00234456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_324_102#_c_341_n 0.0426782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_324_102#_c_342_n 0.00968382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_M1000_g 0.0560989f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.36
cc_17 VNB N_SCE_c_417_n 0.0803146f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.85
cc_18 VNB N_SCE_c_418_n 0.0124764f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_19 VNB N_SCE_M1038_g 0.0327551f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.84
cc_20 VNB N_SCE_c_420_n 0.0242052f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_SCE_c_421_n 0.0148024f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_22 VNB N_SCE_c_422_n 0.0351944f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_23 VNB N_SCE_c_423_n 0.00778217f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_24 VNB N_SCE_c_424_n 0.0416244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_SCE_c_425_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB SCE 0.0167958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_SCE_c_427_n 0.0460925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_CLK_M1025_g 0.0417686f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.36
cc_29 VNB CLK 0.0129694f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.17
cc_30 VNB N_CLK_c_507_n 0.049303f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_31 VNB N_A_871_47#_M1019_g 0.05666f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_A_871_47#_M1002_g 0.0362154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_871_47#_c_548_n 0.0133387f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.665
cc_34 VNB N_A_871_47#_c_549_n 0.00740276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_871_47#_c_550_n 0.0438757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_871_47#_c_551_n 0.00808202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1263_31#_c_719_n 0.0191125f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.85
cc_38 VNB N_A_1263_31#_c_720_n 0.00771554f $X=-0.19 $Y=-0.245 $X2=0.387
+ $Y2=1.295
cc_39 VNB N_A_1263_31#_c_721_n 0.00397216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1263_31#_c_722_n 0.0129209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1263_31#_c_723_n 0.0063772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1263_31#_c_724_n 0.0469123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1263_31#_c_725_n 0.0221182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1135_57#_c_797_n 0.00877269f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.84
cc_45 VNB N_A_1135_57#_c_798_n 0.0204386f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_46 VNB N_A_1135_57#_c_799_n 0.0386433f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.295
cc_47 VNB N_A_1135_57#_c_800_n 0.0176987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1135_57#_c_801_n 0.0101211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1135_57#_c_802_n 0.0016324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1135_57#_c_803_n 0.0388521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1135_57#_c_804_n 6.70291e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1135_57#_c_805_n 0.00173893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1135_57#_c_806_n 0.0053428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1135_57#_c_807_n 0.0375281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1135_57#_c_808_n 0.0317288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_SET_B_M1021_g 0.0419588f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_57 VNB N_SET_B_c_913_n 0.00630692f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_58 VNB N_SET_B_c_914_n 0.00893652f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_59 VNB N_SET_B_c_915_n 0.0177913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_SET_B_c_916_n 0.00481352f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.335
cc_61 VNB N_SET_B_c_917_n 0.00943506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_SET_B_c_918_n 0.0131039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_SET_B_c_919_n 0.0477077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_SET_B_c_920_n 0.0475623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_SET_B_c_921_n 0.0128879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_702_47#_c_1013_n 0.0202875f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.85
cc_67 VNB N_A_702_47#_c_1014_n 0.0144089f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.84
cc_68 VNB N_A_702_47#_c_1015_n 0.057814f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_69 VNB N_A_702_47#_M1018_g 0.0402028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_702_47#_c_1017_n 0.0127031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_702_47#_c_1018_n 0.00492455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_702_47#_M1006_g 0.042224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_702_47#_c_1020_n 6.40364e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_702_47#_c_1021_n 0.0330103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_702_47#_c_1022_n 0.0116756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_702_47#_c_1023_n 0.00980583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_702_47#_c_1024_n 0.0272951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_702_47#_c_1025_n 0.00474514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_2158_231#_M1010_g 0.00854796f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.17
cc_80 VNB N_A_2158_231#_c_1194_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_2158_231#_c_1195_n 0.0338522f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.335
cc_82 VNB N_A_2158_231#_c_1196_n 0.0143359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2158_231#_c_1197_n 0.0225699f $X=-0.19 $Y=-0.245 $X2=0.387
+ $Y2=1.665
cc_84 VNB N_A_2158_231#_c_1198_n 0.00328738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2158_231#_c_1199_n 0.00334136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2158_231#_c_1200_n 0.0178249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1912_463#_M1031_g 0.0495488f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_88 VNB N_A_1912_463#_c_1262_n 0.0299001f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.335
cc_89 VNB N_A_1912_463#_M1005_g 0.0374099f $X=-0.19 $Y=-0.245 $X2=0.387
+ $Y2=1.335
cc_90 VNB N_A_1912_463#_c_1264_n 0.015616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1912_463#_c_1265_n 0.00295807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1912_463#_c_1266_n 0.0144958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2598_153#_M1030_g 0.00178937f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_94 VNB N_A_2598_153#_c_1372_n 0.0103842f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.335
cc_95 VNB N_A_2598_153#_c_1373_n 0.00474618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2598_153#_c_1374_n 0.0348188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2598_153#_c_1375_n 0.00416316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2598_153#_c_1376_n 0.0220424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VPWR_c_1445_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_196_128#_c_1609_n 0.0249931f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.335
cc_101 VNB N_A_196_128#_c_1610_n 0.00267042f $X=-0.19 $Y=-0.245 $X2=0.455
+ $Y2=1.335
cc_102 VNB N_A_196_128#_c_1611_n 0.00231152f $X=-0.19 $Y=-0.245 $X2=0.387
+ $Y2=1.335
cc_103 VNB N_A_196_128#_c_1612_n 0.0162629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_196_128#_c_1613_n 0.0031696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB Q 0.00838398f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.335
cc_106 VNB Q 0.0268028f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.17
cc_107 VNB N_Q_c_1817_n 0.0294554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1833_n 0.0138117f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.335
cc_109 VNB N_VGND_c_1834_n 0.0406488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1835_n 0.0130049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1836_n 0.0051258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1837_n 0.0164669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1838_n 0.0165299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1839_n 0.0317542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1840_n 0.0234444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1841_n 0.037444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1842_n 0.00374536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1843_n 0.0215963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1844_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1845_n 0.0486805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1846_n 0.00682834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1847_n 0.0500086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1848_n 0.0579422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1849_n 0.0964865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1850_n 0.0194853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1851_n 0.797091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1852_n 0.00478335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1853_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1854_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VPB N_SCD_M1013_g 0.0304525f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.36
cc_131 VPB N_SCD_c_269_n 0.00152567f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.675
cc_132 VPB N_SCD_c_274_n 0.0183415f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.84
cc_133 VPB SCD 0.0101243f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_134 VPB N_D_M1036_g 0.0214552f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.36
cc_135 VPB D 0.0109836f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.84
cc_136 VPB N_D_c_300_n 0.0160516f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.335
cc_137 VPB N_A_324_102#_M1009_g 0.0393199f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_138 VPB N_A_324_102#_c_341_n 0.0194123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_324_102#_c_342_n 0.00287075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_324_102#_c_346_n 0.00447336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_324_102#_c_347_n 0.0117367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_SCE_M1000_g 0.0293977f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.36
cc_143 VPB N_SCE_M1026_g 0.0301397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_SCE_c_424_n 0.019375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_SCE_c_431_n 0.0279772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_CLK_M1027_g 0.0475772f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.85
cc_147 VPB CLK 0.00355841f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.17
cc_148 VPB N_CLK_c_507_n 0.0227548f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.335
cc_149 VPB N_A_871_47#_M1023_g 0.0395401f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.17
cc_150 VPB N_A_871_47#_M1001_g 0.0252188f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.335
cc_151 VPB N_A_871_47#_M1002_g 0.0092113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_871_47#_c_555_n 0.0198491f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_871_47#_c_549_n 0.00217742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_871_47#_c_557_n 0.00178211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_871_47#_c_550_n 0.0574543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_871_47#_c_559_n 0.00292889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_871_47#_c_560_n 0.00966818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_871_47#_c_561_n 0.00515334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_871_47#_c_562_n 0.00982051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_871_47#_c_563_n 0.00240995f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_871_47#_c_564_n 0.00424637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_871_47#_c_565_n 0.00259585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_871_47#_c_566_n 0.00376813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_871_47#_c_567_n 0.00439691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_871_47#_c_568_n 0.0225356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_871_47#_c_569_n 0.0523733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_1263_31#_c_726_n 0.016082f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.675
cc_168 VPB N_A_1263_31#_c_727_n 0.0228567f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_169 VPB N_A_1263_31#_c_728_n 0.00865833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_1263_31#_c_729_n 0.01267f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.335
cc_171 VPB N_A_1263_31#_c_721_n 0.00469569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_1263_31#_c_722_n 0.0153524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_1263_31#_c_732_n 0.00390942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_1135_57#_c_809_n 0.0163049f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.85
cc_175 VPB N_A_1135_57#_c_797_n 0.0181162f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.84
cc_176 VPB N_A_1135_57#_M1029_g 0.0252419f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.335
cc_177 VPB N_A_1135_57#_c_812_n 0.0129648f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_1135_57#_c_802_n 0.00946738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_1135_57#_c_808_n 0.00962897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_SET_B_M1020_g 0.0332582f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.36
cc_181 VPB N_SET_B_M1035_g 0.0455276f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.335
cc_182 VPB N_SET_B_c_914_n 0.0351966f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.335
cc_183 VPB N_SET_B_c_925_n 2.34762e-19 $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.665
cc_184 VPB N_SET_B_c_917_n 0.00614018f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_SET_B_c_918_n 0.0163468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_702_47#_M1016_g 0.0189527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_702_47#_c_1027_n 0.0243938f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.335
cc_188 VPB N_A_702_47#_c_1028_n 0.0453444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_702_47#_c_1029_n 0.0499745f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.335
cc_190 VPB N_A_702_47#_c_1030_n 0.0106266f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.665
cc_191 VPB N_A_702_47#_M1028_g 0.0307522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_702_47#_c_1032_n 0.327974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_702_47#_c_1033_n 0.0135809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_702_47#_c_1017_n 0.012697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_702_47#_c_1018_n 0.00418405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_702_47#_c_1020_n 0.0103727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_702_47#_c_1037_n 0.0696185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_702_47#_c_1038_n 0.00972873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_702_47#_c_1039_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_702_47#_c_1023_n 0.00441066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_702_47#_c_1041_n 0.0121189f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_702_47#_c_1024_n 0.0329384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_702_47#_c_1043_n 0.00996663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_2158_231#_M1010_g 0.0507518f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.17
cc_205 VPB N_A_2158_231#_c_1198_n 0.020452f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1912_463#_M1011_g 0.0266555f $X=-0.19 $Y=1.655 $X2=0.455
+ $Y2=1.335
cc_207 VPB N_A_1912_463#_c_1262_n 0.0269668f $X=-0.19 $Y=1.655 $X2=0.455
+ $Y2=1.335
cc_208 VPB N_A_1912_463#_c_1269_n 0.0208066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_1912_463#_c_1264_n 0.0115084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_1912_463#_c_1271_n 0.0222698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_1912_463#_c_1265_n 0.00298481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_1912_463#_c_1273_n 0.00151515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_1912_463#_c_1266_n 0.00477913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_1912_463#_c_1275_n 0.0168547f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_1912_463#_c_1276_n 0.00487408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_1912_463#_c_1277_n 0.0177217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_1912_463#_c_1278_n 0.0300523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_1912_463#_c_1279_n 0.00460347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_2598_153#_M1030_g 0.0261157f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_220 VPB N_A_2598_153#_c_1378_n 0.0141385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_27_408#_c_1413_n 0.0239793f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.17
cc_222 VPB N_A_27_408#_c_1414_n 0.0127708f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.84
cc_223 VPB N_A_27_408#_c_1415_n 0.0115399f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_224 VPB N_A_27_408#_c_1416_n 0.00600994f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_225 VPB N_VPWR_c_1446_n 0.0292513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1447_n 0.0177447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1448_n 0.00151893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1449_n 0.0444784f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1450_n 0.00713462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1451_n 0.0178489f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1452_n 0.0126678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1453_n 0.0178977f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1454_n 0.0266097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1455_n 0.0300858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1456_n 0.00450185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1457_n 0.0711919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1458_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1459_n 0.0186462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1460_n 0.0443005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1461_n 0.035709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1462_n 0.019647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1463_n 0.0330628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1464_n 0.0155059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1445_n 0.137015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1466_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1467_n 0.00631764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1468_n 0.00485096f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1469_n 0.00370284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1470_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1471_n 0.00728342f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_196_128#_c_1614_n 0.0124407f $X=-0.19 $Y=1.655 $X2=0.387
+ $Y2=1.295
cc_252 VPB N_A_196_128#_c_1611_n 0.0198756f $X=-0.19 $Y=1.655 $X2=0.387
+ $Y2=1.335
cc_253 VPB N_A_196_128#_c_1616_n 0.0155967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_196_128#_c_1617_n 0.00126396f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_196_128#_c_1618_n 0.00568192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_A_196_128#_c_1612_n 0.0118622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_196_128#_c_1620_n 0.00176303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_196_128#_c_1621_n 0.00916869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_1703_379#_c_1758_n 0.0096613f $X=-0.19 $Y=1.655 $X2=0.455
+ $Y2=1.675
cc_260 VPB N_A_1703_379#_c_1759_n 0.00402302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_1703_379#_c_1760_n 0.0124554f $X=-0.19 $Y=1.655 $X2=0.455
+ $Y2=1.335
cc_262 VPB N_A_1810_463#_c_1791_n 0.0219579f $X=-0.19 $Y=1.655 $X2=0.545
+ $Y2=0.85
cc_263 VPB N_A_1810_463#_c_1792_n 0.00334867f $X=-0.19 $Y=1.655 $X2=0.455
+ $Y2=1.84
cc_264 VPB N_A_1810_463#_c_1793_n 0.0105348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB Q 0.0102656f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.17
cc_266 VPB Q 0.00536733f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.84
cc_267 VPB Q 0.0419152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 SCD D 0.0141279f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_269 N_SCD_M1013_g N_SCE_M1000_g 0.0278965f $X=0.475 $Y=2.36 $X2=0 $Y2=0
cc_270 N_SCD_c_268_n N_SCE_M1000_g 0.079482f $X=0.455 $Y=1.17 $X2=0 $Y2=0
cc_271 SCD N_SCE_M1000_g 0.00284335f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_272 N_SCD_M1013_g N_A_27_408#_c_1413_n 4.68635e-19 $X=0.475 $Y=2.36 $X2=0
+ $Y2=0
cc_273 N_SCD_M1013_g N_A_27_408#_c_1414_n 0.0132878f $X=0.475 $Y=2.36 $X2=0
+ $Y2=0
cc_274 N_SCD_c_274_n N_A_27_408#_c_1414_n 5.47375e-19 $X=0.455 $Y=1.84 $X2=0
+ $Y2=0
cc_275 SCD N_A_27_408#_c_1414_n 0.0176801f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_276 N_SCD_c_274_n N_A_27_408#_c_1415_n 7.79991e-19 $X=0.455 $Y=1.84 $X2=0
+ $Y2=0
cc_277 SCD N_A_27_408#_c_1415_n 0.0214714f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_278 N_SCD_M1013_g N_VPWR_c_1446_n 0.00324707f $X=0.475 $Y=2.36 $X2=0 $Y2=0
cc_279 N_SCD_M1013_g N_VPWR_c_1459_n 0.00402388f $X=0.475 $Y=2.36 $X2=0 $Y2=0
cc_280 N_SCD_M1013_g N_VPWR_c_1445_n 0.00462577f $X=0.475 $Y=2.36 $X2=0 $Y2=0
cc_281 N_SCD_c_268_n N_A_196_128#_c_1622_n 0.0017653f $X=0.455 $Y=1.17 $X2=0
+ $Y2=0
cc_282 SCD N_A_196_128#_c_1622_n 8.73176e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_283 SCD N_A_196_128#_c_1610_n 0.00803839f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_284 N_SCD_c_271_n N_A_196_128#_c_1610_n 4.87567e-19 $X=0.455 $Y=1.335 $X2=0
+ $Y2=0
cc_285 N_SCD_c_268_n N_VGND_c_1834_n 0.0118713f $X=0.455 $Y=1.17 $X2=0 $Y2=0
cc_286 SCD N_VGND_c_1834_n 0.0265885f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_287 N_SCD_c_271_n N_VGND_c_1834_n 0.00123586f $X=0.455 $Y=1.335 $X2=0 $Y2=0
cc_288 N_SCD_c_268_n N_VGND_c_1841_n 0.00338717f $X=0.455 $Y=1.17 $X2=0 $Y2=0
cc_289 N_SCD_c_268_n N_VGND_c_1851_n 0.00390857f $X=0.455 $Y=1.17 $X2=0 $Y2=0
cc_290 N_D_M1003_g N_A_324_102#_c_335_n 0.0485481f $X=1.335 $Y=0.85 $X2=0 $Y2=0
cc_291 N_D_M1003_g N_A_324_102#_c_336_n 0.00975707f $X=1.335 $Y=0.85 $X2=0 $Y2=0
cc_292 D N_A_324_102#_c_336_n 0.00396812f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_293 N_D_c_300_n N_A_324_102#_c_336_n 0.0214495f $X=1.355 $Y=1.695 $X2=0 $Y2=0
cc_294 N_D_M1036_g N_A_324_102#_M1009_g 0.0190663f $X=1.265 $Y=2.36 $X2=0 $Y2=0
cc_295 D N_A_324_102#_M1009_g 0.0135132f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_296 D N_A_324_102#_c_338_n 0.0113712f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_297 N_D_M1003_g N_SCE_M1000_g 0.0296208f $X=1.335 $Y=0.85 $X2=0 $Y2=0
cc_298 D N_SCE_M1000_g 0.00365298f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_299 N_D_c_300_n N_SCE_M1000_g 0.0785416f $X=1.355 $Y=1.695 $X2=0 $Y2=0
cc_300 N_D_M1003_g N_SCE_c_417_n 0.00899345f $X=1.335 $Y=0.85 $X2=0 $Y2=0
cc_301 N_D_M1036_g N_A_27_408#_c_1414_n 0.0148555f $X=1.265 $Y=2.36 $X2=0 $Y2=0
cc_302 D N_A_27_408#_c_1414_n 0.0633776f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_303 N_D_c_300_n N_A_27_408#_c_1414_n 0.00441334f $X=1.355 $Y=1.695 $X2=0
+ $Y2=0
cc_304 N_D_M1036_g N_A_27_408#_c_1416_n 5.34187e-19 $X=1.265 $Y=2.36 $X2=0 $Y2=0
cc_305 D N_A_27_408#_c_1416_n 0.026708f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_306 N_D_M1036_g N_VPWR_c_1446_n 0.00166858f $X=1.265 $Y=2.36 $X2=0 $Y2=0
cc_307 N_D_M1036_g N_VPWR_c_1460_n 0.00402388f $X=1.265 $Y=2.36 $X2=0 $Y2=0
cc_308 N_D_M1036_g N_VPWR_c_1445_n 0.00462577f $X=1.265 $Y=2.36 $X2=0 $Y2=0
cc_309 N_D_M1003_g N_A_196_128#_c_1622_n 0.0103392f $X=1.335 $Y=0.85 $X2=0 $Y2=0
cc_310 N_D_M1003_g N_A_196_128#_c_1609_n 0.0108062f $X=1.335 $Y=0.85 $X2=0 $Y2=0
cc_311 D N_A_196_128#_c_1609_n 0.0723116f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_312 N_D_c_300_n N_A_196_128#_c_1609_n 0.00246626f $X=1.355 $Y=1.695 $X2=0
+ $Y2=0
cc_313 N_D_M1003_g N_A_196_128#_c_1610_n 0.00273135f $X=1.335 $Y=0.85 $X2=0
+ $Y2=0
cc_314 D N_A_196_128#_c_1610_n 0.0232629f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_315 N_D_c_300_n N_A_196_128#_c_1610_n 0.00190367f $X=1.355 $Y=1.695 $X2=0
+ $Y2=0
cc_316 D N_A_196_128#_c_1614_n 0.00234661f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_317 D N_A_196_128#_c_1611_n 0.0256074f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_318 N_D_M1003_g N_VGND_c_1835_n 0.00178013f $X=1.335 $Y=0.85 $X2=0 $Y2=0
cc_319 N_D_M1003_g N_VGND_c_1851_n 9.32216e-19 $X=1.335 $Y=0.85 $X2=0 $Y2=0
cc_320 N_A_324_102#_c_335_n N_SCE_c_417_n 0.00896847f $X=1.695 $Y=1.17 $X2=0
+ $Y2=0
cc_321 N_A_324_102#_c_335_n N_SCE_M1038_g 0.0104466f $X=1.695 $Y=1.17 $X2=0
+ $Y2=0
cc_322 N_A_324_102#_c_336_n N_SCE_M1038_g 0.0013763f $X=1.805 $Y=1.58 $X2=0
+ $Y2=0
cc_323 N_A_324_102#_c_338_n N_SCE_M1038_g 0.00737308f $X=2.695 $Y=1.505 $X2=0
+ $Y2=0
cc_324 N_A_324_102#_c_339_n N_SCE_M1038_g 0.00302799f $X=2.765 $Y=0.915 $X2=0
+ $Y2=0
cc_325 N_A_324_102#_c_340_n N_SCE_M1038_g 0.00234937f $X=2.86 $Y=1.285 $X2=0
+ $Y2=0
cc_326 N_A_324_102#_c_341_n N_SCE_M1038_g 0.00206077f $X=2.86 $Y=1.285 $X2=0
+ $Y2=0
cc_327 N_A_324_102#_c_339_n N_SCE_c_420_n 0.00270245f $X=2.765 $Y=0.915 $X2=0
+ $Y2=0
cc_328 N_A_324_102#_c_339_n N_SCE_c_422_n 0.00351194f $X=2.765 $Y=0.915 $X2=0
+ $Y2=0
cc_329 N_A_324_102#_c_339_n N_SCE_c_423_n 0.00605565f $X=2.765 $Y=0.915 $X2=0
+ $Y2=0
cc_330 N_A_324_102#_c_341_n N_SCE_c_423_n 0.0126942f $X=2.86 $Y=1.285 $X2=0
+ $Y2=0
cc_331 N_A_324_102#_c_347_n N_SCE_M1026_g 0.00637001f $X=3.32 $Y=2.56 $X2=0
+ $Y2=0
cc_332 N_A_324_102#_c_339_n N_SCE_c_424_n 0.00117792f $X=2.765 $Y=0.915 $X2=0
+ $Y2=0
cc_333 N_A_324_102#_c_340_n N_SCE_c_424_n 0.00414674f $X=2.86 $Y=1.285 $X2=0
+ $Y2=0
cc_334 N_A_324_102#_c_341_n N_SCE_c_424_n 0.0361203f $X=2.86 $Y=1.285 $X2=0
+ $Y2=0
cc_335 N_A_324_102#_c_342_n N_SCE_c_424_n 0.0128447f $X=3.225 $Y=1.705 $X2=0
+ $Y2=0
cc_336 N_A_324_102#_c_347_n N_SCE_c_424_n 0.0078591f $X=3.32 $Y=2.56 $X2=0 $Y2=0
cc_337 N_A_324_102#_c_342_n N_SCE_c_431_n 0.00694079f $X=3.225 $Y=1.705 $X2=0
+ $Y2=0
cc_338 N_A_324_102#_c_347_n N_SCE_c_431_n 0.0125401f $X=3.32 $Y=2.56 $X2=0 $Y2=0
cc_339 N_A_324_102#_c_339_n SCE 0.0472747f $X=2.765 $Y=0.915 $X2=0 $Y2=0
cc_340 N_A_324_102#_c_341_n SCE 2.55228e-19 $X=2.86 $Y=1.285 $X2=0 $Y2=0
cc_341 N_A_324_102#_c_339_n N_SCE_c_427_n 7.32916e-19 $X=2.765 $Y=0.915 $X2=0
+ $Y2=0
cc_342 N_A_324_102#_c_341_n N_SCE_c_427_n 0.0013414f $X=2.86 $Y=1.285 $X2=0
+ $Y2=0
cc_343 N_A_324_102#_c_347_n N_CLK_M1027_g 0.00521918f $X=3.32 $Y=2.56 $X2=0
+ $Y2=0
cc_344 N_A_324_102#_c_342_n N_CLK_c_507_n 4.86603e-19 $X=3.225 $Y=1.705 $X2=0
+ $Y2=0
cc_345 N_A_324_102#_c_339_n N_A_702_47#_c_1023_n 0.00713163f $X=2.765 $Y=0.915
+ $X2=0 $Y2=0
cc_346 N_A_324_102#_c_340_n N_A_702_47#_c_1023_n 0.017639f $X=2.86 $Y=1.285
+ $X2=0 $Y2=0
cc_347 N_A_324_102#_c_342_n N_A_702_47#_c_1023_n 0.0143463f $X=3.225 $Y=1.705
+ $X2=0 $Y2=0
cc_348 N_A_324_102#_c_347_n N_A_702_47#_c_1023_n 0.0156751f $X=3.32 $Y=2.56
+ $X2=0 $Y2=0
cc_349 N_A_324_102#_c_347_n N_A_702_47#_c_1043_n 0.0268612f $X=3.32 $Y=2.56
+ $X2=0 $Y2=0
cc_350 N_A_324_102#_M1009_g N_A_27_408#_c_1414_n 0.00893864f $X=1.805 $Y=2.36
+ $X2=0 $Y2=0
cc_351 N_A_324_102#_M1009_g N_A_27_408#_c_1416_n 0.00413415f $X=1.805 $Y=2.36
+ $X2=0 $Y2=0
cc_352 N_A_324_102#_c_338_n N_A_27_408#_c_1416_n 8.86038e-19 $X=2.695 $Y=1.505
+ $X2=0 $Y2=0
cc_353 N_A_324_102#_M1009_g N_VPWR_c_1460_n 0.00314569f $X=1.805 $Y=2.36 $X2=0
+ $Y2=0
cc_354 N_A_324_102#_M1009_g N_VPWR_c_1445_n 0.00462577f $X=1.805 $Y=2.36 $X2=0
+ $Y2=0
cc_355 N_A_324_102#_c_335_n N_A_196_128#_c_1622_n 0.00177595f $X=1.695 $Y=1.17
+ $X2=0 $Y2=0
cc_356 N_A_324_102#_c_336_n N_A_196_128#_c_1609_n 0.0195666f $X=1.805 $Y=1.58
+ $X2=0 $Y2=0
cc_357 N_A_324_102#_c_338_n N_A_196_128#_c_1609_n 0.0103151f $X=2.695 $Y=1.505
+ $X2=0 $Y2=0
cc_358 N_A_324_102#_c_339_n N_A_196_128#_c_1609_n 0.0279632f $X=2.765 $Y=0.915
+ $X2=0 $Y2=0
cc_359 N_A_324_102#_c_340_n N_A_196_128#_c_1609_n 0.0141053f $X=2.86 $Y=1.285
+ $X2=0 $Y2=0
cc_360 N_A_324_102#_c_341_n N_A_196_128#_c_1609_n 0.00431153f $X=2.86 $Y=1.285
+ $X2=0 $Y2=0
cc_361 N_A_324_102#_M1009_g N_A_196_128#_c_1614_n 0.0125325f $X=1.805 $Y=2.36
+ $X2=0 $Y2=0
cc_362 N_A_324_102#_c_336_n N_A_196_128#_c_1611_n 0.00160854f $X=1.805 $Y=1.58
+ $X2=0 $Y2=0
cc_363 N_A_324_102#_M1009_g N_A_196_128#_c_1611_n 0.00794056f $X=1.805 $Y=2.36
+ $X2=0 $Y2=0
cc_364 N_A_324_102#_c_338_n N_A_196_128#_c_1611_n 0.0167715f $X=2.695 $Y=1.505
+ $X2=0 $Y2=0
cc_365 N_A_324_102#_c_340_n N_A_196_128#_c_1611_n 0.0185546f $X=2.86 $Y=1.285
+ $X2=0 $Y2=0
cc_366 N_A_324_102#_c_341_n N_A_196_128#_c_1611_n 0.00681433f $X=2.86 $Y=1.285
+ $X2=0 $Y2=0
cc_367 N_A_324_102#_c_346_n N_A_196_128#_c_1611_n 0.0135765f $X=3.025 $Y=1.705
+ $X2=0 $Y2=0
cc_368 N_A_324_102#_c_347_n N_A_196_128#_c_1611_n 0.0188369f $X=3.32 $Y=2.56
+ $X2=0 $Y2=0
cc_369 N_A_324_102#_c_341_n N_A_196_128#_c_1649_n 0.00294899f $X=2.86 $Y=1.285
+ $X2=0 $Y2=0
cc_370 N_A_324_102#_c_342_n N_A_196_128#_c_1649_n 7.52857e-19 $X=3.225 $Y=1.705
+ $X2=0 $Y2=0
cc_371 N_A_324_102#_c_346_n N_A_196_128#_c_1649_n 0.00650601f $X=3.025 $Y=1.705
+ $X2=0 $Y2=0
cc_372 N_A_324_102#_M1026_d N_A_196_128#_c_1616_n 0.00307724f $X=3.18 $Y=2.405
+ $X2=0 $Y2=0
cc_373 N_A_324_102#_c_347_n N_A_196_128#_c_1616_n 0.015408f $X=3.32 $Y=2.56
+ $X2=0 $Y2=0
cc_374 N_A_324_102#_c_347_n N_A_196_128#_c_1654_n 0.00214508f $X=3.32 $Y=2.56
+ $X2=0 $Y2=0
cc_375 N_A_324_102#_c_347_n N_A_196_128#_c_1655_n 0.00667989f $X=3.32 $Y=2.56
+ $X2=0 $Y2=0
cc_376 N_A_324_102#_c_335_n N_VGND_c_1835_n 0.0103197f $X=1.695 $Y=1.17 $X2=0
+ $Y2=0
cc_377 N_A_324_102#_c_336_n N_VGND_c_1835_n 0.0028757f $X=1.805 $Y=1.58 $X2=0
+ $Y2=0
cc_378 N_A_324_102#_c_339_n N_VGND_c_1835_n 0.0146038f $X=2.765 $Y=0.915 $X2=0
+ $Y2=0
cc_379 N_A_324_102#_c_335_n N_VGND_c_1851_n 7.83062e-19 $X=1.695 $Y=1.17 $X2=0
+ $Y2=0
cc_380 N_A_324_102#_c_339_n N_VGND_c_1851_n 0.00733575f $X=2.765 $Y=0.915 $X2=0
+ $Y2=0
cc_381 N_SCE_c_422_n N_CLK_M1025_g 0.0165584f $X=3.265 $Y=0.805 $X2=0 $Y2=0
cc_382 N_SCE_c_424_n N_CLK_M1027_g 0.00342529f $X=3.34 $Y=2.03 $X2=0 $Y2=0
cc_383 N_SCE_c_424_n N_CLK_c_507_n 0.0165584f $X=3.34 $Y=2.03 $X2=0 $Y2=0
cc_384 N_SCE_c_421_n N_A_702_47#_c_1023_n 0.00195912f $X=2.87 $Y=0.73 $X2=0
+ $Y2=0
cc_385 N_SCE_c_422_n N_A_702_47#_c_1023_n 0.0102191f $X=3.265 $Y=0.805 $X2=0
+ $Y2=0
cc_386 N_SCE_c_424_n N_A_702_47#_c_1023_n 0.0013298f $X=3.34 $Y=2.03 $X2=0 $Y2=0
cc_387 SCE N_A_702_47#_c_1023_n 0.00146321f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_388 SCE N_A_702_47#_c_1025_n 0.0263759f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_389 N_SCE_c_427_n N_A_702_47#_c_1025_n 0.00121229f $X=2.78 $Y=0.195 $X2=0
+ $Y2=0
cc_390 N_SCE_c_424_n N_A_702_47#_c_1043_n 8.73938e-19 $X=3.34 $Y=2.03 $X2=0
+ $Y2=0
cc_391 N_SCE_M1000_g N_A_27_408#_c_1414_n 0.0177786f $X=0.905 $Y=0.85 $X2=0
+ $Y2=0
cc_392 N_SCE_M1000_g N_VPWR_c_1446_n 0.00997021f $X=0.905 $Y=0.85 $X2=0 $Y2=0
cc_393 N_SCE_M1026_g N_VPWR_c_1447_n 0.00391859f $X=3.105 $Y=2.725 $X2=0 $Y2=0
cc_394 N_SCE_M1000_g N_VPWR_c_1460_n 0.00334468f $X=0.905 $Y=0.85 $X2=0 $Y2=0
cc_395 N_SCE_M1026_g N_VPWR_c_1461_n 0.00327695f $X=3.105 $Y=2.725 $X2=0 $Y2=0
cc_396 N_SCE_M1000_g N_VPWR_c_1445_n 0.00388565f $X=0.905 $Y=0.85 $X2=0 $Y2=0
cc_397 N_SCE_M1026_g N_VPWR_c_1445_n 0.00667022f $X=3.105 $Y=2.725 $X2=0 $Y2=0
cc_398 N_SCE_M1000_g N_A_196_128#_c_1622_n 0.0104602f $X=0.905 $Y=0.85 $X2=0
+ $Y2=0
cc_399 N_SCE_c_417_n N_A_196_128#_c_1622_n 0.00332023f $X=2.09 $Y=0.195 $X2=0
+ $Y2=0
cc_400 N_SCE_M1038_g N_A_196_128#_c_1609_n 0.00357386f $X=2.165 $Y=0.85 $X2=0
+ $Y2=0
cc_401 N_SCE_M1000_g N_A_196_128#_c_1610_n 0.00504003f $X=0.905 $Y=0.85 $X2=0
+ $Y2=0
cc_402 N_SCE_c_424_n N_A_196_128#_c_1611_n 7.4941e-19 $X=3.34 $Y=2.03 $X2=0
+ $Y2=0
cc_403 N_SCE_c_431_n N_A_196_128#_c_1611_n 0.00760439f $X=3.34 $Y=2.105 $X2=0
+ $Y2=0
cc_404 N_SCE_M1026_g N_A_196_128#_c_1649_n 0.00724946f $X=3.105 $Y=2.725 $X2=0
+ $Y2=0
cc_405 N_SCE_M1026_g N_A_196_128#_c_1663_n 0.0120842f $X=3.105 $Y=2.725 $X2=0
+ $Y2=0
cc_406 N_SCE_M1026_g N_A_196_128#_c_1616_n 0.0124714f $X=3.105 $Y=2.725 $X2=0
+ $Y2=0
cc_407 N_SCE_M1026_g N_A_196_128#_c_1617_n 0.00352959f $X=3.105 $Y=2.725 $X2=0
+ $Y2=0
cc_408 N_SCE_M1000_g N_VGND_c_1834_n 0.00173511f $X=0.905 $Y=0.85 $X2=0 $Y2=0
cc_409 N_SCE_c_418_n N_VGND_c_1834_n 0.0112941f $X=0.98 $Y=0.195 $X2=0 $Y2=0
cc_410 N_SCE_c_417_n N_VGND_c_1835_n 0.0226633f $X=2.09 $Y=0.195 $X2=0 $Y2=0
cc_411 N_SCE_M1038_g N_VGND_c_1835_n 0.0119039f $X=2.165 $Y=0.85 $X2=0 $Y2=0
cc_412 SCE N_VGND_c_1835_n 0.0173941f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_413 N_SCE_c_418_n N_VGND_c_1841_n 0.0289955f $X=0.98 $Y=0.195 $X2=0 $Y2=0
cc_414 N_SCE_c_417_n N_VGND_c_1847_n 0.026736f $X=2.09 $Y=0.195 $X2=0 $Y2=0
cc_415 N_SCE_c_422_n N_VGND_c_1847_n 0.00307994f $X=3.265 $Y=0.805 $X2=0 $Y2=0
cc_416 SCE N_VGND_c_1847_n 0.0525072f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_417 N_SCE_c_417_n N_VGND_c_1851_n 0.0325009f $X=2.09 $Y=0.195 $X2=0 $Y2=0
cc_418 N_SCE_c_418_n N_VGND_c_1851_n 0.0105985f $X=0.98 $Y=0.195 $X2=0 $Y2=0
cc_419 N_SCE_c_420_n N_VGND_c_1851_n 0.0101953f $X=2.615 $Y=0.195 $X2=0 $Y2=0
cc_420 N_SCE_c_422_n N_VGND_c_1851_n 0.00381819f $X=3.265 $Y=0.805 $X2=0 $Y2=0
cc_421 N_SCE_c_425_n N_VGND_c_1851_n 0.00846667f $X=2.165 $Y=0.195 $X2=0 $Y2=0
cc_422 SCE N_VGND_c_1851_n 0.0297684f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_423 N_SCE_c_427_n N_VGND_c_1851_n 0.0100791f $X=2.78 $Y=0.195 $X2=0 $Y2=0
cc_424 N_CLK_M1025_g N_A_702_47#_c_1013_n 0.019091f $X=3.85 $Y=0.445 $X2=0 $Y2=0
cc_425 N_CLK_M1025_g N_A_702_47#_c_1014_n 0.00282419f $X=3.85 $Y=0.445 $X2=0
+ $Y2=0
cc_426 CLK N_A_702_47#_c_1014_n 0.0211356f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_427 N_CLK_M1027_g N_A_702_47#_M1016_g 0.0270302f $X=4.19 $Y=2.735 $X2=0 $Y2=0
cc_428 CLK N_A_702_47#_c_1021_n 0.0108738f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_429 N_CLK_c_507_n N_A_702_47#_c_1021_n 0.00332682f $X=4.08 $Y=1.32 $X2=0
+ $Y2=0
cc_430 N_CLK_c_507_n N_A_702_47#_c_1022_n 0.0307925f $X=4.08 $Y=1.32 $X2=0 $Y2=0
cc_431 N_CLK_M1025_g N_A_702_47#_c_1023_n 0.0116788f $X=3.85 $Y=0.445 $X2=0
+ $Y2=0
cc_432 N_CLK_M1027_g N_A_702_47#_c_1023_n 0.00337706f $X=4.19 $Y=2.735 $X2=0
+ $Y2=0
cc_433 CLK N_A_702_47#_c_1023_n 0.0762165f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_434 N_CLK_c_507_n N_A_702_47#_c_1023_n 0.015776f $X=4.08 $Y=1.32 $X2=0 $Y2=0
cc_435 N_CLK_M1027_g N_A_702_47#_c_1041_n 0.013038f $X=4.19 $Y=2.735 $X2=0 $Y2=0
cc_436 N_CLK_M1027_g N_A_702_47#_c_1024_n 0.0307925f $X=4.19 $Y=2.735 $X2=0
+ $Y2=0
cc_437 N_CLK_M1025_g N_A_702_47#_c_1025_n 0.00287898f $X=3.85 $Y=0.445 $X2=0
+ $Y2=0
cc_438 N_CLK_M1027_g N_A_702_47#_c_1043_n 0.00538298f $X=4.19 $Y=2.735 $X2=0
+ $Y2=0
cc_439 CLK N_A_702_47#_c_1043_n 0.0265388f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_440 N_CLK_c_507_n N_A_702_47#_c_1043_n 0.00876639f $X=4.08 $Y=1.32 $X2=0
+ $Y2=0
cc_441 N_CLK_M1027_g N_VPWR_c_1448_n 0.00772087f $X=4.19 $Y=2.735 $X2=0 $Y2=0
cc_442 N_CLK_M1027_g N_VPWR_c_1461_n 0.0032999f $X=4.19 $Y=2.735 $X2=0 $Y2=0
cc_443 N_CLK_M1027_g N_VPWR_c_1445_n 0.00504806f $X=4.19 $Y=2.735 $X2=0 $Y2=0
cc_444 N_CLK_M1027_g N_A_196_128#_c_1616_n 0.00329656f $X=4.19 $Y=2.735 $X2=0
+ $Y2=0
cc_445 N_CLK_M1027_g N_A_196_128#_c_1667_n 0.0128287f $X=4.19 $Y=2.735 $X2=0
+ $Y2=0
cc_446 N_CLK_M1027_g N_A_196_128#_c_1620_n 0.00324017f $X=4.19 $Y=2.735 $X2=0
+ $Y2=0
cc_447 CLK N_A_196_128#_c_1613_n 7.46347e-19 $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_448 N_CLK_M1025_g N_VGND_c_1836_n 0.00305839f $X=3.85 $Y=0.445 $X2=0 $Y2=0
cc_449 CLK N_VGND_c_1836_n 0.0184233f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_450 N_CLK_c_507_n N_VGND_c_1836_n 7.658e-19 $X=4.08 $Y=1.32 $X2=0 $Y2=0
cc_451 N_CLK_M1025_g N_VGND_c_1847_n 0.0057945f $X=3.85 $Y=0.445 $X2=0 $Y2=0
cc_452 N_CLK_M1025_g N_VGND_c_1851_n 0.0120209f $X=3.85 $Y=0.445 $X2=0 $Y2=0
cc_453 CLK N_VGND_c_1851_n 0.0038669f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_454 N_A_871_47#_M1019_g N_A_1263_31#_c_719_n 0.0611725f $X=6.03 $Y=0.495
+ $X2=0 $Y2=0
cc_455 N_A_871_47#_c_561_n N_A_1263_31#_c_726_n 0.00200928f $X=6.975 $Y=2.84
+ $X2=0 $Y2=0
cc_456 N_A_871_47#_c_560_n N_A_1263_31#_c_727_n 0.0105904f $X=6.89 $Y=2.03 $X2=0
+ $Y2=0
cc_457 N_A_871_47#_c_561_n N_A_1263_31#_c_727_n 0.00116346f $X=6.975 $Y=2.84
+ $X2=0 $Y2=0
cc_458 N_A_871_47#_M1023_g N_A_1263_31#_c_728_n 0.00136851f $X=5.6 $Y=2.525
+ $X2=0 $Y2=0
cc_459 N_A_871_47#_c_550_n N_A_1263_31#_c_728_n 0.00619375f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_460 N_A_871_47#_c_559_n N_A_1263_31#_c_728_n 0.00653849f $X=6.165 $Y=2.865
+ $X2=0 $Y2=0
cc_461 N_A_871_47#_c_560_n N_A_1263_31#_c_728_n 0.00292247f $X=6.89 $Y=2.03
+ $X2=0 $Y2=0
cc_462 N_A_871_47#_c_566_n N_A_1263_31#_c_728_n 0.00705195f $X=6.245 $Y=2.03
+ $X2=0 $Y2=0
cc_463 N_A_871_47#_c_557_n N_A_1263_31#_c_729_n 0.00340648f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_464 N_A_871_47#_c_560_n N_A_1263_31#_c_729_n 0.00730841f $X=6.89 $Y=2.03
+ $X2=0 $Y2=0
cc_465 N_A_871_47#_M1019_g N_A_1263_31#_c_720_n 6.41757e-19 $X=6.03 $Y=0.495
+ $X2=0 $Y2=0
cc_466 N_A_871_47#_c_557_n N_A_1263_31#_c_721_n 0.0119879f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_467 N_A_871_47#_c_550_n N_A_1263_31#_c_721_n 7.17586e-19 $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_468 N_A_871_47#_c_560_n N_A_1263_31#_c_721_n 0.032978f $X=6.89 $Y=2.03 $X2=0
+ $Y2=0
cc_469 N_A_871_47#_c_557_n N_A_1263_31#_c_722_n 7.31451e-19 $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_470 N_A_871_47#_c_550_n N_A_1263_31#_c_722_n 0.0234027f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_471 N_A_871_47#_c_560_n N_A_1263_31#_c_722_n 0.0038933f $X=6.89 $Y=2.03 $X2=0
+ $Y2=0
cc_472 N_A_871_47#_c_560_n N_A_1263_31#_c_732_n 0.0139542f $X=6.89 $Y=2.03 $X2=0
+ $Y2=0
cc_473 N_A_871_47#_c_561_n N_A_1263_31#_c_732_n 0.014938f $X=6.975 $Y=2.84 $X2=0
+ $Y2=0
cc_474 N_A_871_47#_c_562_n N_A_1263_31#_c_732_n 0.0158143f $X=7.63 $Y=2.925
+ $X2=0 $Y2=0
cc_475 N_A_871_47#_c_564_n N_A_1263_31#_c_732_n 0.049669f $X=7.715 $Y=2.84 $X2=0
+ $Y2=0
cc_476 N_A_871_47#_c_592_p N_A_1263_31#_c_732_n 0.0138437f $X=7.8 $Y=1.9 $X2=0
+ $Y2=0
cc_477 N_A_871_47#_c_550_n N_A_1263_31#_c_724_n 0.00265698f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_478 N_A_871_47#_M1019_g N_A_1263_31#_c_725_n 0.00818237f $X=6.03 $Y=0.495
+ $X2=0 $Y2=0
cc_479 N_A_871_47#_c_562_n N_A_1135_57#_c_809_n 0.0084243f $X=7.63 $Y=2.925
+ $X2=0 $Y2=0
cc_480 N_A_871_47#_c_564_n N_A_1135_57#_c_809_n 5.93975e-19 $X=7.715 $Y=2.84
+ $X2=0 $Y2=0
cc_481 N_A_871_47#_c_560_n N_A_1135_57#_c_797_n 9.08281e-19 $X=6.89 $Y=2.03
+ $X2=0 $Y2=0
cc_482 N_A_871_47#_c_564_n N_A_1135_57#_M1029_g 0.00329302f $X=7.715 $Y=2.84
+ $X2=0 $Y2=0
cc_483 N_A_871_47#_c_567_n N_A_1135_57#_M1029_g 4.17435e-19 $X=9.305 $Y=1.93
+ $X2=0 $Y2=0
cc_484 N_A_871_47#_c_568_n N_A_1135_57#_M1029_g 0.0167437f $X=9.14 $Y=1.96 $X2=0
+ $Y2=0
cc_485 N_A_871_47#_c_569_n N_A_1135_57#_M1029_g 0.0046689f $X=9.52 $Y=1.93 $X2=0
+ $Y2=0
cc_486 N_A_871_47#_c_567_n N_A_1135_57#_c_799_n 6.4502e-19 $X=9.305 $Y=1.93
+ $X2=0 $Y2=0
cc_487 N_A_871_47#_c_568_n N_A_1135_57#_c_799_n 0.0137072f $X=9.14 $Y=1.96 $X2=0
+ $Y2=0
cc_488 N_A_871_47#_c_569_n N_A_1135_57#_c_799_n 0.00595195f $X=9.52 $Y=1.93
+ $X2=0 $Y2=0
cc_489 N_A_871_47#_M1002_g N_A_1135_57#_c_800_n 0.0655513f $X=9.52 $Y=0.945
+ $X2=0 $Y2=0
cc_490 N_A_871_47#_c_560_n N_A_1135_57#_c_812_n 5.524e-19 $X=6.89 $Y=2.03 $X2=0
+ $Y2=0
cc_491 N_A_871_47#_c_561_n N_A_1135_57#_c_812_n 0.00740072f $X=6.975 $Y=2.84
+ $X2=0 $Y2=0
cc_492 N_A_871_47#_c_562_n N_A_1135_57#_c_812_n 3.70052e-19 $X=7.63 $Y=2.925
+ $X2=0 $Y2=0
cc_493 N_A_871_47#_M1019_g N_A_1135_57#_c_801_n 0.00964767f $X=6.03 $Y=0.495
+ $X2=0 $Y2=0
cc_494 N_A_871_47#_M1023_g N_A_1135_57#_c_802_n 0.00920894f $X=5.6 $Y=2.525
+ $X2=0 $Y2=0
cc_495 N_A_871_47#_M1019_g N_A_1135_57#_c_802_n 0.00347747f $X=6.03 $Y=0.495
+ $X2=0 $Y2=0
cc_496 N_A_871_47#_c_555_n N_A_1135_57#_c_802_n 0.0130973f $X=6.08 $Y=2.95 $X2=0
+ $Y2=0
cc_497 N_A_871_47#_c_549_n N_A_1135_57#_c_802_n 0.0293633f $X=5.465 $Y=1.68
+ $X2=0 $Y2=0
cc_498 N_A_871_47#_c_557_n N_A_1135_57#_c_802_n 0.0247317f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_499 N_A_871_47#_c_550_n N_A_1135_57#_c_802_n 0.0257232f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_500 N_A_871_47#_c_559_n N_A_1135_57#_c_802_n 0.0260985f $X=6.165 $Y=2.865
+ $X2=0 $Y2=0
cc_501 N_A_871_47#_c_566_n N_A_1135_57#_c_802_n 0.0138412f $X=6.245 $Y=2.03
+ $X2=0 $Y2=0
cc_502 N_A_871_47#_M1019_g N_A_1135_57#_c_803_n 0.0211209f $X=6.03 $Y=0.495
+ $X2=0 $Y2=0
cc_503 N_A_871_47#_c_557_n N_A_1135_57#_c_803_n 0.0259599f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_504 N_A_871_47#_c_550_n N_A_1135_57#_c_803_n 0.00825997f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_505 N_A_871_47#_c_560_n N_A_1135_57#_c_803_n 0.00730493f $X=6.89 $Y=2.03
+ $X2=0 $Y2=0
cc_506 N_A_871_47#_c_592_p N_A_1135_57#_c_803_n 0.00729897f $X=7.8 $Y=1.9 $X2=0
+ $Y2=0
cc_507 N_A_871_47#_c_568_n N_A_1135_57#_c_803_n 0.022907f $X=9.14 $Y=1.96 $X2=0
+ $Y2=0
cc_508 N_A_871_47#_M1019_g N_A_1135_57#_c_804_n 5.71886e-19 $X=6.03 $Y=0.495
+ $X2=0 $Y2=0
cc_509 N_A_871_47#_c_549_n N_A_1135_57#_c_804_n 0.0480172f $X=5.465 $Y=1.68
+ $X2=0 $Y2=0
cc_510 N_A_871_47#_c_549_n N_A_1135_57#_c_805_n 0.0151475f $X=5.465 $Y=1.68
+ $X2=0 $Y2=0
cc_511 N_A_871_47#_c_568_n N_A_1135_57#_c_806_n 0.0245822f $X=9.14 $Y=1.96 $X2=0
+ $Y2=0
cc_512 N_A_871_47#_c_568_n N_A_1135_57#_c_808_n 0.00434543f $X=9.14 $Y=1.96
+ $X2=0 $Y2=0
cc_513 N_A_871_47#_c_562_n N_SET_B_M1020_g 0.00661329f $X=7.63 $Y=2.925 $X2=0
+ $Y2=0
cc_514 N_A_871_47#_c_564_n N_SET_B_M1020_g 0.0224071f $X=7.715 $Y=2.84 $X2=0
+ $Y2=0
cc_515 N_A_871_47#_c_592_p N_SET_B_M1020_g 0.00314235f $X=7.8 $Y=1.9 $X2=0 $Y2=0
cc_516 N_A_871_47#_c_592_p N_SET_B_c_914_n 0.00697866f $X=7.8 $Y=1.9 $X2=0 $Y2=0
cc_517 N_A_871_47#_c_568_n N_SET_B_c_914_n 0.0094926f $X=9.14 $Y=1.96 $X2=0
+ $Y2=0
cc_518 N_A_871_47#_M1002_g N_SET_B_c_919_n 0.0169016f $X=9.52 $Y=0.945 $X2=0
+ $Y2=0
cc_519 N_A_871_47#_c_548_n N_A_702_47#_c_1015_n 0.0034104f $X=5.37 $Y=0.35 $X2=0
+ $Y2=0
cc_520 N_A_871_47#_c_549_n N_A_702_47#_c_1015_n 0.00911273f $X=5.465 $Y=1.68
+ $X2=0 $Y2=0
cc_521 N_A_871_47#_c_550_n N_A_702_47#_c_1015_n 0.0235188f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_522 N_A_871_47#_M1023_g N_A_702_47#_c_1027_n 0.0190774f $X=5.6 $Y=2.525 $X2=0
+ $Y2=0
cc_523 N_A_871_47#_c_555_n N_A_702_47#_c_1028_n 0.0118769f $X=6.08 $Y=2.95 $X2=0
+ $Y2=0
cc_524 N_A_871_47#_c_565_n N_A_702_47#_c_1028_n 0.00517187f $X=4.835 $Y=2.86
+ $X2=0 $Y2=0
cc_525 N_A_871_47#_M1023_g N_A_702_47#_c_1029_n 0.00882001f $X=5.6 $Y=2.525
+ $X2=0 $Y2=0
cc_526 N_A_871_47#_c_555_n N_A_702_47#_c_1029_n 0.0111222f $X=6.08 $Y=2.95 $X2=0
+ $Y2=0
cc_527 N_A_871_47#_M1019_g N_A_702_47#_M1018_g 0.0283503f $X=6.03 $Y=0.495 $X2=0
+ $Y2=0
cc_528 N_A_871_47#_c_548_n N_A_702_47#_M1018_g 0.00661016f $X=5.37 $Y=0.35 $X2=0
+ $Y2=0
cc_529 N_A_871_47#_c_549_n N_A_702_47#_M1018_g 0.0190038f $X=5.465 $Y=1.68 $X2=0
+ $Y2=0
cc_530 N_A_871_47#_M1023_g N_A_702_47#_M1028_g 0.0116787f $X=5.6 $Y=2.525 $X2=0
+ $Y2=0
cc_531 N_A_871_47#_c_555_n N_A_702_47#_M1028_g 0.0163654f $X=6.08 $Y=2.95 $X2=0
+ $Y2=0
cc_532 N_A_871_47#_c_550_n N_A_702_47#_M1028_g 0.00765996f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_533 N_A_871_47#_c_559_n N_A_702_47#_M1028_g 0.0123291f $X=6.165 $Y=2.865
+ $X2=0 $Y2=0
cc_534 N_A_871_47#_M1001_g N_A_702_47#_c_1032_n 0.00884409f $X=9.485 $Y=2.525
+ $X2=0 $Y2=0
cc_535 N_A_871_47#_c_555_n N_A_702_47#_c_1032_n 0.00133803f $X=6.08 $Y=2.95
+ $X2=0 $Y2=0
cc_536 N_A_871_47#_c_562_n N_A_702_47#_c_1032_n 0.0122281f $X=7.63 $Y=2.925
+ $X2=0 $Y2=0
cc_537 N_A_871_47#_c_563_n N_A_702_47#_c_1032_n 0.00408675f $X=7.06 $Y=2.925
+ $X2=0 $Y2=0
cc_538 N_A_871_47#_M1001_g N_A_702_47#_c_1033_n 0.0224745f $X=9.485 $Y=2.525
+ $X2=0 $Y2=0
cc_539 N_A_871_47#_c_569_n N_A_702_47#_c_1033_n 0.00523121f $X=9.52 $Y=1.93
+ $X2=0 $Y2=0
cc_540 N_A_871_47#_M1002_g N_A_702_47#_c_1018_n 0.00523121f $X=9.52 $Y=0.945
+ $X2=0 $Y2=0
cc_541 N_A_871_47#_c_551_n N_A_702_47#_c_1021_n 0.0110439f $X=4.515 $Y=0.35
+ $X2=0 $Y2=0
cc_542 N_A_871_47#_c_548_n N_A_702_47#_c_1022_n 0.0030209f $X=5.37 $Y=0.35 $X2=0
+ $Y2=0
cc_543 N_A_871_47#_M1023_g N_A_702_47#_c_1024_n 0.0016758f $X=5.6 $Y=2.525 $X2=0
+ $Y2=0
cc_544 N_A_871_47#_c_550_n N_A_702_47#_c_1024_n 0.00660346f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_545 N_A_871_47#_M1001_g N_A_1912_463#_c_1273_n 4.28711e-19 $X=9.485 $Y=2.525
+ $X2=0 $Y2=0
cc_546 N_A_871_47#_c_567_n N_A_1912_463#_c_1273_n 0.0145023f $X=9.305 $Y=1.93
+ $X2=0 $Y2=0
cc_547 N_A_871_47#_c_569_n N_A_1912_463#_c_1273_n 0.00173007f $X=9.52 $Y=1.93
+ $X2=0 $Y2=0
cc_548 N_A_871_47#_M1002_g N_A_1912_463#_c_1266_n 0.0269102f $X=9.52 $Y=0.945
+ $X2=0 $Y2=0
cc_549 N_A_871_47#_c_567_n N_A_1912_463#_c_1266_n 0.0104614f $X=9.305 $Y=1.93
+ $X2=0 $Y2=0
cc_550 N_A_871_47#_c_561_n N_VPWR_M1032_d 0.00667255f $X=6.975 $Y=2.84 $X2=0
+ $Y2=0
cc_551 N_A_871_47#_c_564_n N_VPWR_M1020_d 0.00405471f $X=7.715 $Y=2.84 $X2=0
+ $Y2=0
cc_552 N_A_871_47#_c_568_n N_VPWR_M1020_d 0.00335707f $X=9.14 $Y=1.96 $X2=0
+ $Y2=0
cc_553 N_A_871_47#_c_555_n N_VPWR_c_1449_n 0.0644797f $X=6.08 $Y=2.95 $X2=0
+ $Y2=0
cc_554 N_A_871_47#_c_565_n N_VPWR_c_1449_n 0.0135067f $X=4.835 $Y=2.86 $X2=0
+ $Y2=0
cc_555 N_A_871_47#_c_555_n N_VPWR_c_1450_n 0.013738f $X=6.08 $Y=2.95 $X2=0 $Y2=0
cc_556 N_A_871_47#_c_559_n N_VPWR_c_1450_n 0.0332593f $X=6.165 $Y=2.865 $X2=0
+ $Y2=0
cc_557 N_A_871_47#_c_560_n N_VPWR_c_1450_n 0.0140335f $X=6.89 $Y=2.03 $X2=0
+ $Y2=0
cc_558 N_A_871_47#_c_561_n N_VPWR_c_1450_n 0.0357186f $X=6.975 $Y=2.84 $X2=0
+ $Y2=0
cc_559 N_A_871_47#_c_563_n N_VPWR_c_1450_n 0.0148638f $X=7.06 $Y=2.925 $X2=0
+ $Y2=0
cc_560 N_A_871_47#_c_562_n N_VPWR_c_1451_n 0.0150705f $X=7.63 $Y=2.925 $X2=0
+ $Y2=0
cc_561 N_A_871_47#_c_564_n N_VPWR_c_1451_n 0.0531934f $X=7.715 $Y=2.84 $X2=0
+ $Y2=0
cc_562 N_A_871_47#_c_568_n N_VPWR_c_1451_n 0.0275698f $X=9.14 $Y=1.96 $X2=0
+ $Y2=0
cc_563 N_A_871_47#_c_562_n N_VPWR_c_1455_n 0.0346501f $X=7.63 $Y=2.925 $X2=0
+ $Y2=0
cc_564 N_A_871_47#_c_563_n N_VPWR_c_1455_n 0.00861406f $X=7.06 $Y=2.925 $X2=0
+ $Y2=0
cc_565 N_A_871_47#_c_555_n N_VPWR_c_1445_n 0.040943f $X=6.08 $Y=2.95 $X2=0 $Y2=0
cc_566 N_A_871_47#_c_562_n N_VPWR_c_1445_n 0.0239858f $X=7.63 $Y=2.925 $X2=0
+ $Y2=0
cc_567 N_A_871_47#_c_563_n N_VPWR_c_1445_n 0.00570876f $X=7.06 $Y=2.925 $X2=0
+ $Y2=0
cc_568 N_A_871_47#_c_565_n N_VPWR_c_1445_n 0.00963977f $X=4.835 $Y=2.86 $X2=0
+ $Y2=0
cc_569 N_A_871_47#_c_548_n N_A_196_128#_M1018_s 0.00986476f $X=5.37 $Y=0.35
+ $X2=0 $Y2=0
cc_570 N_A_871_47#_c_549_n N_A_196_128#_M1018_s 0.00758576f $X=5.465 $Y=1.68
+ $X2=0 $Y2=0
cc_571 N_A_871_47#_M1016_d N_A_196_128#_c_1618_n 0.00217487f $X=4.695 $Y=2.415
+ $X2=0 $Y2=0
cc_572 N_A_871_47#_c_555_n N_A_196_128#_c_1618_n 0.00121557f $X=6.08 $Y=2.95
+ $X2=0 $Y2=0
cc_573 N_A_871_47#_c_565_n N_A_196_128#_c_1618_n 0.0186187f $X=4.835 $Y=2.86
+ $X2=0 $Y2=0
cc_574 N_A_871_47#_M1023_g N_A_196_128#_c_1612_n 0.00474207f $X=5.6 $Y=2.525
+ $X2=0 $Y2=0
cc_575 N_A_871_47#_c_549_n N_A_196_128#_c_1612_n 0.0762362f $X=5.465 $Y=1.68
+ $X2=0 $Y2=0
cc_576 N_A_871_47#_c_550_n N_A_196_128#_c_1612_n 0.00362847f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_577 N_A_871_47#_c_548_n N_A_196_128#_c_1613_n 0.0229121f $X=5.37 $Y=0.35
+ $X2=0 $Y2=0
cc_578 N_A_871_47#_c_549_n N_A_196_128#_c_1613_n 0.0154009f $X=5.465 $Y=1.68
+ $X2=0 $Y2=0
cc_579 N_A_871_47#_M1023_g N_A_196_128#_c_1621_n 0.0052867f $X=5.6 $Y=2.525
+ $X2=0 $Y2=0
cc_580 N_A_871_47#_c_555_n N_A_196_128#_c_1621_n 0.0300997f $X=6.08 $Y=2.95
+ $X2=0 $Y2=0
cc_581 N_A_871_47#_c_549_n N_A_196_128#_c_1621_n 0.00719923f $X=5.465 $Y=1.68
+ $X2=0 $Y2=0
cc_582 N_A_871_47#_c_550_n N_A_196_128#_c_1621_n 0.00315721f $X=6.245 $Y=1.68
+ $X2=0 $Y2=0
cc_583 N_A_871_47#_c_559_n A_1221_463# 0.0038329f $X=6.165 $Y=2.865 $X2=-0.19
+ $Y2=-0.245
cc_584 N_A_871_47#_c_568_n N_A_1703_379#_M1029_d 0.00262981f $X=9.14 $Y=1.96
+ $X2=-0.19 $Y2=-0.245
cc_585 N_A_871_47#_M1001_g N_A_1703_379#_c_1758_n 0.00775018f $X=9.485 $Y=2.525
+ $X2=0 $Y2=0
cc_586 N_A_871_47#_c_568_n N_A_1703_379#_c_1758_n 0.0217787f $X=9.14 $Y=1.96
+ $X2=0 $Y2=0
cc_587 N_A_871_47#_M1001_g N_A_1703_379#_c_1759_n 7.8246e-19 $X=9.485 $Y=2.525
+ $X2=0 $Y2=0
cc_588 N_A_871_47#_M1001_g N_A_1703_379#_c_1760_n 0.016507f $X=9.485 $Y=2.525
+ $X2=0 $Y2=0
cc_589 N_A_871_47#_c_567_n N_A_1703_379#_c_1760_n 0.0243991f $X=9.305 $Y=1.93
+ $X2=0 $Y2=0
cc_590 N_A_871_47#_c_568_n N_A_1703_379#_c_1760_n 0.0162274f $X=9.14 $Y=1.96
+ $X2=0 $Y2=0
cc_591 N_A_871_47#_c_569_n N_A_1703_379#_c_1760_n 0.00325237f $X=9.52 $Y=1.93
+ $X2=0 $Y2=0
cc_592 N_A_871_47#_M1001_g N_A_1810_463#_c_1791_n 0.0067365f $X=9.485 $Y=2.525
+ $X2=0 $Y2=0
cc_593 N_A_871_47#_M1001_g N_A_1810_463#_c_1793_n 0.00762358f $X=9.485 $Y=2.525
+ $X2=0 $Y2=0
cc_594 N_A_871_47#_M1019_g N_VGND_c_1837_n 0.00211738f $X=6.03 $Y=0.495 $X2=0
+ $Y2=0
cc_595 N_A_871_47#_M1019_g N_VGND_c_1848_n 0.0053602f $X=6.03 $Y=0.495 $X2=0
+ $Y2=0
cc_596 N_A_871_47#_c_548_n N_VGND_c_1848_n 0.0550731f $X=5.37 $Y=0.35 $X2=0
+ $Y2=0
cc_597 N_A_871_47#_c_551_n N_VGND_c_1848_n 0.0169678f $X=4.515 $Y=0.35 $X2=0
+ $Y2=0
cc_598 N_A_871_47#_M1002_g N_VGND_c_1849_n 5.42344e-19 $X=9.52 $Y=0.945 $X2=0
+ $Y2=0
cc_599 N_A_871_47#_M1037_d N_VGND_c_1851_n 0.00234978f $X=4.355 $Y=0.235 $X2=0
+ $Y2=0
cc_600 N_A_871_47#_M1019_g N_VGND_c_1851_n 0.0103375f $X=6.03 $Y=0.495 $X2=0
+ $Y2=0
cc_601 N_A_871_47#_c_548_n N_VGND_c_1851_n 0.0333804f $X=5.37 $Y=0.35 $X2=0
+ $Y2=0
cc_602 N_A_871_47#_c_551_n N_VGND_c_1851_n 0.0109496f $X=4.515 $Y=0.35 $X2=0
+ $Y2=0
cc_603 N_A_1263_31#_c_726_n N_A_1135_57#_c_809_n 0.00516017f $X=6.39 $Y=2.205
+ $X2=0 $Y2=0
cc_604 N_A_1263_31#_c_732_n N_A_1135_57#_c_809_n 8.9478e-19 $X=7.365 $Y=2.505
+ $X2=0 $Y2=0
cc_605 N_A_1263_31#_c_729_n N_A_1135_57#_c_797_n 0.0065504f $X=6.725 $Y=2.055
+ $X2=0 $Y2=0
cc_606 N_A_1263_31#_c_721_n N_A_1135_57#_c_797_n 0.0109199f $X=7.23 $Y=1.685
+ $X2=0 $Y2=0
cc_607 N_A_1263_31#_c_722_n N_A_1135_57#_c_797_n 0.0217499f $X=6.785 $Y=1.68
+ $X2=0 $Y2=0
cc_608 N_A_1263_31#_c_732_n N_A_1135_57#_c_797_n 0.00682676f $X=7.365 $Y=2.505
+ $X2=0 $Y2=0
cc_609 N_A_1263_31#_c_723_n N_A_1135_57#_c_798_n 0.00105584f $X=7.22 $Y=0.825
+ $X2=0 $Y2=0
cc_610 N_A_1263_31#_c_724_n N_A_1135_57#_c_798_n 0.00496179f $X=6.725 $Y=0.98
+ $X2=0 $Y2=0
cc_611 N_A_1263_31#_c_727_n N_A_1135_57#_c_812_n 0.00620797f $X=6.65 $Y=2.13
+ $X2=0 $Y2=0
cc_612 N_A_1263_31#_c_721_n N_A_1135_57#_c_812_n 0.00315357f $X=7.23 $Y=1.685
+ $X2=0 $Y2=0
cc_613 N_A_1263_31#_c_732_n N_A_1135_57#_c_812_n 0.00500563f $X=7.365 $Y=2.505
+ $X2=0 $Y2=0
cc_614 N_A_1263_31#_c_720_n N_A_1135_57#_c_801_n 0.00745646f $X=7.055 $Y=0.955
+ $X2=0 $Y2=0
cc_615 N_A_1263_31#_c_728_n N_A_1135_57#_c_803_n 9.84913e-19 $X=6.465 $Y=2.13
+ $X2=0 $Y2=0
cc_616 N_A_1263_31#_c_720_n N_A_1135_57#_c_803_n 0.0435546f $X=7.055 $Y=0.955
+ $X2=0 $Y2=0
cc_617 N_A_1263_31#_c_721_n N_A_1135_57#_c_803_n 0.0622112f $X=7.23 $Y=1.685
+ $X2=0 $Y2=0
cc_618 N_A_1263_31#_c_722_n N_A_1135_57#_c_803_n 0.0039599f $X=6.785 $Y=1.68
+ $X2=0 $Y2=0
cc_619 N_A_1263_31#_c_723_n N_A_1135_57#_c_803_n 0.0204274f $X=7.22 $Y=0.825
+ $X2=0 $Y2=0
cc_620 N_A_1263_31#_c_724_n N_A_1135_57#_c_803_n 0.00872059f $X=6.725 $Y=0.98
+ $X2=0 $Y2=0
cc_621 N_A_1263_31#_c_725_n N_A_1135_57#_c_803_n 0.0124383f $X=6.785 $Y=1.515
+ $X2=0 $Y2=0
cc_622 N_A_1263_31#_c_721_n N_A_1135_57#_c_807_n 0.00422989f $X=7.23 $Y=1.685
+ $X2=0 $Y2=0
cc_623 N_A_1263_31#_c_723_n N_A_1135_57#_c_807_n 0.00453428f $X=7.22 $Y=0.825
+ $X2=0 $Y2=0
cc_624 N_A_1263_31#_c_725_n N_A_1135_57#_c_807_n 0.0131061f $X=6.785 $Y=1.515
+ $X2=0 $Y2=0
cc_625 N_A_1263_31#_c_721_n N_SET_B_c_914_n 0.00469461f $X=7.23 $Y=1.685 $X2=0
+ $Y2=0
cc_626 N_A_1263_31#_c_732_n N_SET_B_c_914_n 0.00529027f $X=7.365 $Y=2.505 $X2=0
+ $Y2=0
cc_627 N_A_1263_31#_c_728_n N_A_702_47#_M1028_g 0.0396577f $X=6.465 $Y=2.13
+ $X2=0 $Y2=0
cc_628 N_A_1263_31#_c_726_n N_A_702_47#_c_1032_n 0.0103107f $X=6.39 $Y=2.205
+ $X2=0 $Y2=0
cc_629 N_A_1263_31#_c_726_n N_VPWR_c_1450_n 0.00785818f $X=6.39 $Y=2.205 $X2=0
+ $Y2=0
cc_630 N_A_1263_31#_c_727_n N_VPWR_c_1450_n 0.00566914f $X=6.65 $Y=2.13 $X2=0
+ $Y2=0
cc_631 N_A_1263_31#_c_726_n N_VPWR_c_1445_n 7.88961e-19 $X=6.39 $Y=2.205 $X2=0
+ $Y2=0
cc_632 N_A_1263_31#_c_719_n N_VGND_c_1837_n 0.0131216f $X=6.39 $Y=0.815 $X2=0
+ $Y2=0
cc_633 N_A_1263_31#_c_720_n N_VGND_c_1837_n 0.0213543f $X=7.055 $Y=0.955 $X2=0
+ $Y2=0
cc_634 N_A_1263_31#_c_723_n N_VGND_c_1837_n 2.85702e-19 $X=7.22 $Y=0.825 $X2=0
+ $Y2=0
cc_635 N_A_1263_31#_c_724_n N_VGND_c_1837_n 0.00755333f $X=6.725 $Y=0.98 $X2=0
+ $Y2=0
cc_636 N_A_1263_31#_c_723_n N_VGND_c_1843_n 0.00449161f $X=7.22 $Y=0.825 $X2=0
+ $Y2=0
cc_637 N_A_1263_31#_c_719_n N_VGND_c_1848_n 0.00445056f $X=6.39 $Y=0.815 $X2=0
+ $Y2=0
cc_638 N_A_1263_31#_c_719_n N_VGND_c_1851_n 0.0079903f $X=6.39 $Y=0.815 $X2=0
+ $Y2=0
cc_639 N_A_1263_31#_c_720_n N_VGND_c_1851_n 0.011029f $X=7.055 $Y=0.955 $X2=0
+ $Y2=0
cc_640 N_A_1263_31#_c_723_n N_VGND_c_1851_n 0.00751301f $X=7.22 $Y=0.825 $X2=0
+ $Y2=0
cc_641 N_A_1263_31#_c_724_n N_VGND_c_1851_n 8.04731e-19 $X=6.725 $Y=0.98 $X2=0
+ $Y2=0
cc_642 N_A_1135_57#_c_809_n N_SET_B_M1020_g 0.00995669f $X=7.15 $Y=2.205 $X2=0
+ $Y2=0
cc_643 N_A_1135_57#_M1029_g N_SET_B_M1020_g 0.00920014f $X=8.44 $Y=2.315 $X2=0
+ $Y2=0
cc_644 N_A_1135_57#_c_812_n N_SET_B_M1020_g 0.0139915f $X=7.235 $Y=2.13 $X2=0
+ $Y2=0
cc_645 N_A_1135_57#_c_797_n N_SET_B_M1021_g 0.00158864f $X=7.235 $Y=2.055 $X2=0
+ $Y2=0
cc_646 N_A_1135_57#_c_803_n N_SET_B_M1021_g 0.0137678f $X=8.365 $Y=1.335 $X2=0
+ $Y2=0
cc_647 N_A_1135_57#_c_806_n N_SET_B_M1021_g 0.00177896f $X=8.53 $Y=1.335 $X2=0
+ $Y2=0
cc_648 N_A_1135_57#_c_807_n N_SET_B_M1021_g 0.0171434f $X=7.435 $Y=1.33 $X2=0
+ $Y2=0
cc_649 N_A_1135_57#_c_808_n N_SET_B_M1021_g 0.0133123f $X=8.53 $Y=1.45 $X2=0
+ $Y2=0
cc_650 N_A_1135_57#_c_797_n N_SET_B_c_914_n 0.0179738f $X=7.235 $Y=2.055 $X2=0
+ $Y2=0
cc_651 N_A_1135_57#_M1029_g N_SET_B_c_914_n 0.00591082f $X=8.44 $Y=2.315 $X2=0
+ $Y2=0
cc_652 N_A_1135_57#_c_803_n N_SET_B_c_914_n 0.0091587f $X=8.365 $Y=1.335 $X2=0
+ $Y2=0
cc_653 N_A_1135_57#_c_798_n N_SET_B_c_919_n 4.10826e-19 $X=7.435 $Y=1.165 $X2=0
+ $Y2=0
cc_654 N_A_1135_57#_c_800_n N_SET_B_c_919_n 0.0169016f $X=9.16 $Y=1.375 $X2=0
+ $Y2=0
cc_655 N_A_1135_57#_c_798_n N_SET_B_c_920_n 0.0171434f $X=7.435 $Y=1.165 $X2=0
+ $Y2=0
cc_656 N_A_1135_57#_c_801_n N_A_702_47#_c_1015_n 0.00208478f $X=5.81 $Y=1.245
+ $X2=0 $Y2=0
cc_657 N_A_1135_57#_c_805_n N_A_702_47#_c_1015_n 3.03039e-19 $X=5.81 $Y=1.335
+ $X2=0 $Y2=0
cc_658 N_A_1135_57#_c_804_n N_A_702_47#_M1018_g 0.00208478f $X=5.82 $Y=0.725
+ $X2=0 $Y2=0
cc_659 N_A_1135_57#_c_802_n N_A_702_47#_M1028_g 9.92912e-19 $X=5.815 $Y=2.525
+ $X2=0 $Y2=0
cc_660 N_A_1135_57#_c_809_n N_A_702_47#_c_1032_n 0.00881082f $X=7.15 $Y=2.205
+ $X2=0 $Y2=0
cc_661 N_A_1135_57#_M1029_g N_A_702_47#_c_1032_n 0.0103003f $X=8.44 $Y=2.315
+ $X2=0 $Y2=0
cc_662 N_A_1135_57#_c_809_n N_VPWR_c_1450_n 8.85066e-19 $X=7.15 $Y=2.205 $X2=0
+ $Y2=0
cc_663 N_A_1135_57#_M1029_g N_VPWR_c_1451_n 0.00885457f $X=8.44 $Y=2.315 $X2=0
+ $Y2=0
cc_664 N_A_1135_57#_M1029_g N_VPWR_c_1445_n 9.39239e-19 $X=8.44 $Y=2.315 $X2=0
+ $Y2=0
cc_665 N_A_1135_57#_c_802_n N_A_196_128#_c_1612_n 0.0155552f $X=5.815 $Y=2.525
+ $X2=0 $Y2=0
cc_666 N_A_1135_57#_c_802_n N_A_196_128#_c_1621_n 0.0165939f $X=5.815 $Y=2.525
+ $X2=0 $Y2=0
cc_667 N_A_1135_57#_M1029_g N_A_1703_379#_c_1758_n 0.00757894f $X=8.44 $Y=2.315
+ $X2=0 $Y2=0
cc_668 N_A_1135_57#_M1029_g N_A_1810_463#_c_1793_n 0.00315074f $X=8.44 $Y=2.315
+ $X2=0 $Y2=0
cc_669 N_A_1135_57#_c_798_n N_VGND_c_1837_n 0.00363816f $X=7.435 $Y=1.165 $X2=0
+ $Y2=0
cc_670 N_A_1135_57#_c_803_n N_VGND_c_1837_n 8.14846e-19 $X=8.365 $Y=1.335 $X2=0
+ $Y2=0
cc_671 N_A_1135_57#_c_798_n N_VGND_c_1838_n 0.0118046f $X=7.435 $Y=1.165 $X2=0
+ $Y2=0
cc_672 N_A_1135_57#_c_798_n N_VGND_c_1911_n 0.00512664f $X=7.435 $Y=1.165 $X2=0
+ $Y2=0
cc_673 N_A_1135_57#_c_803_n N_VGND_c_1911_n 0.00891849f $X=8.365 $Y=1.335 $X2=0
+ $Y2=0
cc_674 N_A_1135_57#_c_800_n N_VGND_c_1913_n 0.00724549f $X=9.16 $Y=1.375 $X2=0
+ $Y2=0
cc_675 N_A_1135_57#_c_803_n N_VGND_c_1913_n 0.037858f $X=8.365 $Y=1.335 $X2=0
+ $Y2=0
cc_676 N_A_1135_57#_c_806_n N_VGND_c_1913_n 0.0208245f $X=8.53 $Y=1.335 $X2=0
+ $Y2=0
cc_677 N_A_1135_57#_c_808_n N_VGND_c_1913_n 0.00617033f $X=8.53 $Y=1.45 $X2=0
+ $Y2=0
cc_678 N_A_1135_57#_c_798_n N_VGND_c_1843_n 0.00345209f $X=7.435 $Y=1.165 $X2=0
+ $Y2=0
cc_679 N_A_1135_57#_c_908_p N_VGND_c_1848_n 0.00883235f $X=5.815 $Y=0.49 $X2=0
+ $Y2=0
cc_680 N_A_1135_57#_c_800_n N_VGND_c_1849_n 5.42344e-19 $X=9.16 $Y=1.375 $X2=0
+ $Y2=0
cc_681 N_A_1135_57#_c_798_n N_VGND_c_1851_n 0.00394323f $X=7.435 $Y=1.165 $X2=0
+ $Y2=0
cc_682 N_A_1135_57#_c_908_p N_VGND_c_1851_n 0.00740923f $X=5.815 $Y=0.49 $X2=0
+ $Y2=0
cc_683 N_SET_B_M1020_g N_A_702_47#_c_1032_n 0.00881443f $X=7.595 $Y=2.525 $X2=0
+ $Y2=0
cc_684 N_SET_B_c_916_n N_A_702_47#_M1006_g 0.0266033f $X=10.535 $Y=1.585 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_925_n N_A_702_47#_M1006_g 0.00155285f $X=10.62 $Y=1.675 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_919_n N_A_702_47#_M1006_g 0.0101942f $X=10.45 $Y=0.452 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_925_n N_A_702_47#_c_1020_n 0.00786439f $X=10.62 $Y=1.675 $X2=0
+ $Y2=0
cc_688 N_SET_B_M1035_g N_A_2158_231#_M1010_g 0.0327289f $X=11.44 $Y=2.625 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_916_n N_A_2158_231#_M1010_g 0.00178145f $X=10.535 $Y=1.585
+ $X2=0 $Y2=0
cc_690 N_SET_B_c_917_n N_A_2158_231#_M1010_g 0.0109645f $X=11.495 $Y=1.67 $X2=0
+ $Y2=0
cc_691 N_SET_B_c_921_n N_A_2158_231#_M1010_g 0.0198758f $X=11.495 $Y=1.505 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_913_n N_A_2158_231#_c_1194_n 0.00777177f $X=11.42 $Y=1.245
+ $X2=0 $Y2=0
cc_693 N_SET_B_c_916_n N_A_2158_231#_c_1194_n 0.014225f $X=10.535 $Y=1.585 $X2=0
+ $Y2=0
cc_694 N_SET_B_c_917_n N_A_2158_231#_c_1194_n 0.0623244f $X=11.495 $Y=1.67 $X2=0
+ $Y2=0
cc_695 N_SET_B_c_918_n N_A_2158_231#_c_1194_n 0.00372371f $X=11.495 $Y=1.67
+ $X2=0 $Y2=0
cc_696 N_SET_B_c_921_n N_A_2158_231#_c_1194_n 0.0092215f $X=11.495 $Y=1.505
+ $X2=0 $Y2=0
cc_697 N_SET_B_c_913_n N_A_2158_231#_c_1195_n 0.0318073f $X=11.42 $Y=1.245 $X2=0
+ $Y2=0
cc_698 N_SET_B_c_916_n N_A_2158_231#_c_1195_n 0.00362397f $X=10.535 $Y=1.585
+ $X2=0 $Y2=0
cc_699 N_SET_B_c_917_n N_A_2158_231#_c_1195_n 0.0045386f $X=11.495 $Y=1.67 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_913_n N_A_2158_231#_c_1196_n 3.81939e-19 $X=11.42 $Y=1.245
+ $X2=0 $Y2=0
cc_701 N_SET_B_c_915_n N_A_2158_231#_c_1196_n 7.37156e-19 $X=11.42 $Y=1.155
+ $X2=0 $Y2=0
cc_702 N_SET_B_c_915_n N_A_2158_231#_c_1200_n 0.0318073f $X=11.42 $Y=1.155 $X2=0
+ $Y2=0
cc_703 N_SET_B_c_916_n N_A_2158_231#_c_1200_n 0.00320735f $X=10.535 $Y=1.585
+ $X2=0 $Y2=0
cc_704 N_SET_B_c_919_n N_A_2158_231#_c_1200_n 0.00304235f $X=10.45 $Y=0.452
+ $X2=0 $Y2=0
cc_705 N_SET_B_c_919_n N_A_1912_463#_M1002_d 0.0111435f $X=10.45 $Y=0.452
+ $X2=-0.19 $Y2=-0.245
cc_706 N_SET_B_c_913_n N_A_1912_463#_M1031_g 0.0123378f $X=11.42 $Y=1.245 $X2=0
+ $Y2=0
cc_707 N_SET_B_c_915_n N_A_1912_463#_M1031_g 0.0115826f $X=11.42 $Y=1.155 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_918_n N_A_1912_463#_M1031_g 0.0150183f $X=11.495 $Y=1.67 $X2=0
+ $Y2=0
cc_709 N_SET_B_c_917_n N_A_1912_463#_c_1264_n 6.37061e-19 $X=11.495 $Y=1.67
+ $X2=0 $Y2=0
cc_710 N_SET_B_c_916_n N_A_1912_463#_c_1266_n 0.0614689f $X=10.535 $Y=1.585
+ $X2=0 $Y2=0
cc_711 N_SET_B_c_925_n N_A_1912_463#_c_1266_n 0.0152728f $X=10.62 $Y=1.675 $X2=0
+ $Y2=0
cc_712 N_SET_B_c_919_n N_A_1912_463#_c_1266_n 0.052337f $X=10.45 $Y=0.452 $X2=0
+ $Y2=0
cc_713 N_SET_B_M1035_g N_A_1912_463#_c_1275_n 0.0166957f $X=11.44 $Y=2.625 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_925_n N_A_1912_463#_c_1275_n 0.0132088f $X=10.62 $Y=1.675 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_917_n N_A_1912_463#_c_1275_n 0.0658602f $X=11.495 $Y=1.67 $X2=0
+ $Y2=0
cc_716 N_SET_B_c_918_n N_A_1912_463#_c_1275_n 0.00112175f $X=11.495 $Y=1.67
+ $X2=0 $Y2=0
cc_717 N_SET_B_M1035_g N_A_1912_463#_c_1276_n 0.00719726f $X=11.44 $Y=2.625
+ $X2=0 $Y2=0
cc_718 N_SET_B_M1035_g N_A_1912_463#_c_1298_n 5.03902e-19 $X=11.44 $Y=2.625
+ $X2=0 $Y2=0
cc_719 N_SET_B_c_917_n N_A_1912_463#_c_1298_n 0.00654178f $X=11.495 $Y=1.67
+ $X2=0 $Y2=0
cc_720 N_SET_B_c_918_n N_A_1912_463#_c_1298_n 6.20543e-19 $X=11.495 $Y=1.67
+ $X2=0 $Y2=0
cc_721 N_SET_B_M1035_g N_A_1912_463#_c_1278_n 0.00681144f $X=11.44 $Y=2.625
+ $X2=0 $Y2=0
cc_722 N_SET_B_c_918_n N_A_1912_463#_c_1278_n 0.00328444f $X=11.495 $Y=1.67
+ $X2=0 $Y2=0
cc_723 N_SET_B_M1035_g N_A_1912_463#_c_1279_n 0.0052412f $X=11.44 $Y=2.625 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_917_n N_A_1912_463#_c_1279_n 0.0113367f $X=11.495 $Y=1.67 $X2=0
+ $Y2=0
cc_725 N_SET_B_c_918_n N_A_1912_463#_c_1279_n 0.00355067f $X=11.495 $Y=1.67
+ $X2=0 $Y2=0
cc_726 N_SET_B_M1020_g N_VPWR_c_1451_n 0.00236964f $X=7.595 $Y=2.525 $X2=0 $Y2=0
cc_727 N_SET_B_M1035_g N_VPWR_c_1452_n 0.00198098f $X=11.44 $Y=2.625 $X2=0 $Y2=0
cc_728 N_SET_B_M1035_g N_VPWR_c_1453_n 0.00314114f $X=11.44 $Y=2.625 $X2=0 $Y2=0
cc_729 N_SET_B_M1035_g N_VPWR_c_1462_n 0.00490845f $X=11.44 $Y=2.625 $X2=0 $Y2=0
cc_730 N_SET_B_M1035_g N_VPWR_c_1445_n 0.00506877f $X=11.44 $Y=2.625 $X2=0 $Y2=0
cc_731 N_SET_B_c_919_n N_VGND_M1021_d 0.0163593f $X=10.45 $Y=0.452 $X2=0 $Y2=0
cc_732 N_SET_B_M1021_g N_VGND_c_1838_n 0.00366568f $X=7.945 $Y=0.835 $X2=0 $Y2=0
cc_733 N_SET_B_c_919_n N_VGND_c_1838_n 0.0295558f $X=10.45 $Y=0.452 $X2=0 $Y2=0
cc_734 N_SET_B_c_920_n N_VGND_c_1838_n 0.00422865f $X=8.035 $Y=0.35 $X2=0 $Y2=0
cc_735 N_SET_B_M1021_g N_VGND_c_1913_n 0.0144243f $X=7.945 $Y=0.835 $X2=0 $Y2=0
cc_736 N_SET_B_c_919_n N_VGND_c_1913_n 0.0663901f $X=10.45 $Y=0.452 $X2=0 $Y2=0
cc_737 N_SET_B_c_920_n N_VGND_c_1913_n 8.28729e-19 $X=8.035 $Y=0.35 $X2=0 $Y2=0
cc_738 N_SET_B_c_915_n N_VGND_c_1839_n 0.0039374f $X=11.42 $Y=1.155 $X2=0 $Y2=0
cc_739 N_SET_B_c_915_n N_VGND_c_1849_n 0.00415323f $X=11.42 $Y=1.155 $X2=0 $Y2=0
cc_740 N_SET_B_c_919_n N_VGND_c_1849_n 0.17804f $X=10.45 $Y=0.452 $X2=0 $Y2=0
cc_741 N_SET_B_c_920_n N_VGND_c_1849_n 0.00651318f $X=8.035 $Y=0.35 $X2=0 $Y2=0
cc_742 N_SET_B_c_915_n N_VGND_c_1851_n 0.00469432f $X=11.42 $Y=1.155 $X2=0 $Y2=0
cc_743 N_SET_B_c_919_n N_VGND_c_1851_n 0.104613f $X=10.45 $Y=0.452 $X2=0 $Y2=0
cc_744 N_SET_B_c_920_n N_VGND_c_1851_n 0.0101042f $X=8.035 $Y=0.35 $X2=0 $Y2=0
cc_745 N_SET_B_c_919_n A_1847_125# 0.00403009f $X=10.45 $Y=0.452 $X2=-0.19
+ $Y2=-0.245
cc_746 N_A_702_47#_M1006_g N_A_2158_231#_M1010_g 0.00763123f $X=10.505 $Y=0.835
+ $X2=0 $Y2=0
cc_747 N_A_702_47#_c_1020_n N_A_2158_231#_M1010_g 0.0371178f $X=10.52 $Y=1.875
+ $X2=0 $Y2=0
cc_748 N_A_702_47#_M1006_g N_A_2158_231#_c_1194_n 2.06046e-19 $X=10.505 $Y=0.835
+ $X2=0 $Y2=0
cc_749 N_A_702_47#_M1006_g N_A_2158_231#_c_1195_n 0.0209654f $X=10.505 $Y=0.835
+ $X2=0 $Y2=0
cc_750 N_A_702_47#_M1006_g N_A_2158_231#_c_1200_n 0.0176321f $X=10.505 $Y=0.835
+ $X2=0 $Y2=0
cc_751 N_A_702_47#_c_1033_n N_A_1912_463#_c_1273_n 0.0072012f $X=10.03 $Y=1.785
+ $X2=0 $Y2=0
cc_752 N_A_702_47#_c_1033_n N_A_1912_463#_c_1266_n 0.00477166f $X=10.03 $Y=1.785
+ $X2=0 $Y2=0
cc_753 N_A_702_47#_c_1017_n N_A_1912_463#_c_1266_n 0.0124373f $X=10.43 $Y=1.71
+ $X2=0 $Y2=0
cc_754 N_A_702_47#_c_1018_n N_A_1912_463#_c_1266_n 0.00774344f $X=10.105 $Y=1.71
+ $X2=0 $Y2=0
cc_755 N_A_702_47#_M1006_g N_A_1912_463#_c_1266_n 0.0167813f $X=10.505 $Y=0.835
+ $X2=0 $Y2=0
cc_756 N_A_702_47#_c_1020_n N_A_1912_463#_c_1266_n 0.00252659f $X=10.52 $Y=1.875
+ $X2=0 $Y2=0
cc_757 N_A_702_47#_c_1037_n N_A_1912_463#_c_1266_n 0.00163074f $X=10.52 $Y=3.075
+ $X2=0 $Y2=0
cc_758 N_A_702_47#_c_1017_n N_A_1912_463#_c_1275_n 0.00524794f $X=10.43 $Y=1.71
+ $X2=0 $Y2=0
cc_759 N_A_702_47#_c_1020_n N_A_1912_463#_c_1275_n 7.05812e-19 $X=10.52 $Y=1.875
+ $X2=0 $Y2=0
cc_760 N_A_702_47#_c_1037_n N_A_1912_463#_c_1275_n 0.0163124f $X=10.52 $Y=3.075
+ $X2=0 $Y2=0
cc_761 N_A_702_47#_M1016_g N_VPWR_c_1448_n 0.00734516f $X=4.62 $Y=2.735 $X2=0
+ $Y2=0
cc_762 N_A_702_47#_c_1028_n N_VPWR_c_1448_n 9.9126e-19 $X=5.11 $Y=3.075 $X2=0
+ $Y2=0
cc_763 N_A_702_47#_c_1030_n N_VPWR_c_1448_n 7.40493e-19 $X=5.185 $Y=3.15 $X2=0
+ $Y2=0
cc_764 N_A_702_47#_M1016_g N_VPWR_c_1449_n 0.00452967f $X=4.62 $Y=2.735 $X2=0
+ $Y2=0
cc_765 N_A_702_47#_c_1030_n N_VPWR_c_1449_n 0.0338741f $X=5.185 $Y=3.15 $X2=0
+ $Y2=0
cc_766 N_A_702_47#_M1028_g N_VPWR_c_1450_n 0.00248721f $X=6.03 $Y=2.525 $X2=0
+ $Y2=0
cc_767 N_A_702_47#_c_1032_n N_VPWR_c_1450_n 0.0228957f $X=10.445 $Y=3.15 $X2=0
+ $Y2=0
cc_768 N_A_702_47#_c_1032_n N_VPWR_c_1451_n 0.0267251f $X=10.445 $Y=3.15 $X2=0
+ $Y2=0
cc_769 N_A_702_47#_c_1037_n N_VPWR_c_1452_n 0.00553976f $X=10.52 $Y=3.075 $X2=0
+ $Y2=0
cc_770 N_A_702_47#_c_1032_n N_VPWR_c_1455_n 0.0310838f $X=10.445 $Y=3.15 $X2=0
+ $Y2=0
cc_771 N_A_702_47#_c_1032_n N_VPWR_c_1457_n 0.0561062f $X=10.445 $Y=3.15 $X2=0
+ $Y2=0
cc_772 N_A_702_47#_M1016_g N_VPWR_c_1445_n 0.00443906f $X=4.62 $Y=2.735 $X2=0
+ $Y2=0
cc_773 N_A_702_47#_c_1029_n N_VPWR_c_1445_n 0.0182075f $X=5.955 $Y=3.15 $X2=0
+ $Y2=0
cc_774 N_A_702_47#_c_1030_n N_VPWR_c_1445_n 0.00511492f $X=5.185 $Y=3.15 $X2=0
+ $Y2=0
cc_775 N_A_702_47#_c_1032_n N_VPWR_c_1445_n 0.116413f $X=10.445 $Y=3.15 $X2=0
+ $Y2=0
cc_776 N_A_702_47#_c_1039_n N_VPWR_c_1445_n 0.00372135f $X=6.03 $Y=3.15 $X2=0
+ $Y2=0
cc_777 N_A_702_47#_M1027_s N_A_196_128#_c_1616_n 0.00642117f $X=3.715 $Y=2.105
+ $X2=0 $Y2=0
cc_778 N_A_702_47#_c_1043_n N_A_196_128#_c_1616_n 0.00885048f $X=4.025 $Y=2.155
+ $X2=0 $Y2=0
cc_779 N_A_702_47#_M1027_s N_A_196_128#_c_1654_n 0.00835142f $X=3.715 $Y=2.105
+ $X2=0 $Y2=0
cc_780 N_A_702_47#_c_1041_n N_A_196_128#_c_1667_n 0.0129612f $X=4.67 $Y=2.09
+ $X2=0 $Y2=0
cc_781 N_A_702_47#_M1027_s N_A_196_128#_c_1655_n 0.00525417f $X=3.715 $Y=2.105
+ $X2=0 $Y2=0
cc_782 N_A_702_47#_c_1041_n N_A_196_128#_c_1655_n 0.00178644f $X=4.67 $Y=2.09
+ $X2=0 $Y2=0
cc_783 N_A_702_47#_c_1043_n N_A_196_128#_c_1655_n 0.0108729f $X=4.025 $Y=2.155
+ $X2=0 $Y2=0
cc_784 N_A_702_47#_M1016_g N_A_196_128#_c_1618_n 0.00936113f $X=4.62 $Y=2.735
+ $X2=0 $Y2=0
cc_785 N_A_702_47#_c_1038_n N_A_196_128#_c_1618_n 0.00547575f $X=4.67 $Y=2.18
+ $X2=0 $Y2=0
cc_786 N_A_702_47#_c_1041_n N_A_196_128#_c_1618_n 0.0186421f $X=4.67 $Y=2.09
+ $X2=0 $Y2=0
cc_787 N_A_702_47#_M1016_g N_A_196_128#_c_1612_n 6.8096e-19 $X=4.62 $Y=2.735
+ $X2=0 $Y2=0
cc_788 N_A_702_47#_c_1015_n N_A_196_128#_c_1612_n 0.0181986f $X=5.525 $Y=1.2
+ $X2=0 $Y2=0
cc_789 N_A_702_47#_c_1027_n N_A_196_128#_c_1612_n 0.0107653f $X=5.035 $Y=2.18
+ $X2=0 $Y2=0
cc_790 N_A_702_47#_c_1028_n N_A_196_128#_c_1612_n 8.75586e-19 $X=5.11 $Y=3.075
+ $X2=0 $Y2=0
cc_791 N_A_702_47#_M1018_g N_A_196_128#_c_1612_n 0.00156435f $X=5.6 $Y=0.495
+ $X2=0 $Y2=0
cc_792 N_A_702_47#_c_1021_n N_A_196_128#_c_1612_n 0.00921257f $X=4.58 $Y=0.84
+ $X2=0 $Y2=0
cc_793 N_A_702_47#_c_1041_n N_A_196_128#_c_1612_n 0.0132017f $X=4.67 $Y=2.09
+ $X2=0 $Y2=0
cc_794 N_A_702_47#_c_1024_n N_A_196_128#_c_1612_n 0.0168567f $X=4.67 $Y=2.09
+ $X2=0 $Y2=0
cc_795 N_A_702_47#_M1016_g N_A_196_128#_c_1620_n 0.00653979f $X=4.62 $Y=2.735
+ $X2=0 $Y2=0
cc_796 N_A_702_47#_c_1028_n N_A_196_128#_c_1620_n 5.19516e-19 $X=5.11 $Y=3.075
+ $X2=0 $Y2=0
cc_797 N_A_702_47#_c_1038_n N_A_196_128#_c_1620_n 0.00116014f $X=4.67 $Y=2.18
+ $X2=0 $Y2=0
cc_798 N_A_702_47#_c_1041_n N_A_196_128#_c_1620_n 0.0130816f $X=4.67 $Y=2.09
+ $X2=0 $Y2=0
cc_799 N_A_702_47#_c_1013_n N_A_196_128#_c_1613_n 0.00370481f $X=4.28 $Y=0.765
+ $X2=0 $Y2=0
cc_800 N_A_702_47#_c_1015_n N_A_196_128#_c_1613_n 0.00534529f $X=5.525 $Y=1.2
+ $X2=0 $Y2=0
cc_801 N_A_702_47#_M1018_g N_A_196_128#_c_1613_n 0.00102374f $X=5.6 $Y=0.495
+ $X2=0 $Y2=0
cc_802 N_A_702_47#_c_1021_n N_A_196_128#_c_1613_n 0.00126223f $X=4.58 $Y=0.84
+ $X2=0 $Y2=0
cc_803 N_A_702_47#_M1016_g N_A_196_128#_c_1621_n 0.00130571f $X=4.62 $Y=2.735
+ $X2=0 $Y2=0
cc_804 N_A_702_47#_c_1028_n N_A_196_128#_c_1621_n 0.0151828f $X=5.11 $Y=3.075
+ $X2=0 $Y2=0
cc_805 N_A_702_47#_c_1032_n N_A_1703_379#_c_1758_n 0.00617063f $X=10.445 $Y=3.15
+ $X2=0 $Y2=0
cc_806 N_A_702_47#_c_1033_n N_A_1703_379#_c_1759_n 0.00442771f $X=10.03 $Y=1.785
+ $X2=0 $Y2=0
cc_807 N_A_702_47#_c_1017_n N_A_1703_379#_c_1759_n 7.6011e-19 $X=10.43 $Y=1.71
+ $X2=0 $Y2=0
cc_808 N_A_702_47#_c_1037_n N_A_1703_379#_c_1759_n 0.00740909f $X=10.52 $Y=3.075
+ $X2=0 $Y2=0
cc_809 N_A_702_47#_c_1032_n N_A_1703_379#_c_1760_n 0.0044666f $X=10.445 $Y=3.15
+ $X2=0 $Y2=0
cc_810 N_A_702_47#_c_1033_n N_A_1703_379#_c_1760_n 0.0085671f $X=10.03 $Y=1.785
+ $X2=0 $Y2=0
cc_811 N_A_702_47#_c_1032_n N_A_1810_463#_c_1791_n 0.0177083f $X=10.445 $Y=3.15
+ $X2=0 $Y2=0
cc_812 N_A_702_47#_c_1033_n N_A_1810_463#_c_1791_n 0.0064725f $X=10.03 $Y=1.785
+ $X2=0 $Y2=0
cc_813 N_A_702_47#_c_1037_n N_A_1810_463#_c_1791_n 0.0163977f $X=10.52 $Y=3.075
+ $X2=0 $Y2=0
cc_814 N_A_702_47#_c_1037_n N_A_1810_463#_c_1792_n 0.00623187f $X=10.52 $Y=3.075
+ $X2=0 $Y2=0
cc_815 N_A_702_47#_c_1032_n N_A_1810_463#_c_1793_n 0.00741659f $X=10.445 $Y=3.15
+ $X2=0 $Y2=0
cc_816 N_A_702_47#_c_1013_n N_VGND_c_1836_n 0.00317987f $X=4.28 $Y=0.765 $X2=0
+ $Y2=0
cc_817 N_A_702_47#_c_1025_n N_VGND_c_1847_n 0.0165536f $X=3.635 $Y=0.445 $X2=0
+ $Y2=0
cc_818 N_A_702_47#_c_1013_n N_VGND_c_1848_n 0.00585385f $X=4.28 $Y=0.765 $X2=0
+ $Y2=0
cc_819 N_A_702_47#_M1018_g N_VGND_c_1848_n 0.00501274f $X=5.6 $Y=0.495 $X2=0
+ $Y2=0
cc_820 N_A_702_47#_c_1021_n N_VGND_c_1848_n 3.91805e-19 $X=4.58 $Y=0.84 $X2=0
+ $Y2=0
cc_821 N_A_702_47#_M1006_g N_VGND_c_1849_n 5.57796e-19 $X=10.505 $Y=0.835 $X2=0
+ $Y2=0
cc_822 N_A_702_47#_M1025_s N_VGND_c_1851_n 0.00216892f $X=3.51 $Y=0.235 $X2=0
+ $Y2=0
cc_823 N_A_702_47#_c_1013_n N_VGND_c_1851_n 0.0097283f $X=4.28 $Y=0.765 $X2=0
+ $Y2=0
cc_824 N_A_702_47#_M1018_g N_VGND_c_1851_n 0.010419f $X=5.6 $Y=0.495 $X2=0 $Y2=0
cc_825 N_A_702_47#_c_1021_n N_VGND_c_1851_n 3.40618e-19 $X=4.58 $Y=0.84 $X2=0
+ $Y2=0
cc_826 N_A_702_47#_c_1025_n N_VGND_c_1851_n 0.011696f $X=3.635 $Y=0.445 $X2=0
+ $Y2=0
cc_827 N_A_2158_231#_c_1194_n N_A_1912_463#_M1031_g 0.0126994f $X=11.995
+ $Y=1.325 $X2=0 $Y2=0
cc_828 N_A_2158_231#_c_1196_n N_A_1912_463#_M1031_g 0.0127775f $X=12.16 $Y=0.83
+ $X2=0 $Y2=0
cc_829 N_A_2158_231#_c_1198_n N_A_1912_463#_M1031_g 0.00409326f $X=12.605
+ $Y=2.63 $X2=0 $Y2=0
cc_830 N_A_2158_231#_c_1199_n N_A_1912_463#_M1031_g 0.0052772f $X=12.16 $Y=1.325
+ $X2=0 $Y2=0
cc_831 N_A_2158_231#_c_1198_n N_A_1912_463#_c_1262_n 0.0186816f $X=12.605
+ $Y=2.63 $X2=0 $Y2=0
cc_832 N_A_2158_231#_c_1197_n N_A_1912_463#_M1005_g 4.96823e-19 $X=12.51
+ $Y=1.325 $X2=0 $Y2=0
cc_833 N_A_2158_231#_c_1198_n N_A_1912_463#_M1005_g 6.04727e-19 $X=12.605
+ $Y=2.63 $X2=0 $Y2=0
cc_834 N_A_2158_231#_c_1198_n N_A_1912_463#_c_1269_n 0.00288479f $X=12.605
+ $Y=2.63 $X2=0 $Y2=0
cc_835 N_A_2158_231#_c_1197_n N_A_1912_463#_c_1264_n 0.00754367f $X=12.51
+ $Y=1.325 $X2=0 $Y2=0
cc_836 N_A_2158_231#_c_1199_n N_A_1912_463#_c_1264_n 0.00585776f $X=12.16
+ $Y=1.325 $X2=0 $Y2=0
cc_837 N_A_2158_231#_M1010_g N_A_1912_463#_c_1275_n 0.0157532f $X=11.01 $Y=2.625
+ $X2=0 $Y2=0
cc_838 N_A_2158_231#_c_1194_n N_A_1912_463#_c_1277_n 0.00808059f $X=11.995
+ $Y=1.325 $X2=0 $Y2=0
cc_839 N_A_2158_231#_c_1198_n N_A_1912_463#_c_1277_n 0.0263331f $X=12.605
+ $Y=2.63 $X2=0 $Y2=0
cc_840 N_A_2158_231#_c_1199_n N_A_1912_463#_c_1277_n 0.00370852f $X=12.16
+ $Y=1.325 $X2=0 $Y2=0
cc_841 N_A_2158_231#_c_1197_n N_A_1912_463#_c_1298_n 0.00108398f $X=12.51
+ $Y=1.325 $X2=0 $Y2=0
cc_842 N_A_2158_231#_c_1198_n N_A_1912_463#_c_1298_n 0.026006f $X=12.605 $Y=2.63
+ $X2=0 $Y2=0
cc_843 N_A_2158_231#_c_1199_n N_A_1912_463#_c_1298_n 0.02084f $X=12.16 $Y=1.325
+ $X2=0 $Y2=0
cc_844 N_A_2158_231#_c_1198_n N_A_1912_463#_c_1278_n 0.0212083f $X=12.605
+ $Y=2.63 $X2=0 $Y2=0
cc_845 N_A_2158_231#_c_1194_n N_A_1912_463#_c_1279_n 0.00389895f $X=11.995
+ $Y=1.325 $X2=0 $Y2=0
cc_846 N_A_2158_231#_c_1196_n N_A_2598_153#_c_1372_n 0.0141016f $X=12.16 $Y=0.83
+ $X2=0 $Y2=0
cc_847 N_A_2158_231#_c_1197_n N_A_2598_153#_c_1372_n 0.00499846f $X=12.51
+ $Y=1.325 $X2=0 $Y2=0
cc_848 N_A_2158_231#_c_1198_n N_A_2598_153#_c_1378_n 0.0670897f $X=12.605
+ $Y=2.63 $X2=0 $Y2=0
cc_849 N_A_2158_231#_c_1197_n N_A_2598_153#_c_1375_n 0.0107942f $X=12.51
+ $Y=1.325 $X2=0 $Y2=0
cc_850 N_A_2158_231#_c_1198_n N_A_2598_153#_c_1375_n 0.0170718f $X=12.605
+ $Y=2.63 $X2=0 $Y2=0
cc_851 N_A_2158_231#_M1010_g N_VPWR_c_1452_n 0.00109221f $X=11.01 $Y=2.625 $X2=0
+ $Y2=0
cc_852 N_A_2158_231#_c_1198_n N_VPWR_c_1454_n 0.00974663f $X=12.605 $Y=2.63
+ $X2=0 $Y2=0
cc_853 N_A_2158_231#_M1010_g N_VPWR_c_1457_n 0.00490845f $X=11.01 $Y=2.625 $X2=0
+ $Y2=0
cc_854 N_A_2158_231#_c_1198_n N_VPWR_c_1463_n 0.00618668f $X=12.605 $Y=2.63
+ $X2=0 $Y2=0
cc_855 N_A_2158_231#_M1010_g N_VPWR_c_1445_n 0.00506877f $X=11.01 $Y=2.625 $X2=0
+ $Y2=0
cc_856 N_A_2158_231#_c_1198_n N_VPWR_c_1445_n 0.00842003f $X=12.605 $Y=2.63
+ $X2=0 $Y2=0
cc_857 N_A_2158_231#_M1010_g N_A_1810_463#_c_1791_n 0.00130176f $X=11.01
+ $Y=2.625 $X2=0 $Y2=0
cc_858 N_A_2158_231#_c_1194_n N_VGND_c_1839_n 0.01936f $X=11.995 $Y=1.325 $X2=0
+ $Y2=0
cc_859 N_A_2158_231#_c_1196_n N_VGND_c_1845_n 0.00541646f $X=12.16 $Y=0.83 $X2=0
+ $Y2=0
cc_860 N_A_2158_231#_c_1200_n N_VGND_c_1849_n 0.00415323f $X=10.955 $Y=1.155
+ $X2=0 $Y2=0
cc_861 N_A_2158_231#_c_1196_n N_VGND_c_1851_n 0.00969249f $X=12.16 $Y=0.83 $X2=0
+ $Y2=0
cc_862 N_A_2158_231#_c_1200_n N_VGND_c_1851_n 0.00469432f $X=10.955 $Y=1.155
+ $X2=0 $Y2=0
cc_863 N_A_1912_463#_c_1265_n N_A_2598_153#_M1030_g 0.0144021f $X=13.335 $Y=1.65
+ $X2=0 $Y2=0
cc_864 N_A_1912_463#_M1005_g N_A_2598_153#_c_1372_n 0.00493646f $X=13.33
+ $Y=0.975 $X2=0 $Y2=0
cc_865 N_A_1912_463#_c_1262_n N_A_2598_153#_c_1378_n 0.0115418f $X=13.255
+ $Y=1.65 $X2=0 $Y2=0
cc_866 N_A_1912_463#_c_1269_n N_A_2598_153#_c_1378_n 0.00485692f $X=13.34
+ $Y=1.725 $X2=0 $Y2=0
cc_867 N_A_1912_463#_M1005_g N_A_2598_153#_c_1373_n 0.01341f $X=13.33 $Y=0.975
+ $X2=0 $Y2=0
cc_868 N_A_1912_463#_c_1265_n N_A_2598_153#_c_1373_n 0.00901568f $X=13.335
+ $Y=1.65 $X2=0 $Y2=0
cc_869 N_A_1912_463#_M1005_g N_A_2598_153#_c_1374_n 0.0153226f $X=13.33 $Y=0.975
+ $X2=0 $Y2=0
cc_870 N_A_1912_463#_c_1265_n N_A_2598_153#_c_1374_n 0.0029232f $X=13.335
+ $Y=1.65 $X2=0 $Y2=0
cc_871 N_A_1912_463#_c_1262_n N_A_2598_153#_c_1375_n 0.00735728f $X=13.255
+ $Y=1.65 $X2=0 $Y2=0
cc_872 N_A_1912_463#_M1005_g N_A_2598_153#_c_1375_n 0.00561655f $X=13.33
+ $Y=0.975 $X2=0 $Y2=0
cc_873 N_A_1912_463#_M1005_g N_A_2598_153#_c_1376_n 0.013069f $X=13.33 $Y=0.975
+ $X2=0 $Y2=0
cc_874 N_A_1912_463#_c_1275_n N_VPWR_c_1452_n 0.0103307f $X=11.52 $Y=2.025 $X2=0
+ $Y2=0
cc_875 N_A_1912_463#_M1011_g N_VPWR_c_1453_n 0.0146237f $X=12.39 $Y=2.625 $X2=0
+ $Y2=0
cc_876 N_A_1912_463#_c_1271_n N_VPWR_c_1453_n 0.00152271f $X=12.277 $Y=2.255
+ $X2=0 $Y2=0
cc_877 N_A_1912_463#_c_1276_n N_VPWR_c_1453_n 0.0199993f $X=11.655 $Y=2.63 $X2=0
+ $Y2=0
cc_878 N_A_1912_463#_c_1277_n N_VPWR_c_1453_n 0.022048f $X=12.09 $Y=2.095 $X2=0
+ $Y2=0
cc_879 N_A_1912_463#_c_1269_n N_VPWR_c_1454_n 0.00445975f $X=13.34 $Y=1.725
+ $X2=0 $Y2=0
cc_880 N_A_1912_463#_c_1276_n N_VPWR_c_1462_n 0.00520225f $X=11.655 $Y=2.63
+ $X2=0 $Y2=0
cc_881 N_A_1912_463#_M1011_g N_VPWR_c_1463_n 0.00407914f $X=12.39 $Y=2.625 $X2=0
+ $Y2=0
cc_882 N_A_1912_463#_c_1269_n N_VPWR_c_1463_n 0.00312414f $X=13.34 $Y=1.725
+ $X2=0 $Y2=0
cc_883 N_A_1912_463#_M1011_g N_VPWR_c_1445_n 0.00425776f $X=12.39 $Y=2.625 $X2=0
+ $Y2=0
cc_884 N_A_1912_463#_c_1269_n N_VPWR_c_1445_n 0.00410284f $X=13.34 $Y=1.725
+ $X2=0 $Y2=0
cc_885 N_A_1912_463#_c_1276_n N_VPWR_c_1445_n 0.00776731f $X=11.655 $Y=2.63
+ $X2=0 $Y2=0
cc_886 N_A_1912_463#_c_1273_n N_A_1703_379#_M1017_d 0.00129794f $X=9.96 $Y=1.935
+ $X2=0 $Y2=0
cc_887 N_A_1912_463#_c_1266_n N_A_1703_379#_M1017_d 5.28981e-19 $X=10.115
+ $Y=0.92 $X2=0 $Y2=0
cc_888 N_A_1912_463#_c_1275_n N_A_1703_379#_M1017_d 0.00180341f $X=11.52
+ $Y=2.025 $X2=0 $Y2=0
cc_889 N_A_1912_463#_c_1275_n N_A_1703_379#_c_1759_n 0.0100777f $X=11.52
+ $Y=2.025 $X2=0 $Y2=0
cc_890 N_A_1912_463#_M1001_d N_A_1703_379#_c_1760_n 0.00647441f $X=9.56 $Y=2.315
+ $X2=0 $Y2=0
cc_891 N_A_1912_463#_c_1273_n N_A_1703_379#_c_1760_n 0.0424704f $X=9.96 $Y=1.935
+ $X2=0 $Y2=0
cc_892 N_A_1912_463#_c_1275_n N_A_1810_463#_c_1792_n 0.0129376f $X=11.52
+ $Y=2.025 $X2=0 $Y2=0
cc_893 N_A_1912_463#_M1031_g N_VGND_c_1839_n 0.00584217f $X=11.945 $Y=0.835
+ $X2=0 $Y2=0
cc_894 N_A_1912_463#_M1005_g N_VGND_c_1840_n 0.0130043f $X=13.33 $Y=0.975 $X2=0
+ $Y2=0
cc_895 N_A_1912_463#_M1031_g N_VGND_c_1845_n 0.00400506f $X=11.945 $Y=0.835
+ $X2=0 $Y2=0
cc_896 N_A_1912_463#_M1005_g N_VGND_c_1845_n 0.00336309f $X=13.33 $Y=0.975 $X2=0
+ $Y2=0
cc_897 N_A_1912_463#_M1031_g N_VGND_c_1851_n 0.00469432f $X=11.945 $Y=0.835
+ $X2=0 $Y2=0
cc_898 N_A_1912_463#_M1005_g N_VGND_c_1851_n 0.00420878f $X=13.33 $Y=0.975 $X2=0
+ $Y2=0
cc_899 N_A_2598_153#_M1030_g N_VPWR_c_1454_n 0.0283369f $X=13.925 $Y=2.465 $X2=0
+ $Y2=0
cc_900 N_A_2598_153#_c_1378_n N_VPWR_c_1454_n 0.00321344f $X=13.125 $Y=1.98
+ $X2=0 $Y2=0
cc_901 N_A_2598_153#_c_1373_n N_VPWR_c_1454_n 0.0348304f $X=13.81 $Y=1.46 $X2=0
+ $Y2=0
cc_902 N_A_2598_153#_c_1374_n N_VPWR_c_1454_n 0.00505597f $X=13.81 $Y=1.46 $X2=0
+ $Y2=0
cc_903 N_A_2598_153#_M1030_g N_VPWR_c_1464_n 0.00525069f $X=13.925 $Y=2.465
+ $X2=0 $Y2=0
cc_904 N_A_2598_153#_M1030_g N_VPWR_c_1445_n 0.00979769f $X=13.925 $Y=2.465
+ $X2=0 $Y2=0
cc_905 N_A_2598_153#_c_1378_n N_VPWR_c_1445_n 0.0119997f $X=13.125 $Y=1.98 $X2=0
+ $Y2=0
cc_906 N_A_2598_153#_c_1374_n Q 0.00246766f $X=13.81 $Y=1.46 $X2=0 $Y2=0
cc_907 N_A_2598_153#_c_1373_n Q 0.0269566f $X=13.81 $Y=1.46 $X2=0 $Y2=0
cc_908 N_A_2598_153#_c_1374_n Q 0.0167362f $X=13.81 $Y=1.46 $X2=0 $Y2=0
cc_909 N_A_2598_153#_c_1376_n Q 0.00567283f $X=13.822 $Y=1.295 $X2=0 $Y2=0
cc_910 N_A_2598_153#_c_1376_n N_Q_c_1817_n 0.00208348f $X=13.822 $Y=1.295 $X2=0
+ $Y2=0
cc_911 N_A_2598_153#_c_1373_n N_VGND_c_1840_n 0.0254615f $X=13.81 $Y=1.46 $X2=0
+ $Y2=0
cc_912 N_A_2598_153#_c_1374_n N_VGND_c_1840_n 0.00239906f $X=13.81 $Y=1.46 $X2=0
+ $Y2=0
cc_913 N_A_2598_153#_c_1376_n N_VGND_c_1840_n 0.00769457f $X=13.822 $Y=1.295
+ $X2=0 $Y2=0
cc_914 N_A_2598_153#_c_1376_n N_VGND_c_1850_n 0.00482246f $X=13.822 $Y=1.295
+ $X2=0 $Y2=0
cc_915 N_A_2598_153#_c_1372_n N_VGND_c_1851_n 0.0112547f $X=13.115 $Y=0.975
+ $X2=0 $Y2=0
cc_916 N_A_2598_153#_c_1376_n N_VGND_c_1851_n 0.00995713f $X=13.822 $Y=1.295
+ $X2=0 $Y2=0
cc_917 N_A_27_408#_c_1414_n N_VPWR_M1013_d 0.00176461f $X=1.855 $Y=2.095
+ $X2=-0.19 $Y2=1.655
cc_918 N_A_27_408#_c_1413_n N_VPWR_c_1446_n 0.00155436f $X=0.26 $Y=2.185 $X2=0
+ $Y2=0
cc_919 N_A_27_408#_c_1414_n N_VPWR_c_1446_n 0.0152916f $X=1.855 $Y=2.095 $X2=0
+ $Y2=0
cc_920 N_A_27_408#_c_1413_n N_VPWR_c_1459_n 0.00600261f $X=0.26 $Y=2.185 $X2=0
+ $Y2=0
cc_921 N_A_27_408#_c_1413_n N_VPWR_c_1445_n 0.00893043f $X=0.26 $Y=2.185 $X2=0
+ $Y2=0
cc_922 N_A_27_408#_c_1414_n A_196_408# 0.00366293f $X=1.855 $Y=2.095 $X2=-0.19
+ $Y2=1.655
cc_923 N_A_27_408#_c_1414_n N_A_196_128#_M1036_d 0.00316474f $X=1.855 $Y=2.095
+ $X2=0 $Y2=0
cc_924 N_A_27_408#_c_1414_n N_A_196_128#_c_1610_n 0.00177614f $X=1.855 $Y=2.095
+ $X2=0 $Y2=0
cc_925 N_A_27_408#_M1009_d N_A_196_128#_c_1614_n 0.00696686f $X=1.88 $Y=2.04
+ $X2=0 $Y2=0
cc_926 N_A_27_408#_c_1414_n N_A_196_128#_c_1614_n 0.00588115f $X=1.855 $Y=2.095
+ $X2=0 $Y2=0
cc_927 N_A_27_408#_c_1416_n N_A_196_128#_c_1614_n 0.0206114f $X=2.02 $Y=2.095
+ $X2=0 $Y2=0
cc_928 N_A_27_408#_c_1416_n N_A_196_128#_c_1611_n 0.0168302f $X=2.02 $Y=2.095
+ $X2=0 $Y2=0
cc_929 N_A_27_408#_c_1414_n N_A_196_128#_c_1720_n 0.0209841f $X=1.855 $Y=2.095
+ $X2=0 $Y2=0
cc_930 N_VPWR_M1026_s N_A_196_128#_c_1614_n 5.34856e-19 $X=2.415 $Y=2.405 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1447_n N_A_196_128#_c_1614_n 0.00390681f $X=2.54 $Y=2.905 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1460_n N_A_196_128#_c_1614_n 0.00993038f $X=2.375 $Y=3.33 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1445_n N_A_196_128#_c_1614_n 0.0186253f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_934 N_VPWR_M1026_s N_A_196_128#_c_1611_n 0.00183507f $X=2.415 $Y=2.405 $X2=0
+ $Y2=0
cc_935 N_VPWR_M1026_s N_A_196_128#_c_1649_n 0.0160242f $X=2.415 $Y=2.405 $X2=0
+ $Y2=0
cc_936 N_VPWR_c_1447_n N_A_196_128#_c_1649_n 0.00847404f $X=2.54 $Y=2.905 $X2=0
+ $Y2=0
cc_937 N_VPWR_c_1461_n N_A_196_128#_c_1649_n 0.0027996f $X=4.24 $Y=3.33 $X2=0
+ $Y2=0
cc_938 N_VPWR_c_1445_n N_A_196_128#_c_1649_n 0.00542996f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_939 N_VPWR_M1026_s N_A_196_128#_c_1663_n 0.00736506f $X=2.415 $Y=2.405 $X2=0
+ $Y2=0
cc_940 N_VPWR_c_1447_n N_A_196_128#_c_1663_n 0.00619077f $X=2.54 $Y=2.905 $X2=0
+ $Y2=0
cc_941 N_VPWR_c_1448_n N_A_196_128#_c_1616_n 0.00652315f $X=4.405 $Y=2.93 $X2=0
+ $Y2=0
cc_942 N_VPWR_c_1461_n N_A_196_128#_c_1616_n 0.0615312f $X=4.24 $Y=3.33 $X2=0
+ $Y2=0
cc_943 N_VPWR_c_1445_n N_A_196_128#_c_1616_n 0.0371731f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_944 N_VPWR_M1026_s N_A_196_128#_c_1617_n 0.00170467f $X=2.415 $Y=2.405 $X2=0
+ $Y2=0
cc_945 N_VPWR_c_1447_n N_A_196_128#_c_1617_n 0.013931f $X=2.54 $Y=2.905 $X2=0
+ $Y2=0
cc_946 N_VPWR_c_1461_n N_A_196_128#_c_1617_n 0.0112903f $X=4.24 $Y=3.33 $X2=0
+ $Y2=0
cc_947 N_VPWR_c_1445_n N_A_196_128#_c_1617_n 0.00644478f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_948 N_VPWR_M1027_d N_A_196_128#_c_1667_n 0.00231772f $X=4.265 $Y=2.415 $X2=0
+ $Y2=0
cc_949 N_VPWR_c_1448_n N_A_196_128#_c_1667_n 0.00730491f $X=4.405 $Y=2.93 $X2=0
+ $Y2=0
cc_950 N_VPWR_c_1461_n N_A_196_128#_c_1667_n 0.00239434f $X=4.24 $Y=3.33 $X2=0
+ $Y2=0
cc_951 N_VPWR_c_1445_n N_A_196_128#_c_1667_n 0.00510835f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_952 N_VPWR_c_1445_n N_A_196_128#_c_1618_n 0.00569045f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_953 N_VPWR_c_1460_n N_A_196_128#_c_1720_n 0.00489925f $X=2.375 $Y=3.33 $X2=0
+ $Y2=0
cc_954 N_VPWR_c_1445_n N_A_196_128#_c_1720_n 0.00919153f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_955 N_VPWR_M1026_s N_A_196_128#_c_1746_n 0.00359154f $X=2.415 $Y=2.405 $X2=0
+ $Y2=0
cc_956 N_VPWR_c_1447_n N_A_196_128#_c_1746_n 0.0144703f $X=2.54 $Y=2.905 $X2=0
+ $Y2=0
cc_957 N_VPWR_c_1445_n N_A_196_128#_c_1746_n 7.79863e-19 $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_958 N_VPWR_M1027_d N_A_196_128#_c_1620_n 0.00225122f $X=4.265 $Y=2.415 $X2=0
+ $Y2=0
cc_959 N_VPWR_c_1448_n N_A_196_128#_c_1620_n 0.0083294f $X=4.405 $Y=2.93 $X2=0
+ $Y2=0
cc_960 N_VPWR_c_1445_n N_A_196_128#_c_1620_n 7.61439e-19 $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_961 N_VPWR_c_1451_n N_A_1703_379#_c_1758_n 0.0222675f $X=8.145 $Y=2.25 $X2=0
+ $Y2=0
cc_962 N_VPWR_c_1457_n N_A_1703_379#_c_1758_n 0.00742525f $X=11.09 $Y=3.33 $X2=0
+ $Y2=0
cc_963 N_VPWR_c_1445_n N_A_1703_379#_c_1758_n 0.00901465f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_964 N_VPWR_c_1452_n N_A_1810_463#_c_1791_n 0.0112121f $X=11.225 $Y=2.63 $X2=0
+ $Y2=0
cc_965 N_VPWR_c_1457_n N_A_1810_463#_c_1791_n 0.0606476f $X=11.09 $Y=3.33 $X2=0
+ $Y2=0
cc_966 N_VPWR_c_1445_n N_A_1810_463#_c_1791_n 0.0504644f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_967 N_VPWR_c_1457_n N_A_1810_463#_c_1793_n 0.01313f $X=11.09 $Y=3.33 $X2=0
+ $Y2=0
cc_968 N_VPWR_c_1445_n N_A_1810_463#_c_1793_n 0.0104144f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_969 N_VPWR_c_1445_n N_Q_M1030_d 0.00336915f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_970 N_VPWR_c_1454_n Q 0.00239408f $X=13.555 $Y=1.98 $X2=0 $Y2=0
cc_971 N_VPWR_c_1464_n Q 0.0188828f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_972 N_VPWR_c_1445_n Q 0.010808f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_973 N_A_196_128#_c_1622_n N_VGND_c_1834_n 0.0105391f $X=1.12 $Y=0.85 $X2=0
+ $Y2=0
cc_974 N_A_196_128#_c_1622_n N_VGND_c_1835_n 0.0108738f $X=1.12 $Y=0.85 $X2=0
+ $Y2=0
cc_975 N_A_196_128#_c_1609_n N_VGND_c_1835_n 0.0185794f $X=2.425 $Y=1.275 $X2=0
+ $Y2=0
cc_976 N_A_196_128#_c_1622_n N_VGND_c_1841_n 0.00461379f $X=1.12 $Y=0.85 $X2=0
+ $Y2=0
cc_977 N_A_196_128#_c_1622_n N_VGND_c_1851_n 0.00820409f $X=1.12 $Y=0.85 $X2=0
+ $Y2=0
cc_978 N_A_1703_379#_c_1760_n N_A_1810_463#_M1001_s 0.00438057f $X=10.08
+ $Y=2.455 $X2=-0.19 $Y2=1.655
cc_979 N_A_1703_379#_c_1759_n N_A_1810_463#_c_1791_n 0.0223928f $X=10.245
+ $Y=2.43 $X2=0 $Y2=0
cc_980 N_A_1703_379#_c_1760_n N_A_1810_463#_c_1791_n 0.0279292f $X=10.08
+ $Y=2.455 $X2=0 $Y2=0
cc_981 N_A_1703_379#_c_1759_n N_A_1810_463#_c_1792_n 0.0109733f $X=10.245
+ $Y=2.43 $X2=0 $Y2=0
cc_982 N_A_1703_379#_c_1758_n N_A_1810_463#_c_1793_n 0.0100104f $X=8.655 $Y=2.25
+ $X2=0 $Y2=0
cc_983 N_A_1703_379#_c_1760_n N_A_1810_463#_c_1793_n 0.0253593f $X=10.08
+ $Y=2.455 $X2=0 $Y2=0
cc_984 N_Q_c_1817_n N_VGND_c_1840_n 0.00160995f $X=14.055 $Y=0.49 $X2=0 $Y2=0
cc_985 N_Q_c_1817_n N_VGND_c_1850_n 0.019238f $X=14.055 $Y=0.49 $X2=0 $Y2=0
cc_986 N_Q_c_1817_n N_VGND_c_1851_n 0.0145419f $X=14.055 $Y=0.49 $X2=0 $Y2=0
cc_987 N_VGND_c_1838_n A_1502_125# 0.00227771f $X=7.57 $Y=0.82 $X2=-0.19
+ $Y2=-0.245
cc_988 N_VGND_c_1911_n A_1502_125# 0.00111485f $X=7.655 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_989 N_VGND_c_1913_n A_1502_125# 0.00505734f $X=8.69 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
