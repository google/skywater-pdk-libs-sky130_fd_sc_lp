* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand2_2 A B VGND VNB VPB VPWR Y
M1000 Y A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=1.0206e+12p ps=9.18e+06u
M1001 a_27_65# B VGND VNB nshort w=840000u l=150000u
+  ad=7.476e+11p pd=6.82e+06u as=2.352e+11p ps=2.24e+06u
M1002 Y A a_27_65# VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1003 VPWR B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND B a_27_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_65# A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
