* File: sky130_fd_sc_lp__a21o_0.pex.spice
* Created: Fri Aug 28 09:50:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21O_0%A_80_275# 1 2 9 11 12 15 19 23 24 29 31 32 35
+ 37 38 39
r66 38 39 8.73571 $w=2.83e-07 $l=1.7e-07 $layer=LI1_cond $X=1.23 $Y=2.055
+ $X2=1.23 $Y2=2.225
r67 37 38 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.12 $Y=1.525
+ $X2=1.12 $Y2=2.055
r68 33 35 14.4668 $w=2.33e-07 $l=2.95e-07 $layer=LI1_cond $X=1.667 $Y=0.74
+ $X2=1.667 $Y2=0.445
r69 31 33 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.667 $Y2=0.74
r70 31 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.55 $Y=0.825
+ $X2=1.205 $Y2=0.825
r71 29 39 11.5244 $w=2.83e-07 $l=2.85e-07 $layer=LI1_cond $X=1.282 $Y=2.51
+ $X2=1.282 $Y2=2.225
r72 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.875
+ $Y=1.02 $X2=0.875 $Y2=1.02
r73 21 37 11.4679 $w=4.93e-07 $l=2.47e-07 $layer=LI1_cond $X=0.957 $Y=1.278
+ $X2=0.957 $Y2=1.525
r74 21 23 6.23411 $w=4.93e-07 $l=2.58e-07 $layer=LI1_cond $X=0.957 $Y=1.278
+ $X2=0.957 $Y2=1.02
r75 20 32 31.6434 $w=9.6e-08 $l=2.87374e-07 $layer=LI1_cond $X=0.957 $Y=0.91
+ $X2=1.205 $Y2=0.825
r76 20 23 2.65795 $w=4.93e-07 $l=1.1e-07 $layer=LI1_cond $X=0.957 $Y=0.91
+ $X2=0.957 $Y2=1.02
r77 19 24 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.875 $Y=1.375
+ $X2=0.875 $Y2=1.02
r78 18 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.875 $Y=0.855
+ $X2=0.875 $Y2=1.02
r79 15 18 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.965 $Y=0.445
+ $X2=0.965 $Y2=0.855
r80 11 19 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.71 $Y=1.45
+ $X2=0.875 $Y2=1.375
r81 11 12 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.71 $Y=1.45
+ $X2=0.55 $Y2=1.45
r82 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=1.525
+ $X2=0.55 $Y2=1.45
r83 7 9 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=0.475 $Y=1.525
+ $X2=0.475 $Y2=2.735
r84 2 29 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.18
+ $Y=2.365 $X2=1.305 $Y2=2.51
r85 1 35 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.235 $X2=1.68 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_0%B1 3 7 11 12 13 14 18 19
c45 7 0 9.24364e-20 $X=1.52 $Y=2.685
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.47
+ $Y=1.245 $X2=1.47 $Y2=1.245
r47 13 14 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.585 $Y=1.295
+ $X2=1.585 $Y2=1.665
r48 13 19 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=1.585 $Y=1.295
+ $X2=1.585 $Y2=1.245
r49 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.47 $Y=1.585
+ $X2=1.47 $Y2=1.245
r50 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.47 $Y=1.585
+ $X2=1.47 $Y2=1.75
r51 10 18 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.47 $Y=1.08
+ $X2=1.47 $Y2=1.245
r52 7 12 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=1.52 $Y=2.685
+ $X2=1.52 $Y2=1.75
r53 3 10 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.455 $Y=0.445
+ $X2=1.455 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_0%A1 3 7 11 12 13 14 15 16 23 40
c49 14 0 9.24364e-20 $X=2.075 $Y=0.84
c50 11 0 1.4009e-19 $X=2.04 $Y=1.66
c51 7 0 1.15658e-19 $X=1.95 $Y=2.685
r52 29 40 1.03882 $w=3.53e-07 $l=3.2e-08 $layer=LI1_cond $X=2.132 $Y=0.957
+ $X2=2.132 $Y2=0.925
r53 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.04
+ $Y=1.32 $X2=2.04 $Y2=1.32
r54 16 24 11.1998 $w=3.53e-07 $l=3.45e-07 $layer=LI1_cond $X=2.132 $Y=1.665
+ $X2=2.132 $Y2=1.32
r55 15 24 0.81158 $w=3.53e-07 $l=2.5e-08 $layer=LI1_cond $X=2.132 $Y=1.295
+ $X2=2.132 $Y2=1.32
r56 14 40 0.876506 $w=3.53e-07 $l=2.7e-08 $layer=LI1_cond $X=2.132 $Y=0.898
+ $X2=2.132 $Y2=0.925
r57 14 38 3.83066 $w=3.53e-07 $l=1.18e-07 $layer=LI1_cond $X=2.132 $Y=0.898
+ $X2=2.132 $Y2=0.78
r58 14 15 10.1285 $w=3.53e-07 $l=3.12e-07 $layer=LI1_cond $X=2.132 $Y=0.983
+ $X2=2.132 $Y2=1.295
r59 14 29 0.844043 $w=3.53e-07 $l=2.6e-08 $layer=LI1_cond $X=2.132 $Y=0.983
+ $X2=2.132 $Y2=0.957
r60 13 38 7.51593 $w=3.43e-07 $l=2.25e-07 $layer=LI1_cond $X=2.127 $Y=0.555
+ $X2=2.127 $Y2=0.78
r61 11 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.04 $Y=1.66
+ $X2=2.04 $Y2=1.32
r62 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.66
+ $X2=2.04 $Y2=1.825
r63 10 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.155
+ $X2=2.04 $Y2=1.32
r64 7 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.95 $Y=2.685
+ $X2=1.95 $Y2=1.825
r65 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.95 $Y=0.445
+ $X2=1.95 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_0%A2 1 3 6 9 13 17 20 21 22 23 28
c43 21 0 3.53624e-21 $X=2.64 $Y=0.925
r44 22 23 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.637 $Y=1.295
+ $X2=2.637 $Y2=1.665
r45 21 22 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.637 $Y=0.925
+ $X2=2.637 $Y2=1.295
r46 21 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.61
+ $Y=1.005 $X2=2.61 $Y2=1.005
r47 19 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.61 $Y=1.345
+ $X2=2.61 $Y2=1.005
r48 19 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=1.345
+ $X2=2.61 $Y2=1.51
r49 15 17 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.38 $Y=2.14
+ $X2=2.52 $Y2=2.14
r50 13 28 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.61 $Y=0.915 $X2=2.61
+ $Y2=1.005
r51 10 13 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.34 $Y=0.84
+ $X2=2.61 $Y2=0.84
r52 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.52 $Y=2.065
+ $X2=2.52 $Y2=2.14
r53 9 20 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.52 $Y=2.065
+ $X2=2.52 $Y2=1.51
r54 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.38 $Y=2.215
+ $X2=2.38 $Y2=2.14
r55 4 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.38 $Y=2.215 $X2=2.38
+ $Y2=2.685
r56 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.34 $Y=0.765
+ $X2=2.34 $Y2=0.84
r57 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.34 $Y=0.765 $X2=2.34
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_0%X 1 2 9 11 12 13 14 15 16 17 26
r20 17 39 7.99275 $w=3.08e-07 $l=2.15e-07 $layer=LI1_cond $X=0.24 $Y=2.775
+ $X2=0.24 $Y2=2.56
r21 16 39 5.76222 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=0.24 $Y=2.405
+ $X2=0.24 $Y2=2.56
r22 15 16 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.405
r23 14 15 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r24 13 14 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r25 12 13 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.295
r26 11 26 3.51922 $w=3.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.445
+ $X2=0.24 $Y2=0.61
r27 11 12 11.1527 $w=3.08e-07 $l=3e-07 $layer=LI1_cond $X=0.24 $Y=0.625 $X2=0.24
+ $Y2=0.925
r28 11 26 0.557634 $w=3.08e-07 $l=1.5e-08 $layer=LI1_cond $X=0.24 $Y=0.625
+ $X2=0.24 $Y2=0.61
r29 7 11 3.30593 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=0.445
+ $X2=0.24 $Y2=0.445
r30 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.395 $Y=0.445
+ $X2=0.75 $Y2=0.445
r31 2 39 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.415 $X2=0.26 $Y2=2.56
r32 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.235 $X2=0.75 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_0%VPWR 1 2 9 13 15 17 22 29 30 33 36
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 27 36 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.167 $Y2=3.33
r39 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 23 33 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.71 $Y2=3.33
r43 23 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 22 36 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=2.167 $Y2=3.33
r45 22 25 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 17 33 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.71 $Y2=3.33
r49 17 19 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 11 36 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.167 $Y=3.245
+ $X2=2.167 $Y2=3.33
r53 11 13 33.2175 $w=2.53e-07 $l=7.35e-07 $layer=LI1_cond $X=2.167 $Y=3.245
+ $X2=2.167 $Y2=2.51
r54 7 33 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=3.245
+ $X2=0.71 $Y2=3.33
r55 7 9 27.2215 $w=2.88e-07 $l=6.85e-07 $layer=LI1_cond $X=0.71 $Y=3.245
+ $X2=0.71 $Y2=2.56
r56 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.025
+ $Y=2.365 $X2=2.165 $Y2=2.51
r57 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.415 $X2=0.69 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_0%A_319_473# 1 2 9 11 12 15
c28 15 0 1.12122e-19 $X=2.595 $Y=2.51
r29 13 15 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=2.612 $Y=2.175
+ $X2=2.612 $Y2=2.51
r30 11 13 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=2.465 $Y=2.09
+ $X2=2.612 $Y2=2.175
r31 11 12 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.465 $Y=2.09
+ $X2=1.87 $Y2=2.09
r32 7 12 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=1.732 $Y=2.175
+ $X2=1.87 $Y2=2.09
r33 7 9 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=1.732 $Y=2.175
+ $X2=1.732 $Y2=2.51
r34 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.455
+ $Y=2.365 $X2=2.595 $Y2=2.51
r35 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=2.365 $X2=1.735 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_0%VGND 1 2 9 11 13 15 17 22 28 32
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r45 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r46 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=0 $X2=1.215
+ $Y2=0
r47 23 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.38 $Y=0 $X2=2.16
+ $Y2=0
r48 22 31 3.9577 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.675
+ $Y2=0
r49 22 25 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.16
+ $Y2=0
r50 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r51 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=1.215
+ $Y2=0
r53 17 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=0.72
+ $Y2=0
r54 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r55 15 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r56 11 31 3.18546 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.675 $Y2=0
r57 11 13 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0.445
r58 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=0.085
+ $X2=1.215 $Y2=0
r59 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.215 $Y=0.085
+ $X2=1.215 $Y2=0.445
r60 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.235 $X2=2.555 $Y2=0.445
r61 1 9 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.235 $X2=1.215 $Y2=0.445
.ends

