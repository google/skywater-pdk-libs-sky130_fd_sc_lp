# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dlxtn_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.190000 1.285000 1.520000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.970000 0.255000 6.195000 1.005000 ;
        RECT 5.970000 1.005000 7.095000 1.175000 ;
        RECT 6.000000 1.685000 7.095000 1.855000 ;
        RECT 6.000000 1.855000 6.225000 3.075000 ;
        RECT 6.860000 1.855000 7.095000 3.075000 ;
        RECT 6.865000 1.175000 7.095000 1.685000 ;
        RECT 6.875000 0.255000 7.095000 1.005000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.280000 1.845000 0.650000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.090000  0.680000 0.470000 1.010000 ;
      RECT 0.090000  1.010000 0.260000 1.700000 ;
      RECT 0.090000  1.700000 2.685000 1.880000 ;
      RECT 0.090000  1.880000 0.410000 3.055000 ;
      RECT 0.580000  2.395000 0.835000 3.245000 ;
      RECT 0.640000  0.085000 0.885000 1.020000 ;
      RECT 1.005000  2.395000 1.305000 2.905000 ;
      RECT 1.005000  2.905000 2.130000 3.075000 ;
      RECT 1.055000  0.820000 1.865000 0.965000 ;
      RECT 1.055000  0.965000 3.410000 1.010000 ;
      RECT 1.530000  2.050000 3.225000 2.220000 ;
      RECT 1.530000  2.220000 1.780000 2.735000 ;
      RECT 1.695000  1.010000 3.410000 1.145000 ;
      RECT 1.695000  1.145000 2.140000 1.530000 ;
      RECT 1.960000  2.400000 3.695000 2.570000 ;
      RECT 1.960000  2.570000 2.130000 2.905000 ;
      RECT 2.035000  0.255000 2.235000 0.625000 ;
      RECT 2.035000  0.625000 3.950000 0.795000 ;
      RECT 2.300000  2.740000 2.560000 3.245000 ;
      RECT 2.355000  1.315000 2.685000 1.700000 ;
      RECT 2.415000  0.085000 2.745000 0.455000 ;
      RECT 2.895000  1.675000 3.225000 2.050000 ;
      RECT 3.020000  2.740000 4.035000 3.020000 ;
      RECT 3.080000  1.145000 3.410000 1.325000 ;
      RECT 3.080000  1.325000 3.695000 1.495000 ;
      RECT 3.250000  0.255000 4.300000 0.455000 ;
      RECT 3.435000  1.495000 3.695000 2.400000 ;
      RECT 3.620000  0.795000 3.950000 1.065000 ;
      RECT 3.865000  1.245000 5.035000 1.415000 ;
      RECT 3.865000  1.415000 4.035000 2.740000 ;
      RECT 4.130000  0.455000 4.300000 1.245000 ;
      RECT 4.205000  1.595000 4.385000 1.675000 ;
      RECT 4.205000  1.675000 5.375000 1.845000 ;
      RECT 4.205000  1.845000 4.415000 2.265000 ;
      RECT 4.205000  2.435000 4.915000 3.245000 ;
      RECT 4.470000  0.085000 4.720000 0.885000 ;
      RECT 4.585000  2.015000 4.915000 2.435000 ;
      RECT 4.705000  1.415000 5.035000 1.505000 ;
      RECT 4.890000  0.255000 5.385000 1.075000 ;
      RECT 5.085000  1.845000 5.375000 3.035000 ;
      RECT 5.205000  1.075000 5.385000 1.345000 ;
      RECT 5.205000  1.345000 6.695000 1.515000 ;
      RECT 5.205000  1.515000 5.375000 1.675000 ;
      RECT 5.545000  1.815000 5.830000 3.245000 ;
      RECT 5.555000  0.085000 5.800000 1.095000 ;
      RECT 6.365000  0.085000 6.695000 0.835000 ;
      RECT 6.395000  2.025000 6.690000 3.245000 ;
      RECT 7.265000  0.085000 7.495000 1.095000 ;
      RECT 7.265000  1.815000 7.585000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__dlxtn_4
