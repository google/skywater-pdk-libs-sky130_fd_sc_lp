* File: sky130_fd_sc_lp__or4_4.spice
* Created: Fri Aug 28 11:25:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4_4.pex.spice"
.subckt sky130_fd_sc_lp__or4_4  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1004 N_A_58_367#_M1004_d N_D_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.5 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_C_M1009_g N_A_58_367#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1806 AS=0.1176 PD=1.27 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1007 N_A_58_367#_M1007_d N_B_M1007_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1806 PD=1.12 PS=1.27 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g N_A_58_367#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1785 AS=0.1176 PD=1.265 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1013_d N_A_58_367#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1785 AS=0.1176 PD=1.265 PS=1.12 NRD=10.704 NRS=0 M=1 R=5.6 SA=75002.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A_58_367#_M1011_g N_X_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1011_d N_A_58_367#_M1014_g N_X_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_A_58_367#_M1015_g N_X_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 A_141_367# N_D_M1000_g N_A_58_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1012 A_213_367# N_C_M1012_g A_141_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1002 A_321_367# N_B_M1002_g A_213_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.2457 PD=1.65 PS=1.65 NRD=21.8867 NRS=21.8867 M=1 R=8.4 SA=75001.1
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g A_321_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.2457 PD=1.685 PS=1.65 NRD=10.1455 NRS=21.8867 M=1 R=8.4
+ SA=75001.6 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1008_d N_A_58_367#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.1764 PD=1.685 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4 SA=75002.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A_58_367#_M1003_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1003_d N_A_58_367#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_A_58_367#_M1010_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__or4_4.pxi.spice"
*
.ends
*
*
