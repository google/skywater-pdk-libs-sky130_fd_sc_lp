* File: sky130_fd_sc_lp__a31o_2.pxi.spice
* Created: Wed Sep  2 09:26:24 2020
* 
x_PM_SKY130_FD_SC_LP__A31O_2%A_85_23# N_A_85_23#_M1011_d N_A_85_23#_M1010_d
+ N_A_85_23#_M1008_g N_A_85_23#_M1002_g N_A_85_23#_c_60_n N_A_85_23#_M1009_g
+ N_A_85_23#_M1007_g N_A_85_23#_c_62_n N_A_85_23#_c_75_p N_A_85_23#_c_136_p
+ N_A_85_23#_c_69_n N_A_85_23#_c_70_n N_A_85_23#_c_141_p N_A_85_23#_c_71_n
+ N_A_85_23#_c_63_n N_A_85_23#_c_64_n N_A_85_23#_c_65_n
+ PM_SKY130_FD_SC_LP__A31O_2%A_85_23#
x_PM_SKY130_FD_SC_LP__A31O_2%A3 N_A3_M1003_g N_A3_M1006_g A3 N_A3_c_160_n
+ N_A3_c_161_n PM_SKY130_FD_SC_LP__A31O_2%A3
x_PM_SKY130_FD_SC_LP__A31O_2%A2 N_A2_M1004_g N_A2_M1005_g A2 N_A2_c_191_n
+ N_A2_c_192_n PM_SKY130_FD_SC_LP__A31O_2%A2
x_PM_SKY130_FD_SC_LP__A31O_2%A1 N_A1_M1011_g N_A1_M1001_g A1 A1 N_A1_c_224_n
+ N_A1_c_225_n PM_SKY130_FD_SC_LP__A31O_2%A1
x_PM_SKY130_FD_SC_LP__A31O_2%B1 N_B1_c_256_n N_B1_M1000_g N_B1_M1010_g B1
+ N_B1_c_259_n PM_SKY130_FD_SC_LP__A31O_2%B1
x_PM_SKY130_FD_SC_LP__A31O_2%VPWR N_VPWR_M1002_d N_VPWR_M1007_d N_VPWR_M1005_d
+ N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n
+ N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n VPWR N_VPWR_c_288_n
+ N_VPWR_c_279_n PM_SKY130_FD_SC_LP__A31O_2%VPWR
x_PM_SKY130_FD_SC_LP__A31O_2%X N_X_M1008_s N_X_M1002_s N_X_c_330_n X X X X X X X
+ N_X_c_352_p X PM_SKY130_FD_SC_LP__A31O_2%X
x_PM_SKY130_FD_SC_LP__A31O_2%A_342_367# N_A_342_367#_M1003_d
+ N_A_342_367#_M1001_d N_A_342_367#_c_357_n N_A_342_367#_c_361_n
+ N_A_342_367#_c_358_n N_A_342_367#_c_359_n N_A_342_367#_c_363_n
+ PM_SKY130_FD_SC_LP__A31O_2%A_342_367#
x_PM_SKY130_FD_SC_LP__A31O_2%VGND N_VGND_M1008_d N_VGND_M1009_d N_VGND_M1000_d
+ N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n
+ VGND N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n N_VGND_c_388_n
+ PM_SKY130_FD_SC_LP__A31O_2%VGND
cc_1 VNB N_A_85_23#_M1008_g 0.0353014f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.665
cc_2 VNB N_A_85_23#_M1002_g 0.00984183f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_3 VNB N_A_85_23#_c_60_n 0.0183471f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.195
cc_4 VNB N_A_85_23#_M1007_g 0.00587376f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=2.465
cc_5 VNB N_A_85_23#_c_62_n 0.00310515f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=1.705
cc_6 VNB N_A_85_23#_c_63_n 0.00361844f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.36
cc_7 VNB N_A_85_23#_c_64_n 0.0583405f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.36
cc_8 VNB N_A_85_23#_c_65_n 0.00199422f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=1.195
cc_9 VNB N_A3_M1003_g 0.00732504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A3 0.00273652f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.665
cc_11 VNB N_A3_c_160_n 0.0293398f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.525
cc_12 VNB N_A3_c_161_n 0.0179696f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_13 VNB N_A2_M1005_g 0.00792256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A2 0.00330576f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.665
cc_15 VNB N_A2_c_191_n 0.0325524f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.525
cc_16 VNB N_A2_c_192_n 0.0169277f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_17 VNB N_A1_M1001_g 0.00792444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A1 0.00774411f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.665
cc_19 VNB N_A1_c_224_n 0.0284516f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_20 VNB N_A1_c_225_n 0.0185641f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.195
cc_21 VNB N_B1_c_256_n 0.0223944f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=0.245
cc_22 VNB N_B1_M1010_g 0.0106005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB B1 0.0213492f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.665
cc_24 VNB N_B1_c_259_n 0.0597663f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_25 VNB N_VPWR_c_279_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.375
cc_26 VNB N_X_c_330_n 0.00143591f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.665
cc_27 VNB X 0.00509068f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_28 VNB N_VGND_c_380_n 0.0112389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_381_n 0.0485381f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.465
cc_30 VNB N_VGND_c_382_n 0.0335703f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.665
cc_31 VNB N_VGND_c_383_n 0.0439209f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=2.465
cc_32 VNB N_VGND_c_384_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=2.465
cc_33 VNB N_VGND_c_385_n 0.0130978f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=1.705
cc_34 VNB N_VGND_c_386_n 0.0123263f $X=-0.19 $Y=-0.245 $X2=3.355 $Y2=1.98
cc_35 VNB N_VGND_c_387_n 0.217693f $X=-0.19 $Y=-0.245 $X2=3.39 $Y2=2.91
cc_36 VNB N_VGND_c_388_n 0.0127692f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.375
cc_37 VPB N_A_85_23#_M1002_g 0.026765f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_38 VPB N_A_85_23#_M1007_g 0.0192202f $X=-0.19 $Y=1.655 $X2=1.125 $Y2=2.465
cc_39 VPB N_A_85_23#_c_62_n 8.40353e-19 $X=-0.19 $Y=1.655 $X2=1.165 $Y2=1.705
cc_40 VPB N_A_85_23#_c_69_n 0.0326639f $X=-0.19 $Y=1.655 $X2=3.26 $Y2=1.79
cc_41 VPB N_A_85_23#_c_70_n 8.22803e-19 $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.79
cc_42 VPB N_A_85_23#_c_71_n 0.0454116f $X=-0.19 $Y=1.655 $X2=3.355 $Y2=1.98
cc_43 VPB N_A3_M1003_g 0.0198643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A2_M1005_g 0.0211137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A1_M1001_g 0.0211336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_B1_M1010_g 0.0249673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_280_n 0.0137153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_281_n 0.0623229f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_49 VPB N_VPWR_c_282_n 0.00509064f $X=-0.19 $Y=1.655 $X2=1.125 $Y2=1.525
cc_50 VPB N_VPWR_c_283_n 0.00511587f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=1.025
cc_51 VPB N_VPWR_c_284_n 0.020139f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.94
cc_52 VPB N_VPWR_c_285_n 0.00632158f $X=-0.19 $Y=1.655 $X2=3.26 $Y2=1.79
cc_53 VPB N_VPWR_c_286_n 0.0185323f $X=-0.19 $Y=1.655 $X2=2.855 $Y2=0.855
cc_54 VPB N_VPWR_c_287_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.855 $Y2=0.395
cc_55 VPB N_VPWR_c_288_n 0.0375814f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.375
cc_56 VPB N_VPWR_c_279_n 0.058064f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=1.375
cc_57 VPB X 0.00112233f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.465
cc_58 N_A_85_23#_M1007_g N_A3_M1003_g 0.0189971f $X=1.125 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A_85_23#_c_62_n N_A3_M1003_g 0.00419855f $X=1.165 $Y=1.705 $X2=0 $Y2=0
cc_60 N_A_85_23#_c_69_n N_A3_M1003_g 0.0154698f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_61 N_A_85_23#_c_75_p A3 0.0184294f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_62 N_A_85_23#_c_69_n A3 0.0211969f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_63 N_A_85_23#_c_63_n A3 0.0260432f $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_64 N_A_85_23#_c_64_n A3 2.97194e-19 $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_65 N_A_85_23#_c_75_p N_A3_c_160_n 0.00522694f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_66 N_A_85_23#_c_69_n N_A3_c_160_n 0.00530517f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_67 N_A_85_23#_c_63_n N_A3_c_160_n 0.0021661f $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_68 N_A_85_23#_c_64_n N_A3_c_160_n 0.0204965f $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_69 N_A_85_23#_c_60_n N_A3_c_161_n 0.00948757f $X=0.93 $Y=1.195 $X2=0 $Y2=0
cc_70 N_A_85_23#_c_75_p N_A3_c_161_n 0.01235f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_71 N_A_85_23#_c_65_n N_A3_c_161_n 0.00349356f $X=1.165 $Y=1.195 $X2=0 $Y2=0
cc_72 N_A_85_23#_c_69_n N_A2_M1005_g 0.0114285f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_73 N_A_85_23#_c_75_p A2 0.0219008f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_74 N_A_85_23#_c_69_n A2 0.0231565f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_75 N_A_85_23#_c_75_p N_A2_c_191_n 0.00113701f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_76 N_A_85_23#_c_69_n N_A2_c_191_n 0.00121144f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_77 N_A_85_23#_c_75_p N_A2_c_192_n 0.0120917f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_78 N_A_85_23#_c_69_n N_A1_M1001_g 0.0118981f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_79 N_A_85_23#_c_75_p A1 0.0375429f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_80 N_A_85_23#_c_69_n A1 0.0389988f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_81 N_A_85_23#_c_75_p N_A1_c_224_n 0.0040905f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_82 N_A_85_23#_c_69_n N_A1_c_224_n 0.00460038f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_83 N_A_85_23#_c_75_p N_A1_c_225_n 0.0105528f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_84 N_A_85_23#_c_69_n N_B1_M1010_g 0.015319f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_85 N_A_85_23#_c_69_n B1 0.0109054f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_86 N_A_85_23#_c_69_n N_B1_c_259_n 0.00851946f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_87 N_A_85_23#_c_69_n N_VPWR_M1007_d 0.00166894f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_88 N_A_85_23#_c_70_n N_VPWR_M1007_d 9.73829e-19 $X=1.345 $Y=1.79 $X2=0 $Y2=0
cc_89 N_A_85_23#_c_69_n N_VPWR_M1005_d 0.0043514f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_90 N_A_85_23#_M1002_g N_VPWR_c_281_n 0.0291207f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_91 N_A_85_23#_c_64_n N_VPWR_c_281_n 0.00164228f $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_92 N_A_85_23#_M1007_g N_VPWR_c_282_n 0.00346341f $X=1.125 $Y=2.465 $X2=0
+ $Y2=0
cc_93 N_A_85_23#_c_69_n N_VPWR_c_282_n 0.0128182f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_94 N_A_85_23#_c_70_n N_VPWR_c_282_n 0.00793424f $X=1.345 $Y=1.79 $X2=0 $Y2=0
cc_95 N_A_85_23#_M1002_g N_VPWR_c_284_n 0.00383824f $X=0.695 $Y=2.465 $X2=0
+ $Y2=0
cc_96 N_A_85_23#_M1007_g N_VPWR_c_284_n 0.00585385f $X=1.125 $Y=2.465 $X2=0
+ $Y2=0
cc_97 N_A_85_23#_c_71_n N_VPWR_c_288_n 0.0178111f $X=3.355 $Y=1.98 $X2=0 $Y2=0
cc_98 N_A_85_23#_M1010_d N_VPWR_c_279_n 0.00371702f $X=3.215 $Y=1.835 $X2=0
+ $Y2=0
cc_99 N_A_85_23#_M1002_g N_VPWR_c_279_n 0.00711366f $X=0.695 $Y=2.465 $X2=0
+ $Y2=0
cc_100 N_A_85_23#_M1007_g N_VPWR_c_279_n 0.0107559f $X=1.125 $Y=2.465 $X2=0
+ $Y2=0
cc_101 N_A_85_23#_c_71_n N_VPWR_c_279_n 0.0100304f $X=3.355 $Y=1.98 $X2=0 $Y2=0
cc_102 N_A_85_23#_c_70_n N_X_M1002_s 4.35515e-19 $X=1.345 $Y=1.79 $X2=0 $Y2=0
cc_103 N_A_85_23#_M1008_g N_X_c_330_n 0.00136696f $X=0.5 $Y=0.665 $X2=0 $Y2=0
cc_104 N_A_85_23#_c_60_n N_X_c_330_n 0.00160342f $X=0.93 $Y=1.195 $X2=0 $Y2=0
cc_105 N_A_85_23#_c_65_n N_X_c_330_n 0.00604125f $X=1.165 $Y=1.195 $X2=0 $Y2=0
cc_106 N_A_85_23#_M1008_g X 0.00593752f $X=0.5 $Y=0.665 $X2=0 $Y2=0
cc_107 N_A_85_23#_M1002_g X 0.0207394f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_85_23#_M1007_g X 8.73308e-19 $X=1.125 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_85_23#_c_70_n X 0.0124936f $X=1.345 $Y=1.79 $X2=0 $Y2=0
cc_110 N_A_85_23#_c_63_n X 0.0379391f $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_111 N_A_85_23#_c_64_n X 0.014472f $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_112 N_A_85_23#_M1002_g X 0.00368408f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_85_23#_c_70_n X 7.21294e-19 $X=1.345 $Y=1.79 $X2=0 $Y2=0
cc_114 N_A_85_23#_c_64_n X 0.00335442f $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_115 N_A_85_23#_M1002_g X 0.0156513f $X=0.695 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_85_23#_c_69_n N_A_342_367#_M1003_d 0.00176461f $X=3.26 $Y=1.79
+ $X2=-0.19 $Y2=-0.245
cc_117 N_A_85_23#_c_69_n N_A_342_367#_M1001_d 0.00176461f $X=3.26 $Y=1.79 $X2=0
+ $Y2=0
cc_118 N_A_85_23#_c_69_n N_A_342_367#_c_357_n 0.0153678f $X=3.26 $Y=1.79 $X2=0
+ $Y2=0
cc_119 N_A_85_23#_c_69_n N_A_342_367#_c_358_n 0.044744f $X=3.26 $Y=1.79 $X2=0
+ $Y2=0
cc_120 N_A_85_23#_c_69_n N_A_342_367#_c_359_n 0.01723f $X=3.26 $Y=1.79 $X2=0
+ $Y2=0
cc_121 N_A_85_23#_c_75_p N_VGND_M1009_d 0.00823621f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_122 N_A_85_23#_c_136_p N_VGND_M1009_d 0.00539699f $X=1.345 $Y=0.94 $X2=0
+ $Y2=0
cc_123 N_A_85_23#_c_65_n N_VGND_M1009_d 0.00142271f $X=1.165 $Y=1.195 $X2=0
+ $Y2=0
cc_124 N_A_85_23#_M1008_g N_VGND_c_381_n 0.0180438f $X=0.5 $Y=0.665 $X2=0 $Y2=0
cc_125 N_A_85_23#_c_60_n N_VGND_c_381_n 6.70942e-19 $X=0.93 $Y=1.195 $X2=0 $Y2=0
cc_126 N_A_85_23#_c_69_n N_VGND_c_382_n 0.00393355f $X=3.26 $Y=1.79 $X2=0 $Y2=0
cc_127 N_A_85_23#_c_141_p N_VGND_c_383_n 0.0212513f $X=2.855 $Y=0.395 $X2=0
+ $Y2=0
cc_128 N_A_85_23#_M1008_g N_VGND_c_385_n 0.00477554f $X=0.5 $Y=0.665 $X2=0 $Y2=0
cc_129 N_A_85_23#_c_60_n N_VGND_c_385_n 0.00479301f $X=0.93 $Y=1.195 $X2=0 $Y2=0
cc_130 N_A_85_23#_M1011_d N_VGND_c_387_n 0.0048164f $X=2.675 $Y=0.245 $X2=0
+ $Y2=0
cc_131 N_A_85_23#_M1008_g N_VGND_c_387_n 0.00825815f $X=0.5 $Y=0.665 $X2=0 $Y2=0
cc_132 N_A_85_23#_c_60_n N_VGND_c_387_n 0.0082582f $X=0.93 $Y=1.195 $X2=0 $Y2=0
cc_133 N_A_85_23#_c_75_p N_VGND_c_387_n 0.033333f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_134 N_A_85_23#_c_136_p N_VGND_c_387_n 6.05226e-19 $X=1.345 $Y=0.94 $X2=0
+ $Y2=0
cc_135 N_A_85_23#_c_141_p N_VGND_c_387_n 0.0127519f $X=2.855 $Y=0.395 $X2=0
+ $Y2=0
cc_136 N_A_85_23#_M1008_g N_VGND_c_388_n 5.67122e-19 $X=0.5 $Y=0.665 $X2=0 $Y2=0
cc_137 N_A_85_23#_c_60_n N_VGND_c_388_n 0.0122166f $X=0.93 $Y=1.195 $X2=0 $Y2=0
cc_138 N_A_85_23#_c_75_p N_VGND_c_388_n 0.0194812f $X=2.69 $Y=0.94 $X2=0 $Y2=0
cc_139 N_A_85_23#_c_136_p N_VGND_c_388_n 0.0149789f $X=1.345 $Y=0.94 $X2=0 $Y2=0
cc_140 N_A_85_23#_c_63_n N_VGND_c_388_n 0.00579414f $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_141 N_A_85_23#_c_64_n N_VGND_c_388_n 0.0011027f $X=1.07 $Y=1.36 $X2=0 $Y2=0
cc_142 N_A_85_23#_c_75_p A_355_49# 0.00561753f $X=2.69 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_85_23#_c_75_p A_427_49# 0.0127782f $X=2.69 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A3_M1003_g N_A2_M1005_g 0.029847f $X=1.635 $Y=2.465 $X2=0 $Y2=0
cc_145 A3 A2 0.0258905f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A3_c_160_n A2 3.77439e-19 $X=1.61 $Y=1.36 $X2=0 $Y2=0
cc_147 A3 N_A2_c_191_n 0.00183055f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A3_c_160_n N_A2_c_191_n 0.0447806f $X=1.61 $Y=1.36 $X2=0 $Y2=0
cc_149 N_A3_c_161_n N_A2_c_192_n 0.0447806f $X=1.61 $Y=1.195 $X2=0 $Y2=0
cc_150 N_A3_M1003_g N_VPWR_c_282_n 0.00212688f $X=1.635 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A3_M1003_g N_VPWR_c_286_n 0.00585385f $X=1.635 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A3_M1003_g N_VPWR_c_279_n 0.0107539f $X=1.635 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A3_c_161_n N_VGND_c_383_n 0.00479301f $X=1.61 $Y=1.195 $X2=0 $Y2=0
cc_154 N_A3_c_161_n N_VGND_c_387_n 0.00444402f $X=1.61 $Y=1.195 $X2=0 $Y2=0
cc_155 N_A3_c_161_n N_VGND_c_388_n 0.0165769f $X=1.61 $Y=1.195 $X2=0 $Y2=0
cc_156 N_A2_M1005_g N_A1_M1001_g 0.0349523f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_157 A2 A1 0.0209146f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A2_c_191_n A1 0.00152088f $X=2.15 $Y=1.36 $X2=0 $Y2=0
cc_159 A2 N_A1_c_224_n 8.63357e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A2_c_191_n N_A1_c_224_n 0.0210528f $X=2.15 $Y=1.36 $X2=0 $Y2=0
cc_161 N_A2_c_192_n N_A1_c_225_n 0.0357984f $X=2.15 $Y=1.195 $X2=0 $Y2=0
cc_162 N_A2_M1005_g N_VPWR_c_283_n 0.00834014f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A2_M1005_g N_VPWR_c_286_n 0.0054895f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A2_M1005_g N_VPWR_c_279_n 0.0105005f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A2_M1005_g N_A_342_367#_c_357_n 7.54694e-19 $X=2.065 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A2_M1005_g N_A_342_367#_c_361_n 0.0120138f $X=2.065 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A2_M1005_g N_A_342_367#_c_358_n 0.0124105f $X=2.065 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A2_M1005_g N_A_342_367#_c_363_n 0.00108543f $X=2.065 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A2_c_192_n N_VGND_c_383_n 0.00575161f $X=2.15 $Y=1.195 $X2=0 $Y2=0
cc_170 N_A2_c_192_n N_VGND_c_387_n 0.00657254f $X=2.15 $Y=1.195 $X2=0 $Y2=0
cc_171 N_A2_c_192_n N_VGND_c_388_n 0.00334197f $X=2.15 $Y=1.195 $X2=0 $Y2=0
cc_172 N_A1_c_225_n N_B1_c_256_n 0.0194313f $X=2.69 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A1_M1001_g N_B1_M1010_g 0.0272015f $X=2.71 $Y=2.465 $X2=0 $Y2=0
cc_174 A1 B1 0.020065f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A1_c_224_n B1 4.13251e-19 $X=2.69 $Y=1.36 $X2=0 $Y2=0
cc_176 A1 N_B1_c_259_n 0.0181378f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A1_c_224_n N_B1_c_259_n 0.0222349f $X=2.69 $Y=1.36 $X2=0 $Y2=0
cc_178 N_A1_M1001_g N_VPWR_c_283_n 0.0100448f $X=2.71 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A1_M1001_g N_VPWR_c_288_n 0.00549284f $X=2.71 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A1_M1001_g N_VPWR_c_279_n 0.010487f $X=2.71 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A1_M1001_g N_A_342_367#_c_361_n 0.00109181f $X=2.71 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A1_M1001_g N_A_342_367#_c_358_n 0.0124105f $X=2.71 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A1_M1001_g N_A_342_367#_c_359_n 7.54694e-19 $X=2.71 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A1_M1001_g N_A_342_367#_c_363_n 0.0121839f $X=2.71 $Y=2.465 $X2=0 $Y2=0
cc_185 A1 N_VGND_c_382_n 0.00183598f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A1_c_225_n N_VGND_c_382_n 0.00101452f $X=2.69 $Y=1.195 $X2=0 $Y2=0
cc_187 N_A1_c_225_n N_VGND_c_383_n 0.00575161f $X=2.69 $Y=1.195 $X2=0 $Y2=0
cc_188 N_A1_c_225_n N_VGND_c_387_n 0.00697924f $X=2.69 $Y=1.195 $X2=0 $Y2=0
cc_189 N_B1_M1010_g N_VPWR_c_288_n 0.00549284f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_190 N_B1_M1010_g N_VPWR_c_279_n 0.0110256f $X=3.14 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B1_M1010_g N_A_342_367#_c_359_n 0.00227309f $X=3.14 $Y=2.465 $X2=0
+ $Y2=0
cc_192 N_B1_M1010_g N_A_342_367#_c_363_n 0.00943908f $X=3.14 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_B1_c_256_n N_VGND_c_382_n 0.0175156f $X=3.14 $Y=1.195 $X2=0 $Y2=0
cc_194 B1 N_VGND_c_382_n 0.0111342f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_195 N_B1_c_259_n N_VGND_c_382_n 0.00769708f $X=3.47 $Y=1.36 $X2=0 $Y2=0
cc_196 N_B1_c_256_n N_VGND_c_383_n 0.00477554f $X=3.14 $Y=1.195 $X2=0 $Y2=0
cc_197 N_B1_c_256_n N_VGND_c_387_n 0.0085718f $X=3.14 $Y=1.195 $X2=0 $Y2=0
cc_198 N_VPWR_c_279_n N_X_M1002_s 0.00223819f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_281_n X 0.0950581f $X=0.37 $Y=1.99 $X2=0 $Y2=0
cc_200 N_VPWR_c_284_n X 0.0232928f $X=1.22 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VPWR_c_279_n X 0.0152794f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_c_279_n N_A_342_367#_M1003_d 0.00258346f $X=3.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_203 N_VPWR_c_279_n N_A_342_367#_M1001_d 0.00223819f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_283_n N_A_342_367#_c_361_n 0.0412283f $X=2.39 $Y=2.57 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_286_n N_A_342_367#_c_361_n 0.0169299f $X=2.225 $Y=3.33 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_279_n N_A_342_367#_c_361_n 0.0112082f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_207 N_VPWR_M1005_d N_A_342_367#_c_358_n 0.0111512f $X=2.14 $Y=1.835 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_283_n N_A_342_367#_c_358_n 0.0221174f $X=2.39 $Y=2.57 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_283_n N_A_342_367#_c_363_n 0.0416706f $X=2.39 $Y=2.57 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_288_n N_A_342_367#_c_363_n 0.0177952f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_211 N_VPWR_c_279_n N_A_342_367#_c_363_n 0.0123247f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_212 N_X_c_330_n N_VGND_c_381_n 0.0322421f $X=0.715 $Y=1.125 $X2=0 $Y2=0
cc_213 N_X_c_352_p N_VGND_c_385_n 0.0124525f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_214 N_X_M1008_s N_VGND_c_387_n 0.00536646f $X=0.575 $Y=0.245 $X2=0 $Y2=0
cc_215 N_X_c_352_p N_VGND_c_387_n 0.00730901f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_216 N_VGND_c_387_n A_355_49# 0.00312872f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_217 N_VGND_c_387_n A_427_49# 0.00581048f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
