* File: sky130_fd_sc_lp__einvn_m.pxi.spice
* Created: Fri Aug 28 10:33:26 2020
* 
x_PM_SKY130_FD_SC_LP__EINVN_M%TE_B N_TE_B_M1004_g N_TE_B_c_43_n N_TE_B_M1002_g
+ N_TE_B_c_44_n N_TE_B_c_45_n N_TE_B_M1005_g N_TE_B_c_46_n TE_B TE_B
+ N_TE_B_c_41_n PM_SKY130_FD_SC_LP__EINVN_M%TE_B
x_PM_SKY130_FD_SC_LP__EINVN_M%A_47_154# N_A_47_154#_M1004_s N_A_47_154#_M1002_s
+ N_A_47_154#_M1000_g N_A_47_154#_c_84_n N_A_47_154#_c_89_n N_A_47_154#_c_85_n
+ N_A_47_154#_c_86_n N_A_47_154#_c_87_n N_A_47_154#_c_88_n
+ PM_SKY130_FD_SC_LP__EINVN_M%A_47_154#
x_PM_SKY130_FD_SC_LP__EINVN_M%A N_A_M1001_g N_A_M1003_g N_A_c_128_n N_A_c_129_n
+ N_A_c_133_n A N_A_c_131_n PM_SKY130_FD_SC_LP__EINVN_M%A
x_PM_SKY130_FD_SC_LP__EINVN_M%VPWR N_VPWR_M1002_d N_VPWR_c_160_n VPWR
+ N_VPWR_c_161_n N_VPWR_c_159_n N_VPWR_c_163_n PM_SKY130_FD_SC_LP__EINVN_M%VPWR
x_PM_SKY130_FD_SC_LP__EINVN_M%Z N_Z_M1001_d N_Z_M1003_d Z Z Z Z Z N_Z_c_187_n
+ PM_SKY130_FD_SC_LP__EINVN_M%Z
x_PM_SKY130_FD_SC_LP__EINVN_M%VGND N_VGND_M1004_d N_VGND_c_205_n N_VGND_c_213_n
+ N_VGND_c_206_n N_VGND_c_207_n VGND N_VGND_c_208_n N_VGND_c_209_n
+ PM_SKY130_FD_SC_LP__EINVN_M%VGND
cc_1 VNB N_TE_B_M1004_g 0.0370475f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.98
cc_2 VNB TE_B 0.0294652f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_3 VNB N_TE_B_c_41_n 0.0422408f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.495
cc_4 VNB N_A_47_154#_M1000_g 0.0296962f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=2.49
cc_5 VNB N_A_47_154#_c_84_n 0.0277154f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_6 VNB N_A_47_154#_c_85_n 0.00356353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_47_154#_c_86_n 0.0054421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_47_154#_c_87_n 2.38365e-19 $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.507
cc_9 VNB N_A_47_154#_c_88_n 0.013555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_M1001_g 0.0179861f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.98
cc_11 VNB N_A_c_128_n 0.0124135f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=2.885
cc_12 VNB N_A_c_129_n 0.015018f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=2.885
cc_13 VNB A 0.0233039f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_14 VNB N_A_c_131_n 0.0440658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_159_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_16 VNB N_Z_c_187_n 0.0323695f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.495
cc_17 VNB N_VGND_c_205_n 0.0150397f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.565
cc_18 VNB N_VGND_c_206_n 0.0278122f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=2.885
cc_19 VNB N_VGND_c_207_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.49
cc_20 VNB N_VGND_c_208_n 0.0216928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_209_n 0.147325f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.66
cc_22 VPB N_TE_B_M1004_g 0.0522719f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.98
cc_23 VPB N_TE_B_c_43_n 0.0190688f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.565
cc_24 VPB N_TE_B_c_44_n 0.0236093f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=2.49
cc_25 VPB N_TE_B_c_45_n 0.0155381f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=2.565
cc_26 VPB N_TE_B_c_46_n 0.0151318f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.49
cc_27 VPB N_A_47_154#_c_89_n 0.0555612f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.495
cc_28 VPB N_A_47_154#_c_85_n 0.00721425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_A_47_154#_c_86_n 0.00226754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_A_47_154#_c_87_n 0.00182907f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.507
cc_31 VPB N_A_47_154#_c_88_n 0.0427471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_c_129_n 0.0526147f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=2.885
cc_33 VPB N_A_c_133_n 0.0317244f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.49
cc_34 VPB N_VPWR_c_160_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=1.01 $Y2=2.49
cc_35 VPB N_VPWR_c_161_n 0.0269588f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.47
cc_36 VPB N_VPWR_c_159_n 0.0493638f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_37 VPB N_VPWR_c_163_n 0.0252934f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.495
cc_38 VPB N_Z_c_187_n 0.051605f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.495
cc_39 TE_B N_A_47_154#_M1000_g 3.13445e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_40 N_TE_B_c_41_n N_A_47_154#_M1000_g 0.0229342f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_41 N_TE_B_M1004_g N_A_47_154#_c_84_n 0.0170491f $X=0.575 $Y=0.98 $X2=0 $Y2=0
cc_42 TE_B N_A_47_154#_c_84_n 0.0253281f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_43 N_TE_B_c_41_n N_A_47_154#_c_84_n 0.00116678f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_44 N_TE_B_M1004_g N_A_47_154#_c_89_n 0.0309586f $X=0.575 $Y=0.98 $X2=0 $Y2=0
cc_45 N_TE_B_c_43_n N_A_47_154#_c_89_n 0.00458376f $X=0.655 $Y=2.565 $X2=0 $Y2=0
cc_46 N_TE_B_c_46_n N_A_47_154#_c_89_n 0.0107758f $X=0.615 $Y=2.49 $X2=0 $Y2=0
cc_47 N_TE_B_M1004_g N_A_47_154#_c_85_n 0.0144354f $X=0.575 $Y=0.98 $X2=0 $Y2=0
cc_48 N_TE_B_M1004_g N_A_47_154#_c_86_n 0.00383478f $X=0.575 $Y=0.98 $X2=0 $Y2=0
cc_49 N_TE_B_M1004_g N_A_47_154#_c_87_n 0.00146961f $X=0.575 $Y=0.98 $X2=0 $Y2=0
cc_50 N_TE_B_c_44_n N_A_47_154#_c_87_n 0.00103702f $X=1.01 $Y=2.49 $X2=0 $Y2=0
cc_51 N_TE_B_M1004_g N_A_47_154#_c_88_n 0.0408314f $X=0.575 $Y=0.98 $X2=0 $Y2=0
cc_52 N_TE_B_c_44_n N_A_47_154#_c_88_n 0.0214535f $X=1.01 $Y=2.49 $X2=0 $Y2=0
cc_53 N_TE_B_c_41_n N_A_M1001_g 4.92795e-19 $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_54 N_TE_B_c_44_n N_A_c_133_n 0.0257604f $X=1.01 $Y=2.49 $X2=0 $Y2=0
cc_55 N_TE_B_c_45_n N_A_c_133_n 0.0257604f $X=1.085 $Y=2.565 $X2=0 $Y2=0
cc_56 N_TE_B_c_41_n N_A_c_131_n 0.002845f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_57 N_TE_B_c_43_n N_VPWR_c_160_n 0.0119415f $X=0.655 $Y=2.565 $X2=0 $Y2=0
cc_58 N_TE_B_c_44_n N_VPWR_c_160_n 0.00354254f $X=1.01 $Y=2.49 $X2=0 $Y2=0
cc_59 N_TE_B_c_45_n N_VPWR_c_160_n 0.00955773f $X=1.085 $Y=2.565 $X2=0 $Y2=0
cc_60 N_TE_B_c_45_n N_VPWR_c_161_n 0.00486043f $X=1.085 $Y=2.565 $X2=0 $Y2=0
cc_61 N_TE_B_c_43_n N_VPWR_c_159_n 0.00950102f $X=0.655 $Y=2.565 $X2=0 $Y2=0
cc_62 N_TE_B_c_45_n N_VPWR_c_159_n 0.00818711f $X=1.085 $Y=2.565 $X2=0 $Y2=0
cc_63 N_TE_B_c_46_n N_VPWR_c_159_n 0.0014965f $X=0.615 $Y=2.49 $X2=0 $Y2=0
cc_64 N_TE_B_c_43_n N_VPWR_c_163_n 0.00486043f $X=0.655 $Y=2.565 $X2=0 $Y2=0
cc_65 N_TE_B_c_46_n N_VPWR_c_163_n 0.00116881f $X=0.615 $Y=2.49 $X2=0 $Y2=0
cc_66 N_TE_B_c_44_n N_Z_c_187_n 0.00248279f $X=1.01 $Y=2.49 $X2=0 $Y2=0
cc_67 N_TE_B_M1004_g N_VGND_c_205_n 9.01787e-19 $X=0.575 $Y=0.98 $X2=0 $Y2=0
cc_68 TE_B N_VGND_c_205_n 0.0285297f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_69 N_TE_B_c_41_n N_VGND_c_205_n 9.09245e-19 $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_70 TE_B N_VGND_c_213_n 0.00837641f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_71 TE_B N_VGND_c_206_n 0.0313238f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_72 N_TE_B_c_41_n N_VGND_c_206_n 0.00735687f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_73 TE_B N_VGND_c_209_n 0.0253668f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_74 N_TE_B_c_41_n N_VGND_c_209_n 0.0106807f $X=0.485 $Y=0.495 $X2=0 $Y2=0
cc_75 N_A_47_154#_M1000_g N_A_M1001_g 0.0330743f $X=1.015 $Y=0.98 $X2=0 $Y2=0
cc_76 N_A_47_154#_M1000_g N_A_c_129_n 0.00485776f $X=1.015 $Y=0.98 $X2=0 $Y2=0
cc_77 N_A_47_154#_c_87_n N_A_c_129_n 0.00192681f $X=1.025 $Y=1.7 $X2=0 $Y2=0
cc_78 N_A_47_154#_c_88_n N_A_c_129_n 0.039754f $X=1.025 $Y=1.7 $X2=0 $Y2=0
cc_79 N_A_47_154#_c_87_n N_VPWR_c_160_n 0.00179539f $X=1.025 $Y=1.7 $X2=0 $Y2=0
cc_80 N_A_47_154#_c_88_n N_VPWR_c_160_n 5.02403e-19 $X=1.025 $Y=1.7 $X2=0 $Y2=0
cc_81 N_A_47_154#_M1002_s N_VPWR_c_159_n 0.0028801f $X=0.315 $Y=2.675 $X2=0
+ $Y2=0
cc_82 N_A_47_154#_c_89_n N_VPWR_c_159_n 0.012144f $X=0.44 $Y=2.82 $X2=0 $Y2=0
cc_83 N_A_47_154#_c_89_n N_VPWR_c_163_n 0.0146615f $X=0.44 $Y=2.82 $X2=0 $Y2=0
cc_84 N_A_47_154#_M1000_g N_Z_c_187_n 0.00205238f $X=1.015 $Y=0.98 $X2=0 $Y2=0
cc_85 N_A_47_154#_c_87_n N_Z_c_187_n 0.0254669f $X=1.025 $Y=1.7 $X2=0 $Y2=0
cc_86 N_A_47_154#_c_88_n N_Z_c_187_n 0.00212006f $X=1.025 $Y=1.7 $X2=0 $Y2=0
cc_87 N_A_47_154#_M1000_g N_VGND_c_205_n 0.00871701f $X=1.015 $Y=0.98 $X2=0
+ $Y2=0
cc_88 N_A_47_154#_M1000_g N_VGND_c_213_n 0.0107469f $X=1.015 $Y=0.98 $X2=0 $Y2=0
cc_89 N_A_47_154#_c_85_n N_VGND_c_213_n 0.00942199f $X=0.94 $Y=1.62 $X2=0 $Y2=0
cc_90 N_A_47_154#_c_87_n N_VGND_c_213_n 0.00713418f $X=1.025 $Y=1.7 $X2=0 $Y2=0
cc_91 N_A_47_154#_c_88_n N_VGND_c_213_n 0.00265109f $X=1.025 $Y=1.7 $X2=0 $Y2=0
cc_92 N_A_47_154#_M1000_g N_VGND_c_206_n 0.00103255f $X=1.015 $Y=0.98 $X2=0
+ $Y2=0
cc_93 N_A_47_154#_M1000_g N_VGND_c_209_n 0.00132218f $X=1.015 $Y=0.98 $X2=0
+ $Y2=0
cc_94 N_A_c_133_n N_VPWR_c_160_n 0.00220193f $X=1.46 $Y=2.565 $X2=0 $Y2=0
cc_95 N_A_c_133_n N_VPWR_c_161_n 0.00553654f $X=1.46 $Y=2.565 $X2=0 $Y2=0
cc_96 N_A_c_133_n N_VPWR_c_159_n 0.010948f $X=1.46 $Y=2.565 $X2=0 $Y2=0
cc_97 N_A_M1001_g N_Z_c_187_n 0.00782799f $X=1.445 $Y=0.98 $X2=0 $Y2=0
cc_98 N_A_c_128_n N_Z_c_187_n 0.00668002f $X=1.46 $Y=1.415 $X2=0 $Y2=0
cc_99 N_A_c_129_n N_Z_c_187_n 0.0429225f $X=1.46 $Y=2.415 $X2=0 $Y2=0
cc_100 N_A_c_133_n N_Z_c_187_n 0.0152489f $X=1.46 $Y=2.565 $X2=0 $Y2=0
cc_101 A N_Z_c_187_n 0.0249411f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_102 N_A_c_131_n N_Z_c_187_n 4.67739e-19 $X=1.465 $Y=0.42 $X2=0 $Y2=0
cc_103 N_A_M1001_g N_VGND_c_205_n 0.00367955f $X=1.445 $Y=0.98 $X2=0 $Y2=0
cc_104 A N_VGND_c_205_n 0.0337552f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_105 N_A_c_131_n N_VGND_c_205_n 0.00449261f $X=1.465 $Y=0.42 $X2=0 $Y2=0
cc_106 N_A_M1001_g N_VGND_c_213_n 0.00255365f $X=1.445 $Y=0.98 $X2=0 $Y2=0
cc_107 A N_VGND_c_208_n 0.0327149f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_108 N_A_c_131_n N_VGND_c_208_n 0.00813345f $X=1.465 $Y=0.42 $X2=0 $Y2=0
cc_109 A N_VGND_c_209_n 0.0186382f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_110 N_A_c_131_n N_VGND_c_209_n 0.011167f $X=1.465 $Y=0.42 $X2=0 $Y2=0
cc_111 N_VPWR_c_159_n A_232_535# 0.00899413f $X=1.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_112 N_VPWR_c_159_n N_Z_M1003_d 0.00235821f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_113 N_VPWR_c_160_n N_Z_c_187_n 0.00267659f $X=0.87 $Y=2.95 $X2=0 $Y2=0
cc_114 N_VPWR_c_161_n N_Z_c_187_n 0.010662f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_115 N_VPWR_c_159_n N_Z_c_187_n 0.0115728f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_116 N_Z_c_187_n N_VGND_c_213_n 0.015402f $X=1.66 $Y=1.02 $X2=0 $Y2=0
cc_117 N_Z_c_187_n N_VGND_c_209_n 9.13886e-19 $X=1.66 $Y=1.02 $X2=0 $Y2=0
cc_118 N_VGND_c_205_n A_218_154# 0.00103787f $X=1.07 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_119 N_VGND_c_213_n A_218_154# 0.00395355f $X=1.07 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
