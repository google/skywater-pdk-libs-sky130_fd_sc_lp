* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a311o_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 a_72_312# C1 a_558_486# VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=1.344e+11p ps=1.7e+06u
M1001 a_72_312# A1 a_330_48# VNB nshort w=420000u l=150000u
+  ad=3.507e+11p pd=3.35e+06u as=1.638e+11p ps=1.62e+06u
M1002 a_558_486# B1 a_224_486# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.84e+11p ps=3.76e+06u
M1003 a_72_312# C1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.814e+11p ps=3.02e+06u
M1004 VPWR a_72_312# X VPB phighvt w=640000u l=150000u
+  ad=5.76e+11p pd=4.36e+06u as=1.824e+11p ps=1.85e+06u
M1005 VPWR A2 a_224_486# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_72_312# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 a_224_486# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_224_486# A3 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_330_48# A2 a_246_48# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1010 VGND B1 a_72_312# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_246_48# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
