* File: sky130_fd_sc_lp__dlygate4s18_1.spice
* Created: Fri Aug 28 10:30:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlygate4s18_1.pex.spice"
.subckt sky130_fd_sc_lp__dlygate4s18_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_27_52#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1491 AS=0.1113 PD=1.13 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_A_288_52#_M1000_d N_A_27_52#_M1000_g N_VGND_M1005_d VNB NSHORT L=0.18
+ W=0.42 AD=0.1113 AS=0.1491 PD=1.37 PS=1.13 NRD=0 NRS=107.136 M=1 R=2.33333
+ SA=90001 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1006 N_VGND_M1006_d N_A_288_52#_M1006_g N_A_405_136#_M1006_s VNB NSHORT L=0.18
+ W=0.42 AD=0.1295 AS=0.1113 PD=1 PS=1.37 NRD=109.992 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001 A=0.0756 P=1.2 MULT=1
MM1001 N_X_M1001_d N_A_405_136#_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.259 PD=2.21 PS=2 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_27_52#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1491 AS=0.1113 PD=1.13 PS=1.37 NRD=21.0987 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_A_288_52#_M1004_d N_A_27_52#_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1113 AS=0.1491 PD=1.37 PS=1.13 NRD=0 NRS=180.57 M=1 R=2.33333
+ SA=90001 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_288_52#_M1007_g N_A_405_136#_M1007_s VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.12495 AS=0.1113 PD=0.96 PS=1.37 NRD=180.57 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001 A=0.0756 P=1.2 MULT=1
MM1002 N_X_M1002_d N_A_405_136#_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.37485 PD=3.05 PS=2.88 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_35 VNB 0 1.65637e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dlygate4s18_1.pxi.spice"
*
.ends
*
*
