* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VPWR A2 a_819_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND A2 a_1201_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Y D1 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 Y C1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_819_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_454_367# B1 a_819_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_819_367# B1 a_454_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_27_367# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_819_367# B1 a_454_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_1201_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_27_367# C1 a_454_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_819_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 Y A1 a_1201_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_27_367# D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 Y D1 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_1201_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_1201_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_819_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_454_367# B1 a_819_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VPWR A2 a_819_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 a_27_367# C1 a_454_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_454_367# C1 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_1201_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 VPWR A1 a_819_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_819_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 Y A1 a_1201_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 VGND A2 a_1201_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 VPWR A1 a_819_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 Y D1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X37 VGND D1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 a_454_367# C1 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
