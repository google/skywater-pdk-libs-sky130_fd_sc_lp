* File: sky130_fd_sc_lp__o2111ai_1.pex.spice
* Created: Wed Sep  2 10:13:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111AI_1%D1 3 6 8 9 13 15
r29 13 16 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.73 $Y=1.35
+ $X2=0.73 $Y2=1.515
r30 13 15 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.73 $Y=1.35
+ $X2=0.73 $Y2=1.185
r31 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.35 $X2=0.72 $Y2=1.35
r32 8 9 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.747 $Y=0.925
+ $X2=0.747 $Y2=1.295
r33 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.83 $Y=2.465
+ $X2=0.83 $Y2=1.515
r34 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.83 $Y=0.655
+ $X2=0.83 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_1%C1 3 6 8 9 10 15 17
c36 8 0 1.48545e-19 $X=1.2 $Y=0.555
c37 6 0 1.09784e-19 $X=1.37 $Y=2.465
r38 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.28 $Y=1.35
+ $X2=1.28 $Y2=1.515
r39 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.28 $Y=1.35
+ $X2=1.28 $Y2=1.185
r40 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.28
+ $Y=1.35 $X2=1.28 $Y2=1.35
r41 9 10 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.21 $Y=0.925 $X2=1.21
+ $Y2=1.295
r42 8 9 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.21 $Y=0.555 $X2=1.21
+ $Y2=0.925
r43 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.37 $Y=2.465
+ $X2=1.37 $Y2=1.515
r44 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.27 $Y=0.655
+ $X2=1.27 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_1%B1 3 7 9 15 16
c32 16 0 1.48545e-19 $X=1.92 $Y=1.51
c33 15 0 5.94326e-20 $X=1.82 $Y=1.51
r34 14 16 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.82 $Y=1.51 $X2=1.92
+ $Y2=1.51
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.51 $X2=1.82 $Y2=1.51
r36 11 14 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.73 $Y=1.51 $X2=1.82
+ $Y2=1.51
r37 9 15 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.72 $Y2=1.51
r38 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.675
+ $X2=1.92 $Y2=1.51
r39 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.92 $Y=1.675 $X2=1.92
+ $Y2=2.465
r40 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.345
+ $X2=1.73 $Y2=1.51
r41 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.73 $Y=1.345 $X2=1.73
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_1%A2 3 7 9 10 18
c31 7 0 5.94326e-20 $X=2.49 $Y=2.465
r32 16 18 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.4 $Y=1.51 $X2=2.49
+ $Y2=1.51
r33 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=1.51 $X2=2.4 $Y2=1.51
r34 13 16 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.28 $Y=1.51 $X2=2.4
+ $Y2=1.51
r35 10 17 6.66473 $w=4.13e-07 $l=2.4e-07 $layer=LI1_cond $X=2.64 $Y=1.552
+ $X2=2.4 $Y2=1.552
r36 9 17 6.66473 $w=4.13e-07 $l=2.4e-07 $layer=LI1_cond $X=2.16 $Y=1.552 $X2=2.4
+ $Y2=1.552
r37 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=1.675
+ $X2=2.49 $Y2=1.51
r38 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.49 $Y=1.675 $X2=2.49
+ $Y2=2.465
r39 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.345
+ $X2=2.28 $Y2=1.51
r40 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.28 $Y=1.345 $X2=2.28
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_1%A1 3 7 9 14 15
r24 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.46 $X2=3.07 $Y2=1.46
r25 11 14 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.85 $Y=1.46
+ $X2=3.07 $Y2=1.46
r26 9 15 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.07 $Y=1.665
+ $X2=3.07 $Y2=1.46
r27 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.625
+ $X2=2.85 $Y2=1.46
r28 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.85 $Y=1.625 $X2=2.85
+ $Y2=2.465
r29 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.295
+ $X2=2.85 $Y2=1.46
r30 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.85 $Y=1.295 $X2=2.85
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_1%VPWR 1 2 3 12 18 20 22 27 28 29 35 39 45
+ 49
r41 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 43 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 40 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.645 $Y2=3.33
r45 40 42 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 39 48 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.9 $Y=3.33 $X2=3.13
+ $Y2=3.33
r47 39 42 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=3.33 $X2=2.64
+ $Y2=3.33
r48 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 35 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=3.33
+ $X2=1.645 $Y2=3.33
r50 35 37 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.48 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 33 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 29 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 29 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 29 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 27 32 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.43 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 27 28 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.43 $Y=3.33
+ $X2=0.605 $Y2=3.33
r58 26 37 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.78 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 26 28 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.78 $Y=3.33
+ $X2=0.605 $Y2=3.33
r60 22 25 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=3.065 $Y=2.01
+ $X2=3.065 $Y2=2.95
r61 20 48 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.13 $Y2=3.33
r62 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.065 $Y2=2.95
r63 16 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=3.245
+ $X2=1.645 $Y2=3.33
r64 16 18 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=1.645 $Y=3.245
+ $X2=1.645 $Y2=2.435
r65 12 15 25.3537 $w=3.48e-07 $l=7.7e-07 $layer=LI1_cond $X=0.605 $Y=2.18
+ $X2=0.605 $Y2=2.95
r66 10 28 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=3.245
+ $X2=0.605 $Y2=3.33
r67 10 15 9.71345 $w=3.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.605 $Y=3.245
+ $X2=0.605 $Y2=2.95
r68 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.835 $X2=3.065 $Y2=2.95
r69 3 22 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.835 $X2=3.065 $Y2=2.01
r70 2 18 300 $w=1.7e-07 $l=6.9282e-07 $layer=licon1_PDIFF $count=2 $X=1.445
+ $Y=1.835 $X2=1.645 $Y2=2.435
r71 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.49
+ $Y=1.835 $X2=0.615 $Y2=2.95
r72 1 12 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.49
+ $Y=1.835 $X2=0.615 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_1%Y 1 2 3 13 14 15 16 18 20 23 28 29 30 51
c44 14 0 1.09784e-19 $X=0.95 $Y=1.805
r45 51 52 2.26693 $w=4.13e-07 $l=6.5e-08 $layer=LI1_cond $X=1.157 $Y=2.035
+ $X2=1.157 $Y2=2.1
r46 47 48 0.97194 $w=4.13e-07 $l=3.5e-08 $layer=LI1_cond $X=1.157 $Y=1.98
+ $X2=1.157 $Y2=2.015
r47 30 40 11.3524 $w=3.33e-07 $l=3.3e-07 $layer=LI1_cond $X=1.117 $Y=2.775
+ $X2=1.117 $Y2=2.445
r48 29 40 1.37605 $w=3.33e-07 $l=4e-08 $layer=LI1_cond $X=1.117 $Y=2.405
+ $X2=1.117 $Y2=2.445
r49 28 51 0.277697 $w=4.13e-07 $l=1e-08 $layer=LI1_cond $X=1.157 $Y=2.025
+ $X2=1.157 $Y2=2.035
r50 28 48 0.277697 $w=4.13e-07 $l=1e-08 $layer=LI1_cond $X=1.157 $Y=2.025
+ $X2=1.157 $Y2=2.015
r51 28 29 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=1.117 $Y=2.11
+ $X2=1.117 $Y2=2.405
r52 28 52 0.344013 $w=3.33e-07 $l=1e-08 $layer=LI1_cond $X=1.117 $Y=2.11
+ $X2=1.117 $Y2=2.1
r53 18 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.1 $X2=2.2
+ $Y2=2.015
r54 18 20 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.2 $Y=2.1 $X2=2.2
+ $Y2=2.485
r55 17 48 6.00275 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=1.365 $Y=2.015
+ $X2=1.157 $Y2=2.015
r56 16 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=2.015
+ $X2=2.2 $Y2=2.015
r57 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.035 $Y=2.015
+ $X2=1.365 $Y2=2.015
r58 14 47 4.8597 $w=4.13e-07 $l=1.75e-07 $layer=LI1_cond $X=1.157 $Y=1.805
+ $X2=1.157 $Y2=1.98
r59 14 15 24.4894 $w=2.38e-07 $l=5.1e-07 $layer=LI1_cond $X=0.95 $Y=1.805
+ $X2=0.44 $Y2=1.805
r60 11 15 7.03987 $w=2.4e-07 $l=2.16852e-07 $layer=LI1_cond $X=0.275 $Y=1.685
+ $X2=0.44 $Y2=1.805
r61 11 13 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.275 $Y=1.685
+ $X2=0.275 $Y2=0.93
r62 10 23 2.08194 $w=3.3e-07 $l=2.08e-07 $layer=LI1_cond $X=0.275 $Y=0.67
+ $X2=0.275 $Y2=0.462
r63 10 13 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.275 $Y=0.67
+ $X2=0.275 $Y2=0.93
r64 3 27 600 $w=1.7e-07 $l=2.80936e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.835 $X2=2.2 $Y2=2.015
r65 3 20 300 $w=1.7e-07 $l=7.45486e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.835 $X2=2.2 $Y2=2.485
r66 2 47 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.835 $X2=1.1 $Y2=1.98
r67 2 40 300 $w=1.7e-07 $l=7.0075e-07 $layer=licon1_PDIFF $count=2 $X=0.905
+ $Y=1.835 $X2=1.1 $Y2=2.445
r68 1 23 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.42
r69 1 13 182 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_1%A_361_47# 1 2 9 11 12 15
r24 13 15 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=3.065 $Y=1.005
+ $X2=3.065 $Y2=0.42
r25 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.9 $Y=1.09
+ $X2=3.065 $Y2=1.005
r26 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.9 $Y=1.09 $X2=2.17
+ $Y2=1.09
r27 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.005 $Y=1.005
+ $X2=2.17 $Y2=1.09
r28 7 9 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=2.005 $Y=1.005
+ $X2=2.005 $Y2=0.42
r29 2 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.925
+ $Y=0.235 $X2=3.065 $Y2=0.42
r30 1 9 91 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_NDIFF $count=2 $X=1.805
+ $Y=0.235 $X2=2.005 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_1%VGND 1 6 8 10 20 21 24
r33 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r34 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r35 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r36 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=0 $X2=2.565
+ $Y2=0
r37 18 20 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.73 $Y=0 $X2=3.12
+ $Y2=0
r38 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r39 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r40 12 16 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r41 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r42 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.565
+ $Y2=0
r43 10 16 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r44 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r45 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r46 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=0.085
+ $X2=2.565 $Y2=0
r47 4 6 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.565 $Y=0.085
+ $X2=2.565 $Y2=0.36
r48 1 6 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=2.355
+ $Y=0.235 $X2=2.565 $Y2=0.36
.ends

