* File: sky130_fd_sc_lp__a31oi_1.pex.spice
* Created: Wed Sep  2 09:26:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31OI_1%A3 3 7 9 10 17
r29 14 17 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.46 $Y=1.375
+ $X2=0.68 $Y2=1.375
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.46
+ $Y=1.375 $X2=0.46 $Y2=1.375
r31 10 15 7.54049 $w=4.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=1.375
r32 9 15 2.08014 $w=4.58e-07 $l=8e-08 $layer=LI1_cond $X=0.315 $Y=1.295
+ $X2=0.315 $Y2=1.375
r33 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.68 $Y=1.54
+ $X2=0.68 $Y2=1.375
r34 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.68 $Y=1.54 $X2=0.68
+ $Y2=2.465
r35 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.68 $Y=1.21
+ $X2=0.68 $Y2=1.375
r36 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.68 $Y=1.21 $X2=0.68
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_1%A2 3 6 8 9 13 15
r36 13 16 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.35
+ $X2=1.135 $Y2=1.515
r37 13 15 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.35
+ $X2=1.135 $Y2=1.185
r38 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.35 $X2=1.14 $Y2=1.35
r39 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.925 $X2=1.2
+ $Y2=1.295
r40 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.11 $Y=2.465
+ $X2=1.11 $Y2=1.515
r41 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.04 $Y=0.655
+ $X2=1.04 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_1%A1 3 6 8 11 13
r35 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.35
+ $X2=1.68 $Y2=1.515
r36 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.35
+ $X2=1.68 $Y2=1.185
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.35 $X2=1.68 $Y2=1.35
r38 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.7 $Y=2.465 $X2=1.7
+ $Y2=1.515
r39 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.59 $Y=0.655
+ $X2=1.59 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_1%B1 1 3 6 9 10 13
r24 10 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.56
+ $Y=1.35 $X2=2.56 $Y2=1.35
r25 8 13 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.205 $Y=1.35
+ $X2=2.56 $Y2=1.35
r26 8 9 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.205 $Y=1.35 $X2=2.13
+ $Y2=1.35
r27 4 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.515
+ $X2=2.13 $Y2=1.35
r28 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.13 $Y=1.515 $X2=2.13
+ $Y2=2.465
r29 1 9 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.185
+ $X2=2.13 $Y2=1.35
r30 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.13 $Y=1.185 $X2=2.13
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_1%VPWR 1 2 9 15 18 19 21 22 23 35 36
r34 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r37 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r39 27 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 23 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 23 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r43 21 29 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=3.33
+ $X2=1.405 $Y2=3.33
r45 20 32 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=1.405 $Y2=3.33
r47 18 26 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=0.3 $Y=3.33 $X2=0.24
+ $Y2=3.33
r48 18 19 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.3 $Y=3.33 $X2=0.43
+ $Y2=3.33
r49 17 29 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 17 19 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.43
+ $Y2=3.33
r51 13 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.405 $Y=3.245
+ $X2=1.405 $Y2=3.33
r52 13 15 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=1.405 $Y=3.245
+ $X2=1.405 $Y2=2.45
r53 9 12 37.0112 $w=2.58e-07 $l=8.35e-07 $layer=LI1_cond $X=0.43 $Y=2.115
+ $X2=0.43 $Y2=2.95
r54 7 19 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.43 $Y=3.245
+ $X2=0.43 $Y2=3.33
r55 7 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.43 $Y=3.245
+ $X2=0.43 $Y2=2.95
r56 2 15 300 $w=1.7e-07 $l=7.16607e-07 $layer=licon1_PDIFF $count=2 $X=1.185
+ $Y=1.835 $X2=1.405 $Y2=2.45
r57 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.34
+ $Y=1.835 $X2=0.465 $Y2=2.95
r58 1 9 400 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_PDIFF $count=1 $X=0.34
+ $Y=1.835 $X2=0.465 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_1%A_151_367# 1 2 7 9 11 13 15
r27 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=2.195
+ $X2=1.915 $Y2=2.11
r28 13 15 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=1.915 $Y=2.195
+ $X2=1.915 $Y2=2.95
r29 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=2.11
+ $X2=0.895 $Y2=2.11
r30 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.75 $Y=2.11
+ $X2=1.915 $Y2=2.11
r31 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.75 $Y=2.11 $X2=1.06
+ $Y2=2.11
r32 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=2.195
+ $X2=0.895 $Y2=2.11
r33 7 9 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.895 $Y=2.195
+ $X2=0.895 $Y2=2.95
r34 2 20 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.775
+ $Y=1.835 $X2=1.915 $Y2=2.11
r35 2 15 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.775
+ $Y=1.835 $X2=1.915 $Y2=2.95
r36 1 18 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=1.835 $X2=0.895 $Y2=2.11
r37 1 9 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.755
+ $Y=1.835 $X2=0.895 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_1%Y 1 2 8 9 10 11 12 16 18 19 20 25
r57 20 33 2.96276 $w=5.43e-07 $l=1.35e-07 $layer=LI1_cond $X=2.522 $Y=2.775
+ $X2=2.522 $Y2=2.91
r58 19 20 8.12016 $w=5.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.522 $Y=2.405
+ $X2=2.522 $Y2=2.775
r59 18 19 8.12016 $w=5.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.522 $Y=2.035
+ $X2=2.522 $Y2=2.405
r60 18 25 1.20705 $w=5.43e-07 $l=5.5e-08 $layer=LI1_cond $X=2.522 $Y=2.035
+ $X2=2.522 $Y2=1.98
r61 17 25 2.7433 $w=5.43e-07 $l=1.25e-07 $layer=LI1_cond $X=2.522 $Y=1.855
+ $X2=2.522 $Y2=1.98
r62 11 17 9.60392 $w=1.7e-07 $l=3.11615e-07 $layer=LI1_cond $X=2.25 $Y=1.77
+ $X2=2.522 $Y2=1.855
r63 11 12 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=2.25 $Y=1.77
+ $X2=0.885 $Y2=1.77
r64 9 16 4.04406 $w=2.75e-07 $l=1.87e-07 $layer=LI1_cond $X=1.635 $Y=0.392
+ $X2=1.822 $Y2=0.392
r65 9 10 31.4303 $w=2.73e-07 $l=7.5e-07 $layer=LI1_cond $X=1.635 $Y=0.392
+ $X2=0.885 $Y2=0.392
r66 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.8 $Y=1.685
+ $X2=0.885 $Y2=1.77
r67 7 10 7.32204 $w=2.75e-07 $l=1.75425e-07 $layer=LI1_cond $X=0.8 $Y=0.53
+ $X2=0.885 $Y2=0.392
r68 7 8 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=0.8 $Y=0.53 $X2=0.8
+ $Y2=1.685
r69 2 33 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.205
+ $Y=1.835 $X2=2.345 $Y2=2.91
r70 2 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.205
+ $Y=1.835 $X2=2.345 $Y2=1.98
r71 1 16 91 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=2 $X=1.665
+ $Y=0.235 $X2=1.845 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_1%VGND 1 2 9 13 16 17 19 20 21 33 34
r34 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r36 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r37 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r38 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 25 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r41 21 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r42 21 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r43 19 30 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.16
+ $Y2=0
r44 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.345
+ $Y2=0
r45 18 33 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.64
+ $Y2=0
r46 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.345
+ $Y2=0
r47 16 24 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.24 $Y2=0
r48 16 17 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.422
+ $Y2=0
r49 15 27 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.72
+ $Y2=0
r50 15 17 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.422
+ $Y2=0
r51 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=0.085
+ $X2=2.345 $Y2=0
r52 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=0.085
+ $X2=2.345 $Y2=0.38
r53 7 17 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.422 $Y=0.085
+ $X2=0.422 $Y2=0
r54 7 9 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=0.422 $Y=0.085
+ $X2=0.422 $Y2=0.38
r55 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.205
+ $Y=0.235 $X2=2.345 $Y2=0.38
r56 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.335
+ $Y=0.235 $X2=0.46 $Y2=0.38
.ends

