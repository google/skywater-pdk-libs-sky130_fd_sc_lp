* File: sky130_fd_sc_lp__xnor2_1.pex.spice
* Created: Fri Aug 28 11:34:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XNOR2_1%B 3 6 10 14 16 17 20 21 23 24 28 30
c81 21 0 2.5595e-19 $X=2.3 $Y=1.51
c82 20 0 1.7733e-19 $X=2.3 $Y=1.51
r83 28 31 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.35
+ $X2=0.385 $Y2=1.515
r84 28 30 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.35
+ $X2=0.385 $Y2=1.185
r85 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.355
+ $Y=1.35 $X2=0.355 $Y2=1.35
r86 24 29 10.2259 $w=3.53e-07 $l=3.15e-07 $layer=LI1_cond $X=0.262 $Y=1.665
+ $X2=0.262 $Y2=1.35
r87 23 29 1.78548 $w=3.53e-07 $l=5.5e-08 $layer=LI1_cond $X=0.262 $Y=1.295
+ $X2=0.262 $Y2=1.35
r88 21 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.51 $X2=2.3
+ $Y2=1.675
r89 21 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.51 $X2=2.3
+ $Y2=1.345
r90 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.3
+ $Y=1.51 $X2=2.3 $Y2=1.51
r91 18 24 8.27811 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.262 $Y=1.92
+ $X2=0.262 $Y2=1.665
r92 17 18 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.44 $Y=2.005
+ $X2=0.262 $Y2=1.92
r93 16 20 12.9592 $w=4.66e-07 $l=6.35157e-07 $layer=LI1_cond $X=1.825 $Y=2.005
+ $X2=2.145 $Y2=1.51
r94 16 17 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=1.825 $Y=2.005
+ $X2=0.44 $Y2=2.005
r95 14 34 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.39 $Y=2.465
+ $X2=2.39 $Y2=1.675
r96 10 33 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.39 $Y=0.655
+ $X2=2.39 $Y2=1.345
r97 6 31 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.505 $Y=2.465
+ $X2=0.505 $Y2=1.515
r98 3 30 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.505 $Y=0.655
+ $X2=0.505 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_1%A 1 3 6 8 10 13 16 17 18 19 20 25
c61 25 0 1.26526e-19 $X=1.49 $Y=1.51
r62 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.49
+ $Y=1.51 $X2=1.49 $Y2=1.51
r63 20 25 10.2833 $w=3.23e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=1.587
+ $X2=1.49 $Y2=1.587
r64 19 20 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.587
+ $X2=1.2 $Y2=1.587
r65 17 24 31.1191 $w=4.9e-07 $l=2.85e-07 $layer=POLY_cond $X=1.775 $Y=1.43
+ $X2=1.49 $Y2=1.43
r66 17 18 9.23259 $w=4.9e-07 $l=7.5e-08 $layer=POLY_cond $X=1.775 $Y=1.43
+ $X2=1.85 $Y2=1.43
r67 15 24 52.411 $w=4.9e-07 $l=4.8e-07 $layer=POLY_cond $X=1.01 $Y=1.43 $X2=1.49
+ $Y2=1.43
r68 15 16 9.23259 $w=4.9e-07 $l=1.1e-07 $layer=POLY_cond $X=1.01 $Y=1.43 $X2=0.9
+ $Y2=1.43
r69 11 18 47.473 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.85 $Y=1.675
+ $X2=1.85 $Y2=1.43
r70 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.85 $Y=1.675
+ $X2=1.85 $Y2=2.465
r71 8 18 47.473 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.85 $Y=1.185
+ $X2=1.85 $Y2=1.43
r72 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.85 $Y=1.185
+ $X2=1.85 $Y2=0.655
r73 4 16 47.473 $w=1.5e-07 $l=2.61916e-07 $layer=POLY_cond $X=0.935 $Y=1.675
+ $X2=0.9 $Y2=1.43
r74 4 6 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.935 $Y=1.675
+ $X2=0.935 $Y2=2.465
r75 1 16 47.473 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=0.9 $Y=1.185 $X2=0.9
+ $Y2=1.43
r76 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.9 $Y=1.185 $X2=0.9
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_1%A_33_47# 1 2 9 13 17 19 21 23 24 25 27 29 30
+ 34 41
c89 29 0 1.31259e-19 $X=2.76 $Y=1.675
c90 25 0 1.29424e-19 $X=2.165 $Y=2.345
c91 13 0 1.7733e-19 $X=2.885 $Y=2.465
r92 41 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.51
+ $X2=2.84 $Y2=1.675
r93 41 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.51
+ $X2=2.84 $Y2=1.345
r94 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.51 $X2=2.84 $Y2=1.51
r95 38 40 19.3832 $w=2.14e-07 $l=3.4e-07 $layer=LI1_cond $X=2.8 $Y=1.17 $X2=2.8
+ $Y2=1.51
r96 34 36 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.25 $Y=2.1 $X2=2.25
+ $Y2=2.345
r97 29 40 9.95691 $w=2.14e-07 $l=1.83916e-07 $layer=LI1_cond $X=2.76 $Y=1.675
+ $X2=2.8 $Y2=1.51
r98 29 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.76 $Y=1.675
+ $X2=2.76 $Y2=2.015
r99 28 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=2.1
+ $X2=2.25 $Y2=2.1
r100 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.675 $Y=2.1
+ $X2=2.76 $Y2=2.015
r101 27 28 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.675 $Y=2.1
+ $X2=2.335 $Y2=2.1
r102 26 33 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.815 $Y=2.345
+ $X2=0.685 $Y2=2.345
r103 25 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=2.345
+ $X2=2.25 $Y2=2.345
r104 25 26 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=2.165 $Y=2.345
+ $X2=0.815 $Y2=2.345
r105 23 38 2.08775 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.675 $Y=1.17
+ $X2=2.8 $Y2=1.17
r106 23 24 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=2.675 $Y=1.17
+ $X2=0.78 $Y2=1.17
r107 19 33 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=2.43
+ $X2=0.685 $Y2=2.345
r108 19 21 21.2759 $w=2.58e-07 $l=4.8e-07 $layer=LI1_cond $X=0.685 $Y=2.43
+ $X2=0.685 $Y2=2.91
r109 15 24 26.6617 $w=2.32e-07 $l=5.62183e-07 $layer=LI1_cond $X=0.29 $Y=1.015
+ $X2=0.78 $Y2=1.17
r110 15 17 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.29 $Y=0.845
+ $X2=0.29 $Y2=0.38
r111 13 44 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.885 $Y=2.465
+ $X2=2.885 $Y2=1.675
r112 9 43 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.885 $Y=0.655
+ $X2=2.885 $Y2=1.345
r113 2 33 600 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.345
r114 2 21 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.91
r115 1 17 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_1%VPWR 1 2 3 10 12 14 16 18 25 35 39 42 47
c46 3 0 1.46742e-19 $X=2.96 $Y=1.835
r47 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 37 39 11.2323 $w=8.13e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=3.007
+ $X2=1.825 $Y2=3.007
r49 34 37 0.660411 $w=8.13e-07 $l=4.5e-08 $layer=LI1_cond $X=1.635 $Y=3.007
+ $X2=1.68 $Y2=3.007
r50 34 35 18.6436 $w=8.13e-07 $l=6.5e-07 $layer=LI1_cond $X=1.635 $Y=3.007
+ $X2=0.985 $Y2=3.007
r51 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 29 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 28 39 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=1.825 $Y2=3.33
r54 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 25 41 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.935 $Y=3.33
+ $X2=3.147 $Y2=3.33
r56 25 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 24 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 23 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=0.985 $Y2=3.33
r60 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 21 31 4.08199 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.192 $Y2=3.33
r62 21 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 18 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 18 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 18 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 14 41 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.1 $Y=3.245
+ $X2=3.147 $Y2=3.33
r67 14 16 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.1 $Y=3.245
+ $X2=3.1 $Y2=2.85
r68 10 31 3.13023 $w=2.6e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.192 $Y2=3.33
r69 10 12 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.425
r70 3 16 600 $w=1.7e-07 $l=1.08274e-06 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.85
r71 2 34 300 $w=1.7e-07 $l=1.16118e-06 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=1.835 $X2=1.635 $Y2=2.725
r72 1 12 300 $w=1.7e-07 $l=6.495e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_1%Y 1 2 7 9 11 18 19 20 21 22 30 37 39 43
c33 43 0 1.46742e-19 $X=3.145 $Y=1.845
r34 36 39 2.65948 $w=2.58e-07 $l=6e-08 $layer=LI1_cond $X=3.145 $Y=1.975
+ $X2=3.145 $Y2=2.035
r35 22 37 3.02975 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=3.145 $Y=2.455
+ $X2=3.145 $Y2=2.355
r36 22 37 0.797845 $w=2.58e-07 $l=1.8e-08 $layer=LI1_cond $X=3.145 $Y=2.337
+ $X2=3.145 $Y2=2.355
r37 21 36 0.576222 $w=2.58e-07 $l=1.3e-08 $layer=LI1_cond $X=3.145 $Y=1.962
+ $X2=3.145 $Y2=1.975
r38 21 43 6.28782 $w=2.58e-07 $l=1.17e-07 $layer=LI1_cond $X=3.145 $Y=1.962
+ $X2=3.145 $Y2=1.845
r39 21 22 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.145 $Y=2.047
+ $X2=3.145 $Y2=2.337
r40 21 39 0.531897 $w=2.58e-07 $l=1.2e-08 $layer=LI1_cond $X=3.145 $Y=2.047
+ $X2=3.145 $Y2=2.035
r41 19 20 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.145 $Y=0.555
+ $X2=3.145 $Y2=0.925
r42 19 30 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=3.145 $Y=0.555
+ $X2=3.145 $Y2=0.42
r43 18 43 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.185 $Y=1.175
+ $X2=3.185 $Y2=1.845
r44 17 20 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=3.145 $Y=1.045
+ $X2=3.145 $Y2=0.925
r45 17 18 6.86404 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.145 $Y=1.045
+ $X2=3.145 $Y2=1.175
r46 12 16 3.93867 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=2.765 $Y=2.455
+ $X2=2.635 $Y2=2.455
r47 11 22 3.93867 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=3.015 $Y=2.455
+ $X2=3.145 $Y2=2.455
r48 11 12 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=3.015 $Y=2.455
+ $X2=2.765 $Y2=2.455
r49 7 16 3.02975 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=2.635 $Y=2.555 $X2=2.635
+ $Y2=2.455
r50 7 9 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=2.635 $Y=2.555
+ $X2=2.635 $Y2=2.91
r51 2 16 600 $w=1.7e-07 $l=7.30342e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.835 $X2=2.67 $Y2=2.47
r52 2 9 600 $w=1.7e-07 $l=1.17303e-06 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.835 $X2=2.67 $Y2=2.91
r53 1 30 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_1%VGND 1 2 9 13 16 17 18 24 30 31 34 39
r47 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r49 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r50 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=0 $X2=2.135
+ $Y2=0
r51 28 30 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.3 $Y=0 $X2=3.12
+ $Y2=0
r52 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=2.135
+ $Y2=0
r53 24 26 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.97 $Y=0 $X2=1.68
+ $Y2=0
r54 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r55 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r56 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r57 18 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r58 18 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r59 16 21 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.72
+ $Y2=0
r60 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.115
+ $Y2=0
r61 15 26 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.68
+ $Y2=0
r62 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.115
+ $Y2=0
r63 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=0.085
+ $X2=2.135 $Y2=0
r64 11 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.135 $Y=0.085
+ $X2=2.135 $Y2=0.455
r65 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0
r66 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.38
r67 2 13 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.135 $Y2=0.455
r68 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.975
+ $Y=0.235 $X2=1.115 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_1%A_302_47# 1 2 9 11 12 13 15
r29 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=0.745 $X2=2.67
+ $Y2=0.83
r30 13 15 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.67 $Y=0.745
+ $X2=2.67 $Y2=0.38
r31 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=0.83
+ $X2=2.67 $Y2=0.83
r32 11 12 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.505 $Y=0.83
+ $X2=1.8 $Y2=0.83
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.635 $Y=0.745
+ $X2=1.8 $Y2=0.83
r34 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.635 $Y=0.745
+ $X2=1.635 $Y2=0.38
r35 2 18 182 $w=1.7e-07 $l=6.89928e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.67 $Y2=0.83
r36 2 15 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=2.465
+ $Y=0.235 $X2=2.67 $Y2=0.38
r37 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.235 $X2=1.635 $Y2=0.38
.ends

