* File: sky130_fd_sc_lp__a31oi_lp.pex.spice
* Created: Fri Aug 28 10:00:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31OI_LP%A3 3 7 9 11 12 13 16 18 19 23 24
c36 24 0 9.33564e-21 $X=0.53 $Y=1.275
r37 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.53
+ $Y=1.275 $X2=0.53 $Y2=1.275
r38 18 19 7.76402 $w=5.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.41 $Y=1.295
+ $X2=0.41 $Y2=1.665
r39 18 24 0.419677 $w=5.68e-07 $l=2e-08 $layer=LI1_cond $X=0.41 $Y=1.295
+ $X2=0.41 $Y2=1.275
r40 14 16 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.62 $Y=0.805
+ $X2=0.8 $Y2=0.805
r41 12 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.53 $Y=1.615
+ $X2=0.53 $Y2=1.275
r42 12 13 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.615
+ $X2=0.53 $Y2=1.78
r43 11 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.11
+ $X2=0.53 $Y2=1.275
r44 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.8 $Y=0.73 $X2=0.8
+ $Y2=0.805
r45 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.8 $Y=0.73 $X2=0.8
+ $Y2=0.445
r46 5 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.62 $Y=0.88 $X2=0.62
+ $Y2=0.805
r47 5 11 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=0.62 $Y=0.88 $X2=0.62
+ $Y2=1.11
r48 3 13 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.57 $Y=2.545
+ $X2=0.57 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_LP%A2 1 3 7 11 12 13 14 15 21
c49 7 0 1.77034e-19 $X=1.19 $Y=0.445
r50 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.1
+ $Y=1.285 $X2=1.1 $Y2=1.285
r51 14 15 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.125 $Y=1.295
+ $X2=1.125 $Y2=1.665
r52 14 22 0.303274 $w=3.78e-07 $l=1e-08 $layer=LI1_cond $X=1.125 $Y=1.295
+ $X2=1.125 $Y2=1.285
r53 13 22 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.125 $Y=0.925
+ $X2=1.125 $Y2=1.285
r54 12 13 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.125 $Y=0.555
+ $X2=1.125 $Y2=0.925
r55 11 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.1 $Y=1.625 $X2=1.1
+ $Y2=1.285
r56 10 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.12 $X2=1.1
+ $Y2=1.285
r57 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.19 $Y=0.445
+ $X2=1.19 $Y2=1.12
r58 1 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.79 $X2=1.1
+ $Y2=1.625
r59 1 3 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.1 $Y=1.79 $X2=1.1
+ $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_LP%A1 3 5 7 11 12 13 17
r40 12 13 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.67 $Y=1.285
+ $X2=1.67 $Y2=1.665
r41 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.67
+ $Y=1.285 $X2=1.67 $Y2=1.285
r42 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.67 $Y=1.625
+ $X2=1.67 $Y2=1.285
r43 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.12
+ $X2=1.67 $Y2=1.285
r44 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.79
+ $X2=1.67 $Y2=1.625
r45 5 7 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.67 $Y=1.79 $X2=1.67
+ $Y2=2.545
r46 3 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.58 $Y=0.445
+ $X2=1.58 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_LP%B1 1 3 8 10 12 16 19 20 21 22 23 27
r49 22 23 12.1647 $w=3.58e-07 $l=3.8e-07 $layer=LI1_cond $X=2.225 $Y=1.285
+ $X2=2.225 $Y2=1.665
r50 22 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.24
+ $Y=1.285 $X2=2.24 $Y2=1.285
r51 20 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.24 $Y=1.625
+ $X2=2.24 $Y2=1.285
r52 20 21 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.24 $Y=1.625
+ $X2=2.24 $Y2=1.79
r53 19 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.24 $Y=1.12
+ $X2=2.24 $Y2=1.285
r54 15 16 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.15 $Y=0.805
+ $X2=2.37 $Y2=0.805
r55 13 15 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.01 $Y=0.805
+ $X2=2.15 $Y2=0.805
r56 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=0.73
+ $X2=2.37 $Y2=0.805
r57 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.37 $Y=0.73 $X2=2.37
+ $Y2=0.445
r58 8 21 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.2 $Y=2.545 $X2=2.2
+ $Y2=1.79
r59 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.15 $Y=0.88 $X2=2.15
+ $Y2=0.805
r60 4 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.15 $Y=0.88 $X2=2.15
+ $Y2=1.12
r61 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.01 $Y=0.73 $X2=2.01
+ $Y2=0.805
r62 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.01 $Y=0.73 $X2=2.01
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_LP%VPWR 1 2 7 9 13 17 19 26 27 33
r35 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r37 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 24 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 23 26 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r41 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 21 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.53 $Y=3.33
+ $X2=1.365 $Y2=3.33
r43 21 23 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.53 $Y=3.33 $X2=1.68
+ $Y2=3.33
r44 19 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 19 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 15 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=3.245
+ $X2=1.365 $Y2=3.33
r47 15 17 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.365 $Y=3.245
+ $X2=1.365 $Y2=2.485
r48 14 30 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=3.33
+ $X2=0.235 $Y2=3.33
r49 13 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=1.365 $Y2=3.33
r50 13 14 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=0.47
+ $Y2=3.33
r51 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.305 $Y=2.19
+ $X2=0.305 $Y2=2.9
r52 7 30 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.235 $Y2=3.33
r53 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.305 $Y2=2.9
r54 2 17 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=1.225
+ $Y=2.045 $X2=1.365 $Y2=2.485
r55 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.045 $X2=0.305 $Y2=2.9
r56 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.045 $X2=0.305 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_LP%A_139_409# 1 2 9 13 14 17
r36 17 19 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.935 $Y=2.19
+ $X2=1.935 $Y2=2.9
r37 15 17 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.935 $Y=2.14
+ $X2=1.935 $Y2=2.19
r38 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.77 $Y=2.055
+ $X2=1.935 $Y2=2.14
r39 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.77 $Y=2.055 $X2=1
+ $Y2=2.055
r40 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.835 $Y=2.19
+ $X2=0.835 $Y2=2.9
r41 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.835 $Y=2.14
+ $X2=1 $Y2=2.055
r42 7 9 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.835 $Y=2.14 $X2=0.835
+ $Y2=2.19
r43 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=2.045 $X2=1.935 $Y2=2.9
r44 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=2.045 $X2=1.935 $Y2=2.19
r45 1 11 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.695
+ $Y=2.045 $X2=0.835 $Y2=2.9
r46 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.695
+ $Y=2.045 $X2=0.835 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_LP%Y 1 2 9 11 12 17 18 19 20
c41 12 0 1.67698e-19 $X=1.96 $Y=0.855
r42 20 28 3.28593 $w=4.53e-07 $l=1.25e-07 $layer=LI1_cond $X=2.527 $Y=2.775
+ $X2=2.527 $Y2=2.9
r43 19 20 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.527 $Y=2.405
+ $X2=2.527 $Y2=2.775
r44 17 18 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=2.527 $Y=2.19
+ $X2=2.527 $Y2=2.025
r45 15 19 4.02198 $w=4.53e-07 $l=1.53e-07 $layer=LI1_cond $X=2.527 $Y=2.252
+ $X2=2.527 $Y2=2.405
r46 15 17 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=2.527 $Y=2.252
+ $X2=2.527 $Y2=2.19
r47 13 18 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=2.67 $Y=0.94
+ $X2=2.67 $Y2=2.025
r48 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.585 $Y=0.855
+ $X2=2.67 $Y2=0.94
r49 11 12 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.585 $Y=0.855
+ $X2=1.96 $Y2=0.855
r50 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.795 $Y=0.77
+ $X2=1.96 $Y2=0.855
r51 7 9 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.795 $Y=0.77 $X2=1.795
+ $Y2=0.47
r52 2 28 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=2.045 $X2=2.465 $Y2=2.9
r53 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=2.045 $X2=2.465 $Y2=2.19
r54 1 9 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.235 $X2=1.795 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A31OI_LP%VGND 1 2 9 11 13 15 17 22 28 32
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r41 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=0 $X2=0.585
+ $Y2=0
r43 23 25 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=0.75 $Y=0 $X2=2.16
+ $Y2=0
r44 22 31 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.65
+ $Y2=0
r45 22 25 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.16
+ $Y2=0
r46 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.42 $Y=0 $X2=0.585
+ $Y2=0
r49 17 19 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.42 $Y=0 $X2=0.24
+ $Y2=0
r50 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r51 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r52 11 31 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.585 $Y=0.085
+ $X2=2.65 $Y2=0
r53 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.585 $Y=0.085
+ $X2=2.585 $Y2=0.4
r54 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.585 $Y=0.085
+ $X2=0.585 $Y2=0
r55 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.585 $Y=0.085
+ $X2=0.585 $Y2=0.445
r56 2 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.445
+ $Y=0.235 $X2=2.585 $Y2=0.4
r57 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.44
+ $Y=0.235 $X2=0.585 $Y2=0.445
.ends

