* File: sky130_fd_sc_lp__sdfbbp_1.pex.spice
* Created: Wed Sep  2 10:33:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%SCD 5 9 13 15 16 17 18 21 22
c41 21 0 3.63052e-20 $X=0.385 $Y=1.38
r42 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.38 $X2=0.385 $Y2=1.38
r43 18 22 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.55
+ $X2=0.385 $Y2=1.55
r44 16 17 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=0.485 $Y=2.12
+ $X2=0.485 $Y2=2.27
r45 15 16 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=0.475 $Y=1.885
+ $X2=0.475 $Y2=2.12
r46 14 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.72
+ $X2=0.385 $Y2=1.38
r47 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.72
+ $X2=0.385 $Y2=1.885
r48 13 21 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.385 $Y=1.31
+ $X2=0.385 $Y2=1.38
r49 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.425 $Y=1.16
+ $X2=0.425 $Y2=1.31
r50 9 12 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=0.555 $Y=0.805
+ $X2=0.555 $Y2=1.16
r51 5 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.495 $Y=2.725
+ $X2=0.495 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%D 3 7 9 15
c43 9 0 3.02992e-19 $X=1.68 $Y=1.665
r44 13 15 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.435 $Y=1.69
+ $X2=1.625 $Y2=1.69
r45 11 13 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.375 $Y=1.69
+ $X2=1.435 $Y2=1.69
r46 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.69 $X2=1.625 $Y2=1.69
r47 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.855
+ $X2=1.435 $Y2=1.69
r48 5 7 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.435 $Y=1.855
+ $X2=1.435 $Y2=2.725
r49 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.525
+ $X2=1.375 $Y2=1.69
r50 1 3 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.375 $Y=1.525
+ $X2=1.375 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_332_93# 1 2 7 9 12 14 15 17 19 22 25 28
+ 30 36 39 40 44
c91 39 0 1.52779e-19 $X=2.49 $Y=1.69
c92 22 0 3.10692e-20 $X=2.075 $Y=2.17
c93 15 0 1.65e-19 $X=1.81 $Y=1.165
c94 14 0 1.50206e-19 $X=2 $Y=1.165
r95 39 42 2.24867 $w=4.08e-07 $l=8e-08 $layer=LI1_cond $X=2.53 $Y=1.69 $X2=2.53
+ $Y2=1.77
r96 39 41 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=1.69
+ $X2=2.53 $Y2=1.525
r97 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.69 $X2=2.49 $Y2=1.69
r98 36 44 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=2.55
+ $X2=3.15 $Y2=2.385
r99 32 44 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.07 $Y=1.855
+ $X2=3.07 $Y2=2.385
r100 31 42 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.735 $Y=1.77
+ $X2=2.53 $Y2=1.77
r101 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.985 $Y=1.77
+ $X2=3.07 $Y2=1.855
r102 30 31 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.985 $Y=1.77
+ $X2=2.735 $Y2=1.77
r103 28 41 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.65 $Y=0.825
+ $X2=2.65 $Y2=1.525
r104 24 40 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.15 $Y=1.69
+ $X2=2.49 $Y2=1.69
r105 24 25 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.15 $Y=1.69
+ $X2=2.075 $Y2=1.69
r106 20 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.865 $Y=2.17
+ $X2=2.075 $Y2=2.17
r107 19 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.075 $Y=2.095
+ $X2=2.075 $Y2=2.17
r108 18 25 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.855
+ $X2=2.075 $Y2=1.69
r109 18 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.075 $Y=1.855
+ $X2=2.075 $Y2=2.095
r110 17 25 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.525
+ $X2=2.075 $Y2=1.69
r111 16 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.075 $Y=1.24
+ $X2=2.075 $Y2=1.525
r112 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2 $Y=1.165
+ $X2=2.075 $Y2=1.24
r113 14 15 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2 $Y=1.165 $X2=1.81
+ $Y2=1.165
r114 10 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.865 $Y=2.245
+ $X2=1.865 $Y2=2.17
r115 10 12 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.865 $Y=2.245
+ $X2=1.865 $Y2=2.725
r116 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.735 $Y=1.09
+ $X2=1.81 $Y2=1.165
r117 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.735 $Y=1.09
+ $X2=1.735 $Y2=0.805
r118 2 36 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.01
+ $Y=2.405 $X2=3.15 $Y2=2.55
r119 1 28 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=2.51
+ $Y=0.595 $X2=2.65 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%SCE 4 9 11 12 16 17 18 21 25 26 27 28 29 32
c97 27 0 1.52779e-19 $X=2.952 $Y=2.095
c98 26 0 3.13616e-19 $X=1.03 $Y=2.245
c99 25 0 1.64649e-19 $X=1.03 $Y=2.095
c100 4 0 1.06923e-19 $X=0.945 $Y=0.805
r101 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.715
+ $X2=0.925 $Y2=1.88
r102 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.715
+ $X2=0.925 $Y2=1.55
r103 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.715 $X2=0.925 $Y2=1.715
r104 29 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.2 $Y=1.715
+ $X2=0.925 $Y2=1.715
r105 27 28 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=2.952 $Y=2.095
+ $X2=2.952 $Y2=2.245
r106 25 26 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.03 $Y=2.095
+ $X2=1.03 $Y2=2.245
r107 25 35 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.015 $Y=2.095
+ $X2=1.015 $Y2=1.88
r108 23 27 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.97 $Y=1.24
+ $X2=2.97 $Y2=2.095
r109 21 28 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.935 $Y=2.725
+ $X2=2.935 $Y2=2.245
r110 17 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.895 $Y=1.165
+ $X2=2.97 $Y2=1.24
r111 17 18 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.895 $Y=1.165
+ $X2=2.51 $Y2=1.165
r112 14 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.435 $Y=1.09
+ $X2=2.51 $Y2=1.165
r113 14 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.435 $Y=1.09
+ $X2=2.435 $Y2=0.805
r114 13 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.435 $Y=0.255
+ $X2=2.435 $Y2=0.805
r115 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.36 $Y=0.18
+ $X2=2.435 $Y2=0.255
r116 11 12 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=2.36 $Y=0.18
+ $X2=1.02 $Y2=0.18
r117 9 26 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.045 $Y=2.725
+ $X2=1.045 $Y2=2.245
r118 4 34 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=0.945 $Y=0.805
+ $X2=0.945 $Y2=1.55
r119 1 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.945 $Y=0.255
+ $X2=1.02 $Y2=0.18
r120 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.945 $Y=0.255
+ $X2=0.945 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%CLK 3 7 12 14 16 17 21
r42 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.61 $Y=1.665
+ $X2=3.61 $Y2=2.035
r43 16 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.61
+ $Y=1.665 $X2=3.61 $Y2=1.665
r44 12 21 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=3.61 $Y=2.02
+ $X2=3.61 $Y2=1.665
r45 12 14 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=3.61 $Y=2.095
+ $X2=3.925 $Y2=2.095
r46 10 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.61 $Y=1.5
+ $X2=3.61 $Y2=1.665
r47 5 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.925 $Y=2.17
+ $X2=3.925 $Y2=2.095
r48 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.925 $Y=2.17
+ $X2=3.925 $Y2=2.69
r49 3 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.7 $Y=0.74 $X2=3.7
+ $Y2=1.5
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_893_101# 1 2 7 8 10 13 15 16 19 21 23 26
+ 29 33 37 39 41 44 48 49 55 59 60 63 64
c175 44 0 1.49262e-19 $X=9.915 $Y=2.25
c176 21 0 1.36771e-19 $X=9.74 $Y=2.455
c177 19 0 6.11734e-20 $X=6.515 $Y=0.445
c178 15 0 7.21799e-20 $X=6.37 $Y=1.165
r179 63 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.775 $Y=1.29
+ $X2=9.775 $Y2=1.125
r180 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.775
+ $Y=1.29 $X2=9.775 $Y2=1.29
r181 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.395
+ $Y=1.58 $X2=5.395 $Y2=1.58
r182 55 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.295
+ $X2=9.84 $Y2=1.295
r183 52 60 7.64176 $w=4.55e-07 $l=3.72552e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.242 $Y2=1.58
r184 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.295
r185 49 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.295
+ $X2=5.04 $Y2=1.295
r186 48 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.295
+ $X2=9.84 $Y2=1.295
r187 48 49 5.58167 $w=1.4e-07 $l=4.51e-06 $layer=MET1_cond $X=9.695 $Y=1.295
+ $X2=5.185 $Y2=1.295
r188 46 64 26.5563 $w=3.43e-07 $l=7.95e-07 $layer=LI1_cond $X=9.782 $Y=2.085
+ $X2=9.782 $Y2=1.29
r189 44 46 4.89723 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=9.827 $Y=2.25
+ $X2=9.827 $Y2=2.085
r190 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.915
+ $Y=2.25 $X2=9.915 $Y2=2.25
r191 40 41 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.865 $Y=2 $X2=4.695
+ $Y2=2
r192 39 60 11.2615 $w=4.55e-07 $l=4.2e-07 $layer=LI1_cond $X=5.242 $Y=2
+ $X2=5.242 $Y2=1.58
r193 39 40 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.045 $Y=2
+ $X2=4.865 $Y2=2
r194 35 41 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=2.085
+ $X2=4.695 $Y2=2
r195 35 37 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=4.695 $Y=2.085
+ $X2=4.695 $Y2=2.43
r196 31 41 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.61 $Y=1.915
+ $X2=4.695 $Y2=2
r197 31 33 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=4.61 $Y=1.915
+ $X2=4.61 $Y2=0.78
r198 28 59 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.395 $Y=1.565
+ $X2=5.395 $Y2=1.58
r199 26 65 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=9.745 $Y=0.605
+ $X2=9.745 $Y2=1.125
r200 21 45 26.034 $w=3.24e-07 $l=2.5807e-07 $layer=POLY_cond $X=9.74 $Y=2.455
+ $X2=9.915 $Y2=2.27
r201 21 23 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=9.74 $Y=2.455
+ $X2=9.74 $Y2=2.785
r202 17 30 5.80308 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.515 $Y=1.06
+ $X2=6.515 $Y2=1.15
r203 17 19 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=6.515 $Y=1.06
+ $X2=6.515 $Y2=0.445
r204 15 30 41.8991 $w=1.7e-07 $l=1.52315e-07 $layer=POLY_cond $X=6.37 $Y=1.165
+ $X2=6.515 $Y2=1.15
r205 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=6.37 $Y=1.165
+ $X2=6.08 $Y2=1.165
r206 11 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.005 $Y=1.565
+ $X2=6.005 $Y2=1.49
r207 11 13 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=6.005 $Y=1.565
+ $X2=6.005 $Y2=2.495
r208 10 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.005 $Y=1.415
+ $X2=6.005 $Y2=1.49
r209 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.005 $Y=1.24
+ $X2=6.08 $Y2=1.165
r210 9 10 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.005 $Y=1.24
+ $X2=6.005 $Y2=1.415
r211 8 28 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.56 $Y=1.49
+ $X2=5.395 $Y2=1.565
r212 7 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.93 $Y=1.49
+ $X2=6.005 $Y2=1.49
r213 7 8 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.93 $Y=1.49 $X2=5.56
+ $Y2=1.49
r214 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=4.555
+ $Y=2.285 $X2=4.7 $Y2=2.43
r215 1 33 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=4.465
+ $Y=0.505 $X2=4.61 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_1297_290# 1 2 9 13 17 19 20 23 26 27 28
+ 29 30 31 34 35 39 40 45 53 55 57
c179 45 0 6.02433e-20 $X=6.65 $Y=1.615
c180 35 0 1.36771e-19 $X=9.03 $Y=2.045
c181 30 0 1.11578e-19 $X=7.63 $Y=2.33
c182 29 0 1.98194e-19 $X=7.63 $Y=2.13
c183 26 0 5.71347e-21 $X=6.57 $Y=2.33
c184 23 0 1.77109e-19 $X=9.325 $Y=0.605
r185 57 58 7.77419 $w=3.1e-07 $l=5e-08 $layer=POLY_cond $X=6.825 $Y=1.615
+ $X2=6.875 $Y2=1.615
r186 51 53 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.11 $Y=0.73
+ $X2=8.26 $Y2=0.73
r187 46 57 27.2097 $w=3.1e-07 $l=1.75e-07 $layer=POLY_cond $X=6.65 $Y=1.615
+ $X2=6.825 $Y2=1.615
r188 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.65
+ $Y=1.615 $X2=6.65 $Y2=1.615
r189 42 45 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=6.57 $Y=1.61 $X2=6.65
+ $Y2=1.61
r190 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.195
+ $Y=1.29 $X2=9.195 $Y2=1.29
r191 37 39 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=9.195 $Y=1.96
+ $X2=9.195 $Y2=1.29
r192 36 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.345 $Y=2.045
+ $X2=8.26 $Y2=2.045
r193 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.03 $Y=2.045
+ $X2=9.195 $Y2=1.96
r194 35 36 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=9.03 $Y=2.045
+ $X2=8.345 $Y2=2.045
r195 34 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.26 $Y=1.96
+ $X2=8.26 $Y2=2.045
r196 33 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.26 $Y=0.815
+ $X2=8.26 $Y2=0.73
r197 33 34 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=8.26 $Y=0.815
+ $X2=8.26 $Y2=1.96
r198 32 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=2.045
+ $X2=7.63 $Y2=2.045
r199 31 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.175 $Y=2.045
+ $X2=8.26 $Y2=2.045
r200 31 32 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.175 $Y=2.045
+ $X2=7.795 $Y2=2.045
r201 29 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.63 $Y=2.13 $X2=7.63
+ $Y2=2.045
r202 29 30 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=7.63 $Y=2.13 $X2=7.63
+ $Y2=2.33
r203 27 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.465 $Y=2.415
+ $X2=7.63 $Y2=2.33
r204 27 28 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=7.465 $Y=2.415
+ $X2=6.655 $Y2=2.415
r205 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.57 $Y=2.33
+ $X2=6.655 $Y2=2.415
r206 25 42 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.57 $Y=1.77
+ $X2=6.57 $Y2=1.61
r207 25 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.57 $Y=1.77
+ $X2=6.57 $Y2=2.33
r208 21 40 38.7026 $w=2.82e-07 $l=2.13014e-07 $layer=POLY_cond $X=9.325 $Y=1.125
+ $X2=9.215 $Y2=1.29
r209 21 23 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=9.325 $Y=1.125
+ $X2=9.325 $Y2=0.605
r210 19 40 52.9858 $w=2.82e-07 $l=3.91727e-07 $layer=POLY_cond $X=9.03 $Y=1.6
+ $X2=9.215 $Y2=1.29
r211 19 20 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=9.03 $Y=1.6 $X2=8.83
+ $Y2=1.6
r212 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.755 $Y=1.675
+ $X2=8.83 $Y2=1.6
r213 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.755 $Y=1.675
+ $X2=8.755 $Y2=2.285
r214 11 58 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.875 $Y=1.45
+ $X2=6.875 $Y2=1.615
r215 11 13 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=6.875 $Y=1.45
+ $X2=6.875 $Y2=0.445
r216 7 57 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=1.78
+ $X2=6.825 $Y2=1.615
r217 7 9 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=6.825 $Y=1.78
+ $X2=6.825 $Y2=2.495
r218 2 49 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=7.49
+ $Y=1.865 $X2=7.63 $Y2=2.125
r219 1 51 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=7.89
+ $Y=0.235 $X2=8.11 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%SET_B 3 7 11 13 15 18 19 21 22 28 32 38 44
c136 38 0 1.48965e-19 $X=11.245 $Y=1.93
c137 28 0 5.60316e-21 $X=11.28 $Y=2.035
c138 22 0 3.09772e-19 $X=7.105 $Y=2.035
c139 11 0 1.26004e-19 $X=11.32 $Y=0.605
c140 7 0 5.15316e-20 $X=7.415 $Y=2.285
r141 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.245
+ $Y=1.93 $X2=11.245 $Y2=1.93
r142 33 46 6.97157 $w=4.03e-07 $l=2.45e-07 $layer=LI1_cond $X=7.325 $Y=1.577
+ $X2=7.08 $Y2=1.577
r143 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.325 $Y=1.54
+ $X2=7.325 $Y2=1.705
r144 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.325 $Y=1.54
+ $X2=7.325 $Y2=1.375
r145 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.325
+ $Y=1.54 $X2=7.325 $Y2=1.54
r146 28 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=2.035
+ $X2=11.28 $Y2=2.035
r147 25 44 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=6.96 $Y=2.05
+ $X2=7.08 $Y2=2.05
r148 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=2.035
+ $X2=6.96 $Y2=2.035
r149 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=2.035
+ $X2=6.96 $Y2=2.035
r150 21 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=11.28 $Y2=2.035
r151 21 22 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=7.105 $Y2=2.035
r152 19 33 3.27237 $w=4.03e-07 $l=1.15e-07 $layer=LI1_cond $X=7.44 $Y=1.577
+ $X2=7.325 $Y2=1.577
r153 18 44 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.08 $Y=1.95 $X2=7.08
+ $Y2=2.05
r154 17 46 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=7.08 $Y=1.78
+ $X2=7.08 $Y2=1.577
r155 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.08 $Y=1.78
+ $X2=7.08 $Y2=1.95
r156 13 37 38.8445 $w=3.55e-07 $l=2.1609e-07 $layer=POLY_cond $X=11.39 $Y=2.095
+ $X2=11.272 $Y2=1.93
r157 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.39 $Y=2.095
+ $X2=11.39 $Y2=2.675
r158 9 37 38.8445 $w=3.55e-07 $l=1.8747e-07 $layer=POLY_cond $X=11.32 $Y=1.765
+ $X2=11.272 $Y2=1.93
r159 9 11 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=11.32 $Y=1.765
+ $X2=11.32 $Y2=0.605
r160 7 35 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.415 $Y=2.285
+ $X2=7.415 $Y2=1.705
r161 3 34 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.385 $Y=0.555
+ $X2=7.385 $Y2=1.375
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_1216_457# 1 2 9 13 17 18 21 25 27 31 33
+ 34
c95 34 0 1.67734e-19 $X=7.865 $Y=1.19
c96 33 0 1.71701e-19 $X=7.865 $Y=1.19
r97 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.865
+ $Y=1.19 $X2=7.865 $Y2=1.19
r98 28 31 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.465 $Y=1.11
+ $X2=6.3 $Y2=1.11
r99 27 33 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.705 $Y=1.11
+ $X2=7.85 $Y2=1.11
r100 27 28 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.705 $Y=1.11
+ $X2=6.465 $Y2=1.11
r101 23 31 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.22 $Y=1.195
+ $X2=6.3 $Y2=1.11
r102 23 25 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=6.22 $Y=1.195
+ $X2=6.22 $Y2=2.495
r103 19 31 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.3 $Y=1.025 $X2=6.3
+ $Y2=1.11
r104 19 21 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=6.3 $Y=1.025
+ $X2=6.3 $Y2=0.47
r105 17 34 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.865 $Y=1.53
+ $X2=7.865 $Y2=1.19
r106 17 18 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.865 $Y=1.53
+ $X2=7.865 $Y2=1.695
r107 16 34 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.865 $Y=1.025
+ $X2=7.865 $Y2=1.19
r108 13 18 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=7.845 $Y=2.285
+ $X2=7.845 $Y2=1.695
r109 9 16 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=7.815 $Y=0.555 $X2=7.815
+ $Y2=1.025
r110 2 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.08
+ $Y=2.285 $X2=6.22 $Y2=2.495
r111 1 21 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=6.16
+ $Y=0.235 $X2=6.3 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_1650_21# 1 2 7 9 12 16 18 20 24 31 32 34
+ 35 37 38 39 41 42 43 44 47 49 51 53 57 62
c173 44 0 1.8236e-19 $X=12.5 $Y=0.915
c174 32 0 1.71701e-19 $X=8.655 $Y=1.15
c175 24 0 1.75295e-19 $X=12.635 $Y=1.785
r176 62 64 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=13.145 $Y=0.815
+ $X2=13.145 $Y2=0.915
r177 53 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.675 $Y=0.915
+ $X2=11.675 $Y2=1.085
r178 52 57 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.8 $Y=0.915
+ $X2=12.65 $Y2=0.915
r179 51 64 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.02 $Y=0.915
+ $X2=13.145 $Y2=0.915
r180 51 52 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=13.02 $Y=0.915
+ $X2=12.8 $Y2=0.915
r181 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.635
+ $Y=1.43 $X2=12.635 $Y2=1.43
r182 47 60 21.187 $w=2.62e-07 $l=4.55e-07 $layer=LI1_cond $X=12.65 $Y=1.935
+ $X2=13.105 $Y2=1.935
r183 47 49 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=12.65 $Y=1.765
+ $X2=12.65 $Y2=1.43
r184 46 57 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.65 $Y=1 $X2=12.65
+ $Y2=0.915
r185 46 49 16.5184 $w=2.98e-07 $l=4.3e-07 $layer=LI1_cond $X=12.65 $Y=1
+ $X2=12.65 $Y2=1.43
r186 45 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.76 $Y=0.915
+ $X2=11.675 $Y2=0.915
r187 44 57 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.5 $Y=0.915
+ $X2=12.65 $Y2=0.915
r188 44 45 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=12.5 $Y=0.915
+ $X2=11.76 $Y2=0.915
r189 42 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.59 $Y=1.085
+ $X2=11.675 $Y2=1.085
r190 42 43 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=11.59 $Y=1.085
+ $X2=10.655 $Y2=1.085
r191 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.57 $Y=1
+ $X2=10.655 $Y2=1.085
r192 40 41 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=10.57 $Y=0.435
+ $X2=10.57 $Y2=1
r193 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.485 $Y=0.35
+ $X2=10.57 $Y2=0.435
r194 38 39 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=10.485 $Y=0.35
+ $X2=9.615 $Y2=0.35
r195 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.53 $Y=0.435
+ $X2=9.615 $Y2=0.35
r196 36 37 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.53 $Y=0.435
+ $X2=9.53 $Y2=0.775
r197 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.445 $Y=0.86
+ $X2=9.53 $Y2=0.775
r198 34 35 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=9.445 $Y=0.86
+ $X2=8.82 $Y2=0.86
r199 32 67 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=8.655 $Y=1.15
+ $X2=8.325 $Y2=1.15
r200 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.655
+ $Y=1.15 $X2=8.655 $Y2=1.15
r201 29 35 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=8.672 $Y=0.945
+ $X2=8.82 $Y2=0.86
r202 29 31 8.0085 $w=2.93e-07 $l=2.05e-07 $layer=LI1_cond $X=8.672 $Y=0.945
+ $X2=8.672 $Y2=1.15
r203 24 50 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=12.635 $Y=1.785
+ $X2=12.635 $Y2=1.43
r204 21 24 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=12.32 $Y=1.86
+ $X2=12.635 $Y2=1.86
r205 18 50 58.4553 $w=2.35e-07 $l=5.54482e-07 $layer=POLY_cond $X=12.35 $Y=1
+ $X2=12.635 $Y2=1.43
r206 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=12.35 $Y=1
+ $X2=12.35 $Y2=0.605
r207 14 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.32 $Y=1.935
+ $X2=12.32 $Y2=1.86
r208 14 16 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.32 $Y=1.935
+ $X2=12.32 $Y2=2.675
r209 10 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.325 $Y=1.315
+ $X2=8.325 $Y2=1.15
r210 10 12 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=8.325 $Y=1.315
+ $X2=8.325 $Y2=2.285
r211 7 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.325 $Y=0.985
+ $X2=8.325 $Y2=1.15
r212 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.325 $Y=0.985
+ $X2=8.325 $Y2=0.555
r213 2 60 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=12.96
+ $Y=1.785 $X2=13.105 $Y2=1.995
r214 1 62 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=12.96
+ $Y=0.655 $X2=13.105 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_755_106# 1 2 7 8 9 11 15 16 18 19 21 22
+ 23 24 26 29 31 36 37 38 41 44 45 49 53 56 58
c159 37 0 1.03084e-19 $X=10.18 $Y=1.77
c160 29 0 1.44251e-20 $X=6.435 $Y=2.495
r161 56 58 31.1954 $w=2.88e-07 $l=7.85e-07 $layer=LI1_cond $X=4.2 $Y=2.515
+ $X2=4.2 $Y2=1.73
r162 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.18
+ $Y=1.225 $X2=4.18 $Y2=1.225
r163 49 52 13.1924 $w=3.78e-07 $l=4.35e-07 $layer=LI1_cond $X=4.155 $Y=0.79
+ $X2=4.155 $Y2=1.225
r164 47 58 6.43709 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=4.155 $Y=1.54
+ $X2=4.155 $Y2=1.73
r165 47 52 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=4.155 $Y=1.54
+ $X2=4.155 $Y2=1.225
r166 43 53 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=4.18 $Y=1.175
+ $X2=4.18 $Y2=1.225
r167 39 41 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=10.255 $Y=1.695
+ $X2=10.255 $Y2=0.715
r168 38 46 69.8667 $w=2.35e-07 $l=3.75566e-07 $layer=POLY_cond $X=9.54 $Y=1.77
+ $X2=9.23 $Y2=1.915
r169 37 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.18 $Y=1.77
+ $X2=10.255 $Y2=1.695
r170 37 38 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=10.18 $Y=1.77
+ $X2=9.54 $Y2=1.77
r171 34 36 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=9.23 $Y=3.075
+ $X2=9.23 $Y2=2.575
r172 33 46 13.2911 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=9.23 $Y=2.065
+ $X2=9.23 $Y2=1.915
r173 33 36 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=9.23 $Y=2.065
+ $X2=9.23 $Y2=2.575
r174 32 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.51 $Y=3.15
+ $X2=6.435 $Y2=3.15
r175 31 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.155 $Y=3.15
+ $X2=9.23 $Y2=3.075
r176 31 32 1356.27 $w=1.5e-07 $l=2.645e-06 $layer=POLY_cond $X=9.155 $Y=3.15
+ $X2=6.51 $Y2=3.15
r177 27 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.435 $Y=3.075
+ $X2=6.435 $Y2=3.15
r178 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.435 $Y=3.075
+ $X2=6.435 $Y2=2.495
r179 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.085 $Y=0.73
+ $X2=6.085 $Y2=0.445
r180 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.01 $Y=0.805
+ $X2=6.085 $Y2=0.73
r181 22 23 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=6.01 $Y=0.805
+ $X2=5.68 $Y2=0.805
r182 20 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.605 $Y=0.88
+ $X2=5.68 $Y2=0.805
r183 20 21 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.605 $Y=0.88
+ $X2=5.605 $Y2=1.025
r184 18 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.36 $Y=3.15
+ $X2=6.435 $Y2=3.15
r185 18 19 702.489 $w=1.5e-07 $l=1.37e-06 $layer=POLY_cond $X=6.36 $Y=3.15
+ $X2=4.99 $Y2=3.15
r186 17 44 12.05 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=4.99 $Y=1.1 $X2=4.87
+ $Y2=1.1
r187 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.53 $Y=1.1
+ $X2=5.605 $Y2=1.025
r188 16 17 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.53 $Y=1.1
+ $X2=4.99 $Y2=1.1
r189 13 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.915 $Y=3.075
+ $X2=4.99 $Y2=3.15
r190 13 15 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.915 $Y=3.075
+ $X2=4.915 $Y2=2.605
r191 12 44 12.05 $w=1.5e-07 $l=9.48683e-08 $layer=POLY_cond $X=4.915 $Y=1.175
+ $X2=4.87 $Y2=1.1
r192 12 15 733.255 $w=1.5e-07 $l=1.43e-06 $layer=POLY_cond $X=4.915 $Y=1.175
+ $X2=4.915 $Y2=2.605
r193 9 44 12.05 $w=1.5e-07 $l=9.48683e-08 $layer=POLY_cond $X=4.825 $Y=1.025
+ $X2=4.87 $Y2=1.1
r194 9 11 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=4.825 $Y=1.025
+ $X2=4.825 $Y2=0.715
r195 8 43 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.345 $Y=1.1
+ $X2=4.18 $Y2=1.175
r196 7 44 12.05 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=4.75 $Y=1.1 $X2=4.87
+ $Y2=1.1
r197 7 8 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.75 $Y=1.1 $X2=4.345
+ $Y2=1.1
r198 2 56 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4
+ $Y=2.37 $X2=4.14 $Y2=2.515
r199 1 49 182 $w=1.7e-07 $l=3.83569e-07 $layer=licon1_NDIFF $count=1 $X=3.775
+ $Y=0.53 $X2=4.05 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_2064_453# 1 2 9 13 17 21 23 27 31 36 40
+ 43 44 46 47 50 53 54 57 59 63 65 69 73
c172 63 0 1.75295e-19 $X=12.235 $Y=1.37
c173 43 0 2.17177e-19 $X=10.705 $Y=1.91
c174 36 0 1.49262e-19 $X=10.705 $Y=2.265
r175 73 74 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=13.8 $Y=1.33
+ $X2=13.8 $Y2=1.255
r176 70 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.8 $Y=1.42
+ $X2=13.8 $Y2=1.585
r177 70 73 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=13.8 $Y=1.42 $X2=13.8
+ $Y2=1.33
r178 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.8
+ $Y=1.42 $X2=13.8 $Y2=1.42
r179 66 69 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=13.695 $Y=1.42
+ $X2=13.8 $Y2=1.42
r180 61 63 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=12.105 $Y=1.37
+ $X2=12.235 $Y2=1.37
r181 56 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.695 $Y=1.585
+ $X2=13.695 $Y2=1.42
r182 56 57 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=13.695 $Y=1.585
+ $X2=13.695 $Y2=2.33
r183 55 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.32 $Y=2.415
+ $X2=12.235 $Y2=2.415
r184 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.61 $Y=2.415
+ $X2=13.695 $Y2=2.33
r185 54 55 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=13.61 $Y=2.415
+ $X2=12.32 $Y2=2.415
r186 53 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.235 $Y=2.33
+ $X2=12.235 $Y2=2.415
r187 52 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.235 $Y=1.535
+ $X2=12.235 $Y2=1.37
r188 52 53 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=12.235 $Y=1.535
+ $X2=12.235 $Y2=2.33
r189 51 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.85 $Y=2.415
+ $X2=11.685 $Y2=2.415
r190 50 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.15 $Y=2.415
+ $X2=12.235 $Y2=2.415
r191 50 51 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.15 $Y=2.415
+ $X2=11.85 $Y2=2.415
r192 46 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.52 $Y=2.415
+ $X2=11.685 $Y2=2.415
r193 46 47 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=11.52 $Y=2.415
+ $X2=10.87 $Y2=2.415
r194 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.705
+ $Y=1.91 $X2=10.705 $Y2=1.91
r195 41 47 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=10.722 $Y=2.33
+ $X2=10.87 $Y2=2.415
r196 41 43 16.4077 $w=2.93e-07 $l=4.2e-07 $layer=LI1_cond $X=10.722 $Y=2.33
+ $X2=10.722 $Y2=1.91
r197 39 44 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.705 $Y=1.745
+ $X2=10.705 $Y2=1.91
r198 36 44 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=10.705 $Y=2.265
+ $X2=10.705 $Y2=1.91
r199 33 36 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=10.395 $Y=2.34
+ $X2=10.705 $Y2=2.34
r200 29 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.82 $Y=1.405
+ $X2=14.82 $Y2=1.33
r201 29 31 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=14.82 $Y=1.405
+ $X2=14.82 $Y2=2.155
r202 25 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.82 $Y=1.255
+ $X2=14.82 $Y2=1.33
r203 25 27 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=14.82 $Y=1.255
+ $X2=14.82 $Y2=0.895
r204 24 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.965 $Y=1.33
+ $X2=13.8 $Y2=1.33
r205 23 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.745 $Y=1.33
+ $X2=14.82 $Y2=1.33
r206 23 24 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=14.745 $Y=1.33
+ $X2=13.965 $Y2=1.33
r207 21 76 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=13.83 $Y=2.415
+ $X2=13.83 $Y2=1.585
r208 17 74 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=13.83 $Y=0.655
+ $X2=13.83 $Y2=1.255
r209 13 39 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=10.645 $Y=0.715
+ $X2=10.645 $Y2=1.745
r210 7 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.395 $Y=2.415
+ $X2=10.395 $Y2=2.34
r211 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.395 $Y=2.415
+ $X2=10.395 $Y2=2.785
r212 2 59 300 $w=1.7e-07 $l=3.32265e-07 $layer=licon1_PDIFF $count=2 $X=11.465
+ $Y=2.255 $X2=11.685 $Y2=2.495
r213 1 61 182 $w=1.7e-07 $l=1.21697e-06 $layer=licon1_NDIFF $count=1 $X=11.825
+ $Y=0.285 $X2=12.105 $Y2=1.37
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_1861_431# 1 2 9 13 15 17 22 24 25 28 29
+ 34 38 39
c121 39 0 5.60316e-21 $X=11.84 $Y=1.88
c122 17 0 1.77109e-19 $X=10.135 $Y=0.78
r123 39 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.84 $Y=1.88
+ $X2=11.84 $Y2=2.045
r124 39 42 47.9601 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=11.84 $Y=1.88
+ $X2=11.84 $Y2=1.705
r125 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.84
+ $Y=1.88 $X2=11.84 $Y2=1.88
r126 35 38 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.675 $Y=1.88
+ $X2=11.84 $Y2=1.88
r127 29 32 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=9.445 $Y=2.68
+ $X2=9.445 $Y2=2.805
r128 28 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.675 $Y=1.715
+ $X2=11.675 $Y2=1.88
r129 27 28 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=11.675 $Y=1.52
+ $X2=11.675 $Y2=1.715
r130 26 34 1.34256 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.395 $Y=1.435
+ $X2=10.265 $Y2=1.435
r131 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.59 $Y=1.435
+ $X2=11.675 $Y2=1.52
r132 25 26 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=11.59 $Y=1.435
+ $X2=10.395 $Y2=1.435
r133 23 34 5.16603 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=10.31 $Y=1.52
+ $X2=10.265 $Y2=1.435
r134 23 24 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=10.31 $Y=1.52
+ $X2=10.31 $Y2=2.595
r135 22 34 5.16603 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=10.22 $Y=1.35
+ $X2=10.265 $Y2=1.435
r136 21 22 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=10.22 $Y=0.945
+ $X2=10.22 $Y2=1.35
r137 17 21 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.135 $Y=0.78
+ $X2=10.22 $Y2=0.945
r138 17 19 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=10.135 $Y=0.78
+ $X2=9.96 $Y2=0.78
r139 16 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.61 $Y=2.68
+ $X2=9.445 $Y2=2.68
r140 15 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.225 $Y=2.68
+ $X2=10.31 $Y2=2.595
r141 15 16 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=10.225 $Y=2.68
+ $X2=9.61 $Y2=2.68
r142 13 43 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=11.9 $Y=2.675
+ $X2=11.9 $Y2=2.045
r143 9 42 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=11.75 $Y=0.605
+ $X2=11.75 $Y2=1.705
r144 2 32 600 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=1 $X=9.305
+ $Y=2.155 $X2=9.445 $Y2=2.805
r145 1 19 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=9.82
+ $Y=0.285 $X2=9.96 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%RESET_B 3 6 8 11 13
r35 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.23 $Y=1.35
+ $X2=13.23 $Y2=1.515
r36 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.23 $Y=1.35
+ $X2=13.23 $Y2=1.185
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.23
+ $Y=1.35 $X2=13.23 $Y2=1.35
r38 6 14 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=13.32 $Y=2.105
+ $X2=13.32 $Y2=1.515
r39 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.32 $Y=0.865
+ $X2=13.32 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_2892_137# 1 2 9 13 17 21 25 26 28
c52 21 0 1.84272e-19 $X=14.605 $Y=1.98
r53 26 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.27 $Y=1.47
+ $X2=15.27 $Y2=1.635
r54 26 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.27 $Y=1.47
+ $X2=15.27 $Y2=1.305
r55 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.27
+ $Y=1.47 $X2=15.27 $Y2=1.47
r56 23 28 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=14.77 $Y=1.47
+ $X2=14.645 $Y2=1.47
r57 23 25 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=14.77 $Y=1.47
+ $X2=15.27 $Y2=1.47
r58 19 28 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=14.645 $Y=1.635
+ $X2=14.645 $Y2=1.47
r59 19 21 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=14.645 $Y=1.635
+ $X2=14.645 $Y2=1.98
r60 15 28 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=14.645 $Y=1.305
+ $X2=14.645 $Y2=1.47
r61 15 17 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=14.645 $Y=1.305
+ $X2=14.645 $Y2=0.895
r62 13 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=15.33 $Y=2.465
+ $X2=15.33 $Y2=1.635
r63 9 30 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=15.33 $Y=0.685
+ $X2=15.33 $Y2=1.305
r64 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=14.46
+ $Y=1.835 $X2=14.605 $Y2=1.98
r65 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=14.46
+ $Y=0.685 $X2=14.605 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_27_481# 1 2 9 11 12 14 15 16 19
c50 16 0 2.49076e-20 $X=1.305 $Y=2.98
c51 9 0 4.55157e-20 $X=0.28 $Y=2.55
r52 17 19 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.16 $Y=2.895
+ $X2=2.16 $Y2=2.55
r53 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.995 $Y=2.98
+ $X2=2.16 $Y2=2.895
r54 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.995 $Y=2.98
+ $X2=1.305 $Y2=2.98
r55 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.22 $Y=2.895
+ $X2=1.305 $Y2=2.98
r56 13 14 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.22 $Y=2.235
+ $X2=1.22 $Y2=2.895
r57 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.135 $Y=2.15
+ $X2=1.22 $Y2=2.235
r58 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.135 $Y=2.15
+ $X2=0.445 $Y2=2.15
r59 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.235
+ $X2=0.445 $Y2=2.15
r60 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.28 $Y=2.235
+ $X2=0.28 $Y2=2.55
r61 2 19 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=1.94
+ $Y=2.405 $X2=2.16 $Y2=2.55
r62 1 9 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.405 $X2=0.28 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 39 43 47 51
+ 55 59 63 67 71 76 77 79 80 82 83 84 86 91 106 110 115 127 136 137 140 143 146
+ 149 152 155 158
r187 158 159 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r188 155 156 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r189 152 153 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r190 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r191 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r192 144 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r193 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r194 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r196 134 137 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.6 $Y2=3.33
r197 134 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=13.68 $Y2=3.33
r198 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r199 131 158 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.78 $Y=3.33
+ $X2=13.615 $Y2=3.33
r200 131 133 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=13.78 $Y=3.33
+ $X2=14.64 $Y2=3.33
r201 130 159 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r202 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r203 127 158 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.45 $Y=3.33
+ $X2=13.615 $Y2=3.33
r204 127 129 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.45 $Y=3.33
+ $X2=13.2 $Y2=3.33
r205 126 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=13.2 $Y2=3.33
r206 126 156 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r207 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r208 123 155 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.34 $Y=3.33
+ $X2=11.175 $Y2=3.33
r209 123 125 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=11.34 $Y=3.33
+ $X2=12.24 $Y2=3.33
r210 122 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r211 121 122 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r212 119 122 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r213 119 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r214 118 121 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r215 118 119 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r216 116 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=3.33
+ $X2=8.54 $Y2=3.33
r217 116 118 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=8.705 $Y=3.33
+ $X2=8.88 $Y2=3.33
r218 115 155 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.01 $Y=3.33
+ $X2=11.175 $Y2=3.33
r219 115 121 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.01 $Y=3.33
+ $X2=10.8 $Y2=3.33
r220 114 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r221 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r222 111 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.285 $Y=3.33
+ $X2=7.12 $Y2=3.33
r223 111 113 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.285 $Y=3.33
+ $X2=7.44 $Y2=3.33
r224 110 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=8.54 $Y2=3.33
r225 110 113 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=7.44 $Y2=3.33
r226 109 150 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.96 $Y2=3.33
r227 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r228 106 149 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=7.12 $Y2=3.33
r229 106 108 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=5.52 $Y2=3.33
r230 105 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r231 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r232 102 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r233 102 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r234 101 104 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r235 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r236 99 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.71 $Y2=3.33
r237 99 101 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.08 $Y2=3.33
r238 98 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r239 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r240 95 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r241 95 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r242 94 97 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r243 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r244 92 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.79 $Y2=3.33
r245 92 94 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.2 $Y2=3.33
r246 91 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.68 $Y2=3.33
r247 91 97 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.16 $Y2=3.33
r248 89 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r249 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r250 86 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.79 $Y2=3.33
r251 86 88 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r252 84 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r253 84 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r254 82 133 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=14.95 $Y=3.33
+ $X2=14.64 $Y2=3.33
r255 82 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.95 $Y=3.33
+ $X2=15.075 $Y2=3.33
r256 81 136 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=15.2 $Y=3.33
+ $X2=15.6 $Y2=3.33
r257 81 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.2 $Y=3.33
+ $X2=15.075 $Y2=3.33
r258 79 125 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=12.37 $Y=3.33
+ $X2=12.24 $Y2=3.33
r259 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.37 $Y=3.33
+ $X2=12.535 $Y2=3.33
r260 78 129 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=12.7 $Y=3.33
+ $X2=13.2 $Y2=3.33
r261 78 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.7 $Y=3.33
+ $X2=12.535 $Y2=3.33
r262 76 104 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=5.04 $Y2=3.33
r263 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=5.21 $Y2=3.33
r264 75 108 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.375 $Y=3.33
+ $X2=5.52 $Y2=3.33
r265 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=3.33
+ $X2=5.21 $Y2=3.33
r266 71 74 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=15.075 $Y=1.98
+ $X2=15.075 $Y2=2.465
r267 69 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.075 $Y=3.245
+ $X2=15.075 $Y2=3.33
r268 69 74 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=15.075 $Y=3.245
+ $X2=15.075 $Y2=2.465
r269 65 158 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.615 $Y=3.245
+ $X2=13.615 $Y2=3.33
r270 65 67 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=13.615 $Y=3.245
+ $X2=13.615 $Y2=2.87
r271 61 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.535 $Y=3.245
+ $X2=12.535 $Y2=3.33
r272 61 63 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=12.535 $Y=3.245
+ $X2=12.535 $Y2=2.895
r273 57 155 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.175 $Y=3.245
+ $X2=11.175 $Y2=3.33
r274 57 59 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=11.175 $Y=3.245
+ $X2=11.175 $Y2=2.895
r275 53 152 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.54 $Y=3.245
+ $X2=8.54 $Y2=3.33
r276 53 55 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=8.54 $Y=3.245
+ $X2=8.54 $Y2=2.515
r277 49 149 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.12 $Y=3.245
+ $X2=7.12 $Y2=3.33
r278 49 51 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=7.12 $Y=3.245 $X2=7.12
+ $Y2=2.845
r279 45 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.21 $Y=3.245
+ $X2=5.21 $Y2=3.33
r280 45 47 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=5.21 $Y=3.245
+ $X2=5.21 $Y2=2.43
r281 41 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=3.33
r282 41 43 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=2.515
r283 40 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.68 $Y2=3.33
r284 39 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=3.71 $Y2=3.33
r285 39 40 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=2.805 $Y2=3.33
r286 35 143 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=3.33
r287 35 37 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=2.55
r288 31 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=3.33
r289 31 33 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=2.74
r290 10 74 300 $w=1.7e-07 $l=7.31779e-07 $layer=licon1_PDIFF $count=2 $X=14.895
+ $Y=1.835 $X2=15.115 $Y2=2.465
r291 10 71 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=14.895
+ $Y=1.835 $X2=15.115 $Y2=1.98
r292 9 67 600 $w=1.7e-07 $l=1.18993e-06 $layer=licon1_PDIFF $count=1 $X=13.395
+ $Y=1.785 $X2=13.615 $Y2=2.87
r293 8 63 600 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=1 $X=12.395
+ $Y=2.255 $X2=12.535 $Y2=2.895
r294 7 59 600 $w=1.7e-07 $l=8.50074e-07 $layer=licon1_PDIFF $count=1 $X=10.47
+ $Y=2.575 $X2=11.175 $Y2=2.895
r295 6 55 600 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=1 $X=8.4
+ $Y=1.865 $X2=8.54 $Y2=2.515
r296 5 51 600 $w=1.7e-07 $l=6.60908e-07 $layer=licon1_PDIFF $count=1 $X=6.9
+ $Y=2.285 $X2=7.12 $Y2=2.845
r297 4 47 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=2.285 $X2=5.21 $Y2=2.43
r298 3 43 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.565
+ $Y=2.37 $X2=3.71 $Y2=2.515
r299 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.575
+ $Y=2.405 $X2=2.72 $Y2=2.55
r300 1 33 600 $w=1.7e-07 $l=4.3119e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.405 $X2=0.79 $Y2=2.74
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_204_119# 1 2 3 4 15 17 18 21 24 26 27 28
+ 30 31 32 34 35 36 38 39 40 43 49 52 55 56 58
c182 56 0 7.21799e-20 $X=5.79 $Y=2.265
c183 49 0 2.47968e-19 $X=2.06 $Y=2.12
c184 43 0 6.11734e-20 $X=5.87 $Y=0.47
c185 24 0 1.50206e-19 $X=2.06 $Y=2.035
c186 21 0 1.8478e-19 $X=1.65 $Y=2.55
c187 18 0 3.63052e-20 $X=1.325 $Y=1.26
r188 55 56 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.79 $Y=2.495
+ $X2=5.79 $Y2=2.265
r189 51 52 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.06 $Y=1.26
+ $X2=2.3 $Y2=1.26
r190 45 58 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.87 $Y=1
+ $X2=5.83 $Y2=0.915
r191 45 56 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=5.87 $Y=1
+ $X2=5.87 $Y2=2.265
r192 41 58 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=0.83 $X2=5.83
+ $Y2=0.915
r193 41 43 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=5.83 $Y=0.83
+ $X2=5.83 $Y2=0.47
r194 39 58 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.705 $Y=0.915
+ $X2=5.83 $Y2=0.915
r195 39 40 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.705 $Y=0.915
+ $X2=5.045 $Y2=0.915
r196 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.96 $Y=0.83
+ $X2=5.045 $Y2=0.915
r197 37 38 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.96 $Y=0.435
+ $X2=4.96 $Y2=0.83
r198 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.875 $Y=0.35
+ $X2=4.96 $Y2=0.435
r199 35 36 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=4.875 $Y=0.35
+ $X2=3.785 $Y2=0.35
r200 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.7 $Y=0.435
+ $X2=3.785 $Y2=0.35
r201 33 34 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.7 $Y=0.435
+ $X2=3.7 $Y2=1.15
r202 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.615 $Y=1.235
+ $X2=3.7 $Y2=1.15
r203 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.615 $Y=1.235
+ $X2=3.085 $Y2=1.235
r204 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3 $Y=1.15
+ $X2=3.085 $Y2=1.235
r205 29 30 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3 $Y=0.435 $X2=3
+ $Y2=1.15
r206 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.915 $Y=0.35
+ $X2=3 $Y2=0.435
r207 27 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.915 $Y=0.35
+ $X2=2.385 $Y2=0.35
r208 26 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=1.175
+ $X2=2.3 $Y2=1.26
r209 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.3 $Y=0.435
+ $X2=2.385 $Y2=0.35
r210 25 26 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.3 $Y=0.435
+ $X2=2.3 $Y2=1.175
r211 24 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=2.035
+ $X2=2.06 $Y2=2.12
r212 23 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=1.345
+ $X2=2.06 $Y2=1.26
r213 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.06 $Y=1.345
+ $X2=2.06 $Y2=2.035
r214 19 49 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.65 $Y=2.12
+ $X2=2.06 $Y2=2.12
r215 19 21 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.65 $Y=2.205
+ $X2=1.65 $Y2=2.55
r216 17 51 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=1.26
+ $X2=2.06 $Y2=1.26
r217 17 18 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.975 $Y=1.26
+ $X2=1.325 $Y2=1.26
r218 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.16 $Y=1.175
+ $X2=1.325 $Y2=1.26
r219 13 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.16 $Y=1.175
+ $X2=1.16 $Y2=0.805
r220 4 55 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.645
+ $Y=2.285 $X2=5.79 $Y2=2.495
r221 3 21 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=2.405 $X2=1.65 $Y2=2.55
r222 2 43 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=5.725
+ $Y=0.235 $X2=5.87 $Y2=0.47
r223 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.595 $X2=1.16 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%Q_N 1 2 9 13 16 17 18 19 20
r34 20 31 4.0579 $w=3.53e-07 $l=1.25e-07 $layer=LI1_cond $X=14.137 $Y=2.775
+ $X2=14.137 $Y2=2.9
r35 19 20 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=14.137 $Y=2.405
+ $X2=14.137 $Y2=2.775
r36 18 19 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=14.137 $Y=2.035
+ $X2=14.137 $Y2=2.405
r37 16 17 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=14.137 $Y=1.93
+ $X2=14.137 $Y2=1.765
r38 14 18 3.01908 $w=3.53e-07 $l=9.3e-08 $layer=LI1_cond $X=14.137 $Y=1.942
+ $X2=14.137 $Y2=2.035
r39 14 16 0.389558 $w=3.53e-07 $l=1.2e-08 $layer=LI1_cond $X=14.137 $Y=1.942
+ $X2=14.137 $Y2=1.93
r40 13 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.23 $Y=1.075
+ $X2=14.23 $Y2=1.765
r41 7 13 10.1875 $w=4.33e-07 $l=2.17e-07 $layer=LI1_cond $X=14.097 $Y=0.858
+ $X2=14.097 $Y2=1.075
r42 7 9 11.339 $w=4.33e-07 $l=4.28e-07 $layer=LI1_cond $X=14.097 $Y=0.858
+ $X2=14.097 $Y2=0.43
r43 2 31 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=13.905
+ $Y=1.785 $X2=14.045 $Y2=2.9
r44 2 16 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.905
+ $Y=1.785 $X2=14.045 $Y2=1.93
r45 1 9 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=13.905
+ $Y=0.235 $X2=14.045 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%Q 1 2 9 14 15 16 17 23 29
r25 21 29 0.467207 $w=3.68e-07 $l=1.5e-08 $layer=LI1_cond $X=15.565 $Y=0.94
+ $X2=15.565 $Y2=0.925
r26 17 31 8.0716 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=15.565 $Y=0.975
+ $X2=15.565 $Y2=1.125
r27 17 21 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=15.565 $Y=0.975
+ $X2=15.565 $Y2=0.94
r28 17 29 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=15.565 $Y=0.89
+ $X2=15.565 $Y2=0.925
r29 16 17 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=15.565 $Y=0.555
+ $X2=15.565 $Y2=0.89
r30 16 23 3.89339 $w=3.68e-07 $l=1.25e-07 $layer=LI1_cond $X=15.565 $Y=0.555
+ $X2=15.565 $Y2=0.43
r31 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=15.665 $Y=1.815
+ $X2=15.665 $Y2=1.125
r32 14 15 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=15.565 $Y=1.98
+ $X2=15.565 $Y2=1.815
r33 7 14 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=15.565 $Y=2 $X2=15.565
+ $Y2=1.98
r34 7 9 28.0324 $w=3.68e-07 $l=9e-07 $layer=LI1_cond $X=15.565 $Y=2 $X2=15.565
+ $Y2=2.9
r35 2 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.405
+ $Y=1.835 $X2=15.545 $Y2=1.98
r36 2 9 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=15.405
+ $Y=1.835 $X2=15.545 $Y2=2.9
r37 1 23 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=15.405
+ $Y=0.265 $X2=15.545 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 54 58 64 69 70 72 73 75 76 78 79 81 82 84 85 87 88 89 128 140 141 147
r184 147 148 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r185 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r186 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r187 138 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.6 $Y2=0
r188 138 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=13.68 $Y2=0
r189 137 138 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r190 135 147 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.7 $Y=0
+ $X2=13.575 $Y2=0
r191 135 137 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=13.7 $Y=0
+ $X2=14.64 $Y2=0
r192 134 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r193 133 134 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r194 131 134 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=13.2 $Y2=0
r195 130 133 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=13.2 $Y2=0
r196 130 131 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r197 128 147 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.45 $Y=0
+ $X2=13.575 $Y2=0
r198 128 133 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.45 $Y=0
+ $X2=13.2 $Y2=0
r199 127 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r200 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r201 124 127 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r202 123 126 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r203 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r204 121 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r205 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r206 117 120 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=7.44 $Y=0
+ $X2=8.88 $Y2=0
r207 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r208 115 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r209 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r210 112 115 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.96 $Y2=0
r211 111 114 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.52 $Y=0
+ $X2=6.96 $Y2=0
r212 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r213 109 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r214 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r215 106 109 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=5.04 $Y2=0
r216 105 108 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0
+ $X2=5.04 $Y2=0
r217 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r218 103 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=3.6 $Y2=0
r219 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r220 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=3.12 $Y2=0
r221 99 102 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r222 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r223 97 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r224 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r225 94 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r226 94 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r227 93 96 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r228 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r229 91 144 4.61231 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.252 $Y2=0
r230 91 93 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.505 $Y=0
+ $X2=0.72 $Y2=0
r231 89 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.88 $Y2=0
r232 89 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r233 87 137 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=14.95 $Y=0
+ $X2=14.64 $Y2=0
r234 87 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.95 $Y=0
+ $X2=15.075 $Y2=0
r235 86 140 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=15.2 $Y=0 $X2=15.6
+ $Y2=0
r236 86 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.2 $Y=0
+ $X2=15.075 $Y2=0
r237 84 126 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=10.86 $Y=0 $X2=10.8
+ $Y2=0
r238 84 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.86 $Y=0
+ $X2=11.025 $Y2=0
r239 83 130 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=11.19 $Y=0 $X2=11.28
+ $Y2=0
r240 83 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.19 $Y=0
+ $X2=11.025 $Y2=0
r241 81 120 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=8.935 $Y=0
+ $X2=8.88 $Y2=0
r242 81 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.935 $Y=0 $X2=9.1
+ $Y2=0
r243 80 123 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=9.265 $Y=0
+ $X2=9.36 $Y2=0
r244 80 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.265 $Y=0 $X2=9.1
+ $Y2=0
r245 78 114 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=6.96 $Y2=0
r246 78 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.005 $Y=0 $X2=7.13
+ $Y2=0
r247 77 117 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.255 $Y=0
+ $X2=7.44 $Y2=0
r248 77 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.255 $Y=0 $X2=7.13
+ $Y2=0
r249 75 108 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.225 $Y=0
+ $X2=5.04 $Y2=0
r250 75 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.35
+ $Y2=0
r251 74 111 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.475 $Y=0
+ $X2=5.52 $Y2=0
r252 74 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.475 $Y=0 $X2=5.35
+ $Y2=0
r253 72 102 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=0
+ $X2=3.12 $Y2=0
r254 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.35
+ $Y2=0
r255 71 105 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0
+ $X2=3.6 $Y2=0
r256 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.35
+ $Y2=0
r257 69 96 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=1.68 $Y2=0
r258 69 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.91
+ $Y2=0
r259 68 99 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=0
+ $X2=2.16 $Y2=0
r260 68 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.91
+ $Y2=0
r261 64 66 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=15.075 $Y=0.41
+ $X2=15.075 $Y2=0.96
r262 62 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.075 $Y=0.085
+ $X2=15.075 $Y2=0
r263 62 64 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=15.075 $Y=0.085
+ $X2=15.075 $Y2=0.41
r264 58 60 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=13.575 $Y=0.38
+ $X2=13.575 $Y2=0.835
r265 56 147 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.575 $Y=0.085
+ $X2=13.575 $Y2=0
r266 56 58 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=13.575 $Y=0.085
+ $X2=13.575 $Y2=0.38
r267 52 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.025 $Y=0.085
+ $X2=11.025 $Y2=0
r268 52 54 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=11.025 $Y=0.085
+ $X2=11.025 $Y2=0.54
r269 48 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.1 $Y=0.085 $X2=9.1
+ $Y2=0
r270 48 50 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.1 $Y=0.085
+ $X2=9.1 $Y2=0.47
r271 44 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.13 $Y=0.085
+ $X2=7.13 $Y2=0
r272 44 46 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=7.13 $Y=0.085
+ $X2=7.13 $Y2=0.53
r273 40 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.35 $Y=0.085
+ $X2=5.35 $Y2=0
r274 40 42 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=5.35 $Y=0.085
+ $X2=5.35 $Y2=0.485
r275 36 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0
r276 36 38 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.35 $Y=0.085
+ $X2=3.35 $Y2=0.74
r277 32 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.91 $Y=0.085
+ $X2=1.91 $Y2=0
r278 32 34 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=1.91 $Y=0.085
+ $X2=1.91 $Y2=0.785
r279 28 144 3.15387 $w=3.3e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.252 $Y2=0
r280 28 30 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.34 $Y2=0.805
r281 9 66 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=14.895
+ $Y=0.685 $X2=15.115 $Y2=0.96
r282 9 64 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=14.895
+ $Y=0.685 $X2=15.115 $Y2=0.41
r283 8 60 182 $w=1.7e-07 $l=2.96648e-07 $layer=licon1_NDIFF $count=1 $X=13.395
+ $Y=0.655 $X2=13.615 $Y2=0.835
r284 8 58 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=13.395
+ $Y=0.655 $X2=13.615 $Y2=0.38
r285 7 54 182 $w=1.7e-07 $l=3.22025e-07 $layer=licon1_NDIFF $count=1 $X=10.72
+ $Y=0.505 $X2=11.025 $Y2=0.54
r286 6 50 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=8.955
+ $Y=0.285 $X2=9.1 $Y2=0.47
r287 5 46 182 $w=1.7e-07 $l=3.89776e-07 $layer=licon1_NDIFF $count=1 $X=6.95
+ $Y=0.235 $X2=7.17 $Y2=0.53
r288 4 42 182 $w=1.7e-07 $l=4.19881e-07 $layer=licon1_NDIFF $count=1 $X=4.9
+ $Y=0.505 $X2=5.31 $Y2=0.485
r289 3 38 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.53 $X2=3.35 $Y2=0.74
r290 2 34 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.81
+ $Y=0.595 $X2=1.95 $Y2=0.785
r291 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.195
+ $Y=0.595 $X2=0.34 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_1492_47# 1 2 7 10 12
c26 12 0 1.67734e-19 $X=8.54 $Y=0.38
r27 10 12 42.9773 $w=1.98e-07 $l=7.75e-07 $layer=LI1_cond $X=7.765 $Y=0.365
+ $X2=8.54 $Y2=0.365
r28 7 10 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=7.6 $Y=0.465
+ $X2=7.765 $Y2=0.365
r29 7 9 3.32727 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.6 $Y=0.465 $X2=7.6
+ $Y2=0.555
r30 2 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.4
+ $Y=0.235 $X2=8.54 $Y2=0.38
r31 1 9 182 $w=1.7e-07 $l=3.83667e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.6 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__SDFBBP_1%A_2279_57# 1 2 7 9 14
c28 7 0 1.19113e-20 $X=12.4 $Y=0.35
c29 2 0 1.8236e-19 $X=12.425 $Y=0.285
r30 14 17 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=12.525 $Y=0.35
+ $X2=12.525 $Y2=0.455
r31 9 12 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=11.535 $Y=0.35
+ $X2=11.535 $Y2=0.455
r32 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.7 $Y=0.35
+ $X2=11.535 $Y2=0.35
r33 7 14 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.4 $Y=0.35
+ $X2=12.525 $Y2=0.35
r34 7 8 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=12.4 $Y=0.35 $X2=11.7
+ $Y2=0.35
r35 2 17 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=12.425
+ $Y=0.285 $X2=12.565 $Y2=0.455
r36 1 12 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=11.395
+ $Y=0.285 $X2=11.535 $Y2=0.455
.ends

