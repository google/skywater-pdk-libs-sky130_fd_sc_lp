* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor2_8 A B VGND VNB VPB VPWR Y
X0 VPWR A a_47_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_47_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_47_367# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_47_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_47_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 Y B a_47_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 Y B a_47_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_47_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VPWR A a_47_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 Y B a_47_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_47_367# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 Y B a_47_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 VPWR A a_47_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VPWR A a_47_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_47_367# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_47_367# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
