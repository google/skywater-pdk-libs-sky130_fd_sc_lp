# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__nor4b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.960000 1.355000 9.030000 1.525000 ;
        RECT 7.735000 1.210000 9.030000 1.355000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.230000 1.355000 6.625000 1.835000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.010000 1.315000 4.700000 1.485000 ;
        RECT 3.885000 1.210000 4.700000 1.315000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.325000 0.550000 1.760000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  2.612400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.095000 0.255000 1.295000 0.965000 ;
        RECT 1.095000 0.965000 5.615000 1.005000 ;
        RECT 1.095000 1.005000 8.235000 1.040000 ;
        RECT 1.095000 1.040000 3.405000 1.145000 ;
        RECT 1.475000 1.665000 5.060000 1.835000 ;
        RECT 1.475000 1.835000 1.805000 2.735000 ;
        RECT 1.965000 0.255000 2.185000 0.965000 ;
        RECT 2.335000 1.835000 2.665000 2.735000 ;
        RECT 3.205000 0.255000 3.395000 0.840000 ;
        RECT 3.205000 0.840000 5.615000 0.965000 ;
        RECT 4.065000 0.255000 4.255000 0.840000 ;
        RECT 4.870000 1.040000 7.425000 1.185000 ;
        RECT 4.870000 1.185000 5.060000 1.665000 ;
        RECT 5.425000 0.255000 5.615000 0.840000 ;
        RECT 6.285000 0.255000 6.475000 1.005000 ;
        RECT 7.145000 0.255000 7.375000 0.870000 ;
        RECT 7.145000 0.870000 8.235000 1.005000 ;
        RECT 8.045000 0.255000 8.235000 0.870000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.095000  1.930000 0.925000 2.100000 ;
      RECT 0.095000  2.100000 0.355000 3.075000 ;
      RECT 0.105000  0.255000 0.365000 0.985000 ;
      RECT 0.105000  0.985000 0.925000 1.155000 ;
      RECT 0.525000  2.270000 0.855000 3.245000 ;
      RECT 0.535000  0.085000 0.865000 0.815000 ;
      RECT 0.720000  1.155000 0.925000 1.315000 ;
      RECT 0.720000  1.315000 2.800000 1.485000 ;
      RECT 0.720000  1.485000 0.925000 1.930000 ;
      RECT 1.095000  1.815000 1.305000 2.905000 ;
      RECT 1.095000  2.905000 4.815000 3.075000 ;
      RECT 1.465000  0.085000 1.795000 0.795000 ;
      RECT 1.975000  2.005000 2.165000 2.905000 ;
      RECT 2.355000  0.085000 3.035000 0.785000 ;
      RECT 2.835000  2.005000 3.025000 2.905000 ;
      RECT 3.195000  2.005000 6.625000 2.185000 ;
      RECT 3.195000  2.185000 3.525000 2.735000 ;
      RECT 3.565000  0.085000 3.895000 0.670000 ;
      RECT 3.695000  2.355000 3.895000 2.905000 ;
      RECT 4.115000  2.185000 4.315000 2.735000 ;
      RECT 4.425000  0.085000 5.255000 0.670000 ;
      RECT 4.485000  2.355000 4.815000 2.905000 ;
      RECT 5.005000  2.355000 5.335000 2.905000 ;
      RECT 5.005000  2.905000 6.985000 3.075000 ;
      RECT 5.505000  2.185000 5.730000 2.735000 ;
      RECT 5.785000  0.085000 6.115000 0.835000 ;
      RECT 5.900000  2.355000 6.125000 2.905000 ;
      RECT 6.295000  2.185000 6.625000 2.735000 ;
      RECT 6.645000  0.085000 6.975000 0.835000 ;
      RECT 6.795000  1.695000 8.775000 1.925000 ;
      RECT 6.795000  1.925000 6.985000 2.905000 ;
      RECT 7.155000  2.105000 7.485000 3.245000 ;
      RECT 7.545000  0.085000 7.875000 0.700000 ;
      RECT 7.655000  1.925000 7.845000 3.075000 ;
      RECT 8.015000  2.105000 8.345000 3.245000 ;
      RECT 8.405000  0.085000 8.735000 1.040000 ;
      RECT 8.515000  1.925000 8.775000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_lp__nor4b_4
