* File: sky130_fd_sc_lp__o2bb2a_lp.pxi.spice
* Created: Fri Aug 28 11:12:09 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%A_86_22# N_A_86_22#_M1012_s N_A_86_22#_M1000_d
+ N_A_86_22#_M1009_g N_A_86_22#_c_80_n N_A_86_22#_M1005_g N_A_86_22#_M1006_g
+ N_A_86_22#_c_83_n N_A_86_22#_c_84_n N_A_86_22#_c_101_p N_A_86_22#_c_146_p
+ N_A_86_22#_c_91_n N_A_86_22#_c_85_n N_A_86_22#_c_86_n N_A_86_22#_c_87_n
+ N_A_86_22#_c_121_p N_A_86_22#_c_88_n PM_SKY130_FD_SC_LP__O2BB2A_LP%A_86_22#
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%A1_N N_A1_N_M1010_g N_A1_N_M1007_g A1_N A1_N
+ N_A1_N_c_180_n PM_SKY130_FD_SC_LP__O2BB2A_LP%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%A2_N N_A2_N_c_222_n N_A2_N_M1011_g
+ N_A2_N_M1004_g N_A2_N_c_223_n N_A2_N_c_224_n N_A2_N_c_225_n N_A2_N_c_230_n
+ A2_N A2_N N_A2_N_c_227_n PM_SKY130_FD_SC_LP__O2BB2A_LP%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%A_298_416# N_A_298_416#_M1011_d
+ N_A_298_416#_M1007_d N_A_298_416#_c_267_n N_A_298_416#_M1000_g
+ N_A_298_416#_c_268_n N_A_298_416#_M1012_g N_A_298_416#_c_275_n
+ N_A_298_416#_c_269_n N_A_298_416#_c_270_n N_A_298_416#_c_276_n
+ N_A_298_416#_c_271_n N_A_298_416#_c_272_n N_A_298_416#_c_273_n
+ PM_SKY130_FD_SC_LP__O2BB2A_LP%A_298_416#
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%B2 N_B2_M1008_g N_B2_M1001_g N_B2_c_342_n
+ N_B2_c_343_n B2 N_B2_c_344_n N_B2_c_345_n N_B2_c_346_n
+ PM_SKY130_FD_SC_LP__O2BB2A_LP%B2
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%B1 N_B1_M1002_g N_B1_M1003_g B1 N_B1_c_391_n
+ PM_SKY130_FD_SC_LP__O2BB2A_LP%B1
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%X N_X_M1009_s N_X_M1005_s X X X X
+ PM_SKY130_FD_SC_LP__O2BB2A_LP%X
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%VPWR N_VPWR_M1005_d N_VPWR_M1004_d
+ N_VPWR_M1002_d N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n
+ VPWR N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n
+ N_VPWR_c_433_n PM_SKY130_FD_SC_LP__O2BB2A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%VGND N_VGND_M1006_d N_VGND_M1001_d
+ N_VGND_c_485_n N_VGND_c_486_n VGND N_VGND_c_487_n N_VGND_c_488_n
+ N_VGND_c_489_n N_VGND_c_490_n N_VGND_c_491_n N_VGND_c_492_n
+ PM_SKY130_FD_SC_LP__O2BB2A_LP%VGND
x_PM_SKY130_FD_SC_LP__O2BB2A_LP%A_604_142# N_A_604_142#_M1012_d
+ N_A_604_142#_M1003_d N_A_604_142#_c_535_n N_A_604_142#_c_536_n
+ N_A_604_142#_c_537_n N_A_604_142#_c_538_n
+ PM_SKY130_FD_SC_LP__O2BB2A_LP%A_604_142#
cc_1 VNB N_A_86_22#_M1009_g 0.0246094f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.45
cc_2 VNB N_A_86_22#_c_80_n 0.0108827f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.555
cc_3 VNB N_A_86_22#_M1005_g 0.00687791f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.58
cc_4 VNB N_A_86_22#_M1006_g 0.0197761f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.45
cc_5 VNB N_A_86_22#_c_83_n 0.0173463f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.43
cc_6 VNB N_A_86_22#_c_84_n 0.00631095f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.49
cc_7 VNB N_A_86_22#_c_85_n 0.00676923f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.945
cc_8 VNB N_A_86_22#_c_86_n 0.00546515f $X=-0.19 $Y=-0.245 $X2=2.67 $Y2=0.96
cc_9 VNB N_A_86_22#_c_87_n 0.0250001f $X=-0.19 $Y=-0.245 $X2=2.505 $Y2=0.962
cc_10 VNB N_A_86_22#_c_88_n 0.0442983f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.025
cc_11 VNB N_A1_N_M1010_g 0.0609631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A1_N 0.00355169f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.45
cc_13 VNB N_A1_N_c_180_n 0.0203892f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.45
cc_14 VNB N_A2_N_c_222_n 0.017521f $X=-0.19 $Y=-0.245 $X2=2.525 $Y2=0.71
cc_15 VNB N_A2_N_c_223_n 0.0167267f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.43
cc_16 VNB N_A2_N_c_224_n 0.0183495f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.58
cc_17 VNB N_A2_N_c_225_n 0.0170602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A2_N 0.0125762f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.45
cc_19 VNB N_A2_N_c_227_n 0.0150895f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.49
cc_20 VNB N_A_298_416#_c_267_n 0.0509905f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.45
cc_21 VNB N_A_298_416#_c_268_n 0.0232782f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.555
cc_22 VNB N_A_298_416#_c_269_n 0.00644008f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.19
cc_23 VNB N_A_298_416#_c_270_n 0.0643124f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.49
cc_24 VNB N_A_298_416#_c_271_n 0.00356283f $X=-0.19 $Y=-0.245 $X2=2.98 $Y2=2.225
cc_25 VNB N_A_298_416#_c_272_n 0.00418204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_298_416#_c_273_n 0.026132f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.19
cc_27 VNB N_B2_c_342_n 0.0150661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B2_c_343_n 0.0120988f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.19
cc_29 VNB N_B2_c_344_n 0.0107449f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.58
cc_30 VNB N_B2_c_345_n 0.00213201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B2_c_346_n 0.0148176f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.86
cc_32 VNB N_B1_M1003_g 0.0449664f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.86
cc_33 VNB B1 0.00779945f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.45
cc_34 VNB N_B1_c_391_n 0.0124328f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.43
cc_35 VNB X 0.0567851f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.86
cc_36 VNB N_VPWR_c_433_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_485_n 0.00321f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.45
cc_38 VNB N_VGND_c_486_n 0.0250089f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.555
cc_39 VNB N_VGND_c_487_n 0.0272205f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.86
cc_40 VNB N_VGND_c_488_n 0.0577777f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.19
cc_41 VNB N_VGND_c_489_n 0.022032f $X=-0.19 $Y=-0.245 $X2=2.98 $Y2=2.225
cc_42 VNB N_VGND_c_490_n 0.25662f $X=-0.19 $Y=-0.245 $X2=2.98 $Y2=2.225
cc_43 VNB N_VGND_c_491_n 0.00445561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_492_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.025
cc_45 VNB N_A_604_142#_c_535_n 0.00417146f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.45
cc_46 VNB N_A_604_142#_c_536_n 0.025076f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.19
cc_47 VNB N_A_604_142#_c_537_n 0.00351278f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.43
cc_48 VNB N_A_604_142#_c_538_n 0.0138987f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.58
cc_49 VPB N_A_86_22#_M1005_g 0.0499345f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.58
cc_50 VPB N_A_86_22#_c_84_n 0.00279221f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.49
cc_51 VPB N_A_86_22#_c_91_n 0.00768923f $X=-0.19 $Y=1.655 $X2=2.98 $Y2=2.225
cc_52 VPB N_A1_N_M1007_g 0.0304869f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.86
cc_53 VPB A1_N 0.00138214f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.45
cc_54 VPB N_A1_N_c_180_n 0.0279565f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.45
cc_55 VPB N_A2_N_M1004_g 0.0310123f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.45
cc_56 VPB N_A2_N_c_225_n 0.00343498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A2_N_c_230_n 0.0121406f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.86
cc_58 VPB A2_N 0.00682571f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.45
cc_59 VPB N_A_298_416#_M1000_g 0.033036f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.19
cc_60 VPB N_A_298_416#_c_275_n 0.00944064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_298_416#_c_276_n 0.00243462f $X=-0.19 $Y=1.655 $X2=2.505 $Y2=0.945
cc_62 VPB N_A_298_416#_c_273_n 0.024365f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.19
cc_63 VPB N_B2_M1008_g 0.0284778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_B2_c_344_n 0.0162589f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.58
cc_65 VPB N_B2_c_345_n 0.00383323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_B1_M1002_g 0.0358714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB B1 0.0137267f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.45
cc_68 VPB N_B1_c_391_n 0.0188255f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.43
cc_69 VPB X 0.0553309f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.86
cc_70 VPB N_VPWR_c_434_n 0.00329211f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.58
cc_71 VPB N_VPWR_c_435_n 0.00329119f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.45
cc_72 VPB N_VPWR_c_436_n 0.0110915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_437_n 0.0448783f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.19
cc_74 VPB N_VPWR_c_438_n 0.0277818f $X=-0.19 $Y=1.655 $X2=2.98 $Y2=2.49
cc_75 VPB N_VPWR_c_439_n 0.0424169f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_440_n 0.0241502f $X=-0.19 $Y=1.655 $X2=2.505 $Y2=0.962
cc_77 VPB N_VPWR_c_441_n 0.0052165f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.025
cc_78 VPB N_VPWR_c_433_n 0.0698416f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 N_A_86_22#_c_80_n N_A1_N_M1010_g 0.00194429f $X=0.555 $Y=1.555 $X2=0 $Y2=0
cc_80 N_A_86_22#_M1006_g N_A1_N_M1010_g 0.0172222f $X=0.865 $Y=0.45 $X2=0 $Y2=0
cc_81 N_A_86_22#_c_83_n N_A1_N_M1010_g 0.00256095f $X=0.555 $Y=1.43 $X2=0 $Y2=0
cc_82 N_A_86_22#_c_84_n N_A1_N_M1010_g 0.0062994f $X=0.72 $Y=2.49 $X2=0 $Y2=0
cc_83 N_A_86_22#_c_85_n N_A1_N_M1010_g 0.00113995f $X=0.8 $Y=0.945 $X2=0 $Y2=0
cc_84 N_A_86_22#_c_87_n N_A1_N_M1010_g 0.0147414f $X=2.505 $Y=0.962 $X2=0 $Y2=0
cc_85 N_A_86_22#_c_88_n N_A1_N_M1010_g 0.017448f $X=0.865 $Y=1.025 $X2=0 $Y2=0
cc_86 N_A_86_22#_M1005_g N_A1_N_M1007_g 0.0201575f $X=0.555 $Y=2.58 $X2=0 $Y2=0
cc_87 N_A_86_22#_c_84_n N_A1_N_M1007_g 0.00647036f $X=0.72 $Y=2.49 $X2=0 $Y2=0
cc_88 N_A_86_22#_c_101_p N_A1_N_M1007_g 0.0244636f $X=2.815 $Y=2.575 $X2=0 $Y2=0
cc_89 N_A_86_22#_c_80_n A1_N 3.43681e-19 $X=0.555 $Y=1.555 $X2=0 $Y2=0
cc_90 N_A_86_22#_M1005_g A1_N 8.54765e-19 $X=0.555 $Y=2.58 $X2=0 $Y2=0
cc_91 N_A_86_22#_c_84_n A1_N 0.0441124f $X=0.72 $Y=2.49 $X2=0 $Y2=0
cc_92 N_A_86_22#_c_101_p A1_N 0.0127041f $X=2.815 $Y=2.575 $X2=0 $Y2=0
cc_93 N_A_86_22#_c_87_n A1_N 0.0107616f $X=2.505 $Y=0.962 $X2=0 $Y2=0
cc_94 N_A_86_22#_c_80_n N_A1_N_c_180_n 0.013043f $X=0.555 $Y=1.555 $X2=0 $Y2=0
cc_95 N_A_86_22#_c_84_n N_A1_N_c_180_n 0.00228665f $X=0.72 $Y=2.49 $X2=0 $Y2=0
cc_96 N_A_86_22#_c_101_p N_A1_N_c_180_n 8.51332e-19 $X=2.815 $Y=2.575 $X2=0
+ $Y2=0
cc_97 N_A_86_22#_c_87_n N_A1_N_c_180_n 0.00470852f $X=2.505 $Y=0.962 $X2=0 $Y2=0
cc_98 N_A_86_22#_c_101_p N_A2_N_M1004_g 0.0184089f $X=2.815 $Y=2.575 $X2=0 $Y2=0
cc_99 N_A_86_22#_c_87_n N_A2_N_c_223_n 0.00776319f $X=2.505 $Y=0.962 $X2=0 $Y2=0
cc_100 N_A_86_22#_c_87_n N_A2_N_c_224_n 0.0084268f $X=2.505 $Y=0.962 $X2=0 $Y2=0
cc_101 N_A_86_22#_c_87_n A2_N 0.0551953f $X=2.505 $Y=0.962 $X2=0 $Y2=0
cc_102 N_A_86_22#_c_87_n N_A2_N_c_227_n 0.00470746f $X=2.505 $Y=0.962 $X2=0
+ $Y2=0
cc_103 N_A_86_22#_c_101_p N_A_298_416#_M1007_d 0.00567691f $X=2.815 $Y=2.575
+ $X2=0 $Y2=0
cc_104 N_A_86_22#_c_86_n N_A_298_416#_c_267_n 0.00587058f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_105 N_A_86_22#_c_87_n N_A_298_416#_c_267_n 0.0166871f $X=2.505 $Y=0.962 $X2=0
+ $Y2=0
cc_106 N_A_86_22#_c_101_p N_A_298_416#_M1000_g 0.0183397f $X=2.815 $Y=2.575
+ $X2=0 $Y2=0
cc_107 N_A_86_22#_c_91_n N_A_298_416#_M1000_g 0.0144644f $X=2.98 $Y=2.225 $X2=0
+ $Y2=0
cc_108 N_A_86_22#_c_121_p N_A_298_416#_M1000_g 0.0156215f $X=2.98 $Y=2.575 $X2=0
+ $Y2=0
cc_109 N_A_86_22#_c_86_n N_A_298_416#_c_268_n 0.00238035f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_110 N_A_86_22#_c_101_p N_A_298_416#_c_275_n 0.0642298f $X=2.815 $Y=2.575
+ $X2=0 $Y2=0
cc_111 N_A_86_22#_c_91_n N_A_298_416#_c_275_n 0.0182455f $X=2.98 $Y=2.225 $X2=0
+ $Y2=0
cc_112 N_A_86_22#_c_86_n N_A_298_416#_c_269_n 0.0230325f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_113 N_A_86_22#_c_87_n N_A_298_416#_c_269_n 0.0225145f $X=2.505 $Y=0.962 $X2=0
+ $Y2=0
cc_114 N_A_86_22#_c_86_n N_A_298_416#_c_270_n 0.00545495f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_115 N_A_86_22#_c_87_n N_A_298_416#_c_271_n 0.0243142f $X=2.505 $Y=0.962 $X2=0
+ $Y2=0
cc_116 N_A_86_22#_c_101_p N_A_298_416#_c_272_n 0.00366717f $X=2.815 $Y=2.575
+ $X2=0 $Y2=0
cc_117 N_A_86_22#_c_86_n N_A_298_416#_c_272_n 0.0133752f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_118 N_A_86_22#_c_87_n N_A_298_416#_c_272_n 0.00179636f $X=2.505 $Y=0.962
+ $X2=0 $Y2=0
cc_119 N_A_86_22#_c_101_p N_A_298_416#_c_273_n 4.71747e-19 $X=2.815 $Y=2.575
+ $X2=0 $Y2=0
cc_120 N_A_86_22#_c_86_n N_A_298_416#_c_273_n 0.00373219f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_121 N_A_86_22#_c_87_n N_A_298_416#_c_273_n 4.33408e-19 $X=2.505 $Y=0.962
+ $X2=0 $Y2=0
cc_122 N_A_86_22#_c_91_n N_B2_M1008_g 0.0100984f $X=2.98 $Y=2.225 $X2=0 $Y2=0
cc_123 N_A_86_22#_c_121_p N_B2_M1008_g 0.0146553f $X=2.98 $Y=2.575 $X2=0 $Y2=0
cc_124 N_A_86_22#_c_91_n N_B2_c_344_n 9.27233e-19 $X=2.98 $Y=2.225 $X2=0 $Y2=0
cc_125 N_A_86_22#_c_91_n N_B2_c_345_n 0.0114317f $X=2.98 $Y=2.225 $X2=0 $Y2=0
cc_126 N_A_86_22#_c_91_n N_B1_M1002_g 0.00184779f $X=2.98 $Y=2.225 $X2=0 $Y2=0
cc_127 N_A_86_22#_c_121_p N_B1_M1002_g 0.0024654f $X=2.98 $Y=2.575 $X2=0 $Y2=0
cc_128 N_A_86_22#_M1009_g X 0.0141339f $X=0.505 $Y=0.45 $X2=0 $Y2=0
cc_129 N_A_86_22#_c_80_n X 0.00461673f $X=0.555 $Y=1.555 $X2=0 $Y2=0
cc_130 N_A_86_22#_M1005_g X 0.0467474f $X=0.555 $Y=2.58 $X2=0 $Y2=0
cc_131 N_A_86_22#_M1006_g X 0.00202736f $X=0.865 $Y=0.45 $X2=0 $Y2=0
cc_132 N_A_86_22#_c_83_n X 0.00742403f $X=0.555 $Y=1.43 $X2=0 $Y2=0
cc_133 N_A_86_22#_c_146_p X 0.0129587f $X=0.805 $Y=2.575 $X2=0 $Y2=0
cc_134 N_A_86_22#_c_85_n X 0.113027f $X=0.8 $Y=0.945 $X2=0 $Y2=0
cc_135 N_A_86_22#_c_88_n X 0.0121819f $X=0.865 $Y=1.025 $X2=0 $Y2=0
cc_136 N_A_86_22#_c_84_n N_VPWR_M1005_d 0.00559067f $X=0.72 $Y=2.49 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_86_22#_c_101_p N_VPWR_M1005_d 0.016769f $X=2.815 $Y=2.575 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_86_22#_c_146_p N_VPWR_M1005_d 7.33924e-19 $X=0.805 $Y=2.575 $X2=-0.19
+ $Y2=-0.245
cc_139 N_A_86_22#_c_101_p N_VPWR_M1004_d 0.0119464f $X=2.815 $Y=2.575 $X2=0
+ $Y2=0
cc_140 N_A_86_22#_M1005_g N_VPWR_c_434_n 0.0104788f $X=0.555 $Y=2.58 $X2=0 $Y2=0
cc_141 N_A_86_22#_c_101_p N_VPWR_c_434_n 0.0130839f $X=2.815 $Y=2.575 $X2=0
+ $Y2=0
cc_142 N_A_86_22#_c_146_p N_VPWR_c_434_n 0.00723599f $X=0.805 $Y=2.575 $X2=0
+ $Y2=0
cc_143 N_A_86_22#_c_101_p N_VPWR_c_435_n 0.0196988f $X=2.815 $Y=2.575 $X2=0
+ $Y2=0
cc_144 N_A_86_22#_c_121_p N_VPWR_c_435_n 0.00808459f $X=2.98 $Y=2.575 $X2=0
+ $Y2=0
cc_145 N_A_86_22#_c_101_p N_VPWR_c_438_n 0.0150487f $X=2.815 $Y=2.575 $X2=0
+ $Y2=0
cc_146 N_A_86_22#_c_101_p N_VPWR_c_439_n 0.00676762f $X=2.815 $Y=2.575 $X2=0
+ $Y2=0
cc_147 N_A_86_22#_c_121_p N_VPWR_c_439_n 0.0177952f $X=2.98 $Y=2.575 $X2=0 $Y2=0
cc_148 N_A_86_22#_M1005_g N_VPWR_c_440_n 0.00798845f $X=0.555 $Y=2.58 $X2=0
+ $Y2=0
cc_149 N_A_86_22#_c_146_p N_VPWR_c_440_n 3.14802e-19 $X=0.805 $Y=2.575 $X2=0
+ $Y2=0
cc_150 N_A_86_22#_M1005_g N_VPWR_c_433_n 0.0138209f $X=0.555 $Y=2.58 $X2=0 $Y2=0
cc_151 N_A_86_22#_c_101_p N_VPWR_c_433_n 0.0404896f $X=2.815 $Y=2.575 $X2=0
+ $Y2=0
cc_152 N_A_86_22#_c_146_p N_VPWR_c_433_n 0.00123907f $X=0.805 $Y=2.575 $X2=0
+ $Y2=0
cc_153 N_A_86_22#_c_121_p N_VPWR_c_433_n 0.0124497f $X=2.98 $Y=2.575 $X2=0 $Y2=0
cc_154 N_A_86_22#_M1009_g N_VGND_c_485_n 0.00236935f $X=0.505 $Y=0.45 $X2=0
+ $Y2=0
cc_155 N_A_86_22#_M1006_g N_VGND_c_485_n 0.0127614f $X=0.865 $Y=0.45 $X2=0 $Y2=0
cc_156 N_A_86_22#_c_85_n N_VGND_c_485_n 0.00369403f $X=0.8 $Y=0.945 $X2=0 $Y2=0
cc_157 N_A_86_22#_c_87_n N_VGND_c_485_n 0.0218886f $X=2.505 $Y=0.962 $X2=0 $Y2=0
cc_158 N_A_86_22#_M1009_g N_VGND_c_487_n 0.00544432f $X=0.505 $Y=0.45 $X2=0
+ $Y2=0
cc_159 N_A_86_22#_M1006_g N_VGND_c_487_n 0.0048178f $X=0.865 $Y=0.45 $X2=0 $Y2=0
cc_160 N_A_86_22#_M1009_g N_VGND_c_490_n 0.0108302f $X=0.505 $Y=0.45 $X2=0 $Y2=0
cc_161 N_A_86_22#_M1006_g N_VGND_c_490_n 0.00443041f $X=0.865 $Y=0.45 $X2=0
+ $Y2=0
cc_162 N_A_86_22#_c_85_n N_VGND_c_490_n 0.00916864f $X=0.8 $Y=0.945 $X2=0 $Y2=0
cc_163 N_A_86_22#_c_87_n N_VGND_c_490_n 0.0170383f $X=2.505 $Y=0.962 $X2=0 $Y2=0
cc_164 N_A_86_22#_c_86_n N_A_604_142#_c_535_n 0.013592f $X=2.67 $Y=0.96 $X2=0
+ $Y2=0
cc_165 N_A1_N_M1010_g N_A2_N_c_222_n 0.0414328f $X=1.295 $Y=0.45 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A1_N_M1007_g N_A2_N_M1004_g 0.044864f $X=1.365 $Y=2.58 $X2=0 $Y2=0
cc_167 A1_N N_A2_N_M1004_g 8.67877e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A1_N_M1010_g N_A2_N_c_224_n 0.0217587f $X=1.295 $Y=0.45 $X2=0 $Y2=0
cc_169 A1_N N_A2_N_c_225_n 2.52415e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A1_N_c_180_n N_A2_N_c_225_n 0.0176933f $X=1.365 $Y=1.715 $X2=0 $Y2=0
cc_171 N_A1_N_M1010_g A2_N 0.00930274f $X=1.295 $Y=0.45 $X2=0 $Y2=0
cc_172 A1_N A2_N 0.0208734f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_173 N_A1_N_c_180_n A2_N 0.00325314f $X=1.365 $Y=1.715 $X2=0 $Y2=0
cc_174 A1_N N_A_298_416#_c_275_n 0.00400986f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A1_N_M1010_g N_A_298_416#_c_271_n 0.00116561f $X=1.295 $Y=0.45 $X2=0
+ $Y2=0
cc_176 A1_N N_VPWR_M1005_d 0.003952f $X=1.115 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_177 N_A1_N_M1007_g N_VPWR_c_434_n 0.0080455f $X=1.365 $Y=2.58 $X2=0 $Y2=0
cc_178 N_A1_N_M1007_g N_VPWR_c_435_n 0.00182395f $X=1.365 $Y=2.58 $X2=0 $Y2=0
cc_179 N_A1_N_M1007_g N_VPWR_c_438_n 0.00695957f $X=1.365 $Y=2.58 $X2=0 $Y2=0
cc_180 N_A1_N_M1007_g N_VPWR_c_433_n 0.00953065f $X=1.365 $Y=2.58 $X2=0 $Y2=0
cc_181 N_A1_N_M1010_g N_VGND_c_485_n 0.0130241f $X=1.295 $Y=0.45 $X2=0 $Y2=0
cc_182 N_A1_N_M1010_g N_VGND_c_488_n 0.0048178f $X=1.295 $Y=0.45 $X2=0 $Y2=0
cc_183 N_A1_N_M1010_g N_VGND_c_490_n 0.00455744f $X=1.295 $Y=0.45 $X2=0 $Y2=0
cc_184 N_A2_N_c_223_n N_A_298_416#_c_267_n 0.0143365f $X=1.805 $Y=0.81 $X2=0
+ $Y2=0
cc_185 A2_N N_A_298_416#_c_267_n 0.0126029f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_186 N_A2_N_c_227_n N_A_298_416#_c_267_n 0.0162204f $X=1.895 $Y=1.375 $X2=0
+ $Y2=0
cc_187 N_A2_N_M1004_g N_A_298_416#_M1000_g 0.0237215f $X=1.925 $Y=2.58 $X2=0
+ $Y2=0
cc_188 N_A2_N_c_230_n N_A_298_416#_M1000_g 8.687e-19 $X=1.895 $Y=1.88 $X2=0
+ $Y2=0
cc_189 N_A2_N_M1004_g N_A_298_416#_c_275_n 0.0177538f $X=1.925 $Y=2.58 $X2=0
+ $Y2=0
cc_190 N_A2_N_c_230_n N_A_298_416#_c_275_n 0.00210689f $X=1.895 $Y=1.88 $X2=0
+ $Y2=0
cc_191 A2_N N_A_298_416#_c_275_n 0.0563158f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_192 N_A2_N_c_222_n N_A_298_416#_c_270_n 0.0037342f $X=1.685 $Y=0.735 $X2=0
+ $Y2=0
cc_193 N_A2_N_M1004_g N_A_298_416#_c_276_n 0.00319443f $X=1.925 $Y=2.58 $X2=0
+ $Y2=0
cc_194 N_A2_N_c_222_n N_A_298_416#_c_271_n 0.00795073f $X=1.685 $Y=0.735 $X2=0
+ $Y2=0
cc_195 N_A2_N_c_223_n N_A_298_416#_c_271_n 0.00371883f $X=1.805 $Y=0.81 $X2=0
+ $Y2=0
cc_196 N_A2_N_c_225_n N_A_298_416#_c_272_n 2.31274e-19 $X=1.895 $Y=1.715 $X2=0
+ $Y2=0
cc_197 A2_N N_A_298_416#_c_272_n 0.0307f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A2_N_c_225_n N_A_298_416#_c_273_n 0.0162204f $X=1.895 $Y=1.715 $X2=0
+ $Y2=0
cc_199 N_A2_N_M1004_g N_VPWR_c_435_n 0.0106975f $X=1.925 $Y=2.58 $X2=0 $Y2=0
cc_200 N_A2_N_M1004_g N_VPWR_c_438_n 0.00625647f $X=1.925 $Y=2.58 $X2=0 $Y2=0
cc_201 N_A2_N_M1004_g N_VPWR_c_433_n 0.00722795f $X=1.925 $Y=2.58 $X2=0 $Y2=0
cc_202 N_A2_N_c_222_n N_VGND_c_485_n 0.00237422f $X=1.685 $Y=0.735 $X2=0 $Y2=0
cc_203 N_A2_N_c_222_n N_VGND_c_488_n 0.00542974f $X=1.685 $Y=0.735 $X2=0 $Y2=0
cc_204 N_A2_N_c_222_n N_VGND_c_490_n 0.00760646f $X=1.685 $Y=0.735 $X2=0 $Y2=0
cc_205 N_A_298_416#_M1000_g N_B2_M1008_g 0.0294952f $X=2.715 $Y=2.58 $X2=0 $Y2=0
cc_206 N_A_298_416#_c_276_n N_B2_M1008_g 7.90473e-19 $X=2.54 $Y=2.06 $X2=0 $Y2=0
cc_207 N_A_298_416#_c_270_n N_B2_c_342_n 0.00922856f $X=2.67 $Y=0.43 $X2=0 $Y2=0
cc_208 N_A_298_416#_c_268_n N_B2_c_343_n 0.00300598f $X=2.945 $Y=0.595 $X2=0
+ $Y2=0
cc_209 N_A_298_416#_c_272_n N_B2_c_344_n 2.85737e-19 $X=2.62 $Y=1.665 $X2=0
+ $Y2=0
cc_210 N_A_298_416#_c_273_n N_B2_c_344_n 0.0178647f $X=2.715 $Y=1.665 $X2=0
+ $Y2=0
cc_211 N_A_298_416#_c_268_n N_B2_c_345_n 4.17882e-19 $X=2.945 $Y=0.595 $X2=0
+ $Y2=0
cc_212 N_A_298_416#_c_276_n N_B2_c_345_n 0.00205953f $X=2.54 $Y=2.06 $X2=0 $Y2=0
cc_213 N_A_298_416#_c_272_n N_B2_c_345_n 0.0185845f $X=2.62 $Y=1.665 $X2=0 $Y2=0
cc_214 N_A_298_416#_c_273_n N_B2_c_345_n 0.00248433f $X=2.715 $Y=1.665 $X2=0
+ $Y2=0
cc_215 N_A_298_416#_c_272_n N_B2_c_346_n 2.54124e-19 $X=2.62 $Y=1.665 $X2=0
+ $Y2=0
cc_216 N_A_298_416#_c_273_n N_B2_c_346_n 0.00165604f $X=2.715 $Y=1.665 $X2=0
+ $Y2=0
cc_217 N_A_298_416#_c_275_n N_VPWR_M1004_d 0.00700057f $X=2.455 $Y=2.185 $X2=0
+ $Y2=0
cc_218 N_A_298_416#_M1000_g N_VPWR_c_435_n 0.00520855f $X=2.715 $Y=2.58 $X2=0
+ $Y2=0
cc_219 N_A_298_416#_M1000_g N_VPWR_c_439_n 0.00686123f $X=2.715 $Y=2.58 $X2=0
+ $Y2=0
cc_220 N_A_298_416#_M1000_g N_VPWR_c_433_n 0.00930969f $X=2.715 $Y=2.58 $X2=0
+ $Y2=0
cc_221 N_A_298_416#_c_271_n N_VGND_c_485_n 0.0137212f $X=2.065 $Y=0.472 $X2=0
+ $Y2=0
cc_222 N_A_298_416#_c_269_n N_VGND_c_486_n 0.010097f $X=2.67 $Y=0.43 $X2=0 $Y2=0
cc_223 N_A_298_416#_c_270_n N_VGND_c_486_n 0.00755746f $X=2.67 $Y=0.43 $X2=0
+ $Y2=0
cc_224 N_A_298_416#_c_270_n N_VGND_c_488_n 0.0152335f $X=2.67 $Y=0.43 $X2=0
+ $Y2=0
cc_225 N_A_298_416#_c_271_n N_VGND_c_488_n 0.0670212f $X=2.065 $Y=0.472 $X2=0
+ $Y2=0
cc_226 N_A_298_416#_M1011_d N_VGND_c_490_n 0.00231257f $X=1.76 $Y=0.24 $X2=0
+ $Y2=0
cc_227 N_A_298_416#_c_270_n N_VGND_c_490_n 0.0174904f $X=2.67 $Y=0.43 $X2=0
+ $Y2=0
cc_228 N_A_298_416#_c_271_n N_VGND_c_490_n 0.0414983f $X=2.065 $Y=0.472 $X2=0
+ $Y2=0
cc_229 N_A_298_416#_c_267_n N_A_604_142#_c_535_n 7.58573e-19 $X=2.375 $Y=1.5
+ $X2=0 $Y2=0
cc_230 N_A_298_416#_c_268_n N_A_604_142#_c_535_n 0.00709118f $X=2.945 $Y=0.595
+ $X2=0 $Y2=0
cc_231 N_A_298_416#_c_267_n N_A_604_142#_c_537_n 0.00325921f $X=2.375 $Y=1.5
+ $X2=0 $Y2=0
cc_232 N_A_298_416#_c_268_n N_A_604_142#_c_537_n 0.00194636f $X=2.945 $Y=0.595
+ $X2=0 $Y2=0
cc_233 N_B2_M1008_g N_B1_M1002_g 0.0631084f $X=3.245 $Y=2.58 $X2=0 $Y2=0
cc_234 N_B2_c_342_n N_B1_M1003_g 0.0183466f $X=3.365 $Y=1.205 $X2=0 $Y2=0
cc_235 N_B2_c_346_n N_B1_M1003_g 0.00814396f $X=3.245 $Y=1.55 $X2=0 $Y2=0
cc_236 N_B2_c_344_n B1 4.17281e-19 $X=3.245 $Y=1.715 $X2=0 $Y2=0
cc_237 N_B2_c_345_n B1 0.0199435f $X=3.245 $Y=1.715 $X2=0 $Y2=0
cc_238 N_B2_c_344_n N_B1_c_391_n 0.0181729f $X=3.245 $Y=1.715 $X2=0 $Y2=0
cc_239 N_B2_c_345_n N_B1_c_391_n 4.19061e-19 $X=3.245 $Y=1.715 $X2=0 $Y2=0
cc_240 N_B2_M1008_g N_VPWR_c_437_n 0.00521606f $X=3.245 $Y=2.58 $X2=0 $Y2=0
cc_241 N_B2_M1008_g N_VPWR_c_439_n 0.00914935f $X=3.245 $Y=2.58 $X2=0 $Y2=0
cc_242 N_B2_M1008_g N_VPWR_c_433_n 0.0161749f $X=3.245 $Y=2.58 $X2=0 $Y2=0
cc_243 N_B2_c_342_n N_VGND_c_486_n 0.00750773f $X=3.365 $Y=1.205 $X2=0 $Y2=0
cc_244 N_B2_c_342_n N_VGND_c_488_n 0.00310242f $X=3.365 $Y=1.205 $X2=0 $Y2=0
cc_245 N_B2_c_342_n N_VGND_c_490_n 0.00375113f $X=3.365 $Y=1.205 $X2=0 $Y2=0
cc_246 N_B2_c_342_n N_A_604_142#_c_535_n 0.0012088f $X=3.365 $Y=1.205 $X2=0
+ $Y2=0
cc_247 N_B2_c_342_n N_A_604_142#_c_536_n 0.00574613f $X=3.365 $Y=1.205 $X2=0
+ $Y2=0
cc_248 N_B2_c_343_n N_A_604_142#_c_536_n 0.00623324f $X=3.365 $Y=1.355 $X2=0
+ $Y2=0
cc_249 N_B2_c_345_n N_A_604_142#_c_536_n 0.00985854f $X=3.245 $Y=1.715 $X2=0
+ $Y2=0
cc_250 N_B2_c_346_n N_A_604_142#_c_536_n 0.00238339f $X=3.245 $Y=1.55 $X2=0
+ $Y2=0
cc_251 N_B2_c_343_n N_A_604_142#_c_537_n 0.00258469f $X=3.365 $Y=1.355 $X2=0
+ $Y2=0
cc_252 N_B2_c_344_n N_A_604_142#_c_537_n 0.00471146f $X=3.245 $Y=1.715 $X2=0
+ $Y2=0
cc_253 N_B2_c_345_n N_A_604_142#_c_537_n 0.0204432f $X=3.245 $Y=1.715 $X2=0
+ $Y2=0
cc_254 N_B2_c_346_n N_A_604_142#_c_537_n 2.6903e-19 $X=3.245 $Y=1.55 $X2=0 $Y2=0
cc_255 N_B2_c_342_n N_A_604_142#_c_538_n 4.81543e-19 $X=3.365 $Y=1.205 $X2=0
+ $Y2=0
cc_256 N_B1_M1002_g N_VPWR_c_437_n 0.0274481f $X=3.775 $Y=2.58 $X2=0 $Y2=0
cc_257 B1 N_VPWR_c_437_n 0.0273201f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_258 N_B1_c_391_n N_VPWR_c_437_n 0.00185447f $X=3.815 $Y=1.715 $X2=0 $Y2=0
cc_259 N_B1_M1002_g N_VPWR_c_439_n 0.00853443f $X=3.775 $Y=2.58 $X2=0 $Y2=0
cc_260 N_B1_M1002_g N_VPWR_c_433_n 0.0144982f $X=3.775 $Y=2.58 $X2=0 $Y2=0
cc_261 N_B1_M1003_g N_VGND_c_486_n 0.00331843f $X=3.825 $Y=0.92 $X2=0 $Y2=0
cc_262 N_B1_M1003_g N_VGND_c_489_n 0.00373213f $X=3.825 $Y=0.92 $X2=0 $Y2=0
cc_263 N_B1_M1003_g N_VGND_c_490_n 0.00446563f $X=3.825 $Y=0.92 $X2=0 $Y2=0
cc_264 N_B1_M1003_g N_A_604_142#_c_536_n 0.0151674f $X=3.825 $Y=0.92 $X2=0 $Y2=0
cc_265 B1 N_A_604_142#_c_536_n 0.0425975f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_266 N_B1_c_391_n N_A_604_142#_c_536_n 0.00445386f $X=3.815 $Y=1.715 $X2=0
+ $Y2=0
cc_267 N_B1_M1003_g N_A_604_142#_c_538_n 0.00705273f $X=3.825 $Y=0.92 $X2=0
+ $Y2=0
cc_268 X N_VPWR_c_434_n 0.0148254f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_269 X N_VPWR_c_440_n 0.019758f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_270 X N_VPWR_c_433_n 0.0125705f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_271 X N_VGND_c_485_n 0.0138848f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_272 X N_VGND_c_487_n 0.0197885f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_273 N_X_M1009_s N_VGND_c_490_n 0.0023122f $X=0.145 $Y=0.24 $X2=0 $Y2=0
cc_274 X N_VGND_c_490_n 0.0125808f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_275 A_116_48# N_VGND_c_490_n 0.00470202f $X=0.58 $Y=0.24 $X2=4.08 $Y2=0
cc_276 N_VGND_c_490_n A_274_48# 0.00359358f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_277 N_VGND_c_486_n N_A_604_142#_c_535_n 0.0120629f $X=3.61 $Y=0.855 $X2=0
+ $Y2=0
cc_278 N_VGND_c_488_n N_A_604_142#_c_535_n 0.00449032f $X=3.445 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_490_n N_A_604_142#_c_535_n 0.007221f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_c_486_n N_A_604_142#_c_536_n 0.0169767f $X=3.61 $Y=0.855 $X2=0
+ $Y2=0
cc_281 N_VGND_c_490_n N_A_604_142#_c_538_n 0.0123586f $X=4.08 $Y=0 $X2=0 $Y2=0
