* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__lsbuf_lp A DESTPWR DESTVPB VGND VPB VPWR X
X0 VPWR A a_206_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X1 DESTPWR a_193_718# a_434_1085# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X2 a_206_446# A a_278_47# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_276_718# A VGND VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_434_1085# a_193_718# a_246_987# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X5 a_206_47# A a_278_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X6 a_276_1085# a_246_987# DESTPWR DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X7 VGND A a_206_446# VGND sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_193_718# a_246_987# a_276_1085# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X9 a_193_718# A a_276_718# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_712_718# a_193_718# X VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND a_278_47# a_434_718# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_712_1085# a_193_718# X DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 DESTPWR a_193_718# a_712_1085# DESTVPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X14 VGND a_193_718# a_712_718# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_434_718# a_278_47# a_246_987# VGND sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
