* File: sky130_fd_sc_lp__nand2_lp2.pxi.spice
* Created: Wed Sep  2 10:03:04 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2_LP2%B N_B_M1003_g N_B_M1001_g B B N_B_c_34_n
+ N_B_c_35_n PM_SKY130_FD_SC_LP__NAND2_LP2%B
x_PM_SKY130_FD_SC_LP__NAND2_LP2%A N_A_M1000_g N_A_c_63_n N_A_M1002_g N_A_c_65_n
+ A N_A_c_66_n N_A_c_67_n PM_SKY130_FD_SC_LP__NAND2_LP2%A
x_PM_SKY130_FD_SC_LP__NAND2_LP2%VPWR N_VPWR_M1003_s N_VPWR_M1002_d N_VPWR_c_99_n
+ N_VPWR_c_100_n N_VPWR_c_101_n N_VPWR_c_102_n N_VPWR_c_103_n VPWR
+ N_VPWR_c_104_n N_VPWR_c_98_n PM_SKY130_FD_SC_LP__NAND2_LP2%VPWR
x_PM_SKY130_FD_SC_LP__NAND2_LP2%Y N_Y_M1000_d N_Y_M1003_d N_Y_c_123_n
+ N_Y_c_124_n N_Y_c_125_n N_Y_c_121_n Y Y PM_SKY130_FD_SC_LP__NAND2_LP2%Y
x_PM_SKY130_FD_SC_LP__NAND2_LP2%VGND N_VGND_M1001_s N_VGND_c_154_n
+ N_VGND_c_155_n N_VGND_c_156_n VGND N_VGND_c_157_n N_VGND_c_158_n
+ PM_SKY130_FD_SC_LP__NAND2_LP2%VGND
cc_1 VNB N_B_M1001_g 0.0446218f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.495
cc_2 VNB N_B_c_34_n 0.0677065f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_3 VNB N_B_c_35_n 0.031314f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_4 VNB N_A_M1000_g 0.0223227f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.545
cc_5 VNB N_A_c_63_n 0.0153207f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.11
cc_6 VNB N_A_M1002_g 0.00969693f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.495
cc_7 VNB N_A_c_65_n 0.026828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_c_66_n 0.0182104f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.275
cc_9 VNB N_A_c_67_n 0.00237362f $X=-0.19 $Y=-0.245 $X2=0.487 $Y2=1.11
cc_10 VNB N_VPWR_c_98_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_Y_c_121_n 0.0488869f $X=-0.19 $Y=-0.245 $X2=0.487 $Y2=1.11
cc_12 VNB Y 0.0319887f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.275
cc_13 VNB N_VGND_c_154_n 0.0251828f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.495
cc_14 VNB N_VGND_c_155_n 0.0116899f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_VGND_c_156_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_VGND_c_157_n 0.0368502f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_17 VNB N_VGND_c_158_n 0.152443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VPB N_B_M1003_g 0.0405011f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.545
cc_19 VPB N_B_c_34_n 0.0207617f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_20 VPB N_B_c_35_n 0.011116f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_21 VPB N_A_M1002_g 0.0478789f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.495
cc_22 VPB N_VPWR_c_99_n 0.0140682f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.495
cc_23 VPB N_VPWR_c_100_n 0.0463954f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_24 VPB N_VPWR_c_101_n 0.0433017f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_25 VPB N_VPWR_c_102_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.295
cc_26 VPB N_VPWR_c_103_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_104_n 0.0126445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_98_n 0.0593457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_Y_c_123_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_30 VPB N_Y_c_124_n 0.0304119f $X=-0.19 $Y=1.655 $X2=0.487 $Y2=1.275
cc_31 VPB N_Y_c_125_n 0.0100597f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.275
cc_32 VPB N_Y_c_121_n 0.00227167f $X=-0.19 $Y=1.655 $X2=0.487 $Y2=1.11
cc_33 N_B_M1001_g N_A_M1000_g 0.0367696f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_34 N_B_c_34_n N_A_M1002_g 0.0316273f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_35 N_B_c_35_n N_A_M1002_g 8.45303e-19 $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_36 N_B_c_34_n N_A_c_65_n 0.0367696f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_37 N_B_c_35_n N_A_c_65_n 0.00110392f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_38 N_B_M1001_g N_A_c_67_n 0.0035211f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_39 N_B_c_35_n N_A_c_67_n 0.0143724f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_40 N_B_M1003_g N_VPWR_c_100_n 0.0237672f $X=0.63 $Y=2.545 $X2=0 $Y2=0
cc_41 N_B_c_34_n N_VPWR_c_100_n 0.00213795f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_42 N_B_c_35_n N_VPWR_c_100_n 0.0221614f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_43 N_B_M1003_g N_VPWR_c_101_n 9.32056e-19 $X=0.63 $Y=2.545 $X2=0 $Y2=0
cc_44 N_B_M1003_g N_VPWR_c_102_n 0.00769046f $X=0.63 $Y=2.545 $X2=0 $Y2=0
cc_45 N_B_M1003_g N_VPWR_c_98_n 0.0134474f $X=0.63 $Y=2.545 $X2=0 $Y2=0
cc_46 N_B_M1003_g N_Y_c_123_n 0.0275305f $X=0.63 $Y=2.545 $X2=0 $Y2=0
cc_47 N_B_M1003_g N_Y_c_125_n 0.00535934f $X=0.63 $Y=2.545 $X2=0 $Y2=0
cc_48 N_B_c_34_n N_Y_c_125_n 0.00363299f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_49 N_B_c_35_n N_Y_c_125_n 0.00621187f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_50 N_B_M1001_g Y 0.00121001f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_51 N_B_M1001_g N_VGND_c_154_n 0.0150742f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_52 N_B_c_34_n N_VGND_c_154_n 0.00390484f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_53 N_B_c_35_n N_VGND_c_154_n 0.0119653f $X=0.385 $Y=1.275 $X2=0 $Y2=0
cc_54 N_B_M1001_g N_VGND_c_157_n 0.00445056f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_55 N_B_M1001_g N_VGND_c_158_n 0.00804604f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_56 N_A_M1002_g N_VPWR_c_100_n 9.45383e-19 $X=1.16 $Y=2.545 $X2=0 $Y2=0
cc_57 N_A_M1002_g N_VPWR_c_101_n 0.0228842f $X=1.16 $Y=2.545 $X2=0 $Y2=0
cc_58 N_A_M1002_g N_VPWR_c_102_n 0.00769046f $X=1.16 $Y=2.545 $X2=0 $Y2=0
cc_59 N_A_M1002_g N_VPWR_c_98_n 0.0134474f $X=1.16 $Y=2.545 $X2=0 $Y2=0
cc_60 N_A_M1002_g N_Y_c_123_n 0.0282068f $X=1.16 $Y=2.545 $X2=0 $Y2=0
cc_61 N_A_c_63_n N_Y_c_124_n 2.68303e-19 $X=1.16 $Y=1.52 $X2=0 $Y2=0
cc_62 N_A_M1002_g N_Y_c_124_n 0.0196736f $X=1.16 $Y=2.545 $X2=0 $Y2=0
cc_63 N_A_c_67_n N_Y_c_124_n 0.0192947f $X=1.16 $Y=1.015 $X2=0 $Y2=0
cc_64 N_A_c_63_n N_Y_c_125_n 3.02817e-19 $X=1.16 $Y=1.52 $X2=0 $Y2=0
cc_65 N_A_M1002_g N_Y_c_125_n 0.00277178f $X=1.16 $Y=2.545 $X2=0 $Y2=0
cc_66 N_A_c_67_n N_Y_c_125_n 0.00534367f $X=1.16 $Y=1.015 $X2=0 $Y2=0
cc_67 N_A_M1000_g N_Y_c_121_n 0.00442487f $X=1.07 $Y=0.495 $X2=0 $Y2=0
cc_68 N_A_M1002_g N_Y_c_121_n 0.00542577f $X=1.16 $Y=2.545 $X2=0 $Y2=0
cc_69 N_A_c_66_n N_Y_c_121_n 0.0136805f $X=1.16 $Y=1.015 $X2=0 $Y2=0
cc_70 N_A_c_67_n N_Y_c_121_n 0.0329161f $X=1.16 $Y=1.015 $X2=0 $Y2=0
cc_71 N_A_M1000_g Y 0.00940558f $X=1.07 $Y=0.495 $X2=0 $Y2=0
cc_72 N_A_c_66_n Y 0.00116454f $X=1.16 $Y=1.015 $X2=0 $Y2=0
cc_73 N_A_c_67_n Y 0.0162244f $X=1.16 $Y=1.015 $X2=0 $Y2=0
cc_74 N_A_M1000_g N_VGND_c_154_n 0.00222856f $X=1.07 $Y=0.495 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_VGND_c_157_n 0.00452629f $X=1.07 $Y=0.495 $X2=0 $Y2=0
cc_76 N_A_M1000_g N_VGND_c_158_n 0.00638091f $X=1.07 $Y=0.495 $X2=0 $Y2=0
cc_77 N_A_c_67_n N_VGND_c_158_n 0.00315634f $X=1.16 $Y=1.015 $X2=0 $Y2=0
cc_78 N_VPWR_c_100_n N_Y_c_123_n 0.0685263f $X=0.365 $Y=2.19 $X2=0 $Y2=0
cc_79 N_VPWR_c_101_n N_Y_c_123_n 0.066879f $X=1.425 $Y=2.215 $X2=0 $Y2=0
cc_80 N_VPWR_c_102_n N_Y_c_123_n 0.021949f $X=1.26 $Y=3.33 $X2=0 $Y2=0
cc_81 N_VPWR_c_98_n N_Y_c_123_n 0.0124703f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_82 N_VPWR_c_101_n N_Y_c_124_n 0.0233986f $X=1.425 $Y=2.215 $X2=0 $Y2=0
cc_83 Y N_VGND_c_154_n 0.0142378f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_84 Y N_VGND_c_157_n 0.0343546f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_85 Y N_VGND_c_158_n 0.0254496f $X=1.595 $Y=0.47 $X2=0 $Y2=0
