* File: sky130_fd_sc_lp__nand4bb_4.spice
* Created: Wed Sep  2 10:06:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4bb_4.pex.spice"
.subckt sky130_fd_sc_lp__nand4bb_4  VNB VPB A_N B_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1032 N_VGND_M1032_d N_A_N_M1032_g N_A_44_69#_M1032_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=2.856 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1004 N_A_217_69#_M1004_d N_B_N_M1004_g N_VGND_M1032_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1015 N_Y_M1015_d N_A_44_69#_M1015_g N_A_324_45#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.3679 PD=1.12 PS=2.7 NRD=0 NRS=17.136 M=1 R=5.6
+ SA=75000.3 SB=75003.5 A=0.126 P=1.98 MULT=1
MM1016 N_Y_M1015_d N_A_44_69#_M1016_g N_A_324_45#_M1016_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75000.8 SB=75003.1 A=0.126 P=1.98 MULT=1
MM1028 N_Y_M1028_d N_A_44_69#_M1028_g N_A_324_45#_M1016_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75001.3 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1029 N_Y_M1028_d N_A_44_69#_M1029_g N_A_324_45#_M1029_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75001.8 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1000 N_A_324_45#_M1029_s N_A_217_69#_M1000_g N_A_842_67#_M1000_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.20075 AS=0.1176 PD=1.39 PS=1.12 NRD=12.132 NRS=0 M=1 R=5.6
+ SA=75002.4 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1012 N_A_324_45#_M1012_d N_A_217_69#_M1012_g N_A_842_67#_M1000_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75002.8 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1022 N_A_324_45#_M1012_d N_A_217_69#_M1022_g N_A_842_67#_M1022_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75003.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1030 N_A_324_45#_M1030_d N_A_217_69#_M1030_g N_A_842_67#_M1022_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75003.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_842_67#_M1001_d N_C_M1001_g N_A_1251_47#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1013 N_A_842_67#_M1001_d N_C_M1013_g N_A_1251_47#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1017 N_A_842_67#_M1017_d N_C_M1017_g N_A_1251_47#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1019 N_A_842_67#_M1017_d N_C_M1019_g N_A_1251_47#_M1019_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1008 N_A_1251_47#_M1019_s N_D_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1010 N_A_1251_47#_M1010_d N_D_M1010_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1024 N_A_1251_47#_M1010_d N_D_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1034 N_A_1251_47#_M1034_d N_D_M1034_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_N_M1002_g N_A_44_69#_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1011 N_A_217_69#_M1011_d N_B_N_M1011_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A_44_69#_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75007.5 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A_44_69#_M1014_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75007.1 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1014_d N_A_44_69#_M1025_g N_Y_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75006.7 A=0.189 P=2.82 MULT=1
MM1035 N_VPWR_M1035_d N_A_44_69#_M1035_g N_Y_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75006.2 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_217_69#_M1005_g N_VPWR_M1035_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75005.8 A=0.189 P=2.82 MULT=1
MM1018 N_Y_M1005_d N_A_217_69#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75005.4 A=0.189 P=2.82 MULT=1
MM1023 N_Y_M1023_d N_A_217_69#_M1023_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8 SB=75005
+ A=0.189 P=2.82 MULT=1
MM1031 N_Y_M1023_d N_A_217_69#_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.7434 PD=1.54 PS=2.44 NRD=0 NRS=70.3487 M=1 R=8.4 SA=75003.2
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1031_s N_C_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.7434 AS=0.1764 PD=2.44 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_C_M1009_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005 SB=75002.8
+ A=0.189 P=2.82 MULT=1
MM1020 N_VPWR_M1009_d N_C_M1020_g N_Y_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.4
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1033 N_VPWR_M1033_d N_C_M1033_g N_Y_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.8
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_D_M1003_g N_VPWR_M1033_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1021 N_Y_M1003_d N_D_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.7
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1026 N_Y_M1026_d N_D_M1026_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_Y_M1026_d N_D_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75007.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX36_noxref VNB VPB NWDIODE A=19.5079 P=24.65
*
.include "sky130_fd_sc_lp__nand4bb_4.pxi.spice"
*
.ends
*
*
