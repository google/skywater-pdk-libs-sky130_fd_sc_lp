* File: sky130_fd_sc_lp__sdfstp_2.pex.spice
* Created: Wed Sep  2 10:35:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%SCD 3 5 7 11 14 15 16 20
r33 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.3 $X2=0.385 $Y2=1.3
r34 16 21 9.38857 $w=4.63e-07 $l=3.65e-07 $layer=LI1_cond $X=0.317 $Y=1.665
+ $X2=0.317 $Y2=1.3
r35 15 21 0.128611 $w=4.63e-07 $l=5e-09 $layer=LI1_cond $X=0.317 $Y=1.295
+ $X2=0.317 $Y2=1.3
r36 13 20 44.2071 $w=3.9e-07 $l=3.1e-07 $layer=POLY_cond $X=0.415 $Y=1.61
+ $X2=0.415 $Y2=1.3
r37 13 14 49.7341 $w=3.9e-07 $l=1.95e-07 $layer=POLY_cond $X=0.415 $Y=1.61
+ $X2=0.415 $Y2=1.805
r38 9 20 2.13905 $w=3.9e-07 $l=1.5e-08 $layer=POLY_cond $X=0.415 $Y=1.285
+ $X2=0.415 $Y2=1.3
r39 9 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.415 $Y=1.21
+ $X2=0.785 $Y2=1.21
r40 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.785 $Y=1.135
+ $X2=0.785 $Y2=1.21
r41 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.785 $Y=1.135
+ $X2=0.785 $Y2=0.815
r42 3 14 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=0.535 $Y=2.725
+ $X2=0.535 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%D 1 3 7 9 10 11 12 13
r42 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.415
+ $Y=2.08 $X2=1.415 $Y2=2.08
r43 12 13 20.1154 $w=2.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.087
+ $X2=2.16 $Y2=2.087
r44 12 21 11.1054 $w=2.73e-07 $l=2.65e-07 $layer=LI1_cond $X=1.68 $Y=2.087
+ $X2=1.415 $Y2=2.087
r45 11 21 9.01001 $w=2.73e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=2.087
+ $X2=1.415 $Y2=2.087
r46 10 11 20.1154 $w=2.73e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=2.087
+ $X2=1.2 $Y2=2.087
r47 9 10 20.1154 $w=2.73e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=2.087
+ $X2=0.72 $Y2=2.087
r48 5 20 65.0101 $w=2.92e-07 $l=3.82426e-07 $layer=POLY_cond $X=1.575 $Y=1.755
+ $X2=1.45 $Y2=2.08
r49 5 7 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.575 $Y=1.755 $X2=1.575
+ $Y2=0.815
r50 1 20 38.5991 $w=2.92e-07 $l=2.18746e-07 $layer=POLY_cond $X=1.325 $Y=2.245
+ $X2=1.45 $Y2=2.08
r51 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.325 $Y=2.245
+ $X2=1.325 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_358_429# 1 2 9 12 16 18 19 20 23 25 26 32
+ 34
r73 30 32 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=3.66 $Y=1.78
+ $X2=3.66 $Y2=2.465
r74 29 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.125 $Y=1.645
+ $X2=3.125 $Y2=1.555
r75 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.125
+ $Y=1.645 $X2=3.125 $Y2=1.645
r76 26 28 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=3.085 $Y=1.665
+ $X2=3.125 $Y2=1.665
r77 25 30 6.8319 $w=2.3e-07 $l=1.73205e-07 $layer=LI1_cond $X=3.535 $Y=1.665
+ $X2=3.66 $Y2=1.78
r78 25 28 20.5435 $w=2.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.535 $Y=1.665
+ $X2=3.125 $Y2=1.665
r79 21 26 6.95328 $w=2.3e-07 $l=1.97292e-07 $layer=LI1_cond $X=2.937 $Y=1.55
+ $X2=3.085 $Y2=1.665
r80 21 23 28.7134 $w=2.93e-07 $l=7.35e-07 $layer=LI1_cond $X=2.937 $Y=1.55
+ $X2=2.937 $Y2=0.815
r81 18 19 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.9 $Y=2.145 $X2=1.9
+ $Y2=2.295
r82 17 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.01 $Y=1.555
+ $X2=1.935 $Y2=1.555
r83 16 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.96 $Y=1.555
+ $X2=3.125 $Y2=1.555
r84 16 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.96 $Y=1.555
+ $X2=2.01 $Y2=1.555
r85 14 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.935 $Y=1.63
+ $X2=1.935 $Y2=1.555
r86 14 18 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.935 $Y=1.63
+ $X2=1.935 $Y2=2.145
r87 10 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.935 $Y=1.48
+ $X2=1.935 $Y2=1.555
r88 10 12 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=1.935 $Y=1.48
+ $X2=1.935 $Y2=0.815
r89 9 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.865 $Y=2.725
+ $X2=1.865 $Y2=2.295
r90 2 32 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=2.31 $X2=3.62 $Y2=2.465
r91 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.78
+ $Y=0.605 $X2=2.92 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%SCE 3 8 9 10 13 15 17 19 21 24 26 29 33 34
+ 35 36 41 42
c85 13 0 6.49935e-20 $X=2.705 $Y=0.815
r86 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.6 $Y=0.43
+ $X2=3.6 $Y2=0.43
r87 35 36 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=0.925 $X2=3.6
+ $Y2=1.295
r88 34 35 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=0.555 $X2=3.6
+ $Y2=0.925
r89 34 42 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.6 $Y=0.555
+ $X2=3.6 $Y2=0.43
r90 32 41 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.6 $Y=0.77 $X2=3.6
+ $Y2=0.43
r91 32 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=0.77 $X2=3.6
+ $Y2=0.935
r92 31 41 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=0.265
+ $X2=3.6 $Y2=0.43
r93 27 29 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.405 $Y=2.125
+ $X2=3.69 $Y2=2.125
r94 22 24 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.965 $Y=1.6
+ $X2=1.145 $Y2=1.6
r95 21 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.69 $Y=2.05
+ $X2=3.69 $Y2=2.125
r96 21 33 571.734 $w=1.5e-07 $l=1.115e-06 $layer=POLY_cond $X=3.69 $Y=2.05
+ $X2=3.69 $Y2=0.935
r97 17 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.405 $Y=2.2
+ $X2=3.405 $Y2=2.125
r98 17 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.405 $Y=2.2
+ $X2=3.405 $Y2=2.63
r99 16 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.78 $Y=0.19
+ $X2=2.705 $Y2=0.19
r100 15 31 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.435 $Y=0.19
+ $X2=3.6 $Y2=0.265
r101 15 16 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=3.435 $Y=0.19
+ $X2=2.78 $Y2=0.19
r102 11 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.705 $Y=0.265
+ $X2=2.705 $Y2=0.19
r103 11 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.705 $Y=0.265
+ $X2=2.705 $Y2=0.815
r104 9 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.63 $Y=0.19
+ $X2=2.705 $Y2=0.19
r105 9 10 723 $w=1.5e-07 $l=1.41e-06 $layer=POLY_cond $X=2.63 $Y=0.19 $X2=1.22
+ $Y2=0.19
r106 6 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.145 $Y=1.525
+ $X2=1.145 $Y2=1.6
r107 6 8 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.145 $Y=1.525
+ $X2=1.145 $Y2=0.815
r108 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.145 $Y=0.265
+ $X2=1.22 $Y2=0.19
r109 5 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.145 $Y=0.265
+ $X2=1.145 $Y2=0.815
r110 1 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.965 $Y=1.675
+ $X2=0.965 $Y2=1.6
r111 1 3 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.965 $Y=1.675
+ $X2=0.965 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%CLK 3 7 11 12 13 14 15 20
c40 11 0 1.4009e-19 $X=4.4 $Y=1.66
r41 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.4 $Y=1.32
+ $X2=4.4 $Y2=1.32
r42 15 21 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=4.495 $Y=1.665
+ $X2=4.495 $Y2=1.32
r43 14 21 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=4.495 $Y=1.295
+ $X2=4.495 $Y2=1.32
r44 13 14 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.495 $Y=0.925
+ $X2=4.495 $Y2=1.295
r45 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.4 $Y=1.66 $X2=4.4
+ $Y2=1.32
r46 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.4 $Y=1.66 $X2=4.4
+ $Y2=1.825
r47 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.4 $Y=1.155
+ $X2=4.4 $Y2=1.32
r48 7 12 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.45 $Y=2.735
+ $X2=4.45 $Y2=1.825
r49 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.31 $Y=0.445
+ $X2=4.31 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_963_47# 1 2 9 13 17 21 23 27 32 33 36 37
+ 38 40 41 42 44 45 46 47 53 55 57 58 65 70
c176 70 0 1.91871e-19 $X=9.95 $Y=1.93
c177 58 0 1.62957e-19 $X=9.76 $Y=1.82
c178 53 0 1.4273e-19 $X=5.995 $Y=1.54
c179 46 0 6.69659e-20 $X=8.35 $Y=1.82
c180 42 0 1.47232e-19 $X=7.65 $Y=2.65
r181 69 70 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=9.915 $Y=1.93
+ $X2=9.95 $Y2=1.93
r182 65 66 53.4108 $w=3.7e-07 $l=4.1e-07 $layer=POLY_cond $X=6.13 $Y=1.41
+ $X2=6.54 $Y2=1.41
r183 62 69 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=9.775 $Y=1.93
+ $X2=9.915 $Y2=1.93
r184 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.775
+ $Y=1.93 $X2=9.775 $Y2=1.93
r185 58 61 4.22562 $w=2.98e-07 $l=1.1e-07 $layer=LI1_cond $X=9.76 $Y=1.82
+ $X2=9.76 $Y2=1.93
r186 54 65 17.5865 $w=3.7e-07 $l=1.35e-07 $layer=POLY_cond $X=5.995 $Y=1.41
+ $X2=6.13 $Y2=1.41
r187 53 56 8.97179 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=5.985 $Y=1.54
+ $X2=5.985 $Y2=1.705
r188 53 55 8.83798 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=5.985 $Y=1.54
+ $X2=5.985 $Y2=1.375
r189 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.995
+ $Y=1.54 $X2=5.995 $Y2=1.54
r190 47 50 4.10192 $w=2.93e-07 $l=1.05e-07 $layer=LI1_cond $X=4.972 $Y=0.34
+ $X2=4.972 $Y2=0.445
r191 45 58 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=9.61 $Y=1.82 $X2=9.76
+ $Y2=1.82
r192 45 46 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=9.61 $Y=1.82
+ $X2=8.35 $Y2=1.82
r193 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.265 $Y=1.905
+ $X2=8.35 $Y2=1.82
r194 43 44 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.265 $Y=1.905
+ $X2=8.265 $Y2=2.565
r195 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.18 $Y=2.65
+ $X2=8.265 $Y2=2.565
r196 41 42 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.18 $Y=2.65
+ $X2=7.65 $Y2=2.65
r197 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.565 $Y=2.565
+ $X2=7.65 $Y2=2.65
r198 39 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.565 $Y=2.105
+ $X2=7.565 $Y2=2.565
r199 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.48 $Y=2.02
+ $X2=7.565 $Y2=2.105
r200 37 38 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.48 $Y=2.02
+ $X2=6.79 $Y2=2.02
r201 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.705 $Y=2.105
+ $X2=6.79 $Y2=2.02
r202 35 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.705 $Y=2.105
+ $X2=6.705 $Y2=2.705
r203 34 57 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.09 $Y=2.87 $X2=6
+ $Y2=2.87
r204 33 36 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.62 $Y=2.87
+ $X2=6.705 $Y2=2.705
r205 33 34 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=6.62 $Y=2.87
+ $X2=6.09 $Y2=2.87
r206 32 57 3.59259 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=2.705 $X2=6
+ $Y2=2.87
r207 32 56 61.6162 $w=1.78e-07 $l=1e-06 $layer=LI1_cond $X=6 $Y=2.705 $X2=6
+ $Y2=1.705
r208 29 55 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=5.975 $Y=0.425
+ $X2=5.975 $Y2=1.375
r209 28 47 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=5.12 $Y=0.34
+ $X2=4.972 $Y2=0.34
r210 27 29 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.88 $Y=0.34
+ $X2=5.975 $Y2=0.425
r211 27 28 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.88 $Y=0.34
+ $X2=5.12 $Y2=0.34
r212 23 57 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.91 $Y=2.87 $X2=6
+ $Y2=2.87
r213 23 25 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=5.91 $Y=2.87
+ $X2=5.095 $Y2=2.87
r214 19 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.95 $Y=1.765
+ $X2=9.95 $Y2=1.93
r215 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=9.95 $Y=1.765
+ $X2=9.95 $Y2=0.945
r216 15 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.915 $Y=2.095
+ $X2=9.915 $Y2=1.93
r217 15 17 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.915 $Y=2.095
+ $X2=9.915 $Y2=2.525
r218 11 66 23.9667 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=6.54 $Y=1.115
+ $X2=6.54 $Y2=1.41
r219 11 13 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=6.54 $Y=1.115
+ $X2=6.54 $Y2=0.485
r220 7 65 23.9667 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=6.13 $Y=1.705
+ $X2=6.13 $Y2=1.41
r221 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.13 $Y=1.705
+ $X2=6.13 $Y2=2.285
r222 2 25 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=4.955
+ $Y=2.415 $X2=5.095 $Y2=2.87
r223 1 50 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.815
+ $Y=0.235 $X2=4.955 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_1365_29# 1 2 9 14 18 21 23 26 30 33 36
c61 18 0 9.66906e-20 $X=6.99 $Y=0.97
c62 14 0 2.25861e-19 $X=6.92 $Y=2.285
r63 34 36 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.92 $Y=1.135
+ $X2=6.92 $Y2=1.505
r64 28 30 26.5598 $w=1.88e-07 $l=4.55e-07 $layer=LI1_cond $X=7.915 $Y=1.765
+ $X2=7.915 $Y2=2.22
r65 26 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.01 $Y=1.67
+ $X2=7.01 $Y2=1.835
r66 26 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.01 $Y=1.67
+ $X2=7.01 $Y2=1.505
r67 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.01
+ $Y=1.67 $X2=7.01 $Y2=1.67
r68 23 28 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=7.82 $Y=1.675
+ $X2=7.915 $Y2=1.765
r69 23 25 49.9091 $w=1.78e-07 $l=8.1e-07 $layer=LI1_cond $X=7.82 $Y=1.675
+ $X2=7.01 $Y2=1.675
r70 18 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.99 $Y=0.97
+ $X2=6.99 $Y2=1.135
r71 18 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.99 $Y=0.97
+ $X2=6.99 $Y2=0.805
r72 17 21 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=6.99 $Y=0.89
+ $X2=7.71 $Y2=0.89
r73 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.99
+ $Y=0.97 $X2=6.99 $Y2=0.97
r74 14 37 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.92 $Y=2.285
+ $X2=6.92 $Y2=1.835
r75 9 33 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.9 $Y=0.485 $X2=6.9
+ $Y2=0.805
r76 2 30 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=2.075 $X2=7.915 $Y2=2.22
r77 1 21 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=7.585
+ $Y=0.625 $X2=7.71 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_1237_55# 1 2 9 11 13 16 18 20 22 25 28 31
+ 36 38 41 42 49
c96 41 0 1.80425e-19 $X=6.335 $Y=0.715
c97 31 0 7.86288e-20 $X=6.345 $Y=2.22
c98 28 0 9.66906e-20 $X=6.345 $Y=1.225
c99 11 0 1.35218e-19 $X=7.965 $Y=1.155
c100 9 0 6.69659e-20 $X=7.7 $Y=2.285
r101 39 49 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.92 $Y=1.34
+ $X2=9.085 $Y2=1.34
r102 39 46 14.0362 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=8.92 $Y=1.34 $X2=8.83
+ $Y2=1.34
r103 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.92
+ $Y=1.32 $X2=8.92 $Y2=1.32
r104 36 43 7.77419 $w=2.79e-07 $l=4.5e-08 $layer=POLY_cond $X=7.745 $Y=1.32
+ $X2=7.7 $Y2=1.32
r105 35 38 68.5885 $w=1.88e-07 $l=1.175e-06 $layer=LI1_cond $X=7.745 $Y=1.32
+ $X2=8.92 $Y2=1.32
r106 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.745
+ $Y=1.32 $X2=7.745 $Y2=1.32
r107 33 42 1.14861 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=6.45 $Y=1.32
+ $X2=6.355 $Y2=1.32
r108 33 35 75.5933 $w=1.88e-07 $l=1.295e-06 $layer=LI1_cond $X=6.45 $Y=1.32
+ $X2=7.745 $Y2=1.32
r109 29 42 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.355 $Y=1.415
+ $X2=6.355 $Y2=1.32
r110 29 31 46.9904 $w=1.88e-07 $l=8.05e-07 $layer=LI1_cond $X=6.355 $Y=1.415
+ $X2=6.355 $Y2=2.22
r111 28 42 5.40251 $w=1.8e-07 $l=9.98749e-08 $layer=LI1_cond $X=6.345 $Y=1.225
+ $X2=6.355 $Y2=1.32
r112 28 41 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.345 $Y=1.225
+ $X2=6.345 $Y2=0.715
r113 23 41 5.69365 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=6.335 $Y=0.62
+ $X2=6.335 $Y2=0.715
r114 23 25 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=6.335 $Y=0.62
+ $X2=6.335 $Y2=0.49
r115 20 22 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.59 $Y=1.375
+ $X2=9.59 $Y2=0.945
r116 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.515 $Y=1.45
+ $X2=9.59 $Y2=1.375
r117 18 49 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.515 $Y=1.45
+ $X2=9.085 $Y2=1.45
r118 14 46 23.9667 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=8.83 $Y=1.525
+ $X2=8.83 $Y2=1.34
r119 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.83 $Y=1.525
+ $X2=8.83 $Y2=2.315
r120 11 36 38.0072 $w=2.79e-07 $l=2.91033e-07 $layer=POLY_cond $X=7.965 $Y=1.155
+ $X2=7.745 $Y2=1.32
r121 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.965 $Y=1.155
+ $X2=7.965 $Y2=0.835
r122 7 43 17.2686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.7 $Y=1.485
+ $X2=7.7 $Y2=1.32
r123 7 9 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=7.7 $Y=1.485 $X2=7.7
+ $Y2=2.285
r124 2 31 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=2.075 $X2=6.345 $Y2=2.22
r125 1 25 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=6.185
+ $Y=0.275 $X2=6.325 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%SET_B 3 8 11 13 15 19 22 23 25 28 29 30 31
+ 32 41 45
c96 45 0 1.35218e-19 $X=9.738 $Y=0.452
c97 28 0 1.62831e-19 $X=10.87 $Y=0.382
c98 25 0 1.6681e-19 $X=11.925 $Y=1.67
c99 23 0 1.40857e-19 $X=11.04 $Y=1.675
r100 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.48
+ $Y=0.35 $X2=8.48 $Y2=0.35
r101 38 41 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=8.325 $Y=0.35
+ $X2=8.48 $Y2=0.35
r102 32 45 3.13464 $w=3.73e-07 $l=1.02e-07 $layer=LI1_cond $X=9.84 $Y=0.452
+ $X2=9.738 $Y2=0.452
r103 31 45 11.6166 $w=3.73e-07 $l=3.78e-07 $layer=LI1_cond $X=9.36 $Y=0.452
+ $X2=9.738 $Y2=0.452
r104 30 31 14.7513 $w=3.73e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=0.452
+ $X2=9.36 $Y2=0.452
r105 30 42 12.2927 $w=3.73e-07 $l=4e-07 $layer=LI1_cond $X=8.88 $Y=0.452
+ $X2=8.48 $Y2=0.452
r106 29 42 2.45854 $w=3.73e-07 $l=8e-08 $layer=LI1_cond $X=8.4 $Y=0.452 $X2=8.48
+ $Y2=0.452
r107 28 32 41.2722 $w=2.63e-07 $l=9.45e-07 $layer=LI1_cond $X=10.87 $Y=0.382
+ $X2=9.925 $Y2=0.382
r108 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.925
+ $Y=1.67 $X2=11.925 $Y2=1.67
r109 23 25 54.5303 $w=1.78e-07 $l=8.85e-07 $layer=LI1_cond $X=11.04 $Y=1.675
+ $X2=11.925 $Y2=1.675
r110 22 23 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=10.955 $Y=1.585
+ $X2=11.04 $Y2=1.675
r111 21 28 7.04737 $w=2.35e-07 $l=1.54771e-07 $layer=LI1_cond $X=10.955 $Y=0.5
+ $X2=10.87 $Y2=0.382
r112 21 22 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=10.955 $Y=0.5
+ $X2=10.955 $Y2=1.585
r113 17 19 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=8.225 $Y=1.62
+ $X2=8.325 $Y2=1.62
r114 13 26 38.7444 $w=2.79e-07 $l=1.90526e-07 $layer=POLY_cond $X=11.87 $Y=1.835
+ $X2=11.925 $Y2=1.67
r115 13 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=11.87 $Y=1.835
+ $X2=11.87 $Y2=2.385
r116 9 26 68.1135 $w=2.79e-07 $l=3.77326e-07 $layer=POLY_cond $X=11.835 $Y=1.335
+ $X2=11.925 $Y2=1.67
r117 9 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=11.835 $Y=1.335
+ $X2=11.835 $Y2=0.835
r118 6 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.325 $Y=1.545
+ $X2=8.325 $Y2=1.62
r119 6 8 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=8.325 $Y=1.545
+ $X2=8.325 $Y2=0.835
r120 5 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.325 $Y=0.515
+ $X2=8.325 $Y2=0.35
r121 5 8 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.325 $Y=0.515
+ $X2=8.325 $Y2=0.835
r122 1 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.225 $Y=1.695
+ $X2=8.225 $Y2=1.62
r123 1 3 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.225 $Y=1.695
+ $X2=8.225 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_794_47# 1 2 7 9 12 15 16 18 19 22 26 28
+ 30 32 35 38 39 41 43 46 47 49 51 52 55 62 65
c169 47 0 3.09915e-20 $X=4.855 $Y=2.09
c170 43 0 1.62957e-19 $X=10.72 $Y=1.755
c171 22 0 1.80425e-19 $X=6.11 $Y=0.485
c172 16 0 1.4273e-19 $X=6.035 $Y=1.06
c173 12 0 1.88293e-19 $X=4.88 $Y=2.735
r174 65 66 12.9577 $w=6.4e-07 $layer=POLY_cond $X=5.125 $Y=2.09 $X2=5.125
+ $Y2=2.09
r175 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.97
+ $Y=2.09 $X2=4.97 $Y2=2.09
r176 61 62 7.81899 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=2.16
+ $X2=4.305 $Y2=2.16
r177 58 61 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.05 $Y=2.16 $X2=4.14
+ $Y2=2.16
r178 55 57 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=4.097 $Y=0.445
+ $X2=4.097 $Y2=0.61
r179 52 66 43.8891 $w=6.4e-07 $l=6.8e-07 $layer=POLY_cond $X=5.125 $Y=1.41
+ $X2=5.125 $Y2=2.09
r180 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.97
+ $Y=1.41 $X2=4.97 $Y2=1.41
r181 49 64 2.88909 $w=2.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.995 $Y=1.995
+ $X2=4.995 $Y2=2.09
r182 49 51 24.0778 $w=2.78e-07 $l=5.85e-07 $layer=LI1_cond $X=4.995 $Y=1.995
+ $X2=4.995 $Y2=1.41
r183 47 64 4.25761 $w=1.9e-07 $l=1.4e-07 $layer=LI1_cond $X=4.855 $Y=2.09
+ $X2=4.995 $Y2=2.09
r184 47 62 32.1053 $w=1.88e-07 $l=5.5e-07 $layer=LI1_cond $X=4.855 $Y=2.09
+ $X2=4.305 $Y2=2.09
r185 46 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=1.995
+ $X2=4.05 $Y2=2.16
r186 46 57 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=4.05 $Y=1.995
+ $X2=4.05 $Y2=0.61
r187 43 44 64.8304 $w=1.71e-07 $l=2.3e-07 $layer=POLY_cond $X=10.72 $Y=1.755
+ $X2=10.95 $Y2=1.755
r188 39 52 22.9895 $w=6.4e-07 $l=2.75e-07 $layer=POLY_cond $X=5.125 $Y=1.135
+ $X2=5.125 $Y2=1.41
r189 39 40 12.1186 $w=6.4e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.125 $Y=1.135
+ $X2=5.2 $Y2=1.06
r190 37 44 5.94057 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=10.95 $Y=1.875
+ $X2=10.95 $Y2=1.755
r191 37 38 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=10.95 $Y=1.875
+ $X2=10.95 $Y2=3.075
r192 33 43 5.94057 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=10.72 $Y=1.635
+ $X2=10.72 $Y2=1.755
r193 33 35 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=10.72 $Y=1.635
+ $X2=10.72 $Y2=0.835
r194 30 43 73.2866 $w=1.71e-07 $l=2.6e-07 $layer=POLY_cond $X=10.46 $Y=1.755
+ $X2=10.72 $Y2=1.755
r195 30 32 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.46 $Y=1.785
+ $X2=10.46 $Y2=2.315
r196 29 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.635 $Y=3.15
+ $X2=6.56 $Y2=3.15
r197 28 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.875 $Y=3.15
+ $X2=10.95 $Y2=3.075
r198 28 29 2174.13 $w=1.5e-07 $l=4.24e-06 $layer=POLY_cond $X=10.875 $Y=3.15
+ $X2=6.635 $Y2=3.15
r199 24 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.56 $Y=3.075
+ $X2=6.56 $Y2=3.15
r200 24 26 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.56 $Y=3.075
+ $X2=6.56 $Y2=2.285
r201 20 22 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.11 $Y=0.985
+ $X2=6.11 $Y2=0.485
r202 18 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.485 $Y=3.15
+ $X2=6.56 $Y2=3.15
r203 18 19 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=6.485 $Y=3.15
+ $X2=5.445 $Y2=3.15
r204 17 40 26.1659 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=5.445 $Y=1.06
+ $X2=5.2 $Y2=1.06
r205 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.035 $Y=1.06
+ $X2=6.11 $Y2=0.985
r206 16 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.035 $Y=1.06
+ $X2=5.445 $Y2=1.06
r207 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.37 $Y=3.075
+ $X2=5.445 $Y2=3.15
r208 14 65 28.0482 $w=3.2e-07 $l=3.16938e-07 $layer=POLY_cond $X=5.37 $Y=2.255
+ $X2=5.125 $Y2=2.09
r209 14 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.37 $Y=2.255
+ $X2=5.37 $Y2=3.075
r210 10 65 28.0482 $w=3.2e-07 $l=3.16938e-07 $layer=POLY_cond $X=4.88 $Y=2.255
+ $X2=5.125 $Y2=2.09
r211 10 12 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.88 $Y=2.255
+ $X2=4.88 $Y2=2.735
r212 7 40 55.1563 $w=4.05e-07 $l=5.89322e-07 $layer=POLY_cond $X=4.74 $Y=0.765
+ $X2=5.2 $Y2=1.06
r213 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.74 $Y=0.765
+ $X2=4.74 $Y2=0.445
r214 2 61 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=2.085 $X2=4.14 $Y2=2.23
r215 1 55 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.97
+ $Y=0.235 $X2=4.095 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_2214_99# 1 2 7 9 12 14 17 21 23 25
c62 12 0 1.75145e-19 $X=11.44 $Y=2.385
c63 7 0 1.62831e-19 $X=11.145 $Y=1.155
r64 23 25 51.6465 $w=2.68e-07 $l=1.21e-06 $layer=LI1_cond $X=13.065 $Y=1.415
+ $X2=13.065 $Y2=2.625
r65 19 23 29.2677 $w=1.78e-07 $l=4.75e-07 $layer=LI1_cond $X=12.59 $Y=1.325
+ $X2=13.065 $Y2=1.325
r66 19 21 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=12.59 $Y=1.235
+ $X2=12.59 $Y2=0.83
r67 17 32 9.71062 $w=2.73e-07 $l=5.5e-08 $layer=POLY_cond $X=11.385 $Y=1.32
+ $X2=11.44 $Y2=1.32
r68 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.385
+ $Y=1.32 $X2=11.385 $Y2=1.32
r69 14 19 10.1667 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=12.425 $Y=1.325
+ $X2=12.59 $Y2=1.325
r70 14 16 64.0808 $w=1.78e-07 $l=1.04e-06 $layer=LI1_cond $X=12.425 $Y=1.325
+ $X2=11.385 $Y2=1.325
r71 10 32 16.7618 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.44 $Y=1.485
+ $X2=11.44 $Y2=1.32
r72 10 12 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=11.44 $Y=1.485
+ $X2=11.44 $Y2=2.385
r73 7 17 42.3736 $w=2.73e-07 $l=3.11769e-07 $layer=POLY_cond $X=11.145 $Y=1.155
+ $X2=11.385 $Y2=1.32
r74 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.145 $Y=1.155
+ $X2=11.145 $Y2=0.835
r75 2 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=12.895
+ $Y=2.415 $X2=13.035 $Y2=2.625
r76 1 21 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=12.45
+ $Y=0.625 $X2=12.59 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_1998_463# 1 2 3 12 16 18 22 24 26 28 30
+ 31 32 34 36 40 41 46
c99 41 0 1.6681e-19 $X=12.665 $Y=1.75
c100 34 0 1.75145e-19 $X=10.505 $Y=0.8
r101 46 47 15.535 $w=4.28e-07 $l=5.45e-07 $layer=LI1_cond $X=12.085 $Y=2.242
+ $X2=12.63 $Y2=2.242
r102 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.665
+ $Y=1.75 $X2=12.665 $Y2=1.75
r103 38 47 3.65327 $w=2.6e-07 $l=3.07e-07 $layer=LI1_cond $X=12.63 $Y=1.935
+ $X2=12.63 $Y2=2.242
r104 38 40 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=12.63 $Y=1.935
+ $X2=12.63 $Y2=1.75
r105 37 44 7.64692 $w=1.7e-07 $l=3.1496e-07 $layer=LI1_cond $X=10.7 $Y=2.02
+ $X2=10.39 $Y2=2.01
r106 36 46 8.29179 $w=4.28e-07 $l=2.79542e-07 $layer=LI1_cond $X=11.955 $Y=2.02
+ $X2=12.085 $Y2=2.242
r107 36 37 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=11.955 $Y=2.02
+ $X2=10.7 $Y2=2.02
r108 32 44 2.43745 $w=6.05e-07 $l=9.84378e-08 $layer=LI1_cond $X=10.397 $Y=1.915
+ $X2=10.39 $Y2=2.01
r109 32 34 22.0434 $w=6.03e-07 $l=1.115e-06 $layer=LI1_cond $X=10.397 $Y=1.915
+ $X2=10.397 $Y2=0.8
r110 29 41 43.3659 $w=3.95e-07 $l=3.08e-07 $layer=POLY_cond $X=12.697 $Y=2.058
+ $X2=12.697 $Y2=1.75
r111 29 30 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=12.697 $Y=2.058
+ $X2=12.697 $Y2=2.255
r112 27 41 3.51996 $w=3.95e-07 $l=2.5e-08 $layer=POLY_cond $X=12.697 $Y=1.725
+ $X2=12.697 $Y2=1.75
r113 27 28 12.1181 $w=2.72e-07 $l=1.32288e-07 $layer=POLY_cond $X=12.697
+ $Y=1.725 $X2=12.597 $Y2=1.65
r114 24 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.77 $Y=1.725
+ $X2=13.77 $Y2=1.65
r115 24 26 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=13.77 $Y=1.725
+ $X2=13.77 $Y2=2.155
r116 20 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.77 $Y=1.575
+ $X2=13.77 $Y2=1.65
r117 20 22 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=13.77 $Y=1.575
+ $X2=13.77 $Y2=0.865
r118 19 28 14.0569 $w=1.5e-07 $l=2.98e-07 $layer=POLY_cond $X=12.895 $Y=1.65
+ $X2=12.597 $Y2=1.65
r119 18 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.695 $Y=1.65
+ $X2=13.77 $Y2=1.65
r120 18 19 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=13.695 $Y=1.65
+ $X2=12.895 $Y2=1.65
r121 16 30 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=12.82 $Y=2.625
+ $X2=12.82 $Y2=2.255
r122 10 28 12.1181 $w=2.72e-07 $l=2.56776e-07 $layer=POLY_cond $X=12.375
+ $Y=1.575 $X2=12.597 $Y2=1.65
r123 10 12 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.375 $Y=1.575
+ $X2=12.375 $Y2=0.835
r124 3 46 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.945
+ $Y=2.175 $X2=12.085 $Y2=2.385
r125 2 44 600 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_PDIFF $count=1 $X=9.99
+ $Y=2.315 $X2=10.245 $Y2=2.02
r126 1 34 91 $w=1.7e-07 $l=5.60714e-07 $layer=licon1_NDIFF $count=2 $X=10.025
+ $Y=0.625 $X2=10.505 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_2686_131# 1 2 9 13 15 19 23 25 28 32 36
+ 39 40
r67 40 41 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=14.25 $Y=1.39
+ $X2=14.25 $Y2=1.315
r68 37 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=14.25 $Y=1.48
+ $X2=14.25 $Y2=1.645
r69 37 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=14.25 $Y=1.48
+ $X2=14.25 $Y2=1.39
r70 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.25
+ $Y=1.48 $X2=14.25 $Y2=1.48
r71 34 39 0.851123 $w=3.3e-07 $l=1.48e-07 $layer=LI1_cond $X=13.685 $Y=1.48
+ $X2=13.537 $Y2=1.48
r72 34 36 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=13.685 $Y=1.48
+ $X2=14.25 $Y2=1.48
r73 30 39 5.78497 $w=2.87e-07 $l=1.65e-07 $layer=LI1_cond $X=13.537 $Y=1.645
+ $X2=13.537 $Y2=1.48
r74 30 32 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=13.537 $Y=1.645
+ $X2=13.537 $Y2=1.98
r75 26 39 5.78497 $w=2.87e-07 $l=1.68464e-07 $layer=LI1_cond $X=13.53 $Y=1.315
+ $X2=13.537 $Y2=1.48
r76 26 28 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=13.53 $Y=1.315
+ $X2=13.53 $Y2=0.865
r77 21 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.71 $Y=1.465
+ $X2=14.71 $Y2=1.39
r78 21 23 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=14.71 $Y=1.465
+ $X2=14.71 $Y2=2.465
r79 17 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.71 $Y=1.315
+ $X2=14.71 $Y2=1.39
r80 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.71 $Y=1.315
+ $X2=14.71 $Y2=0.655
r81 16 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.415 $Y=1.39
+ $X2=14.25 $Y2=1.39
r82 15 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.635 $Y=1.39
+ $X2=14.71 $Y2=1.39
r83 15 16 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=14.635 $Y=1.39
+ $X2=14.415 $Y2=1.39
r84 13 43 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=14.28 $Y=2.465
+ $X2=14.28 $Y2=1.645
r85 9 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.28 $Y=0.655
+ $X2=14.28 $Y2=1.315
r86 2 32 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=13.43
+ $Y=1.835 $X2=13.555 $Y2=1.98
r87 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=13.43
+ $Y=0.655 $X2=13.555 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_39_481# 1 2 7 9 13
r24 11 16 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=0.415 $Y=2.52
+ $X2=0.285 $Y2=2.52
r25 11 13 76.7527 $w=2.48e-07 $l=1.665e-06 $layer=LI1_cond $X=0.415 $Y=2.52
+ $X2=2.08 $Y2=2.52
r26 7 16 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=0.285 $Y=2.645
+ $X2=0.285 $Y2=2.52
r27 7 9 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.285 $Y=2.645
+ $X2=0.285 $Y2=2.9
r28 2 13 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=2.405 $X2=2.08 $Y2=2.55
r29 1 16 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=2.405 $X2=0.32 $Y2=2.56
r30 1 9 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=2.405 $X2=0.32 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 58 62 64 69 70 72 73 75 76 78 79 81 82 83 85 97 120 128 133 136 139 143
c169 38 0 3.09915e-20 $X=4.665 $Y=2.93
r170 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r171 139 140 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r172 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r173 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r174 131 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r175 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r176 128 142 4.48049 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=14.76 $Y=3.33
+ $X2=15.06 $Y2=3.33
r177 128 130 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=14.76 $Y=3.33
+ $X2=14.64 $Y2=3.33
r178 127 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.64 $Y2=3.33
r179 127 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=12.72 $Y2=3.33
r180 126 127 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r181 124 139 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.76 $Y=3.33
+ $X2=12.6 $Y2=3.33
r182 124 126 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=12.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r183 123 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r184 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r185 120 139 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.44 $Y=3.33
+ $X2=12.6 $Y2=3.33
r186 120 122 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=12.44 $Y=3.33
+ $X2=12.24 $Y2=3.33
r187 119 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r188 118 119 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r189 116 119 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=11.28 $Y2=3.33
r190 115 118 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=11.28 $Y2=3.33
r191 115 116 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r192 113 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r193 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 109 112 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r195 109 110 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r196 107 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r197 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r198 104 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r199 104 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r200 103 106 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r201 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r202 101 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=3.33
+ $X2=4.665 $Y2=3.33
r203 101 103 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.83 $Y=3.33
+ $X2=5.04 $Y2=3.33
r204 100 137 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r205 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r206 97 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.5 $Y=3.33
+ $X2=4.665 $Y2=3.33
r207 97 99 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.5 $Y=3.33
+ $X2=3.12 $Y2=3.33
r208 96 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r209 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r210 93 96 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r211 93 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r212 92 95 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r213 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r214 90 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=0.75 $Y2=3.33
r215 90 92 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=1.2 $Y2=3.33
r216 88 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r217 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r218 85 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.75 $Y2=3.33
r219 85 87 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.24 $Y2=3.33
r220 83 113 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=8.4 $Y2=3.33
r221 83 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=7.44 $Y2=3.33
r222 81 126 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=13.855 $Y=3.33
+ $X2=13.68 $Y2=3.33
r223 81 82 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=13.855 $Y=3.33
+ $X2=14.037 $Y2=3.33
r224 80 130 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=14.22 $Y=3.33
+ $X2=14.64 $Y2=3.33
r225 80 82 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=14.22 $Y=3.33
+ $X2=14.037 $Y2=3.33
r226 78 118 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=11.53 $Y=3.33
+ $X2=11.28 $Y2=3.33
r227 78 79 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=11.53 $Y=3.33
+ $X2=11.657 $Y2=3.33
r228 77 122 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=11.785 $Y=3.33
+ $X2=12.24 $Y2=3.33
r229 77 79 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=11.785 $Y=3.33
+ $X2=11.657 $Y2=3.33
r230 75 112 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r231 75 76 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=8.52 $Y=3.33
+ $X2=8.632 $Y2=3.33
r232 74 115 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=8.745 $Y=3.33
+ $X2=8.88 $Y2=3.33
r233 74 76 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=8.745 $Y=3.33
+ $X2=8.632 $Y2=3.33
r234 72 106 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.98 $Y=3.33
+ $X2=6.96 $Y2=3.33
r235 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.98 $Y=3.33
+ $X2=7.145 $Y2=3.33
r236 71 109 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.31 $Y=3.33
+ $X2=7.44 $Y2=3.33
r237 71 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.31 $Y=3.33
+ $X2=7.145 $Y2=3.33
r238 69 95 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=2.64 $Y2=3.33
r239 69 70 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=2.895 $Y2=3.33
r240 68 99 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.025 $Y=3.33
+ $X2=3.12 $Y2=3.33
r241 68 70 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.025 $Y=3.33
+ $X2=2.895 $Y2=3.33
r242 64 67 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=14.925 $Y=2.25
+ $X2=14.925 $Y2=2.95
r243 62 142 3.28569 $w=3.3e-07 $l=1.72337e-07 $layer=LI1_cond $X=14.925 $Y=3.245
+ $X2=15.06 $Y2=3.33
r244 62 67 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=14.925 $Y=3.245
+ $X2=14.925 $Y2=2.95
r245 58 61 14.9975 $w=3.63e-07 $l=4.75e-07 $layer=LI1_cond $X=14.037 $Y=1.99
+ $X2=14.037 $Y2=2.465
r246 56 82 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=14.037 $Y=3.245
+ $X2=14.037 $Y2=3.33
r247 56 61 24.6275 $w=3.63e-07 $l=7.8e-07 $layer=LI1_cond $X=14.037 $Y=3.245
+ $X2=14.037 $Y2=2.465
r248 52 139 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=12.6 $Y=3.245
+ $X2=12.6 $Y2=3.33
r249 52 54 22.3286 $w=3.18e-07 $l=6.2e-07 $layer=LI1_cond $X=12.6 $Y=3.245
+ $X2=12.6 $Y2=2.625
r250 48 79 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=11.657 $Y=3.245
+ $X2=11.657 $Y2=3.33
r251 48 50 36.381 $w=2.53e-07 $l=8.05e-07 $layer=LI1_cond $X=11.657 $Y=3.245
+ $X2=11.657 $Y2=2.44
r252 44 76 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=8.632 $Y=3.245
+ $X2=8.632 $Y2=3.33
r253 44 46 51.4758 $w=2.23e-07 $l=1.005e-06 $layer=LI1_cond $X=8.632 $Y=3.245
+ $X2=8.632 $Y2=2.24
r254 40 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.145 $Y=3.245
+ $X2=7.145 $Y2=3.33
r255 40 42 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=7.145 $Y=3.245
+ $X2=7.145 $Y2=2.37
r256 36 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=3.245
+ $X2=4.665 $Y2=3.33
r257 36 38 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.665 $Y=3.245
+ $X2=4.665 $Y2=2.93
r258 32 70 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=3.245
+ $X2=2.895 $Y2=3.33
r259 32 34 34.5733 $w=2.58e-07 $l=7.8e-07 $layer=LI1_cond $X=2.895 $Y=3.245
+ $X2=2.895 $Y2=2.465
r260 28 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=3.245
+ $X2=0.75 $Y2=3.33
r261 28 30 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.75 $Y=3.245
+ $X2=0.75 $Y2=2.92
r262 9 67 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=14.785
+ $Y=1.835 $X2=14.925 $Y2=2.95
r263 9 64 400 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_PDIFF $count=1 $X=14.785
+ $Y=1.835 $X2=14.925 $Y2=2.25
r264 8 61 300 $w=1.7e-07 $l=7.31779e-07 $layer=licon1_PDIFF $count=2 $X=13.845
+ $Y=1.835 $X2=14.065 $Y2=2.465
r265 8 58 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=13.845
+ $Y=1.835 $X2=13.985 $Y2=1.99
r266 7 54 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=12.48
+ $Y=2.415 $X2=12.605 $Y2=2.625
r267 6 50 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=11.515
+ $Y=2.175 $X2=11.655 $Y2=2.44
r268 5 46 300 $w=1.7e-07 $l=4.77179e-07 $layer=licon1_PDIFF $count=2 $X=8.3
+ $Y=1.895 $X2=8.615 $Y2=2.24
r269 4 42 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=6.995
+ $Y=2.075 $X2=7.145 $Y2=2.37
r270 3 38 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=4.525
+ $Y=2.415 $X2=4.665 $Y2=2.93
r271 2 34 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.795
+ $Y=2.31 $X2=2.93 $Y2=2.465
r272 1 30 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=2.405 $X2=0.75 $Y2=2.92
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_244_121# 1 2 3 4 15 17 21 22 24 26 27 30
+ 31 32 33 35 39 41 42 46 51
c138 33 0 1.88293e-19 $X=4.66 $Y=2.58
c139 21 0 6.49935e-20 $X=2.425 $Y=1.277
r140 51 53 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=5.56 $Y=2.35 $X2=5.56
+ $Y2=2.44
r141 51 52 5.38305 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.56 $Y=2.35
+ $X2=5.56 $Y2=2.185
r142 46 48 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.745 $Y=2.44
+ $X2=4.745 $Y2=2.58
r143 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.235 $Y=2.58
+ $X2=4.235 $Y2=2.885
r144 39 52 51.8599 $w=3.28e-07 $l=1.485e-06 $layer=LI1_cond $X=5.545 $Y=0.7
+ $X2=5.545 $Y2=2.185
r145 36 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.83 $Y=2.44
+ $X2=4.745 $Y2=2.44
r146 35 53 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.38 $Y=2.44
+ $X2=5.56 $Y2=2.44
r147 35 36 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.38 $Y=2.44
+ $X2=4.83 $Y2=2.44
r148 34 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.32 $Y=2.58
+ $X2=4.235 $Y2=2.58
r149 33 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=2.58
+ $X2=4.745 $Y2=2.58
r150 33 34 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.66 $Y=2.58
+ $X2=4.32 $Y2=2.58
r151 31 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.15 $Y=2.885
+ $X2=4.235 $Y2=2.885
r152 31 32 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=4.15 $Y=2.885
+ $X2=3.365 $Y2=2.885
r153 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.28 $Y=2.8
+ $X2=3.365 $Y2=2.885
r154 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.28 $Y=2.12
+ $X2=3.28 $Y2=2.8
r155 28 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=2.035
+ $X2=2.51 $Y2=2.035
r156 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.195 $Y=2.035
+ $X2=3.28 $Y2=2.12
r157 27 28 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.195 $Y=2.035
+ $X2=2.595 $Y2=2.035
r158 25 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=2.12
+ $X2=2.51 $Y2=2.035
r159 25 26 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.51 $Y=2.12
+ $X2=2.51 $Y2=2.815
r160 24 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.95
+ $X2=2.51 $Y2=2.035
r161 23 24 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.51 $Y=1.405
+ $X2=2.51 $Y2=1.95
r162 21 23 7.17723 $w=2.55e-07 $l=1.65118e-07 $layer=LI1_cond $X=2.425 $Y=1.277
+ $X2=2.51 $Y2=1.405
r163 21 22 40.6745 $w=2.53e-07 $l=9e-07 $layer=LI1_cond $X=2.425 $Y=1.277
+ $X2=1.525 $Y2=1.277
r164 17 26 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.425 $Y=2.945
+ $X2=2.51 $Y2=2.815
r165 17 19 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=2.425 $Y=2.945
+ $X2=1.595 $Y2=2.945
r166 13 22 6.96323 $w=2.55e-07 $l=2.19499e-07 $layer=LI1_cond $X=1.36 $Y=1.15
+ $X2=1.525 $Y2=1.277
r167 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.36 $Y=1.15
+ $X2=1.36 $Y2=0.815
r168 4 51 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=5.52
+ $Y=2.075 $X2=5.645 $Y2=2.35
r169 3 19 600 $w=1.7e-07 $l=6.0469e-07 $layer=licon1_PDIFF $count=1 $X=1.4
+ $Y=2.405 $X2=1.595 $Y2=2.92
r170 2 39 182 $w=1.7e-07 $l=4.92189e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.275 $X2=5.545 $Y2=0.7
r171 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.22
+ $Y=0.605 $X2=1.36 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_1781_379# 1 2 9 12 14 15
c36 12 0 1.91871e-19 $X=9.045 $Y=2.24
r37 15 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=10.675 $Y=2.36
+ $X2=10.675 $Y2=2.45
r38 12 14 4.6879 $w=2.93e-07 $l=1.2e-07 $layer=LI1_cond $X=9.062 $Y=2.24
+ $X2=9.062 $Y2=2.36
r39 10 14 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=9.21 $Y=2.36
+ $X2=9.062 $Y2=2.36
r40 9 15 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.51 $Y=2.36
+ $X2=10.675 $Y2=2.36
r41 9 10 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=10.51 $Y=2.36
+ $X2=9.21 $Y2=2.36
r42 2 18 600 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=1 $X=10.535
+ $Y=1.895 $X2=10.675 $Y2=2.45
r43 1 12 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=8.905
+ $Y=1.895 $X2=9.045 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%A_1888_463# 1 2 7 11 14
r26 14 16 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=9.585 $Y=2.72
+ $X2=9.585 $Y2=2.88
r27 9 11 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=11.21 $Y=2.795
+ $X2=11.21 $Y2=2.44
r28 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.75 $Y=2.88
+ $X2=9.585 $Y2=2.88
r29 7 9 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=11.06 $Y=2.88
+ $X2=11.21 $Y2=2.795
r30 7 8 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=11.06 $Y=2.88
+ $X2=9.75 $Y2=2.88
r31 2 11 600 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_PDIFF $count=1 $X=11.1
+ $Y=2.175 $X2=11.225 $Y2=2.44
r32 1 14 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=9.44
+ $Y=2.315 $X2=9.585 $Y2=2.72
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%Q 1 2 9 13 17 20 23
r31 21 23 8.80447 $w=7.18e-07 $l=5.3e-07 $layer=LI1_cond $X=14.915 $Y=1.825
+ $X2=14.915 $Y2=1.295
r32 20 22 8.75285 $w=8.83e-07 $l=5e-09 $layer=LI1_cond $X=14.832 $Y=1.99
+ $X2=14.832 $Y2=1.995
r33 20 21 2.73456 $w=8.83e-07 $l=1.65e-07 $layer=LI1_cond $X=14.832 $Y=1.99
+ $X2=14.832 $Y2=1.825
r34 17 23 2.65795 $w=7.18e-07 $l=1.6e-07 $layer=LI1_cond $X=14.915 $Y=1.135
+ $X2=14.915 $Y2=1.295
r35 16 17 9.83367 $w=7.18e-07 $l=1.7e-07 $layer=LI1_cond $X=14.832 $Y=0.965
+ $X2=14.832 $Y2=1.135
r36 13 22 50.7409 $w=1.98e-07 $l=9.15e-07 $layer=LI1_cond $X=14.49 $Y=2.91
+ $X2=14.49 $Y2=1.995
r37 9 16 30.2227 $w=1.98e-07 $l=5.45e-07 $layer=LI1_cond $X=14.49 $Y=0.42
+ $X2=14.49 $Y2=0.965
r38 2 20 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=14.355
+ $Y=1.835 $X2=14.495 $Y2=1.99
r39 2 13 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=14.355
+ $Y=1.835 $X2=14.495 $Y2=2.91
r40 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=14.355
+ $Y=0.235 $X2=14.495 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_2%VGND 1 2 3 4 5 6 7 8 27 31 35 39 42 43 47
+ 51 55 59 61 64 65 67 68 70 71 72 74 79 84 92 113 118 121 124 127 131
r154 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r155 127 128 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r156 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r157 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r158 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r159 116 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r160 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r161 113 130 4.48049 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=14.76 $Y=0 $X2=15.06
+ $Y2=0
r162 113 115 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=14.76 $Y=0
+ $X2=14.64 $Y2=0
r163 112 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.64 $Y2=0
r164 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r165 109 112 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.68 $Y2=0
r166 108 111 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.68 $Y2=0
r167 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r168 106 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r169 105 106 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r170 103 106 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=11.76 $Y2=0
r171 102 105 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=8.4 $Y=0
+ $X2=11.76 $Y2=0
r172 102 103 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r173 100 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r174 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r175 97 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.28 $Y=0
+ $X2=7.115 $Y2=0
r176 97 99 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=7.28 $Y=0 $X2=7.92
+ $Y2=0
r177 96 128 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r178 96 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r179 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r180 93 124 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.655 $Y=0
+ $X2=4.527 $Y2=0
r181 93 95 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.655 $Y=0
+ $X2=5.04 $Y2=0
r182 92 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.95 $Y=0
+ $X2=7.115 $Y2=0
r183 92 95 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=6.95 $Y=0 $X2=5.04
+ $Y2=0
r184 91 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r185 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r186 88 91 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.08 $Y2=0
r187 88 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r188 87 90 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r189 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r190 85 121 12.9614 $w=1.7e-07 $l=3.18e-07 $layer=LI1_cond $X=2.62 $Y=0
+ $X2=2.302 $Y2=0
r191 85 87 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.62 $Y=0 $X2=2.64
+ $Y2=0
r192 84 124 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.4 $Y=0 $X2=4.527
+ $Y2=0
r193 84 90 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.4 $Y=0 $X2=4.08
+ $Y2=0
r194 83 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r195 83 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=0.72 $Y2=0
r196 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r197 80 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=0
+ $X2=0.57 $Y2=0
r198 80 82 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=0.735 $Y=0
+ $X2=1.68 $Y2=0
r199 79 121 12.9614 $w=1.7e-07 $l=3.17e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=2.302 $Y2=0
r200 79 82 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=1.68 $Y2=0
r201 77 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r202 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r203 74 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.405 $Y=0
+ $X2=0.57 $Y2=0
r204 74 76 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.405 $Y=0
+ $X2=0.24 $Y2=0
r205 72 100 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=7.92 $Y2=0
r206 72 128 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=6.96 $Y2=0
r207 70 111 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=13.84 $Y=0
+ $X2=13.68 $Y2=0
r208 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.84 $Y=0
+ $X2=14.005 $Y2=0
r209 69 115 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=14.17 $Y=0
+ $X2=14.64 $Y2=0
r210 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.17 $Y=0
+ $X2=14.005 $Y2=0
r211 67 105 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=11.885 $Y=0
+ $X2=11.76 $Y2=0
r212 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.885 $Y=0
+ $X2=12.05 $Y2=0
r213 66 108 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=12.215 $Y=0
+ $X2=12.24 $Y2=0
r214 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.215 $Y=0
+ $X2=12.05 $Y2=0
r215 64 99 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.965 $Y=0 $X2=7.92
+ $Y2=0
r216 64 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.965 $Y=0 $X2=8.05
+ $Y2=0
r217 63 102 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.135 $Y=0
+ $X2=8.4 $Y2=0
r218 63 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.135 $Y=0 $X2=8.05
+ $Y2=0
r219 59 130 3.28569 $w=3.3e-07 $l=1.72337e-07 $layer=LI1_cond $X=14.925 $Y=0.085
+ $X2=15.06 $Y2=0
r220 59 61 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=14.925 $Y=0.085
+ $X2=14.925 $Y2=0.36
r221 55 57 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=14.005 $Y=0.41
+ $X2=14.005 $Y2=0.93
r222 53 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.005 $Y=0.085
+ $X2=14.005 $Y2=0
r223 53 55 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=14.005 $Y=0.085
+ $X2=14.005 $Y2=0.41
r224 49 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.05 $Y=0.085
+ $X2=12.05 $Y2=0
r225 49 51 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=12.05 $Y=0.085
+ $X2=12.05 $Y2=0.83
r226 45 47 46.3045 $w=1.98e-07 $l=8.35e-07 $layer=LI1_cond $X=8.54 $Y=0.91
+ $X2=9.375 $Y2=0.91
r227 43 45 22.4591 $w=1.98e-07 $l=4.05e-07 $layer=LI1_cond $X=8.135 $Y=0.91
+ $X2=8.54 $Y2=0.91
r228 42 43 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=8.05 $Y=0.81
+ $X2=8.135 $Y2=0.91
r229 41 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.05 $Y=0.085
+ $X2=8.05 $Y2=0
r230 41 42 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.05 $Y=0.085
+ $X2=8.05 $Y2=0.81
r231 37 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.115 $Y=0.085
+ $X2=7.115 $Y2=0
r232 37 39 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=7.115 $Y=0.085
+ $X2=7.115 $Y2=0.445
r233 33 124 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.527 $Y=0.085
+ $X2=4.527 $Y2=0
r234 33 35 16.2698 $w=2.53e-07 $l=3.6e-07 $layer=LI1_cond $X=4.527 $Y=0.085
+ $X2=4.527 $Y2=0.445
r235 29 121 2.65008 $w=6.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.302 $Y=0.085
+ $X2=2.302 $Y2=0
r236 29 31 13.7502 $w=6.33e-07 $l=7.3e-07 $layer=LI1_cond $X=2.302 $Y=0.085
+ $X2=2.302 $Y2=0.815
r237 25 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.57 $Y=0.085
+ $X2=0.57 $Y2=0
r238 25 27 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=0.57 $Y=0.085
+ $X2=0.57 $Y2=0.815
r239 8 61 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=14.785
+ $Y=0.235 $X2=14.925 $Y2=0.36
r240 7 57 182 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_NDIFF $count=1 $X=13.845
+ $Y=0.655 $X2=14.005 $Y2=0.93
r241 7 55 182 $w=1.7e-07 $l=3.37528e-07 $layer=licon1_NDIFF $count=1 $X=13.845
+ $Y=0.655 $X2=14.065 $Y2=0.41
r242 6 51 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=11.91
+ $Y=0.625 $X2=12.05 $Y2=0.83
r243 5 47 121.333 $w=1.7e-07 $l=1.10618e-06 $layer=licon1_NDIFF $count=1 $X=8.4
+ $Y=0.625 $X2=9.375 $Y2=0.905
r244 5 45 121.333 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=8.4
+ $Y=0.625 $X2=8.54 $Y2=0.905
r245 4 39 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=6.975
+ $Y=0.275 $X2=7.115 $Y2=0.445
r246 3 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.235 $X2=4.525 $Y2=0.445
r247 2 31 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.605 $X2=2.49 $Y2=0.815
r248 1 27 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.445
+ $Y=0.605 $X2=0.57 $Y2=0.815
.ends

