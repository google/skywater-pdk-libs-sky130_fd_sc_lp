* File: sky130_fd_sc_lp__nor3b_m.pxi.spice
* Created: Fri Aug 28 10:56:58 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3B_M%C_N N_C_N_c_67_n N_C_N_M1005_g N_C_N_c_61_n
+ N_C_N_M1003_g N_C_N_c_62_n N_C_N_c_63_n N_C_N_c_64_n C_N C_N N_C_N_c_66_n
+ PM_SKY130_FD_SC_LP__NOR3B_M%C_N
x_PM_SKY130_FD_SC_LP__NOR3B_M%A N_A_M1000_g N_A_M1004_g N_A_c_100_n N_A_c_101_n
+ A A N_A_c_102_n N_A_c_103_n PM_SKY130_FD_SC_LP__NOR3B_M%A
x_PM_SKY130_FD_SC_LP__NOR3B_M%B N_B_c_147_n N_B_M1001_g N_B_M1006_g N_B_c_144_n
+ N_B_c_149_n B B N_B_c_146_n PM_SKY130_FD_SC_LP__NOR3B_M%B
x_PM_SKY130_FD_SC_LP__NOR3B_M%A_27_439# N_A_27_439#_M1003_s N_A_27_439#_M1005_s
+ N_A_27_439#_M1007_g N_A_27_439#_c_186_n N_A_27_439#_M1002_g
+ N_A_27_439#_c_187_n N_A_27_439#_c_194_n N_A_27_439#_c_188_n
+ N_A_27_439#_c_189_n N_A_27_439#_c_195_n N_A_27_439#_c_190_n
+ N_A_27_439#_c_197_n N_A_27_439#_c_198_n N_A_27_439#_c_199_n
+ N_A_27_439#_c_191_n N_A_27_439#_c_240_p N_A_27_439#_c_200_n
+ N_A_27_439#_c_201_n PM_SKY130_FD_SC_LP__NOR3B_M%A_27_439#
x_PM_SKY130_FD_SC_LP__NOR3B_M%VPWR N_VPWR_M1005_d N_VPWR_c_269_n VPWR
+ N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_268_n N_VPWR_c_273_n
+ PM_SKY130_FD_SC_LP__NOR3B_M%VPWR
x_PM_SKY130_FD_SC_LP__NOR3B_M%Y N_Y_M1004_d N_Y_M1002_d N_Y_M1007_d N_Y_c_295_n
+ Y Y Y Y Y PM_SKY130_FD_SC_LP__NOR3B_M%Y
x_PM_SKY130_FD_SC_LP__NOR3B_M%VGND N_VGND_M1003_d N_VGND_M1006_d N_VGND_c_329_n
+ N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n VGND
+ N_VGND_c_334_n N_VGND_c_335_n N_VGND_c_336_n PM_SKY130_FD_SC_LP__NOR3B_M%VGND
cc_1 VNB N_C_N_c_61_n 0.0190963f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.795
cc_2 VNB N_C_N_c_62_n 0.0216955f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.215
cc_3 VNB N_C_N_c_63_n 0.0240876f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.72
cc_4 VNB N_C_N_c_64_n 0.029165f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.87
cc_5 VNB C_N 0.0257366f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_C_N_c_66_n 0.0196146f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_7 VNB N_A_M1004_g 0.0326366f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.495
cc_8 VNB N_A_c_100_n 0.0236905f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.72
cc_9 VNB N_A_c_101_n 0.00315406f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=0.87
cc_10 VNB N_A_c_102_n 0.0173358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_103_n 0.00714969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_M1006_g 0.0350658f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.795
cc_13 VNB N_B_c_144_n 0.00592118f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_14 VNB B 0.00533186f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.87
cc_15 VNB N_B_c_146_n 0.0370796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_439#_c_186_n 0.0198176f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.72
cc_17 VNB N_A_27_439#_c_187_n 0.0411724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_439#_c_188_n 0.0218213f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_19 VNB N_A_27_439#_c_189_n 0.0194252f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.665
cc_20 VNB N_A_27_439#_c_190_n 0.0123097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_439#_c_191_n 0.0156462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_268_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_23 VNB N_Y_c_295_n 0.0209826f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=0.87
cc_24 VNB Y 0.0289671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB Y 0.0272754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_329_n 0.00617492f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.38
cc_27 VNB N_VGND_c_330_n 0.019416f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.72
cc_28 VNB N_VGND_c_331_n 0.00626661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_332_n 0.0236734f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_30 VNB N_VGND_c_333_n 0.00362871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_334_n 0.0169445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_335_n 0.165042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_336_n 0.00401277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_C_N_c_67_n 0.020591f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.12
cc_35 VPB N_C_N_c_63_n 0.0560359f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.72
cc_36 VPB C_N 0.0112827f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_37 VPB N_A_M1000_g 0.0343476f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.12
cc_38 VPB N_A_c_101_n 0.0135039f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=0.87
cc_39 VPB N_A_c_103_n 0.00380662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_B_c_147_n 0.0151442f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=0.945
cc_41 VPB N_B_c_144_n 0.0178267f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.38
cc_42 VPB N_B_c_149_n 0.0177405f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=0.87
cc_43 VPB B 0.00377893f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.87
cc_44 VPB N_A_27_439#_M1007_g 0.0191427f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.215
cc_45 VPB N_A_27_439#_c_187_n 0.0178035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_27_439#_c_194_n 0.0295983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_27_439#_c_195_n 0.00185509f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_27_439#_c_190_n 0.00741223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_27_439#_c_197_n 0.00784371f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_27_439#_c_198_n 0.00248194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_27_439#_c_199_n 0.0183763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_27_439#_c_200_n 0.0219315f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_27_439#_c_201_n 0.0475215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_269_n 0.0395751f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.795
cc_55 VPB N_VPWR_c_270_n 0.0210774f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.215
cc_56 VPB N_VPWR_c_271_n 0.0457141f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.38
cc_57 VPB N_VPWR_c_268_n 0.0802623f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.38
cc_58 VPB N_VPWR_c_273_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB Y 0.0366705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 N_C_N_c_63_n N_A_M1000_g 0.0190531f $X=0.27 $Y=1.72 $X2=0 $Y2=0
cc_61 N_C_N_c_61_n N_A_M1004_g 0.0191366f $X=0.635 $Y=0.795 $X2=0 $Y2=0
cc_62 N_C_N_c_62_n N_A_M1004_g 0.0021227f $X=0.27 $Y=1.215 $X2=0 $Y2=0
cc_63 N_C_N_c_66_n N_A_c_100_n 0.00466505f $X=0.27 $Y=1.38 $X2=0 $Y2=0
cc_64 N_C_N_c_63_n N_A_c_101_n 0.00466505f $X=0.27 $Y=1.72 $X2=0 $Y2=0
cc_65 N_C_N_c_62_n N_A_c_102_n 0.00466505f $X=0.27 $Y=1.215 $X2=0 $Y2=0
cc_66 N_C_N_c_61_n N_A_27_439#_c_189_n 0.00286136f $X=0.635 $Y=0.795 $X2=0 $Y2=0
cc_67 N_C_N_c_64_n N_A_27_439#_c_189_n 0.00742642f $X=0.635 $Y=0.87 $X2=0 $Y2=0
cc_68 N_C_N_c_67_n N_A_27_439#_c_195_n 0.00832603f $X=0.475 $Y=2.12 $X2=0 $Y2=0
cc_69 N_C_N_c_63_n N_A_27_439#_c_195_n 0.00637268f $X=0.27 $Y=1.72 $X2=0 $Y2=0
cc_70 C_N N_A_27_439#_c_195_n 6.85577e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 N_C_N_c_62_n N_A_27_439#_c_190_n 0.0116665f $X=0.27 $Y=1.215 $X2=0 $Y2=0
cc_72 N_C_N_c_63_n N_A_27_439#_c_190_n 0.00219282f $X=0.27 $Y=1.72 $X2=0 $Y2=0
cc_73 N_C_N_c_64_n N_A_27_439#_c_190_n 9.95341e-19 $X=0.635 $Y=0.87 $X2=0 $Y2=0
cc_74 C_N N_A_27_439#_c_190_n 0.0546211f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_C_N_c_67_n N_A_27_439#_c_199_n 0.00706427f $X=0.475 $Y=2.12 $X2=0 $Y2=0
cc_76 N_C_N_c_63_n N_A_27_439#_c_199_n 0.00794076f $X=0.27 $Y=1.72 $X2=0 $Y2=0
cc_77 C_N N_A_27_439#_c_199_n 0.0264307f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_C_N_c_62_n N_A_27_439#_c_191_n 0.0039479f $X=0.27 $Y=1.215 $X2=0 $Y2=0
cc_79 N_C_N_c_64_n N_A_27_439#_c_191_n 0.0163796f $X=0.635 $Y=0.87 $X2=0 $Y2=0
cc_80 C_N N_A_27_439#_c_191_n 0.0138836f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_C_N_c_67_n N_VPWR_c_269_n 0.00498548f $X=0.475 $Y=2.12 $X2=0 $Y2=0
cc_82 N_C_N_c_67_n N_VPWR_c_270_n 0.00370896f $X=0.475 $Y=2.12 $X2=0 $Y2=0
cc_83 N_C_N_c_67_n N_VPWR_c_268_n 0.00445256f $X=0.475 $Y=2.12 $X2=0 $Y2=0
cc_84 N_C_N_c_61_n Y 6.67093e-19 $X=0.635 $Y=0.795 $X2=0 $Y2=0
cc_85 N_C_N_c_61_n N_VGND_c_329_n 0.00290325f $X=0.635 $Y=0.795 $X2=0 $Y2=0
cc_86 N_C_N_c_61_n N_VGND_c_332_n 0.0053602f $X=0.635 $Y=0.795 $X2=0 $Y2=0
cc_87 N_C_N_c_61_n N_VGND_c_335_n 0.00650215f $X=0.635 $Y=0.795 $X2=0 $Y2=0
cc_88 N_C_N_c_64_n N_VGND_c_335_n 7.53157e-19 $X=0.635 $Y=0.87 $X2=0 $Y2=0
cc_89 N_A_M1004_g N_B_M1006_g 0.0284093f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_90 N_A_c_102_n N_B_M1006_g 0.0123535f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_91 N_A_c_103_n N_B_M1006_g 0.00636821f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_92 N_A_M1000_g N_B_c_144_n 0.0069703f $X=1.015 $Y=2.405 $X2=0 $Y2=0
cc_93 N_A_c_101_n N_B_c_144_n 0.0123535f $X=1.03 $Y=1.775 $X2=0 $Y2=0
cc_94 N_A_M1000_g N_B_c_149_n 0.0479865f $X=1.015 $Y=2.405 $X2=0 $Y2=0
cc_95 N_A_c_103_n N_B_c_149_n 0.00101965f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_96 N_A_c_102_n B 5.0476e-19 $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_97 N_A_c_103_n B 0.0494619f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_98 N_A_c_100_n N_B_c_146_n 0.0123535f $X=1.03 $Y=1.61 $X2=0 $Y2=0
cc_99 N_A_M1000_g N_A_27_439#_c_190_n 0.00480985f $X=1.015 $Y=2.405 $X2=0 $Y2=0
cc_100 N_A_M1004_g N_A_27_439#_c_190_n 0.00252687f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_101 N_A_c_102_n N_A_27_439#_c_190_n 0.00625632f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_102 N_A_c_103_n N_A_27_439#_c_190_n 0.0584981f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_103 N_A_M1000_g N_A_27_439#_c_197_n 0.0149818f $X=1.015 $Y=2.405 $X2=0 $Y2=0
cc_104 N_A_c_101_n N_A_27_439#_c_197_n 0.00330292f $X=1.03 $Y=1.775 $X2=0 $Y2=0
cc_105 N_A_c_103_n N_A_27_439#_c_197_n 0.0301339f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_106 N_A_M1000_g N_A_27_439#_c_199_n 6.53268e-19 $X=1.015 $Y=2.405 $X2=0 $Y2=0
cc_107 N_A_M1004_g N_A_27_439#_c_191_n 0.00233011f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_108 N_A_M1000_g N_VPWR_c_269_n 0.00387667f $X=1.015 $Y=2.405 $X2=0 $Y2=0
cc_109 N_A_M1000_g N_VPWR_c_271_n 0.00370896f $X=1.015 $Y=2.405 $X2=0 $Y2=0
cc_110 N_A_M1000_g N_VPWR_c_268_n 0.00445256f $X=1.015 $Y=2.405 $X2=0 $Y2=0
cc_111 N_A_c_103_n Y 0.00475788f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_112 N_A_M1004_g Y 0.0108314f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_113 N_A_c_102_n Y 4.14396e-19 $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_114 N_A_c_103_n Y 0.019464f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_115 N_A_M1004_g N_VGND_c_329_n 0.00280551f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_116 N_A_c_102_n N_VGND_c_329_n 0.00228717f $X=1.03 $Y=1.27 $X2=0 $Y2=0
cc_117 N_A_M1004_g N_VGND_c_330_n 0.00507086f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_118 N_A_M1004_g N_VGND_c_335_n 0.00945726f $X=1.065 $Y=0.495 $X2=0 $Y2=0
cc_119 N_B_c_147_n N_A_27_439#_M1007_g 0.0176783f $X=1.375 $Y=2.12 $X2=0 $Y2=0
cc_120 N_B_c_149_n N_A_27_439#_M1007_g 0.00511192f $X=1.495 $Y=2.045 $X2=0 $Y2=0
cc_121 N_B_M1006_g N_A_27_439#_c_186_n 0.0215315f $X=1.495 $Y=0.495 $X2=0 $Y2=0
cc_122 N_B_M1006_g N_A_27_439#_c_187_n 0.00460661f $X=1.495 $Y=0.495 $X2=0 $Y2=0
cc_123 N_B_c_144_n N_A_27_439#_c_187_n 0.00862219f $X=1.495 $Y=1.97 $X2=0 $Y2=0
cc_124 B N_A_27_439#_c_187_n 0.00216863f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_B_c_146_n N_A_27_439#_c_187_n 0.0197331f $X=1.625 $Y=1.345 $X2=0 $Y2=0
cc_126 N_B_c_144_n N_A_27_439#_c_194_n 0.00511192f $X=1.495 $Y=1.97 $X2=0 $Y2=0
cc_127 N_B_c_147_n N_A_27_439#_c_197_n 0.0101584f $X=1.375 $Y=2.12 $X2=0 $Y2=0
cc_128 N_B_c_149_n N_A_27_439#_c_197_n 0.0132312f $X=1.495 $Y=2.045 $X2=0 $Y2=0
cc_129 B N_A_27_439#_c_197_n 0.0199524f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_B_c_146_n N_A_27_439#_c_197_n 9.46968e-19 $X=1.625 $Y=1.345 $X2=0 $Y2=0
cc_131 N_B_c_147_n N_A_27_439#_c_198_n 0.0107414f $X=1.375 $Y=2.12 $X2=0 $Y2=0
cc_132 N_B_c_147_n N_VPWR_c_271_n 0.00370896f $X=1.375 $Y=2.12 $X2=0 $Y2=0
cc_133 N_B_c_147_n N_VPWR_c_268_n 0.00445256f $X=1.375 $Y=2.12 $X2=0 $Y2=0
cc_134 N_B_M1006_g Y 0.00232786f $X=1.495 $Y=0.495 $X2=0 $Y2=0
cc_135 N_B_c_144_n Y 0.00287276f $X=1.495 $Y=1.97 $X2=0 $Y2=0
cc_136 B Y 0.0471601f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_137 N_B_c_146_n Y 0.00116364f $X=1.625 $Y=1.345 $X2=0 $Y2=0
cc_138 N_B_M1006_g Y 0.0219752f $X=1.495 $Y=0.495 $X2=0 $Y2=0
cc_139 B Y 0.0252256f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B_c_146_n Y 0.00160297f $X=1.625 $Y=1.345 $X2=0 $Y2=0
cc_141 N_B_M1006_g N_VGND_c_330_n 0.00438487f $X=1.495 $Y=0.495 $X2=0 $Y2=0
cc_142 N_B_M1006_g N_VGND_c_331_n 0.00284292f $X=1.495 $Y=0.495 $X2=0 $Y2=0
cc_143 N_B_M1006_g N_VGND_c_335_n 0.00711361f $X=1.495 $Y=0.495 $X2=0 $Y2=0
cc_144 N_A_27_439#_c_197_n N_VPWR_M1005_d 0.00113743f $X=1.655 $Y=2.14 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_27_439#_c_240_p N_VPWR_M1005_d 0.00190894f $X=0.69 $Y=2.14 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_27_439#_c_197_n N_VPWR_c_269_n 0.00875025f $X=1.655 $Y=2.14 $X2=0
+ $Y2=0
cc_147 N_A_27_439#_c_240_p N_VPWR_c_269_n 0.0151472f $X=0.69 $Y=2.14 $X2=0 $Y2=0
cc_148 N_A_27_439#_c_200_n N_VPWR_c_271_n 0.0213969f $X=1.825 $Y=2.945 $X2=0
+ $Y2=0
cc_149 N_A_27_439#_c_201_n N_VPWR_c_271_n 0.00606749f $X=1.825 $Y=2.945 $X2=0
+ $Y2=0
cc_150 N_A_27_439#_c_199_n N_VPWR_c_268_n 0.0118826f $X=0.267 $Y=2.14 $X2=0
+ $Y2=0
cc_151 N_A_27_439#_c_200_n N_VPWR_c_268_n 0.0112432f $X=1.825 $Y=2.945 $X2=0
+ $Y2=0
cc_152 N_A_27_439#_c_201_n N_VPWR_c_268_n 0.00840148f $X=1.825 $Y=2.945 $X2=0
+ $Y2=0
cc_153 N_A_27_439#_c_197_n A_218_439# 0.00366293f $X=1.655 $Y=2.14 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_27_439#_c_197_n A_290_439# 0.00560887f $X=1.655 $Y=2.14 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_27_439#_c_198_n A_290_439# 0.00462479f $X=1.74 $Y=2.78 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_27_439#_c_186_n N_Y_c_295_n 0.00326899f $X=1.925 $Y=0.815 $X2=0 $Y2=0
cc_157 N_A_27_439#_M1007_g Y 0.00251199f $X=1.895 $Y=2.405 $X2=0 $Y2=0
cc_158 N_A_27_439#_c_187_n Y 0.033583f $X=2.105 $Y=1.935 $X2=0 $Y2=0
cc_159 N_A_27_439#_c_194_n Y 0.0117263f $X=2.105 $Y=2.01 $X2=0 $Y2=0
cc_160 N_A_27_439#_c_197_n Y 0.0121725f $X=1.655 $Y=2.14 $X2=0 $Y2=0
cc_161 N_A_27_439#_c_186_n Y 0.00634851f $X=1.925 $Y=0.815 $X2=0 $Y2=0
cc_162 N_A_27_439#_c_187_n Y 0.00209759f $X=2.105 $Y=1.935 $X2=0 $Y2=0
cc_163 N_A_27_439#_c_188_n Y 0.016001f $X=2.105 $Y=0.89 $X2=0 $Y2=0
cc_164 N_A_27_439#_c_189_n Y 0.00496162f $X=0.42 $Y=0.495 $X2=0 $Y2=0
cc_165 N_A_27_439#_c_191_n Y 0.00591099f $X=0.69 $Y=0.905 $X2=0 $Y2=0
cc_166 N_A_27_439#_c_191_n N_VGND_c_329_n 0.00109477f $X=0.69 $Y=0.905 $X2=0
+ $Y2=0
cc_167 N_A_27_439#_c_186_n N_VGND_c_331_n 0.00269517f $X=1.925 $Y=0.815 $X2=0
+ $Y2=0
cc_168 N_A_27_439#_c_189_n N_VGND_c_332_n 0.0119771f $X=0.42 $Y=0.495 $X2=0
+ $Y2=0
cc_169 N_A_27_439#_c_186_n N_VGND_c_334_n 0.00439066f $X=1.925 $Y=0.815 $X2=0
+ $Y2=0
cc_170 N_A_27_439#_c_186_n N_VGND_c_335_n 0.0075491f $X=1.925 $Y=0.815 $X2=0
+ $Y2=0
cc_171 N_A_27_439#_c_189_n N_VGND_c_335_n 0.00991124f $X=0.42 $Y=0.495 $X2=0
+ $Y2=0
cc_172 N_A_27_439#_c_191_n N_VGND_c_335_n 0.0067504f $X=0.69 $Y=0.905 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_268_n Y 0.0119058f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_174 Y N_VGND_c_330_n 0.00945977f $X=2.16 $Y=0.925 $X2=0 $Y2=0
cc_175 N_Y_c_295_n N_VGND_c_331_n 0.00151731f $X=2.14 $Y=0.43 $X2=0 $Y2=0
cc_176 Y N_VGND_c_331_n 0.0153252f $X=2.16 $Y=0.925 $X2=0 $Y2=0
cc_177 N_Y_c_295_n N_VGND_c_334_n 0.0200925f $X=2.14 $Y=0.43 $X2=0 $Y2=0
cc_178 Y N_VGND_c_334_n 0.001622f $X=2.16 $Y=0.925 $X2=0 $Y2=0
cc_179 N_Y_c_295_n N_VGND_c_335_n 0.0115306f $X=2.14 $Y=0.43 $X2=0 $Y2=0
cc_180 Y N_VGND_c_335_n 0.0174675f $X=2.16 $Y=0.925 $X2=0 $Y2=0
