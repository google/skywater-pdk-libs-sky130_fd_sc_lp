* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__bufbuf_16 A VGND VNB VPB VPWR X
X0 X a_610_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR a_610_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR a_610_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND a_27_49# a_196_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_610_47# a_196_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_27_49# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_610_47# a_196_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VPWR a_27_49# a_196_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND a_196_49# a_610_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VGND a_610_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 X a_610_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 X a_610_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VPWR a_610_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 X a_610_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VPWR a_610_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR a_610_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 X a_610_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VGND a_610_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 VPWR a_610_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 X a_610_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_610_47# a_196_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 X a_610_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 X a_610_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_27_49# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VPWR a_196_49# a_610_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VGND a_610_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 X a_610_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_196_49# a_27_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VPWR a_27_49# a_196_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_610_47# a_196_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 VGND a_610_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 X a_610_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 VPWR a_610_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 X a_610_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 X a_610_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 VGND a_196_49# a_610_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X36 X a_610_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X37 a_610_47# a_196_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 VGND a_610_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 VPWR a_196_49# a_610_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X40 VGND a_610_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X41 VGND a_610_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X42 X a_610_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X43 X a_610_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X44 VGND a_27_49# a_196_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X45 a_610_47# a_196_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X46 a_196_49# a_27_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X47 VPWR a_196_49# a_610_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X48 VPWR a_610_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X49 VGND a_610_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X50 VGND a_196_49# a_610_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X51 X a_610_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
