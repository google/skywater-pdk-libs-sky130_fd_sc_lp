* File: sky130_fd_sc_lp__dlclkp_2.pex.spice
* Created: Fri Aug 28 10:25:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%A_78_269# 1 2 9 13 15 18 19 21 22 24 27 30
+ 31 35 39
c105 35 0 1.79399e-19 $X=1.155 $Y=1.645
c106 31 0 1.62138e-19 $X=0.555 $Y=1.51
r107 36 39 9.60369 $w=2.38e-07 $l=2e-07 $layer=LI1_cond $X=1.59 $Y=0.725
+ $X2=1.79 $Y2=0.725
r108 31 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.51
+ $X2=0.555 $Y2=1.675
r109 31 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.51
+ $X2=0.555 $Y2=1.345
r110 30 33 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.59 $Y=1.51
+ $X2=0.59 $Y2=1.645
r111 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.555
+ $Y=1.51 $X2=0.555 $Y2=1.51
r112 25 27 4.93904 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=1.685 $Y=2.45
+ $X2=1.685 $Y2=2.57
r113 23 36 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.59 $Y=0.845
+ $X2=1.59 $Y2=0.725
r114 23 24 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.59 $Y=0.845
+ $X2=1.59 $Y2=1.56
r115 21 25 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.545 $Y=2.365
+ $X2=1.685 $Y2=2.45
r116 21 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.545 $Y=2.365
+ $X2=1.24 $Y2=2.365
r117 20 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=1.645
+ $X2=1.155 $Y2=1.645
r118 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.505 $Y=1.645
+ $X2=1.59 $Y2=1.56
r119 19 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.505 $Y=1.645
+ $X2=1.24 $Y2=1.645
r120 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.155 $Y=2.28
+ $X2=1.24 $Y2=2.365
r121 17 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=1.73
+ $X2=1.155 $Y2=1.645
r122 17 18 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.155 $Y=1.73
+ $X2=1.155 $Y2=2.28
r123 16 33 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.645
+ $X2=0.59 $Y2=1.645
r124 15 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=1.645
+ $X2=1.155 $Y2=1.645
r125 15 16 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=1.645
+ $X2=0.72 $Y2=1.645
r126 13 42 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.525 $Y=0.655
+ $X2=0.525 $Y2=1.345
r127 9 43 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.51 $Y=2.465
+ $X2=0.51 $Y2=1.675
r128 2 27 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=2.325 $X2=1.71 $Y2=2.57
r129 1 39 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=0.405 $X2=1.79 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%GATE 3 7 9 12
c52 12 0 4.99354e-20 $X=1.125 $Y=1.295
c53 9 0 1.62138e-19 $X=1.2 $Y=1.295
c54 3 0 1.75443e-19 $X=1.135 $Y=2.645
r55 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.125 $Y=1.295
+ $X2=1.125 $Y2=1.46
r56 12 14 54.0802 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.125 $Y=1.295
+ $X2=1.125 $Y2=1.085
r57 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.125
+ $Y=1.295 $X2=1.125 $Y2=1.295
r58 7 14 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.215 $Y=0.615 $X2=1.215
+ $Y2=1.085
r59 3 15 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=1.135 $Y=2.645
+ $X2=1.135 $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%A_284_367# 1 2 9 13 14 17 20 23 25 28 32 33
+ 35 39 42 43 48
c120 32 0 1.03708e-19 $X=2.025 $Y=1.1
c121 14 0 1.61721e-19 $X=1.855 $Y=2.005
c122 9 0 6.18699e-20 $X=1.495 $Y=2.645
r123 41 43 8.37256 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=2.052
+ $X2=3.4 $Y2=2.052
r124 41 42 8.59491 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=2.052
+ $X2=3.07 $Y2=2.052
r125 37 39 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=0.59
+ $X2=3.4 $Y2=0.59
r126 33 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.025 $Y=1.1
+ $X2=2.025 $Y2=0.935
r127 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.025
+ $Y=1.1 $X2=2.025 $Y2=1.1
r128 29 32 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=1.14
+ $X2=2.025 $Y2=1.14
r129 27 28 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.62 $Y=0.695
+ $X2=4.62 $Y2=1.985
r130 25 28 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.535 $Y=2.08
+ $X2=4.62 $Y2=1.985
r131 25 43 66.2536 $w=1.88e-07 $l=1.135e-06 $layer=LI1_cond $X=4.535 $Y=2.08
+ $X2=3.4 $Y2=2.08
r132 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.535 $Y=0.61
+ $X2=4.62 $Y2=0.695
r133 23 39 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=4.535 $Y=0.61
+ $X2=3.4 $Y2=0.61
r134 22 35 4.60183 $w=1.95e-07 $l=9.21954e-08 $layer=LI1_cond $X=2.025 $Y=2.02
+ $X2=1.94 $Y2=2.005
r135 22 42 64.3889 $w=1.78e-07 $l=1.045e-06 $layer=LI1_cond $X=2.025 $Y=2.02
+ $X2=3.07 $Y2=2.02
r136 20 35 1.84097 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.94 $Y=1.9
+ $X2=1.94 $Y2=2.005
r137 19 29 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.94 $Y=1.265
+ $X2=1.94 $Y2=1.14
r138 19 20 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.94 $Y=1.265
+ $X2=1.94 $Y2=1.9
r139 17 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=2
+ $X2=1.585 $Y2=2.165
r140 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=2 $X2=1.585 $Y2=2
r141 14 35 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=2.005
+ $X2=1.94 $Y2=2.005
r142 14 16 14.2597 $w=2.08e-07 $l=2.7e-07 $layer=LI1_cond $X=1.855 $Y=2.005
+ $X2=1.585 $Y2=2.005
r143 13 48 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.005 $Y=0.615
+ $X2=2.005 $Y2=0.935
r144 9 46 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.495 $Y=2.645
+ $X2=1.495 $Y2=2.165
r145 2 41 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=1.955 $X2=3.235 $Y2=2.08
r146 1 37 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.095
+ $Y=0.405 $X2=3.235 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%A_300_55# 1 2 9 11 12 15 19 22 25 27 28 29
+ 30 33 38 39 40 41 46
c112 41 0 3.33623e-19 $X=3.235 $Y=0.97
c113 12 0 1.61721e-19 $X=1.65 $Y=1.55
c114 11 0 1.03708e-19 $X=1.96 $Y=1.55
r115 44 46 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=4.2 $Y=1.065
+ $X2=4.2 $Y2=1.73
r116 41 43 43.488 $w=1.88e-07 $l=7.45e-07 $layer=LI1_cond $X=3.235 $Y=0.97
+ $X2=3.98 $Y2=0.97
r117 40 44 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=4.035 $Y=0.97
+ $X2=4.2 $Y2=1.065
r118 40 43 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=4.035 $Y=0.97
+ $X2=3.98 $Y2=0.97
r119 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.11
+ $Y=1.1 $X2=3.11 $Y2=1.1
r120 36 38 19.8052 $w=2.08e-07 $l=3.75e-07 $layer=LI1_cond $X=3.13 $Y=1.475
+ $X2=3.13 $Y2=1.1
r121 35 41 6.83868 $w=1.9e-07 $l=1.44914e-07 $layer=LI1_cond $X=3.13 $Y=1.065
+ $X2=3.235 $Y2=0.97
r122 35 38 1.84848 $w=2.08e-07 $l=3.5e-08 $layer=LI1_cond $X=3.13 $Y=1.065
+ $X2=3.13 $Y2=1.1
r123 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=1.64 $X2=2.37 $Y2=1.64
r124 30 36 7.02201 $w=2.85e-07 $l=1.87281e-07 $layer=LI1_cond $X=3.025 $Y=1.617
+ $X2=3.13 $Y2=1.475
r125 30 32 26.486 $w=2.83e-07 $l=6.55e-07 $layer=LI1_cond $X=3.025 $Y=1.617
+ $X2=2.37 $Y2=1.617
r126 28 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.11 $Y=1.44
+ $X2=3.11 $Y2=1.1
r127 28 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.44
+ $X2=3.11 $Y2=1.605
r128 27 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=0.935
+ $X2=3.11 $Y2=1.1
r129 24 33 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=2.11 $Y=1.64
+ $X2=2.37 $Y2=1.64
r130 24 25 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=2.11 $Y=1.64
+ $X2=2.035 $Y2=1.64
r131 22 29 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=3.02 $Y=2.275
+ $X2=3.02 $Y2=1.605
r132 19 27 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.02 $Y=0.615
+ $X2=3.02 $Y2=0.935
r133 13 25 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.035 $Y=1.805
+ $X2=2.035 $Y2=1.64
r134 13 15 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.035 $Y=1.805
+ $X2=2.035 $Y2=2.535
r135 11 25 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.96 $Y=1.55
+ $X2=2.035 $Y2=1.64
r136 11 12 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.96 $Y=1.55
+ $X2=1.65 $Y2=1.55
r137 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.575 $Y=1.475
+ $X2=1.65 $Y2=1.55
r138 7 9 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.575 $Y=1.475
+ $X2=1.575 $Y2=0.615
r139 2 46 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.605 $X2=4.2 $Y2=1.73
r140 1 43 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.665 $X2=3.98 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%A_33_47# 1 2 9 13 14 15 18 22 26 31 32 34
+ 37 38 39 40 43 44 45 47 50 51 53 56 57 59 60 62 68 69 72 79 80 82 84
c230 84 0 1.90112e-19 $X=2.565 $Y=0.935
c231 80 0 1.43511e-19 $X=2.565 $Y=1.1
c232 62 0 4.99354e-20 $X=0.287 $Y=0.75
c233 45 0 6.18699e-20 $X=2.165 $Y=2.43
c234 40 0 1.75443e-19 $X=1.995 $Y=2.99
r235 80 84 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.565 $Y=1.1
+ $X2=2.565 $Y2=0.935
r236 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.565
+ $Y=1.1 $X2=2.565 $Y2=1.1
r237 76 79 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.445 $Y=1.1
+ $X2=2.565 $Y2=1.1
r238 72 74 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.235 $Y=2.715
+ $X2=1.235 $Y2=2.99
r239 68 69 6.43819 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=0.29 $Y=2.015
+ $X2=0.29 $Y2=1.91
r240 66 69 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=0.205 $Y=1.095
+ $X2=0.205 $Y2=1.91
r241 65 66 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.287 $Y=0.93
+ $X2=0.287 $Y2=1.095
r242 62 65 6.19223 $w=3.33e-07 $l=1.8e-07 $layer=LI1_cond $X=0.287 $Y=0.75
+ $X2=0.287 $Y2=0.93
r243 62 63 3.21382 $w=3.33e-07 $l=8.5e-08 $layer=LI1_cond $X=0.287 $Y=0.75
+ $X2=0.287 $Y2=0.665
r244 60 92 11.9307 $w=3.03e-07 $l=7.5e-08 $layer=POLY_cond $X=5.57 $Y=1.41
+ $X2=5.645 $Y2=1.41
r245 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.57
+ $Y=1.44 $X2=5.57 $Y2=1.44
r246 57 59 30.6459 $w=1.88e-07 $l=5.25e-07 $layer=LI1_cond $X=5.045 $Y=1.44
+ $X2=5.57 $Y2=1.44
r247 55 57 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.96 $Y=1.535
+ $X2=5.045 $Y2=1.44
r248 55 56 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=4.96 $Y=1.535
+ $X2=4.96 $Y2=2.345
r249 54 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=2.43
+ $X2=3.5 $Y2=2.43
r250 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.875 $Y=2.43
+ $X2=4.96 $Y2=2.345
r251 53 54 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=4.875 $Y=2.43
+ $X2=3.665 $Y2=2.43
r252 51 88 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.5 $Y=2.94 $X2=3.5
+ $Y2=3.055
r253 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.5
+ $Y=2.94 $X2=3.5 $Y2=2.94
r254 48 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=2.515 $X2=3.5
+ $Y2=2.43
r255 48 50 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=3.5 $Y=2.515
+ $X2=3.5 $Y2=2.94
r256 47 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0.935
+ $X2=2.445 $Y2=1.1
r257 46 47 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.445 $Y=0.435
+ $X2=2.445 $Y2=0.935
r258 44 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=2.43
+ $X2=3.5 $Y2=2.43
r259 44 45 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=3.335 $Y=2.43
+ $X2=2.165 $Y2=2.43
r260 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.08 $Y=2.515
+ $X2=2.165 $Y2=2.43
r261 42 43 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.08 $Y=2.515
+ $X2=2.08 $Y2=2.905
r262 41 74 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=2.99
+ $X2=1.235 $Y2=2.99
r263 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.995 $Y=2.99
+ $X2=2.08 $Y2=2.905
r264 40 41 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.995 $Y=2.99
+ $X2=1.32 $Y2=2.99
r265 38 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=0.35
+ $X2=2.445 $Y2=0.435
r266 38 39 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.36 $Y=0.35
+ $X2=1.255 $Y2=0.35
r267 36 39 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.165 $Y=0.435
+ $X2=1.255 $Y2=0.35
r268 36 37 14.1717 $w=1.78e-07 $l=2.3e-07 $layer=LI1_cond $X=1.165 $Y=0.435
+ $X2=1.165 $Y2=0.665
r269 35 71 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.46 $Y=2.715
+ $X2=0.29 $Y2=2.715
r270 34 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=2.715
+ $X2=1.235 $Y2=2.715
r271 34 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.15 $Y=2.715
+ $X2=0.46 $Y2=2.715
r272 33 62 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.455 $Y=0.75
+ $X2=0.287 $Y2=0.75
r273 32 37 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.075 $Y=0.75
+ $X2=1.165 $Y2=0.665
r274 32 33 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.075 $Y=0.75
+ $X2=0.455 $Y2=0.75
r275 31 71 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.29 $Y=2.63
+ $X2=0.29 $Y2=2.715
r276 30 68 2.2032 $w=3.38e-07 $l=6.5e-08 $layer=LI1_cond $X=0.29 $Y=2.08
+ $X2=0.29 $Y2=2.015
r277 30 31 18.6425 $w=3.38e-07 $l=5.5e-07 $layer=LI1_cond $X=0.29 $Y=2.08
+ $X2=0.29 $Y2=2.63
r278 26 63 9.90697 $w=2.83e-07 $l=2.45e-07 $layer=LI1_cond $X=0.262 $Y=0.42
+ $X2=0.262 $Y2=0.665
r279 20 92 19.2026 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=5.645 $Y=1.605
+ $X2=5.645 $Y2=1.41
r280 20 22 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.645 $Y=1.605
+ $X2=5.645 $Y2=2.155
r281 16 60 43.7459 $w=3.03e-07 $l=3.59514e-07 $layer=POLY_cond $X=5.295 $Y=1.215
+ $X2=5.57 $Y2=1.41
r282 16 18 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.295 $Y=1.215
+ $X2=5.295 $Y2=0.875
r283 14 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.335 $Y=3.055
+ $X2=3.5 $Y2=3.055
r284 14 15 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=3.335 $Y=3.055
+ $X2=2.47 $Y2=3.055
r285 13 84 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.475 $Y=0.615
+ $X2=2.475 $Y2=0.935
r286 7 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.395 $Y=2.98
+ $X2=2.47 $Y2=3.055
r287 7 9 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.395 $Y=2.98
+ $X2=2.395 $Y2=2.535
r288 2 71 400 $w=1.7e-07 $l=9.2038e-07 $layer=licon1_PDIFF $count=1 $X=0.17
+ $Y=1.835 $X2=0.295 $Y2=2.695
r289 2 68 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.17
+ $Y=1.835 $X2=0.295 $Y2=2.015
r290 1 65 182 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.93
r291 1 26 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%CLK 1 5 7 9 12 14 16 19 21 23 27
c63 14 0 1.82504e-19 $X=5.12 $Y=1.725
r64 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.68
+ $Y=1.545 $X2=3.68 $Y2=1.545
r65 23 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.68 $Y=1.455 $X2=3.68
+ $Y2=1.545
r66 21 27 3.373 $w=4.08e-07 $l=1.2e-07 $layer=LI1_cond $X=3.64 $Y=1.665 $X2=3.64
+ $Y2=1.545
r67 18 19 74.5076 $w=2.62e-07 $l=4.05e-07 $layer=POLY_cond $X=4.53 $Y=1.552
+ $X2=4.935 $Y2=1.552
r68 14 19 34.0344 $w=2.62e-07 $l=2.57352e-07 $layer=POLY_cond $X=5.12 $Y=1.725
+ $X2=4.935 $Y2=1.552
r69 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.12 $Y=1.725
+ $X2=5.12 $Y2=2.155
r70 10 19 15.8058 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=4.935 $Y=1.38
+ $X2=4.935 $Y2=1.552
r71 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.935 $Y=1.38
+ $X2=4.935 $Y2=0.875
r72 7 18 15.8058 $w=1.5e-07 $l=1.73e-07 $layer=POLY_cond $X=4.53 $Y=1.725
+ $X2=4.53 $Y2=1.552
r73 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.53 $Y=1.725 $X2=4.53
+ $Y2=2.155
r74 3 18 40.4733 $w=2.62e-07 $l=2.93666e-07 $layer=POLY_cond $X=4.31 $Y=1.38
+ $X2=4.53 $Y2=1.552
r75 3 5 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.31 $Y=1.38 $X2=4.31
+ $Y2=0.875
r76 2 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.455
+ $X2=3.68 $Y2=1.455
r77 1 3 22.5321 $w=2.62e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.235 $Y=1.455
+ $X2=4.31 $Y2=1.38
r78 1 2 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.235 $Y=1.455
+ $X2=3.845 $Y2=1.455
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%A_1039_367# 1 2 9 13 15 19 23 25 28 30 31
+ 32 37 40 44
c75 28 0 1.82504e-19 $X=5.385 $Y=1.98
r76 44 45 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=6.132 $Y=1.42
+ $X2=6.132 $Y2=1.345
r77 40 42 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=5.51 $Y=0.875
+ $X2=5.51 $Y2=1.09
r78 38 47 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.132 $Y=1.51
+ $X2=6.132 $Y2=1.675
r79 38 44 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=6.132 $Y=1.51
+ $X2=6.132 $Y2=1.42
r80 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.11
+ $Y=1.51 $X2=6.11 $Y2=1.51
r81 35 37 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=6.07 $Y=1.705
+ $X2=6.07 $Y2=1.51
r82 34 37 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.07 $Y=1.175
+ $X2=6.07 $Y2=1.51
r83 33 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.675 $Y=1.09
+ $X2=5.51 $Y2=1.09
r84 32 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.945 $Y=1.09
+ $X2=6.07 $Y2=1.175
r85 32 33 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.945 $Y=1.09
+ $X2=5.675 $Y2=1.09
r86 30 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.945 $Y=1.79
+ $X2=6.07 $Y2=1.705
r87 30 31 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.945 $Y=1.79
+ $X2=5.55 $Y2=1.79
r88 26 31 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=5.382 $Y=1.875
+ $X2=5.55 $Y2=1.79
r89 26 28 3.61213 $w=3.33e-07 $l=1.05e-07 $layer=LI1_cond $X=5.382 $Y=1.875
+ $X2=5.382 $Y2=1.98
r90 21 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.675 $Y=1.495
+ $X2=6.675 $Y2=1.42
r91 21 23 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=6.675 $Y=1.495
+ $X2=6.675 $Y2=2.465
r92 17 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.675 $Y=1.345
+ $X2=6.675 $Y2=1.42
r93 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.675 $Y=1.345
+ $X2=6.675 $Y2=0.655
r94 16 44 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=6.32 $Y=1.42
+ $X2=6.132 $Y2=1.42
r95 15 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.6 $Y=1.42
+ $X2=6.675 $Y2=1.42
r96 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.6 $Y=1.42 $X2=6.32
+ $Y2=1.42
r97 13 47 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.245 $Y=2.465
+ $X2=6.245 $Y2=1.675
r98 9 45 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.245 $Y=0.655
+ $X2=6.245 $Y2=1.345
r99 2 28 300 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=2 $X=5.195
+ $Y=1.835 $X2=5.385 $Y2=1.98
r100 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.37
+ $Y=0.665 $X2=5.51 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%VPWR 1 2 3 4 5 20 24 28 32 34 39 40 41 43
+ 55 59 65 68 72 75 79
r86 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r87 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r88 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r90 65 68 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.805 $Y=3.065
+ $X2=0.805 $Y2=3.33
r91 63 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r92 63 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r93 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r94 60 75 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=5.985 $Y2=3.33
r95 60 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=6.48 $Y2=3.33
r96 59 78 4.14267 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=6.785 $Y=3.33
+ $X2=6.992 $Y2=3.33
r97 59 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.785 $Y=3.33
+ $X2=6.48 $Y2=3.33
r98 58 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r99 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r100 55 75 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.775 $Y=3.33
+ $X2=5.985 $Y2=3.33
r101 55 57 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.775 $Y=3.33
+ $X2=5.52 $Y2=3.33
r102 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r103 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r104 51 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 50 53 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r106 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r107 48 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=2.725 $Y2=3.33
r108 48 50 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=3.12 $Y2=3.33
r109 47 73 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 47 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r112 44 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.805 $Y2=3.33
r113 44 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.2 $Y2=3.33
r114 43 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=2.725 $Y2=3.33
r115 43 46 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r116 41 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r117 41 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r118 39 53 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.66 $Y=3.33 $X2=4.56
+ $Y2=3.33
r119 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=3.33
+ $X2=4.825 $Y2=3.33
r120 38 57 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.99 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.99 $Y=3.33
+ $X2=4.825 $Y2=3.33
r122 34 37 41.4026 $w=2.68e-07 $l=9.7e-07 $layer=LI1_cond $X=6.92 $Y=1.98
+ $X2=6.92 $Y2=2.95
r123 32 78 3.14202 $w=2.7e-07 $l=1.15521e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.992 $Y2=3.33
r124 32 37 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=2.95
r125 28 31 11.25 $w=4.18e-07 $l=4.1e-07 $layer=LI1_cond $X=5.985 $Y=2.13
+ $X2=5.985 $Y2=2.54
r126 26 75 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=3.33
r127 26 31 19.3446 $w=4.18e-07 $l=7.05e-07 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=2.54
r128 22 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.825 $Y=3.245
+ $X2=4.825 $Y2=3.33
r129 22 24 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.825 $Y=3.245
+ $X2=4.825 $Y2=2.78
r130 18 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=3.33
r131 18 20 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=2.78
r132 5 37 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.75
+ $Y=1.835 $X2=6.89 $Y2=2.95
r133 5 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.75
+ $Y=1.835 $X2=6.89 $Y2=1.98
r134 4 31 300 $w=1.7e-07 $l=8.45917e-07 $layer=licon1_PDIFF $count=2 $X=5.72
+ $Y=1.835 $X2=6.03 $Y2=2.54
r135 4 28 600 $w=1.7e-07 $l=3.89776e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.835 $X2=5.94 $Y2=2.13
r136 3 24 600 $w=1.7e-07 $l=1.04925e-06 $layer=licon1_PDIFF $count=1 $X=4.605
+ $Y=1.835 $X2=4.825 $Y2=2.78
r137 2 20 600 $w=1.7e-07 $l=5.68375e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=2.325 $X2=2.725 $Y2=2.78
r138 1 65 600 $w=1.7e-07 $l=1.33548e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.835 $X2=0.805 $Y2=3.065
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%GCLK 1 2 7 8 9 10 11 12 13 22
r18 13 40 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=6.477 $Y=2.775
+ $X2=6.477 $Y2=2.91
r19 12 13 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=6.477 $Y=2.405
+ $X2=6.477 $Y2=2.775
r20 11 12 21.7684 $w=2.23e-07 $l=4.25e-07 $layer=LI1_cond $X=6.477 $Y=1.98
+ $X2=6.477 $Y2=2.405
r21 10 11 16.1342 $w=2.23e-07 $l=3.15e-07 $layer=LI1_cond $X=6.477 $Y=1.665
+ $X2=6.477 $Y2=1.98
r22 9 10 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=6.477 $Y=1.295
+ $X2=6.477 $Y2=1.665
r23 8 9 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=6.477 $Y=0.925
+ $X2=6.477 $Y2=1.295
r24 7 8 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=6.477 $Y=0.555
+ $X2=6.477 $Y2=0.925
r25 7 22 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=6.477 $Y=0.555
+ $X2=6.477 $Y2=0.42
r26 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.91
r27 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=1.98
r28 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.32
+ $Y=0.235 $X2=6.46 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_2%VGND 1 2 3 4 5 18 22 26 28 30 33 34 35 37
+ 49 56 61 67 71 77 81
r80 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r81 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r82 71 74 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=4.605 $Y=0 $X2=4.605
+ $Y2=0.26
r83 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r84 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r85 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r86 65 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r87 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r88 62 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6.03
+ $Y2=0
r89 62 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6.48
+ $Y2=0
r90 61 80 4.352 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=6.76 $Y=0 $X2=6.98
+ $Y2=0
r91 61 64 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.76 $Y=0 $X2=6.48
+ $Y2=0
r92 60 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r93 60 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r94 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r95 57 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.77 $Y=0 $X2=4.605
+ $Y2=0
r96 57 59 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=4.77 $Y=0 $X2=5.52
+ $Y2=0
r97 56 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=6.03
+ $Y2=0
r98 56 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.865 $Y=0 $X2=5.52
+ $Y2=0
r99 55 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r100 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r101 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r102 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r103 49 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.605
+ $Y2=0
r104 49 54 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.44 $Y=0 $X2=4.08
+ $Y2=0
r105 48 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r106 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r107 45 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r108 45 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r109 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r110 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r111 42 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.74
+ $Y2=0
r112 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.2
+ $Y2=0
r113 40 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r114 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r115 37 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.74
+ $Y2=0
r116 37 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0
+ $X2=0.24 $Y2=0
r117 35 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r118 35 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r119 33 47 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.64
+ $Y2=0
r120 33 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.795
+ $Y2=0
r121 32 51 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.12
+ $Y2=0
r122 32 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.795
+ $Y2=0
r123 28 80 3.12553 $w=2.95e-07 $l=1.15888e-07 $layer=LI1_cond $X=6.907 $Y=0.085
+ $X2=6.98 $Y2=0
r124 28 30 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=6.907 $Y=0.085
+ $X2=6.907 $Y2=0.38
r125 24 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0
r126 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.03 $Y=0.085
+ $X2=6.03 $Y2=0.38
r127 20 34 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0
r128 20 22 30.0622 $w=1.88e-07 $l=5.15e-07 $layer=LI1_cond $X=2.795 $Y=0.085
+ $X2=2.795 $Y2=0.6
r129 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r130 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.39
r131 5 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.75
+ $Y=0.235 $X2=6.89 $Y2=0.38
r132 4 26 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.905
+ $Y=0.235 $X2=6.03 $Y2=0.38
r133 3 74 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.665 $X2=4.605 $Y2=0.26
r134 2 22 182 $w=1.7e-07 $l=3.17884e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.405 $X2=2.785 $Y2=0.6
r135 1 18 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.39
.ends

