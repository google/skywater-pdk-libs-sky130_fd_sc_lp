* NGSPICE file created from sky130_fd_sc_lp__a221oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_27_367# B1 a_303_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3734e+12p pd=1.226e+07u as=1.7766e+12p ps=1.542e+07u
M1001 Y A1 a_760_47# VNB nshort w=840000u l=150000u
+  ad=7.056e+11p pd=6.72e+06u as=4.704e+11p ps=4.48e+06u
M1002 a_384_47# B1 Y VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1003 Y C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.386e+12p ps=1.002e+07u
M1004 a_384_47# B2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_367# C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1006 a_303_367# B1 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_760_47# A1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_303_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=8.442e+11p pd=6.38e+06u as=0p ps=0u
M1010 VGND B2 a_384_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_760_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A2 a_303_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y B1 a_384_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_303_367# B2 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A2 a_760_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_303_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_367# B2 a_303_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y C1 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_303_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

