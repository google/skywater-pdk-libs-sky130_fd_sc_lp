* File: sky130_fd_sc_lp__or4_1.pxi.spice
* Created: Wed Sep  2 10:31:49 2020
* 
x_PM_SKY130_FD_SC_LP__OR4_1%D N_D_M1003_g N_D_M1006_g D D D N_D_c_67_n
+ PM_SKY130_FD_SC_LP__OR4_1%D
x_PM_SKY130_FD_SC_LP__OR4_1%C N_C_M1004_g N_C_M1001_g N_C_c_99_n N_C_c_100_n C C
+ N_C_c_101_n N_C_c_102_n PM_SKY130_FD_SC_LP__OR4_1%C
x_PM_SKY130_FD_SC_LP__OR4_1%B N_B_M1005_g N_B_c_137_n N_B_M1000_g B B
+ N_B_c_139_n N_B_c_140_n PM_SKY130_FD_SC_LP__OR4_1%B
x_PM_SKY130_FD_SC_LP__OR4_1%A N_A_c_184_n N_A_M1008_g N_A_c_185_n N_A_c_186_n
+ N_A_c_187_n N_A_M1002_g A N_A_c_183_n N_A_c_189_n PM_SKY130_FD_SC_LP__OR4_1%A
x_PM_SKY130_FD_SC_LP__OR4_1%A_40_480# N_A_40_480#_M1003_d N_A_40_480#_M1000_d
+ N_A_40_480#_M1006_s N_A_40_480#_c_237_n N_A_40_480#_M1009_g
+ N_A_40_480#_M1007_g N_A_40_480#_c_248_n N_A_40_480#_c_249_n
+ N_A_40_480#_c_336_p N_A_40_480#_c_239_n N_A_40_480#_c_240_n
+ N_A_40_480#_c_284_n N_A_40_480#_c_241_n N_A_40_480#_c_242_n
+ N_A_40_480#_c_243_n N_A_40_480#_c_250_n N_A_40_480#_c_244_n
+ N_A_40_480#_c_245_n N_A_40_480#_c_252_n N_A_40_480#_c_253_n
+ N_A_40_480#_c_246_n PM_SKY130_FD_SC_LP__OR4_1%A_40_480#
x_PM_SKY130_FD_SC_LP__OR4_1%VPWR N_VPWR_M1008_d VPWR N_VPWR_c_343_n
+ N_VPWR_c_344_n N_VPWR_c_345_n N_VPWR_c_342_n PM_SKY130_FD_SC_LP__OR4_1%VPWR
x_PM_SKY130_FD_SC_LP__OR4_1%X N_X_M1009_d N_X_M1007_d X X X X X X X X
+ N_X_c_371_n PM_SKY130_FD_SC_LP__OR4_1%X
x_PM_SKY130_FD_SC_LP__OR4_1%VGND N_VGND_M1003_s N_VGND_M1001_d N_VGND_M1002_d
+ N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n N_VGND_c_390_n N_VGND_c_391_n
+ VGND N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n N_VGND_c_395_n
+ PM_SKY130_FD_SC_LP__OR4_1%VGND
cc_1 VNB N_D_M1003_g 0.0268967f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.445
cc_2 VNB N_D_M1006_g 0.00682453f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.61
cc_3 VNB D 0.0371684f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_4 VNB N_D_c_67_n 0.084293f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_5 VNB N_C_M1004_g 0.00342898f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.445
cc_6 VNB N_C_M1001_g 0.0256893f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.61
cc_7 VNB N_C_c_99_n 0.0208936f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_C_c_100_n 0.0153087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C_c_101_n 0.0162259f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=0.84
cc_10 VNB N_C_c_102_n 0.0025276f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.51
cc_11 VNB N_B_c_137_n 0.0351868f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.61
cc_12 VNB N_B_M1000_g 0.03216f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_13 VNB N_B_c_139_n 0.0247549f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_14 VNB N_B_c_140_n 0.00233251f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_15 VNB N_A_M1002_g 0.0459397f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_A_c_183_n 0.0270587f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.005
cc_17 VNB N_A_40_480#_c_237_n 0.0202184f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_A_40_480#_M1007_g 0.00792626f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.005
cc_19 VNB N_A_40_480#_c_239_n 0.0130494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_40_480#_c_240_n 0.00399566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_40_480#_c_241_n 0.00221475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_40_480#_c_242_n 0.0149952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_40_480#_c_243_n 0.00361616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_40_480#_c_244_n 9.79898e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_40_480#_c_245_n 0.00450934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_40_480#_c_246_n 0.041599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_342_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB X 0.0400938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_371_n 0.0354295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_387_n 0.012093f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_31 VNB N_VGND_c_388_n 0.0191613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_389_n 0.00622594f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_33 VNB N_VGND_c_390_n 0.0154881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_391_n 0.00470919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_392_n 0.0230408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_393_n 0.189726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_394_n 0.0139508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_395_n 0.0122121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_D_M1006_g 0.059094f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.61
cc_40 VPB D 0.0145027f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_41 VPB N_C_M1004_g 0.0423944f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.445
cc_42 VPB N_C_c_102_n 0.00485806f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.51
cc_43 VPB N_B_M1005_g 0.0327641f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.445
cc_44 VPB N_B_c_137_n 0.0392273f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.61
cc_45 VPB N_B_c_140_n 0.0031443f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_46 VPB N_A_c_184_n 0.0204154f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.84
cc_47 VPB N_A_c_185_n 0.0291097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_c_186_n 0.00707373f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.51
cc_49 VPB N_A_c_187_n 0.0317758f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.61
cc_50 VPB N_A_c_183_n 0.00666538f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.005
cc_51 VPB N_A_c_189_n 0.00237127f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_52 VPB N_A_40_480#_M1007_g 0.0259084f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.005
cc_53 VPB N_A_40_480#_c_248_n 0.020798f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.51
cc_54 VPB N_A_40_480#_c_249_n 0.0144455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_40_480#_c_250_n 0.0113875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_40_480#_c_244_n 0.00206767f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_40_480#_c_252_n 0.038131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_40_480#_c_253_n 0.0052352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_343_n 0.0535747f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.61
cc_60 VPB N_VPWR_c_344_n 0.0443772f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_61 VPB N_VPWR_c_345_n 0.0152759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_342_n 0.0856816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB X 0.0571021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 N_D_M1003_g N_C_M1001_g 0.0153358f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_65 D N_C_M1001_g 2.74829e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_66 N_D_c_67_n N_C_M1001_g 0.00372919f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_67 N_D_M1006_g N_C_c_100_n 0.0657384f $X=0.54 $Y=2.61 $X2=0 $Y2=0
cc_68 D N_C_c_101_n 6.91353e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_69 N_D_c_67_n N_C_c_101_n 0.0657384f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_70 N_D_M1006_g N_C_c_102_n 0.00685638f $X=0.54 $Y=2.61 $X2=0 $Y2=0
cc_71 D N_C_c_102_n 0.0658523f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_72 N_D_c_67_n N_C_c_102_n 0.0146797f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_73 N_D_M1006_g N_A_40_480#_c_248_n 0.0123831f $X=0.54 $Y=2.61 $X2=0 $Y2=0
cc_74 N_D_M1006_g N_A_40_480#_c_249_n 0.00716284f $X=0.54 $Y=2.61 $X2=0 $Y2=0
cc_75 D N_A_40_480#_c_249_n 0.0233305f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_76 N_D_c_67_n N_A_40_480#_c_249_n 0.00291471f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_77 N_D_M1003_g N_A_40_480#_c_240_n 0.00449694f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_78 D N_A_40_480#_c_240_n 0.00285604f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_79 N_D_c_67_n N_A_40_480#_c_240_n 4.82886e-19 $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_80 N_D_M1006_g N_A_40_480#_c_252_n 0.015901f $X=0.54 $Y=2.61 $X2=0 $Y2=0
cc_81 N_D_M1006_g N_VPWR_c_343_n 0.00462485f $X=0.54 $Y=2.61 $X2=0 $Y2=0
cc_82 N_D_M1006_g N_VPWR_c_342_n 0.00502397f $X=0.54 $Y=2.61 $X2=0 $Y2=0
cc_83 N_D_M1003_g N_VGND_c_388_n 0.00369789f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_84 D N_VGND_c_388_n 0.0234756f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_85 N_D_c_67_n N_VGND_c_388_n 0.00176905f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_86 N_D_M1003_g N_VGND_c_393_n 0.0117894f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_87 D N_VGND_c_393_n 0.00297929f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_88 N_D_c_67_n N_VGND_c_393_n 5.23483e-19 $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_89 N_D_M1003_g N_VGND_c_394_n 0.00585385f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_90 N_D_M1003_g N_VGND_c_395_n 5.80076e-19 $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_91 N_C_M1004_g N_B_c_137_n 0.0804049f $X=0.9 $Y=2.61 $X2=0 $Y2=0
cc_92 N_C_c_99_n N_B_c_137_n 0.0177211f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_93 N_C_c_102_n N_B_c_137_n 0.00217131f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_94 N_C_M1001_g N_B_M1000_g 0.00771567f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_95 N_C_c_101_n N_B_M1000_g 0.00318479f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_96 N_C_c_101_n N_B_c_139_n 0.0177211f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_97 N_C_c_102_n N_B_c_139_n 0.00211076f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_98 N_C_M1004_g N_B_c_140_n 2.32959e-19 $X=0.9 $Y=2.61 $X2=0 $Y2=0
cc_99 N_C_c_101_n N_B_c_140_n 0.00189036f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_100 N_C_c_102_n N_B_c_140_n 0.0506018f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_101 N_C_M1004_g N_A_40_480#_c_248_n 0.00257991f $X=0.9 $Y=2.61 $X2=0 $Y2=0
cc_102 N_C_M1001_g N_A_40_480#_c_239_n 0.0125964f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_103 N_C_c_101_n N_A_40_480#_c_239_n 0.00516389f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_104 N_C_c_102_n N_A_40_480#_c_239_n 0.0261144f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_105 N_C_c_102_n N_A_40_480#_c_240_n 0.0201834f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_106 N_C_M1004_g N_A_40_480#_c_252_n 0.0173202f $X=0.9 $Y=2.61 $X2=0 $Y2=0
cc_107 N_C_c_100_n N_A_40_480#_c_252_n 7.26127e-19 $X=0.99 $Y=1.575 $X2=0 $Y2=0
cc_108 N_C_c_102_n N_A_40_480#_c_252_n 0.0478813f $X=0.99 $Y=1.07 $X2=0 $Y2=0
cc_109 N_C_M1004_g N_VPWR_c_343_n 0.00481372f $X=0.9 $Y=2.61 $X2=0 $Y2=0
cc_110 N_C_M1004_g N_VPWR_c_342_n 0.00502397f $X=0.9 $Y=2.61 $X2=0 $Y2=0
cc_111 N_C_M1001_g N_VGND_c_393_n 0.00422351f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_112 N_C_M1001_g N_VGND_c_394_n 0.00354752f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_113 N_C_M1001_g N_VGND_c_395_n 0.0078322f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_114 N_B_M1005_g N_A_c_186_n 0.0508449f $X=1.26 $Y=2.61 $X2=0 $Y2=0
cc_115 N_B_c_137_n N_A_c_186_n 0.00519856f $X=1.575 $Y=1.465 $X2=0 $Y2=0
cc_116 N_B_c_140_n N_A_c_186_n 7.33922e-19 $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_117 N_B_M1005_g N_A_c_187_n 0.00308937f $X=1.26 $Y=2.61 $X2=0 $Y2=0
cc_118 N_B_c_137_n N_A_c_187_n 0.00634885f $X=1.575 $Y=1.465 $X2=0 $Y2=0
cc_119 N_B_c_140_n N_A_c_187_n 0.00238698f $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_120 N_B_M1000_g N_A_M1002_g 0.0349349f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_121 N_B_c_140_n N_A_M1002_g 8.42914e-19 $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_122 N_B_c_137_n N_A_c_183_n 0.0210419f $X=1.575 $Y=1.465 $X2=0 $Y2=0
cc_123 N_B_c_140_n N_A_c_183_n 0.00141213f $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_124 N_B_c_137_n N_A_c_189_n 9.91218e-19 $X=1.575 $Y=1.465 $X2=0 $Y2=0
cc_125 N_B_c_140_n N_A_c_189_n 0.0209832f $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_126 N_B_M1000_g N_A_40_480#_c_239_n 0.0134722f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_127 N_B_c_139_n N_A_40_480#_c_239_n 0.00288398f $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_128 N_B_c_140_n N_A_40_480#_c_239_n 0.0272335f $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_129 N_B_M1000_g N_A_40_480#_c_241_n 0.00447228f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_130 N_B_c_140_n N_A_40_480#_c_241_n 0.00528059f $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_131 N_B_c_139_n N_A_40_480#_c_243_n 0.00130402f $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_132 N_B_c_140_n N_A_40_480#_c_243_n 0.0144378f $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_133 N_B_M1005_g N_A_40_480#_c_252_n 0.0230177f $X=1.26 $Y=2.61 $X2=0 $Y2=0
cc_134 N_B_c_137_n N_A_40_480#_c_252_n 0.00729108f $X=1.575 $Y=1.465 $X2=0 $Y2=0
cc_135 N_B_c_140_n N_A_40_480#_c_252_n 0.0323335f $X=1.56 $Y=1.17 $X2=0 $Y2=0
cc_136 N_B_M1005_g N_VPWR_c_343_n 0.00481372f $X=1.26 $Y=2.61 $X2=0 $Y2=0
cc_137 N_B_M1005_g N_VPWR_c_344_n 0.00250715f $X=1.26 $Y=2.61 $X2=0 $Y2=0
cc_138 N_B_M1005_g N_VPWR_c_342_n 0.00502397f $X=1.26 $Y=2.61 $X2=0 $Y2=0
cc_139 N_B_M1000_g N_VGND_c_390_n 0.00354752f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_140 N_B_M1000_g N_VGND_c_393_n 0.00427489f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_141 N_B_M1000_g N_VGND_c_395_n 0.00801045f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_M1002_g N_A_40_480#_c_237_n 0.0238321f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A_c_187_n N_A_40_480#_M1007_g 0.00722679f $X=2.07 $Y=2.145 $X2=0 $Y2=0
cc_144 N_A_c_183_n N_A_40_480#_M1007_g 0.00309564f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_145 N_A_c_189_n N_A_40_480#_M1007_g 3.80618e-19 $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_146 N_A_M1002_g N_A_40_480#_c_284_n 0.00411011f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_M1002_g N_A_40_480#_c_241_n 0.00601097f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A_M1002_g N_A_40_480#_c_242_n 0.0110897f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_c_183_n N_A_40_480#_c_242_n 0.00221896f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A_c_189_n N_A_40_480#_c_242_n 0.014647f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A_M1002_g N_A_40_480#_c_243_n 0.00222409f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_152 N_A_c_183_n N_A_40_480#_c_243_n 0.00270344f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_153 N_A_c_189_n N_A_40_480#_c_243_n 0.00952969f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_154 N_A_c_187_n N_A_40_480#_c_244_n 0.003469f $X=2.07 $Y=2.145 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_A_40_480#_c_244_n 5.99721e-19 $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_156 N_A_c_183_n N_A_40_480#_c_244_n 0.00225255f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A_c_189_n N_A_40_480#_c_244_n 0.0200465f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A_M1002_g N_A_40_480#_c_245_n 0.00391645f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_c_185_n N_A_40_480#_c_252_n 0.013891f $X=1.995 $Y=2.22 $X2=0 $Y2=0
cc_160 N_A_c_186_n N_A_40_480#_c_252_n 0.0104663f $X=1.695 $Y=2.22 $X2=0 $Y2=0
cc_161 N_A_c_187_n N_A_40_480#_c_252_n 0.0102866f $X=2.07 $Y=2.145 $X2=0 $Y2=0
cc_162 N_A_c_189_n N_A_40_480#_c_252_n 0.00963813f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_163 N_A_c_187_n N_A_40_480#_c_253_n 0.00255223f $X=2.07 $Y=2.145 $X2=0 $Y2=0
cc_164 N_A_c_183_n N_A_40_480#_c_253_n 9.39532e-19 $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A_c_189_n N_A_40_480#_c_253_n 0.0133149f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_166 N_A_M1002_g N_A_40_480#_c_246_n 0.00626879f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A_c_183_n N_A_40_480#_c_246_n 0.00949866f $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_168 N_A_c_189_n N_A_40_480#_c_246_n 3.42781e-19 $X=2.16 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A_c_184_n N_VPWR_c_343_n 0.00400048f $X=1.62 $Y=2.295 $X2=0 $Y2=0
cc_170 N_A_c_184_n N_VPWR_c_344_n 0.013872f $X=1.62 $Y=2.295 $X2=0 $Y2=0
cc_171 N_A_c_185_n N_VPWR_c_344_n 0.0102073f $X=1.995 $Y=2.22 $X2=0 $Y2=0
cc_172 N_A_c_184_n N_VPWR_c_342_n 0.00418664f $X=1.62 $Y=2.295 $X2=0 $Y2=0
cc_173 N_A_M1002_g N_VGND_c_389_n 0.00570283f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_174 N_A_M1002_g N_VGND_c_390_n 0.00542362f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_175 N_A_M1002_g N_VGND_c_393_n 0.0100279f $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_176 N_A_M1002_g N_VGND_c_395_n 5.42397e-19 $X=2.16 $Y=0.445 $X2=0 $Y2=0
cc_177 N_A_40_480#_c_250_n N_VPWR_M1008_d 0.00404168f $X=2.565 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A_40_480#_c_244_n N_VPWR_M1008_d 0.00174518f $X=2.73 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A_40_480#_c_248_n N_VPWR_c_343_n 0.00696076f $X=0.325 $Y=2.61 $X2=0
+ $Y2=0
cc_180 N_A_40_480#_M1007_g N_VPWR_c_344_n 0.017989f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_40_480#_c_250_n N_VPWR_c_344_n 0.0318616f $X=2.565 $Y=2.04 $X2=0
+ $Y2=0
cc_182 N_A_40_480#_c_252_n N_VPWR_c_344_n 0.0489829f $X=2.165 $Y=2.095 $X2=0
+ $Y2=0
cc_183 N_A_40_480#_M1007_g N_VPWR_c_345_n 0.00486043f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_40_480#_M1007_g N_VPWR_c_342_n 0.00913103f $X=2.885 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_A_40_480#_c_248_n N_VPWR_c_342_n 0.0105112f $X=0.325 $Y=2.61 $X2=0
+ $Y2=0
cc_186 N_A_40_480#_c_242_n N_X_M1009_d 9.95962e-19 $X=2.565 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A_40_480#_c_237_n X 0.00443379f $X=2.65 $Y=1.185 $X2=0 $Y2=0
cc_188 N_A_40_480#_c_242_n X 0.0134242f $X=2.565 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_40_480#_c_244_n X 0.0444127f $X=2.73 $Y=1.35 $X2=0 $Y2=0
cc_190 N_A_40_480#_c_246_n X 0.0193206f $X=2.885 $Y=1.35 $X2=0 $Y2=0
cc_191 N_A_40_480#_c_237_n N_X_c_371_n 0.00831149f $X=2.65 $Y=1.185 $X2=0 $Y2=0
cc_192 N_A_40_480#_c_242_n N_X_c_371_n 0.00751764f $X=2.565 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_40_480#_c_246_n N_X_c_371_n 0.00656419f $X=2.885 $Y=1.35 $X2=0 $Y2=0
cc_194 N_A_40_480#_c_239_n N_VGND_M1001_d 0.0053212f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_195 N_A_40_480#_c_242_n N_VGND_M1002_d 4.51105e-19 $X=2.565 $Y=1.16 $X2=0
+ $Y2=0
cc_196 N_A_40_480#_c_237_n N_VGND_c_389_n 0.00296604f $X=2.65 $Y=1.185 $X2=0
+ $Y2=0
cc_197 N_A_40_480#_c_241_n N_VGND_c_389_n 0.0065956f $X=2.03 $Y=1.075 $X2=0
+ $Y2=0
cc_198 N_A_40_480#_c_242_n N_VGND_c_389_n 0.0196424f $X=2.565 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_40_480#_c_245_n N_VGND_c_389_n 0.0135111f $X=1.972 $Y=0.73 $X2=0
+ $Y2=0
cc_200 N_A_40_480#_c_239_n N_VGND_c_390_n 0.00241405f $X=1.83 $Y=0.73 $X2=0
+ $Y2=0
cc_201 N_A_40_480#_c_284_n N_VGND_c_390_n 0.0149298f $X=1.945 $Y=0.445 $X2=0
+ $Y2=0
cc_202 N_A_40_480#_c_237_n N_VGND_c_392_n 0.0054895f $X=2.65 $Y=1.185 $X2=0
+ $Y2=0
cc_203 N_A_40_480#_M1003_d N_VGND_c_393_n 0.00261603f $X=0.585 $Y=0.235 $X2=0
+ $Y2=0
cc_204 N_A_40_480#_M1000_d N_VGND_c_393_n 0.00258129f $X=1.785 $Y=0.235 $X2=0
+ $Y2=0
cc_205 N_A_40_480#_c_237_n N_VGND_c_393_n 0.011021f $X=2.65 $Y=1.185 $X2=0 $Y2=0
cc_206 N_A_40_480#_c_336_p N_VGND_c_393_n 0.00831597f $X=0.725 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_40_480#_c_239_n N_VGND_c_393_n 0.0113118f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_208 N_A_40_480#_c_284_n N_VGND_c_393_n 0.0106937f $X=1.945 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_A_40_480#_c_336_p N_VGND_c_394_n 0.0114892f $X=0.725 $Y=0.445 $X2=0
+ $Y2=0
cc_210 N_A_40_480#_c_239_n N_VGND_c_394_n 0.00241405f $X=1.83 $Y=0.73 $X2=0
+ $Y2=0
cc_211 N_A_40_480#_c_239_n N_VGND_c_395_n 0.0419672f $X=1.83 $Y=0.73 $X2=0 $Y2=0
cc_212 N_VPWR_c_342_n N_X_M1007_d 0.00371702f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_345_n X 0.018528f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_c_342_n X 0.0104192f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_215 N_X_c_371_n N_VGND_c_392_n 0.0385528f $X=2.865 $Y=0.38 $X2=0 $Y2=0
cc_216 N_X_M1009_d N_VGND_c_393_n 0.00215158f $X=2.725 $Y=0.235 $X2=0 $Y2=0
cc_217 N_X_c_371_n N_VGND_c_393_n 0.02208f $X=2.865 $Y=0.38 $X2=0 $Y2=0
