* File: sky130_fd_sc_lp__clkbuflp_16.pxi.spice
* Created: Fri Aug 28 10:15:35 2020
* 
x_PM_SKY130_FD_SC_LP__CLKBUFLP_16%A N_A_c_166_n N_A_M1018_g N_A_M1005_g
+ N_A_c_168_n N_A_M1002_g N_A_M1016_g N_A_c_170_n N_A_M1007_g N_A_M1025_g
+ N_A_c_172_n N_A_M1009_g N_A_c_173_n N_A_M1021_g N_A_M1029_g N_A_c_175_n
+ N_A_M1033_g N_A_M1046_g N_A_c_177_n N_A_M1038_g N_A_M1047_g N_A_c_179_n
+ N_A_M1035_g A A A N_A_c_181_n PM_SKY130_FD_SC_LP__CLKBUFLP_16%A
x_PM_SKY130_FD_SC_LP__CLKBUFLP_16%A_130_417# N_A_130_417#_M1002_d
+ N_A_130_417#_M1033_d N_A_130_417#_M1005_s N_A_130_417#_M1025_s
+ N_A_130_417#_M1046_s N_A_130_417#_M1010_g N_A_130_417#_M1004_g
+ N_A_130_417#_M1000_g N_A_130_417#_M1006_g N_A_130_417#_M1001_g
+ N_A_130_417#_M1012_g N_A_130_417#_M1008_g N_A_130_417#_M1040_g
+ N_A_130_417#_M1013_g N_A_130_417#_M1003_g N_A_130_417#_M1017_g
+ N_A_130_417#_M1049_g N_A_130_417#_M1022_g N_A_130_417#_M1011_g
+ N_A_130_417#_M1019_g N_A_130_417#_M1023_g N_A_130_417#_M1014_g
+ N_A_130_417#_M1026_g N_A_130_417#_M1030_g N_A_130_417#_M1037_g
+ N_A_130_417#_M1015_g N_A_130_417#_M1020_g N_A_130_417#_M1039_g
+ N_A_130_417#_M1032_g N_A_130_417#_M1041_g N_A_130_417#_M1027_g
+ N_A_130_417#_M1042_g N_A_130_417#_M1024_g N_A_130_417#_M1031_g
+ N_A_130_417#_M1043_g N_A_130_417#_M1028_g N_A_130_417#_M1044_g
+ N_A_130_417#_M1036_g N_A_130_417#_M1045_g N_A_130_417#_M1034_g
+ N_A_130_417#_M1048_g N_A_130_417#_c_355_n N_A_130_417#_c_357_n
+ N_A_130_417#_c_363_n N_A_130_417#_c_364_n N_A_130_417#_c_369_n
+ N_A_130_417#_c_374_n N_A_130_417#_c_351_n N_A_130_417#_c_326_n
+ N_A_130_417#_c_388_n N_A_130_417#_c_390_n N_A_130_417#_c_391_n
+ N_A_130_417#_c_392_n N_A_130_417#_c_327_n N_A_130_417#_c_328_n
+ N_A_130_417#_c_329_n N_A_130_417#_c_330_n N_A_130_417#_c_331_n
+ N_A_130_417#_c_332_n N_A_130_417#_c_333_n N_A_130_417#_c_334_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_16%A_130_417#
x_PM_SKY130_FD_SC_LP__CLKBUFLP_16%VPWR N_VPWR_M1005_d N_VPWR_M1016_d
+ N_VPWR_M1029_d N_VPWR_M1047_d N_VPWR_M1006_d N_VPWR_M1013_d N_VPWR_M1022_d
+ N_VPWR_M1026_d N_VPWR_M1039_d N_VPWR_M1042_d N_VPWR_M1044_d N_VPWR_M1048_d
+ N_VPWR_c_722_n N_VPWR_c_723_n N_VPWR_c_724_n N_VPWR_c_725_n N_VPWR_c_726_n
+ N_VPWR_c_727_n N_VPWR_c_728_n N_VPWR_c_729_n N_VPWR_c_730_n N_VPWR_c_731_n
+ N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_735_n N_VPWR_c_736_n
+ N_VPWR_c_737_n N_VPWR_c_738_n N_VPWR_c_739_n N_VPWR_c_740_n N_VPWR_c_741_n
+ N_VPWR_c_742_n N_VPWR_c_743_n N_VPWR_c_744_n N_VPWR_c_745_n N_VPWR_c_746_n
+ VPWR N_VPWR_c_747_n N_VPWR_c_748_n N_VPWR_c_749_n N_VPWR_c_750_n
+ N_VPWR_c_751_n N_VPWR_c_721_n N_VPWR_c_753_n N_VPWR_c_754_n N_VPWR_c_755_n
+ N_VPWR_c_756_n N_VPWR_c_757_n N_VPWR_c_758_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_16%VPWR
x_PM_SKY130_FD_SC_LP__CLKBUFLP_16%X N_X_M1000_d N_X_M1003_d N_X_M1014_d
+ N_X_M1032_d N_X_M1028_d N_X_M1004_s N_X_M1012_s N_X_M1017_s N_X_M1023_s
+ N_X_M1037_s N_X_M1041_s N_X_M1043_s N_X_M1045_s N_X_c_954_n N_X_c_935_n
+ N_X_c_968_n N_X_c_972_n N_X_c_936_n N_X_c_982_n N_X_c_986_n N_X_c_937_n
+ N_X_c_938_n N_X_c_939_n N_X_c_940_n X N_X_c_945_n N_X_c_946_n N_X_c_1043_n
+ N_X_c_1046_n N_X_c_947_n N_X_c_948_n N_X_c_1062_n N_X_c_949_n N_X_c_950_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_16%X
x_PM_SKY130_FD_SC_LP__CLKBUFLP_16%VGND N_VGND_M1018_s N_VGND_M1009_s
+ N_VGND_M1035_s N_VGND_M1008_s N_VGND_M1011_s N_VGND_M1015_s N_VGND_M1024_s
+ N_VGND_M1034_s N_VGND_c_1173_n N_VGND_c_1174_n N_VGND_c_1175_n N_VGND_c_1176_n
+ N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n N_VGND_c_1180_n
+ N_VGND_c_1181_n N_VGND_c_1182_n N_VGND_c_1183_n N_VGND_c_1184_n
+ N_VGND_c_1185_n VGND N_VGND_c_1186_n N_VGND_c_1187_n N_VGND_c_1188_n
+ N_VGND_c_1189_n N_VGND_c_1190_n N_VGND_c_1191_n N_VGND_c_1192_n
+ N_VGND_c_1193_n N_VGND_c_1194_n N_VGND_c_1195_n N_VGND_c_1196_n
+ N_VGND_c_1197_n PM_SKY130_FD_SC_LP__CLKBUFLP_16%VGND
cc_1 VNB N_A_c_166_n 0.0179343f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.895
cc_2 VNB N_A_M1005_g 0.00588564f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.585
cc_3 VNB N_A_c_168_n 0.0149762f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.895
cc_4 VNB N_A_M1016_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.585
cc_5 VNB N_A_c_170_n 0.0149941f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=0.895
cc_6 VNB N_A_M1025_g 0.00509213f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.585
cc_7 VNB N_A_c_172_n 0.0152614f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=0.895
cc_8 VNB N_A_c_173_n 0.0152614f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=0.895
cc_9 VNB N_A_M1029_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.585
cc_10 VNB N_A_c_175_n 0.0149941f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=0.895
cc_11 VNB N_A_M1046_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.585
cc_12 VNB N_A_c_177_n 0.0149957f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=0.895
cc_13 VNB N_A_M1047_g 0.00527519f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.585
cc_14 VNB N_A_c_179_n 0.0156424f $X=-0.19 $Y=-0.245 $X2=3.205 $Y2=0.895
cc_15 VNB A 0.0397639f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_A_c_181_n 0.266876f $X=-0.19 $Y=-0.245 $X2=3.205 $Y2=1.23
cc_17 VNB N_A_130_417#_M1010_g 0.0307422f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=1.565
cc_18 VNB N_A_130_417#_M1004_g 0.00689281f $X=-0.19 $Y=-0.245 $X2=1.625
+ $Y2=0.895
cc_19 VNB N_A_130_417#_M1000_g 0.0283879f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=0.51
cc_20 VNB N_A_130_417#_M1006_g 0.00578869f $X=-0.19 $Y=-0.245 $X2=2.115
+ $Y2=2.585
cc_21 VNB N_A_130_417#_M1001_g 0.0283982f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=0.51
cc_22 VNB N_A_130_417#_M1012_g 0.00668071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_130_417#_M1008_g 0.0298646f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=1.565
cc_24 VNB N_A_130_417#_M1040_g 0.0298646f $X=-0.19 $Y=-0.245 $X2=3.205 $Y2=0.895
cc_25 VNB N_A_130_417#_M1013_g 0.0066789f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_26 VNB N_A_130_417#_M1003_g 0.0284115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_130_417#_M1017_g 0.00578869f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.23
cc_28 VNB N_A_130_417#_M1049_g 0.028362f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.23
cc_29 VNB N_A_130_417#_M1022_g 0.00624034f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=1.23
cc_30 VNB N_A_130_417#_M1011_g 0.029872f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=1.23
cc_31 VNB N_A_130_417#_M1019_g 0.0298687f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=0.925
cc_32 VNB N_A_130_417#_M1023_g 0.00624034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_130_417#_M1014_g 0.028362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_130_417#_M1026_g 0.00578869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_130_417#_M1030_g 0.0284115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_130_417#_M1037_g 0.00668246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_130_417#_M1015_g 0.0298646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_130_417#_M1020_g 0.0298502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_130_417#_M1039_g 0.00667696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_130_417#_M1032_g 0.0284115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_130_417#_M1041_g 0.00578869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_130_417#_M1027_g 0.0283664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_130_417#_M1042_g 0.00624034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_130_417#_M1024_g 0.0298577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_130_417#_M1031_g 0.0298688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_130_417#_M1043_g 0.00624031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_130_417#_M1028_g 0.028362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_130_417#_M1044_g 0.00624442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_130_417#_M1036_g 0.0284012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_130_417#_M1045_g 0.00668415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_130_417#_M1034_g 0.0439353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_130_417#_M1048_g 0.0102035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_130_417#_c_326_n 8.32813e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_130_417#_c_327_n 0.00913155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_130_417#_c_328_n 0.00548966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_130_417#_c_329_n 0.00241669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_130_417#_c_330_n 0.0054933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_130_417#_c_331_n 0.00224443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_130_417#_c_332_n 0.0930195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_130_417#_c_333_n 0.42179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_130_417#_c_334_n 0.0235889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VPWR_c_721_n 0.521925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_X_c_935_n 0.00241701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_X_c_936_n 5.57045e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_X_c_937_n 0.00777018f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=1.23
cc_66 VNB N_X_c_938_n 0.00616132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_X_c_939_n 0.00931594f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.06
cc_68 VNB N_X_c_940_n 0.00402829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1173_n 0.0107201f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=0.895
cc_70 VNB N_VGND_c_1174_n 0.016276f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=0.51
cc_71 VNB N_VGND_c_1175_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1176_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.565
cc_73 VNB N_VGND_c_1177_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=0.895
cc_74 VNB N_VGND_c_1178_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.585
cc_75 VNB N_VGND_c_1179_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=3.205 $Y2=0.51
cc_76 VNB N_VGND_c_1180_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_77 VNB N_VGND_c_1181_n 0.0173614f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.23
cc_78 VNB N_VGND_c_1182_n 0.0344559f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.23
cc_79 VNB N_VGND_c_1183_n 0.00436918f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.06
cc_80 VNB N_VGND_c_1184_n 0.0345943f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.23
cc_81 VNB N_VGND_c_1185_n 0.00436918f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.23
cc_82 VNB N_VGND_c_1186_n 0.0344559f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.23
cc_83 VNB N_VGND_c_1187_n 0.0352307f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.295
cc_84 VNB N_VGND_c_1188_n 0.0345943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1189_n 0.0345943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1190_n 0.0345943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1191_n 0.0331697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1192_n 0.604587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1193_n 0.00436918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1194_n 0.00436918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1195_n 0.00436918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1196_n 0.00436918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1197_n 0.00510891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VPB N_A_M1005_g 0.0532342f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.585
cc_95 VPB N_A_M1016_g 0.0405497f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.585
cc_96 VPB N_A_M1025_g 0.0402651f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.585
cc_97 VPB N_A_M1029_g 0.0403586f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.585
cc_98 VPB N_A_M1046_g 0.0403586f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.585
cc_99 VPB N_A_M1047_g 0.0411978f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=2.585
cc_100 VPB A 0.0102435f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_101 VPB N_A_130_417#_M1004_g 0.0413889f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=0.895
cc_102 VPB N_A_130_417#_M1006_g 0.0387555f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.585
cc_103 VPB N_A_130_417#_M1012_g 0.0407434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_130_417#_M1013_g 0.0407878f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_105 VPB N_A_130_417#_M1017_g 0.0391333f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.23
cc_106 VPB N_A_130_417#_M1022_g 0.0396878f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=1.23
cc_107 VPB N_A_130_417#_M1023_g 0.0396878f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_130_417#_M1026_g 0.0391333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_130_417#_M1037_g 0.0407922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_130_417#_M1039_g 0.0407682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_130_417#_M1041_g 0.0391375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_130_417#_M1042_g 0.0396878f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_130_417#_M1043_g 0.0396704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_130_417#_M1044_g 0.0396978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_130_417#_M1045_g 0.0407943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_130_417#_M1048_g 0.0574004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_130_417#_c_351_n 0.0057534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_130_417#_c_326_n 0.00349467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_722_n 0.0103398f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.585
cc_120 VPB N_VPWR_c_723_n 0.0468912f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=0.895
cc_121 VPB N_VPWR_c_724_n 0.00581683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_725_n 0.00268334f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_123 VPB N_VPWR_c_726_n 0.00308897f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.23
cc_124 VPB N_VPWR_c_727_n 0.00263836f $X=-0.19 $Y=1.655 $X2=1.265 $Y2=1.23
cc_125 VPB N_VPWR_c_728_n 0.00263836f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=1.23
cc_126 VPB N_VPWR_c_729_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_730_n 0.00192114f $X=-0.19 $Y=1.655 $X2=0.41 $Y2=1.295
cc_128 VPB N_VPWR_c_731_n 0.00258651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_732_n 0.00250384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_733_n 0.00192114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_734_n 0.00249606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_735_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_736_n 0.0494031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_737_n 0.0198321f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_738_n 0.00375865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_739_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_740_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_741_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_742_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_743_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_744_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_745_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_746_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_747_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_748_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_749_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_750_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_751_n 0.014713f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_721_n 0.0572293f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_753_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_754_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_755_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_756_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_757_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_758_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_X_c_935_n 0.00616477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_X_c_937_n 0.00206422f $X=-0.19 $Y=1.655 $X2=2.845 $Y2=1.23
cc_158 VPB N_X_c_938_n 0.00174467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_X_c_939_n 0.00288582f $X=-0.19 $Y=1.655 $X2=0.41 $Y2=1.06
cc_160 VPB N_X_c_945_n 6.79904e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_X_c_946_n 0.00195079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_X_c_947_n 0.00195079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_X_c_948_n 6.44256e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_X_c_949_n 0.00195407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_X_c_950_n 0.0222756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 N_A_c_179_n N_A_130_417#_M1010_g 0.0181566f $X=3.205 $Y=0.895 $X2=0 $Y2=0
cc_167 N_A_c_181_n N_A_130_417#_M1010_g 0.0324925f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_168 N_A_M1005_g N_A_130_417#_c_355_n 0.0164409f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_169 N_A_M1016_g N_A_130_417#_c_355_n 0.0172367f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_170 N_A_c_166_n N_A_130_417#_c_357_n 0.00187286f $X=0.475 $Y=0.895 $X2=0
+ $Y2=0
cc_171 N_A_c_168_n N_A_130_417#_c_357_n 0.0129284f $X=0.835 $Y=0.895 $X2=0 $Y2=0
cc_172 N_A_c_170_n N_A_130_417#_c_357_n 0.0144779f $X=1.265 $Y=0.895 $X2=0 $Y2=0
cc_173 N_A_c_172_n N_A_130_417#_c_357_n 0.00244168f $X=1.625 $Y=0.895 $X2=0
+ $Y2=0
cc_174 A N_A_130_417#_c_357_n 0.0314936f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A_c_181_n N_A_130_417#_c_357_n 0.0317654f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_176 N_A_c_181_n N_A_130_417#_c_363_n 0.0503827f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_177 N_A_M1016_g N_A_130_417#_c_364_n 0.00162903f $X=1.055 $Y=2.585 $X2=0
+ $Y2=0
cc_178 N_A_M1025_g N_A_130_417#_c_364_n 0.0340433f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_179 N_A_M1029_g N_A_130_417#_c_364_n 0.0335321f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_180 N_A_M1046_g N_A_130_417#_c_364_n 0.00223092f $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_181 N_A_c_181_n N_A_130_417#_c_364_n 0.00558636f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_182 N_A_c_173_n N_A_130_417#_c_369_n 0.00244168f $X=2.055 $Y=0.895 $X2=0
+ $Y2=0
cc_183 N_A_c_175_n N_A_130_417#_c_369_n 0.0144779f $X=2.415 $Y=0.895 $X2=0 $Y2=0
cc_184 N_A_c_177_n N_A_130_417#_c_369_n 0.0137574f $X=2.845 $Y=0.895 $X2=0 $Y2=0
cc_185 N_A_c_179_n N_A_130_417#_c_369_n 0.0023736f $X=3.205 $Y=0.895 $X2=0 $Y2=0
cc_186 N_A_c_181_n N_A_130_417#_c_369_n 0.0392067f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_187 N_A_M1029_g N_A_130_417#_c_374_n 0.00223092f $X=2.115 $Y=2.585 $X2=0
+ $Y2=0
cc_188 N_A_M1046_g N_A_130_417#_c_374_n 0.0335321f $X=2.645 $Y=2.585 $X2=0 $Y2=0
cc_189 N_A_M1047_g N_A_130_417#_c_374_n 0.0335321f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_190 N_A_c_181_n N_A_130_417#_c_374_n 0.00653214f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_191 N_A_M1005_g N_A_130_417#_c_351_n 0.00807709f $X=0.525 $Y=2.585 $X2=0
+ $Y2=0
cc_192 N_A_M1016_g N_A_130_417#_c_351_n 0.00576474f $X=1.055 $Y=2.585 $X2=0
+ $Y2=0
cc_193 N_A_M1025_g N_A_130_417#_c_351_n 2.92044e-19 $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_194 A N_A_130_417#_c_351_n 0.00399643f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A_c_181_n N_A_130_417#_c_351_n 0.00360216f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_196 N_A_M1005_g N_A_130_417#_c_326_n 0.00609732f $X=0.525 $Y=2.585 $X2=0
+ $Y2=0
cc_197 N_A_M1016_g N_A_130_417#_c_326_n 0.0147265f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_198 N_A_M1025_g N_A_130_417#_c_326_n 0.00166752f $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_199 A N_A_130_417#_c_326_n 0.0105986f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_200 N_A_c_181_n N_A_130_417#_c_326_n 0.00167458f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_201 A N_A_130_417#_c_388_n 0.0251886f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_202 N_A_c_181_n N_A_130_417#_c_388_n 0.0248096f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_203 N_A_c_181_n N_A_130_417#_c_390_n 0.0194179f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_204 N_A_c_181_n N_A_130_417#_c_391_n 0.0474044f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_205 N_A_c_181_n N_A_130_417#_c_392_n 0.0485554f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_206 N_A_c_181_n N_A_130_417#_c_327_n 0.0270022f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_207 N_A_c_181_n N_A_130_417#_c_332_n 0.0125638f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_208 N_A_M1047_g N_A_130_417#_c_333_n 0.0324925f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_209 N_A_M1005_g N_VPWR_c_723_n 0.0234468f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_210 N_A_M1016_g N_VPWR_c_723_n 0.00115344f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_211 A N_VPWR_c_723_n 0.0191914f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_212 N_A_M1016_g N_VPWR_c_724_n 0.00321157f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_213 N_A_M1025_g N_VPWR_c_724_n 0.0227327f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_214 N_A_M1029_g N_VPWR_c_724_n 0.00117568f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_215 N_A_c_181_n N_VPWR_c_724_n 0.00217526f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_216 N_A_M1025_g N_VPWR_c_725_n 9.25377e-19 $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_217 N_A_M1029_g N_VPWR_c_725_n 0.0227384f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_218 N_A_M1046_g N_VPWR_c_725_n 0.0227384f $X=2.645 $Y=2.585 $X2=0 $Y2=0
cc_219 N_A_M1047_g N_VPWR_c_725_n 9.25377e-19 $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_220 N_A_c_181_n N_VPWR_c_725_n 0.00214033f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_221 N_A_M1046_g N_VPWR_c_726_n 9.25377e-19 $X=2.645 $Y=2.585 $X2=0 $Y2=0
cc_222 N_A_M1047_g N_VPWR_c_726_n 0.022713f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_223 N_A_M1005_g N_VPWR_c_737_n 0.00794322f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_224 N_A_M1016_g N_VPWR_c_737_n 0.00787395f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_225 N_A_M1025_g N_VPWR_c_739_n 0.00839865f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_226 N_A_M1029_g N_VPWR_c_739_n 0.00839865f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_227 N_A_M1046_g N_VPWR_c_741_n 0.00839865f $X=2.645 $Y=2.585 $X2=0 $Y2=0
cc_228 N_A_M1047_g N_VPWR_c_741_n 0.00839865f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_229 N_A_M1005_g N_VPWR_c_721_n 0.012523f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_230 N_A_M1016_g N_VPWR_c_721_n 0.0123608f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_231 N_A_M1025_g N_VPWR_c_721_n 0.0136348f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_232 N_A_M1029_g N_VPWR_c_721_n 0.0136348f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_233 N_A_M1046_g N_VPWR_c_721_n 0.0136348f $X=2.645 $Y=2.585 $X2=0 $Y2=0
cc_234 N_A_M1047_g N_VPWR_c_721_n 0.0136348f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_235 N_A_M1047_g N_X_c_935_n 7.18504e-19 $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_236 N_A_M1047_g N_X_c_945_n 0.00139237f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_237 N_A_M1047_g N_X_c_950_n 7.33163e-19 $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_238 A N_VGND_M1018_s 0.00230452f $X=0.155 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_239 N_A_c_166_n N_VGND_c_1174_n 0.0122997f $X=0.475 $Y=0.895 $X2=0 $Y2=0
cc_240 N_A_c_168_n N_VGND_c_1174_n 0.00219969f $X=0.835 $Y=0.895 $X2=0 $Y2=0
cc_241 A N_VGND_c_1174_n 0.0209431f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_242 N_A_c_170_n N_VGND_c_1175_n 0.00219945f $X=1.265 $Y=0.895 $X2=0 $Y2=0
cc_243 N_A_c_172_n N_VGND_c_1175_n 0.0114626f $X=1.625 $Y=0.895 $X2=0 $Y2=0
cc_244 N_A_c_173_n N_VGND_c_1175_n 0.0114624f $X=2.055 $Y=0.895 $X2=0 $Y2=0
cc_245 N_A_c_175_n N_VGND_c_1175_n 0.00219945f $X=2.415 $Y=0.895 $X2=0 $Y2=0
cc_246 N_A_c_181_n N_VGND_c_1175_n 0.00282316f $X=3.205 $Y=1.23 $X2=0 $Y2=0
cc_247 N_A_c_177_n N_VGND_c_1176_n 0.00220741f $X=2.845 $Y=0.895 $X2=0 $Y2=0
cc_248 N_A_c_179_n N_VGND_c_1176_n 0.0115825f $X=3.205 $Y=0.895 $X2=0 $Y2=0
cc_249 N_A_c_173_n N_VGND_c_1182_n 0.00486043f $X=2.055 $Y=0.895 $X2=0 $Y2=0
cc_250 N_A_c_175_n N_VGND_c_1182_n 0.00526721f $X=2.415 $Y=0.895 $X2=0 $Y2=0
cc_251 N_A_c_177_n N_VGND_c_1182_n 0.00549284f $X=2.845 $Y=0.895 $X2=0 $Y2=0
cc_252 N_A_c_179_n N_VGND_c_1182_n 0.00486043f $X=3.205 $Y=0.895 $X2=0 $Y2=0
cc_253 N_A_c_166_n N_VGND_c_1186_n 0.00486043f $X=0.475 $Y=0.895 $X2=0 $Y2=0
cc_254 N_A_c_168_n N_VGND_c_1186_n 0.00549284f $X=0.835 $Y=0.895 $X2=0 $Y2=0
cc_255 N_A_c_170_n N_VGND_c_1186_n 0.00526721f $X=1.265 $Y=0.895 $X2=0 $Y2=0
cc_256 N_A_c_172_n N_VGND_c_1186_n 0.00486043f $X=1.625 $Y=0.895 $X2=0 $Y2=0
cc_257 N_A_c_166_n N_VGND_c_1192_n 0.00426996f $X=0.475 $Y=0.895 $X2=0 $Y2=0
cc_258 N_A_c_168_n N_VGND_c_1192_n 0.00987174f $X=0.835 $Y=0.895 $X2=0 $Y2=0
cc_259 N_A_c_170_n N_VGND_c_1192_n 0.009316f $X=1.265 $Y=0.895 $X2=0 $Y2=0
cc_260 N_A_c_172_n N_VGND_c_1192_n 0.00814425f $X=1.625 $Y=0.895 $X2=0 $Y2=0
cc_261 N_A_c_173_n N_VGND_c_1192_n 0.00814425f $X=2.055 $Y=0.895 $X2=0 $Y2=0
cc_262 N_A_c_175_n N_VGND_c_1192_n 0.009316f $X=2.415 $Y=0.895 $X2=0 $Y2=0
cc_263 N_A_c_177_n N_VGND_c_1192_n 0.00987174f $X=2.845 $Y=0.895 $X2=0 $Y2=0
cc_264 N_A_c_179_n N_VGND_c_1192_n 0.00814425f $X=3.205 $Y=0.895 $X2=0 $Y2=0
cc_265 A N_VGND_c_1192_n 0.0115239f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_266 A A_110_47# 0.00206043f $X=0.155 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_267 N_A_130_417#_c_351_n N_VPWR_c_723_n 0.0777308f $X=0.79 $Y=2.23 $X2=0
+ $Y2=0
cc_268 N_A_130_417#_c_363_n N_VPWR_c_724_n 0.0090108f $X=1.685 $Y=1.37 $X2=0
+ $Y2=0
cc_269 N_A_130_417#_c_364_n N_VPWR_c_724_n 0.065356f $X=1.85 $Y=2.23 $X2=0 $Y2=0
cc_270 N_A_130_417#_c_351_n N_VPWR_c_724_n 0.0405957f $X=0.79 $Y=2.23 $X2=0
+ $Y2=0
cc_271 N_A_130_417#_c_364_n N_VPWR_c_725_n 0.0652318f $X=1.85 $Y=2.23 $X2=0
+ $Y2=0
cc_272 N_A_130_417#_c_374_n N_VPWR_c_725_n 0.0652318f $X=2.91 $Y=2.23 $X2=0
+ $Y2=0
cc_273 N_A_130_417#_c_392_n N_VPWR_c_725_n 0.00852535f $X=2.45 $Y=1.357 $X2=0
+ $Y2=0
cc_274 N_A_130_417#_M1004_g N_VPWR_c_726_n 0.022677f $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_275 N_A_130_417#_M1006_g N_VPWR_c_726_n 9.25377e-19 $X=4.235 $Y=2.585 $X2=0
+ $Y2=0
cc_276 N_A_130_417#_c_374_n N_VPWR_c_726_n 0.0652318f $X=2.91 $Y=2.23 $X2=0
+ $Y2=0
cc_277 N_A_130_417#_c_327_n N_VPWR_c_726_n 0.0097636f $X=3.6 $Y=1.295 $X2=0
+ $Y2=0
cc_278 N_A_130_417#_M1004_g N_VPWR_c_727_n 9.25377e-19 $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_279 N_A_130_417#_M1006_g N_VPWR_c_727_n 0.0219427f $X=4.235 $Y=2.585 $X2=0
+ $Y2=0
cc_280 N_A_130_417#_M1012_g N_VPWR_c_727_n 0.0221625f $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_281 N_A_130_417#_M1013_g N_VPWR_c_727_n 9.25377e-19 $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_282 N_A_130_417#_c_328_n N_VPWR_c_727_n 9.52051e-19 $X=5.04 $Y=1.295 $X2=0
+ $Y2=0
cc_283 N_A_130_417#_c_333_n N_VPWR_c_727_n 0.00249543f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_284 N_A_130_417#_M1012_g N_VPWR_c_728_n 9.25377e-19 $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_285 N_A_130_417#_M1013_g N_VPWR_c_728_n 0.0222781f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_286 N_A_130_417#_M1017_g N_VPWR_c_728_n 0.022015f $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_287 N_A_130_417#_M1022_g N_VPWR_c_728_n 9.25377e-19 $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_288 N_A_130_417#_c_333_n N_VPWR_c_728_n 0.00249543f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_289 N_A_130_417#_M1017_g N_VPWR_c_729_n 0.00839865f $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_290 N_A_130_417#_M1022_g N_VPWR_c_729_n 0.00839865f $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_291 N_A_130_417#_M1017_g N_VPWR_c_730_n 9.25377e-19 $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_292 N_A_130_417#_M1022_g N_VPWR_c_730_n 0.0222379f $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_293 N_A_130_417#_M1023_g N_VPWR_c_730_n 0.0221625f $X=6.885 $Y=2.585 $X2=0
+ $Y2=0
cc_294 N_A_130_417#_M1026_g N_VPWR_c_730_n 9.25377e-19 $X=7.415 $Y=2.585 $X2=0
+ $Y2=0
cc_295 N_A_130_417#_c_329_n N_VPWR_c_730_n 0.00426821f $X=6.635 $Y=1.295 $X2=0
+ $Y2=0
cc_296 N_A_130_417#_c_333_n N_VPWR_c_730_n 0.00167771f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_297 N_A_130_417#_M1023_g N_VPWR_c_731_n 9.25377e-19 $X=6.885 $Y=2.585 $X2=0
+ $Y2=0
cc_298 N_A_130_417#_M1026_g N_VPWR_c_731_n 0.022015f $X=7.415 $Y=2.585 $X2=0
+ $Y2=0
cc_299 N_A_130_417#_M1037_g N_VPWR_c_731_n 0.0221625f $X=7.945 $Y=2.585 $X2=0
+ $Y2=0
cc_300 N_A_130_417#_M1039_g N_VPWR_c_731_n 9.25377e-19 $X=8.475 $Y=2.585 $X2=0
+ $Y2=0
cc_301 N_A_130_417#_c_330_n N_VPWR_c_731_n 0.00116707f $X=8.4 $Y=1.295 $X2=0
+ $Y2=0
cc_302 N_A_130_417#_c_333_n N_VPWR_c_731_n 0.00249543f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_303 N_A_130_417#_M1037_g N_VPWR_c_732_n 9.25377e-19 $X=7.945 $Y=2.585 $X2=0
+ $Y2=0
cc_304 N_A_130_417#_M1039_g N_VPWR_c_732_n 0.0222781f $X=8.475 $Y=2.585 $X2=0
+ $Y2=0
cc_305 N_A_130_417#_M1041_g N_VPWR_c_732_n 0.0220157f $X=9.005 $Y=2.585 $X2=0
+ $Y2=0
cc_306 N_A_130_417#_M1042_g N_VPWR_c_732_n 9.25377e-19 $X=9.535 $Y=2.585 $X2=0
+ $Y2=0
cc_307 N_A_130_417#_c_333_n N_VPWR_c_732_n 0.00249543f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_308 N_A_130_417#_M1041_g N_VPWR_c_733_n 9.25377e-19 $X=9.005 $Y=2.585 $X2=0
+ $Y2=0
cc_309 N_A_130_417#_M1042_g N_VPWR_c_733_n 0.0222379f $X=9.535 $Y=2.585 $X2=0
+ $Y2=0
cc_310 N_A_130_417#_M1043_g N_VPWR_c_733_n 0.0221625f $X=10.065 $Y=2.585 $X2=0
+ $Y2=0
cc_311 N_A_130_417#_M1044_g N_VPWR_c_733_n 9.25377e-19 $X=10.595 $Y=2.585 $X2=0
+ $Y2=0
cc_312 N_A_130_417#_c_331_n N_VPWR_c_733_n 0.00426821f $X=9.84 $Y=1.295 $X2=0
+ $Y2=0
cc_313 N_A_130_417#_c_333_n N_VPWR_c_733_n 0.00172943f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_314 N_A_130_417#_M1043_g N_VPWR_c_734_n 9.25377e-19 $X=10.065 $Y=2.585 $X2=0
+ $Y2=0
cc_315 N_A_130_417#_M1044_g N_VPWR_c_734_n 0.0220722f $X=10.595 $Y=2.585 $X2=0
+ $Y2=0
cc_316 N_A_130_417#_M1045_g N_VPWR_c_734_n 0.0221628f $X=11.125 $Y=2.585 $X2=0
+ $Y2=0
cc_317 N_A_130_417#_M1048_g N_VPWR_c_734_n 9.25377e-19 $X=11.655 $Y=2.585 $X2=0
+ $Y2=0
cc_318 N_A_130_417#_c_333_n N_VPWR_c_734_n 0.00249543f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_319 N_A_130_417#_c_334_n N_VPWR_c_734_n 0.00147753f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_320 N_A_130_417#_M1045_g N_VPWR_c_735_n 0.00839865f $X=11.125 $Y=2.585 $X2=0
+ $Y2=0
cc_321 N_A_130_417#_M1048_g N_VPWR_c_735_n 0.00839865f $X=11.655 $Y=2.585 $X2=0
+ $Y2=0
cc_322 N_A_130_417#_M1045_g N_VPWR_c_736_n 9.25377e-19 $X=11.125 $Y=2.585 $X2=0
+ $Y2=0
cc_323 N_A_130_417#_M1048_g N_VPWR_c_736_n 0.0238638f $X=11.655 $Y=2.585 $X2=0
+ $Y2=0
cc_324 N_A_130_417#_c_333_n N_VPWR_c_736_n 0.00232557f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_325 N_A_130_417#_c_334_n N_VPWR_c_736_n 0.00410842f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_326 N_A_130_417#_c_355_n N_VPWR_c_737_n 0.027786f $X=0.79 $Y=2.91 $X2=0 $Y2=0
cc_327 N_A_130_417#_c_364_n N_VPWR_c_739_n 0.0189236f $X=1.85 $Y=2.23 $X2=0
+ $Y2=0
cc_328 N_A_130_417#_c_374_n N_VPWR_c_741_n 0.0189236f $X=2.91 $Y=2.23 $X2=0
+ $Y2=0
cc_329 N_A_130_417#_M1023_g N_VPWR_c_743_n 0.00839865f $X=6.885 $Y=2.585 $X2=0
+ $Y2=0
cc_330 N_A_130_417#_M1026_g N_VPWR_c_743_n 0.00839865f $X=7.415 $Y=2.585 $X2=0
+ $Y2=0
cc_331 N_A_130_417#_M1037_g N_VPWR_c_745_n 0.00839865f $X=7.945 $Y=2.585 $X2=0
+ $Y2=0
cc_332 N_A_130_417#_M1039_g N_VPWR_c_745_n 0.00839865f $X=8.475 $Y=2.585 $X2=0
+ $Y2=0
cc_333 N_A_130_417#_M1004_g N_VPWR_c_747_n 0.00839865f $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_334 N_A_130_417#_M1006_g N_VPWR_c_747_n 0.00839865f $X=4.235 $Y=2.585 $X2=0
+ $Y2=0
cc_335 N_A_130_417#_M1012_g N_VPWR_c_748_n 0.00839865f $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_336 N_A_130_417#_M1013_g N_VPWR_c_748_n 0.00839865f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_337 N_A_130_417#_M1041_g N_VPWR_c_749_n 0.00839865f $X=9.005 $Y=2.585 $X2=0
+ $Y2=0
cc_338 N_A_130_417#_M1042_g N_VPWR_c_749_n 0.00839865f $X=9.535 $Y=2.585 $X2=0
+ $Y2=0
cc_339 N_A_130_417#_M1043_g N_VPWR_c_750_n 0.00839865f $X=10.065 $Y=2.585 $X2=0
+ $Y2=0
cc_340 N_A_130_417#_M1044_g N_VPWR_c_750_n 0.00839865f $X=10.595 $Y=2.585 $X2=0
+ $Y2=0
cc_341 N_A_130_417#_M1005_s N_VPWR_c_721_n 0.00223559f $X=0.65 $Y=2.085 $X2=0
+ $Y2=0
cc_342 N_A_130_417#_M1025_s N_VPWR_c_721_n 0.00223559f $X=1.71 $Y=2.085 $X2=0
+ $Y2=0
cc_343 N_A_130_417#_M1046_s N_VPWR_c_721_n 0.00223559f $X=2.77 $Y=2.085 $X2=0
+ $Y2=0
cc_344 N_A_130_417#_M1004_g N_VPWR_c_721_n 0.0136348f $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_345 N_A_130_417#_M1006_g N_VPWR_c_721_n 0.0136348f $X=4.235 $Y=2.585 $X2=0
+ $Y2=0
cc_346 N_A_130_417#_M1012_g N_VPWR_c_721_n 0.0136348f $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_347 N_A_130_417#_M1013_g N_VPWR_c_721_n 0.0136348f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_348 N_A_130_417#_M1017_g N_VPWR_c_721_n 0.0136348f $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_349 N_A_130_417#_M1022_g N_VPWR_c_721_n 0.0136348f $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_350 N_A_130_417#_M1023_g N_VPWR_c_721_n 0.0136348f $X=6.885 $Y=2.585 $X2=0
+ $Y2=0
cc_351 N_A_130_417#_M1026_g N_VPWR_c_721_n 0.0136348f $X=7.415 $Y=2.585 $X2=0
+ $Y2=0
cc_352 N_A_130_417#_M1037_g N_VPWR_c_721_n 0.0136348f $X=7.945 $Y=2.585 $X2=0
+ $Y2=0
cc_353 N_A_130_417#_M1039_g N_VPWR_c_721_n 0.0136348f $X=8.475 $Y=2.585 $X2=0
+ $Y2=0
cc_354 N_A_130_417#_M1041_g N_VPWR_c_721_n 0.0136348f $X=9.005 $Y=2.585 $X2=0
+ $Y2=0
cc_355 N_A_130_417#_M1042_g N_VPWR_c_721_n 0.0136348f $X=9.535 $Y=2.585 $X2=0
+ $Y2=0
cc_356 N_A_130_417#_M1043_g N_VPWR_c_721_n 0.0136348f $X=10.065 $Y=2.585 $X2=0
+ $Y2=0
cc_357 N_A_130_417#_M1044_g N_VPWR_c_721_n 0.0136348f $X=10.595 $Y=2.585 $X2=0
+ $Y2=0
cc_358 N_A_130_417#_M1045_g N_VPWR_c_721_n 0.0136348f $X=11.125 $Y=2.585 $X2=0
+ $Y2=0
cc_359 N_A_130_417#_M1048_g N_VPWR_c_721_n 0.0136348f $X=11.655 $Y=2.585 $X2=0
+ $Y2=0
cc_360 N_A_130_417#_c_355_n N_VPWR_c_721_n 0.0168452f $X=0.79 $Y=2.91 $X2=0
+ $Y2=0
cc_361 N_A_130_417#_c_364_n N_VPWR_c_721_n 0.0123859f $X=1.85 $Y=2.23 $X2=0
+ $Y2=0
cc_362 N_A_130_417#_c_374_n N_VPWR_c_721_n 0.0123859f $X=2.91 $Y=2.23 $X2=0
+ $Y2=0
cc_363 N_A_130_417#_M1010_g N_X_c_954_n 0.0030895f $X=3.655 $Y=0.51 $X2=0 $Y2=0
cc_364 N_A_130_417#_M1000_g N_X_c_954_n 0.0131183f $X=4.015 $Y=0.51 $X2=0 $Y2=0
cc_365 N_A_130_417#_M1001_g N_X_c_954_n 0.0130014f $X=4.445 $Y=0.51 $X2=0 $Y2=0
cc_366 N_A_130_417#_M1008_g N_X_c_954_n 0.00380366f $X=4.805 $Y=0.51 $X2=0 $Y2=0
cc_367 N_A_130_417#_M1010_g N_X_c_935_n 7.39268e-19 $X=3.655 $Y=0.51 $X2=0 $Y2=0
cc_368 N_A_130_417#_M1004_g N_X_c_935_n 0.00947745f $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_369 N_A_130_417#_M1000_g N_X_c_935_n 0.00447372f $X=4.015 $Y=0.51 $X2=0 $Y2=0
cc_370 N_A_130_417#_M1006_g N_X_c_935_n 0.0165207f $X=4.235 $Y=2.585 $X2=0 $Y2=0
cc_371 N_A_130_417#_M1001_g N_X_c_935_n 0.00467303f $X=4.445 $Y=0.51 $X2=0 $Y2=0
cc_372 N_A_130_417#_M1012_g N_X_c_935_n 0.00759698f $X=4.765 $Y=2.585 $X2=0
+ $Y2=0
cc_373 N_A_130_417#_c_327_n N_X_c_935_n 0.0319389f $X=3.6 $Y=1.295 $X2=0 $Y2=0
cc_374 N_A_130_417#_c_328_n N_X_c_935_n 0.0206481f $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_375 N_A_130_417#_c_332_n N_X_c_935_n 0.041021f $X=11.76 $Y=1.295 $X2=0 $Y2=0
cc_376 N_A_130_417#_c_333_n N_X_c_935_n 0.0253813f $X=11.755 $Y=1.37 $X2=0 $Y2=0
cc_377 N_A_130_417#_M1040_g N_X_c_968_n 0.00380579f $X=5.235 $Y=0.51 $X2=0 $Y2=0
cc_378 N_A_130_417#_M1003_g N_X_c_968_n 0.0217998f $X=5.595 $Y=0.51 $X2=0 $Y2=0
cc_379 N_A_130_417#_M1049_g N_X_c_968_n 0.0217998f $X=6.025 $Y=0.51 $X2=0 $Y2=0
cc_380 N_A_130_417#_M1011_g N_X_c_968_n 0.00375611f $X=6.385 $Y=0.51 $X2=0 $Y2=0
cc_381 N_A_130_417#_M1019_g N_X_c_972_n 0.00375611f $X=6.815 $Y=0.51 $X2=0 $Y2=0
cc_382 N_A_130_417#_M1014_g N_X_c_972_n 0.0217998f $X=7.175 $Y=0.51 $X2=0 $Y2=0
cc_383 N_A_130_417#_M1030_g N_X_c_972_n 0.0217998f $X=7.605 $Y=0.51 $X2=0 $Y2=0
cc_384 N_A_130_417#_M1015_g N_X_c_972_n 0.00380584f $X=7.965 $Y=0.51 $X2=0 $Y2=0
cc_385 N_A_130_417#_M1020_g N_X_c_936_n 0.00375925f $X=8.395 $Y=0.51 $X2=0 $Y2=0
cc_386 N_A_130_417#_M1032_g N_X_c_936_n 0.0219027f $X=8.755 $Y=0.51 $X2=0 $Y2=0
cc_387 N_A_130_417#_M1027_g N_X_c_936_n 0.0219027f $X=9.185 $Y=0.51 $X2=0 $Y2=0
cc_388 N_A_130_417#_M1024_g N_X_c_936_n 0.00375925f $X=9.545 $Y=0.51 $X2=0 $Y2=0
cc_389 N_A_130_417#_c_332_n N_X_c_936_n 0.00874f $X=11.76 $Y=1.295 $X2=0 $Y2=0
cc_390 N_A_130_417#_c_333_n N_X_c_936_n 0.00107711f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_391 N_A_130_417#_M1031_g N_X_c_982_n 0.00375611f $X=9.975 $Y=0.51 $X2=0 $Y2=0
cc_392 N_A_130_417#_M1028_g N_X_c_982_n 0.0217998f $X=10.335 $Y=0.51 $X2=0 $Y2=0
cc_393 N_A_130_417#_M1036_g N_X_c_982_n 0.0217998f $X=10.765 $Y=0.51 $X2=0 $Y2=0
cc_394 N_A_130_417#_M1034_g N_X_c_982_n 0.0038152f $X=11.125 $Y=0.51 $X2=0 $Y2=0
cc_395 N_A_130_417#_M1000_g N_X_c_986_n 0.00518482f $X=4.015 $Y=0.51 $X2=0 $Y2=0
cc_396 N_A_130_417#_M1001_g N_X_c_986_n 0.00483909f $X=4.445 $Y=0.51 $X2=0 $Y2=0
cc_397 N_A_130_417#_c_332_n N_X_c_986_n 4.57783e-19 $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_398 N_A_130_417#_M1013_g N_X_c_937_n 0.00619305f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_399 N_A_130_417#_M1003_g N_X_c_937_n 7.83167e-19 $X=5.595 $Y=0.51 $X2=0 $Y2=0
cc_400 N_A_130_417#_M1017_g N_X_c_937_n 0.0137996f $X=5.825 $Y=2.585 $X2=0 $Y2=0
cc_401 N_A_130_417#_M1049_g N_X_c_937_n 0.00757137f $X=6.025 $Y=0.51 $X2=0 $Y2=0
cc_402 N_A_130_417#_M1022_g N_X_c_937_n 0.00816497f $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_403 N_A_130_417#_M1011_g N_X_c_937_n 4.48848e-19 $X=6.385 $Y=0.51 $X2=0 $Y2=0
cc_404 N_A_130_417#_M1023_g N_X_c_937_n 0.00266239f $X=6.885 $Y=2.585 $X2=0
+ $Y2=0
cc_405 N_A_130_417#_c_328_n N_X_c_937_n 0.0156828f $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_406 N_A_130_417#_c_329_n N_X_c_937_n 0.018301f $X=6.635 $Y=1.295 $X2=0 $Y2=0
cc_407 N_A_130_417#_c_332_n N_X_c_937_n 0.0681569f $X=11.76 $Y=1.295 $X2=0 $Y2=0
cc_408 N_A_130_417#_c_333_n N_X_c_937_n 0.0361723f $X=11.755 $Y=1.37 $X2=0 $Y2=0
cc_409 N_A_130_417#_M1022_g N_X_c_938_n 0.00266332f $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_410 N_A_130_417#_M1019_g N_X_c_938_n 4.04842e-19 $X=6.815 $Y=0.51 $X2=0 $Y2=0
cc_411 N_A_130_417#_M1023_g N_X_c_938_n 0.00812776f $X=6.885 $Y=2.585 $X2=0
+ $Y2=0
cc_412 N_A_130_417#_M1014_g N_X_c_938_n 0.00753665f $X=7.175 $Y=0.51 $X2=0 $Y2=0
cc_413 N_A_130_417#_M1026_g N_X_c_938_n 0.0134633f $X=7.415 $Y=2.585 $X2=0 $Y2=0
cc_414 N_A_130_417#_M1030_g N_X_c_938_n 7.57428e-19 $X=7.605 $Y=0.51 $X2=0 $Y2=0
cc_415 N_A_130_417#_M1037_g N_X_c_938_n 0.00582966f $X=7.945 $Y=2.585 $X2=0
+ $Y2=0
cc_416 N_A_130_417#_c_329_n N_X_c_938_n 0.021111f $X=6.635 $Y=1.295 $X2=0 $Y2=0
cc_417 N_A_130_417#_c_330_n N_X_c_938_n 0.020471f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_418 N_A_130_417#_c_332_n N_X_c_938_n 0.0634073f $X=11.76 $Y=1.295 $X2=0 $Y2=0
cc_419 N_A_130_417#_c_333_n N_X_c_938_n 0.0336373f $X=11.755 $Y=1.37 $X2=0 $Y2=0
cc_420 N_A_130_417#_M1039_g N_X_c_939_n 0.00636771f $X=8.475 $Y=2.585 $X2=0
+ $Y2=0
cc_421 N_A_130_417#_M1032_g N_X_c_939_n 8.28923e-19 $X=8.755 $Y=0.51 $X2=0 $Y2=0
cc_422 N_A_130_417#_M1041_g N_X_c_939_n 0.0139748f $X=9.005 $Y=2.585 $X2=0 $Y2=0
cc_423 N_A_130_417#_M1027_g N_X_c_939_n 0.00761198f $X=9.185 $Y=0.51 $X2=0 $Y2=0
cc_424 N_A_130_417#_M1042_g N_X_c_939_n 0.00824263f $X=9.535 $Y=2.585 $X2=0
+ $Y2=0
cc_425 N_A_130_417#_M1024_g N_X_c_939_n 4.37272e-19 $X=9.545 $Y=0.51 $X2=0 $Y2=0
cc_426 N_A_130_417#_M1043_g N_X_c_939_n 0.00103838f $X=10.065 $Y=2.585 $X2=0
+ $Y2=0
cc_427 N_A_130_417#_c_330_n N_X_c_939_n 0.0160863f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_428 N_A_130_417#_c_331_n N_X_c_939_n 0.0184068f $X=9.84 $Y=1.295 $X2=0 $Y2=0
cc_429 N_A_130_417#_c_332_n N_X_c_939_n 0.0532058f $X=11.76 $Y=1.295 $X2=0 $Y2=0
cc_430 N_A_130_417#_c_333_n N_X_c_939_n 0.0351674f $X=11.755 $Y=1.37 $X2=0 $Y2=0
cc_431 N_A_130_417#_M1042_g N_X_c_940_n 0.00266381f $X=9.535 $Y=2.585 $X2=0
+ $Y2=0
cc_432 N_A_130_417#_M1031_g N_X_c_940_n 3.89318e-19 $X=9.975 $Y=0.51 $X2=0 $Y2=0
cc_433 N_A_130_417#_M1043_g N_X_c_940_n 0.00815297f $X=10.065 $Y=2.585 $X2=0
+ $Y2=0
cc_434 N_A_130_417#_M1028_g N_X_c_940_n 0.00751767f $X=10.335 $Y=0.51 $X2=0
+ $Y2=0
cc_435 N_A_130_417#_M1044_g N_X_c_940_n 0.0160033f $X=10.595 $Y=2.585 $X2=0
+ $Y2=0
cc_436 N_A_130_417#_M1036_g N_X_c_940_n 7.51268e-19 $X=10.765 $Y=0.51 $X2=0
+ $Y2=0
cc_437 N_A_130_417#_M1045_g N_X_c_940_n 0.00158263f $X=11.125 $Y=2.585 $X2=0
+ $Y2=0
cc_438 N_A_130_417#_c_331_n N_X_c_940_n 0.0210876f $X=9.84 $Y=1.295 $X2=0 $Y2=0
cc_439 N_A_130_417#_c_332_n N_X_c_940_n 0.0614893f $X=11.76 $Y=1.295 $X2=0 $Y2=0
cc_440 N_A_130_417#_c_333_n N_X_c_940_n 0.0326487f $X=11.755 $Y=1.37 $X2=0 $Y2=0
cc_441 N_A_130_417#_c_334_n N_X_c_940_n 0.0204188f $X=11.755 $Y=1.37 $X2=0 $Y2=0
cc_442 N_A_130_417#_M1004_g N_X_c_945_n 0.0236913f $X=3.705 $Y=2.585 $X2=0 $Y2=0
cc_443 N_A_130_417#_M1006_g N_X_c_945_n 0.0236913f $X=4.235 $Y=2.585 $X2=0 $Y2=0
cc_444 N_A_130_417#_M1012_g N_X_c_945_n 0.0012576f $X=4.765 $Y=2.585 $X2=0 $Y2=0
cc_445 N_A_130_417#_M1006_g N_X_c_946_n 0.00106399f $X=4.235 $Y=2.585 $X2=0
+ $Y2=0
cc_446 N_A_130_417#_M1012_g N_X_c_946_n 0.0225373f $X=4.765 $Y=2.585 $X2=0 $Y2=0
cc_447 N_A_130_417#_M1013_g N_X_c_946_n 0.0225373f $X=5.295 $Y=2.585 $X2=0 $Y2=0
cc_448 N_A_130_417#_M1017_g N_X_c_946_n 0.00106399f $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_449 N_A_130_417#_c_328_n N_X_c_946_n 0.00854418f $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_450 N_A_130_417#_c_332_n N_X_c_946_n 4.08285e-19 $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_451 N_A_130_417#_c_333_n N_X_c_946_n 0.00193921f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_452 N_A_130_417#_M1013_g N_X_c_1043_n 0.00162105f $X=5.295 $Y=2.585 $X2=0
+ $Y2=0
cc_453 N_A_130_417#_M1017_g N_X_c_1043_n 0.0263299f $X=5.825 $Y=2.585 $X2=0
+ $Y2=0
cc_454 N_A_130_417#_M1022_g N_X_c_1043_n 0.0263299f $X=6.355 $Y=2.585 $X2=0
+ $Y2=0
cc_455 N_A_130_417#_M1023_g N_X_c_1046_n 0.0263299f $X=6.885 $Y=2.585 $X2=0
+ $Y2=0
cc_456 N_A_130_417#_M1026_g N_X_c_1046_n 0.0263299f $X=7.415 $Y=2.585 $X2=0
+ $Y2=0
cc_457 N_A_130_417#_M1037_g N_X_c_1046_n 0.00162105f $X=7.945 $Y=2.585 $X2=0
+ $Y2=0
cc_458 N_A_130_417#_M1026_g N_X_c_947_n 0.00106399f $X=7.415 $Y=2.585 $X2=0
+ $Y2=0
cc_459 N_A_130_417#_M1037_g N_X_c_947_n 0.0225373f $X=7.945 $Y=2.585 $X2=0 $Y2=0
cc_460 N_A_130_417#_M1039_g N_X_c_947_n 0.0225373f $X=8.475 $Y=2.585 $X2=0 $Y2=0
cc_461 N_A_130_417#_M1041_g N_X_c_947_n 0.00106399f $X=9.005 $Y=2.585 $X2=0
+ $Y2=0
cc_462 N_A_130_417#_c_330_n N_X_c_947_n 0.00854418f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_463 N_A_130_417#_c_332_n N_X_c_947_n 4.08285e-19 $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_464 N_A_130_417#_c_333_n N_X_c_947_n 0.00200044f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_465 N_A_130_417#_M1039_g N_X_c_948_n 0.00162331f $X=8.475 $Y=2.585 $X2=0
+ $Y2=0
cc_466 N_A_130_417#_M1041_g N_X_c_948_n 0.0264375f $X=9.005 $Y=2.585 $X2=0 $Y2=0
cc_467 N_A_130_417#_M1042_g N_X_c_948_n 0.0264375f $X=9.535 $Y=2.585 $X2=0 $Y2=0
cc_468 N_A_130_417#_M1043_g N_X_c_948_n 0.00162331f $X=10.065 $Y=2.585 $X2=0
+ $Y2=0
cc_469 N_A_130_417#_c_332_n N_X_c_948_n 2.5788e-19 $X=11.76 $Y=1.295 $X2=0 $Y2=0
cc_470 N_A_130_417#_c_333_n N_X_c_948_n 3.83988e-19 $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_471 N_A_130_417#_M1043_g N_X_c_1062_n 0.0263299f $X=10.065 $Y=2.585 $X2=0
+ $Y2=0
cc_472 N_A_130_417#_M1044_g N_X_c_1062_n 0.0263299f $X=10.595 $Y=2.585 $X2=0
+ $Y2=0
cc_473 N_A_130_417#_M1045_g N_X_c_1062_n 0.00162105f $X=11.125 $Y=2.585 $X2=0
+ $Y2=0
cc_474 N_A_130_417#_M1044_g N_X_c_949_n 0.00106399f $X=10.595 $Y=2.585 $X2=0
+ $Y2=0
cc_475 N_A_130_417#_M1045_g N_X_c_949_n 0.0225379f $X=11.125 $Y=2.585 $X2=0
+ $Y2=0
cc_476 N_A_130_417#_M1048_g N_X_c_949_n 0.0232394f $X=11.655 $Y=2.585 $X2=0
+ $Y2=0
cc_477 N_A_130_417#_c_332_n N_X_c_949_n 4.08767e-19 $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_478 N_A_130_417#_c_333_n N_X_c_949_n 0.00190916f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_479 N_A_130_417#_c_334_n N_X_c_949_n 0.00851652f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_480 N_A_130_417#_M1004_g N_X_c_950_n 0.00377467f $X=3.705 $Y=2.585 $X2=0
+ $Y2=0
cc_481 N_A_130_417#_M1006_g N_X_c_950_n 0.0119838f $X=4.235 $Y=2.585 $X2=0 $Y2=0
cc_482 N_A_130_417#_M1012_g N_X_c_950_n 0.0128326f $X=4.765 $Y=2.585 $X2=0 $Y2=0
cc_483 N_A_130_417#_M1013_g N_X_c_950_n 0.0129913f $X=5.295 $Y=2.585 $X2=0 $Y2=0
cc_484 N_A_130_417#_M1017_g N_X_c_950_n 0.0120518f $X=5.825 $Y=2.585 $X2=0 $Y2=0
cc_485 N_A_130_417#_M1022_g N_X_c_950_n 0.0136791f $X=6.355 $Y=2.585 $X2=0 $Y2=0
cc_486 N_A_130_417#_M1023_g N_X_c_950_n 0.0135255f $X=6.885 $Y=2.585 $X2=0 $Y2=0
cc_487 N_A_130_417#_M1026_g N_X_c_950_n 0.0120518f $X=7.415 $Y=2.585 $X2=0 $Y2=0
cc_488 N_A_130_417#_M1037_g N_X_c_950_n 0.0128326f $X=7.945 $Y=2.585 $X2=0 $Y2=0
cc_489 N_A_130_417#_M1039_g N_X_c_950_n 0.0130681f $X=8.475 $Y=2.585 $X2=0 $Y2=0
cc_490 N_A_130_417#_M1041_g N_X_c_950_n 0.0120618f $X=9.005 $Y=2.585 $X2=0 $Y2=0
cc_491 N_A_130_417#_M1042_g N_X_c_950_n 0.0136791f $X=9.535 $Y=2.585 $X2=0 $Y2=0
cc_492 N_A_130_417#_M1043_g N_X_c_950_n 0.0135255f $X=10.065 $Y=2.585 $X2=0
+ $Y2=0
cc_493 N_A_130_417#_M1044_g N_X_c_950_n 0.012096f $X=10.595 $Y=2.585 $X2=0 $Y2=0
cc_494 N_A_130_417#_M1045_g N_X_c_950_n 0.0128347f $X=11.125 $Y=2.585 $X2=0
+ $Y2=0
cc_495 N_A_130_417#_M1048_g N_X_c_950_n 0.00752702f $X=11.655 $Y=2.585 $X2=0
+ $Y2=0
cc_496 N_A_130_417#_c_328_n N_X_c_950_n 0.0108655f $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_497 N_A_130_417#_c_329_n N_X_c_950_n 0.00362452f $X=6.635 $Y=1.295 $X2=0
+ $Y2=0
cc_498 N_A_130_417#_c_330_n N_X_c_950_n 0.0107029f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_499 N_A_130_417#_c_331_n N_X_c_950_n 0.00362452f $X=9.84 $Y=1.295 $X2=0 $Y2=0
cc_500 N_A_130_417#_c_332_n N_X_c_950_n 0.36091f $X=11.76 $Y=1.295 $X2=0 $Y2=0
cc_501 N_A_130_417#_c_333_n N_X_c_950_n 0.0124913f $X=11.755 $Y=1.37 $X2=0 $Y2=0
cc_502 N_A_130_417#_c_334_n N_X_c_950_n 0.00704358f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_503 N_A_130_417#_c_357_n N_VGND_c_1174_n 0.0113319f $X=1.05 $Y=0.44 $X2=0
+ $Y2=0
cc_504 N_A_130_417#_c_357_n N_VGND_c_1175_n 0.0117425f $X=1.05 $Y=0.44 $X2=0
+ $Y2=0
cc_505 N_A_130_417#_c_363_n N_VGND_c_1175_n 2.39408e-19 $X=1.685 $Y=1.37 $X2=0
+ $Y2=0
cc_506 N_A_130_417#_c_369_n N_VGND_c_1175_n 0.0117425f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_507 N_A_130_417#_c_390_n N_VGND_c_1175_n 0.0081747f $X=1.85 $Y=1.37 $X2=0
+ $Y2=0
cc_508 N_A_130_417#_M1010_g N_VGND_c_1176_n 0.00990949f $X=3.655 $Y=0.51 $X2=0
+ $Y2=0
cc_509 N_A_130_417#_M1000_g N_VGND_c_1176_n 0.00212931f $X=4.015 $Y=0.51 $X2=0
+ $Y2=0
cc_510 N_A_130_417#_c_369_n N_VGND_c_1176_n 0.0114143f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_511 N_A_130_417#_c_327_n N_VGND_c_1176_n 0.00510807f $X=3.6 $Y=1.295 $X2=0
+ $Y2=0
cc_512 N_A_130_417#_c_332_n N_VGND_c_1176_n 0.00716823f $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_513 N_A_130_417#_M1001_g N_VGND_c_1177_n 0.00220741f $X=4.445 $Y=0.51 $X2=0
+ $Y2=0
cc_514 N_A_130_417#_M1008_g N_VGND_c_1177_n 0.0115246f $X=4.805 $Y=0.51 $X2=0
+ $Y2=0
cc_515 N_A_130_417#_M1040_g N_VGND_c_1177_n 0.0115246f $X=5.235 $Y=0.51 $X2=0
+ $Y2=0
cc_516 N_A_130_417#_M1003_g N_VGND_c_1177_n 0.00220741f $X=5.595 $Y=0.51 $X2=0
+ $Y2=0
cc_517 N_A_130_417#_c_328_n N_VGND_c_1177_n 0.00508451f $X=5.04 $Y=1.295 $X2=0
+ $Y2=0
cc_518 N_A_130_417#_c_332_n N_VGND_c_1177_n 0.00245528f $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_519 N_A_130_417#_c_333_n N_VGND_c_1177_n 6.10932e-19 $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_520 N_A_130_417#_M1049_g N_VGND_c_1178_n 0.00220741f $X=6.025 $Y=0.51 $X2=0
+ $Y2=0
cc_521 N_A_130_417#_M1011_g N_VGND_c_1178_n 0.0115226f $X=6.385 $Y=0.51 $X2=0
+ $Y2=0
cc_522 N_A_130_417#_M1019_g N_VGND_c_1178_n 0.0115246f $X=6.815 $Y=0.51 $X2=0
+ $Y2=0
cc_523 N_A_130_417#_M1014_g N_VGND_c_1178_n 0.00220741f $X=7.175 $Y=0.51 $X2=0
+ $Y2=0
cc_524 N_A_130_417#_c_329_n N_VGND_c_1178_n 0.00463148f $X=6.635 $Y=1.295 $X2=0
+ $Y2=0
cc_525 N_A_130_417#_c_332_n N_VGND_c_1178_n 0.00331917f $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_526 N_A_130_417#_c_333_n N_VGND_c_1178_n 6.10573e-19 $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_527 N_A_130_417#_M1030_g N_VGND_c_1179_n 0.00220741f $X=7.605 $Y=0.51 $X2=0
+ $Y2=0
cc_528 N_A_130_417#_M1015_g N_VGND_c_1179_n 0.0115246f $X=7.965 $Y=0.51 $X2=0
+ $Y2=0
cc_529 N_A_130_417#_M1020_g N_VGND_c_1179_n 0.0115246f $X=8.395 $Y=0.51 $X2=0
+ $Y2=0
cc_530 N_A_130_417#_M1032_g N_VGND_c_1179_n 0.00220741f $X=8.755 $Y=0.51 $X2=0
+ $Y2=0
cc_531 N_A_130_417#_c_330_n N_VGND_c_1179_n 0.00508451f $X=8.4 $Y=1.295 $X2=0
+ $Y2=0
cc_532 N_A_130_417#_c_332_n N_VGND_c_1179_n 0.00245528f $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_533 N_A_130_417#_c_333_n N_VGND_c_1179_n 6.10214e-19 $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_534 N_A_130_417#_M1027_g N_VGND_c_1180_n 0.00220741f $X=9.185 $Y=0.51 $X2=0
+ $Y2=0
cc_535 N_A_130_417#_M1024_g N_VGND_c_1180_n 0.0115226f $X=9.545 $Y=0.51 $X2=0
+ $Y2=0
cc_536 N_A_130_417#_M1031_g N_VGND_c_1180_n 0.0115246f $X=9.975 $Y=0.51 $X2=0
+ $Y2=0
cc_537 N_A_130_417#_M1028_g N_VGND_c_1180_n 0.00220741f $X=10.335 $Y=0.51 $X2=0
+ $Y2=0
cc_538 N_A_130_417#_c_331_n N_VGND_c_1180_n 0.00444328f $X=9.84 $Y=1.295 $X2=0
+ $Y2=0
cc_539 N_A_130_417#_c_332_n N_VGND_c_1180_n 0.0039156f $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_540 N_A_130_417#_c_333_n N_VGND_c_1180_n 6.09855e-19 $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_541 N_A_130_417#_M1036_g N_VGND_c_1181_n 0.00220741f $X=10.765 $Y=0.51 $X2=0
+ $Y2=0
cc_542 N_A_130_417#_M1034_g N_VGND_c_1181_n 0.0126793f $X=11.125 $Y=0.51 $X2=0
+ $Y2=0
cc_543 N_A_130_417#_c_332_n N_VGND_c_1181_n 0.00726742f $X=11.76 $Y=1.295 $X2=0
+ $Y2=0
cc_544 N_A_130_417#_c_333_n N_VGND_c_1181_n 0.00161407f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_545 N_A_130_417#_c_334_n N_VGND_c_1181_n 0.0058429f $X=11.755 $Y=1.37 $X2=0
+ $Y2=0
cc_546 N_A_130_417#_c_369_n N_VGND_c_1182_n 0.0187546f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_547 N_A_130_417#_M1019_g N_VGND_c_1184_n 0.00486043f $X=6.815 $Y=0.51 $X2=0
+ $Y2=0
cc_548 N_A_130_417#_M1014_g N_VGND_c_1184_n 0.00549284f $X=7.175 $Y=0.51 $X2=0
+ $Y2=0
cc_549 N_A_130_417#_M1030_g N_VGND_c_1184_n 0.00549284f $X=7.605 $Y=0.51 $X2=0
+ $Y2=0
cc_550 N_A_130_417#_M1015_g N_VGND_c_1184_n 0.00486043f $X=7.965 $Y=0.51 $X2=0
+ $Y2=0
cc_551 N_A_130_417#_c_357_n N_VGND_c_1186_n 0.0187546f $X=1.05 $Y=0.44 $X2=0
+ $Y2=0
cc_552 N_A_130_417#_M1010_g N_VGND_c_1187_n 0.00564095f $X=3.655 $Y=0.51 $X2=0
+ $Y2=0
cc_553 N_A_130_417#_M1000_g N_VGND_c_1187_n 0.00549284f $X=4.015 $Y=0.51 $X2=0
+ $Y2=0
cc_554 N_A_130_417#_M1001_g N_VGND_c_1187_n 0.00549284f $X=4.445 $Y=0.51 $X2=0
+ $Y2=0
cc_555 N_A_130_417#_M1008_g N_VGND_c_1187_n 0.00486043f $X=4.805 $Y=0.51 $X2=0
+ $Y2=0
cc_556 N_A_130_417#_M1040_g N_VGND_c_1188_n 0.00486043f $X=5.235 $Y=0.51 $X2=0
+ $Y2=0
cc_557 N_A_130_417#_M1003_g N_VGND_c_1188_n 0.00549284f $X=5.595 $Y=0.51 $X2=0
+ $Y2=0
cc_558 N_A_130_417#_M1049_g N_VGND_c_1188_n 0.00549284f $X=6.025 $Y=0.51 $X2=0
+ $Y2=0
cc_559 N_A_130_417#_M1011_g N_VGND_c_1188_n 0.00486043f $X=6.385 $Y=0.51 $X2=0
+ $Y2=0
cc_560 N_A_130_417#_M1020_g N_VGND_c_1189_n 0.00486043f $X=8.395 $Y=0.51 $X2=0
+ $Y2=0
cc_561 N_A_130_417#_M1032_g N_VGND_c_1189_n 0.00549284f $X=8.755 $Y=0.51 $X2=0
+ $Y2=0
cc_562 N_A_130_417#_M1027_g N_VGND_c_1189_n 0.00549284f $X=9.185 $Y=0.51 $X2=0
+ $Y2=0
cc_563 N_A_130_417#_M1024_g N_VGND_c_1189_n 0.00486043f $X=9.545 $Y=0.51 $X2=0
+ $Y2=0
cc_564 N_A_130_417#_M1031_g N_VGND_c_1190_n 0.00486043f $X=9.975 $Y=0.51 $X2=0
+ $Y2=0
cc_565 N_A_130_417#_M1028_g N_VGND_c_1190_n 0.00549284f $X=10.335 $Y=0.51 $X2=0
+ $Y2=0
cc_566 N_A_130_417#_M1036_g N_VGND_c_1190_n 0.00549284f $X=10.765 $Y=0.51 $X2=0
+ $Y2=0
cc_567 N_A_130_417#_M1034_g N_VGND_c_1190_n 0.00486043f $X=11.125 $Y=0.51 $X2=0
+ $Y2=0
cc_568 N_A_130_417#_M1002_d N_VGND_c_1192_n 0.00223819f $X=0.91 $Y=0.235 $X2=0
+ $Y2=0
cc_569 N_A_130_417#_M1033_d N_VGND_c_1192_n 0.00223819f $X=2.49 $Y=0.235 $X2=0
+ $Y2=0
cc_570 N_A_130_417#_M1010_g N_VGND_c_1192_n 0.0093799f $X=3.655 $Y=0.51 $X2=0
+ $Y2=0
cc_571 N_A_130_417#_M1000_g N_VGND_c_1192_n 0.00987174f $X=4.015 $Y=0.51 $X2=0
+ $Y2=0
cc_572 N_A_130_417#_M1001_g N_VGND_c_1192_n 0.00987174f $X=4.445 $Y=0.51 $X2=0
+ $Y2=0
cc_573 N_A_130_417#_M1008_g N_VGND_c_1192_n 0.00814425f $X=4.805 $Y=0.51 $X2=0
+ $Y2=0
cc_574 N_A_130_417#_M1040_g N_VGND_c_1192_n 0.00814425f $X=5.235 $Y=0.51 $X2=0
+ $Y2=0
cc_575 N_A_130_417#_M1003_g N_VGND_c_1192_n 0.00987174f $X=5.595 $Y=0.51 $X2=0
+ $Y2=0
cc_576 N_A_130_417#_M1049_g N_VGND_c_1192_n 0.00987174f $X=6.025 $Y=0.51 $X2=0
+ $Y2=0
cc_577 N_A_130_417#_M1011_g N_VGND_c_1192_n 0.00814425f $X=6.385 $Y=0.51 $X2=0
+ $Y2=0
cc_578 N_A_130_417#_M1019_g N_VGND_c_1192_n 0.00814425f $X=6.815 $Y=0.51 $X2=0
+ $Y2=0
cc_579 N_A_130_417#_M1014_g N_VGND_c_1192_n 0.00987174f $X=7.175 $Y=0.51 $X2=0
+ $Y2=0
cc_580 N_A_130_417#_M1030_g N_VGND_c_1192_n 0.00987174f $X=7.605 $Y=0.51 $X2=0
+ $Y2=0
cc_581 N_A_130_417#_M1015_g N_VGND_c_1192_n 0.00814425f $X=7.965 $Y=0.51 $X2=0
+ $Y2=0
cc_582 N_A_130_417#_M1020_g N_VGND_c_1192_n 0.00814425f $X=8.395 $Y=0.51 $X2=0
+ $Y2=0
cc_583 N_A_130_417#_M1032_g N_VGND_c_1192_n 0.00987174f $X=8.755 $Y=0.51 $X2=0
+ $Y2=0
cc_584 N_A_130_417#_M1027_g N_VGND_c_1192_n 0.00987174f $X=9.185 $Y=0.51 $X2=0
+ $Y2=0
cc_585 N_A_130_417#_M1024_g N_VGND_c_1192_n 0.00814425f $X=9.545 $Y=0.51 $X2=0
+ $Y2=0
cc_586 N_A_130_417#_M1031_g N_VGND_c_1192_n 0.00814425f $X=9.975 $Y=0.51 $X2=0
+ $Y2=0
cc_587 N_A_130_417#_M1028_g N_VGND_c_1192_n 0.00987174f $X=10.335 $Y=0.51 $X2=0
+ $Y2=0
cc_588 N_A_130_417#_M1036_g N_VGND_c_1192_n 0.00987174f $X=10.765 $Y=0.51 $X2=0
+ $Y2=0
cc_589 N_A_130_417#_M1034_g N_VGND_c_1192_n 0.00814425f $X=11.125 $Y=0.51 $X2=0
+ $Y2=0
cc_590 N_A_130_417#_c_357_n N_VGND_c_1192_n 0.012836f $X=1.05 $Y=0.44 $X2=0
+ $Y2=0
cc_591 N_A_130_417#_c_369_n N_VGND_c_1192_n 0.012836f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_721_n N_X_M1004_s 0.00223559f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_593 N_VPWR_c_721_n N_X_M1012_s 0.00223559f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_594 N_VPWR_c_721_n N_X_M1017_s 0.00223559f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_595 N_VPWR_c_721_n N_X_M1023_s 0.00223559f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_596 N_VPWR_c_721_n N_X_M1037_s 0.00223559f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_597 N_VPWR_c_721_n N_X_M1041_s 0.00223559f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_598 N_VPWR_c_721_n N_X_M1043_s 0.00223559f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_599 N_VPWR_c_721_n N_X_M1045_s 0.00223559f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_600 N_VPWR_c_727_n N_X_c_935_n 0.00243974f $X=4.5 $Y=2.23 $X2=0 $Y2=0
cc_601 N_VPWR_c_728_n N_X_c_937_n 0.00245303f $X=5.56 $Y=2.23 $X2=0 $Y2=0
cc_602 N_VPWR_c_731_n N_X_c_938_n 0.00125115f $X=7.68 $Y=2.23 $X2=0 $Y2=0
cc_603 N_VPWR_c_732_n N_X_c_939_n 0.00321135f $X=8.74 $Y=2.23 $X2=0 $Y2=0
cc_604 N_VPWR_c_734_n N_X_c_940_n 6.11785e-19 $X=10.86 $Y=2.23 $X2=0 $Y2=0
cc_605 N_VPWR_c_726_n N_X_c_945_n 0.0643692f $X=3.44 $Y=2.23 $X2=0 $Y2=0
cc_606 N_VPWR_c_727_n N_X_c_945_n 0.0644905f $X=4.5 $Y=2.23 $X2=0 $Y2=0
cc_607 N_VPWR_c_747_n N_X_c_945_n 0.0189236f $X=4.335 $Y=3.33 $X2=0 $Y2=0
cc_608 N_VPWR_c_721_n N_X_c_945_n 0.0123859f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_609 N_VPWR_c_727_n N_X_c_946_n 0.0644905f $X=4.5 $Y=2.23 $X2=0 $Y2=0
cc_610 N_VPWR_c_728_n N_X_c_946_n 0.0644905f $X=5.56 $Y=2.23 $X2=0 $Y2=0
cc_611 N_VPWR_c_748_n N_X_c_946_n 0.0189236f $X=5.395 $Y=3.33 $X2=0 $Y2=0
cc_612 N_VPWR_c_721_n N_X_c_946_n 0.0123859f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_613 N_VPWR_c_728_n N_X_c_1043_n 0.0644905f $X=5.56 $Y=2.23 $X2=0 $Y2=0
cc_614 N_VPWR_c_729_n N_X_c_1043_n 0.0189236f $X=6.455 $Y=3.33 $X2=0 $Y2=0
cc_615 N_VPWR_c_730_n N_X_c_1043_n 0.0644905f $X=6.62 $Y=2.23 $X2=0 $Y2=0
cc_616 N_VPWR_c_721_n N_X_c_1043_n 0.0123859f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_617 N_VPWR_c_730_n N_X_c_1046_n 0.0644905f $X=6.62 $Y=2.23 $X2=0 $Y2=0
cc_618 N_VPWR_c_731_n N_X_c_1046_n 0.0644905f $X=7.68 $Y=2.23 $X2=0 $Y2=0
cc_619 N_VPWR_c_743_n N_X_c_1046_n 0.0189236f $X=7.515 $Y=3.33 $X2=0 $Y2=0
cc_620 N_VPWR_c_721_n N_X_c_1046_n 0.0123859f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_621 N_VPWR_c_731_n N_X_c_947_n 0.0644905f $X=7.68 $Y=2.23 $X2=0 $Y2=0
cc_622 N_VPWR_c_732_n N_X_c_947_n 0.0644905f $X=8.74 $Y=2.23 $X2=0 $Y2=0
cc_623 N_VPWR_c_745_n N_X_c_947_n 0.0189236f $X=8.575 $Y=3.33 $X2=0 $Y2=0
cc_624 N_VPWR_c_721_n N_X_c_947_n 0.0123859f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_625 N_VPWR_c_732_n N_X_c_948_n 0.0644905f $X=8.74 $Y=2.23 $X2=0 $Y2=0
cc_626 N_VPWR_c_733_n N_X_c_948_n 0.0644905f $X=9.8 $Y=2.23 $X2=0 $Y2=0
cc_627 N_VPWR_c_749_n N_X_c_948_n 0.0189236f $X=9.635 $Y=3.33 $X2=0 $Y2=0
cc_628 N_VPWR_c_721_n N_X_c_948_n 0.0123859f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_629 N_VPWR_c_733_n N_X_c_1062_n 0.0644905f $X=9.8 $Y=2.23 $X2=0 $Y2=0
cc_630 N_VPWR_c_734_n N_X_c_1062_n 0.0644905f $X=10.86 $Y=2.23 $X2=0 $Y2=0
cc_631 N_VPWR_c_750_n N_X_c_1062_n 0.0189236f $X=10.695 $Y=3.33 $X2=0 $Y2=0
cc_632 N_VPWR_c_721_n N_X_c_1062_n 0.0123859f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_633 N_VPWR_c_734_n N_X_c_949_n 0.0644905f $X=10.86 $Y=2.23 $X2=0 $Y2=0
cc_634 N_VPWR_c_735_n N_X_c_949_n 0.0189236f $X=11.755 $Y=3.33 $X2=0 $Y2=0
cc_635 N_VPWR_c_736_n N_X_c_949_n 0.0643692f $X=11.92 $Y=2.23 $X2=0 $Y2=0
cc_636 N_VPWR_c_721_n N_X_c_949_n 0.0123859f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_637 N_VPWR_c_726_n N_X_c_950_n 0.00184902f $X=3.44 $Y=2.23 $X2=0 $Y2=0
cc_638 N_VPWR_c_727_n N_X_c_950_n 0.028524f $X=4.5 $Y=2.23 $X2=0 $Y2=0
cc_639 N_VPWR_c_728_n N_X_c_950_n 0.0289694f $X=5.56 $Y=2.23 $X2=0 $Y2=0
cc_640 N_VPWR_c_730_n N_X_c_950_n 0.0268429f $X=6.62 $Y=2.23 $X2=0 $Y2=0
cc_641 N_VPWR_c_731_n N_X_c_950_n 0.0289017f $X=7.68 $Y=2.23 $X2=0 $Y2=0
cc_642 N_VPWR_c_732_n N_X_c_950_n 0.0287191f $X=8.74 $Y=2.23 $X2=0 $Y2=0
cc_643 N_VPWR_c_733_n N_X_c_950_n 0.0268429f $X=9.8 $Y=2.23 $X2=0 $Y2=0
cc_644 N_VPWR_c_734_n N_X_c_950_n 0.0289063f $X=10.86 $Y=2.23 $X2=0 $Y2=0
cc_645 N_VPWR_c_736_n N_X_c_950_n 0.00184902f $X=11.92 $Y=2.23 $X2=0 $Y2=0
cc_646 N_X_c_954_n N_VGND_c_1176_n 0.0109656f $X=4.23 $Y=0.44 $X2=0 $Y2=0
cc_647 N_X_c_954_n N_VGND_c_1177_n 0.0113755f $X=4.23 $Y=0.44 $X2=0 $Y2=0
cc_648 N_X_c_968_n N_VGND_c_1177_n 0.0113755f $X=5.81 $Y=0.44 $X2=0 $Y2=0
cc_649 N_X_c_968_n N_VGND_c_1178_n 0.0113755f $X=5.81 $Y=0.44 $X2=0 $Y2=0
cc_650 N_X_c_972_n N_VGND_c_1178_n 0.0113755f $X=7.39 $Y=0.44 $X2=0 $Y2=0
cc_651 N_X_c_972_n N_VGND_c_1179_n 0.0113755f $X=7.39 $Y=0.44 $X2=0 $Y2=0
cc_652 N_X_c_936_n N_VGND_c_1179_n 0.0113755f $X=8.97 $Y=0.44 $X2=0 $Y2=0
cc_653 N_X_c_936_n N_VGND_c_1180_n 0.0113755f $X=8.97 $Y=0.44 $X2=0 $Y2=0
cc_654 N_X_c_982_n N_VGND_c_1180_n 0.0113755f $X=10.55 $Y=0.44 $X2=0 $Y2=0
cc_655 N_X_c_982_n N_VGND_c_1181_n 0.0113755f $X=10.55 $Y=0.44 $X2=0 $Y2=0
cc_656 N_X_c_972_n N_VGND_c_1184_n 0.0177952f $X=7.39 $Y=0.44 $X2=0 $Y2=0
cc_657 N_X_c_954_n N_VGND_c_1187_n 0.0177952f $X=4.23 $Y=0.44 $X2=0 $Y2=0
cc_658 N_X_c_968_n N_VGND_c_1188_n 0.0177952f $X=5.81 $Y=0.44 $X2=0 $Y2=0
cc_659 N_X_c_936_n N_VGND_c_1189_n 0.0177952f $X=8.97 $Y=0.44 $X2=0 $Y2=0
cc_660 N_X_c_982_n N_VGND_c_1190_n 0.0177952f $X=10.55 $Y=0.44 $X2=0 $Y2=0
cc_661 N_X_M1000_d N_VGND_c_1192_n 0.00223819f $X=4.09 $Y=0.235 $X2=0 $Y2=0
cc_662 N_X_M1003_d N_VGND_c_1192_n 0.00223819f $X=5.67 $Y=0.235 $X2=0 $Y2=0
cc_663 N_X_M1014_d N_VGND_c_1192_n 0.00223819f $X=7.25 $Y=0.235 $X2=0 $Y2=0
cc_664 N_X_M1032_d N_VGND_c_1192_n 0.00223819f $X=8.83 $Y=0.235 $X2=0 $Y2=0
cc_665 N_X_M1028_d N_VGND_c_1192_n 0.00223819f $X=10.41 $Y=0.235 $X2=0 $Y2=0
cc_666 N_X_c_954_n N_VGND_c_1192_n 0.0123247f $X=4.23 $Y=0.44 $X2=0 $Y2=0
cc_667 N_X_c_968_n N_VGND_c_1192_n 0.0123247f $X=5.81 $Y=0.44 $X2=0 $Y2=0
cc_668 N_X_c_972_n N_VGND_c_1192_n 0.0123247f $X=7.39 $Y=0.44 $X2=0 $Y2=0
cc_669 N_X_c_936_n N_VGND_c_1192_n 0.0123247f $X=8.97 $Y=0.44 $X2=0 $Y2=0
cc_670 N_X_c_982_n N_VGND_c_1192_n 0.0123247f $X=10.55 $Y=0.44 $X2=0 $Y2=0
cc_671 N_VGND_c_1192_n A_110_47# 0.00476829f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_672 N_VGND_c_1192_n A_584_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_673 N_VGND_c_1192_n A_268_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_674 N_VGND_c_1192_n A_426_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_675 N_VGND_c_1192_n A_1378_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_676 N_VGND_c_1192_n A_2010_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_677 N_VGND_c_1192_n A_1852_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_678 N_VGND_c_1192_n A_746_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_679 N_VGND_c_1192_n A_904_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_680 N_VGND_c_1192_n A_1536_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_681 N_VGND_c_1192_n A_2168_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_682 N_VGND_c_1192_n A_1062_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_683 N_VGND_c_1192_n A_1220_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
cc_684 N_VGND_c_1192_n A_1694_47# 0.00899413f $X=12.24 $Y=0 $X2=-0.19 $Y2=-0.245
