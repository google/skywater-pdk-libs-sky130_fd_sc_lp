* File: sky130_fd_sc_lp__nor4b_2.pxi.spice
* Created: Wed Sep  2 10:11:01 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4B_2%D_N N_D_N_M1012_g N_D_N_c_90_n N_D_N_M1008_g D_N
+ N_D_N_c_92_n PM_SKY130_FD_SC_LP__NOR4B_2%D_N
x_PM_SKY130_FD_SC_LP__NOR4B_2%C N_C_c_116_n N_C_M1003_g N_C_M1015_g N_C_M1009_g
+ N_C_M1017_g N_C_c_119_n N_C_c_120_n N_C_c_121_n C N_C_c_122_n N_C_c_123_n
+ N_C_c_124_n N_C_c_125_n PM_SKY130_FD_SC_LP__NOR4B_2%C
x_PM_SKY130_FD_SC_LP__NOR4B_2%A_27_535# N_A_27_535#_M1008_s N_A_27_535#_M1012_s
+ N_A_27_535#_M1002_g N_A_27_535#_M1004_g N_A_27_535#_M1014_g
+ N_A_27_535#_M1010_g N_A_27_535#_c_214_n N_A_27_535#_c_207_n
+ N_A_27_535#_c_208_n N_A_27_535#_c_216_n N_A_27_535#_c_217_n
+ N_A_27_535#_c_209_n N_A_27_535#_c_210_n N_A_27_535#_c_211_n
+ PM_SKY130_FD_SC_LP__NOR4B_2%A_27_535#
x_PM_SKY130_FD_SC_LP__NOR4B_2%B N_B_M1001_g N_B_M1000_g N_B_c_292_n N_B_M1005_g
+ N_B_M1016_g N_B_c_294_n N_B_c_295_n B B N_B_c_297_n N_B_c_298_n N_B_c_299_n
+ PM_SKY130_FD_SC_LP__NOR4B_2%B
x_PM_SKY130_FD_SC_LP__NOR4B_2%A N_A_c_370_n N_A_M1007_g N_A_M1006_g N_A_c_372_n
+ N_A_M1011_g N_A_M1013_g A A N_A_c_375_n PM_SKY130_FD_SC_LP__NOR4B_2%A
x_PM_SKY130_FD_SC_LP__NOR4B_2%VPWR N_VPWR_M1012_d N_VPWR_M1006_s N_VPWR_c_422_n
+ N_VPWR_c_423_n N_VPWR_c_424_n VPWR N_VPWR_c_425_n N_VPWR_c_426_n
+ N_VPWR_c_427_n N_VPWR_c_421_n VPWR PM_SKY130_FD_SC_LP__NOR4B_2%VPWR
x_PM_SKY130_FD_SC_LP__NOR4B_2%A_229_367# N_A_229_367#_M1015_d
+ N_A_229_367#_M1017_d N_A_229_367#_M1016_d N_A_229_367#_c_485_n
+ N_A_229_367#_c_489_n N_A_229_367#_c_500_n N_A_229_367#_c_486_n
+ N_A_229_367#_c_487_n N_A_229_367#_c_504_n N_A_229_367#_c_505_n
+ N_A_229_367#_c_508_n PM_SKY130_FD_SC_LP__NOR4B_2%A_229_367#
x_PM_SKY130_FD_SC_LP__NOR4B_2%A_312_367# N_A_312_367#_M1015_s
+ N_A_312_367#_M1010_d N_A_312_367#_c_543_n
+ PM_SKY130_FD_SC_LP__NOR4B_2%A_312_367#
x_PM_SKY130_FD_SC_LP__NOR4B_2%Y N_Y_M1003_d N_Y_M1014_d N_Y_M1000_d N_Y_M1011_s
+ N_Y_M1004_s N_Y_c_563_n N_Y_c_565_n N_Y_c_566_n N_Y_c_567_n N_Y_c_568_n
+ N_Y_c_559_n N_Y_c_557_n N_Y_c_598_n N_Y_c_599_n N_Y_c_558_n N_Y_c_639_p
+ N_Y_c_578_n Y Y Y N_Y_c_561_n Y N_Y_c_562_n PM_SKY130_FD_SC_LP__NOR4B_2%Y
x_PM_SKY130_FD_SC_LP__NOR4B_2%A_672_367# N_A_672_367#_M1001_s
+ N_A_672_367#_M1013_d N_A_672_367#_c_651_n N_A_672_367#_c_652_n
+ N_A_672_367#_c_653_n PM_SKY130_FD_SC_LP__NOR4B_2%A_672_367#
x_PM_SKY130_FD_SC_LP__NOR4B_2%VGND N_VGND_M1008_d N_VGND_M1002_s N_VGND_M1009_s
+ N_VGND_M1007_d N_VGND_M1005_s N_VGND_c_675_n N_VGND_c_676_n N_VGND_c_677_n
+ N_VGND_c_678_n N_VGND_c_679_n N_VGND_c_680_n VGND N_VGND_c_681_n
+ N_VGND_c_682_n N_VGND_c_683_n N_VGND_c_684_n N_VGND_c_685_n N_VGND_c_686_n
+ N_VGND_c_687_n N_VGND_c_688_n N_VGND_c_689_n N_VGND_c_690_n VGND
+ PM_SKY130_FD_SC_LP__NOR4B_2%VGND
cc_1 VNB N_D_N_M1012_g 0.0127387f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_2 VNB N_D_N_c_90_n 0.0259489f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.185
cc_3 VNB D_N 0.0190916f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_D_N_c_92_n 0.0491873f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.35
cc_5 VNB N_C_c_116_n 0.0199427f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.515
cc_6 VNB N_C_M1015_g 0.00817268f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.865
cc_7 VNB N_C_M1017_g 0.00788071f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.35
cc_8 VNB N_C_c_119_n 0.0608465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C_c_120_n 0.010804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_C_c_121_n 0.00456254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_c_122_n 0.0317146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C_c_123_n 0.00684189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C_c_124_n 0.017698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_C_c_125_n 0.0161757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_535#_M1002_g 0.0229546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_535#_M1014_g 0.0224707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_535#_c_207_n 0.00947935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_535#_c_208_n 0.00507193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_535#_c_209_n 0.00151092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_535#_c_210_n 0.00581427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_535#_c_211_n 0.0318358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_M1000_g 0.0272465f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.865
cc_23 VNB N_B_c_292_n 0.0214535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_M1016_g 0.00860293f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.35
cc_25 VNB N_B_c_294_n 0.0093816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_c_295_n 0.00100467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB B 0.0195108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_297_n 0.0320968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B_c_298_n 0.0455495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_c_299_n 0.0016291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_c_370_n 0.016218f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.515
cc_32 VNB N_A_M1006_g 0.00649923f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.865
cc_33 VNB N_A_c_372_n 0.0162428f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_A_M1013_g 0.00688502f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.35
cc_35 VNB A 0.00713233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_c_375_n 0.0345625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_421_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_557_n 0.00507063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_558_n 0.0055464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_675_n 0.0216477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_676_n 4.10922e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_677_n 0.00564356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_678_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_679_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_680_n 0.0330576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_681_n 0.0296693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_682_n 0.0148157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_683_n 0.0167396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_684_n 0.017071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_685_n 0.012974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_686_n 0.00961405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_687_n 0.00436768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_688_n 0.00632057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_689_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_690_n 0.28401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VPB N_D_N_M1012_g 0.0880408f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_57 VPB N_C_M1015_g 0.0247941f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=0.865
cc_58 VPB N_C_M1017_g 0.0209809f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.35
cc_59 VPB N_A_27_535#_M1004_g 0.0187302f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.35
cc_60 VPB N_A_27_535#_M1010_g 0.0187183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_27_535#_c_214_n 0.0588086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_27_535#_c_208_n 9.47055e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_27_535#_c_216_n 0.0250426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_27_535#_c_217_n 0.0173185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_27_535#_c_209_n 7.75299e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_27_535#_c_211_n 0.00439329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_B_M1001_g 0.0213095f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_68 VPB N_B_M1016_g 0.0250067f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.35
cc_69 VPB N_B_c_294_n 0.00797833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_B_c_295_n 0.00407419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_B_c_297_n 0.0100807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_B_c_299_n 0.00903533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_M1006_g 0.0209403f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=0.865
cc_74 VPB N_A_M1013_g 0.0188867f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.35
cc_75 VPB N_VPWR_c_422_n 0.00826164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_423_n 0.00949009f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.35
cc_77 VPB N_VPWR_c_424_n 0.0311969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_425_n 0.0154916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_426_n 0.100667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_427_n 0.00510915f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_421_n 0.0549449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_229_367#_c_485_n 0.00752302f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.35
cc_83 VPB N_A_229_367#_c_486_n 0.0125091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_229_367#_c_487_n 0.0074629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_Y_c_559_n 0.00447594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_Y_c_557_n 0.00147222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_Y_c_561_n 0.00678215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_Y_c_562_n 0.00128371f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 N_D_N_c_92_n N_C_c_119_n 0.0186602f $X=0.475 $Y=1.35 $X2=0 $Y2=0
cc_90 N_D_N_c_90_n N_C_c_121_n 5.68741e-19 $X=0.53 $Y=1.185 $X2=0 $Y2=0
cc_91 N_D_N_c_92_n N_C_c_121_n 3.09133e-19 $X=0.475 $Y=1.35 $X2=0 $Y2=0
cc_92 N_D_N_M1012_g N_A_27_535#_c_214_n 0.0337093f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_93 N_D_N_c_90_n N_A_27_535#_c_207_n 0.0127568f $X=0.53 $Y=1.185 $X2=0 $Y2=0
cc_94 D_N N_A_27_535#_c_207_n 0.0147661f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_95 N_D_N_c_92_n N_A_27_535#_c_207_n 0.00447104f $X=0.475 $Y=1.35 $X2=0 $Y2=0
cc_96 N_D_N_M1012_g N_A_27_535#_c_208_n 0.0103854f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_97 N_D_N_c_90_n N_A_27_535#_c_208_n 0.0108102f $X=0.53 $Y=1.185 $X2=0 $Y2=0
cc_98 D_N N_A_27_535#_c_208_n 0.0231913f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_99 N_D_N_c_92_n N_A_27_535#_c_208_n 0.00904358f $X=0.475 $Y=1.35 $X2=0 $Y2=0
cc_100 N_D_N_M1012_g N_A_27_535#_c_217_n 0.0219129f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_101 D_N N_A_27_535#_c_217_n 0.0187736f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_102 N_D_N_c_92_n N_A_27_535#_c_217_n 0.00360399f $X=0.475 $Y=1.35 $X2=0 $Y2=0
cc_103 N_D_N_M1012_g N_A_27_535#_c_209_n 0.00104351f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_104 N_D_N_M1012_g N_VPWR_c_422_n 0.01261f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_105 N_D_N_M1012_g N_VPWR_c_425_n 0.00486043f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_106 N_D_N_M1012_g N_VPWR_c_421_n 0.0093594f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_107 N_D_N_M1012_g N_A_229_367#_c_487_n 0.0165118f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_108 N_D_N_c_90_n N_VGND_c_675_n 0.0103286f $X=0.53 $Y=1.185 $X2=0 $Y2=0
cc_109 N_D_N_c_90_n N_VGND_c_681_n 0.00399858f $X=0.53 $Y=1.185 $X2=0 $Y2=0
cc_110 N_D_N_c_90_n N_VGND_c_690_n 0.0046122f $X=0.53 $Y=1.185 $X2=0 $Y2=0
cc_111 N_C_c_116_n N_A_27_535#_M1002_g 0.0305173f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_112 N_C_c_125_n N_A_27_535#_M1002_g 0.010446f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_113 N_C_M1015_g N_A_27_535#_M1004_g 0.0305173f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_114 N_C_c_122_n N_A_27_535#_M1014_g 0.0207201f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_115 N_C_c_123_n N_A_27_535#_M1014_g 0.00530336f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_116 N_C_c_124_n N_A_27_535#_M1014_g 0.0146789f $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_117 N_C_c_125_n N_A_27_535#_M1014_g 0.0114971f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_118 N_C_c_119_n N_A_27_535#_c_208_n 0.00231463f $X=1.41 $Y=1.35 $X2=0 $Y2=0
cc_119 N_C_c_121_n N_A_27_535#_c_208_n 0.031508f $X=0.965 $Y=1.17 $X2=0 $Y2=0
cc_120 N_C_M1015_g N_A_27_535#_c_216_n 8.54853e-19 $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_121 N_C_c_119_n N_A_27_535#_c_216_n 0.00781199f $X=1.41 $Y=1.35 $X2=0 $Y2=0
cc_122 N_C_c_121_n N_A_27_535#_c_216_n 0.0146135f $X=0.965 $Y=1.17 $X2=0 $Y2=0
cc_123 N_C_c_125_n N_A_27_535#_c_216_n 0.006321f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_124 N_C_M1015_g N_A_27_535#_c_209_n 0.00975692f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_125 N_C_c_119_n N_A_27_535#_c_209_n 0.00833871f $X=1.41 $Y=1.35 $X2=0 $Y2=0
cc_126 N_C_c_120_n N_A_27_535#_c_209_n 3.03422e-19 $X=1.485 $Y=1.35 $X2=0 $Y2=0
cc_127 N_C_c_121_n N_A_27_535#_c_209_n 0.0059007f $X=0.965 $Y=1.17 $X2=0 $Y2=0
cc_128 N_C_c_125_n N_A_27_535#_c_209_n 0.0122704f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_129 N_C_M1015_g N_A_27_535#_c_210_n 0.00993202f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_130 N_C_M1017_g N_A_27_535#_c_210_n 6.00642e-19 $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_131 N_C_c_120_n N_A_27_535#_c_210_n 0.00483228f $X=1.485 $Y=1.35 $X2=0 $Y2=0
cc_132 N_C_c_123_n N_A_27_535#_c_210_n 0.00751423f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_133 N_C_c_125_n N_A_27_535#_c_210_n 0.0655412f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_134 N_C_M1017_g N_A_27_535#_c_211_n 0.0616026f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_135 N_C_c_120_n N_A_27_535#_c_211_n 0.0305173f $X=1.485 $Y=1.35 $X2=0 $Y2=0
cc_136 N_C_c_125_n N_A_27_535#_c_211_n 0.00246472f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_137 N_C_c_122_n N_B_M1000_g 0.00270603f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_138 N_C_c_124_n N_B_M1000_g 0.0167766f $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_139 N_C_M1017_g N_B_c_297_n 0.0354381f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_140 N_C_c_122_n N_B_c_297_n 0.00842231f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_141 N_C_M1015_g N_VPWR_c_422_n 0.00271901f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_142 N_C_M1015_g N_VPWR_c_426_n 0.00585385f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_143 N_C_M1017_g N_VPWR_c_426_n 0.00535386f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_144 N_C_M1015_g N_VPWR_c_421_n 0.0077284f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_145 N_C_M1017_g N_VPWR_c_421_n 0.00653988f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_146 N_C_M1015_g N_A_229_367#_c_489_n 0.0147f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_147 N_C_M1017_g N_A_229_367#_c_489_n 0.0114506f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_148 N_C_M1015_g N_A_229_367#_c_487_n 0.00437029f $X=1.485 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_C_c_119_n N_A_229_367#_c_487_n 7.6621e-19 $X=1.41 $Y=1.35 $X2=0 $Y2=0
cc_150 N_C_M1017_g N_A_312_367#_c_543_n 0.00473961f $X=2.775 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_C_c_116_n N_Y_c_563_n 0.00215121f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_152 N_C_c_125_n N_Y_c_563_n 0.0181602f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_153 N_C_c_116_n N_Y_c_565_n 0.00559302f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_154 N_C_c_125_n N_Y_c_566_n 0.0402256f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_155 N_C_c_124_n N_Y_c_567_n 0.0116765f $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_156 N_C_c_122_n N_Y_c_568_n 0.00227939f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_157 N_C_c_123_n N_Y_c_568_n 0.0103865f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_158 N_C_c_124_n N_Y_c_568_n 0.0100805f $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_159 N_C_M1017_g N_Y_c_559_n 0.0085509f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_160 N_C_c_122_n N_Y_c_559_n 0.0032621f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_161 N_C_M1017_g N_Y_c_557_n 0.00591549f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_162 N_C_c_122_n N_Y_c_557_n 0.00276043f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_163 N_C_c_123_n N_Y_c_557_n 0.0251002f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_164 N_C_c_123_n N_Y_c_558_n 0.00796797f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_165 N_C_c_124_n N_Y_c_558_n 0.00532954f $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_166 N_C_c_122_n N_Y_c_578_n 2.87881e-19 $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_167 N_C_c_124_n N_Y_c_578_n 7.17169e-19 $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_168 N_C_c_125_n N_Y_c_578_n 0.0194512f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_169 N_C_M1015_g N_Y_c_561_n 0.00163288f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_170 N_C_c_123_n N_Y_c_561_n 0.0207557f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_171 N_C_c_125_n N_Y_c_561_n 0.00517824f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_172 N_C_M1017_g N_Y_c_562_n 0.00934979f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_173 N_C_c_122_n N_Y_c_562_n 0.001478f $X=2.795 $Y=1.35 $X2=0 $Y2=0
cc_174 N_C_c_116_n N_VGND_c_675_n 0.0164138f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_175 N_C_c_119_n N_VGND_c_675_n 0.00303328f $X=1.41 $Y=1.35 $X2=0 $Y2=0
cc_176 N_C_c_121_n N_VGND_c_675_n 0.0175843f $X=0.965 $Y=1.17 $X2=0 $Y2=0
cc_177 N_C_c_125_n N_VGND_c_675_n 0.0242303f $X=2.49 $Y=1.3 $X2=0 $Y2=0
cc_178 N_C_c_116_n N_VGND_c_676_n 4.78045e-19 $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_179 N_C_c_124_n N_VGND_c_676_n 0.00109224f $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_180 N_C_c_124_n N_VGND_c_677_n 0.00667942f $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_181 N_C_c_116_n N_VGND_c_682_n 0.0054895f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_182 N_C_c_124_n N_VGND_c_683_n 0.00428252f $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_183 N_C_c_116_n N_VGND_c_690_n 0.011298f $X=1.485 $Y=1.185 $X2=0 $Y2=0
cc_184 N_C_c_124_n N_VGND_c_690_n 0.00674292f $X=2.795 $Y=1.185 $X2=0 $Y2=0
cc_185 N_A_27_535#_c_214_n N_VPWR_c_425_n 0.0153489f $X=0.26 $Y=2.885 $X2=0
+ $Y2=0
cc_186 N_A_27_535#_M1004_g N_VPWR_c_426_n 0.00371105f $X=1.915 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_27_535#_M1010_g N_VPWR_c_426_n 0.00371105f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_27_535#_M1012_s N_VPWR_c_421_n 0.00376753f $X=0.135 $Y=2.675 $X2=0
+ $Y2=0
cc_189 N_A_27_535#_M1004_g N_VPWR_c_421_n 0.00547858f $X=1.915 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A_27_535#_M1010_g N_VPWR_c_421_n 0.00547858f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A_27_535#_c_214_n N_VPWR_c_421_n 0.00990863f $X=0.26 $Y=2.885 $X2=0
+ $Y2=0
cc_192 N_A_27_535#_c_216_n N_A_229_367#_M1015_d 0.00126943f $X=1.245 $Y=1.78
+ $X2=-0.19 $Y2=-0.245
cc_193 N_A_27_535#_c_209_n N_A_229_367#_M1015_d 0.00124998f $X=1.415 $Y=1.53
+ $X2=-0.19 $Y2=-0.245
cc_194 N_A_27_535#_M1004_g N_A_229_367#_c_489_n 0.0104404f $X=1.915 $Y=2.465
+ $X2=0 $Y2=0
cc_195 N_A_27_535#_M1010_g N_A_229_367#_c_489_n 0.0104404f $X=2.345 $Y=2.465
+ $X2=0 $Y2=0
cc_196 N_A_27_535#_M1004_g N_A_229_367#_c_487_n 9.57644e-19 $X=1.915 $Y=2.465
+ $X2=0 $Y2=0
cc_197 N_A_27_535#_c_216_n N_A_229_367#_c_487_n 0.0114298f $X=1.245 $Y=1.78
+ $X2=0 $Y2=0
cc_198 N_A_27_535#_c_209_n N_A_229_367#_c_487_n 0.00963114f $X=1.415 $Y=1.53
+ $X2=0 $Y2=0
cc_199 N_A_27_535#_M1004_g N_A_312_367#_c_543_n 0.0129864f $X=1.915 $Y=2.465
+ $X2=0 $Y2=0
cc_200 N_A_27_535#_M1010_g N_A_312_367#_c_543_n 0.0128886f $X=2.345 $Y=2.465
+ $X2=0 $Y2=0
cc_201 N_A_27_535#_M1002_g N_Y_c_566_n 0.00993147f $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_202 N_A_27_535#_M1014_g N_Y_c_566_n 0.00993147f $X=2.345 $Y=0.655 $X2=0 $Y2=0
cc_203 N_A_27_535#_M1004_g N_Y_c_561_n 0.012546f $X=1.915 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A_27_535#_M1010_g N_Y_c_561_n 0.014514f $X=2.345 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A_27_535#_c_209_n N_Y_c_561_n 0.00331434f $X=1.415 $Y=1.53 $X2=0 $Y2=0
cc_206 N_A_27_535#_c_210_n N_Y_c_561_n 0.056631f $X=2.155 $Y=1.51 $X2=0 $Y2=0
cc_207 N_A_27_535#_c_211_n N_Y_c_561_n 0.00239121f $X=2.345 $Y=1.51 $X2=0 $Y2=0
cc_208 N_A_27_535#_c_207_n N_VGND_M1008_d 0.00597441f $X=0.525 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_209 N_A_27_535#_c_208_n N_VGND_M1008_d 0.00263273f $X=0.61 $Y=1.695 $X2=-0.19
+ $Y2=-0.245
cc_210 N_A_27_535#_c_207_n N_VGND_c_675_n 0.010356f $X=0.525 $Y=0.9 $X2=0 $Y2=0
cc_211 N_A_27_535#_M1002_g N_VGND_c_676_n 0.00796021f $X=1.915 $Y=0.655 $X2=0
+ $Y2=0
cc_212 N_A_27_535#_M1014_g N_VGND_c_676_n 0.00899467f $X=2.345 $Y=0.655 $X2=0
+ $Y2=0
cc_213 N_A_27_535#_M1002_g N_VGND_c_682_n 0.00366311f $X=1.915 $Y=0.655 $X2=0
+ $Y2=0
cc_214 N_A_27_535#_M1014_g N_VGND_c_683_n 0.00366311f $X=2.345 $Y=0.655 $X2=0
+ $Y2=0
cc_215 N_A_27_535#_M1002_g N_VGND_c_690_n 0.00436859f $X=1.915 $Y=0.655 $X2=0
+ $Y2=0
cc_216 N_A_27_535#_M1014_g N_VGND_c_690_n 0.00436859f $X=2.345 $Y=0.655 $X2=0
+ $Y2=0
cc_217 N_A_27_535#_c_207_n N_VGND_c_690_n 0.0201098f $X=0.525 $Y=0.9 $X2=0 $Y2=0
cc_218 N_B_M1000_g N_A_c_370_n 0.0208077f $X=3.515 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_219 N_B_M1001_g N_A_M1006_g 0.0294456f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_220 N_B_c_294_n N_A_M1006_g 0.0107352f $X=4.815 $Y=1.7 $X2=0 $Y2=0
cc_221 N_B_c_292_n N_A_c_372_n 0.0314439f $X=4.805 $Y=1.185 $X2=0 $Y2=0
cc_222 N_B_M1016_g N_A_M1013_g 0.0314439f $X=4.805 $Y=2.465 $X2=0 $Y2=0
cc_223 N_B_c_294_n N_A_M1013_g 0.0106984f $X=4.815 $Y=1.7 $X2=0 $Y2=0
cc_224 N_B_M1000_g A 5.32413e-19 $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_225 N_B_c_294_n A 0.05642f $X=4.815 $Y=1.7 $X2=0 $Y2=0
cc_226 N_B_c_295_n A 0.00655445f $X=3.495 $Y=1.51 $X2=0 $Y2=0
cc_227 B A 0.0198391f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_228 N_B_c_297_n A 3.64801e-19 $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_229 N_B_c_298_n A 0.00200965f $X=4.98 $Y=1.35 $X2=0 $Y2=0
cc_230 N_B_c_294_n N_A_c_375_n 0.00243542f $X=4.815 $Y=1.7 $X2=0 $Y2=0
cc_231 N_B_c_295_n N_A_c_375_n 0.00133434f $X=3.495 $Y=1.51 $X2=0 $Y2=0
cc_232 B N_A_c_375_n 0.00129495f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_233 N_B_c_297_n N_A_c_375_n 0.0219675f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_234 N_B_c_298_n N_A_c_375_n 0.0314439f $X=4.98 $Y=1.35 $X2=0 $Y2=0
cc_235 N_B_M1016_g N_VPWR_c_423_n 0.0149637f $X=4.805 $Y=2.465 $X2=0 $Y2=0
cc_236 N_B_c_299_n N_VPWR_c_423_n 3.54275e-19 $X=5.005 $Y=1.615 $X2=0 $Y2=0
cc_237 N_B_M1016_g N_VPWR_c_424_n 0.0127212f $X=4.805 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B_M1001_g N_VPWR_c_426_n 0.0054895f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B_M1016_g N_VPWR_c_426_n 0.00417534f $X=4.805 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B_M1001_g N_VPWR_c_421_n 0.0107458f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B_M1016_g N_VPWR_c_421_n 0.00682364f $X=4.805 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B_M1001_g N_A_229_367#_c_500_n 0.00680984f $X=3.285 $Y=2.465 $X2=0
+ $Y2=0
cc_243 N_B_M1016_g N_A_229_367#_c_486_n 0.011598f $X=4.805 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B_c_298_n N_A_229_367#_c_486_n 9.73221e-19 $X=4.98 $Y=1.35 $X2=0 $Y2=0
cc_245 N_B_c_299_n N_A_229_367#_c_486_n 0.0238207f $X=5.005 $Y=1.615 $X2=0 $Y2=0
cc_246 N_B_M1001_g N_A_229_367#_c_504_n 0.00486069f $X=3.285 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_B_M1001_g N_A_229_367#_c_505_n 0.0164934f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B_c_295_n N_A_229_367#_c_505_n 0.0110913f $X=3.495 $Y=1.51 $X2=0 $Y2=0
cc_249 N_B_c_297_n N_A_229_367#_c_505_n 0.00114548f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_250 N_B_M1001_g N_A_229_367#_c_508_n 0.00360326f $X=3.285 $Y=2.465 $X2=0
+ $Y2=0
cc_251 N_B_c_294_n N_A_229_367#_c_508_n 0.0620214f $X=4.815 $Y=1.7 $X2=0 $Y2=0
cc_252 N_B_c_295_n N_A_229_367#_c_508_n 9.71555e-19 $X=3.495 $Y=1.51 $X2=0 $Y2=0
cc_253 N_B_M1001_g N_Y_c_559_n 0.00664543f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_254 N_B_M1001_g N_Y_c_557_n 0.00264626f $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_255 N_B_M1000_g N_Y_c_557_n 0.00227903f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_256 N_B_c_295_n N_Y_c_557_n 0.0312303f $X=3.495 $Y=1.51 $X2=0 $Y2=0
cc_257 N_B_c_297_n N_Y_c_557_n 0.00801018f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_258 N_B_M1000_g N_Y_c_598_n 0.0120137f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_259 N_B_c_294_n N_Y_c_599_n 0.00115217f $X=4.815 $Y=1.7 $X2=0 $Y2=0
cc_260 N_B_M1000_g N_Y_c_558_n 0.0197091f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_261 N_B_c_294_n N_Y_c_558_n 0.00580735f $X=4.815 $Y=1.7 $X2=0 $Y2=0
cc_262 N_B_c_295_n N_Y_c_558_n 0.0211483f $X=3.495 $Y=1.51 $X2=0 $Y2=0
cc_263 N_B_c_297_n N_Y_c_558_n 0.00849494f $X=3.515 $Y=1.51 $X2=0 $Y2=0
cc_264 N_B_M1001_g N_Y_c_562_n 5.39933e-19 $X=3.285 $Y=2.465 $X2=0 $Y2=0
cc_265 N_B_M1001_g N_A_672_367#_c_651_n 0.00263789f $X=3.285 $Y=2.465 $X2=0
+ $Y2=0
cc_266 N_B_M1001_g N_A_672_367#_c_652_n 0.00359192f $X=3.285 $Y=2.465 $X2=0
+ $Y2=0
cc_267 N_B_M1016_g N_A_672_367#_c_653_n 0.00314718f $X=4.805 $Y=2.465 $X2=0
+ $Y2=0
cc_268 N_B_M1000_g N_VGND_c_677_n 0.00676345f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_269 N_B_M1000_g N_VGND_c_678_n 0.00124765f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_270 N_B_c_292_n N_VGND_c_678_n 5.80819e-19 $X=4.805 $Y=1.185 $X2=0 $Y2=0
cc_271 N_B_c_292_n N_VGND_c_680_n 0.0163657f $X=4.805 $Y=1.185 $X2=0 $Y2=0
cc_272 B N_VGND_c_680_n 0.0259713f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_273 N_B_c_298_n N_VGND_c_680_n 0.00192467f $X=4.98 $Y=1.35 $X2=0 $Y2=0
cc_274 N_B_M1000_g N_VGND_c_684_n 0.0042814f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_275 N_B_c_292_n N_VGND_c_685_n 0.00486043f $X=4.805 $Y=1.185 $X2=0 $Y2=0
cc_276 N_B_M1000_g N_VGND_c_690_n 0.00674084f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_277 N_B_c_292_n N_VGND_c_690_n 0.0082726f $X=4.805 $Y=1.185 $X2=0 $Y2=0
cc_278 N_A_M1006_g N_VPWR_c_423_n 0.00345464f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_279 N_A_M1013_g N_VPWR_c_423_n 0.00944188f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_280 N_A_M1006_g N_VPWR_c_426_n 0.00357877f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_281 N_A_M1013_g N_VPWR_c_426_n 0.00357877f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_282 N_A_M1006_g N_VPWR_c_421_n 0.00594089f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_283 N_A_M1013_g N_VPWR_c_421_n 0.00537654f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_284 N_A_M1006_g N_A_229_367#_c_486_n 0.0176599f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_285 N_A_M1013_g N_A_229_367#_c_486_n 0.0149546f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A_M1006_g N_A_229_367#_c_504_n 8.79421e-19 $X=3.945 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_A_M1006_g N_Y_c_559_n 7.27507e-19 $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_288 A N_Y_c_557_n 0.00384127f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_289 N_A_c_370_n N_Y_c_599_n 0.0122129f $X=3.945 $Y=1.185 $X2=0 $Y2=0
cc_290 N_A_c_372_n N_Y_c_599_n 0.0122595f $X=4.375 $Y=1.185 $X2=0 $Y2=0
cc_291 A N_Y_c_599_n 0.0507175f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_292 N_A_c_375_n N_Y_c_599_n 0.00230884f $X=4.375 $Y=1.35 $X2=0 $Y2=0
cc_293 N_A_c_370_n N_Y_c_558_n 0.00353079f $X=3.945 $Y=1.185 $X2=0 $Y2=0
cc_294 N_A_M1006_g N_A_672_367#_c_652_n 0.00661539f $X=3.945 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_M1006_g N_A_672_367#_c_653_n 0.0150609f $X=3.945 $Y=2.465 $X2=0 $Y2=0
cc_296 N_A_M1013_g N_A_672_367#_c_653_n 0.0095355f $X=4.375 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A_c_370_n N_VGND_c_678_n 0.011763f $X=3.945 $Y=1.185 $X2=0 $Y2=0
cc_298 N_A_c_372_n N_VGND_c_678_n 0.0106438f $X=4.375 $Y=1.185 $X2=0 $Y2=0
cc_299 N_A_c_372_n N_VGND_c_680_n 6.29195e-19 $X=4.375 $Y=1.185 $X2=0 $Y2=0
cc_300 N_A_c_370_n N_VGND_c_684_n 0.00486043f $X=3.945 $Y=1.185 $X2=0 $Y2=0
cc_301 N_A_c_372_n N_VGND_c_685_n 0.00486043f $X=4.375 $Y=1.185 $X2=0 $Y2=0
cc_302 N_A_c_370_n N_VGND_c_690_n 0.0082726f $X=3.945 $Y=1.185 $X2=0 $Y2=0
cc_303 N_A_c_372_n N_VGND_c_690_n 0.0082726f $X=4.375 $Y=1.185 $X2=0 $Y2=0
cc_304 N_VPWR_c_421_n N_A_229_367#_M1015_d 0.00215158f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_305 N_VPWR_c_421_n N_A_229_367#_M1017_d 0.00324785f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_423_n N_A_229_367#_M1016_d 0.00329544f $X=4.935 $Y=2.56 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_424_n N_A_229_367#_M1016_d 0.00372718f $X=5.065 $Y=3.245 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_421_n N_A_229_367#_M1016_d 6.51481e-19 $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_422_n N_A_229_367#_c_485_n 0.0224616f $X=0.69 $Y=2.885 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_426_n N_A_229_367#_c_485_n 0.0193729f $X=4.935 $Y=3.33 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_421_n N_A_229_367#_c_485_n 0.0117747f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_421_n N_A_229_367#_c_489_n 0.011165f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_313 N_VPWR_c_426_n N_A_229_367#_c_500_n 0.0209582f $X=4.935 $Y=3.33 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_421_n N_A_229_367#_c_500_n 0.0125636f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_315 N_VPWR_M1006_s N_A_229_367#_c_486_n 0.00366015f $X=4.02 $Y=1.835 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_423_n N_A_229_367#_c_486_n 0.0696091f $X=4.935 $Y=2.56 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_421_n N_A_312_367#_M1015_s 0.0024313f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_318 N_VPWR_c_421_n N_A_312_367#_M1010_d 0.00230064f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_426_n N_A_312_367#_c_543_n 0.0468076f $X=4.935 $Y=3.33 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_421_n N_A_312_367#_c_543_n 0.0409108f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_421_n N_Y_M1004_s 0.00230064f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_322 N_VPWR_c_421_n N_A_672_367#_M1001_s 0.00693476f $X=5.04 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_323 N_VPWR_c_423_n N_A_672_367#_M1013_d 0.00350091f $X=4.935 $Y=2.56 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_421_n N_A_672_367#_M1013_d 0.00223577f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_426_n N_A_672_367#_c_651_n 0.0229651f $X=4.935 $Y=3.33 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_421_n N_A_672_367#_c_651_n 0.0127825f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_423_n N_A_672_367#_c_652_n 0.0118737f $X=4.935 $Y=2.56 $X2=0
+ $Y2=0
cc_328 N_VPWR_M1006_s N_A_672_367#_c_653_n 0.00336331f $X=4.02 $Y=1.835 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_423_n N_A_672_367#_c_653_n 0.0373318f $X=4.935 $Y=2.56 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_426_n N_A_672_367#_c_653_n 0.0547501f $X=4.935 $Y=3.33 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_421_n N_A_672_367#_c_653_n 0.0356838f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_332 N_A_229_367#_c_489_n N_A_312_367#_M1015_s 0.00351441f $X=2.905 $Y=2.4
+ $X2=-0.19 $Y2=1.655
cc_333 N_A_229_367#_c_489_n N_A_312_367#_M1010_d 0.00351441f $X=2.905 $Y=2.4
+ $X2=0 $Y2=0
cc_334 N_A_229_367#_c_489_n N_A_312_367#_c_543_n 0.060791f $X=2.905 $Y=2.4 $X2=0
+ $Y2=0
cc_335 N_A_229_367#_c_489_n N_Y_M1004_s 0.00343263f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_336 N_A_229_367#_M1017_d N_Y_c_559_n 0.00264495f $X=2.85 $Y=1.835 $X2=0 $Y2=0
cc_337 N_A_229_367#_c_489_n N_Y_c_559_n 0.0044528f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_338 N_A_229_367#_c_504_n N_Y_c_559_n 0.0224048f $X=3.07 $Y=2.23 $X2=0 $Y2=0
cc_339 N_A_229_367#_c_489_n N_Y_c_561_n 0.0620124f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_340 N_A_229_367#_c_505_n N_A_672_367#_M1001_s 0.00697751f $X=3.645 $Y=2.16
+ $X2=-0.19 $Y2=1.655
cc_341 N_A_229_367#_c_508_n N_A_672_367#_M1001_s 0.00700284f $X=3.815 $Y=2.16
+ $X2=-0.19 $Y2=1.655
cc_342 N_A_229_367#_c_486_n N_A_672_367#_M1013_d 0.00380671f $X=5.02 $Y=2.17
+ $X2=0 $Y2=0
cc_343 N_A_229_367#_c_500_n N_A_672_367#_c_651_n 0.0171513f $X=3.07 $Y=2.6 $X2=0
+ $Y2=0
cc_344 N_A_229_367#_c_500_n N_A_672_367#_c_652_n 0.0234565f $X=3.07 $Y=2.6 $X2=0
+ $Y2=0
cc_345 N_A_229_367#_c_505_n N_A_672_367#_c_652_n 0.0267679f $X=3.645 $Y=2.16
+ $X2=0 $Y2=0
cc_346 N_A_229_367#_c_486_n N_A_672_367#_c_653_n 0.00344783f $X=5.02 $Y=2.17
+ $X2=0 $Y2=0
cc_347 N_A_229_367#_c_508_n N_A_672_367#_c_653_n 0.00144624f $X=3.815 $Y=2.16
+ $X2=0 $Y2=0
cc_348 N_A_312_367#_c_543_n N_Y_M1004_s 0.0036349f $X=2.56 $Y=2.82 $X2=1.485
+ $Y2=2.465
cc_349 N_A_312_367#_M1015_s N_Y_c_561_n 0.00252346f $X=1.56 $Y=1.835 $X2=0 $Y2=0
cc_350 N_A_312_367#_M1010_d N_Y_c_561_n 9.47075e-19 $X=2.42 $Y=1.835 $X2=0 $Y2=0
cc_351 N_A_312_367#_M1010_d N_Y_c_562_n 8.49102e-19 $X=2.42 $Y=1.835 $X2=0 $Y2=0
cc_352 N_Y_c_566_n N_VGND_M1002_s 0.00335318f $X=2.465 $Y=0.83 $X2=0 $Y2=0
cc_353 N_Y_c_568_n N_VGND_M1009_s 0.0069943f $X=3.06 $Y=0.83 $X2=0 $Y2=0
cc_354 N_Y_c_558_n N_VGND_M1009_s 0.0100133f $X=3.825 $Y=0.955 $X2=0 $Y2=0
cc_355 N_Y_c_599_n N_VGND_M1007_d 0.00329816f $X=4.495 $Y=0.955 $X2=0 $Y2=0
cc_356 N_Y_c_566_n N_VGND_c_676_n 0.0165001f $X=2.465 $Y=0.83 $X2=0 $Y2=0
cc_357 N_Y_c_567_n N_VGND_c_677_n 0.0176269f $X=2.56 $Y=0.42 $X2=0 $Y2=0
cc_358 N_Y_c_568_n N_VGND_c_677_n 0.00578381f $X=3.06 $Y=0.83 $X2=0 $Y2=0
cc_359 N_Y_c_598_n N_VGND_c_677_n 0.0181626f $X=3.73 $Y=0.42 $X2=0 $Y2=0
cc_360 N_Y_c_558_n N_VGND_c_677_n 0.0218303f $X=3.825 $Y=0.955 $X2=0 $Y2=0
cc_361 N_Y_c_599_n N_VGND_c_678_n 0.0170777f $X=4.495 $Y=0.955 $X2=0 $Y2=0
cc_362 N_Y_c_565_n N_VGND_c_682_n 0.0156591f $X=1.7 $Y=0.42 $X2=0 $Y2=0
cc_363 N_Y_c_566_n N_VGND_c_682_n 0.00191958f $X=2.465 $Y=0.83 $X2=0 $Y2=0
cc_364 N_Y_c_566_n N_VGND_c_683_n 0.00191958f $X=2.465 $Y=0.83 $X2=0 $Y2=0
cc_365 N_Y_c_567_n N_VGND_c_683_n 0.0156591f $X=2.56 $Y=0.42 $X2=0 $Y2=0
cc_366 N_Y_c_568_n N_VGND_c_683_n 0.00309081f $X=3.06 $Y=0.83 $X2=0 $Y2=0
cc_367 N_Y_c_598_n N_VGND_c_684_n 0.015688f $X=3.73 $Y=0.42 $X2=0 $Y2=0
cc_368 N_Y_c_558_n N_VGND_c_684_n 0.00313464f $X=3.825 $Y=0.955 $X2=0 $Y2=0
cc_369 N_Y_c_639_p N_VGND_c_685_n 0.0117038f $X=4.59 $Y=0.43 $X2=0 $Y2=0
cc_370 N_Y_M1003_d N_VGND_c_690_n 0.00245675f $X=1.56 $Y=0.235 $X2=0 $Y2=0
cc_371 N_Y_M1014_d N_VGND_c_690_n 0.00245675f $X=2.42 $Y=0.235 $X2=0 $Y2=0
cc_372 N_Y_M1000_d N_VGND_c_690_n 0.00380103f $X=3.59 $Y=0.235 $X2=0 $Y2=0
cc_373 N_Y_M1011_s N_VGND_c_690_n 0.00536823f $X=4.45 $Y=0.235 $X2=0 $Y2=0
cc_374 N_Y_c_565_n N_VGND_c_690_n 0.00983963f $X=1.7 $Y=0.42 $X2=0 $Y2=0
cc_375 N_Y_c_566_n N_VGND_c_690_n 0.00882814f $X=2.465 $Y=0.83 $X2=0 $Y2=0
cc_376 N_Y_c_567_n N_VGND_c_690_n 0.00983963f $X=2.56 $Y=0.42 $X2=0 $Y2=0
cc_377 N_Y_c_568_n N_VGND_c_690_n 0.0065039f $X=3.06 $Y=0.83 $X2=0 $Y2=0
cc_378 N_Y_c_598_n N_VGND_c_690_n 0.00984745f $X=3.73 $Y=0.42 $X2=0 $Y2=0
cc_379 N_Y_c_558_n N_VGND_c_690_n 0.00729747f $X=3.825 $Y=0.955 $X2=0 $Y2=0
cc_380 N_Y_c_639_p N_VGND_c_690_n 0.00727431f $X=4.59 $Y=0.43 $X2=0 $Y2=0
