# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlybuf4s15kapwr_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlybuf4s15kapwr_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.550000 1.860000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.445200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.210000 0.310000 3.750000 0.640000 ;
        RECT 3.230000 1.815000 3.750000 3.075000 ;
        RECT 3.515000 0.640000 3.750000 1.815000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.595000 2.380000 0.925000 3.075000 ;
        RECT 2.710000 2.165000 3.040000 3.075000 ;
      LAYER mcon ;
        RECT 0.675000 2.725000 0.845000 2.895000 ;
        RECT 2.790000 2.725000 2.960000 2.895000 ;
      LAYER met1 ;
        RECT 0.070000 2.690000 3.770000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
        RECT 0.580000  0.085000 0.910000 0.650000 ;
        RECT 2.710000  0.085000 3.040000 0.670000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 3.840000 3.415000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.305000 0.410000 0.820000 ;
      RECT 0.095000 0.820000 1.265000 1.020000 ;
      RECT 0.095000 2.030000 1.265000 2.205000 ;
      RECT 0.095000 2.205000 0.425000 3.075000 ;
      RECT 0.910000 1.020000 1.265000 1.600000 ;
      RECT 0.910000 1.600000 1.500000 1.930000 ;
      RECT 0.910000 1.930000 1.265000 2.030000 ;
      RECT 1.385000 2.395000 1.840000 3.075000 ;
      RECT 1.435000 0.270000 1.840000 1.280000 ;
      RECT 1.445000 2.100000 1.840000 2.395000 ;
      RECT 1.670000 1.280000 1.840000 1.385000 ;
      RECT 1.670000 1.385000 2.685000 1.655000 ;
      RECT 1.670000 1.655000 1.840000 2.100000 ;
      RECT 2.010000 0.270000 2.260000 0.980000 ;
      RECT 2.010000 0.980000 3.025000 1.215000 ;
      RECT 2.010000 2.080000 2.540000 2.250000 ;
      RECT 2.010000 2.250000 2.260000 3.075000 ;
      RECT 2.370000 1.825000 3.025000 1.995000 ;
      RECT 2.370000 1.995000 2.540000 2.080000 ;
      RECT 2.855000 1.215000 3.025000 1.295000 ;
      RECT 2.855000 1.295000 3.345000 1.625000 ;
      RECT 2.855000 1.625000 3.025000 1.825000 ;
  END
END sky130_fd_sc_lp__dlybuf4s15kapwr_1
