* File: sky130_fd_sc_lp__nand2b_2.pxi.spice
* Created: Fri Aug 28 10:48:12 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2B_2%A_N N_A_N_c_53_n N_A_N_M1008_g N_A_N_c_54_n
+ N_A_N_M1001_g A_N PM_SKY130_FD_SC_LP__NAND2B_2%A_N
x_PM_SKY130_FD_SC_LP__NAND2B_2%B N_B_M1000_g N_B_M1002_g N_B_M1009_g N_B_M1007_g
+ N_B_c_84_n N_B_c_85_n N_B_c_86_n B N_B_c_87_n N_B_c_88_n N_B_c_89_n N_B_c_90_n
+ PM_SKY130_FD_SC_LP__NAND2B_2%B
x_PM_SKY130_FD_SC_LP__NAND2B_2%A_27_131# N_A_27_131#_M1008_s N_A_27_131#_M1001_s
+ N_A_27_131#_M1003_g N_A_27_131#_M1004_g N_A_27_131#_M1005_g
+ N_A_27_131#_M1006_g N_A_27_131#_c_167_n N_A_27_131#_c_162_n
+ N_A_27_131#_c_168_n N_A_27_131#_c_163_n N_A_27_131#_c_170_n
+ N_A_27_131#_c_164_n PM_SKY130_FD_SC_LP__NAND2B_2%A_27_131#
x_PM_SKY130_FD_SC_LP__NAND2B_2%VPWR N_VPWR_M1001_d N_VPWR_M1004_d N_VPWR_M1007_d
+ N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n VPWR
+ N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_234_n N_VPWR_c_242_n N_VPWR_c_243_n
+ N_VPWR_c_244_n PM_SKY130_FD_SC_LP__NAND2B_2%VPWR
x_PM_SKY130_FD_SC_LP__NAND2B_2%Y N_Y_M1003_d N_Y_M1002_s N_Y_M1006_s N_Y_c_293_n
+ N_Y_c_306_n N_Y_c_274_n N_Y_c_308_n N_Y_c_275_n N_Y_c_286_n Y Y Y N_Y_c_277_n
+ N_Y_c_296_n N_Y_c_278_n PM_SKY130_FD_SC_LP__NAND2B_2%Y
x_PM_SKY130_FD_SC_LP__NAND2B_2%VGND N_VGND_M1008_d N_VGND_M1009_d N_VGND_c_332_n
+ N_VGND_c_324_n N_VGND_c_325_n VGND N_VGND_c_326_n N_VGND_c_327_n
+ N_VGND_c_328_n N_VGND_c_329_n N_VGND_c_330_n N_VGND_c_331_n
+ PM_SKY130_FD_SC_LP__NAND2B_2%VGND
x_PM_SKY130_FD_SC_LP__NAND2B_2%A_229_47# N_A_229_47#_M1000_s N_A_229_47#_M1005_s
+ N_A_229_47#_c_366_n N_A_229_47#_c_367_n N_A_229_47#_c_371_n
+ PM_SKY130_FD_SC_LP__NAND2B_2%A_229_47#
cc_1 VNB N_A_N_c_53_n 0.0220883f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_A_N_c_54_n 0.0340998f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.515
cc_3 VNB N_A_N_M1001_g 0.00871108f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.045
cc_4 VNB A_N 0.00471009f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_B_M1002_g 0.00780581f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.045
cc_6 VNB N_B_M1007_g 0.00811201f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.35
cc_7 VNB N_B_c_84_n 0.0187618f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_8 VNB N_B_c_85_n 0.00316584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B_c_86_n 0.0355322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_87_n 0.0316047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_88_n 0.0196613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_c_89_n 0.0196625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_90_n 0.00399605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_131#_M1003_g 0.023619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_131#_M1005_g 0.023679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_131#_c_162_n 0.0132059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_131#_c_163_n 0.0302778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_131#_c_164_n 0.0374788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_234_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_274_n 0.0208582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_275_n 0.046278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_324_n 0.0175498f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.35
cc_23 VNB N_VGND_c_325_n 0.0173644f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.35
cc_24 VNB N_VGND_c_326_n 0.017784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_327_n 0.0381222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_328_n 0.0176385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_329_n 0.199796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_330_n 0.00817107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_331_n 0.00497021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_A_N_M1001_g 0.0290214f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.045
cc_31 VPB N_B_M1002_g 0.0220541f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.045
cc_32 VPB N_B_M1007_g 0.0231284f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.35
cc_33 VPB N_A_27_131#_M1004_g 0.0172018f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.35
cc_34 VPB N_A_27_131#_M1006_g 0.0187408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_27_131#_c_167_n 0.00949618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A_27_131#_c_168_n 0.0361166f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_27_131#_c_163_n 0.00199429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_27_131#_c_170_n 0.00209803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_131#_c_164_n 0.00725013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_235_n 0.0346281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_236_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_237_n 3.16049e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_238_n 0.0340406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_239_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_240_n 0.0193272f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_234_n 0.0861051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_242_n 0.0310026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_243_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_244_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_Y_c_275_n 0.0436895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_Y_c_277_n 0.0121397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_Y_c_278_n 0.0033961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 N_A_N_M1001_g N_B_M1002_g 0.0213891f $X=0.625 $Y=2.045 $X2=0 $Y2=0
cc_54 N_A_N_c_54_n N_B_c_87_n 0.0176596f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_55 A_N N_B_c_87_n 0.00234853f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_56 N_A_N_c_53_n N_B_c_88_n 0.00993698f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_57 N_A_N_c_53_n N_B_c_90_n 5.91657e-19 $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_58 N_A_N_c_54_n N_B_c_90_n 2.80441e-19 $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_59 A_N N_B_c_90_n 0.0262432f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_60 N_A_N_c_54_n N_A_27_131#_c_167_n 0.00117784f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_61 N_A_N_M1001_g N_A_27_131#_c_167_n 0.0148069f $X=0.625 $Y=2.045 $X2=0 $Y2=0
cc_62 A_N N_A_27_131#_c_167_n 0.0241331f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A_N_c_54_n N_A_27_131#_c_168_n 0.00525075f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_64 N_A_N_M1001_g N_A_27_131#_c_168_n 0.00151602f $X=0.625 $Y=2.045 $X2=0
+ $Y2=0
cc_65 A_N N_A_27_131#_c_168_n 0.00505266f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A_N_c_53_n N_A_27_131#_c_163_n 0.00547137f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_67 N_A_N_c_54_n N_A_27_131#_c_163_n 0.0081318f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_68 N_A_N_M1001_g N_A_27_131#_c_163_n 0.00539031f $X=0.625 $Y=2.045 $X2=0
+ $Y2=0
cc_69 A_N N_A_27_131#_c_163_n 0.0240707f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A_N_M1001_g N_VPWR_c_235_n 0.012245f $X=0.625 $Y=2.045 $X2=0 $Y2=0
cc_71 N_A_N_c_53_n N_VGND_c_332_n 0.00357562f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_72 N_A_N_c_54_n N_VGND_c_332_n 0.00363588f $X=0.625 $Y=1.515 $X2=0 $Y2=0
cc_73 A_N N_VGND_c_332_n 0.0219939f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_N_c_53_n N_VGND_c_324_n 0.00975614f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_75 N_A_N_c_53_n N_VGND_c_326_n 0.00332367f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_76 N_A_N_c_53_n N_VGND_c_329_n 0.00387424f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_77 N_B_c_84_n N_A_27_131#_M1003_g 0.0120029f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B_c_87_n N_A_27_131#_M1003_g 0.0209638f $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_79 N_B_c_88_n N_A_27_131#_M1003_g 0.0139011f $X=1.095 $Y=1.185 $X2=0 $Y2=0
cc_80 N_B_c_90_n N_A_27_131#_M1003_g 0.00464285f $X=1.155 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B_M1002_g N_A_27_131#_M1004_g 0.0221076f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_82 N_B_c_84_n N_A_27_131#_M1005_g 0.0131899f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_83 N_B_c_85_n N_A_27_131#_M1005_g 7.40643e-19 $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B_c_89_n N_A_27_131#_M1005_g 0.0429482f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_85 N_B_M1007_g N_A_27_131#_M1006_g 0.018833f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_86 N_B_M1002_g N_A_27_131#_c_167_n 0.0151631f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_87 N_B_c_84_n N_A_27_131#_c_167_n 0.00653336f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_88 N_B_c_87_n N_A_27_131#_c_167_n 0.003756f $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_89 N_B_c_90_n N_A_27_131#_c_167_n 0.0208968f $X=1.155 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B_M1002_g N_A_27_131#_c_170_n 0.00160719f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B_c_84_n N_A_27_131#_c_170_n 0.0248146f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_92 N_B_c_85_n N_A_27_131#_c_170_n 0.00279025f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B_c_86_n N_A_27_131#_c_170_n 7.56781e-19 $X=2.53 $Y=1.35 $X2=0 $Y2=0
cc_94 N_B_c_90_n N_A_27_131#_c_170_n 0.00783335f $X=1.155 $Y=1.16 $X2=0 $Y2=0
cc_95 N_B_M1002_g N_A_27_131#_c_164_n 0.00931265f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_96 N_B_c_84_n N_A_27_131#_c_164_n 0.00578226f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B_c_85_n N_A_27_131#_c_164_n 0.0010181f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_98 N_B_c_86_n N_A_27_131#_c_164_n 0.0215874f $X=2.53 $Y=1.35 $X2=0 $Y2=0
cc_99 N_B_M1002_g N_VPWR_c_235_n 0.00554853f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_100 N_B_M1002_g N_VPWR_c_236_n 0.00585385f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_101 N_B_M1002_g N_VPWR_c_237_n 6.64182e-19 $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_102 N_B_M1007_g N_VPWR_c_237_n 6.47957e-19 $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_103 N_B_M1007_g N_VPWR_c_238_n 0.0163543f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_104 N_B_M1007_g N_VPWR_c_239_n 0.00486043f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_105 N_B_M1002_g N_VPWR_c_234_n 0.0118611f $X=1.15 $Y=2.465 $X2=0 $Y2=0
cc_106 N_B_M1007_g N_VPWR_c_234_n 0.0082726f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_107 N_B_c_85_n N_Y_c_274_n 0.0230126f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_108 N_B_c_86_n N_Y_c_274_n 8.54812e-19 $X=2.53 $Y=1.35 $X2=0 $Y2=0
cc_109 N_B_c_89_n N_Y_c_274_n 0.0144913f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_110 N_B_M1007_g N_Y_c_275_n 0.00975236f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_111 N_B_c_85_n N_Y_c_275_n 0.0343353f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_112 N_B_c_86_n N_Y_c_275_n 0.00751394f $X=2.53 $Y=1.35 $X2=0 $Y2=0
cc_113 N_B_c_89_n N_Y_c_275_n 0.00580904f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_114 N_B_c_84_n N_Y_c_286_n 0.0460258f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_115 N_B_c_89_n N_Y_c_286_n 3.37063e-19 $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_116 N_B_M1007_g N_Y_c_277_n 0.0200375f $X=2.44 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B_c_85_n N_Y_c_277_n 0.0160051f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_118 N_B_c_86_n N_Y_c_277_n 0.00117498f $X=2.53 $Y=1.35 $X2=0 $Y2=0
cc_119 N_B_c_84_n N_Y_c_278_n 0.0124255f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B_c_85_n N_VGND_M1009_d 0.00195953f $X=2.53 $Y=1.16 $X2=0 $Y2=0
cc_121 N_B_c_87_n N_VGND_c_332_n 5.32026e-19 $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_122 N_B_c_88_n N_VGND_c_332_n 0.00235903f $X=1.095 $Y=1.185 $X2=0 $Y2=0
cc_123 N_B_c_88_n N_VGND_c_324_n 0.00549395f $X=1.095 $Y=1.185 $X2=0 $Y2=0
cc_124 N_B_c_89_n N_VGND_c_325_n 0.00459147f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_125 N_B_c_88_n N_VGND_c_327_n 0.00547432f $X=1.095 $Y=1.185 $X2=0 $Y2=0
cc_126 N_B_c_89_n N_VGND_c_327_n 0.00424523f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_127 N_B_c_88_n N_VGND_c_329_n 0.0111586f $X=1.095 $Y=1.185 $X2=0 $Y2=0
cc_128 N_B_c_89_n N_VGND_c_329_n 0.00713961f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_129 N_B_c_90_n N_A_229_47#_M1000_s 0.00168172f $X=1.155 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_130 N_B_c_88_n N_A_229_47#_c_366_n 0.00265698f $X=1.095 $Y=1.185 $X2=0 $Y2=0
cc_131 N_B_c_84_n N_A_229_47#_c_367_n 0.0106712f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_132 N_B_c_87_n N_A_229_47#_c_367_n 5.43363e-19 $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_133 N_B_c_88_n N_A_229_47#_c_367_n 0.00525137f $X=1.095 $Y=1.185 $X2=0 $Y2=0
cc_134 N_B_c_90_n N_A_229_47#_c_367_n 0.0127696f $X=1.155 $Y=1.16 $X2=0 $Y2=0
cc_135 N_B_c_84_n N_A_229_47#_c_371_n 0.00418809f $X=2.365 $Y=1.16 $X2=0 $Y2=0
cc_136 N_B_c_89_n N_A_229_47#_c_371_n 0.00304519f $X=2.53 $Y=1.185 $X2=0 $Y2=0
cc_137 N_A_27_131#_c_167_n N_VPWR_M1001_d 0.00279856f $X=1.47 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_27_131#_c_170_n N_VPWR_M1004_d 0.00120595f $X=1.635 $Y=1.51 $X2=0
+ $Y2=0
cc_139 N_A_27_131#_c_167_n N_VPWR_c_235_n 0.0230207f $X=1.47 $Y=1.78 $X2=0 $Y2=0
cc_140 N_A_27_131#_M1004_g N_VPWR_c_236_n 0.00486043f $X=1.58 $Y=2.465 $X2=0
+ $Y2=0
cc_141 N_A_27_131#_M1004_g N_VPWR_c_237_n 0.0123843f $X=1.58 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_27_131#_M1006_g N_VPWR_c_237_n 0.0122924f $X=2.01 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_27_131#_M1006_g N_VPWR_c_238_n 6.72004e-19 $X=2.01 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_27_131#_M1006_g N_VPWR_c_239_n 0.00486043f $X=2.01 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_27_131#_M1004_g N_VPWR_c_234_n 0.0082726f $X=1.58 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_27_131#_M1006_g N_VPWR_c_234_n 0.0082726f $X=2.01 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_27_131#_c_167_n N_Y_M1002_s 0.00176461f $X=1.47 $Y=1.78 $X2=0 $Y2=0
cc_148 N_A_27_131#_c_167_n N_Y_c_293_n 0.0135055f $X=1.47 $Y=1.78 $X2=0 $Y2=0
cc_149 N_A_27_131#_M1005_g N_Y_c_274_n 0.00788184f $X=2.01 $Y=0.655 $X2=0 $Y2=0
cc_150 N_A_27_131#_M1005_g N_Y_c_286_n 0.00233574f $X=2.01 $Y=0.655 $X2=0 $Y2=0
cc_151 N_A_27_131#_M1004_g N_Y_c_296_n 0.01223f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_27_131#_M1006_g N_Y_c_296_n 0.00477152f $X=2.01 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_27_131#_c_170_n N_Y_c_296_n 0.0178538f $X=1.635 $Y=1.51 $X2=0 $Y2=0
cc_154 N_A_27_131#_c_164_n N_Y_c_296_n 0.00165473f $X=2.01 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A_27_131#_M1004_g N_Y_c_278_n 0.0010124f $X=1.58 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A_27_131#_M1006_g N_Y_c_278_n 0.0157648f $X=2.01 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_27_131#_c_170_n N_Y_c_278_n 0.00280776f $X=1.635 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A_27_131#_c_164_n N_Y_c_278_n 0.00156561f $X=2.01 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A_27_131#_c_162_n N_VGND_c_326_n 0.00429694f $X=0.26 $Y=0.85 $X2=0
+ $Y2=0
cc_160 N_A_27_131#_M1003_g N_VGND_c_327_n 0.00357877f $X=1.545 $Y=0.655 $X2=0
+ $Y2=0
cc_161 N_A_27_131#_M1005_g N_VGND_c_327_n 0.00357877f $X=2.01 $Y=0.655 $X2=0
+ $Y2=0
cc_162 N_A_27_131#_M1003_g N_VGND_c_329_n 0.00557672f $X=1.545 $Y=0.655 $X2=0
+ $Y2=0
cc_163 N_A_27_131#_M1005_g N_VGND_c_329_n 0.00547177f $X=2.01 $Y=0.655 $X2=0
+ $Y2=0
cc_164 N_A_27_131#_c_162_n N_VGND_c_329_n 0.00748852f $X=0.26 $Y=0.85 $X2=0
+ $Y2=0
cc_165 N_A_27_131#_M1003_g N_A_229_47#_c_371_n 0.0115727f $X=1.545 $Y=0.655
+ $X2=0 $Y2=0
cc_166 N_A_27_131#_M1005_g N_A_229_47#_c_371_n 0.00989781f $X=2.01 $Y=0.655
+ $X2=0 $Y2=0
cc_167 N_VPWR_c_234_n N_Y_M1002_s 0.00397496f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_168 N_VPWR_c_234_n N_Y_M1006_s 0.00536646f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_169 N_VPWR_c_236_n N_Y_c_306_n 0.0138717f $X=1.63 $Y=3.33 $X2=0 $Y2=0
cc_170 N_VPWR_c_234_n N_Y_c_306_n 0.00886411f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_171 N_VPWR_c_239_n N_Y_c_308_n 0.0124525f $X=2.49 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_234_n N_Y_c_308_n 0.00730901f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_173 N_VPWR_M1007_d N_Y_c_277_n 0.0035839f $X=2.515 $Y=1.835 $X2=0 $Y2=0
cc_174 N_VPWR_c_238_n N_Y_c_277_n 0.0228284f $X=2.655 $Y=2.41 $X2=0 $Y2=0
cc_175 N_VPWR_M1004_d N_Y_c_296_n 0.00448436f $X=1.655 $Y=1.835 $X2=0 $Y2=0
cc_176 N_VPWR_c_237_n N_Y_c_296_n 0.0170777f $X=1.795 $Y=2.485 $X2=0 $Y2=0
cc_177 N_Y_c_274_n N_VGND_M1009_d 0.00736545f $X=2.875 $Y=0.815 $X2=0 $Y2=0
cc_178 N_Y_c_274_n N_VGND_c_325_n 0.0195099f $X=2.875 $Y=0.815 $X2=0 $Y2=0
cc_179 N_Y_c_274_n N_VGND_c_327_n 0.00201765f $X=2.875 $Y=0.815 $X2=0 $Y2=0
cc_180 N_Y_c_274_n N_VGND_c_328_n 0.00761636f $X=2.875 $Y=0.815 $X2=0 $Y2=0
cc_181 N_Y_M1003_d N_VGND_c_329_n 0.00253334f $X=1.62 $Y=0.235 $X2=0 $Y2=0
cc_182 N_Y_c_274_n N_VGND_c_329_n 0.0186652f $X=2.875 $Y=0.815 $X2=0 $Y2=0
cc_183 N_Y_c_274_n N_A_229_47#_M1005_s 0.00377356f $X=2.875 $Y=0.815 $X2=0 $Y2=0
cc_184 N_Y_M1003_d N_A_229_47#_c_371_n 0.0040671f $X=1.62 $Y=0.235 $X2=0 $Y2=0
cc_185 N_Y_c_274_n N_A_229_47#_c_371_n 0.0160872f $X=2.875 $Y=0.815 $X2=0 $Y2=0
cc_186 N_Y_c_286_n N_A_229_47#_c_371_n 0.0162882f $X=1.96 $Y=0.78 $X2=0 $Y2=0
cc_187 N_VGND_c_329_n N_A_229_47#_M1000_s 0.00259748f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_188 N_VGND_c_329_n N_A_229_47#_M1005_s 0.00223577f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_189 N_VGND_c_327_n N_A_229_47#_c_366_n 0.0197886f $X=2.56 $Y=0 $X2=0 $Y2=0
cc_190 N_VGND_c_329_n N_A_229_47#_c_366_n 0.012627f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_191 N_VGND_c_327_n N_A_229_47#_c_371_n 0.052801f $X=2.56 $Y=0 $X2=0 $Y2=0
cc_192 N_VGND_c_329_n N_A_229_47#_c_371_n 0.0338748f $X=3.12 $Y=0 $X2=0 $Y2=0
