* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__bufbuf_8 A VGND VNB VPB VPWR X
X0 VPWR A a_1217_23# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VGND a_117_265# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 X a_117_265# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 X a_117_265# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 X a_117_265# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND a_117_265# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_837_23# a_1217_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VPWR a_117_265# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND a_117_265# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR a_117_265# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 X a_117_265# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 X a_117_265# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_837_23# a_1217_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VPWR a_837_23# a_117_265# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VPWR a_837_23# a_117_265# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR a_117_265# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VPWR a_117_265# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 X a_117_265# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VGND A a_1217_23# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_837_23# a_117_265# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VGND a_837_23# a_117_265# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_117_265# a_837_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_117_265# a_837_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 X a_117_265# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VGND a_117_265# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 X a_117_265# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
