* File: sky130_fd_sc_lp__or4_lp.pxi.spice
* Created: Wed Sep  2 10:32:11 2020
* 
x_PM_SKY130_FD_SC_LP__OR4_LP%D N_D_c_88_n N_D_M1004_g N_D_c_89_n N_D_M1001_g
+ N_D_c_91_n N_D_c_92_n N_D_M1014_g N_D_c_93_n N_D_c_94_n D N_D_c_95_n
+ N_D_c_96_n N_D_c_97_n PM_SKY130_FD_SC_LP__OR4_LP%D
x_PM_SKY130_FD_SC_LP__OR4_LP%C N_C_M1009_g N_C_c_140_n N_C_M1005_g N_C_c_141_n
+ N_C_c_142_n N_C_M1006_g N_C_c_143_n N_C_c_144_n N_C_c_145_n N_C_c_146_n C C C
+ C N_C_c_147_n N_C_c_148_n PM_SKY130_FD_SC_LP__OR4_LP%C
x_PM_SKY130_FD_SC_LP__OR4_LP%B N_B_M1007_g N_B_c_208_n N_B_M1011_g N_B_c_210_n
+ N_B_M1010_g N_B_c_212_n B B B N_B_c_213_n N_B_c_214_n
+ PM_SKY130_FD_SC_LP__OR4_LP%B
x_PM_SKY130_FD_SC_LP__OR4_LP%A N_A_M1012_g N_A_M1003_g N_A_M1000_g A A A
+ N_A_c_259_n N_A_c_260_n PM_SKY130_FD_SC_LP__OR4_LP%A
x_PM_SKY130_FD_SC_LP__OR4_LP%A_27_47# N_A_27_47#_M1004_s N_A_27_47#_M1006_d
+ N_A_27_47#_M1010_d N_A_27_47#_M1001_s N_A_27_47#_M1008_g N_A_27_47#_c_302_n
+ N_A_27_47#_M1002_g N_A_27_47#_c_303_n N_A_27_47#_M1013_g N_A_27_47#_c_304_n
+ N_A_27_47#_c_305_n N_A_27_47#_c_306_n N_A_27_47#_c_307_n N_A_27_47#_c_308_n
+ N_A_27_47#_c_309_n N_A_27_47#_c_310_n N_A_27_47#_c_311_n N_A_27_47#_c_312_n
+ N_A_27_47#_c_313_n N_A_27_47#_c_321_n N_A_27_47#_c_314_n N_A_27_47#_c_315_n
+ N_A_27_47#_c_316_n N_A_27_47#_c_317_n N_A_27_47#_c_318_n N_A_27_47#_c_319_n
+ PM_SKY130_FD_SC_LP__OR4_LP%A_27_47#
x_PM_SKY130_FD_SC_LP__OR4_LP%VPWR N_VPWR_M1012_d N_VPWR_c_442_n VPWR
+ N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_441_n N_VPWR_c_446_n
+ PM_SKY130_FD_SC_LP__OR4_LP%VPWR
x_PM_SKY130_FD_SC_LP__OR4_LP%X N_X_M1013_d N_X_M1008_d X X X X X X X X
+ PM_SKY130_FD_SC_LP__OR4_LP%X
x_PM_SKY130_FD_SC_LP__OR4_LP%VGND N_VGND_M1014_d N_VGND_M1011_s N_VGND_M1000_d
+ N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n N_VGND_c_502_n N_VGND_c_503_n
+ N_VGND_c_504_n VGND N_VGND_c_505_n N_VGND_c_506_n N_VGND_c_507_n
+ N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n PM_SKY130_FD_SC_LP__OR4_LP%VGND
cc_1 VNB N_D_c_88_n 0.0168862f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.73
cc_2 VNB N_D_c_89_n 0.0211205f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.7
cc_3 VNB N_D_M1001_g 0.00124935f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.595
cc_4 VNB N_D_c_91_n 0.0168434f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_5 VNB N_D_c_92_n 0.0135809f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_6 VNB N_D_c_93_n 0.00621403f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_7 VNB N_D_c_94_n 0.00453673f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.875
cc_8 VNB N_D_c_95_n 0.016166f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.37
cc_9 VNB N_D_c_96_n 0.00870305f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.37
cc_10 VNB N_D_c_97_n 0.0174604f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.205
cc_11 VNB N_C_c_140_n 0.0135729f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.7
cc_12 VNB N_C_c_141_n 0.0213147f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.595
cc_13 VNB N_C_c_142_n 0.0169272f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_14 VNB N_C_c_143_n 0.0276624f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_15 VNB N_C_c_144_n 0.0279605f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_16 VNB N_C_c_145_n 0.0102538f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.875
cc_17 VNB N_C_c_146_n 0.00647836f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB N_C_c_147_n 0.017834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_C_c_148_n 0.00190845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_c_208_n 0.0174119f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.205
cc_21 VNB N_B_M1011_g 0.0310043f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.595
cc_22 VNB N_B_c_210_n 0.0308227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_M1010_g 0.0294483f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_24 VNB N_B_c_212_n 0.00803211f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_25 VNB N_B_c_213_n 0.0277183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_c_214_n 0.00353287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_M1003_g 0.0268006f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.7
cc_28 VNB N_A_M1000_g 0.026127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_c_259_n 0.00648756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_c_260_n 0.00250966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_302_n 0.0158118f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.805
cc_32 VNB N_A_27_47#_c_303_n 0.019213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_c_304_n 0.00879304f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.205
cc_34 VNB N_A_27_47#_c_305_n 0.024222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_47#_c_306_n 6.54552e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_47#_c_307_n 0.0074432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_47#_c_308_n 0.0151673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_309_n 0.00481328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_47#_c_310_n 0.00559019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_47#_c_311_n 0.0172845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_47#_c_312_n 0.0175689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_47#_c_313_n 0.00786683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_47#_c_314_n 0.0298366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_47#_c_315_n 0.00938688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_47#_c_316_n 0.00112931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_47#_c_317_n 0.00253742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_47#_c_318_n 0.00636813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_47#_c_319_n 0.0309092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VPWR_c_441_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB X 0.0568716f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.7
cc_51 VNB N_VGND_c_499_n 0.00277613f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.805
cc_52 VNB N_VGND_c_500_n 0.00720572f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_53 VNB N_VGND_c_501_n 0.0291649f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_54 VNB N_VGND_c_502_n 0.0375687f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.37
cc_55 VNB N_VGND_c_503_n 0.0269126f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.37
cc_56 VNB N_VGND_c_504_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_505_n 0.0266387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_506_n 0.0352588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_507_n 0.028795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_508_n 0.298575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_509_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_510_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VPB N_D_c_89_n 0.00206778f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.7
cc_64 VPB N_D_M1001_g 0.0318737f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.595
cc_65 VPB N_D_c_94_n 0.011038f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.875
cc_66 VPB N_D_c_96_n 7.83792e-19 $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.37
cc_67 VPB N_C_M1009_g 0.0248978f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_68 VPB N_C_c_145_n 0.00367169f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.875
cc_69 VPB N_C_c_148_n 0.00110089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_B_M1007_g 0.0294186f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_71 VPB N_B_c_213_n 0.00379131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_B_c_214_n 0.00433323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_M1012_g 0.0314082f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_74 VPB N_A_c_259_n 0.0386787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_c_260_n 0.00705216f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_M1008_g 0.0496893f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_77 VPB N_A_27_47#_c_321_n 0.0520253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_314_n 0.0203848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_318_n 0.00100377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_319_n 0.0125695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_442_n 0.00766473f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.38
cc_82 VPB N_VPWR_c_443_n 0.0986188f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.805
cc_83 VPB N_VPWR_c_444_n 0.0255218f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_84 VPB N_VPWR_c_441_n 0.0500147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_446_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.37
cc_86 VPB X 0.0232352f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.7
cc_87 VPB X 0.054324f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=0.805
cc_88 N_D_M1001_g N_C_M1009_g 0.0264609f $X=0.645 $Y=2.595 $X2=0 $Y2=0
cc_89 N_D_c_92_n N_C_c_140_n 0.010654f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_90 N_D_c_95_n N_C_c_143_n 0.00143487f $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_91 N_D_c_96_n N_C_c_143_n 0.00122713f $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_92 N_D_c_97_n N_C_c_143_n 0.00290622f $X=0.595 $Y=1.205 $X2=0 $Y2=0
cc_93 N_D_c_89_n N_C_c_144_n 0.0264609f $X=0.595 $Y=1.7 $X2=0 $Y2=0
cc_94 N_D_c_94_n N_C_c_145_n 0.0264609f $X=0.595 $Y=1.875 $X2=0 $Y2=0
cc_95 N_D_c_91_n N_C_c_146_n 0.00896817f $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_96 N_D_c_95_n N_C_c_147_n 0.0264609f $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_97 N_D_c_96_n N_C_c_147_n 0.0037481f $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_98 N_D_M1001_g N_C_c_148_n 0.00461062f $X=0.645 $Y=2.595 $X2=0 $Y2=0
cc_99 N_D_c_95_n N_C_c_148_n 6.8793e-19 $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_100 N_D_c_96_n N_C_c_148_n 0.0467984f $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_101 N_D_c_88_n N_A_27_47#_c_304_n 0.00686503f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_102 N_D_c_91_n N_A_27_47#_c_305_n 0.0138352f $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_103 N_D_c_93_n N_A_27_47#_c_305_n 0.00419478f $X=0.495 $Y=0.805 $X2=0 $Y2=0
cc_104 N_D_c_95_n N_A_27_47#_c_305_n 6.57544e-19 $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_105 N_D_c_96_n N_A_27_47#_c_305_n 0.029436f $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_106 N_D_c_97_n N_A_27_47#_c_305_n 0.00876313f $X=0.595 $Y=1.205 $X2=0 $Y2=0
cc_107 N_D_c_91_n N_A_27_47#_c_306_n 4.90656e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_108 N_D_c_88_n N_A_27_47#_c_312_n 0.00763597f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_109 N_D_c_92_n N_A_27_47#_c_312_n 0.00111532f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_110 N_D_M1001_g N_A_27_47#_c_321_n 0.0255898f $X=0.645 $Y=2.595 $X2=0 $Y2=0
cc_111 N_D_c_94_n N_A_27_47#_c_321_n 0.00158954f $X=0.595 $Y=1.875 $X2=0 $Y2=0
cc_112 N_D_c_96_n N_A_27_47#_c_321_n 0.00799993f $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_113 N_D_M1001_g N_A_27_47#_c_314_n 0.00656371f $X=0.645 $Y=2.595 $X2=0 $Y2=0
cc_114 N_D_c_96_n N_A_27_47#_c_314_n 0.0487791f $X=0.605 $Y=1.37 $X2=0 $Y2=0
cc_115 N_D_c_97_n N_A_27_47#_c_314_n 0.0222725f $X=0.595 $Y=1.205 $X2=0 $Y2=0
cc_116 N_D_M1001_g N_VPWR_c_443_n 0.00939541f $X=0.645 $Y=2.595 $X2=0 $Y2=0
cc_117 N_D_M1001_g N_VPWR_c_441_n 0.0171501f $X=0.645 $Y=2.595 $X2=0 $Y2=0
cc_118 N_D_c_88_n N_VGND_c_499_n 0.00239794f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_119 N_D_c_92_n N_VGND_c_499_n 0.0127761f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_120 N_D_c_88_n N_VGND_c_505_n 0.00549284f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_121 N_D_c_91_n N_VGND_c_505_n 4.87571e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_122 N_D_c_92_n N_VGND_c_505_n 0.00486043f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_123 N_D_c_88_n N_VGND_c_508_n 0.00720061f $X=0.495 $Y=0.73 $X2=0 $Y2=0
cc_124 N_D_c_91_n N_VGND_c_508_n 6.51792e-19 $X=0.78 $Y=0.805 $X2=0 $Y2=0
cc_125 N_D_c_92_n N_VGND_c_508_n 0.00443987f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_126 N_C_M1009_g N_B_M1007_g 0.051978f $X=1.135 $Y=2.595 $X2=0 $Y2=0
cc_127 N_C_c_148_n N_B_M1007_g 0.00354792f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_128 N_C_c_141_n N_B_M1011_g 0.00207594f $X=1.57 $Y=0.805 $X2=0 $Y2=0
cc_129 N_C_c_144_n N_B_c_213_n 0.0181726f $X=1.175 $Y=1.77 $X2=0 $Y2=0
cc_130 N_C_c_148_n N_B_c_213_n 8.52047e-19 $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_131 N_C_M1009_g N_B_c_214_n 0.00112585f $X=1.135 $Y=2.595 $X2=0 $Y2=0
cc_132 N_C_c_144_n N_B_c_214_n 0.00172928f $X=1.175 $Y=1.77 $X2=0 $Y2=0
cc_133 N_C_c_148_n N_B_c_214_n 0.0552513f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_134 N_C_c_141_n N_A_27_47#_c_305_n 0.0068275f $X=1.57 $Y=0.805 $X2=0 $Y2=0
cc_135 N_C_c_143_n N_A_27_47#_c_305_n 0.0106496f $X=1.175 $Y=1.265 $X2=0 $Y2=0
cc_136 N_C_c_146_n N_A_27_47#_c_305_n 0.00457635f $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_137 N_C_c_147_n N_A_27_47#_c_305_n 0.00115978f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_138 N_C_c_148_n N_A_27_47#_c_305_n 0.0196313f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_139 N_C_c_140_n N_A_27_47#_c_306_n 0.00110574f $X=1.285 $Y=0.73 $X2=0 $Y2=0
cc_140 N_C_c_141_n N_A_27_47#_c_306_n 0.00614559f $X=1.57 $Y=0.805 $X2=0 $Y2=0
cc_141 N_C_c_142_n N_A_27_47#_c_306_n 0.00236045f $X=1.645 $Y=0.73 $X2=0 $Y2=0
cc_142 N_C_c_143_n N_A_27_47#_c_307_n 0.00942903f $X=1.175 $Y=1.265 $X2=0 $Y2=0
cc_143 N_C_c_148_n N_A_27_47#_c_307_n 0.00428316f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_144 N_C_c_141_n N_A_27_47#_c_308_n 6.67655e-19 $X=1.57 $Y=0.805 $X2=0 $Y2=0
cc_145 N_C_c_147_n N_A_27_47#_c_309_n 0.00392071f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_146 N_C_c_148_n N_A_27_47#_c_309_n 0.0136967f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_147 N_C_M1009_g N_A_27_47#_c_321_n 0.00278509f $X=1.135 $Y=2.595 $X2=0 $Y2=0
cc_148 N_C_c_148_n N_A_27_47#_c_321_n 0.0276764f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_149 N_C_c_140_n N_A_27_47#_c_315_n 0.00115811f $X=1.285 $Y=0.73 $X2=0 $Y2=0
cc_150 N_C_c_142_n N_A_27_47#_c_315_n 0.017989f $X=1.645 $Y=0.73 $X2=0 $Y2=0
cc_151 N_C_c_141_n N_A_27_47#_c_316_n 0.00470634f $X=1.57 $Y=0.805 $X2=0 $Y2=0
cc_152 N_C_c_148_n A_252_419# 0.00809094f $X=1.175 $Y=1.43 $X2=-0.19 $Y2=-0.245
cc_153 N_C_M1009_g N_VPWR_c_443_n 0.00656883f $X=1.135 $Y=2.595 $X2=0 $Y2=0
cc_154 N_C_c_148_n N_VPWR_c_443_n 0.00914393f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_155 N_C_M1009_g N_VPWR_c_441_n 0.00824494f $X=1.135 $Y=2.595 $X2=0 $Y2=0
cc_156 N_C_c_148_n N_VPWR_c_441_n 0.0101955f $X=1.175 $Y=1.43 $X2=0 $Y2=0
cc_157 N_C_c_140_n N_VGND_c_499_n 0.0113789f $X=1.285 $Y=0.73 $X2=0 $Y2=0
cc_158 N_C_c_142_n N_VGND_c_499_n 0.00168537f $X=1.645 $Y=0.73 $X2=0 $Y2=0
cc_159 N_C_c_146_n N_VGND_c_499_n 6.29884e-19 $X=1.275 $Y=0.805 $X2=0 $Y2=0
cc_160 N_C_c_143_n N_VGND_c_500_n 6.86331e-19 $X=1.175 $Y=1.265 $X2=0 $Y2=0
cc_161 N_C_c_141_n N_VGND_c_501_n 3.39508e-19 $X=1.57 $Y=0.805 $X2=0 $Y2=0
cc_162 N_C_c_142_n N_VGND_c_501_n 0.00566916f $X=1.645 $Y=0.73 $X2=0 $Y2=0
cc_163 N_C_c_140_n N_VGND_c_503_n 0.00486043f $X=1.285 $Y=0.73 $X2=0 $Y2=0
cc_164 N_C_c_141_n N_VGND_c_503_n 4.87571e-19 $X=1.57 $Y=0.805 $X2=0 $Y2=0
cc_165 N_C_c_142_n N_VGND_c_503_n 0.00359964f $X=1.645 $Y=0.73 $X2=0 $Y2=0
cc_166 N_C_c_140_n N_VGND_c_508_n 0.00443987f $X=1.285 $Y=0.73 $X2=0 $Y2=0
cc_167 N_C_c_141_n N_VGND_c_508_n 6.51792e-19 $X=1.57 $Y=0.805 $X2=0 $Y2=0
cc_168 N_C_c_142_n N_VGND_c_508_n 0.00661248f $X=1.645 $Y=0.73 $X2=0 $Y2=0
cc_169 N_B_M1010_g N_A_M1003_g 0.0238235f $X=2.725 $Y=1.045 $X2=0 $Y2=0
cc_170 N_B_c_210_n N_A_c_259_n 0.00950942f $X=2.65 $Y=1.68 $X2=0 $Y2=0
cc_171 N_B_M1007_g N_A_c_260_n 0.00325001f $X=1.705 $Y=2.595 $X2=0 $Y2=0
cc_172 N_B_c_210_n N_A_c_260_n 0.0149604f $X=2.65 $Y=1.68 $X2=0 $Y2=0
cc_173 N_B_c_213_n N_A_c_260_n 6.92659e-19 $X=1.745 $Y=1.68 $X2=0 $Y2=0
cc_174 N_B_c_214_n N_A_c_260_n 0.0827977f $X=1.745 $Y=1.77 $X2=0 $Y2=0
cc_175 N_B_M1011_g N_A_27_47#_c_306_n 2.16691e-19 $X=2.25 $Y=1.135 $X2=0 $Y2=0
cc_176 N_B_M1011_g N_A_27_47#_c_307_n 0.00309178f $X=2.25 $Y=1.135 $X2=0 $Y2=0
cc_177 N_B_M1011_g N_A_27_47#_c_308_n 0.0141147f $X=2.25 $Y=1.135 $X2=0 $Y2=0
cc_178 N_B_c_210_n N_A_27_47#_c_308_n 0.00475759f $X=2.65 $Y=1.68 $X2=0 $Y2=0
cc_179 N_B_M1010_g N_A_27_47#_c_308_n 0.0112536f $X=2.725 $Y=1.045 $X2=0 $Y2=0
cc_180 N_B_c_213_n N_A_27_47#_c_308_n 0.0113383f $X=1.745 $Y=1.68 $X2=0 $Y2=0
cc_181 N_B_c_214_n N_A_27_47#_c_308_n 0.044191f $X=1.745 $Y=1.77 $X2=0 $Y2=0
cc_182 N_B_c_213_n N_A_27_47#_c_309_n 0.00323735f $X=1.745 $Y=1.68 $X2=0 $Y2=0
cc_183 N_B_c_214_n N_A_27_47#_c_309_n 0.0106482f $X=1.745 $Y=1.77 $X2=0 $Y2=0
cc_184 N_B_M1011_g N_A_27_47#_c_310_n 0.00116053f $X=2.25 $Y=1.135 $X2=0 $Y2=0
cc_185 N_B_M1010_g N_A_27_47#_c_310_n 0.00981896f $X=2.725 $Y=1.045 $X2=0 $Y2=0
cc_186 N_B_M1011_g N_A_27_47#_c_316_n 6.79925e-19 $X=2.25 $Y=1.135 $X2=0 $Y2=0
cc_187 N_B_M1010_g N_A_27_47#_c_317_n 0.0027409f $X=2.725 $Y=1.045 $X2=0 $Y2=0
cc_188 N_B_c_214_n A_366_419# 0.0274295f $X=1.745 $Y=1.77 $X2=-0.19 $Y2=-0.245
cc_189 N_B_M1007_g N_VPWR_c_443_n 0.00655603f $X=1.705 $Y=2.595 $X2=0 $Y2=0
cc_190 N_B_c_214_n N_VPWR_c_443_n 0.0209526f $X=1.745 $Y=1.77 $X2=0 $Y2=0
cc_191 N_B_M1007_g N_VPWR_c_441_n 0.00975774f $X=1.705 $Y=2.595 $X2=0 $Y2=0
cc_192 N_B_c_214_n N_VPWR_c_441_n 0.0234398f $X=1.745 $Y=1.77 $X2=0 $Y2=0
cc_193 N_B_M1011_g N_VGND_c_500_n 0.0124523f $X=2.25 $Y=1.135 $X2=0 $Y2=0
cc_194 N_B_M1010_g N_VGND_c_500_n 0.00213765f $X=2.725 $Y=1.045 $X2=0 $Y2=0
cc_195 N_B_M1011_g N_VGND_c_501_n 0.00380794f $X=2.25 $Y=1.135 $X2=0 $Y2=0
cc_196 N_B_M1010_g N_VGND_c_501_n 0.00399215f $X=2.725 $Y=1.045 $X2=0 $Y2=0
cc_197 N_B_M1010_g N_VGND_c_506_n 0.00320058f $X=2.725 $Y=1.045 $X2=0 $Y2=0
cc_198 N_B_M1011_g N_VGND_c_508_n 0.00291506f $X=2.25 $Y=1.135 $X2=0 $Y2=0
cc_199 N_B_M1010_g N_VGND_c_508_n 0.00415093f $X=2.725 $Y=1.045 $X2=0 $Y2=0
cc_200 N_A_M1012_g N_A_27_47#_M1008_g 0.01253f $X=3.165 $Y=2.595 $X2=0 $Y2=0
cc_201 N_A_c_259_n N_A_27_47#_M1008_g 0.00840646f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_202 N_A_c_260_n N_A_27_47#_M1008_g 0.00575118f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_203 N_A_M1000_g N_A_27_47#_c_302_n 0.0152538f $X=3.515 $Y=1.045 $X2=0 $Y2=0
cc_204 N_A_c_260_n N_A_27_47#_c_308_n 0.0185092f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_205 N_A_M1003_g N_A_27_47#_c_310_n 0.0103174f $X=3.155 $Y=1.045 $X2=0 $Y2=0
cc_206 N_A_M1000_g N_A_27_47#_c_310_n 0.00179788f $X=3.515 $Y=1.045 $X2=0 $Y2=0
cc_207 N_A_M1003_g N_A_27_47#_c_311_n 0.0104907f $X=3.155 $Y=1.045 $X2=0 $Y2=0
cc_208 N_A_M1000_g N_A_27_47#_c_311_n 0.0165958f $X=3.515 $Y=1.045 $X2=0 $Y2=0
cc_209 N_A_c_259_n N_A_27_47#_c_311_n 7.25569e-19 $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_210 N_A_c_260_n N_A_27_47#_c_311_n 0.0196975f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_211 N_A_M1003_g N_A_27_47#_c_317_n 0.0027409f $X=3.155 $Y=1.045 $X2=0 $Y2=0
cc_212 N_A_c_259_n N_A_27_47#_c_317_n 0.00117535f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_213 N_A_c_260_n N_A_27_47#_c_317_n 0.0290435f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_214 N_A_M1000_g N_A_27_47#_c_318_n 0.00142322f $X=3.515 $Y=1.045 $X2=0 $Y2=0
cc_215 N_A_c_260_n N_A_27_47#_c_318_n 6.89066e-19 $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_216 N_A_M1000_g N_A_27_47#_c_319_n 0.0178875f $X=3.515 $Y=1.045 $X2=0 $Y2=0
cc_217 N_A_c_260_n A_366_419# 0.0307802f $X=3.205 $Y=1.77 $X2=-0.19 $Y2=-0.245
cc_218 N_A_c_260_n N_VPWR_M1012_d 0.00830291f $X=3.205 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_219 N_A_M1012_g N_VPWR_c_442_n 0.0099193f $X=3.165 $Y=2.595 $X2=0 $Y2=0
cc_220 N_A_c_259_n N_VPWR_c_442_n 0.00106846f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_221 N_A_c_260_n N_VPWR_c_442_n 0.0662953f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_222 N_A_M1012_g N_VPWR_c_443_n 0.00655603f $X=3.165 $Y=2.595 $X2=0 $Y2=0
cc_223 N_A_c_260_n N_VPWR_c_443_n 0.0245902f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_224 N_A_M1012_g N_VPWR_c_441_n 0.0102422f $X=3.165 $Y=2.595 $X2=0 $Y2=0
cc_225 N_A_c_260_n N_VPWR_c_441_n 0.0281468f $X=3.205 $Y=1.77 $X2=0 $Y2=0
cc_226 N_A_M1003_g N_VGND_c_502_n 0.00144992f $X=3.155 $Y=1.045 $X2=0 $Y2=0
cc_227 N_A_M1000_g N_VGND_c_502_n 0.0096192f $X=3.515 $Y=1.045 $X2=0 $Y2=0
cc_228 N_A_M1003_g N_VGND_c_506_n 0.00320058f $X=3.155 $Y=1.045 $X2=0 $Y2=0
cc_229 N_A_M1000_g N_VGND_c_506_n 0.00266097f $X=3.515 $Y=1.045 $X2=0 $Y2=0
cc_230 N_A_M1003_g N_VGND_c_508_n 0.00415093f $X=3.155 $Y=1.045 $X2=0 $Y2=0
cc_231 N_A_M1000_g N_VGND_c_508_n 0.00348678f $X=3.515 $Y=1.045 $X2=0 $Y2=0
cc_232 N_A_27_47#_M1008_g N_VPWR_c_442_n 0.0246713f $X=3.98 $Y=2.595 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_311_n N_VPWR_c_442_n 0.010409f $X=3.845 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_318_n N_VPWR_c_442_n 0.00143312f $X=4.01 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_321_n N_VPWR_c_443_n 0.0281861f $X=0.38 $Y=2.24 $X2=0 $Y2=0
cc_236 N_A_27_47#_M1008_g N_VPWR_c_444_n 0.00838695f $X=3.98 $Y=2.595 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_M1001_s N_VPWR_c_441_n 0.0023218f $X=0.235 $Y=2.095 $X2=0
+ $Y2=0
cc_238 N_A_27_47#_M1008_g N_VPWR_c_441_n 0.0146536f $X=3.98 $Y=2.595 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_321_n N_VPWR_c_441_n 0.0173447f $X=0.38 $Y=2.24 $X2=0 $Y2=0
cc_240 N_A_27_47#_M1008_g X 0.013629f $X=3.98 $Y=2.595 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_302_n X 0.00213114f $X=3.945 $Y=1.365 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_303_n X 0.0164317f $X=4.305 $Y=1.365 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_318_n X 0.0266514f $X=4.01 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_319_n X 0.0127997f $X=4.305 $Y=1.53 $X2=0 $Y2=0
cc_245 N_A_27_47#_M1008_g X 0.025213f $X=3.98 $Y=2.595 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_318_n X 0.00428474f $X=4.01 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_319_n X 0.00749752f $X=4.305 $Y=1.53 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_308_n N_VGND_M1011_s 0.00259881f $X=2.775 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_305_n N_VGND_c_499_n 0.0254874f $X=1.52 $Y=0.94 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_312_n N_VGND_c_499_n 0.0137946f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_315_n N_VGND_c_499_n 0.0107298f $X=1.94 $Y=0.47 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_307_n N_VGND_c_500_n 0.00949579f $X=1.605 $Y=1.325 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_308_n N_VGND_c_500_n 0.0336211f $X=2.775 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_310_n N_VGND_c_500_n 0.0125448f $X=2.94 $Y=1.045 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_315_n N_VGND_c_500_n 0.0162752f $X=1.94 $Y=0.47 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_316_n N_VGND_c_500_n 0.0114739f $X=1.605 $Y=0.94 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_306_n N_VGND_c_501_n 0.00475325f $X=1.605 $Y=0.855 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_310_n N_VGND_c_501_n 0.00363959f $X=2.94 $Y=1.045 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_315_n N_VGND_c_501_n 0.0326819f $X=1.94 $Y=0.47 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_316_n N_VGND_c_501_n 0.00113417f $X=1.605 $Y=0.94 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_302_n N_VGND_c_502_n 0.00946746f $X=3.945 $Y=1.365 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_303_n N_VGND_c_502_n 0.0011976f $X=4.305 $Y=1.365 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_310_n N_VGND_c_502_n 0.0110409f $X=2.94 $Y=1.045 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_311_n N_VGND_c_502_n 0.0181022f $X=3.845 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_318_n N_VGND_c_502_n 0.00279839f $X=4.01 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_315_n N_VGND_c_503_n 0.0335499f $X=1.94 $Y=0.47 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_312_n N_VGND_c_505_n 0.0211775f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_302_n N_VGND_c_507_n 0.00266097f $X=3.945 $Y=1.365 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_303_n N_VGND_c_507_n 0.00275863f $X=4.305 $Y=1.365 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_M1004_s N_VGND_c_508_n 0.00232985f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1006_d N_VGND_c_508_n 0.0030013f $X=1.72 $Y=0.235 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_302_n N_VGND_c_508_n 0.00348678f $X=3.945 $Y=1.365 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_303_n N_VGND_c_508_n 0.00348678f $X=4.305 $Y=1.365 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_305_n N_VGND_c_508_n 0.0228112f $X=1.52 $Y=0.94 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_310_n N_VGND_c_508_n 0.0130316f $X=2.94 $Y=1.045 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_312_n N_VGND_c_508_n 0.0134543f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_315_n N_VGND_c_508_n 0.0216319f $X=1.94 $Y=0.47 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_308_n A_465_185# 0.00536262f $X=2.775 $Y=1.41 $X2=-0.19
+ $Y2=-0.245
cc_279 A_154_419# N_VPWR_c_441_n 0.010279f $X=0.77 $Y=2.095 $X2=4.56 $Y2=3.33
cc_280 A_252_419# N_VPWR_c_441_n 0.010571f $X=1.26 $Y=2.095 $X2=1.115 $Y2=1.58
cc_281 A_366_419# N_VPWR_c_441_n 0.0198216f $X=1.83 $Y=2.095 $X2=1.595 $Y2=2.69
cc_282 N_VPWR_c_441_n N_X_M1008_d 0.0023218f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_283 N_VPWR_c_442_n X 0.068131f $X=3.715 $Y=2.24 $X2=0 $Y2=0
cc_284 N_VPWR_c_444_n X 0.028866f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_285 N_VPWR_c_441_n X 0.022162f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_286 X N_VGND_c_502_n 0.0258123f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_287 X N_VGND_c_507_n 0.0107254f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_288 X N_VGND_c_508_n 0.0114362f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_289 A_114_47# N_VGND_c_508_n 0.00312872f $X=0.57 $Y=0.235 $X2=4.56 $Y2=0
cc_290 N_VGND_c_508_n A_272_47# 0.00277835f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
cc_291 N_VGND_c_500_n A_465_185# 0.00358252f $X=2.285 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_292 N_VGND_c_501_n A_465_185# 6.45569e-19 $X=2.37 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
