* File: sky130_fd_sc_lp__o311ai_4.pex.spice
* Created: Wed Sep  2 10:23:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311AI_4%A1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 52
r78 50 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.69 $Y=1.35 $X2=1.78
+ $Y2=1.35
r79 47 50 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.35 $Y=1.35
+ $X2=1.69 $Y2=1.35
r80 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=1.35 $X2=1.35 $Y2=1.35
r81 45 47 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.92 $Y=1.35
+ $X2=1.35 $Y2=1.35
r82 43 45 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.67 $Y=1.35
+ $X2=0.92 $Y2=1.35
r83 41 43 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.49 $Y=1.35 $X2=0.67
+ $Y2=1.35
r84 38 41 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.33 $Y=1.35
+ $X2=0.49 $Y2=1.35
r85 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.33
+ $Y=1.35 $X2=0.33 $Y2=1.35
r86 32 48 14.914 $w=2.53e-07 $l=3.3e-07 $layer=LI1_cond $X=1.68 $Y=1.307
+ $X2=1.35 $Y2=1.307
r87 32 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.35 $X2=1.69 $Y2=1.35
r88 31 48 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=1.2 $Y=1.307
+ $X2=1.35 $Y2=1.307
r89 30 31 23.9527 $w=2.53e-07 $l=5.3e-07 $layer=LI1_cond $X=0.67 $Y=1.307
+ $X2=1.2 $Y2=1.307
r90 30 39 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.67 $Y=1.307
+ $X2=0.33 $Y2=1.307
r91 30 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.35 $X2=0.67 $Y2=1.35
r92 29 39 4.06745 $w=2.53e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=1.307 $X2=0.33
+ $Y2=1.307
r93 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.515
+ $X2=1.78 $Y2=1.35
r94 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.78 $Y=1.515
+ $X2=1.78 $Y2=2.465
r95 22 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.185
+ $X2=1.78 $Y2=1.35
r96 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.78 $Y=1.185
+ $X2=1.78 $Y2=0.655
r97 18 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.515
+ $X2=1.35 $Y2=1.35
r98 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.35 $Y=1.515
+ $X2=1.35 $Y2=2.465
r99 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.185
+ $X2=1.35 $Y2=1.35
r100 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.35 $Y=1.185
+ $X2=1.35 $Y2=0.655
r101 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.515
+ $X2=0.92 $Y2=1.35
r102 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.92 $Y=1.515
+ $X2=0.92 $Y2=2.465
r103 8 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.185
+ $X2=0.92 $Y2=1.35
r104 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.92 $Y=1.185
+ $X2=0.92 $Y2=0.655
r105 4 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.515
+ $X2=0.49 $Y2=1.35
r106 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.49 $Y=1.515
+ $X2=0.49 $Y2=2.465
r107 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.185
+ $X2=0.49 $Y2=1.35
r108 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.49 $Y=1.185
+ $X2=0.49 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 49
r94 47 49 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.32 $Y=1.35 $X2=3.5
+ $Y2=1.35
r95 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.32
+ $Y=1.35 $X2=3.32 $Y2=1.35
r96 45 47 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.07 $Y=1.35
+ $X2=3.32 $Y2=1.35
r97 43 45 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.98 $Y=1.35 $X2=3.07
+ $Y2=1.35
r98 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.98
+ $Y=1.35 $X2=2.98 $Y2=1.35
r99 40 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.64 $Y=1.35
+ $X2=2.98 $Y2=1.35
r100 37 40 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.21 $Y=1.35
+ $X2=2.64 $Y2=1.35
r101 32 48 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=3.6 $Y=1.307
+ $X2=3.32 $Y2=1.307
r102 31 48 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=3.12 $Y=1.307
+ $X2=3.32 $Y2=1.307
r103 31 44 6.32714 $w=2.53e-07 $l=1.4e-07 $layer=LI1_cond $X=3.12 $Y=1.307
+ $X2=2.98 $Y2=1.307
r104 30 44 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=2.64 $Y=1.307
+ $X2=2.98 $Y2=1.307
r105 30 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.64
+ $Y=1.35 $X2=2.64 $Y2=1.35
r106 29 30 21.693 $w=2.53e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.307
+ $X2=2.64 $Y2=1.307
r107 25 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.5 $Y=1.515
+ $X2=3.5 $Y2=1.35
r108 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.5 $Y=1.515
+ $X2=3.5 $Y2=2.465
r109 22 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.5 $Y=1.185
+ $X2=3.5 $Y2=1.35
r110 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.5 $Y=1.185
+ $X2=3.5 $Y2=0.655
r111 18 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.515
+ $X2=3.07 $Y2=1.35
r112 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.07 $Y=1.515
+ $X2=3.07 $Y2=2.465
r113 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.185
+ $X2=3.07 $Y2=1.35
r114 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.07 $Y=1.185
+ $X2=3.07 $Y2=0.655
r115 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=1.515
+ $X2=2.64 $Y2=1.35
r116 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.64 $Y=1.515
+ $X2=2.64 $Y2=2.465
r117 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=1.185
+ $X2=2.64 $Y2=1.35
r118 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.64 $Y=1.185
+ $X2=2.64 $Y2=0.655
r119 4 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.515
+ $X2=2.21 $Y2=1.35
r120 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.21 $Y=1.515
+ $X2=2.21 $Y2=2.465
r121 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.185
+ $X2=2.21 $Y2=1.35
r122 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.21 $Y=1.185
+ $X2=2.21 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%A3 3 6 9 13 17 21 25 29 33 35 36 37 38 44
+ 58
c92 58 0 1.96662e-19 $X=5.75 $Y=1.51
r93 56 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.66 $Y=1.51 $X2=5.75
+ $Y2=1.51
r94 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.66
+ $Y=1.51 $X2=5.66 $Y2=1.51
r95 53 56 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.32 $Y=1.51
+ $X2=5.66 $Y2=1.51
r96 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.32
+ $Y=1.51 $X2=5.32 $Y2=1.51
r97 51 53 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=5.22 $Y=1.51 $X2=5.32
+ $Y2=1.51
r98 50 51 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=4.89 $Y=1.51
+ $X2=5.22 $Y2=1.51
r99 49 50 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.79 $Y=1.51 $X2=4.89
+ $Y2=1.51
r100 47 49 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.64 $Y=1.51
+ $X2=4.79 $Y2=1.51
r101 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.64
+ $Y=1.51 $X2=4.64 $Y2=1.51
r102 45 47 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.46 $Y=1.51
+ $X2=4.64 $Y2=1.51
r103 43 45 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.36 $Y=1.51 $X2=4.46
+ $Y2=1.51
r104 43 44 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.36 $Y=1.51
+ $X2=4.285 $Y2=1.51
r105 38 57 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=6 $Y=1.587 $X2=5.66
+ $Y2=1.587
r106 37 57 4.96437 $w=3.23e-07 $l=1.4e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.66 $Y2=1.587
r107 37 54 7.09196 $w=3.23e-07 $l=2e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.32 $Y2=1.587
r108 36 54 9.92874 $w=3.23e-07 $l=2.8e-07 $layer=LI1_cond $X=5.04 $Y=1.587
+ $X2=5.32 $Y2=1.587
r109 36 48 14.1839 $w=3.23e-07 $l=4e-07 $layer=LI1_cond $X=5.04 $Y=1.587
+ $X2=4.64 $Y2=1.587
r110 35 48 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.64 $Y2=1.587
r111 31 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.75 $Y=1.675
+ $X2=5.75 $Y2=1.51
r112 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.75 $Y=1.675
+ $X2=5.75 $Y2=2.465
r113 27 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=1.675
+ $X2=5.32 $Y2=1.51
r114 27 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.32 $Y=1.675
+ $X2=5.32 $Y2=2.465
r115 23 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.22 $Y=1.345
+ $X2=5.22 $Y2=1.51
r116 23 25 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.22 $Y=1.345
+ $X2=5.22 $Y2=0.655
r117 19 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.675
+ $X2=4.89 $Y2=1.51
r118 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.89 $Y=1.675
+ $X2=4.89 $Y2=2.465
r119 15 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=1.345
+ $X2=4.79 $Y2=1.51
r120 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.79 $Y=1.345
+ $X2=4.79 $Y2=0.655
r121 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.46 $Y=1.675
+ $X2=4.46 $Y2=1.51
r122 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.46 $Y=1.675
+ $X2=4.46 $Y2=2.465
r123 7 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.36 $Y=1.345
+ $X2=4.36 $Y2=1.51
r124 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.36 $Y=1.345
+ $X2=4.36 $Y2=0.655
r125 6 44 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.005 $Y=1.42
+ $X2=4.285 $Y2=1.42
r126 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.93 $Y=1.345
+ $X2=4.005 $Y2=1.42
r127 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.93 $Y=1.345
+ $X2=3.93 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 46 47
c72 47 0 1.29791e-19 $X=7.47 $Y=1.535
c73 46 0 1.96662e-19 $X=7.45 $Y=1.51
r74 47 48 8.9734 $w=3.76e-07 $l=7e-08 $layer=POLY_cond $X=7.47 $Y=1.535 $X2=7.54
+ $Y2=1.535
r75 45 47 2.56383 $w=3.76e-07 $l=2e-08 $layer=POLY_cond $X=7.45 $Y=1.535
+ $X2=7.47 $Y2=1.535
r76 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.45
+ $Y=1.51 $X2=7.45 $Y2=1.51
r77 43 45 51.2766 $w=3.76e-07 $l=4e-07 $layer=POLY_cond $X=7.05 $Y=1.535
+ $X2=7.45 $Y2=1.535
r78 42 43 1.28191 $w=3.76e-07 $l=1e-08 $layer=POLY_cond $X=7.04 $Y=1.535
+ $X2=7.05 $Y2=1.535
r79 41 42 53.8404 $w=3.76e-07 $l=4.2e-07 $layer=POLY_cond $X=6.62 $Y=1.535
+ $X2=7.04 $Y2=1.535
r80 40 41 1.28191 $w=3.76e-07 $l=1e-08 $layer=POLY_cond $X=6.61 $Y=1.535
+ $X2=6.62 $Y2=1.535
r81 38 40 23.0745 $w=3.76e-07 $l=1.8e-07 $layer=POLY_cond $X=6.43 $Y=1.535
+ $X2=6.61 $Y2=1.535
r82 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.43
+ $Y=1.51 $X2=6.43 $Y2=1.51
r83 36 38 30.766 $w=3.76e-07 $l=2.4e-07 $layer=POLY_cond $X=6.19 $Y=1.535
+ $X2=6.43 $Y2=1.535
r84 35 36 1.28191 $w=3.76e-07 $l=1e-08 $layer=POLY_cond $X=6.18 $Y=1.535
+ $X2=6.19 $Y2=1.535
r85 31 46 0.354598 $w=3.23e-07 $l=1e-08 $layer=LI1_cond $X=7.44 $Y=1.587
+ $X2=7.45 $Y2=1.587
r86 30 31 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.587
+ $X2=7.44 $Y2=1.587
r87 29 30 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.587
+ $X2=6.96 $Y2=1.587
r88 29 39 1.77299 $w=3.23e-07 $l=5e-08 $layer=LI1_cond $X=6.48 $Y=1.587 $X2=6.43
+ $Y2=1.587
r89 25 48 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.54 $Y=1.345
+ $X2=7.54 $Y2=1.535
r90 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.54 $Y=1.345 $X2=7.54
+ $Y2=0.745
r91 22 47 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.47 $Y=1.725
+ $X2=7.47 $Y2=1.535
r92 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.47 $Y=1.725
+ $X2=7.47 $Y2=2.465
r93 18 43 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.05 $Y=1.345
+ $X2=7.05 $Y2=1.535
r94 18 20 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.05 $Y=1.345 $X2=7.05
+ $Y2=0.745
r95 15 42 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.04 $Y=1.725
+ $X2=7.04 $Y2=1.535
r96 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.04 $Y=1.725
+ $X2=7.04 $Y2=2.465
r97 11 41 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.62 $Y=1.345
+ $X2=6.62 $Y2=1.535
r98 11 13 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.62 $Y=1.345 $X2=6.62
+ $Y2=0.745
r99 8 40 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.61 $Y=1.725 $X2=6.61
+ $Y2=1.535
r100 8 10 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.61 $Y=1.725
+ $X2=6.61 $Y2=2.465
r101 4 36 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.19 $Y=1.345
+ $X2=6.19 $Y2=1.535
r102 4 6 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.19 $Y=1.345 $X2=6.19
+ $Y2=0.745
r103 1 35 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.18 $Y=1.725
+ $X2=6.18 $Y2=1.535
r104 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.18 $Y=1.725
+ $X2=6.18 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%C1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 33 52
r79 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.69
+ $Y=1.51 $X2=9.69 $Y2=1.51
r80 52 54 27.7315 $w=3.65e-07 $l=2.1e-07 $layer=POLY_cond $X=9.48 $Y=1.535
+ $X2=9.69 $Y2=1.535
r81 51 52 38.2959 $w=3.65e-07 $l=2.9e-07 $layer=POLY_cond $X=9.19 $Y=1.535
+ $X2=9.48 $Y2=1.535
r82 49 51 23.7699 $w=3.65e-07 $l=1.8e-07 $layer=POLY_cond $X=9.01 $Y=1.535
+ $X2=9.19 $Y2=1.535
r83 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.01
+ $Y=1.51 $X2=9.01 $Y2=1.51
r84 47 49 3.96164 $w=3.65e-07 $l=3e-08 $layer=POLY_cond $X=8.98 $Y=1.535
+ $X2=9.01 $Y2=1.535
r85 46 47 29.0521 $w=3.65e-07 $l=2.2e-07 $layer=POLY_cond $X=8.76 $Y=1.535
+ $X2=8.98 $Y2=1.535
r86 45 46 30.3726 $w=3.65e-07 $l=2.3e-07 $layer=POLY_cond $X=8.53 $Y=1.535
+ $X2=8.76 $Y2=1.535
r87 44 45 26.411 $w=3.65e-07 $l=2e-07 $layer=POLY_cond $X=8.33 $Y=1.535 $X2=8.53
+ $Y2=1.535
r88 42 44 44.8986 $w=3.65e-07 $l=3.4e-07 $layer=POLY_cond $X=7.99 $Y=1.535
+ $X2=8.33 $Y2=1.535
r89 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.99
+ $Y=1.51 $X2=7.99 $Y2=1.51
r90 40 42 1.32055 $w=3.65e-07 $l=1e-08 $layer=POLY_cond $X=7.98 $Y=1.535
+ $X2=7.99 $Y2=1.535
r91 39 40 10.5644 $w=3.65e-07 $l=8e-08 $layer=POLY_cond $X=7.9 $Y=1.535 $X2=7.98
+ $Y2=1.535
r92 33 55 5.31897 $w=3.23e-07 $l=1.5e-07 $layer=LI1_cond $X=9.84 $Y=1.587
+ $X2=9.69 $Y2=1.587
r93 32 55 11.7017 $w=3.23e-07 $l=3.3e-07 $layer=LI1_cond $X=9.36 $Y=1.587
+ $X2=9.69 $Y2=1.587
r94 32 50 12.4109 $w=3.23e-07 $l=3.5e-07 $layer=LI1_cond $X=9.36 $Y=1.587
+ $X2=9.01 $Y2=1.587
r95 31 50 4.60977 $w=3.23e-07 $l=1.3e-07 $layer=LI1_cond $X=8.88 $Y=1.587
+ $X2=9.01 $Y2=1.587
r96 30 31 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.587
+ $X2=8.88 $Y2=1.587
r97 30 43 14.5385 $w=3.23e-07 $l=4.1e-07 $layer=LI1_cond $X=8.4 $Y=1.587
+ $X2=7.99 $Y2=1.587
r98 29 43 2.48218 $w=3.23e-07 $l=7e-08 $layer=LI1_cond $X=7.92 $Y=1.587 $X2=7.99
+ $Y2=1.587
r99 25 52 23.6381 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.48 $Y=1.345
+ $X2=9.48 $Y2=1.535
r100 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=9.48 $Y=1.345 $X2=9.48
+ $Y2=0.745
r101 22 51 23.6381 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.19 $Y=1.725
+ $X2=9.19 $Y2=1.535
r102 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.19 $Y=1.725
+ $X2=9.19 $Y2=2.465
r103 18 47 23.6381 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.98 $Y=1.345
+ $X2=8.98 $Y2=1.535
r104 18 20 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.98 $Y=1.345 $X2=8.98
+ $Y2=0.745
r105 15 46 23.6381 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.76 $Y=1.725
+ $X2=8.76 $Y2=1.535
r106 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.76 $Y=1.725
+ $X2=8.76 $Y2=2.465
r107 11 45 23.6381 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.53 $Y=1.345
+ $X2=8.53 $Y2=1.535
r108 11 13 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.53 $Y=1.345 $X2=8.53
+ $Y2=0.745
r109 8 44 23.6381 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.33 $Y=1.725
+ $X2=8.33 $Y2=1.535
r110 8 10 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.33 $Y=1.725
+ $X2=8.33 $Y2=2.465
r111 4 40 23.6381 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.98 $Y=1.345
+ $X2=7.98 $Y2=1.535
r112 4 6 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.98 $Y=1.345 $X2=7.98
+ $Y2=0.745
r113 1 39 23.6381 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=7.9 $Y=1.725 $X2=7.9
+ $Y2=1.535
r114 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.9 $Y=1.725 $X2=7.9
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%A_30_367# 1 2 3 4 5 18 22 23 26 30 34 38 42
+ 44 48 50 51 52
r76 46 48 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=3.75 $Y=1.775
+ $X2=3.75 $Y2=1.98
r77 45 52 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.95 $Y=1.69
+ $X2=2.855 $Y2=1.69
r78 44 46 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.62 $Y=1.69
+ $X2=3.75 $Y2=1.775
r79 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.62 $Y=1.69
+ $X2=2.95 $Y2=1.69
r80 40 52 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=1.775
+ $X2=2.855 $Y2=1.69
r81 40 42 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=2.855 $Y=1.775
+ $X2=2.855 $Y2=1.98
r82 39 51 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.09 $Y=1.69
+ $X2=1.995 $Y2=1.69
r83 38 52 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.76 $Y=1.69
+ $X2=2.855 $Y2=1.69
r84 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.76 $Y=1.69
+ $X2=2.09 $Y2=1.69
r85 34 36 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.995 $Y=1.98
+ $X2=1.995 $Y2=2.91
r86 32 51 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=1.775
+ $X2=1.995 $Y2=1.69
r87 32 34 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=1.995 $Y=1.775
+ $X2=1.995 $Y2=1.98
r88 31 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.23 $Y=1.69
+ $X2=1.135 $Y2=1.69
r89 30 51 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.9 $Y=1.69 $X2=1.995
+ $Y2=1.69
r90 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.9 $Y=1.69 $X2=1.23
+ $Y2=1.69
r91 26 28 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.135 $Y=1.98
+ $X2=1.135 $Y2=2.91
r92 24 50 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=1.775
+ $X2=1.135 $Y2=1.69
r93 24 26 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=1.135 $Y=1.775
+ $X2=1.135 $Y2=1.98
r94 22 50 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.04 $Y=1.69
+ $X2=1.135 $Y2=1.69
r95 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.04 $Y=1.69
+ $X2=0.37 $Y2=1.69
r96 18 20 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.24 $Y=1.98 $X2=0.24
+ $Y2=2.91
r97 16 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.24 $Y=1.775
+ $X2=0.37 $Y2=1.69
r98 16 18 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=0.24 $Y=1.775
+ $X2=0.24 $Y2=1.98
r99 5 48 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.575
+ $Y=1.835 $X2=3.715 $Y2=1.98
r100 4 42 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.715
+ $Y=1.835 $X2=2.855 $Y2=1.98
r101 3 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=1.995 $Y2=2.91
r102 3 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=1.995 $Y2=1.98
r103 2 28 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.91
r104 2 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=1.98
r105 1 20 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.91
r106 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%VPWR 1 2 3 4 5 6 21 27 33 37 41 43 47 50 51
+ 53 54 55 56 57 59 64 81 82 85 88 91
r137 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r138 88 89 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r139 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 82 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r141 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r142 79 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.14 $Y=3.33
+ $X2=8.975 $Y2=3.33
r143 79 81 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=9.14 $Y=3.33 $X2=9.84
+ $Y2=3.33
r144 78 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r145 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r146 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r147 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r148 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r149 71 72 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r150 69 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=1.565 $Y2=3.33
r151 69 71 278.578 $w=1.68e-07 $l=4.27e-06 $layer=LI1_cond $X=1.73 $Y=3.33 $X2=6
+ $Y2=3.33
r152 68 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r153 68 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r155 65 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.87 $Y=3.33
+ $X2=0.705 $Y2=3.33
r156 65 67 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.87 $Y=3.33
+ $X2=1.2 $Y2=3.33
r157 64 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=3.33
+ $X2=1.565 $Y2=3.33
r158 64 67 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r159 62 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r160 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r161 59 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.54 $Y=3.33
+ $X2=0.705 $Y2=3.33
r162 59 61 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.54 $Y=3.33 $X2=0.24
+ $Y2=3.33
r163 57 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r164 57 89 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r165 55 77 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=7.95 $Y=3.33 $X2=7.92
+ $Y2=3.33
r166 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.95 $Y=3.33
+ $X2=8.115 $Y2=3.33
r167 53 74 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.09 $Y=3.33
+ $X2=6.96 $Y2=3.33
r168 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.09 $Y=3.33
+ $X2=7.255 $Y2=3.33
r169 52 77 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=7.42 $Y=3.33 $X2=7.92
+ $Y2=3.33
r170 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.42 $Y=3.33
+ $X2=7.255 $Y2=3.33
r171 50 71 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.23 $Y=3.33 $X2=6
+ $Y2=3.33
r172 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=3.33
+ $X2=6.395 $Y2=3.33
r173 49 74 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.56 $Y=3.33 $X2=6.96
+ $Y2=3.33
r174 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.56 $Y=3.33
+ $X2=6.395 $Y2=3.33
r175 45 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.975 $Y=3.245
+ $X2=8.975 $Y2=3.33
r176 45 47 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=8.975 $Y=3.245
+ $X2=8.975 $Y2=2.345
r177 44 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=3.33
+ $X2=8.115 $Y2=3.33
r178 43 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.975 $Y2=3.33
r179 43 44 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.28 $Y2=3.33
r180 39 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=3.245
+ $X2=8.115 $Y2=3.33
r181 39 41 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=8.115 $Y=3.245
+ $X2=8.115 $Y2=2.345
r182 35 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.255 $Y=3.245
+ $X2=7.255 $Y2=3.33
r183 35 37 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=7.255 $Y=3.245
+ $X2=7.255 $Y2=2.345
r184 31 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.395 $Y=3.245
+ $X2=6.395 $Y2=3.33
r185 31 33 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.395 $Y=3.245
+ $X2=6.395 $Y2=2.375
r186 27 30 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=1.565 $Y=2.03
+ $X2=1.565 $Y2=2.95
r187 25 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=3.245
+ $X2=1.565 $Y2=3.33
r188 25 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.565 $Y=3.245
+ $X2=1.565 $Y2=2.95
r189 21 24 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=0.705 $Y=2.03
+ $X2=0.705 $Y2=2.95
r190 19 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=3.245
+ $X2=0.705 $Y2=3.33
r191 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.705 $Y=3.245
+ $X2=0.705 $Y2=2.95
r192 6 47 300 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=2 $X=8.835
+ $Y=1.835 $X2=8.975 $Y2=2.345
r193 5 41 300 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=2 $X=7.975
+ $Y=1.835 $X2=8.115 $Y2=2.345
r194 4 37 300 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=2 $X=7.115
+ $Y=1.835 $X2=7.255 $Y2=2.345
r195 3 33 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=6.255
+ $Y=1.835 $X2=6.395 $Y2=2.375
r196 2 30 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=2.95
r197 2 27 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=2.03
r198 1 24 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.95
r199 1 21 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.03
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%A_457_367# 1 2 3 4 13 15 17 21 23 27 29 33
+ 38 39
r56 31 33 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=5.535 $Y=2.905
+ $X2=5.535 $Y2=2.375
r57 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=2.99
+ $X2=4.675 $Y2=2.99
r58 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.37 $Y=2.99
+ $X2=5.535 $Y2=2.905
r59 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.37 $Y=2.99
+ $X2=4.84 $Y2=2.99
r60 25 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.675 $Y=2.905
+ $X2=4.675 $Y2=2.99
r61 25 27 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=4.675 $Y=2.905
+ $X2=4.675 $Y2=2.375
r62 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=2.99
+ $X2=3.285 $Y2=2.99
r63 23 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.51 $Y=2.99
+ $X2=4.675 $Y2=2.99
r64 23 24 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=4.51 $Y=2.99
+ $X2=3.45 $Y2=2.99
r65 19 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=2.905
+ $X2=3.285 $Y2=2.99
r66 19 21 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=3.285 $Y=2.905
+ $X2=3.285 $Y2=2.03
r67 18 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=2.99
+ $X2=2.425 $Y2=2.99
r68 17 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=2.99
+ $X2=3.285 $Y2=2.99
r69 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.12 $Y=2.99
+ $X2=2.59 $Y2=2.99
r70 13 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=2.905
+ $X2=2.425 $Y2=2.99
r71 13 15 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=2.425 $Y=2.905
+ $X2=2.425 $Y2=2.03
r72 4 33 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=5.395
+ $Y=1.835 $X2=5.535 $Y2=2.375
r73 3 27 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=4.535
+ $Y=1.835 $X2=4.675 $Y2=2.375
r74 2 38 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=1.835 $X2=3.285 $Y2=2.95
r75 2 21 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=1.835 $X2=3.285 $Y2=2.03
r76 1 36 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.835 $X2=2.425 $Y2=2.95
r77 1 15 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.835 $X2=2.425 $Y2=2.03
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%Y 1 2 3 4 5 6 7 8 9 29 32 34 35 38 40 44 46
+ 50 52 56 58 62 64 66 70 71 73 75 76 78 81 82 83 91 93 101 106
c139 75 0 1.29791e-19 $X=7.685 $Y=2.005
r140 83 93 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=5.965 $Y=2.02 $X2=5.87
+ $Y2=2.02
r141 83 97 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=5.965 $Y=2.02 $X2=6.06
+ $Y2=2.02
r142 83 106 14.0097 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=5.965 $Y=2.12
+ $X2=5.965 $Y2=2.465
r143 83 97 0.665455 $w=1.98e-07 $l=1.2e-08 $layer=LI1_cond $X=6.072 $Y=2.02
+ $X2=6.06 $Y2=2.02
r144 82 93 19.4091 $w=1.98e-07 $l=3.5e-07 $layer=LI1_cond $X=5.52 $Y=2.02
+ $X2=5.87 $Y2=2.02
r145 82 94 17.7455 $w=1.98e-07 $l=3.2e-07 $layer=LI1_cond $X=5.52 $Y=2.02
+ $X2=5.2 $Y2=2.02
r146 81 91 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=5.105 $Y=2.02 $X2=5.01
+ $Y2=2.02
r147 81 94 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=5.105 $Y=2.02 $X2=5.2
+ $Y2=2.02
r148 81 101 18.6323 $w=3.03e-07 $l=4.5e-07 $layer=LI1_cond $X=5.105 $Y=2.12
+ $X2=5.105 $Y2=2.57
r149 81 91 1.55273 $w=1.98e-07 $l=2.8e-08 $layer=LI1_cond $X=4.982 $Y=2.02
+ $X2=5.01 $Y2=2.02
r150 71 83 36.4891 $w=1.98e-07 $l=6.58e-07 $layer=LI1_cond $X=6.73 $Y=2.02
+ $X2=6.072 $Y2=2.02
r151 71 73 5.28167 $w=1.85e-07 $l=9.5e-08 $layer=LI1_cond $X=6.73 $Y=2.02
+ $X2=6.825 $Y2=2.02
r152 68 81 35.6018 $w=1.98e-07 $l=6.42e-07 $layer=LI1_cond $X=4.34 $Y=2.02
+ $X2=4.982 $Y2=2.02
r153 68 70 1.9681 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=4.34 $Y=2.02 $X2=4.21
+ $Y2=2.02
r154 64 80 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.44 $Y=2.09
+ $X2=9.44 $Y2=2.005
r155 64 66 16.6218 $w=2.58e-07 $l=3.75e-07 $layer=LI1_cond $X=9.44 $Y=2.09
+ $X2=9.44 $Y2=2.465
r156 60 62 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=9.265 $Y=1.085
+ $X2=9.265 $Y2=0.68
r157 59 78 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.64 $Y=2.005
+ $X2=8.545 $Y2=2.005
r158 58 80 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.31 $Y=2.005
+ $X2=9.44 $Y2=2.005
r159 58 59 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.31 $Y=2.005
+ $X2=8.64 $Y2=2.005
r160 54 78 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.545 $Y=2.09
+ $X2=8.545 $Y2=2.005
r161 54 56 21.89 $w=1.88e-07 $l=3.75e-07 $layer=LI1_cond $X=8.545 $Y=2.09
+ $X2=8.545 $Y2=2.465
r162 53 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.43 $Y=1.17
+ $X2=8.265 $Y2=1.17
r163 52 60 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.1 $Y=1.17
+ $X2=9.265 $Y2=1.085
r164 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.1 $Y=1.17
+ $X2=8.43 $Y2=1.17
r165 48 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.265 $Y=1.085
+ $X2=8.265 $Y2=1.17
r166 48 50 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=8.265 $Y=1.085
+ $X2=8.265 $Y2=0.68
r167 47 75 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.78 $Y=2.005
+ $X2=7.685 $Y2=2.005
r168 46 78 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.45 $Y=2.005
+ $X2=8.545 $Y2=2.005
r169 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.45 $Y=2.005
+ $X2=7.78 $Y2=2.005
r170 42 75 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=2.09
+ $X2=7.685 $Y2=2.005
r171 42 44 21.89 $w=1.88e-07 $l=3.75e-07 $layer=LI1_cond $X=7.685 $Y=2.09
+ $X2=7.685 $Y2=2.465
r172 41 73 5.28167 $w=1.85e-07 $l=1.02225e-07 $layer=LI1_cond $X=6.92 $Y=2.005
+ $X2=6.825 $Y2=2.02
r173 40 75 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.59 $Y=2.005
+ $X2=7.685 $Y2=2.005
r174 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.59 $Y=2.005
+ $X2=6.92 $Y2=2.005
r175 36 73 1.24671 $w=1.9e-07 $l=1e-07 $layer=LI1_cond $X=6.825 $Y=2.12
+ $X2=6.825 $Y2=2.02
r176 36 38 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=6.825 $Y=2.12
+ $X2=6.825 $Y2=2.465
r177 34 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.1 $Y=1.17
+ $X2=8.265 $Y2=1.17
r178 34 35 248.241 $w=1.68e-07 $l=3.805e-06 $layer=LI1_cond $X=8.1 $Y=1.17
+ $X2=4.295 $Y2=1.17
r179 30 70 4.4674 $w=2.37e-07 $l=1e-07 $layer=LI1_cond $X=4.21 $Y=2.12 $X2=4.21
+ $Y2=2.02
r180 30 32 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=4.21 $Y=2.12
+ $X2=4.21 $Y2=2.57
r181 29 70 4.4674 $w=2.37e-07 $l=1.10905e-07 $layer=LI1_cond $X=4.187 $Y=1.92
+ $X2=4.21 $Y2=2.02
r182 28 35 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=4.187 $Y=1.255
+ $X2=4.295 $Y2=1.17
r183 28 29 35.6453 $w=2.13e-07 $l=6.65e-07 $layer=LI1_cond $X=4.187 $Y=1.255
+ $X2=4.187 $Y2=1.92
r184 9 80 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=9.265
+ $Y=1.835 $X2=9.405 $Y2=2.005
r185 9 66 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=9.265
+ $Y=1.835 $X2=9.405 $Y2=2.465
r186 8 78 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=8.405
+ $Y=1.835 $X2=8.545 $Y2=2.005
r187 8 56 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=8.405
+ $Y=1.835 $X2=8.545 $Y2=2.465
r188 7 75 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=7.545
+ $Y=1.835 $X2=7.685 $Y2=2.005
r189 7 44 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=7.545
+ $Y=1.835 $X2=7.685 $Y2=2.465
r190 6 73 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=6.685
+ $Y=1.835 $X2=6.825 $Y2=2.005
r191 6 38 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=6.685
+ $Y=1.835 $X2=6.825 $Y2=2.465
r192 5 83 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=5.825
+ $Y=1.835 $X2=5.965 $Y2=2.005
r193 5 106 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=5.825
+ $Y=1.835 $X2=5.965 $Y2=2.465
r194 4 81 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.835 $X2=5.105 $Y2=2.005
r195 4 101 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.835 $X2=5.105 $Y2=2.57
r196 3 70 600 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=1.835 $X2=4.245 $Y2=2.005
r197 3 32 600 $w=1.7e-07 $l=7.95047e-07 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=1.835 $X2=4.245 $Y2=2.57
r198 2 62 91 $w=1.7e-07 $l=4.47856e-07 $layer=licon1_NDIFF $count=2 $X=9.055
+ $Y=0.325 $X2=9.265 $Y2=0.68
r199 1 50 91 $w=1.7e-07 $l=4.47856e-07 $layer=licon1_NDIFF $count=2 $X=8.055
+ $Y=0.325 $X2=8.265 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 38 42 46
+ 50 53 54 55 56 57 59 71 76 83 84 90 93 96 99
r145 99 100 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r146 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r147 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r148 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r149 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r150 84 100 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=5.52 $Y2=0
r151 83 84 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r152 81 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.6 $Y=0 $X2=5.435
+ $Y2=0
r153 81 83 276.62 $w=1.68e-07 $l=4.24e-06 $layer=LI1_cond $X=5.6 $Y=0 $X2=9.84
+ $Y2=0
r154 77 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.575
+ $Y2=0
r155 77 79 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=5.04
+ $Y2=0
r156 76 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=0 $X2=5.435
+ $Y2=0
r157 76 79 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.27 $Y=0 $X2=5.04
+ $Y2=0
r158 75 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r159 75 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r160 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r161 72 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=3.715
+ $Y2=0
r162 72 74 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=4.08
+ $Y2=0
r163 71 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=4.575
+ $Y2=0
r164 71 74 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=4.08
+ $Y2=0
r165 70 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r166 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r167 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r168 67 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r169 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r170 64 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.135
+ $Y2=0
r171 64 66 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.68
+ $Y2=0
r172 63 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r173 63 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r174 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r175 60 87 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r176 60 62 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.72
+ $Y2=0
r177 59 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.135
+ $Y2=0
r178 59 62 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.72
+ $Y2=0
r179 57 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r180 57 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r181 57 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r182 55 69 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.64
+ $Y2=0
r183 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.855
+ $Y2=0
r184 53 66 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.68
+ $Y2=0
r185 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.995
+ $Y2=0
r186 52 69 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r187 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.995
+ $Y2=0
r188 48 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=0.085
+ $X2=5.435 $Y2=0
r189 48 50 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.435 $Y=0.085
+ $X2=5.435 $Y2=0.44
r190 44 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=0.085
+ $X2=4.575 $Y2=0
r191 44 46 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.575 $Y=0.085
+ $X2=4.575 $Y2=0.45
r192 40 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=0.085
+ $X2=3.715 $Y2=0
r193 40 42 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.715 $Y=0.085
+ $X2=3.715 $Y2=0.45
r194 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=2.855
+ $Y2=0
r195 38 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.715
+ $Y2=0
r196 38 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.55 $Y=0 $X2=3.02
+ $Y2=0
r197 34 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0
r198 34 36 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0.545
r199 30 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0
r200 30 32 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0.545
r201 26 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0
r202 26 28 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0.545
r203 22 87 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r204 22 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.38
r205 7 50 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.235 $X2=5.435 $Y2=0.44
r206 6 46 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=4.435
+ $Y=0.235 $X2=4.575 $Y2=0.45
r207 5 42 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=3.575
+ $Y=0.235 $X2=3.715 $Y2=0.45
r208 4 36 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.855 $Y2=0.545
r209 3 32 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=1.855
+ $Y=0.235 $X2=1.995 $Y2=0.545
r210 2 28 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.235 $X2=1.135 $Y2=0.545
r211 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%A_113_47# 1 2 3 4 5 6 7 8 27 29 30 33 35 39
+ 41 45 47 51 53 54 57 63 66 68 70 74
r91 61 63 50.201 $w=1.88e-07 $l=8.6e-07 $layer=LI1_cond $X=6.405 $Y=0.82
+ $X2=7.265 $Y2=0.82
r92 59 74 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.1 $Y=0.82 $X2=5.005
+ $Y2=0.82
r93 59 61 76.177 $w=1.88e-07 $l=1.305e-06 $layer=LI1_cond $X=5.1 $Y=0.82
+ $X2=6.405 $Y2=0.82
r94 55 74 1.14861 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=5.005 $Y=0.725
+ $X2=5.005 $Y2=0.82
r95 55 57 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=5.005 $Y=0.725
+ $X2=5.005 $Y2=0.42
r96 54 72 6.14599 $w=1.97e-07 $l=1.16146e-07 $layer=LI1_cond $X=4.24 $Y=0.83
+ $X2=4.145 $Y2=0.877
r97 53 74 5.40251 $w=1.8e-07 $l=9.98749e-08 $layer=LI1_cond $X=4.91 $Y=0.83
+ $X2=5.005 $Y2=0.82
r98 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.91 $Y=0.83
+ $X2=4.24 $Y2=0.83
r99 49 72 0.936144 $w=1.9e-07 $l=1.32e-07 $layer=LI1_cond $X=4.145 $Y=0.745
+ $X2=4.145 $Y2=0.877
r100 49 51 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=4.145 $Y=0.745
+ $X2=4.145 $Y2=0.42
r101 48 70 4.6098 $w=2.17e-07 $l=9.5e-08 $layer=LI1_cond $X=3.38 $Y=0.877
+ $X2=3.285 $Y2=0.877
r102 47 72 17.725 $w=2.65e-07 $l=3.67e-07 $layer=LI1_cond $X=3.778 $Y=0.877
+ $X2=4.145 $Y2=0.877
r103 47 48 17.3084 $w=2.63e-07 $l=3.98e-07 $layer=LI1_cond $X=3.778 $Y=0.877
+ $X2=3.38 $Y2=0.877
r104 43 70 1.83355 $w=1.9e-07 $l=1.32e-07 $layer=LI1_cond $X=3.285 $Y=0.745
+ $X2=3.285 $Y2=0.877
r105 43 45 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=3.285 $Y=0.745
+ $X2=3.285 $Y2=0.42
r106 42 68 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.52 $Y=0.925
+ $X2=2.425 $Y2=0.925
r107 41 70 4.6098 $w=2.17e-07 $l=1.16555e-07 $layer=LI1_cond $X=3.19 $Y=0.925
+ $X2=3.285 $Y2=0.877
r108 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.19 $Y=0.925
+ $X2=2.52 $Y2=0.925
r109 37 68 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=0.84
+ $X2=2.425 $Y2=0.925
r110 37 39 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=2.425 $Y=0.84
+ $X2=2.425 $Y2=0.42
r111 36 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.66 $Y=0.925
+ $X2=1.565 $Y2=0.925
r112 35 68 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.33 $Y=0.925
+ $X2=2.425 $Y2=0.925
r113 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.33 $Y=0.925
+ $X2=1.66 $Y2=0.925
r114 31 66 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=0.84
+ $X2=1.565 $Y2=0.925
r115 31 33 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=1.565 $Y=0.84
+ $X2=1.565 $Y2=0.42
r116 29 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.47 $Y=0.925
+ $X2=1.565 $Y2=0.925
r117 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.47 $Y=0.925
+ $X2=0.8 $Y2=0.925
r118 25 30 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.705 $Y=0.84
+ $X2=0.8 $Y2=0.925
r119 25 27 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=0.705 $Y=0.84
+ $X2=0.705 $Y2=0.42
r120 8 63 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=7.125
+ $Y=0.325 $X2=7.265 $Y2=0.82
r121 7 61 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=6.265
+ $Y=0.325 $X2=6.405 $Y2=0.82
r122 6 74 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.235 $X2=5.005 $Y2=0.83
r123 6 57 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.235 $X2=5.005 $Y2=0.42
r124 5 72 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.145 $Y2=0.83
r125 5 51 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.005
+ $Y=0.235 $X2=4.145 $Y2=0.42
r126 4 70 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.235 $X2=3.285 $Y2=0.925
r127 4 45 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.235 $X2=3.285 $Y2=0.42
r128 3 68 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=2.285
+ $Y=0.235 $X2=2.425 $Y2=0.925
r129 3 39 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.285
+ $Y=0.235 $X2=2.425 $Y2=0.42
r130 2 66 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=1.425
+ $Y=0.235 $X2=1.565 $Y2=0.925
r131 2 33 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.425
+ $Y=0.235 $X2=1.565 $Y2=0.42
r132 1 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.705 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_4%A_1166_65# 1 2 3 4 5 16 24 28 30 34 37 38
r58 32 34 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=9.73 $Y=0.425
+ $X2=9.73 $Y2=0.47
r59 31 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.93 $Y=0.34
+ $X2=8.765 $Y2=0.34
r60 30 32 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.6 $Y=0.34
+ $X2=9.73 $Y2=0.425
r61 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.6 $Y=0.34 $X2=8.93
+ $Y2=0.34
r62 26 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=0.425
+ $X2=8.765 $Y2=0.34
r63 26 28 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=8.765 $Y=0.425
+ $X2=8.765 $Y2=0.465
r64 25 37 6.7841 $w=2.35e-07 $l=1.94808e-07 $layer=LI1_cond $X=7.93 $Y=0.34
+ $X2=7.765 $Y2=0.405
r65 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.6 $Y=0.34
+ $X2=8.765 $Y2=0.34
r66 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.6 $Y=0.34 $X2=7.93
+ $Y2=0.34
r67 18 21 33.0367 $w=2.98e-07 $l=8.6e-07 $layer=LI1_cond $X=5.975 $Y=0.405
+ $X2=6.835 $Y2=0.405
r68 16 37 6.7841 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=7.6 $Y=0.405
+ $X2=7.765 $Y2=0.405
r69 16 21 29.3873 $w=2.98e-07 $l=7.65e-07 $layer=LI1_cond $X=7.6 $Y=0.405
+ $X2=6.835 $Y2=0.405
r70 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.555
+ $Y=0.325 $X2=9.695 $Y2=0.47
r71 4 28 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=8.605
+ $Y=0.325 $X2=8.765 $Y2=0.465
r72 3 37 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=7.615
+ $Y=0.325 $X2=7.765 $Y2=0.47
r73 2 21 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=6.695
+ $Y=0.325 $X2=6.835 $Y2=0.45
r74 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.83
+ $Y=0.325 $X2=5.975 $Y2=0.45
.ends

