* File: sky130_fd_sc_lp__or4bb_m.spice
* Created: Wed Sep  2 10:33:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4bb_m.pex.spice"
.subckt sky130_fd_sc_lp__or4bb_m  VNB VPB C_N D_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_C_N_M1010_g N_A_27_530#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_196_530#_M1001_d N_D_N_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_336_439#_M1002_d N_A_196_530#_M1002_g N_VGND_M1002_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_27_530#_M1009_g N_A_336_439#_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_336_439#_M1013_d N_B_M1013_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=17.136 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_336_439#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07455 AS=0.0588 PD=0.775 PS=0.7 NRD=21.42 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1012 N_X_M1012_d N_A_336_439#_M1012_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.07455 PD=1.37 PS=0.775 NRD=0 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_C_N_M1011_g N_A_27_530#_M1011_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_196_530#_M1006_d N_D_N_M1006_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_419_439# N_A_196_530#_M1004_g N_A_336_439#_M1004_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 A_491_439# N_A_27_530#_M1005_g A_419_439# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0917 AS=0.0441 PD=1.01 PS=0.63 NRD=76.5936 NRS=23.443 M=1 R=2.8
+ SA=75000.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 A_593_485# N_B_M1007_g A_491_439# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0917 PD=0.63 PS=1.01 NRD=23.443 NRS=76.5936 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g A_593_485# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.08925 AS=0.0441 PD=0.845 PS=0.63 NRD=39.8531 NRS=23.443 M=1 R=2.8
+ SA=75000.9 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_336_439#_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.08925 PD=1.37 PS=0.845 NRD=0 NRS=28.1316 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
c_97 VPB 0 9.03474e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__or4bb_m.pxi.spice"
*
.ends
*
*
