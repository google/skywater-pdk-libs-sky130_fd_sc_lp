* File: sky130_fd_sc_lp__nor2b_m.pxi.spice
* Created: Fri Aug 28 10:54:59 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2B_M%B_N N_B_N_M1003_g N_B_N_M1004_g N_B_N_c_52_n
+ N_B_N_c_57_n B_N B_N B_N B_N B_N N_B_N_c_54_n PM_SKY130_FD_SC_LP__NOR2B_M%B_N
x_PM_SKY130_FD_SC_LP__NOR2B_M%A N_A_M1005_g N_A_c_93_n N_A_c_100_n N_A_M1001_g
+ N_A_c_94_n N_A_c_95_n N_A_c_96_n N_A_c_101_n A A A A N_A_c_98_n
+ PM_SKY130_FD_SC_LP__NOR2B_M%A
x_PM_SKY130_FD_SC_LP__NOR2B_M%A_47_70# N_A_47_70#_M1003_s N_A_47_70#_M1004_s
+ N_A_47_70#_c_153_n N_A_47_70#_M1002_g N_A_47_70#_M1000_g N_A_47_70#_c_160_n
+ N_A_47_70#_c_155_n N_A_47_70#_c_162_n N_A_47_70#_c_163_n N_A_47_70#_c_156_n
+ N_A_47_70#_c_157_n PM_SKY130_FD_SC_LP__NOR2B_M%A_47_70#
x_PM_SKY130_FD_SC_LP__NOR2B_M%VPWR N_VPWR_M1004_d N_VPWR_c_215_n VPWR
+ N_VPWR_c_216_n N_VPWR_c_217_n N_VPWR_c_214_n N_VPWR_c_219_n
+ PM_SKY130_FD_SC_LP__NOR2B_M%VPWR
x_PM_SKY130_FD_SC_LP__NOR2B_M%Y N_Y_M1005_d N_Y_M1000_d N_Y_c_237_n N_Y_c_238_n
+ N_Y_c_239_n N_Y_c_247_n Y Y Y Y Y Y PM_SKY130_FD_SC_LP__NOR2B_M%Y
x_PM_SKY130_FD_SC_LP__NOR2B_M%VGND N_VGND_M1003_d N_VGND_M1002_d N_VGND_c_267_n
+ N_VGND_c_268_n N_VGND_c_269_n N_VGND_c_270_n N_VGND_c_271_n N_VGND_c_272_n
+ VGND N_VGND_c_273_n N_VGND_c_274_n PM_SKY130_FD_SC_LP__NOR2B_M%VGND
cc_1 VNB N_B_N_M1003_g 0.0445423f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.56
cc_2 VNB N_B_N_c_52_n 0.0164237f $X=-0.19 $Y=-0.245 $X2=0.777 $Y2=1.79
cc_3 VNB B_N 0.00420834f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_4 VNB N_B_N_c_54_n 0.0232211f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.435
cc_5 VNB N_A_c_93_n 0.00514649f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.457
cc_6 VNB N_A_c_94_n 0.0194655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_c_95_n 0.0250611f $X=-0.19 $Y=-0.245 $X2=0.777 $Y2=1.79
cc_8 VNB N_A_c_96_n 0.0172243f $X=-0.19 $Y=-0.245 $X2=0.777 $Y2=1.94
cc_9 VNB A 0.00264092f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_10 VNB N_A_c_98_n 0.0176843f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.27
cc_11 VNB N_A_47_70#_c_153_n 0.0141362f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.67
cc_12 VNB N_A_47_70#_M1002_g 0.043225f $X=-0.19 $Y=-0.245 $X2=0.777 $Y2=1.79
cc_13 VNB N_A_47_70#_c_155_n 0.0421907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_47_70#_c_156_n 9.54519e-19 $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.27
cc_15 VNB N_A_47_70#_c_157_n 0.021299f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.555
cc_16 VNB N_VPWR_c_214_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_237_n 6.55785e-19 $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.67
cc_18 VNB N_Y_c_238_n 0.00730591f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.67
cc_19 VNB N_Y_c_239_n 0.00530539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB Y 0.0119972f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_21 VNB Y 0.031984f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_22 VNB N_VGND_c_267_n 0.00781271f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.67
cc_23 VNB N_VGND_c_268_n 0.0105404f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_24 VNB N_VGND_c_269_n 0.0312063f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_25 VNB N_VGND_c_270_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_26 VNB N_VGND_c_271_n 0.0202814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_272_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_273_n 0.0131219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_274_n 0.175778f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.295
cc_30 VPB N_B_N_M1004_g 0.0453237f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.67
cc_31 VPB N_B_N_c_52_n 0.0115859f $X=-0.19 $Y=1.655 $X2=0.777 $Y2=1.79
cc_32 VPB N_B_N_c_57_n 0.0364148f $X=-0.19 $Y=1.655 $X2=0.777 $Y2=1.94
cc_33 VPB B_N 0.00467776f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_34 VPB N_A_c_93_n 0.0263799f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.457
cc_35 VPB N_A_c_100_n 0.0161998f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.79
cc_36 VPB N_A_c_101_n 0.0279046f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_37 VPB A 0.00480944f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_38 VPB N_A_47_70#_c_153_n 0.00934428f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.67
cc_39 VPB N_A_47_70#_M1000_g 0.0400361f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_40 VPB N_A_47_70#_c_160_n 0.0212328f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_41 VPB N_A_47_70#_c_155_n 0.0321217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_47_70#_c_162_n 0.00419629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_47_70#_c_163_n 0.0317913f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.435
cc_44 VPB N_A_47_70#_c_156_n 0.00308984f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.27
cc_45 VPB N_VPWR_c_215_n 0.0166508f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.79
cc_46 VPB N_VPWR_c_216_n 0.0353157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_217_n 0.0321687f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_48 VPB N_VPWR_c_214_n 0.0767019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_219_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB Y 0.0383688f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_51 N_B_N_c_52_n N_A_c_93_n 0.00660192f $X=0.777 $Y=1.79 $X2=0 $Y2=0
cc_52 N_B_N_c_57_n N_A_c_93_n 0.0176192f $X=0.777 $Y=1.94 $X2=0 $Y2=0
cc_53 B_N N_A_c_93_n 3.4034e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_54 N_B_N_M1004_g N_A_c_100_n 0.0146336f $X=0.98 $Y=2.67 $X2=0 $Y2=0
cc_55 N_B_N_M1003_g N_A_c_94_n 0.00733379f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_56 B_N N_A_c_94_n 0.00347904f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_57 B_N N_A_c_95_n 8.95359e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_58 N_B_N_c_54_n N_A_c_95_n 0.0087395f $X=0.71 $Y=1.435 $X2=0 $Y2=0
cc_59 N_B_N_c_52_n N_A_c_96_n 0.0087395f $X=0.777 $Y=1.79 $X2=0 $Y2=0
cc_60 N_B_N_M1004_g N_A_c_101_n 0.0176192f $X=0.98 $Y=2.67 $X2=0 $Y2=0
cc_61 N_B_N_M1003_g A 5.12028e-19 $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_62 N_B_N_c_52_n A 0.00199273f $X=0.777 $Y=1.79 $X2=0 $Y2=0
cc_63 N_B_N_c_57_n A 0.00287237f $X=0.777 $Y=1.94 $X2=0 $Y2=0
cc_64 B_N A 0.0596628f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_65 N_B_N_c_54_n A 9.99899e-19 $X=0.71 $Y=1.435 $X2=0 $Y2=0
cc_66 N_B_N_M1003_g N_A_c_98_n 0.00911775f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_67 B_N N_A_c_98_n 0.00306928f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_68 N_B_N_M1003_g N_A_47_70#_c_155_n 0.029171f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_69 N_B_N_M1004_g N_A_47_70#_c_155_n 0.0048371f $X=0.98 $Y=2.67 $X2=0 $Y2=0
cc_70 B_N N_A_47_70#_c_155_n 0.104058f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_71 N_B_N_M1004_g N_A_47_70#_c_162_n 0.0140155f $X=0.98 $Y=2.67 $X2=0 $Y2=0
cc_72 N_B_N_M1004_g N_A_47_70#_c_163_n 0.00806715f $X=0.98 $Y=2.67 $X2=0 $Y2=0
cc_73 N_B_N_c_57_n N_A_47_70#_c_163_n 0.00884935f $X=0.777 $Y=1.94 $X2=0 $Y2=0
cc_74 B_N N_A_47_70#_c_163_n 0.0154245f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_75 N_B_N_M1004_g N_VPWR_c_215_n 0.00531583f $X=0.98 $Y=2.67 $X2=0 $Y2=0
cc_76 N_B_N_M1004_g N_VPWR_c_216_n 0.00516473f $X=0.98 $Y=2.67 $X2=0 $Y2=0
cc_77 N_B_N_M1004_g N_VPWR_c_214_n 0.00520574f $X=0.98 $Y=2.67 $X2=0 $Y2=0
cc_78 B_N N_VGND_M1003_d 0.00475422f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_79 N_B_N_M1003_g N_VGND_c_267_n 0.00502529f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_80 B_N N_VGND_c_267_n 0.0132831f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_81 N_B_N_M1003_g N_VGND_c_269_n 0.0045258f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_82 B_N N_VGND_c_269_n 0.00434621f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_83 N_B_N_M1003_g N_VGND_c_274_n 0.00890586f $X=0.575 $Y=0.56 $X2=0 $Y2=0
cc_84 B_N N_VGND_c_274_n 0.0059602f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_85 N_A_c_96_n N_A_47_70#_c_153_n 0.0136247f $X=1.25 $Y=1.55 $X2=0 $Y2=0
cc_86 N_A_c_94_n N_A_47_70#_M1002_g 0.0113451f $X=1.25 $Y=0.88 $X2=0 $Y2=0
cc_87 A N_A_47_70#_M1002_g 0.0016924f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A_c_98_n N_A_47_70#_M1002_g 0.0234965f $X=1.25 $Y=1.045 $X2=0 $Y2=0
cc_89 N_A_c_93_n N_A_47_70#_M1000_g 0.00531448f $X=1.34 $Y=2.2 $X2=0 $Y2=0
cc_90 N_A_c_101_n N_A_47_70#_M1000_g 0.0498977f $X=1.565 $Y=2.275 $X2=0 $Y2=0
cc_91 N_A_c_93_n N_A_47_70#_c_160_n 0.0136247f $X=1.34 $Y=2.2 $X2=0 $Y2=0
cc_92 N_A_c_101_n N_A_47_70#_c_160_n 0.00100631f $X=1.565 $Y=2.275 $X2=0 $Y2=0
cc_93 N_A_c_100_n N_A_47_70#_c_162_n 0.00811985f $X=1.565 $Y=2.35 $X2=0 $Y2=0
cc_94 N_A_c_101_n N_A_47_70#_c_162_n 0.0190042f $X=1.565 $Y=2.275 $X2=0 $Y2=0
cc_95 A N_A_47_70#_c_162_n 0.0171039f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_96 N_A_c_100_n N_A_47_70#_c_163_n 8.0156e-19 $X=1.565 $Y=2.35 $X2=0 $Y2=0
cc_97 N_A_c_93_n N_A_47_70#_c_156_n 0.0027192f $X=1.34 $Y=2.2 $X2=0 $Y2=0
cc_98 N_A_c_95_n N_A_47_70#_c_156_n 0.00201221f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_99 N_A_c_101_n N_A_47_70#_c_156_n 0.00231725f $X=1.565 $Y=2.275 $X2=0 $Y2=0
cc_100 A N_A_47_70#_c_156_n 0.0312602f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_101 N_A_c_95_n N_A_47_70#_c_157_n 0.0136247f $X=1.25 $Y=1.385 $X2=0 $Y2=0
cc_102 A N_A_47_70#_c_157_n 0.0022216f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_103 N_A_c_100_n N_VPWR_c_215_n 0.0075343f $X=1.565 $Y=2.35 $X2=0 $Y2=0
cc_104 N_A_c_101_n N_VPWR_c_215_n 8.99183e-19 $X=1.565 $Y=2.275 $X2=0 $Y2=0
cc_105 N_A_c_100_n N_VPWR_c_217_n 0.00520566f $X=1.565 $Y=2.35 $X2=0 $Y2=0
cc_106 N_A_c_100_n N_VPWR_c_214_n 0.00520574f $X=1.565 $Y=2.35 $X2=0 $Y2=0
cc_107 N_A_c_94_n N_Y_c_237_n 0.00346412f $X=1.25 $Y=0.88 $X2=0 $Y2=0
cc_108 N_A_c_94_n N_Y_c_239_n 2.66831e-19 $X=1.25 $Y=0.88 $X2=0 $Y2=0
cc_109 A N_Y_c_239_n 0.0133285f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_110 N_A_c_98_n N_Y_c_239_n 9.73224e-19 $X=1.25 $Y=1.045 $X2=0 $Y2=0
cc_111 N_A_c_94_n N_Y_c_247_n 0.00367907f $X=1.25 $Y=0.88 $X2=0 $Y2=0
cc_112 N_A_c_94_n N_VGND_c_267_n 0.00340989f $X=1.25 $Y=0.88 $X2=0 $Y2=0
cc_113 A N_VGND_c_267_n 0.00320933f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_114 N_A_c_98_n N_VGND_c_267_n 0.00167293f $X=1.25 $Y=1.045 $X2=0 $Y2=0
cc_115 N_A_c_94_n N_VGND_c_271_n 0.00451107f $X=1.25 $Y=0.88 $X2=0 $Y2=0
cc_116 N_A_c_94_n N_VGND_c_274_n 0.00490041f $X=1.25 $Y=0.88 $X2=0 $Y2=0
cc_117 A N_VGND_c_274_n 0.00628429f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_118 N_A_47_70#_c_162_n N_VPWR_M1004_d 0.00358685f $X=1.705 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_47_70#_c_162_n N_VPWR_c_215_n 0.0233554f $X=1.705 $Y=2.385 $X2=0
+ $Y2=0
cc_120 N_A_47_70#_c_163_n N_VPWR_c_216_n 0.00584962f $X=0.91 $Y=2.385 $X2=0
+ $Y2=0
cc_121 N_A_47_70#_M1000_g N_VPWR_c_217_n 0.00520566f $X=1.925 $Y=2.67 $X2=0
+ $Y2=0
cc_122 N_A_47_70#_M1000_g N_VPWR_c_214_n 0.00520574f $X=1.925 $Y=2.67 $X2=0
+ $Y2=0
cc_123 N_A_47_70#_c_162_n N_VPWR_c_214_n 0.0223611f $X=1.705 $Y=2.385 $X2=0
+ $Y2=0
cc_124 N_A_47_70#_c_163_n N_VPWR_c_214_n 0.0218152f $X=0.91 $Y=2.385 $X2=0 $Y2=0
cc_125 N_A_47_70#_c_162_n A_328_492# 0.00226847f $X=1.705 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_126 N_A_47_70#_M1002_g N_Y_c_237_n 0.00836761f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_127 N_A_47_70#_M1002_g N_Y_c_238_n 0.010153f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_128 N_A_47_70#_c_156_n N_Y_c_238_n 0.0088971f $X=1.79 $Y=1.455 $X2=0 $Y2=0
cc_129 N_A_47_70#_c_157_n N_Y_c_238_n 0.00517662f $X=1.79 $Y=1.455 $X2=0 $Y2=0
cc_130 N_A_47_70#_M1002_g N_Y_c_239_n 0.00381387f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_131 N_A_47_70#_c_157_n N_Y_c_239_n 5.90962e-19 $X=1.79 $Y=1.455 $X2=0 $Y2=0
cc_132 N_A_47_70#_M1002_g N_Y_c_247_n 0.0033503f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_133 N_A_47_70#_M1002_g Y 0.00874092f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_134 N_A_47_70#_c_162_n Y 0.0127049f $X=1.705 $Y=2.385 $X2=0 $Y2=0
cc_135 N_A_47_70#_c_156_n Y 0.069685f $X=1.79 $Y=1.455 $X2=0 $Y2=0
cc_136 N_A_47_70#_c_157_n Y 0.0299866f $X=1.79 $Y=1.455 $X2=0 $Y2=0
cc_137 N_A_47_70#_M1002_g N_VGND_c_268_n 0.00745405f $X=1.715 $Y=0.56 $X2=0
+ $Y2=0
cc_138 N_A_47_70#_c_155_n N_VGND_c_269_n 0.0055846f $X=0.36 $Y=0.625 $X2=0 $Y2=0
cc_139 N_A_47_70#_M1002_g N_VGND_c_271_n 0.0042958f $X=1.715 $Y=0.56 $X2=0 $Y2=0
cc_140 N_A_47_70#_M1002_g N_VGND_c_274_n 0.00490994f $X=1.715 $Y=0.56 $X2=0
+ $Y2=0
cc_141 N_A_47_70#_c_155_n N_VGND_c_274_n 0.00645943f $X=0.36 $Y=0.625 $X2=0
+ $Y2=0
cc_142 N_VPWR_c_217_n Y 0.00542534f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_143 N_VPWR_c_214_n Y 0.00641516f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_144 N_Y_c_238_n N_VGND_c_268_n 0.0145161f $X=2.055 $Y=0.925 $X2=0 $Y2=0
cc_145 N_Y_c_247_n N_VGND_c_268_n 0.0149539f $X=1.6 $Y=0.555 $X2=0 $Y2=0
cc_146 N_Y_c_247_n N_VGND_c_271_n 0.00842964f $X=1.6 $Y=0.555 $X2=0 $Y2=0
cc_147 N_Y_c_238_n N_VGND_c_274_n 0.00610754f $X=2.055 $Y=0.925 $X2=0 $Y2=0
cc_148 N_Y_c_247_n N_VGND_c_274_n 0.0112338f $X=1.6 $Y=0.555 $X2=0 $Y2=0
cc_149 Y N_VGND_c_274_n 0.00749171f $X=2.075 $Y=0.84 $X2=0 $Y2=0
