* File: sky130_fd_sc_lp__a2bb2o_0.spice
* Created: Wed Sep  2 09:23:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2o_0.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2o_0  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_59_194#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1239 PD=0.7 PS=1.43 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_237_47#_M1009_d N_A1_N_M1009_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0609 AS=0.0588 PD=0.71 PS=0.7 NRD=2.856 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A2_N_M1001_g N_A_237_47#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0861 AS=0.0609 PD=0.83 PS=0.71 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_59_194#_M1006_d N_A_237_47#_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0861 PD=0.7 PS=0.83 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75001.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1007 A_523_47# N_B2_M1007_g N_A_59_194#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_B1_M1008_g A_523_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_59_194#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.138023 AS=0.1696 PD=1.24981 PS=1.81 NRD=17.6906 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1004 A_223_490# N_A1_N_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0905774 PD=0.66 PS=0.820189 NRD=30.4759 NRS=28.1316 M=1 R=2.8
+ SA=75000.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_237_47#_M1010_d N_A2_N_M1010_g A_223_490# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_516_535#_M1011_d N_A_237_47#_M1011_g N_A_59_194#_M1011_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_B2_M1005_g N_A_516_535#_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_516_535#_M1002_d N_B1_M1002_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_94 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a2bb2o_0.pxi.spice"
*
.ends
*
*
