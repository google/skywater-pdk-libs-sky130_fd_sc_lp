* File: sky130_fd_sc_lp__a211o_lp.pex.spice
* Created: Fri Aug 28 09:47:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211O_LP%A1 1 3 7 9 10 15
r30 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.32
+ $Y=1.12 $X2=0.32 $Y2=1.12
r31 9 10 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.305 $Y=1.295
+ $X2=0.305 $Y2=1.665
r32 9 15 5.60215 $w=3.58e-07 $l=1.75e-07 $layer=LI1_cond $X=0.305 $Y=1.295
+ $X2=0.305 $Y2=1.12
r33 5 14 40.8239 $w=4.56e-07 $l=2.30857e-07 $layer=POLY_cond $X=0.575 $Y=0.955
+ $X2=0.417 $Y2=1.12
r34 5 7 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.575 $Y=0.955
+ $X2=0.575 $Y2=0.495
r35 1 14 76.3572 $w=4.56e-07 $l=6.95586e-07 $layer=POLY_cond $X=0.555 $Y=1.75
+ $X2=0.417 $Y2=1.12
r36 1 3 197.521 $w=2.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.555 $Y=1.75
+ $X2=0.555 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_LP%A2 3 6 9 11 12 13 17
r38 17 19 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.335
+ $X2=1.075 $Y2=1.17
r39 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.095
+ $Y=1.335 $X2=1.095 $Y2=1.335
r40 13 18 9.87808 $w=3.83e-07 $l=3.3e-07 $layer=LI1_cond $X=1.122 $Y=1.665
+ $X2=1.122 $Y2=1.335
r41 12 18 1.19734 $w=3.83e-07 $l=4e-08 $layer=LI1_cond $X=1.122 $Y=1.295
+ $X2=1.122 $Y2=1.335
r42 9 11 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.135 $Y=2.545
+ $X2=1.135 $Y2=1.84
r43 6 11 34.9505 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=1.075 $Y=1.655
+ $X2=1.075 $Y2=1.84
r44 5 17 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=1.075 $Y=1.355
+ $X2=1.075 $Y2=1.335
r45 5 6 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=1.075 $Y=1.355 $X2=1.075
+ $Y2=1.655
r46 3 19 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.965 $Y=0.495
+ $X2=0.965 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_LP%B1 1 3 4 6 8 10 15 18 19 23
r48 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.665 $Y=1.295
+ $X2=1.665 $Y2=1.665
r49 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.665
+ $Y=1.335 $X2=1.665 $Y2=1.335
r50 17 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.665 $Y=1.675
+ $X2=1.665 $Y2=1.335
r51 14 23 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=1.665 $Y=0.93
+ $X2=1.665 $Y2=1.335
r52 14 15 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.665 $Y=0.855
+ $X2=1.755 $Y2=0.855
r53 11 14 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.395 $Y=0.855
+ $X2=1.665 $Y2=0.855
r54 8 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.755 $Y=0.78
+ $X2=1.755 $Y2=0.855
r55 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.755 $Y=0.78
+ $X2=1.755 $Y2=0.495
r56 4 17 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.84
+ $X2=1.665 $Y2=1.675
r57 4 6 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.665 $Y=1.84
+ $X2=1.665 $Y2=2.545
r58 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=0.78
+ $X2=1.395 $Y2=0.855
r59 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.395 $Y=0.78 $X2=1.395
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_LP%C1 3 7 11 17 20 21 22 26
r50 21 22 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.222 $Y=1.295
+ $X2=2.222 $Y2=1.665
r51 21 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.235
+ $Y=1.335 $X2=2.235 $Y2=1.335
r52 19 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.235 $Y=1.675
+ $X2=2.235 $Y2=1.335
r53 19 20 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.675
+ $X2=2.235 $Y2=1.84
r54 16 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.235 $Y=1.32
+ $X2=2.235 $Y2=1.335
r55 16 17 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=2.235 $Y=1.245
+ $X2=2.545 $Y2=1.245
r56 13 16 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=2.185 $Y=1.245
+ $X2=2.235 $Y2=1.245
r57 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.545 $Y=1.17
+ $X2=2.545 $Y2=1.245
r58 9 11 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.545 $Y=1.17
+ $X2=2.545 $Y2=0.495
r59 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.185 $Y=1.17
+ $X2=2.185 $Y2=1.245
r60 5 7 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.185 $Y=1.17
+ $X2=2.185 $Y2=0.495
r61 3 20 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.195 $Y=2.545
+ $X2=2.195 $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_LP%A_43_57# 1 2 3 10 12 15 17 19 20 24 26 32
+ 34 35 36 37 39 41 43 46 47
r94 46 49 65.7961 $w=5.35e-07 $l=5.05e-07 $layer=POLY_cond $X=3.142 $Y=0.985
+ $X2=3.142 $Y2=1.49
r95 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.04
+ $Y=0.985 $X2=3.04 $Y2=0.985
r96 39 47 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.96 $Y=2.02
+ $X2=2.96 $Y2=1.49
r97 37 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=1.325
+ $X2=3.04 $Y2=1.49
r98 36 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=0.99 $X2=3.04
+ $Y2=0.905
r99 36 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.04 $Y=0.99
+ $X2=3.04 $Y2=1.325
r100 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.875 $Y=2.105
+ $X2=2.96 $Y2=2.02
r101 34 35 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.875 $Y=2.105
+ $X2=2.625 $Y2=2.105
r102 30 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.46 $Y=2.19
+ $X2=2.625 $Y2=2.105
r103 30 32 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.46 $Y=2.19
+ $X2=2.46 $Y2=2.9
r104 27 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0.905
+ $X2=1.97 $Y2=0.905
r105 26 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0.905
+ $X2=3.04 $Y2=0.905
r106 26 27 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.875 $Y=0.905
+ $X2=2.135 $Y2=0.905
r107 22 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=0.82
+ $X2=1.97 $Y2=0.905
r108 22 24 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.97 $Y=0.82
+ $X2=1.97 $Y2=0.495
r109 21 41 14.5407 $w=3.44e-07 $l=5.47083e-07 $layer=LI1_cond $X=0.835 $Y=0.905
+ $X2=0.515 $Y2=0.495
r110 20 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0.905
+ $X2=1.97 $Y2=0.905
r111 20 21 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.805 $Y=0.905
+ $X2=0.835 $Y2=0.905
r112 17 46 31.8222 $w=2.67e-07 $l=2.62857e-07 $layer=POLY_cond $X=3.335 $Y=0.82
+ $X2=3.142 $Y2=0.985
r113 17 19 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.335 $Y=0.82
+ $X2=3.335 $Y2=0.495
r114 15 49 262.119 $w=2.5e-07 $l=1.055e-06 $layer=POLY_cond $X=3.285 $Y=2.545
+ $X2=3.285 $Y2=1.49
r115 10 46 31.8222 $w=2.67e-07 $l=2.35465e-07 $layer=POLY_cond $X=2.975 $Y=0.82
+ $X2=3.142 $Y2=0.985
r116 10 12 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.975 $Y=0.82
+ $X2=2.975 $Y2=0.495
r117 3 32 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=2.045 $X2=2.46 $Y2=2.9
r118 3 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=2.045 $X2=2.46 $Y2=2.19
r119 2 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.83
+ $Y=0.285 $X2=1.97 $Y2=0.495
r120 1 41 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.285 $X2=0.36 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_LP%A_29_409# 1 2 11 13 14 19
r30 17 19 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.4 $Y=2.19 $X2=1.4
+ $Y2=2.9
r31 13 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.235 $Y=2.105
+ $X2=1.4 $Y2=2.19
r32 13 14 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.235 $Y=2.105
+ $X2=0.455 $Y2=2.105
r33 9 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.29 $Y=2.19
+ $X2=0.455 $Y2=2.105
r34 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.29 $Y=2.19 $X2=0.29
+ $Y2=2.9
r35 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.26
+ $Y=2.045 $X2=1.4 $Y2=2.9
r36 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.26
+ $Y=2.045 $X2=1.4 $Y2=2.19
r37 1 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=2.045 $X2=0.29 $Y2=2.9
r38 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=2.045 $X2=0.29 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_LP%VPWR 1 2 11 15 18 19 20 30 31 34
r38 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r40 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r41 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.82 $Y2=3.33
r46 22 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 18 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.02 $Y2=3.33
r51 17 30 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.02 $Y2=3.33
r53 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=3.33
r54 13 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=2.535
r55 9 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245 $X2=0.82
+ $Y2=3.33
r56 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.82 $Y=3.245 $X2=0.82
+ $Y2=2.535
r57 2 15 300 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_PDIFF $count=2 $X=2.875
+ $Y=2.045 $X2=3.02 $Y2=2.535
r58 1 11 300 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=2 $X=0.68
+ $Y=2.045 $X2=0.82 $Y2=2.535
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_LP%X 1 2 7 8 9 10 11 12 13
r16 13 40 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.55 $Y=2.775
+ $X2=3.55 $Y2=2.9
r17 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.55 $Y=2.405
+ $X2=3.55 $Y2=2.775
r18 12 34 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.55 $Y=2.405
+ $X2=3.55 $Y2=2.19
r19 11 34 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.55 $Y=2.035
+ $X2=3.55 $Y2=2.19
r20 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=2.035
r21 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.55 $Y=1.295
+ $X2=3.55 $Y2=1.665
r22 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.55 $Y=0.925 $X2=3.55
+ $Y2=1.295
r23 7 8 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.55 $Y=0.495 $X2=3.55
+ $Y2=0.925
r24 2 40 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.045 $X2=3.55 $Y2=2.9
r25 2 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.045 $X2=3.55 $Y2=2.19
r26 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.285 $X2=3.55 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r50 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r51 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r53 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r54 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=2.76
+ $Y2=0
r55 27 29 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.6
+ $Y2=0
r56 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r57 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r58 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.18
+ $Y2=0
r59 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.68
+ $Y2=0
r60 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.76
+ $Y2=0
r61 22 25 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=1.68
+ $Y2=0
r62 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r63 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r64 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.18
+ $Y2=0
r65 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.72
+ $Y2=0
r66 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r67 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r68 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0
r69 11 13 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0.45
r70 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085 $X2=1.18
+ $Y2=0
r71 7 9 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.45
r72 2 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.285 $X2=2.76 $Y2=0.45
r73 1 9 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.285 $X2=1.18 $Y2=0.45
.ends

