* File: sky130_fd_sc_lp__and2_0.pex.spice
* Created: Wed Sep  2 09:30:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2_0%A 2 5 9 11 12 13 14 19
r34 19 21 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.512 $Y=1.375
+ $X2=0.512 $Y2=1.21
r35 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.46
+ $Y=1.375 $X2=0.46 $Y2=1.375
r36 13 14 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=2.035
r37 13 20 7.54049 $w=4.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=1.375
r38 12 20 2.08014 $w=4.58e-07 $l=8e-08 $layer=LI1_cond $X=0.315 $Y=1.295
+ $X2=0.315 $Y2=1.375
r39 9 11 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=0.655 $Y=2.605
+ $X2=0.655 $Y2=1.88
r40 5 21 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.655 $Y=0.445
+ $X2=0.655 $Y2=1.21
r41 2 11 53.1843 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=0.512 $Y=1.663
+ $X2=0.512 $Y2=1.88
r42 1 19 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=0.512 $Y=1.427
+ $X2=0.512 $Y2=1.375
r43 1 2 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=0.512 $Y=1.427
+ $X2=0.512 $Y2=1.663
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_0%B 3 6 9 11 12 13 17
c39 3 0 1.56886e-19 $X=1.015 $Y=0.445
r40 17 19 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.132 $Y=1.7
+ $X2=1.132 $Y2=1.535
r41 12 13 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.235 $Y=1.665
+ $X2=1.235 $Y2=2.035
r42 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16 $Y=1.7
+ $X2=1.16 $Y2=1.7
r43 9 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.085 $Y=2.605
+ $X2=1.085 $Y2=2.205
r44 6 11 41.2193 $w=3.85e-07 $l=1.92e-07 $layer=POLY_cond $X=1.132 $Y=2.013
+ $X2=1.132 $Y2=2.205
r45 5 17 3.9003 $w=3.85e-07 $l=2.7e-08 $layer=POLY_cond $X=1.132 $Y=1.727
+ $X2=1.132 $Y2=1.7
r46 5 6 41.3143 $w=3.85e-07 $l=2.86e-07 $layer=POLY_cond $X=1.132 $Y=1.727
+ $X2=1.132 $Y2=2.013
r47 3 19 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=1.015 $Y=0.445
+ $X2=1.015 $Y2=1.535
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_0%A_63_47# 1 2 7 9 10 12 16 20 21 22 24 31 32
r63 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=0.93 $X2=1.73 $Y2=0.93
r64 31 32 8.36808 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.847 $Y=2.605
+ $X2=0.847 $Y2=2.44
r65 25 36 28.6003 $w=5.73e-07 $l=3.4e-07 $layer=POLY_cond $X=1.687 $Y=1.27
+ $X2=1.687 $Y2=0.93
r66 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.27 $X2=1.73 $Y2=1.27
r67 22 35 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=1.015 $X2=1.73
+ $Y2=0.93
r68 22 24 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.73 $Y=1.015
+ $X2=1.73 $Y2=1.27
r69 21 29 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.895 $Y=0.93
+ $X2=0.805 $Y2=0.93
r70 20 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=0.93
+ $X2=1.73 $Y2=0.93
r71 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=0.93
+ $X2=0.895 $Y2=0.93
r72 18 29 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=1.015
+ $X2=0.805 $Y2=0.93
r73 18 32 87.803 $w=1.78e-07 $l=1.425e-06 $layer=LI1_cond $X=0.805 $Y=1.015
+ $X2=0.805 $Y2=2.44
r74 14 29 23.0299 $w=1.68e-07 $l=3.53e-07 $layer=LI1_cond $X=0.452 $Y=0.93
+ $X2=0.805 $Y2=0.93
r75 14 16 15.114 $w=3.03e-07 $l=4e-07 $layer=LI1_cond $X=0.452 $Y=0.845
+ $X2=0.452 $Y2=0.445
r76 10 25 43.8576 $w=5.73e-07 $l=2.36525e-07 $layer=POLY_cond $X=1.855 $Y=1.435
+ $X2=1.687 $Y2=1.27
r77 10 12 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=1.855 $Y=1.435
+ $X2=1.855 $Y2=2.715
r78 7 36 43.8576 $w=5.73e-07 $l=3.13838e-07 $layer=POLY_cond $X=1.445 $Y=0.765
+ $X2=1.687 $Y2=0.93
r79 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.445 $Y=0.765
+ $X2=1.445 $Y2=0.445
r80 2 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.73
+ $Y=2.395 $X2=0.87 $Y2=2.605
r81 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.315
+ $Y=0.235 $X2=0.44 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_0%VPWR 1 2 9 11 15 18 19 20 27 28 31
r29 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r30 28 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r31 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 25 31 12.7338 $w=1.7e-07 $l=3.08e-07 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=1.457 $Y2=3.33
r33 25 27 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.765 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 20 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 20 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 20 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 18 23 2.51176 $w=1.7e-07 $l=3.5e-08 $layer=LI1_cond $X=0.275 $Y=3.33
+ $X2=0.24 $Y2=3.33
r39 18 19 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.275 $Y=3.33
+ $X2=0.41 $Y2=3.33
r40 13 31 2.57756 $w=6.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.457 $Y=3.245
+ $X2=1.457 $Y2=3.33
r41 13 15 13.5167 $w=6.13e-07 $l=6.95e-07 $layer=LI1_cond $X=1.457 $Y=3.245
+ $X2=1.457 $Y2=2.55
r42 12 19 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.41 $Y2=3.33
r43 11 31 12.7338 $w=1.7e-07 $l=3.07e-07 $layer=LI1_cond $X=1.15 $Y=3.33
+ $X2=1.457 $Y2=3.33
r44 11 12 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.15 $Y=3.33
+ $X2=0.545 $Y2=3.33
r45 7 19 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.41 $Y=3.245
+ $X2=0.41 $Y2=3.33
r46 7 9 27.3172 $w=2.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.41 $Y=3.245 $X2=0.41
+ $Y2=2.605
r47 2 15 400 $w=1.7e-07 $l=5.52087e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=2.395 $X2=1.64 $Y2=2.55
r48 2 15 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=2.395 $X2=1.3 $Y2=2.55
r49 1 9 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=2.395 $X2=0.44 $Y2=2.605
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_0%X 1 2 7 8 9 10 11 12 13 14 24 30 48
c25 24 0 1.56886e-19 $X=2.065 $Y=0.477
r26 48 49 1.95568 $w=3.78e-07 $l=2e-08 $layer=LI1_cond $X=2.125 $Y=2.405
+ $X2=2.125 $Y2=2.385
r27 41 52 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.125 $Y=2.575
+ $X2=2.125 $Y2=2.55
r28 14 41 6.06549 $w=3.78e-07 $l=2e-07 $layer=LI1_cond $X=2.125 $Y=2.775
+ $X2=2.125 $Y2=2.575
r29 13 52 3.427 $w=3.78e-07 $l=1.13e-07 $layer=LI1_cond $X=2.125 $Y=2.437
+ $X2=2.125 $Y2=2.55
r30 13 48 0.970478 $w=3.78e-07 $l=3.2e-08 $layer=LI1_cond $X=2.125 $Y=2.437
+ $X2=2.125 $Y2=2.405
r31 13 49 1.52122 $w=2.48e-07 $l=3.3e-08 $layer=LI1_cond $X=2.19 $Y=2.352
+ $X2=2.19 $Y2=2.385
r32 12 13 14.613 $w=2.48e-07 $l=3.17e-07 $layer=LI1_cond $X=2.19 $Y=2.035
+ $X2=2.19 $Y2=2.352
r33 11 12 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.19 $Y=1.665
+ $X2=2.19 $Y2=2.035
r34 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.19 $Y=1.295
+ $X2=2.19 $Y2=1.665
r35 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.19 $Y=0.925
+ $X2=2.19 $Y2=1.295
r36 9 30 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.19 $Y=0.925
+ $X2=2.19 $Y2=0.675
r37 8 30 4.45921 $w=2.5e-07 $l=1.98e-07 $layer=LI1_cond $X=2.19 $Y=0.477
+ $X2=2.19 $Y2=0.675
r38 8 24 2.81516 $w=3.95e-07 $l=1.25e-07 $layer=LI1_cond $X=2.19 $Y=0.477
+ $X2=2.065 $Y2=0.477
r39 7 24 11.2327 $w=3.93e-07 $l=3.85e-07 $layer=LI1_cond $X=1.68 $Y=0.477
+ $X2=2.065 $Y2=0.477
r40 7 26 0.583515 $w=3.93e-07 $l=2e-08 $layer=LI1_cond $X=1.68 $Y=0.477 $X2=1.66
+ $Y2=0.477
r41 2 52 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=2.395 $X2=2.07 $Y2=2.55
r42 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.235 $X2=1.66 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_0%VGND 1 6 8 10 17 18 21
r27 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r28 15 21 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.207
+ $Y2=0
r29 15 17 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=2.16
+ $Y2=0
r30 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r31 10 21 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.207
+ $Y2=0
r32 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r33 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r34 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r35 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r36 4 21 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.207 $Y=0.085
+ $X2=1.207 $Y2=0
r37 4 6 14.5572 $w=2.83e-07 $l=3.6e-07 $layer=LI1_cond $X=1.207 $Y=0.085
+ $X2=1.207 $Y2=0.445
r38 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.445
.ends

