* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 a_1275_367# a_762_107# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND a_1275_367# GCLK VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR a_1275_367# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_110_468# GATE a_134_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VPWR a_252_361# a_335_70# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_634_133# a_252_361# a_720_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_720_463# a_762_107# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND SCE a_134_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_252_361# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 GCLK a_1275_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR SCE a_110_468# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_1216_47# a_762_107# a_1275_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VGND a_252_361# a_335_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_720_133# a_762_107# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND a_1275_367# GCLK VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_252_361# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_134_70# a_335_70# a_634_133# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_634_133# a_335_70# a_720_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_1275_367# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 GCLK a_1275_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 GCLK a_1275_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 VGND CLK a_1216_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_134_70# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR a_634_133# a_762_107# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_134_70# a_252_361# a_634_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_634_133# a_762_107# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 VPWR CLK a_1275_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 GCLK a_1275_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
