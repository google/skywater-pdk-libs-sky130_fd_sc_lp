# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nor2_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nor2_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.500000 1.415000 2.245000 1.770000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.415000 1.425000 7.100000 1.750000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  3.292800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.680000 0.315000 0.885000 1.075000 ;
        RECT 0.680000 1.075000 2.605000 1.210000 ;
        RECT 0.680000 1.210000 4.325000 1.245000 ;
        RECT 1.555000 0.315000 1.745000 1.075000 ;
        RECT 2.415000 0.305000 2.605000 1.075000 ;
        RECT 2.425000 1.245000 4.325000 1.360000 ;
        RECT 2.425000 1.360000 5.245000 1.485000 ;
        RECT 3.275000 0.305000 3.465000 1.210000 ;
        RECT 4.065000 1.485000 5.245000 1.920000 ;
        RECT 4.065000 1.920000 7.595000 2.090000 ;
        RECT 4.065000 2.090000 4.395000 2.735000 ;
        RECT 4.135000 0.305000 4.325000 1.210000 ;
        RECT 4.925000 2.090000 5.255000 2.735000 ;
        RECT 4.995000 0.305000 5.185000 1.085000 ;
        RECT 4.995000 1.085000 7.595000 1.255000 ;
        RECT 4.995000 1.255000 5.245000 1.360000 ;
        RECT 5.785000 2.090000 6.115000 2.725000 ;
        RECT 5.855000 0.305000 6.045000 1.085000 ;
        RECT 6.645000 2.090000 6.975000 2.725000 ;
        RECT 6.715000 0.305000 6.905000 1.085000 ;
        RECT 7.425000 1.255000 7.595000 1.920000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.680000 0.085000 ;
        RECT 0.185000  0.085000 0.510000 1.185000 ;
        RECT 1.055000  0.085000 1.385000 0.905000 ;
        RECT 1.915000  0.085000 2.245000 0.905000 ;
        RECT 2.775000  0.085000 3.105000 1.040000 ;
        RECT 3.635000  0.085000 3.965000 1.040000 ;
        RECT 4.495000  0.085000 4.825000 1.190000 ;
        RECT 5.355000  0.085000 5.685000 0.915000 ;
        RECT 6.215000  0.085000 6.545000 0.915000 ;
        RECT 7.075000  0.085000 7.405000 0.915000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.680000 3.415000 ;
        RECT 0.625000 2.280000 0.955000 3.245000 ;
        RECT 1.485000 2.280000 1.815000 3.245000 ;
        RECT 2.345000 2.280000 2.675000 3.245000 ;
        RECT 3.205000 2.095000 3.535000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.185000 1.940000 3.035000 2.110000 ;
      RECT 0.185000 2.110000 0.455000 3.075000 ;
      RECT 1.125000 2.110000 1.315000 3.075000 ;
      RECT 1.985000 2.110000 2.175000 3.075000 ;
      RECT 2.830000 1.700000 3.895000 1.925000 ;
      RECT 2.830000 1.925000 3.035000 1.940000 ;
      RECT 2.845000 2.110000 3.035000 3.075000 ;
      RECT 3.705000 1.925000 3.895000 2.905000 ;
      RECT 3.705000 2.905000 7.405000 3.075000 ;
      RECT 4.565000 2.260000 4.755000 2.905000 ;
      RECT 5.425000 2.260000 5.615000 2.895000 ;
      RECT 5.425000 2.895000 7.405000 2.905000 ;
      RECT 6.285000 2.260000 6.475000 2.895000 ;
      RECT 7.145000 2.260000 7.405000 2.895000 ;
  END
END sky130_fd_sc_lp__nor2_8
