* File: sky130_fd_sc_lp__a22o_1.spice
* Created: Fri Aug 28 09:54:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22o_1.pex.spice"
.subckt sky130_fd_sc_lp__a22o_1  VNB VPB B2 B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_80_246#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2898 AS=0.2226 PD=1.53 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1003 A_294_56# N_B2_M1003_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.2898 PD=1.08 PS=1.53 NRD=9.276 NRS=0 M=1 R=5.6 SA=75001 SB=75001.7
+ A=0.126 P=1.98 MULT=1
MM1004 N_A_80_246#_M1004_d N_B1_M1004_g A_294_56# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1008 PD=1.23 PS=1.08 NRD=8.568 NRS=9.276 M=1 R=5.6 SA=75001.4
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1007 A_480_56# N_A1_M1007_g N_A_80_246#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75002
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_480_56# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6 SA=75002.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_A_80_246#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_A_80_246#_M1002_d N_B2_M1002_g N_A_217_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.189 AS=0.3339 PD=1.56 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1005 N_A_217_367#_M1005_d N_B1_M1005_g N_A_80_246#_M1002_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.189 AS=0.189 PD=1.56 PS=1.56 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75000.6
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_217_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.189 PD=1.65 PS=1.56 NRD=9.3772 NRS=3.1126 M=1 R=8.4
+ SA=75001.1 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1000 N_A_217_367#_M1000_d N_A2_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.6 SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_34 VNB 0 3.30696e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__a22o_1.pxi.spice"
*
.ends
*
*
