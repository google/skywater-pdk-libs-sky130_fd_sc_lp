* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__buflp_1 A VGND VNB VPB VPWR X
X0 a_116_367# a_86_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_308_131# A a_86_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A a_308_403# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_116_47# a_86_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 X a_86_21# a_116_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 X a_86_21# a_116_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_308_403# A a_86_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VGND A a_308_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
