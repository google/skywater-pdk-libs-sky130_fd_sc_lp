* File: sky130_fd_sc_lp__bufinv_16.spice
* Created: Fri Aug 28 10:11:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__bufinv_16.pex.spice"
.subckt sky130_fd_sc_lp__bufinv_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_A_63_49#_M1006_d N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75010.6 A=0.126 P=1.98 MULT=1
MM1017 N_A_63_49#_M1017_d N_A_M1017_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75010.1 A=0.126 P=1.98 MULT=1
MM1040 N_A_63_49#_M1017_d N_A_M1040_g N_VGND_M1040_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1365 PD=1.12 PS=1.165 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75009.7 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1040_s N_A_63_49#_M1001_g N_A_413_49#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1365 AS=0.1176 PD=1.165 PS=1.12 NRD=6.42 NRS=0 M=1 R=5.6
+ SA=75001.5 SB=75009.2 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A_63_49#_M1005_g N_A_413_49#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002
+ SB=75008.8 A=0.126 P=1.98 MULT=1
MM1020 N_VGND_M1005_d N_A_63_49#_M1020_g N_A_413_49#_M1020_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75008.4 A=0.126 P=1.98 MULT=1
MM1035 N_VGND_M1035_d N_A_63_49#_M1035_g N_A_413_49#_M1020_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75007.9 A=0.126 P=1.98 MULT=1
MM1037 N_VGND_M1035_d N_A_63_49#_M1037_g N_A_413_49#_M1037_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75007.5 A=0.126 P=1.98 MULT=1
MM1041 N_VGND_M1041_d N_A_63_49#_M1041_g N_A_413_49#_M1037_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.7
+ SB=75007.1 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1041_d N_A_413_49#_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.1
+ SB=75006.6 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_A_413_49#_M1003_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.5
+ SB=75006.2 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1003_d N_A_413_49#_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005 SB=75005.8
+ A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_413_49#_M1013_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.4
+ SB=75005.3 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1013_d N_A_413_49#_M1014_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.8
+ SB=75004.9 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1016_d N_A_413_49#_M1016_g N_Y_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.3
+ SB=75004.5 A=0.126 P=1.98 MULT=1
MM1021 N_VGND_M1016_d N_A_413_49#_M1021_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.7
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1023 N_VGND_M1023_d N_A_413_49#_M1023_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75007.1
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1030 N_VGND_M1023_d N_A_413_49#_M1030_g N_Y_M1030_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75007.5
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1031 N_VGND_M1031_d N_A_413_49#_M1031_g N_Y_M1030_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75008 SB=75002.8
+ A=0.126 P=1.98 MULT=1
MM1032 N_VGND_M1031_d N_A_413_49#_M1032_g N_Y_M1032_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75008.4
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1036 N_VGND_M1036_d N_A_413_49#_M1036_g N_Y_M1032_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75008.8
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1038 N_VGND_M1036_d N_A_413_49#_M1038_g N_Y_M1038_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75009.3
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1044 N_VGND_M1044_d N_A_413_49#_M1044_g N_Y_M1038_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75009.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1045 N_VGND_M1044_d N_A_413_49#_M1045_g N_Y_M1045_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75010.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1048 N_VGND_M1048_d N_A_413_49#_M1048_g N_Y_M1045_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75010.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_A_63_49#_M1008_d N_A_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75010.6 A=0.189 P=2.82 MULT=1
MM1022 N_A_63_49#_M1022_d N_A_M1022_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75010.1 A=0.189 P=2.82 MULT=1
MM1026 N_A_63_49#_M1022_d N_A_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.20475 PD=1.54 PS=1.585 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75001.1
+ SB=75009.7 A=0.189 P=2.82 MULT=1
MM1004 N_A_413_49#_M1004_d N_A_63_49#_M1004_g N_VPWR_M1026_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.20475 PD=1.54 PS=1.585 NRD=0 NRS=3.9006 M=1 R=8.4
+ SA=75001.5 SB=75009.2 A=0.189 P=2.82 MULT=1
MM1010 N_A_413_49#_M1004_d N_A_63_49#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002
+ SB=75008.8 A=0.189 P=2.82 MULT=1
MM1018 N_A_413_49#_M1018_d N_A_63_49#_M1018_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75008.4 A=0.189 P=2.82 MULT=1
MM1033 N_A_413_49#_M1018_d N_A_63_49#_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75007.9 A=0.189 P=2.82 MULT=1
MM1042 N_A_413_49#_M1042_d N_A_63_49#_M1042_g N_VPWR_M1033_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75007.5 A=0.189 P=2.82 MULT=1
MM1049 N_A_413_49#_M1042_d N_A_63_49#_M1049_g N_VPWR_M1049_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75007.1 A=0.189 P=2.82 MULT=1
MM1000 N_Y_M1000_d N_A_413_49#_M1000_g N_VPWR_M1049_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75006.6 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1000_d N_A_413_49#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75006.2 A=0.189 P=2.82 MULT=1
MM1009 N_Y_M1009_d N_A_413_49#_M1009_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005 SB=75005.8
+ A=0.189 P=2.82 MULT=1
MM1012 N_Y_M1009_d N_A_413_49#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.4
+ SB=75005.3 A=0.189 P=2.82 MULT=1
MM1015 N_Y_M1015_d N_A_413_49#_M1015_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.8
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1019 N_Y_M1015_d N_A_413_49#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.3
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1024 N_Y_M1024_d N_A_413_49#_M1024_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.7
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1025 N_Y_M1024_d N_A_413_49#_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.1
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1027 N_Y_M1027_d N_A_413_49#_M1027_g N_VPWR_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.5
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1028 N_Y_M1027_d N_A_413_49#_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008 SB=75002.8
+ A=0.189 P=2.82 MULT=1
MM1029 N_Y_M1029_d N_A_413_49#_M1029_g N_VPWR_M1028_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.4
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1034 N_Y_M1029_d N_A_413_49#_M1034_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.8
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1039 N_Y_M1039_d N_A_413_49#_M1039_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75009.3
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1043 N_Y_M1039_d N_A_413_49#_M1043_g N_VPWR_M1043_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75009.7
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1046 N_Y_M1046_d N_A_413_49#_M1046_g N_VPWR_M1043_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75010.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1047 N_Y_M1046_d N_A_413_49#_M1047_g N_VPWR_M1047_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75010.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX50_noxref VNB VPB NWDIODE A=22.1935 P=27.53
*
.include "sky130_fd_sc_lp__bufinv_16.pxi.spice"
*
.ends
*
*
