* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_480_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND A3 a_480_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_83_23# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR A1 a_1108_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_1108_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_83_23# B1 a_480_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND A2 a_480_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_480_47# A4 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND a_83_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 X a_83_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR a_83_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_480_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VGND A1 a_480_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VPWR a_83_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_652_345# A3 a_907_345# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_83_23# A4 a_652_345# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VGND A4 a_480_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 X a_83_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR B1 a_83_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_907_345# A3 a_652_345# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 X a_83_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_652_345# A4 a_83_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_907_345# A2 a_1108_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 VGND a_83_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_480_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_1108_367# A2 a_907_345# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 X a_83_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_480_47# B1 a_83_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
