* File: sky130_fd_sc_lp__a2111oi_m.spice
* Created: Wed Sep  2 09:17:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111oi_m.pex.spice"
.subckt sky130_fd_sc_lp__a2111oi_m  VNB VPB D1 C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1009 N_Y_M1009_d N_D1_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1596 PD=0.7 PS=1.6 NRD=0 NRS=32.856 M=1 R=2.8 SA=75000.3
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_C1_M1003_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0903 AS=0.0588 PD=0.85 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0903 PD=0.7 PS=0.85 NRD=0 NRS=37.14 M=1 R=2.8 SA=75001.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 A_443_47# N_A1_M1005_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g A_443_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 A_155_533# N_D1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.2058 PD=0.63 PS=1.82 NRD=23.443 NRS=105.533 M=1 R=2.8 SA=75000.4 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1007 A_227_533# N_C1_M1007_g A_155_533# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.8
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_299_533#_M1008_d N_B1_M1008_g A_227_533# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.1
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_299_533#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.105 AS=0.0588 PD=0.92 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1006 N_A_299_533#_M1006_d N_A2_M1006_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.105 PD=1.37 PS=0.92 NRD=0 NRS=93.7917 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_69 VPB 0 1.69038e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a2111oi_m.pxi.spice"
*
.ends
*
*
