* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_304_463# a_28_108# a_603_191# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_804_328# a_28_108# a_1245_128# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 VPWR a_28_108# a_197_108# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_1796_139# a_1245_128# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_1796_139# a_1245_128# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_1245_128# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_1420_128# a_1440_304# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_789_463# a_804_328# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR RESET_B a_603_191# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_28_108# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 VPWR RESET_B a_1440_304# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_1578_128# a_1245_128# a_1440_304# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_1796_139# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_1245_128# a_28_108# a_1420_128# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 Q a_1796_139# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND a_1245_128# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VPWR D a_304_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 VGND a_28_108# a_197_108# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1440_304# a_1245_128# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VGND a_603_191# a_804_328# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_1245_128# a_197_108# a_1398_472# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_28_108# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_762_191# a_804_328# a_848_191# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_423_191# D a_304_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_804_328# a_197_108# a_1245_128# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_1398_472# a_1440_304# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 VGND RESET_B a_1578_128# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_304_463# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_603_191# a_28_108# a_789_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VGND RESET_B a_423_191# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_603_191# a_197_108# a_762_191# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_304_463# a_197_108# a_603_191# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VPWR a_603_191# a_804_328# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X33 a_848_191# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
