* NGSPICE file created from sky130_fd_sc_lp__bufinv_8.ext - technology: sky130A

.subckt sky130_fd_sc_lp__bufinv_8 A VGND VNB VPB VPWR Y
M1000 Y a_82_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.4112e+12p pd=1.232e+07u as=2.4318e+12p ps=2.15e+07u
M1001 VPWR a_876_23# a_82_23# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=6.867e+11p ps=6.13e+06u
M1002 a_82_23# a_876_23# VGND VNB nshort w=840000u l=150000u
+  ad=4.662e+11p pd=4.47e+06u as=1.6212e+12p ps=1.562e+07u
M1003 Y a_82_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_82_23# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=9.408e+11p ps=8.96e+06u
M1005 Y a_82_23# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_82_23# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_82_23# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_876_23# a_82_23# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_82_23# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_82_23# a_876_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_82_23# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_876_23# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1013 VGND a_82_23# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_82_23# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_876_23# a_82_23# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_82_23# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_82_23# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_876_23# A VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1019 Y a_82_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y a_82_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_876_23# a_82_23# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y a_82_23# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_82_23# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

