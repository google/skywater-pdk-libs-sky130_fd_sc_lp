* File: sky130_fd_sc_lp__a32o_1.pex.spice
* Created: Fri Aug 28 10:00:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32O_1%A_80_21# 1 2 7 9 12 15 17 18 19 20 21 24 27
+ 31 38
c90 12 0 8.17141e-21 $X=0.665 $Y=2.465
r91 31 33 9.85006 $w=6.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.58 $Y=0.38
+ $X2=2.58 $Y2=0.94
r92 28 38 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=0.6 $Y=1.35 $X2=0.665
+ $Y2=1.35
r93 28 35 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.6 $Y=1.35
+ $X2=0.475 $Y2=1.35
r94 27 29 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.7 $Y=1.35 $X2=0.7
+ $Y2=1.515
r95 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.35 $X2=0.6 $Y2=1.35
r96 22 24 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.085 $Y=1.875
+ $X2=3.085 $Y2=1.98
r97 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.92 $Y=1.79
+ $X2=3.085 $Y2=1.875
r98 20 21 132.765 $w=1.68e-07 $l=2.035e-06 $layer=LI1_cond $X=2.92 $Y=1.79
+ $X2=0.885 $Y2=1.79
r99 18 33 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=2.24 $Y=0.94 $X2=2.58
+ $Y2=0.94
r100 18 19 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=2.24 $Y=0.94
+ $X2=0.885 $Y2=0.94
r101 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.8 $Y=1.705
+ $X2=0.885 $Y2=1.79
r102 17 29 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.8 $Y=1.705
+ $X2=0.8 $Y2=1.515
r103 15 27 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=0.7 $Y=1.33 $X2=0.7
+ $Y2=1.35
r104 14 19 8.10976 $w=1.7e-07 $l=2.23495e-07 $layer=LI1_cond $X=0.7 $Y=1.025
+ $X2=0.885 $Y2=0.94
r105 14 15 9.49987 $w=3.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.7 $Y=1.025
+ $X2=0.7 $Y2=1.33
r106 10 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.515
+ $X2=0.665 $Y2=1.35
r107 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.665 $Y=1.515
+ $X2=0.665 $Y2=2.465
r108 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=1.35
r109 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.655
r110 2 24 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.835 $X2=3.085 $Y2=1.98
r111 1 31 45.5 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=4 $X=2.265
+ $Y=0.235 $X2=2.755 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_1%A3 3 7 8 11 13
c37 8 0 8.17141e-21 $X=1.2 $Y=1.295
r38 11 14 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.36
+ $X2=1.145 $Y2=1.525
r39 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.36
+ $X2=1.145 $Y2=1.195
r40 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.36 $X2=1.15 $Y2=1.36
r41 7 13 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.24 $Y=0.655 $X2=1.24
+ $Y2=1.195
r42 3 14 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.17 $Y=2.465 $X2=1.17
+ $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_1%A2 3 7 8 11 13
c33 3 0 2.23288e-20 $X=1.6 $Y=2.465
r34 11 14 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.35 $X2=1.7
+ $Y2=1.515
r35 11 13 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.7 $Y=1.35 $X2=1.7
+ $Y2=1.185
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.695
+ $Y=1.35 $X2=1.695 $Y2=1.35
r37 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.705 $Y=0.655
+ $X2=1.705 $Y2=1.185
r38 3 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.6 $Y=2.465 $X2=1.6
+ $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_1%A1 1 3 6 8 14 15
c34 14 0 6.30552e-20 $X=2.28 $Y=1.36
r35 13 15 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.28 $Y=1.36
+ $X2=2.43 $Y2=1.36
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.36 $X2=2.28 $Y2=1.36
r37 10 13 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.19 $Y=1.36 $X2=2.28
+ $Y2=1.36
r38 8 14 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.16 $Y=1.36 $X2=2.28
+ $Y2=1.36
r39 4 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=1.525
+ $X2=2.43 $Y2=1.36
r40 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.43 $Y=1.525 $X2=2.43
+ $Y2=2.465
r41 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.195
+ $X2=2.19 $Y2=1.36
r42 1 3 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.19 $Y=1.195 $X2=2.19
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_1%B1 3 7 8 9 13 15
c32 3 0 1.50208e-19 $X=2.86 $Y=2.465
r33 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.35
+ $X2=2.88 $Y2=1.515
r34 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.35
+ $X2=2.88 $Y2=1.185
r35 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=1.35 $X2=2.88 $Y2=1.35
r36 9 14 8.64332 $w=3.18e-07 $l=2.4e-07 $layer=LI1_cond $X=3.12 $Y=1.355
+ $X2=2.88 $Y2=1.355
r37 8 14 8.64332 $w=3.18e-07 $l=2.4e-07 $layer=LI1_cond $X=2.64 $Y=1.355
+ $X2=2.88 $Y2=1.355
r38 7 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.97 $Y=0.655
+ $X2=2.97 $Y2=1.185
r39 3 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.86 $Y=2.465
+ $X2=2.86 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_1%B2 3 7 9 10 16
c25 9 0 1.09482e-19 $X=3.6 $Y=1.295
r26 13 16 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.33 $Y=1.375
+ $X2=3.555 $Y2=1.375
r27 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=1.295
+ $X2=3.587 $Y2=1.665
r28 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.555
+ $Y=1.375 $X2=3.555 $Y2=1.375
r29 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.54
+ $X2=3.33 $Y2=1.375
r30 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.33 $Y=1.54 $X2=3.33
+ $Y2=2.465
r31 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.21
+ $X2=3.33 $Y2=1.375
r32 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.33 $Y=1.21 $X2=3.33
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_1%X 1 2 7 8 9 10 11 12 13 24 48
r16 46 48 0.53159 $w=4.48e-07 $l=2e-08 $layer=LI1_cond $X=0.32 $Y=2.015 $X2=0.32
+ $Y2=2.035
r17 34 48 1.06318 $w=4.48e-07 $l=4e-08 $layer=LI1_cond $X=0.32 $Y=2.075 $X2=0.32
+ $Y2=2.035
r18 13 41 3.58824 $w=4.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.32 $Y=2.775
+ $X2=0.32 $Y2=2.91
r19 12 13 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=2.405
+ $X2=0.32 $Y2=2.775
r20 11 46 0.0797386 $w=4.48e-07 $l=3e-09 $layer=LI1_cond $X=0.32 $Y=2.012
+ $X2=0.32 $Y2=2.015
r21 11 44 6.65016 $w=4.48e-07 $l=1.62e-07 $layer=LI1_cond $X=0.32 $Y=2.012
+ $X2=0.32 $Y2=1.85
r22 11 12 8.18649 $w=4.48e-07 $l=3.08e-07 $layer=LI1_cond $X=0.32 $Y=2.097
+ $X2=0.32 $Y2=2.405
r23 11 34 0.584749 $w=4.48e-07 $l=2.2e-08 $layer=LI1_cond $X=0.32 $Y=2.097
+ $X2=0.32 $Y2=2.075
r24 10 44 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=1.85
r25 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.665
r26 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.925 $X2=0.22
+ $Y2=1.295
r27 7 8 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.555 $X2=0.22
+ $Y2=0.925
r28 7 24 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=0.555
+ $X2=0.22 $Y2=0.42
r29 2 46 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.45 $Y2=2.015
r30 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.45 $Y2=2.91
r31 1 24 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_1%VPWR 1 2 11 15 19 21 28 29 32 35
r48 35 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 33 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 26 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 26 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 23 35 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.015 $Y2=3.33
r58 23 25 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 21 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 21 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 17 35 2.94957 $w=7.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=3.245
+ $X2=2.015 $Y2=3.33
r62 17 19 12.2066 $w=7.28e-07 $l=7.45e-07 $layer=LI1_cond $X=2.015 $Y=3.245
+ $X2=2.015 $Y2=2.5
r63 16 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.05 $Y=3.33
+ $X2=0.885 $Y2=3.33
r64 15 35 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=2.015 $Y2=3.33
r65 15 16 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.65 $Y=3.33 $X2=1.05
+ $Y2=3.33
r66 11 14 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.885 $Y=2.19
+ $X2=0.885 $Y2=2.95
r67 9 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=3.245
+ $X2=0.885 $Y2=3.33
r68 9 14 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.885 $Y=3.245
+ $X2=0.885 $Y2=2.95
r69 2 19 150 $w=1.7e-07 $l=8.95168e-07 $layer=licon1_PDIFF $count=4 $X=1.675
+ $Y=1.835 $X2=2.215 $Y2=2.5
r70 1 14 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.74
+ $Y=1.835 $X2=0.885 $Y2=2.95
r71 1 11 400 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=0.74
+ $Y=1.835 $X2=0.885 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_1%A_249_367# 1 2 3 10 12 14 17 20 22 24
r29 22 31 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.565 $Y=2.905
+ $X2=3.565 $Y2=2.99
r30 22 24 32.1889 $w=2.88e-07 $l=8.1e-07 $layer=LI1_cond $X=3.565 $Y=2.905
+ $X2=3.565 $Y2=2.095
r31 21 29 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.75 $Y=2.99 $X2=2.65
+ $Y2=2.99
r32 20 31 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.42 $Y=2.99
+ $X2=3.565 $Y2=2.99
r33 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.42 $Y=2.99
+ $X2=2.75 $Y2=2.99
r34 17 29 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=2.905 $X2=2.65
+ $Y2=2.99
r35 17 19 37.9864 $w=1.98e-07 $l=6.85e-07 $layer=LI1_cond $X=2.65 $Y=2.905
+ $X2=2.65 $Y2=2.22
r36 16 19 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=2.65 $Y=2.215
+ $X2=2.65 $Y2=2.22
r37 15 27 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.48 $Y=2.13 $X2=1.35
+ $Y2=2.13
r38 14 16 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.55 $Y=2.13
+ $X2=2.65 $Y2=2.215
r39 14 15 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=2.55 $Y=2.13
+ $X2=1.48 $Y2=2.13
r40 10 27 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=2.215
+ $X2=1.35 $Y2=2.13
r41 10 12 13.7407 $w=2.58e-07 $l=3.1e-07 $layer=LI1_cond $X=1.35 $Y=2.215
+ $X2=1.35 $Y2=2.525
r42 3 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.835 $X2=3.545 $Y2=2.91
r43 3 24 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.835 $X2=3.545 $Y2=2.095
r44 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.835 $X2=2.645 $Y2=2.91
r45 2 19 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.835 $X2=2.645 $Y2=2.22
r46 1 27 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.835 $X2=1.385 $Y2=2.13
r47 1 12 300 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=2 $X=1.245
+ $Y=1.835 $X2=1.385 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_1%VGND 1 2 7 9 11 13 18 28 35
r43 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 28 31 6.99246 $w=6.48e-07 $l=3.8e-07 $layer=LI1_cond $X=0.87 $Y=0 $X2=0.87
+ $Y2=0.38
r45 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r47 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 22 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r49 21 24 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r50 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 19 28 8.83581 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=0.87
+ $Y2=0
r52 19 21 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.2
+ $Y2=0
r53 18 34 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.61
+ $Y2=0
r54 18 24 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.12
+ $Y2=0
r55 16 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r56 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 13 28 8.83581 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.87
+ $Y2=0
r58 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r59 11 25 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r60 11 22 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r61 7 34 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.61 $Y2=0
r62 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0.38
r63 2 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.235 $X2=3.545 $Y2=0.38
r64 1 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

