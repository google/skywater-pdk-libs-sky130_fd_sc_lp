* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21ai_lp A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_155_409# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=5.7e+11p ps=5.14e+06u
M1001 VGND A1 a_64_57# VNB nshort w=420000u l=150000u
+  ad=1.848e+11p pd=1.72e+06u as=2.373e+11p ps=2.81e+06u
M1002 VPWR B1 Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1003 a_64_57# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A2 a_155_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B1 a_64_57# VNB nshort w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=0p ps=0u
.ends
