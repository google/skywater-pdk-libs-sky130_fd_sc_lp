* File: sky130_fd_sc_lp__a221oi_m.pxi.spice
* Created: Fri Aug 28 09:53:46 2020
* 
x_PM_SKY130_FD_SC_LP__A221OI_M%C1 N_C1_M1009_g N_C1_c_74_n N_C1_M1007_g
+ N_C1_c_71_n C1 C1 C1 N_C1_c_73_n PM_SKY130_FD_SC_LP__A221OI_M%C1
x_PM_SKY130_FD_SC_LP__A221OI_M%B2 N_B2_M1001_g N_B2_M1005_g B2 N_B2_c_114_n
+ PM_SKY130_FD_SC_LP__A221OI_M%B2
x_PM_SKY130_FD_SC_LP__A221OI_M%B1 N_B1_M1002_g N_B1_M1003_g N_B1_c_159_n
+ N_B1_c_153_n N_B1_c_161_n N_B1_c_154_n N_B1_c_155_n B1 B1 N_B1_c_157_n
+ N_B1_c_164_n PM_SKY130_FD_SC_LP__A221OI_M%B1
x_PM_SKY130_FD_SC_LP__A221OI_M%A1 N_A1_M1000_g N_A1_M1004_g N_A1_c_219_n
+ N_A1_c_224_n A1 N_A1_c_221_n PM_SKY130_FD_SC_LP__A221OI_M%A1
x_PM_SKY130_FD_SC_LP__A221OI_M%A2 N_A2_c_264_n N_A2_M1006_g N_A2_M1008_g
+ N_A2_c_265_n N_A2_c_270_n A2 A2 N_A2_c_267_n PM_SKY130_FD_SC_LP__A221OI_M%A2
x_PM_SKY130_FD_SC_LP__A221OI_M%Y N_Y_M1009_s N_Y_M1002_d N_Y_M1007_s N_Y_c_313_n
+ N_Y_c_314_n N_Y_c_308_n Y Y Y Y Y N_Y_c_310_n N_Y_c_311_n N_Y_c_312_n
+ PM_SKY130_FD_SC_LP__A221OI_M%Y
x_PM_SKY130_FD_SC_LP__A221OI_M%A_210_535# N_A_210_535#_M1007_d
+ N_A_210_535#_M1003_d N_A_210_535#_c_364_n N_A_210_535#_c_365_n
+ N_A_210_535#_c_366_n N_A_210_535#_c_367_n
+ PM_SKY130_FD_SC_LP__A221OI_M%A_210_535#
x_PM_SKY130_FD_SC_LP__A221OI_M%A_296_535# N_A_296_535#_M1005_d
+ N_A_296_535#_M1008_d N_A_296_535#_c_404_n N_A_296_535#_c_400_n
+ N_A_296_535#_c_401_n N_A_296_535#_c_407_n
+ PM_SKY130_FD_SC_LP__A221OI_M%A_296_535#
x_PM_SKY130_FD_SC_LP__A221OI_M%VPWR N_VPWR_M1000_d N_VPWR_c_425_n VPWR
+ N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_424_n N_VPWR_c_429_n
+ PM_SKY130_FD_SC_LP__A221OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A221OI_M%VGND N_VGND_M1009_d N_VGND_M1006_d N_VGND_c_463_n
+ N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n N_VGND_c_467_n N_VGND_c_468_n
+ VGND N_VGND_c_469_n N_VGND_c_470_n PM_SKY130_FD_SC_LP__A221OI_M%VGND
cc_1 VNB N_C1_M1009_g 0.0577068f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.485
cc_2 VNB N_C1_c_71_n 0.00279723f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.955
cc_3 VNB C1 0.00845633f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C1_c_73_n 0.0171821f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.615
cc_5 VNB N_B2_M1001_g 0.058998f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.485
cc_6 VNB B2 0.00346735f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.885
cc_7 VNB N_B1_M1002_g 0.0306543f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.485
cc_8 VNB N_B1_c_153_n 0.00411784f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.45
cc_9 VNB N_B1_c_154_n 0.00286132f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_10 VNB N_B1_c_155_n 0.0330873f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_11 VNB B1 0.011045f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.615
cc_12 VNB N_B1_c_157_n 0.0323766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1004_g 0.0366644f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.4
cc_14 VNB N_A1_c_219_n 0.00796785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A1 0.00385216f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_16 VNB N_A1_c_221_n 0.0299407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_264_n 0.021054f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.45
cc_18 VNB N_A2_c_265_n 0.0329372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB A2 0.0290634f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.955
cc_20 VNB N_A2_c_267_n 0.0552303f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_21 VNB N_Y_c_308_n 0.0309824f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.325
cc_22 VNB Y 0.00805645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_310_n 0.0175624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_311_n 0.0375227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_312_n 0.00658565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_424_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.615
cc_27 VNB N_VGND_c_463_n 0.00606944f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.885
cc_28 VNB N_VGND_c_464_n 0.00685879f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.955
cc_29 VNB N_VGND_c_465_n 0.0217261f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_30 VNB N_VGND_c_466_n 0.00401244f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_31 VNB N_VGND_c_467_n 0.0415065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_468_n 0.00401309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_469_n 0.0252142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_470_n 0.211838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_C1_c_74_n 0.0263506f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=2.325
cc_36 VPB N_C1_M1007_g 0.0310938f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.885
cc_37 VPB N_C1_c_71_n 0.0594777f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.955
cc_38 VPB C1 0.0066134f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_39 VPB N_B2_M1001_g 0.00152321f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.485
cc_40 VPB N_B2_M1005_g 0.0470221f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.4
cc_41 VPB N_B2_c_114_n 0.0482545f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_42 VPB N_B1_M1003_g 0.051545f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.4
cc_43 VPB N_B1_c_159_n 0.0194826f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_B1_c_153_n 0.00173513f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.45
cc_45 VPB N_B1_c_161_n 0.00370442f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.325
cc_46 VPB B1 0.0156171f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.615
cc_47 VPB N_B1_c_157_n 0.0168471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_B1_c_164_n 0.0163937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A1_M1000_g 0.0571547f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.485
cc_50 VPB N_A1_c_219_n 0.00148239f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A1_c_224_n 0.0174335f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.955
cc_52 VPB N_A2_M1008_g 0.053008f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.325
cc_53 VPB N_A2_c_265_n 0.00544365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A2_c_270_n 0.00971755f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.615
cc_55 VPB N_Y_c_313_n 0.0169439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_Y_c_314_n 0.0168599f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.45
cc_57 VPB N_Y_c_308_n 0.0498715f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.325
cc_58 VPB N_A_210_535#_c_364_n 0.00785228f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.885
cc_59 VPB N_A_210_535#_c_365_n 0.0330811f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.615
cc_60 VPB N_A_210_535#_c_366_n 0.00390674f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.45
cc_61 VPB N_A_210_535#_c_367_n 0.0172421f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_62 VPB N_A_296_535#_c_400_n 0.0144666f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.615
cc_63 VPB N_A_296_535#_c_401_n 0.00346808f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.45
cc_64 VPB N_VPWR_c_425_n 0.00564356f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.325
cc_65 VPB N_VPWR_c_426_n 0.0547576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_427_n 0.0311859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_424_n 0.0505319f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.615
cc_68 VPB N_VPWR_c_429_n 0.00631563f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.295
cc_69 N_C1_M1009_g N_B2_M1001_g 0.0343728f $X=0.625 $Y=0.485 $X2=0 $Y2=0
cc_70 C1 N_B2_M1001_g 0.011129f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_C1_c_74_n N_B2_M1005_g 0.0262547f $X=0.9 $Y=2.325 $X2=0 $Y2=0
cc_72 N_C1_c_71_n N_B2_M1005_g 0.00328431f $X=0.535 $Y=1.955 $X2=0 $Y2=0
cc_73 C1 N_B2_M1005_g 0.00194964f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_C1_c_74_n B2 4.08045e-19 $X=0.9 $Y=2.325 $X2=0 $Y2=0
cc_75 C1 B2 0.0266541f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_C1_c_73_n B2 3.68517e-19 $X=0.535 $Y=1.615 $X2=0 $Y2=0
cc_77 N_C1_c_74_n N_B2_c_114_n 0.00474155f $X=0.9 $Y=2.325 $X2=0 $Y2=0
cc_78 N_C1_c_73_n N_B2_c_114_n 0.0343728f $X=0.535 $Y=1.615 $X2=0 $Y2=0
cc_79 C1 N_B1_c_154_n 0.0050001f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_80 N_C1_M1007_g N_Y_c_314_n 4.64138e-19 $X=0.975 $Y=2.885 $X2=0 $Y2=0
cc_81 N_C1_c_71_n N_Y_c_314_n 0.0114792f $X=0.535 $Y=1.955 $X2=0 $Y2=0
cc_82 C1 N_Y_c_314_n 0.0128703f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 N_C1_M1009_g N_Y_c_308_n 0.00738727f $X=0.625 $Y=0.485 $X2=0 $Y2=0
cc_84 N_C1_M1007_g N_Y_c_308_n 0.00540252f $X=0.975 $Y=2.885 $X2=0 $Y2=0
cc_85 N_C1_c_71_n N_Y_c_308_n 0.00923365f $X=0.535 $Y=1.955 $X2=0 $Y2=0
cc_86 C1 N_Y_c_308_n 0.0668059f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 N_C1_c_73_n N_Y_c_308_n 0.0163648f $X=0.535 $Y=1.615 $X2=0 $Y2=0
cc_88 N_C1_M1009_g N_Y_c_310_n 0.0167454f $X=0.625 $Y=0.485 $X2=0 $Y2=0
cc_89 C1 N_Y_c_310_n 0.0211352f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 N_C1_M1009_g N_Y_c_311_n 0.00513899f $X=0.625 $Y=0.485 $X2=0 $Y2=0
cc_91 C1 N_Y_c_311_n 0.00522615f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_92 N_C1_c_73_n N_Y_c_311_n 0.00316451f $X=0.535 $Y=1.615 $X2=0 $Y2=0
cc_93 N_C1_c_74_n N_A_210_535#_c_364_n 0.00893527f $X=0.9 $Y=2.325 $X2=0 $Y2=0
cc_94 N_C1_c_74_n N_A_210_535#_c_366_n 0.00219856f $X=0.9 $Y=2.325 $X2=0 $Y2=0
cc_95 N_C1_c_71_n N_A_210_535#_c_366_n 0.0024978f $X=0.535 $Y=1.955 $X2=0 $Y2=0
cc_96 N_C1_M1007_g N_VPWR_c_426_n 0.00585385f $X=0.975 $Y=2.885 $X2=0 $Y2=0
cc_97 N_C1_M1007_g N_VPWR_c_424_n 0.0124078f $X=0.975 $Y=2.885 $X2=0 $Y2=0
cc_98 N_C1_M1009_g N_VGND_c_463_n 0.00290284f $X=0.625 $Y=0.485 $X2=0 $Y2=0
cc_99 N_C1_M1009_g N_VGND_c_465_n 0.00406911f $X=0.625 $Y=0.485 $X2=0 $Y2=0
cc_100 N_C1_M1009_g N_VGND_c_470_n 0.00650419f $X=0.625 $Y=0.485 $X2=0 $Y2=0
cc_101 N_B2_M1001_g N_B1_M1002_g 0.0816602f $X=1.055 $Y=0.485 $X2=0 $Y2=0
cc_102 N_B2_M1001_g N_B1_c_153_n 0.00471063f $X=1.055 $Y=0.485 $X2=0 $Y2=0
cc_103 B2 N_B1_c_153_n 0.01237f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B2_c_114_n N_B1_c_153_n 6.40306e-19 $X=1.405 $Y=1.845 $X2=0 $Y2=0
cc_105 B2 N_B1_c_161_n 0.0142412f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_106 N_B2_c_114_n N_B1_c_161_n 0.00309079f $X=1.405 $Y=1.845 $X2=0 $Y2=0
cc_107 N_B2_M1001_g N_B1_c_154_n 6.95913e-19 $X=1.055 $Y=0.485 $X2=0 $Y2=0
cc_108 N_B2_c_114_n N_B1_c_154_n 8.99181e-19 $X=1.405 $Y=1.845 $X2=0 $Y2=0
cc_109 N_B2_c_114_n N_B1_c_155_n 0.00940209f $X=1.405 $Y=1.845 $X2=0 $Y2=0
cc_110 N_B2_M1005_g N_A1_M1000_g 0.0274436f $X=1.405 $Y=2.885 $X2=0 $Y2=0
cc_111 N_B2_c_114_n N_A1_c_224_n 0.0274436f $X=1.405 $Y=1.845 $X2=0 $Y2=0
cc_112 N_B2_M1001_g N_Y_c_310_n 0.0171578f $X=1.055 $Y=0.485 $X2=0 $Y2=0
cc_113 B2 N_Y_c_310_n 0.010499f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_114 N_B2_c_114_n N_Y_c_310_n 0.00150367f $X=1.405 $Y=1.845 $X2=0 $Y2=0
cc_115 N_B2_M1001_g N_Y_c_312_n 0.00130123f $X=1.055 $Y=0.485 $X2=0 $Y2=0
cc_116 N_B2_M1005_g N_A_210_535#_c_364_n 0.00604149f $X=1.405 $Y=2.885 $X2=0
+ $Y2=0
cc_117 N_B2_M1005_g N_A_210_535#_c_365_n 0.0193848f $X=1.405 $Y=2.885 $X2=0
+ $Y2=0
cc_118 B2 N_A_210_535#_c_365_n 0.00117525f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_119 N_B2_c_114_n N_A_210_535#_c_365_n 0.00107575f $X=1.405 $Y=1.845 $X2=0
+ $Y2=0
cc_120 B2 N_A_210_535#_c_366_n 0.0149683f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_121 N_B2_c_114_n N_A_210_535#_c_366_n 0.00544926f $X=1.405 $Y=1.845 $X2=0
+ $Y2=0
cc_122 N_B2_M1005_g N_A_296_535#_c_401_n 0.00161321f $X=1.405 $Y=2.885 $X2=0
+ $Y2=0
cc_123 N_B2_M1005_g N_VPWR_c_426_n 0.00585385f $X=1.405 $Y=2.885 $X2=0 $Y2=0
cc_124 N_B2_M1005_g N_VPWR_c_424_n 0.0110354f $X=1.405 $Y=2.885 $X2=0 $Y2=0
cc_125 N_B2_M1001_g N_VGND_c_463_n 0.00290284f $X=1.055 $Y=0.485 $X2=0 $Y2=0
cc_126 N_B2_M1001_g N_VGND_c_467_n 0.00406911f $X=1.055 $Y=0.485 $X2=0 $Y2=0
cc_127 N_B2_M1001_g N_VGND_c_470_n 0.00557894f $X=1.055 $Y=0.485 $X2=0 $Y2=0
cc_128 N_B1_c_164_n N_A1_M1000_g 0.0075632f $X=2.555 $Y=1.71 $X2=0 $Y2=0
cc_129 N_B1_M1002_g N_A1_M1004_g 0.025122f $X=1.415 $Y=0.485 $X2=0 $Y2=0
cc_130 N_B1_c_154_n N_A1_M1004_g 6.34754e-19 $X=1.505 $Y=1.275 $X2=0 $Y2=0
cc_131 N_B1_c_155_n N_A1_M1004_g 0.0212221f $X=1.505 $Y=1.275 $X2=0 $Y2=0
cc_132 B1 N_A1_c_219_n 0.00103776f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_133 N_B1_c_153_n N_A1_c_224_n 0.00161873f $X=1.585 $Y=1.75 $X2=0 $Y2=0
cc_134 N_B1_c_164_n N_A1_c_224_n 0.0153171f $X=2.555 $Y=1.71 $X2=0 $Y2=0
cc_135 N_B1_c_153_n A1 0.00790063f $X=1.585 $Y=1.75 $X2=0 $Y2=0
cc_136 N_B1_c_154_n A1 0.00794455f $X=1.505 $Y=1.275 $X2=0 $Y2=0
cc_137 N_B1_c_155_n A1 4.37045e-19 $X=1.505 $Y=1.275 $X2=0 $Y2=0
cc_138 B1 A1 0.00359273f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_139 N_B1_c_164_n A1 0.0175542f $X=2.555 $Y=1.71 $X2=0 $Y2=0
cc_140 N_B1_c_153_n N_A1_c_221_n 0.00728651f $X=1.585 $Y=1.75 $X2=0 $Y2=0
cc_141 N_B1_c_164_n N_A1_c_221_n 0.00391568f $X=2.555 $Y=1.71 $X2=0 $Y2=0
cc_142 N_B1_c_159_n N_A2_M1008_g 0.0450332f $X=2.975 $Y=2.045 $X2=0 $Y2=0
cc_143 N_B1_c_164_n N_A2_M1008_g 0.00418796f $X=2.555 $Y=1.71 $X2=0 $Y2=0
cc_144 B1 N_A2_c_265_n 0.00899438f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_145 N_B1_c_157_n N_A2_c_265_n 0.0149214f $X=2.975 $Y=1.54 $X2=0 $Y2=0
cc_146 N_B1_c_164_n N_A2_c_265_n 0.0055047f $X=2.555 $Y=1.71 $X2=0 $Y2=0
cc_147 N_B1_c_159_n N_A2_c_270_n 0.0149214f $X=2.975 $Y=2.045 $X2=0 $Y2=0
cc_148 B1 N_A2_c_270_n 0.00196947f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_149 N_B1_c_164_n N_A2_c_270_n 0.00573628f $X=2.555 $Y=1.71 $X2=0 $Y2=0
cc_150 B1 A2 0.0337092f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_151 N_B1_c_157_n A2 0.00863643f $X=2.975 $Y=1.54 $X2=0 $Y2=0
cc_152 N_B1_c_164_n A2 0.00136436f $X=2.555 $Y=1.71 $X2=0 $Y2=0
cc_153 B1 N_A2_c_267_n 0.00378101f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_154 N_B1_M1002_g Y 2.17641e-19 $X=1.415 $Y=0.485 $X2=0 $Y2=0
cc_155 N_B1_M1002_g N_Y_c_310_n 0.0111955f $X=1.415 $Y=0.485 $X2=0 $Y2=0
cc_156 N_B1_c_154_n N_Y_c_310_n 0.00837858f $X=1.505 $Y=1.275 $X2=0 $Y2=0
cc_157 N_B1_M1002_g N_Y_c_312_n 0.0109404f $X=1.415 $Y=0.485 $X2=0 $Y2=0
cc_158 N_B1_c_154_n N_Y_c_312_n 0.0153614f $X=1.505 $Y=1.275 $X2=0 $Y2=0
cc_159 N_B1_c_155_n N_Y_c_312_n 0.00455835f $X=1.505 $Y=1.275 $X2=0 $Y2=0
cc_160 N_B1_M1003_g N_A_210_535#_c_365_n 0.0163103f $X=2.885 $Y=2.885 $X2=0
+ $Y2=0
cc_161 N_B1_c_159_n N_A_210_535#_c_365_n 0.00524895f $X=2.975 $Y=2.045 $X2=0
+ $Y2=0
cc_162 N_B1_c_161_n N_A_210_535#_c_365_n 0.0135672f $X=1.67 $Y=1.857 $X2=0 $Y2=0
cc_163 B1 N_A_210_535#_c_365_n 0.01777f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_164 N_B1_c_164_n N_A_210_535#_c_365_n 0.0960688f $X=2.555 $Y=1.71 $X2=0 $Y2=0
cc_165 N_B1_M1003_g N_A_210_535#_c_367_n 0.0115115f $X=2.885 $Y=2.885 $X2=0
+ $Y2=0
cc_166 N_B1_M1003_g N_A_296_535#_c_400_n 0.00161321f $X=2.885 $Y=2.885 $X2=0
+ $Y2=0
cc_167 N_B1_M1003_g N_VPWR_c_427_n 0.00585385f $X=2.885 $Y=2.885 $X2=0 $Y2=0
cc_168 N_B1_M1003_g N_VPWR_c_424_n 0.0120125f $X=2.885 $Y=2.885 $X2=0 $Y2=0
cc_169 N_B1_M1002_g N_VGND_c_467_n 0.00401603f $X=1.415 $Y=0.485 $X2=0 $Y2=0
cc_170 N_B1_M1002_g N_VGND_c_470_n 0.00582181f $X=1.415 $Y=0.485 $X2=0 $Y2=0
cc_171 N_A1_M1004_g N_A2_c_264_n 0.0510569f $X=1.955 $Y=0.485 $X2=-0.19
+ $Y2=-0.245
cc_172 N_A1_c_219_n N_A2_c_265_n 0.00781511f $X=1.955 $Y=1.68 $X2=0 $Y2=0
cc_173 A1 N_A2_c_265_n 0.00618673f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A1_c_221_n N_A2_c_265_n 0.0195472f $X=2.045 $Y=1.36 $X2=0 $Y2=0
cc_175 N_A1_M1000_g N_A2_c_270_n 0.0333426f $X=1.835 $Y=2.885 $X2=0 $Y2=0
cc_176 N_A1_c_224_n N_A2_c_270_n 0.00218923f $X=1.955 $Y=1.755 $X2=0 $Y2=0
cc_177 N_A1_M1004_g A2 7.62088e-19 $X=1.955 $Y=0.485 $X2=0 $Y2=0
cc_178 N_A1_M1004_g N_A2_c_267_n 0.00802267f $X=1.955 $Y=0.485 $X2=0 $Y2=0
cc_179 N_A1_M1004_g Y 0.0168691f $X=1.955 $Y=0.485 $X2=0 $Y2=0
cc_180 N_A1_c_224_n Y 0.0022023f $X=1.955 $Y=1.755 $X2=0 $Y2=0
cc_181 A1 Y 0.0206676f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A1_c_221_n Y 0.00404133f $X=2.045 $Y=1.36 $X2=0 $Y2=0
cc_183 N_A1_M1004_g N_Y_c_312_n 0.00670525f $X=1.955 $Y=0.485 $X2=0 $Y2=0
cc_184 N_A1_c_224_n N_Y_c_312_n 9.52387e-19 $X=1.955 $Y=1.755 $X2=0 $Y2=0
cc_185 N_A1_M1000_g N_A_210_535#_c_365_n 0.0114097f $X=1.835 $Y=2.885 $X2=0
+ $Y2=0
cc_186 N_A1_c_224_n N_A_210_535#_c_365_n 5.95815e-19 $X=1.955 $Y=1.755 $X2=0
+ $Y2=0
cc_187 N_A1_M1000_g N_A_296_535#_c_404_n 2.1266e-19 $X=1.835 $Y=2.885 $X2=0
+ $Y2=0
cc_188 N_A1_M1000_g N_A_296_535#_c_400_n 0.0124817f $X=1.835 $Y=2.885 $X2=0
+ $Y2=0
cc_189 N_A1_M1000_g N_VPWR_c_425_n 0.00763401f $X=1.835 $Y=2.885 $X2=0 $Y2=0
cc_190 N_A1_M1000_g N_VPWR_c_426_n 0.00429465f $X=1.835 $Y=2.885 $X2=0 $Y2=0
cc_191 N_A1_M1000_g N_VPWR_c_424_n 0.00649311f $X=1.835 $Y=2.885 $X2=0 $Y2=0
cc_192 N_A1_M1004_g N_VGND_c_467_n 0.00406911f $X=1.955 $Y=0.485 $X2=0 $Y2=0
cc_193 N_A1_M1004_g N_VGND_c_470_n 0.00594019f $X=1.955 $Y=0.485 $X2=0 $Y2=0
cc_194 N_A2_c_264_n Y 0.00316694f $X=2.315 $Y=0.805 $X2=0 $Y2=0
cc_195 A2 Y 0.0122843f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_196 N_A2_c_267_n Y 0.00464681f $X=2.495 $Y=0.97 $X2=0 $Y2=0
cc_197 N_A2_M1008_g N_A_210_535#_c_365_n 0.0114097f $X=2.455 $Y=2.885 $X2=0
+ $Y2=0
cc_198 N_A2_c_270_n N_A_210_535#_c_365_n 2.59782e-19 $X=2.475 $Y=1.915 $X2=0
+ $Y2=0
cc_199 N_A2_M1008_g N_A_296_535#_c_400_n 0.0124817f $X=2.455 $Y=2.885 $X2=0
+ $Y2=0
cc_200 N_A2_M1008_g N_A_296_535#_c_407_n 2.1266e-19 $X=2.455 $Y=2.885 $X2=0
+ $Y2=0
cc_201 N_A2_M1008_g N_VPWR_c_425_n 0.00763401f $X=2.455 $Y=2.885 $X2=0 $Y2=0
cc_202 N_A2_M1008_g N_VPWR_c_427_n 0.00429465f $X=2.455 $Y=2.885 $X2=0 $Y2=0
cc_203 N_A2_M1008_g N_VPWR_c_424_n 0.00649311f $X=2.455 $Y=2.885 $X2=0 $Y2=0
cc_204 N_A2_c_264_n N_VGND_c_464_n 0.00468315f $X=2.315 $Y=0.805 $X2=0 $Y2=0
cc_205 A2 N_VGND_c_464_n 0.00862023f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_206 N_A2_c_267_n N_VGND_c_464_n 0.00618643f $X=2.495 $Y=0.97 $X2=0 $Y2=0
cc_207 N_A2_c_264_n N_VGND_c_467_n 0.00540927f $X=2.315 $Y=0.805 $X2=0 $Y2=0
cc_208 N_A2_c_264_n N_VGND_c_470_n 0.0110879f $X=2.315 $Y=0.805 $X2=0 $Y2=0
cc_209 A2 N_VGND_c_470_n 0.0216755f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_210 N_A2_c_267_n N_VGND_c_470_n 0.00346594f $X=2.495 $Y=0.97 $X2=0 $Y2=0
cc_211 N_Y_c_314_n N_A_210_535#_c_364_n 0.00128496f $X=0.76 $Y=2.82 $X2=0 $Y2=0
cc_212 N_Y_c_313_n N_VPWR_c_426_n 0.00769639f $X=0.27 $Y=2.82 $X2=0 $Y2=0
cc_213 N_Y_c_314_n N_VPWR_c_426_n 0.0249437f $X=0.76 $Y=2.82 $X2=0 $Y2=0
cc_214 N_Y_M1007_s N_VPWR_c_424_n 0.00344799f $X=0.635 $Y=2.675 $X2=0 $Y2=0
cc_215 N_Y_c_313_n N_VPWR_c_424_n 0.00628456f $X=0.27 $Y=2.82 $X2=0 $Y2=0
cc_216 N_Y_c_314_n N_VPWR_c_424_n 0.021514f $X=0.76 $Y=2.82 $X2=0 $Y2=0
cc_217 N_Y_c_310_n N_VGND_c_463_n 0.0145168f $X=1.465 $Y=0.877 $X2=0 $Y2=0
cc_218 N_Y_c_310_n N_VGND_c_465_n 0.00303106f $X=1.465 $Y=0.877 $X2=0 $Y2=0
cc_219 N_Y_c_311_n N_VGND_c_465_n 0.0154689f $X=0.41 $Y=0.55 $X2=0 $Y2=0
cc_220 Y N_VGND_c_467_n 0.00651177f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_221 N_Y_c_310_n N_VGND_c_467_n 0.00732988f $X=1.465 $Y=0.877 $X2=0 $Y2=0
cc_222 N_Y_c_312_n N_VGND_c_467_n 0.00868209f $X=1.63 $Y=0.57 $X2=0 $Y2=0
cc_223 Y N_VGND_c_470_n 0.0112495f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_224 N_Y_c_310_n N_VGND_c_470_n 0.0185424f $X=1.465 $Y=0.877 $X2=0 $Y2=0
cc_225 N_Y_c_311_n N_VGND_c_470_n 0.0149004f $X=0.41 $Y=0.55 $X2=0 $Y2=0
cc_226 N_Y_c_312_n N_VGND_c_470_n 0.0110115f $X=1.63 $Y=0.57 $X2=0 $Y2=0
cc_227 N_A_210_535#_c_364_n N_A_296_535#_c_404_n 5.51144e-19 $X=1.19 $Y=2.82
+ $X2=0 $Y2=0
cc_228 N_A_210_535#_c_365_n N_A_296_535#_c_400_n 0.0749918f $X=2.995 $Y=2.23
+ $X2=0 $Y2=0
cc_229 N_A_210_535#_c_367_n N_A_296_535#_c_400_n 0.0121358f $X=3.1 $Y=2.82 $X2=0
+ $Y2=0
cc_230 N_A_210_535#_c_364_n N_A_296_535#_c_401_n 0.0121358f $X=1.19 $Y=2.82
+ $X2=0 $Y2=0
cc_231 N_A_210_535#_c_365_n N_A_296_535#_c_401_n 0.0165841f $X=2.995 $Y=2.23
+ $X2=0 $Y2=0
cc_232 N_A_210_535#_c_367_n N_A_296_535#_c_407_n 5.51144e-19 $X=3.1 $Y=2.82
+ $X2=0 $Y2=0
cc_233 N_A_210_535#_c_364_n N_VPWR_c_426_n 0.00833885f $X=1.19 $Y=2.82 $X2=0
+ $Y2=0
cc_234 N_A_210_535#_c_367_n N_VPWR_c_427_n 0.00877924f $X=3.1 $Y=2.82 $X2=0
+ $Y2=0
cc_235 N_A_210_535#_M1007_d N_VPWR_c_424_n 0.00481916f $X=1.05 $Y=2.675 $X2=0
+ $Y2=0
cc_236 N_A_210_535#_M1003_d N_VPWR_c_424_n 0.0042053f $X=2.96 $Y=2.675 $X2=0
+ $Y2=0
cc_237 N_A_210_535#_c_364_n N_VPWR_c_424_n 0.00770513f $X=1.19 $Y=2.82 $X2=0
+ $Y2=0
cc_238 N_A_210_535#_c_367_n N_VPWR_c_424_n 0.00770513f $X=3.1 $Y=2.82 $X2=0
+ $Y2=0
cc_239 N_A_296_535#_c_400_n N_VPWR_c_425_n 0.0243929f $X=2.565 $Y=2.58 $X2=0
+ $Y2=0
cc_240 N_A_296_535#_c_404_n N_VPWR_c_426_n 0.0081737f $X=1.62 $Y=2.82 $X2=0
+ $Y2=0
cc_241 N_A_296_535#_c_400_n N_VPWR_c_426_n 0.00406811f $X=2.565 $Y=2.58 $X2=0
+ $Y2=0
cc_242 N_A_296_535#_c_400_n N_VPWR_c_427_n 0.00406811f $X=2.565 $Y=2.58 $X2=0
+ $Y2=0
cc_243 N_A_296_535#_c_407_n N_VPWR_c_427_n 0.0081737f $X=2.67 $Y=2.82 $X2=0
+ $Y2=0
cc_244 N_A_296_535#_M1005_d N_VPWR_c_424_n 0.00369956f $X=1.48 $Y=2.675 $X2=0
+ $Y2=0
cc_245 N_A_296_535#_M1008_d N_VPWR_c_424_n 0.00369956f $X=2.53 $Y=2.675 $X2=0
+ $Y2=0
cc_246 N_A_296_535#_c_404_n N_VPWR_c_424_n 0.00762225f $X=1.62 $Y=2.82 $X2=0
+ $Y2=0
cc_247 N_A_296_535#_c_400_n N_VPWR_c_424_n 0.0142305f $X=2.565 $Y=2.58 $X2=0
+ $Y2=0
cc_248 N_A_296_535#_c_407_n N_VPWR_c_424_n 0.00762225f $X=2.67 $Y=2.82 $X2=0
+ $Y2=0
