# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxbp_lp2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlxbp_lp2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.110000 0.835000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.705000 0.265000 7.270000 0.595000 ;
        RECT 7.100000 0.595000 7.270000 1.180000 ;
        RECT 7.100000 1.180000 7.555000 2.890000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.375000 2.025000 9.965000 2.890000 ;
        RECT 9.375000 2.890000 9.705000 3.065000 ;
        RECT 9.635000 0.440000 9.965000 2.025000 ;
    END
  END Q_N
  PIN GATE
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.175000 1.895000 1.845000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
        RECT 0.905000  0.085000  1.235000 0.645000 ;
        RECT 3.075000  0.085000  3.405000 0.635000 ;
        RECT 5.035000  0.085000  5.365000 0.715000 ;
        RECT 7.495000  0.085000  7.825000 0.725000 ;
        RECT 8.845000  0.085000  9.175000 0.900000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
        RECT 9.755000 -0.085000 9.925000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.080000 3.415000 ;
        RECT 0.755000 2.885000  1.085000 3.245000 ;
        RECT 3.030000 2.535000  3.360000 3.245000 ;
        RECT 5.490000 1.985000  5.820000 3.245000 ;
        RECT 7.755000 1.815000  8.085000 3.245000 ;
        RECT 8.845000 2.025000  9.175000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
        RECT 9.755000 3.245000 9.925000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.265000 0.445000 0.725000 ;
      RECT 0.115000 0.725000 0.285000 2.025000 ;
      RECT 0.115000 2.025000 0.475000 2.535000 ;
      RECT 0.115000 2.535000 2.280000 2.705000 ;
      RECT 0.115000 2.705000 0.475000 3.065000 ;
      RECT 1.215000 0.825000 2.055000 0.995000 ;
      RECT 1.215000 0.995000 1.385000 2.025000 ;
      RECT 1.215000 2.025000 1.695000 2.185000 ;
      RECT 1.215000 2.185000 3.100000 2.355000 ;
      RECT 1.725000 0.265000 2.055000 0.825000 ;
      RECT 1.950000 2.705000 2.280000 3.065000 ;
      RECT 2.285000 0.265000 2.615000 0.815000 ;
      RECT 2.285000 0.815000 4.505000 0.985000 ;
      RECT 2.285000 0.985000 2.455000 1.675000 ;
      RECT 2.285000 1.675000 2.750000 2.005000 ;
      RECT 2.770000 1.165000 3.100000 1.425000 ;
      RECT 2.770000 1.425000 4.155000 1.495000 ;
      RECT 2.930000 1.495000 4.155000 1.755000 ;
      RECT 2.930000 1.755000 3.100000 2.185000 ;
      RECT 3.740000 0.985000 4.505000 1.145000 ;
      RECT 3.975000 0.335000 4.855000 0.635000 ;
      RECT 4.130000 1.945000 4.460000 2.815000 ;
      RECT 4.130000 2.815000 5.310000 2.985000 ;
      RECT 4.335000 1.145000 4.505000 1.475000 ;
      RECT 4.335000 1.475000 4.960000 1.645000 ;
      RECT 4.640000 1.645000 4.960000 1.805000 ;
      RECT 4.685000 0.635000 4.855000 1.125000 ;
      RECT 4.685000 1.125000 6.350000 1.295000 ;
      RECT 5.140000 1.295000 5.310000 2.815000 ;
      RECT 5.490000 1.475000 5.810000 1.635000 ;
      RECT 5.490000 1.635000 6.760000 1.805000 ;
      RECT 6.020000 1.295000 6.350000 1.455000 ;
      RECT 6.145000 0.265000 6.475000 0.775000 ;
      RECT 6.145000 0.775000 6.760000 0.895000 ;
      RECT 6.145000 0.895000 6.920000 0.945000 ;
      RECT 6.275000 1.805000 6.605000 2.985000 ;
      RECT 6.590000 0.945000 6.920000 1.565000 ;
      RECT 6.590000 1.565000 6.760000 1.635000 ;
      RECT 8.285000 0.265000 8.615000 1.590000 ;
      RECT 8.285000 1.590000 9.195000 1.760000 ;
      RECT 8.285000 1.760000 8.615000 2.855000 ;
      RECT 8.865000 1.090000 9.195000 1.590000 ;
  END
END sky130_fd_sc_lp__dlxbp_lp2
