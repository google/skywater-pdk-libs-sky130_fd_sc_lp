* File: sky130_fd_sc_lp__mux2i_1.spice
* Created: Wed Sep  2 10:01:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2i_1.pex.spice"
.subckt sky130_fd_sc_lp__mux2i_1  VNB VPB A0 A1 S Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1005 N_Y_M1005_d N_A0_M1005_g N_A_29_73#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1386 AS=0.2394 PD=1.17 PS=2.25 NRD=0 NRS=2.856 M=1 R=5.6 SA=75000.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1000 N_A_212_73#_M1000_d N_A1_M1000_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2478 AS=0.1386 PD=2.27 PS=1.17 NRD=2.856 NRS=7.14 M=1 R=5.6 SA=75000.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A_304_237#_M1006_g N_A_29_73#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_A_212_73#_M1008_d N_S_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_S_M1003_g N_A_304_237#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1002_d N_A0_M1002_g N_A_52_367#_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2079 AS=0.3654 PD=1.59 PS=3.1 NRD=0 NRS=1.3002 M=1 R=8.4 SA=75000.2
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1007 A_236_367# N_A1_M1007_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=1.26 AD=0.2142
+ AS=0.2079 PD=1.6 PS=1.59 NRD=17.9664 NRS=7.8012 M=1 R=8.4 SA=75000.7
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A_304_237#_M1004_g A_236_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2961 AS=0.2142 PD=1.73 PS=1.6 NRD=23.443 NRS=17.9664 M=1 R=8.4 SA=75001.2
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1009 N_A_52_367#_M1009_d N_S_M1009_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2961 PD=3.05 PS=1.73 NRD=0 NRS=6.2449 M=1 R=8.4 SA=75001.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_S_M1001_g N_A_304_237#_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__mux2i_1.pxi.spice"
*
.ends
*
*
