* File: sky130_fd_sc_lp__nand2_4.spice
* Created: Fri Aug 28 10:47:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2_4.pex.spice"
.subckt sky130_fd_sc_lp__nand2_4  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1005 N_A_63_65#_M1005_d N_B_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1006 N_A_63_65#_M1006_d N_B_M1006_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1013 N_A_63_65#_M1006_d N_B_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1015 N_A_63_65#_M1015_d N_B_M1015_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1002 N_A_63_65#_M1015_d N_A_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1003 N_A_63_65#_M1003_d N_A_M1003_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1848 AS=0.1176 PD=1.28 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1009 N_A_63_65#_M1003_d N_A_M1009_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1848 AS=0.1176 PD=1.28 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1011 N_A_63_65#_M1011_d N_A_M1011_g N_Y_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.5229 AS=0.1764 PD=3.35 PS=1.54 NRD=9.3772 NRS=0 M=1 R=8.4 SA=75000.3
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1001_d N_B_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.2
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_B_M1010_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1010_d N_A_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.1
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2772 AS=0.1764 PD=1.7 PS=1.54 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1007_d N_A_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2772 AS=0.1764 PD=1.7 PS=1.54 NRD=14.8341 NRS=0 M=1 R=8.4 SA=75003.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_Y_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__nand2_4.pxi.spice"
*
.ends
*
*
