* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__invlp_2 A VGND VNB VPB VPWR Y
M1000 VPWR A a_116_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=8.064e+11p pd=6.32e+06u as=7.056e+11p ps=6.16e+06u
M1001 VGND A a_116_55# VNB nshort w=840000u l=150000u
+  ad=4.788e+11p pd=4.5e+06u as=5.292e+11p ps=4.62e+06u
M1002 a_116_55# A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1003 a_116_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_116_367# A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1005 Y A a_116_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_116_55# A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A a_116_55# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
