* File: sky130_fd_sc_lp__a21boi_lp.pxi.spice
* Created: Wed Sep  2 09:19:36 2020
* 
x_PM_SKY130_FD_SC_LP__A21BOI_LP%A2 N_A2_M1002_g N_A2_M1003_g A2 A2 N_A2_c_64_n
+ PM_SKY130_FD_SC_LP__A21BOI_LP%A2
x_PM_SKY130_FD_SC_LP__A21BOI_LP%A1 N_A1_M1005_g N_A1_M1004_g A1 A1 A1
+ N_A1_c_91_n PM_SKY130_FD_SC_LP__A21BOI_LP%A1
x_PM_SKY130_FD_SC_LP__A21BOI_LP%A_298_318# N_A_298_318#_M1008_d
+ N_A_298_318#_M1001_d N_A_298_318#_M1000_g N_A_298_318#_M1009_g
+ N_A_298_318#_c_128_n N_A_298_318#_c_129_n N_A_298_318#_M1006_g
+ N_A_298_318#_c_131_n N_A_298_318#_c_132_n N_A_298_318#_c_133_n
+ N_A_298_318#_c_134_n N_A_298_318#_c_140_n N_A_298_318#_c_141_n
+ N_A_298_318#_c_142_n N_A_298_318#_c_135_n N_A_298_318#_c_136_n
+ N_A_298_318#_c_144_n PM_SKY130_FD_SC_LP__A21BOI_LP%A_298_318#
x_PM_SKY130_FD_SC_LP__A21BOI_LP%B1_N N_B1_N_M1007_g N_B1_N_c_213_n
+ N_B1_N_M1001_g N_B1_N_M1008_g N_B1_N_c_210_n B1_N N_B1_N_c_211_n
+ N_B1_N_c_212_n PM_SKY130_FD_SC_LP__A21BOI_LP%B1_N
x_PM_SKY130_FD_SC_LP__A21BOI_LP%A_29_409# N_A_29_409#_M1002_s
+ N_A_29_409#_M1005_d N_A_29_409#_c_249_n N_A_29_409#_c_253_n
+ N_A_29_409#_c_250_n N_A_29_409#_c_251_n
+ PM_SKY130_FD_SC_LP__A21BOI_LP%A_29_409#
x_PM_SKY130_FD_SC_LP__A21BOI_LP%VPWR N_VPWR_M1002_d N_VPWR_M1001_s
+ N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n VPWR
+ N_VPWR_c_279_n N_VPWR_c_274_n N_VPWR_c_281_n
+ PM_SKY130_FD_SC_LP__A21BOI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A21BOI_LP%Y N_Y_M1004_d N_Y_M1000_d N_Y_c_312_n
+ N_Y_c_314_n N_Y_c_313_n Y PM_SKY130_FD_SC_LP__A21BOI_LP%Y
x_PM_SKY130_FD_SC_LP__A21BOI_LP%VGND N_VGND_M1003_s N_VGND_M1006_d
+ N_VGND_c_353_n N_VGND_c_354_n VGND N_VGND_c_355_n N_VGND_c_356_n
+ N_VGND_c_357_n N_VGND_c_358_n N_VGND_c_359_n N_VGND_c_360_n
+ PM_SKY130_FD_SC_LP__A21BOI_LP%VGND
cc_1 VNB N_A2_M1002_g 0.0451086f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.545
cc_2 VNB N_A2_M1003_g 0.0246732f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.445
cc_3 VNB A2 0.0239035f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_4 VNB N_A2_c_64_n 0.0428718f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.975
cc_5 VNB N_A1_M1004_g 0.0563593f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.445
cc_6 VNB A1 0.0202117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A1_c_91_n 0.0230488f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.975
cc_8 VNB N_A_298_318#_M1009_g 0.0283629f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.975
cc_9 VNB N_A_298_318#_c_128_n 0.00742322f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.975
cc_10 VNB N_A_298_318#_c_129_n 0.00691396f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=0.975
cc_11 VNB N_A_298_318#_M1006_g 0.0322096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_298_318#_c_131_n 0.0145448f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.975
cc_13 VNB N_A_298_318#_c_132_n 0.0108432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_298_318#_c_133_n 0.00770432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_298_318#_c_134_n 0.0233688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_298_318#_c_135_n 0.0476872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_298_318#_c_136_n 0.0145699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_N_M1007_g 0.0196902f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.545
cc_19 VNB N_B1_N_M1008_g 0.0227387f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.975
cc_20 VNB N_B1_N_c_210_n 0.0111102f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.975
cc_21 VNB N_B1_N_c_211_n 0.0757592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_N_c_212_n 0.00221721f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.975
cc_23 VNB N_VPWR_c_274_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_312_n 0.0118304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_313_n 0.00951199f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.975
cc_26 VNB N_VGND_c_353_n 0.0177827f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_27 VNB N_VGND_c_354_n 0.010217f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.975
cc_28 VNB N_VGND_c_355_n 0.0150312f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.975
cc_29 VNB N_VGND_c_356_n 0.03452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_357_n 0.0314166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_358_n 0.194307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_359_n 0.00511011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_360_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_A2_M1002_g 0.0510324f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.545
cc_35 VPB N_A1_M1005_g 0.0319685f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.545
cc_36 VPB A1 0.0147487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A1_c_91_n 0.0104568f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.975
cc_38 VPB N_A_298_318#_M1000_g 0.0418617f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_39 VPB N_A_298_318#_c_131_n 0.0211889f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.975
cc_40 VPB N_A_298_318#_c_133_n 2.58564e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_298_318#_c_140_n 0.0184714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_298_318#_c_141_n 0.010044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_298_318#_c_142_n 0.0493899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_298_318#_c_135_n 8.60962e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_298_318#_c_144_n 0.0134941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_B1_N_c_213_n 0.0118736f $X=-0.19 $Y=1.655 $X2=0.785 $Y2=0.445
cc_47 VPB N_B1_N_M1001_g 0.0388473f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_48 VPB N_B1_N_c_210_n 0.00560497f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.975
cc_49 VPB N_A_29_409#_c_249_n 0.0237458f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_50 VPB N_A_29_409#_c_250_n 0.0213282f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.975
cc_51 VPB N_A_29_409#_c_251_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=0.975
cc_52 VPB N_VPWR_c_275_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_276_n 0.0174132f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.975
cc_54 VPB N_VPWR_c_277_n 0.0370557f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=0.975
cc_55 VPB N_VPWR_c_278_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_279_n 0.0194022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_274_n 0.0688697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_281_n 0.0242092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_Y_c_314_n 0.0118354f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB Y 0.00808508f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=0.975
cc_61 N_A2_M1002_g N_A1_M1005_g 0.0497804f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_62 N_A2_M1002_g N_A1_M1004_g 0.0116723f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_63 N_A2_M1003_g N_A1_M1004_g 0.0549706f $X=0.785 $Y=0.445 $X2=0 $Y2=0
cc_64 A2 N_A1_M1004_g 0.00124679f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_65 N_A2_M1002_g A1 0.0290738f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_66 A2 A1 0.035364f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A2_c_64_n A1 0.00456523f $X=0.785 $Y=0.975 $X2=0 $Y2=0
cc_68 N_A2_M1002_g N_A1_c_91_n 0.0181444f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_69 N_A2_M1002_g N_A_29_409#_c_249_n 0.0106493f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_70 N_A2_M1002_g N_A_29_409#_c_253_n 0.0168628f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_71 N_A2_M1002_g N_A_29_409#_c_250_n 0.00788277f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_72 N_A2_M1002_g N_A_29_409#_c_251_n 8.67045e-19 $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_73 N_A2_M1002_g N_VPWR_c_275_n 0.0120252f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_74 N_A2_M1002_g N_VPWR_c_274_n 0.0080522f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_75 N_A2_M1002_g N_VPWR_c_281_n 0.00769046f $X=0.555 $Y=2.545 $X2=0 $Y2=0
cc_76 A2 N_Y_c_312_n 0.00919219f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_77 N_A2_M1003_g N_Y_c_313_n 0.00124735f $X=0.785 $Y=0.445 $X2=0 $Y2=0
cc_78 N_A2_M1003_g N_VGND_c_353_n 0.0131198f $X=0.785 $Y=0.445 $X2=0 $Y2=0
cc_79 A2 N_VGND_c_353_n 0.0228504f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_80 N_A2_c_64_n N_VGND_c_353_n 0.00728544f $X=0.785 $Y=0.975 $X2=0 $Y2=0
cc_81 N_A2_M1003_g N_VGND_c_356_n 0.00486043f $X=0.785 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A2_M1003_g N_VGND_c_358_n 0.0052289f $X=0.785 $Y=0.445 $X2=0 $Y2=0
cc_83 A2 N_VGND_c_358_n 0.0147313f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A1_M1005_g N_A_298_318#_M1000_g 0.0319694f $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_85 N_A1_M1004_g N_A_298_318#_M1009_g 0.031904f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_86 A1 N_A_298_318#_c_131_n 0.00140023f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_87 N_A1_c_91_n N_A_298_318#_c_131_n 0.0109234f $X=1.085 $Y=1.625 $X2=0 $Y2=0
cc_88 N_A1_M1004_g N_A_298_318#_c_134_n 0.00237083f $X=1.175 $Y=0.445 $X2=0
+ $Y2=0
cc_89 N_A1_M1005_g N_A_29_409#_c_253_n 0.0162684f $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_90 A1 N_A_29_409#_c_253_n 0.0200668f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A1_M1005_g N_A_29_409#_c_250_n 0.00214146f $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_92 A1 N_A_29_409#_c_250_n 0.0229033f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_93 N_A1_M1005_g N_A_29_409#_c_251_n 0.0117109f $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_94 A1 N_A_29_409#_c_251_n 0.00346429f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A1_M1005_g N_VPWR_c_275_n 0.0112475f $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_96 N_A1_M1005_g N_VPWR_c_277_n 0.00769046f $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_97 N_A1_M1005_g N_VPWR_c_274_n 0.00740844f $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_98 N_A1_M1005_g N_Y_c_312_n 8.50173e-19 $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_99 N_A1_M1004_g N_Y_c_312_n 0.0131483f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_100 A1 N_Y_c_312_n 0.0258104f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A1_c_91_n N_Y_c_312_n 8.8197e-19 $X=1.085 $Y=1.625 $X2=0 $Y2=0
cc_102 N_A1_M1005_g N_Y_c_314_n 9.25956e-19 $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_103 N_A1_M1004_g N_Y_c_313_n 0.00862747f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A1_M1005_g Y 0.00149861f $X=1.085 $Y=2.545 $X2=0 $Y2=0
cc_105 N_A1_M1004_g N_VGND_c_353_n 0.00227125f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A1_M1004_g N_VGND_c_356_n 0.00547815f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A1_M1004_g N_VGND_c_358_n 0.0100007f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_298_318#_M1006_g N_B1_N_M1007_g 0.0252009f $X=1.965 $Y=0.445 $X2=0
+ $Y2=0
cc_109 N_A_298_318#_c_136_n N_B1_N_M1007_g 0.00108861f $X=3.065 $Y=0.455 $X2=0
+ $Y2=0
cc_110 N_A_298_318#_c_131_n N_B1_N_c_213_n 0.0023267f $X=2.01 $Y=1.59 $X2=0
+ $Y2=0
cc_111 N_A_298_318#_c_140_n N_B1_N_c_213_n 0.0142977f $X=2.9 $Y=1.76 $X2=0 $Y2=0
cc_112 N_A_298_318#_c_142_n N_B1_N_c_213_n 9.07767e-19 $X=3.065 $Y=2.19 $X2=0
+ $Y2=0
cc_113 N_A_298_318#_c_144_n N_B1_N_c_213_n 0.00257949f $X=3.065 $Y=1.76 $X2=0
+ $Y2=0
cc_114 N_A_298_318#_c_142_n N_B1_N_M1001_g 0.0297969f $X=3.065 $Y=2.19 $X2=0
+ $Y2=0
cc_115 N_A_298_318#_c_135_n N_B1_N_M1008_g 0.0220224f $X=3.145 $Y=1.675 $X2=0
+ $Y2=0
cc_116 N_A_298_318#_c_136_n N_B1_N_M1008_g 0.00796321f $X=3.065 $Y=0.455 $X2=0
+ $Y2=0
cc_117 N_A_298_318#_c_133_n N_B1_N_c_210_n 0.0033235f $X=2.01 $Y=1.235 $X2=0
+ $Y2=0
cc_118 N_A_298_318#_c_134_n N_B1_N_c_210_n 0.0023267f $X=2.01 $Y=1.235 $X2=0
+ $Y2=0
cc_119 N_A_298_318#_c_140_n N_B1_N_c_210_n 0.00519665f $X=2.9 $Y=1.76 $X2=0
+ $Y2=0
cc_120 N_A_298_318#_c_135_n N_B1_N_c_210_n 0.00413475f $X=3.145 $Y=1.675 $X2=0
+ $Y2=0
cc_121 N_A_298_318#_c_132_n N_B1_N_c_211_n 0.0232701f $X=2.01 $Y=1.145 $X2=0
+ $Y2=0
cc_122 N_A_298_318#_c_133_n N_B1_N_c_211_n 0.00334982f $X=2.01 $Y=1.235 $X2=0
+ $Y2=0
cc_123 N_A_298_318#_c_140_n N_B1_N_c_211_n 0.00662933f $X=2.9 $Y=1.76 $X2=0
+ $Y2=0
cc_124 N_A_298_318#_c_144_n N_B1_N_c_211_n 7.00424e-19 $X=3.065 $Y=1.76 $X2=0
+ $Y2=0
cc_125 N_A_298_318#_M1006_g N_B1_N_c_212_n 0.00117133f $X=1.965 $Y=0.445 $X2=0
+ $Y2=0
cc_126 N_A_298_318#_c_132_n N_B1_N_c_212_n 4.32133e-19 $X=2.01 $Y=1.145 $X2=0
+ $Y2=0
cc_127 N_A_298_318#_c_133_n N_B1_N_c_212_n 0.0217144f $X=2.01 $Y=1.235 $X2=0
+ $Y2=0
cc_128 N_A_298_318#_c_140_n N_B1_N_c_212_n 0.0245014f $X=2.9 $Y=1.76 $X2=0 $Y2=0
cc_129 N_A_298_318#_c_135_n N_B1_N_c_212_n 0.0437465f $X=3.145 $Y=1.675 $X2=0
+ $Y2=0
cc_130 N_A_298_318#_M1000_g N_A_29_409#_c_251_n 0.0132025f $X=1.615 $Y=2.545
+ $X2=0 $Y2=0
cc_131 N_A_298_318#_M1000_g N_VPWR_c_275_n 7.76705e-19 $X=1.615 $Y=2.545 $X2=0
+ $Y2=0
cc_132 N_A_298_318#_M1000_g N_VPWR_c_276_n 0.00384804f $X=1.615 $Y=2.545 $X2=0
+ $Y2=0
cc_133 N_A_298_318#_c_140_n N_VPWR_c_276_n 0.0264017f $X=2.9 $Y=1.76 $X2=0 $Y2=0
cc_134 N_A_298_318#_c_142_n N_VPWR_c_276_n 0.0685263f $X=3.065 $Y=2.19 $X2=0
+ $Y2=0
cc_135 N_A_298_318#_M1000_g N_VPWR_c_277_n 0.00798857f $X=1.615 $Y=2.545 $X2=0
+ $Y2=0
cc_136 N_A_298_318#_c_142_n N_VPWR_c_279_n 0.0220321f $X=3.065 $Y=2.19 $X2=0
+ $Y2=0
cc_137 N_A_298_318#_M1000_g N_VPWR_c_274_n 0.0150632f $X=1.615 $Y=2.545 $X2=0
+ $Y2=0
cc_138 N_A_298_318#_c_142_n N_VPWR_c_274_n 0.0125808f $X=3.065 $Y=2.19 $X2=0
+ $Y2=0
cc_139 N_A_298_318#_M1000_g N_Y_c_312_n 0.00876749f $X=1.615 $Y=2.545 $X2=0
+ $Y2=0
cc_140 N_A_298_318#_M1009_g N_Y_c_312_n 0.0122183f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A_298_318#_c_129_n N_Y_c_312_n 0.00660182f $X=1.68 $Y=1.145 $X2=0 $Y2=0
cc_142 N_A_298_318#_M1006_g N_Y_c_312_n 0.00255593f $X=1.965 $Y=0.445 $X2=0
+ $Y2=0
cc_143 N_A_298_318#_c_131_n N_Y_c_312_n 0.0080292f $X=2.01 $Y=1.59 $X2=0 $Y2=0
cc_144 N_A_298_318#_c_133_n N_Y_c_312_n 0.0429424f $X=2.01 $Y=1.235 $X2=0 $Y2=0
cc_145 N_A_298_318#_c_134_n N_Y_c_312_n 0.00184074f $X=2.01 $Y=1.235 $X2=0 $Y2=0
cc_146 N_A_298_318#_c_141_n N_Y_c_312_n 0.00937694f $X=2.215 $Y=1.76 $X2=0 $Y2=0
cc_147 N_A_298_318#_M1000_g N_Y_c_314_n 0.0177664f $X=1.615 $Y=2.545 $X2=0 $Y2=0
cc_148 N_A_298_318#_M1009_g N_Y_c_313_n 0.0105938f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_298_318#_M1006_g N_Y_c_313_n 0.00132927f $X=1.965 $Y=0.445 $X2=0
+ $Y2=0
cc_150 N_A_298_318#_M1000_g Y 0.021842f $X=1.615 $Y=2.545 $X2=0 $Y2=0
cc_151 N_A_298_318#_c_129_n Y 3.04314e-19 $X=1.68 $Y=1.145 $X2=0 $Y2=0
cc_152 N_A_298_318#_c_131_n Y 0.00575062f $X=2.01 $Y=1.59 $X2=0 $Y2=0
cc_153 N_A_298_318#_c_141_n Y 0.012582f $X=2.215 $Y=1.76 $X2=0 $Y2=0
cc_154 N_A_298_318#_M1009_g N_VGND_c_354_n 0.00232946f $X=1.605 $Y=0.445 $X2=0
+ $Y2=0
cc_155 N_A_298_318#_M1006_g N_VGND_c_354_n 0.0122725f $X=1.965 $Y=0.445 $X2=0
+ $Y2=0
cc_156 N_A_298_318#_c_132_n N_VGND_c_354_n 9.4696e-19 $X=2.01 $Y=1.145 $X2=0
+ $Y2=0
cc_157 N_A_298_318#_c_133_n N_VGND_c_354_n 0.0094495f $X=2.01 $Y=1.235 $X2=0
+ $Y2=0
cc_158 N_A_298_318#_c_136_n N_VGND_c_354_n 0.0116648f $X=3.065 $Y=0.455 $X2=0
+ $Y2=0
cc_159 N_A_298_318#_M1009_g N_VGND_c_356_n 0.00382506f $X=1.605 $Y=0.445 $X2=0
+ $Y2=0
cc_160 N_A_298_318#_M1006_g N_VGND_c_356_n 0.00486043f $X=1.965 $Y=0.445 $X2=0
+ $Y2=0
cc_161 N_A_298_318#_c_136_n N_VGND_c_357_n 0.0194886f $X=3.065 $Y=0.455 $X2=0
+ $Y2=0
cc_162 N_A_298_318#_M1008_d N_VGND_c_358_n 0.00232985f $X=2.925 $Y=0.235 $X2=0
+ $Y2=0
cc_163 N_A_298_318#_M1009_g N_VGND_c_358_n 0.00578672f $X=1.605 $Y=0.445 $X2=0
+ $Y2=0
cc_164 N_A_298_318#_M1006_g N_VGND_c_358_n 0.00814425f $X=1.965 $Y=0.445 $X2=0
+ $Y2=0
cc_165 N_A_298_318#_c_136_n N_VGND_c_358_n 0.0124792f $X=3.065 $Y=0.455 $X2=0
+ $Y2=0
cc_166 N_B1_N_M1001_g N_VPWR_c_276_n 0.0249777f $X=2.8 $Y=2.545 $X2=0 $Y2=0
cc_167 N_B1_N_M1001_g N_VPWR_c_279_n 0.00769046f $X=2.8 $Y=2.545 $X2=0 $Y2=0
cc_168 N_B1_N_M1001_g N_VPWR_c_274_n 0.0140941f $X=2.8 $Y=2.545 $X2=0 $Y2=0
cc_169 N_B1_N_M1001_g N_Y_c_314_n 0.00192699f $X=2.8 $Y=2.545 $X2=0 $Y2=0
cc_170 N_B1_N_M1001_g Y 3.23659e-19 $X=2.8 $Y=2.545 $X2=0 $Y2=0
cc_171 N_B1_N_M1007_g N_VGND_c_354_n 0.00977713f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_172 N_B1_N_M1007_g N_VGND_c_357_n 0.00585385f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_173 N_B1_N_M1008_g N_VGND_c_357_n 0.00549284f $X=2.85 $Y=0.445 $X2=0 $Y2=0
cc_174 N_B1_N_M1007_g N_VGND_c_358_n 0.00977956f $X=2.49 $Y=0.445 $X2=0 $Y2=0
cc_175 N_B1_N_M1008_g N_VGND_c_358_n 0.00855583f $X=2.85 $Y=0.445 $X2=0 $Y2=0
cc_176 N_B1_N_c_212_n N_VGND_c_358_n 0.0113504f $X=2.69 $Y=0.99 $X2=0 $Y2=0
cc_177 N_A_29_409#_c_253_n N_VPWR_M1002_d 0.00490489f $X=1.185 $Y=2.415
+ $X2=-0.19 $Y2=1.655
cc_178 N_A_29_409#_c_249_n N_VPWR_c_275_n 0.0253679f $X=0.29 $Y=2.9 $X2=0 $Y2=0
cc_179 N_A_29_409#_c_253_n N_VPWR_c_275_n 0.0159108f $X=1.185 $Y=2.415 $X2=0
+ $Y2=0
cc_180 N_A_29_409#_c_251_n N_VPWR_c_275_n 0.0253679f $X=1.35 $Y=2.495 $X2=0
+ $Y2=0
cc_181 N_A_29_409#_c_251_n N_VPWR_c_277_n 0.021949f $X=1.35 $Y=2.495 $X2=0 $Y2=0
cc_182 N_A_29_409#_c_249_n N_VPWR_c_274_n 0.0125808f $X=0.29 $Y=2.9 $X2=0 $Y2=0
cc_183 N_A_29_409#_c_253_n N_VPWR_c_274_n 0.0121913f $X=1.185 $Y=2.415 $X2=0
+ $Y2=0
cc_184 N_A_29_409#_c_251_n N_VPWR_c_274_n 0.0124703f $X=1.35 $Y=2.495 $X2=0
+ $Y2=0
cc_185 N_A_29_409#_c_249_n N_VPWR_c_281_n 0.0220321f $X=0.29 $Y=2.9 $X2=0 $Y2=0
cc_186 N_A_29_409#_c_251_n N_Y_c_314_n 0.0536621f $X=1.35 $Y=2.495 $X2=0 $Y2=0
cc_187 N_A_29_409#_c_251_n Y 0.00157587f $X=1.35 $Y=2.495 $X2=0 $Y2=0
cc_188 N_VPWR_c_276_n N_Y_c_314_n 0.0488392f $X=2.535 $Y=2.19 $X2=0 $Y2=0
cc_189 N_VPWR_c_277_n N_Y_c_314_n 0.0233113f $X=2.37 $Y=3.33 $X2=0 $Y2=0
cc_190 N_VPWR_c_274_n N_Y_c_314_n 0.0132625f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_191 N_VPWR_c_276_n Y 0.00692915f $X=2.535 $Y=2.19 $X2=0 $Y2=0
cc_192 N_Y_c_313_n N_VGND_c_353_n 0.0118164f $X=1.58 $Y=0.47 $X2=0 $Y2=0
cc_193 N_Y_c_313_n N_VGND_c_354_n 0.0175876f $X=1.58 $Y=0.47 $X2=0 $Y2=0
cc_194 N_Y_c_313_n N_VGND_c_356_n 0.0241159f $X=1.58 $Y=0.47 $X2=0 $Y2=0
cc_195 N_Y_M1004_d N_VGND_c_358_n 0.00225465f $X=1.25 $Y=0.235 $X2=0 $Y2=0
cc_196 N_Y_c_313_n N_VGND_c_358_n 0.016053f $X=1.58 $Y=0.47 $X2=0 $Y2=0
cc_197 N_VGND_c_358_n A_172_47# 0.010279f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_198 N_VGND_c_358_n A_336_47# 0.00899413f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_199 N_VGND_c_358_n A_513_47# 0.00303139f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
