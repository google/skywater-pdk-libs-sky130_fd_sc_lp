# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__lsbuf_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__lsbuf_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  6.660000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.678000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 1.530000 1.245000 2.135000 ;
        RECT 1.075000 2.135000 1.245000 2.775000 ;
        RECT 1.075000 2.775000 1.910000 3.075000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.487600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.895000 3.585000 4.225000 6.405000 ;
    END
  END X
  PIN DESTPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 6.415000 4.800000 6.905000 ;
    END
  END DESTPWR
  PIN DESTVPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.090000 5.220000 0.390000 6.395000 ;
        RECT 4.410000 5.220000 4.710000 6.395000 ;
    END
  END DESTVPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.265000 0.390000 1.440000 ;
        RECT 4.410000 0.265000 4.710000 1.440000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 1.995000 3.415000 ;
      RECT 0.000000  6.575000 4.800000 6.745000 ;
      RECT 0.090000  1.890000 0.390000 3.245000 ;
      RECT 0.090000  3.415000 0.390000 4.770000 ;
      RECT 0.575000  0.085000 0.905000 1.175000 ;
      RECT 0.575000  2.305000 0.905000 3.245000 ;
      RECT 0.925000  3.585000 1.205000 4.650000 ;
      RECT 0.925000  4.650000 2.040000 4.820000 ;
      RECT 0.925000  4.820000 1.180000 5.435000 ;
      RECT 0.925000  5.435000 1.275000 6.405000 ;
      RECT 1.350000  4.990000 1.680000 5.265000 ;
      RECT 1.365000  0.265000 1.715000 1.360000 ;
      RECT 1.415000  1.360000 1.715000 2.435000 ;
      RECT 1.415000  2.435000 2.335000 2.605000 ;
      RECT 1.510000  5.265000 1.680000 5.355000 ;
      RECT 1.510000  5.355000 2.835000 5.525000 ;
      RECT 1.715000  3.415000 1.995000 4.480000 ;
      RECT 1.715000  5.695000 2.045000 6.575000 ;
      RECT 1.870000  4.820000 2.040000 5.010000 ;
      RECT 1.870000  5.010000 2.280000 5.185000 ;
      RECT 2.165000  2.605000 2.335000 4.310000 ;
      RECT 2.165000  4.310000 2.380000 4.480000 ;
      RECT 2.210000  4.480000 2.380000 4.610000 ;
      RECT 2.210000  4.610000 2.595000 4.740000 ;
      RECT 2.210000  4.740000 2.820000 4.840000 ;
      RECT 2.450000  4.840000 2.820000 4.990000 ;
      RECT 2.505000  3.245000 4.800000 3.415000 ;
      RECT 2.505000  3.585000 2.935000 4.140000 ;
      RECT 2.505000  5.525000 2.835000 6.395000 ;
      RECT 2.550000  4.140000 2.935000 4.400000 ;
      RECT 2.550000  4.400000 3.160000 4.440000 ;
      RECT 2.665000  5.160000 3.160000 5.330000 ;
      RECT 2.665000  5.330000 2.835000 5.355000 ;
      RECT 2.765000  4.440000 3.160000 4.570000 ;
      RECT 2.990000  4.570000 3.160000 5.160000 ;
      RECT 3.105000  3.415000 3.435000 4.230000 ;
      RECT 3.105000  5.500000 3.435000 6.575000 ;
      RECT 4.410000  1.890000 4.710000 3.245000 ;
      RECT 4.410000  3.415000 4.710000 4.770000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.155000  6.575000 0.325000 6.745000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 0.635000  6.575000 0.805000 6.745000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.115000  6.575000 1.285000 6.745000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 1.595000  6.575000 1.765000 6.745000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  6.575000 2.245000 6.745000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 2.555000  6.575000 2.725000 6.745000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.035000  6.575000 3.205000 6.745000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.515000  6.575000 3.685000 6.745000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 3.995000  6.575000 4.165000 6.745000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.475000  6.575000 4.645000 6.745000 ;
  END
END sky130_fd_sc_lp__lsbuf_lp
END LIBRARY
