* File: sky130_fd_sc_lp__o22a_4.spice
* Created: Wed Sep  2 10:20:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22a_4.pex.spice"
.subckt sky130_fd_sc_lp__o22a_4  VNB VPB B1 B2 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1005 N_X_M1005_d N_A_86_23#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1011 N_X_M1005_d N_A_86_23#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1015 N_X_M1015_d N_A_86_23#_M1015_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1016 N_X_M1015_d N_A_86_23#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_A_86_23#_M1010_d N_B1_M1010_g N_A_525_47#_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1006 N_A_86_23#_M1010_d N_B2_M1006_g N_A_525_47#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1021 N_A_86_23#_M1021_d N_B2_M1021_g N_A_525_47#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1019 N_A_86_23#_M1021_d N_B1_M1019_g N_A_525_47#_M1019_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6
+ SA=75001.5 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A1_M1000_g N_A_525_47#_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.1512 PD=1.19 PS=1.2 NRD=4.284 NRS=0 M=1 R=5.6 SA=75002
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1000_d N_A2_M1004_g N_A_525_47#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=5.712 NRS=0 M=1 R=5.6 SA=75002.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1020 N_VGND_M1020_d N_A2_M1020_g N_A_525_47#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1020_d N_A1_M1012_g N_A_525_47#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_86_23#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.1 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_86_23#_M1009_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1009_d N_A_86_23#_M1014_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_A_86_23#_M1022_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.22365 AS=0.1764 PD=1.615 PS=1.54 NRD=5.4569 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.9 A=0.189 P=2.82 MULT=1
MM1003 N_A_608_367#_M1003_d N_B1_M1003_g N_VPWR_M1022_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.22365 PD=1.54 PS=1.615 NRD=0 NRS=6.2449 M=1 R=8.4
+ SA=75002 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1008 N_A_608_367#_M1003_d N_B2_M1008_g N_A_86_23#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1018 N_A_608_367#_M1018_d N_B2_M1018_g N_A_86_23#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1023 N_A_608_367#_M1018_d N_B1_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2709 PD=1.54 PS=1.69 NRD=0 NRS=11.7215 M=1 R=8.4
+ SA=75003.3 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1023_s N_A1_M1007_g N_A_982_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2709 AS=0.1764 PD=1.69 PS=1.54 NRD=11.7215 NRS=0 M=1 R=8.4
+ SA=75003.9 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1001 N_A_86_23#_M1001_d N_A2_M1001_g N_A_982_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1017 N_A_86_23#_M1001_d N_A2_M1017_g N_A_982_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.7
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A1_M1013_g N_A_982_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.2415 P=17.93
*
.include "sky130_fd_sc_lp__o22a_4.pxi.spice"
*
.ends
*
*
