* File: sky130_fd_sc_lp__a2111oi_lp.pex.spice
* Created: Fri Aug 28 09:47:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111OI_LP%A1 3 7 11 12 13 15 22
r33 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.49
+ $Y=1.34 $X2=0.49 $Y2=1.34
r34 15 23 4.10594 $w=6.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.72 $Y=1.51
+ $X2=0.49 $Y2=1.51
r35 13 23 4.46298 $w=6.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.24 $Y=1.51
+ $X2=0.49 $Y2=1.51
r36 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.49 $Y=1.68
+ $X2=0.49 $Y2=1.34
r37 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.68
+ $X2=0.49 $Y2=1.845
r38 10 22 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.175
+ $X2=0.49 $Y2=1.34
r39 7 10 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.55 $Y=0.495
+ $X2=0.55 $Y2=1.175
r40 3 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.53 $Y=2.545 $X2=0.53
+ $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_LP%A2 3 7 9 11 18
r39 18 21 68.5216 $w=4.8e-07 $l=5.05e-07 $layer=POLY_cond $X=1.105 $Y=1.34
+ $X2=1.105 $Y2=1.845
r40 18 20 45.9721 $w=4.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.34
+ $X2=1.105 $Y2=1.175
r41 9 11 8.92596 $w=6.68e-07 $l=5e-07 $layer=LI1_cond $X=1.18 $Y=1.51 $X2=1.68
+ $Y2=1.51
r42 9 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.18 $Y=1.34
+ $X2=1.18 $Y2=1.34
r43 7 21 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.06 $Y=2.545 $X2=1.06
+ $Y2=1.845
r44 3 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.94 $Y=0.495
+ $X2=0.94 $Y2=1.175
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_LP%B1 1 3 4 5 6 8 10 11 12 13 15 16 18 19 21
+ 28
c62 11 0 1.62152e-19 $X=2.265 $Y=1.25
r63 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.43
+ $Y=1.34 $X2=2.43 $Y2=1.34
r64 21 29 3.7489 $w=6.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.64 $Y=1.51 $X2=2.43
+ $Y2=1.51
r65 19 29 4.82002 $w=6.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.16 $Y=1.51
+ $X2=2.43 $Y2=1.51
r66 18 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.43 $Y=1.68
+ $X2=2.43 $Y2=1.34
r67 17 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.43 $Y=1.325
+ $X2=2.43 $Y2=1.34
r68 13 18 47.383 $w=2.95e-07 $l=3.53129e-07 $layer=POLY_cond $X=2.57 $Y=1.97
+ $X2=2.43 $Y2=1.68
r69 13 15 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.57 $Y=1.97
+ $X2=2.57 $Y2=2.545
r70 11 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.265 $Y=1.25
+ $X2=2.43 $Y2=1.325
r71 11 12 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.265 $Y=1.25
+ $X2=1.805 $Y2=1.25
r72 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.73 $Y=1.175
+ $X2=1.805 $Y2=1.25
r73 9 16 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.73 $Y=0.93 $X2=1.73
+ $Y2=0.855
r74 9 10 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.73 $Y=0.93
+ $X2=1.73 $Y2=1.175
r75 6 16 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.73 $Y=0.78 $X2=1.73
+ $Y2=0.855
r76 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.73 $Y=0.78 $X2=1.73
+ $Y2=0.495
r77 4 16 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.655 $Y=0.855
+ $X2=1.73 $Y2=0.855
r78 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.655 $Y=0.855
+ $X2=1.445 $Y2=0.855
r79 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.37 $Y=0.78
+ $X2=1.445 $Y2=0.855
r80 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.37 $Y=0.78 $X2=1.37
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_LP%C1 1 3 4 5 8 10 12 16 17 18 19 20 21 22
+ 23 24 31
c66 31 0 1.26081e-19 $X=3.1 $Y=1.345
c67 16 0 2.58109e-19 $X=3.1 $Y=1.18
r68 23 24 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=2.405 $X2=3.1
+ $Y2=2.775
r69 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=2.035 $X2=3.1
+ $Y2=2.405
r70 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=1.665 $X2=3.1
+ $Y2=2.035
r71 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=1.295 $X2=3.1
+ $Y2=1.665
r72 20 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.1
+ $Y=1.345 $X2=3.1 $Y2=1.345
r73 17 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.1 $Y=1.685 $X2=3.1
+ $Y2=1.345
r74 17 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.685
+ $X2=3.1 $Y2=1.85
r75 16 31 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.18 $X2=3.1
+ $Y2=1.345
r76 13 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.05 $Y=0.88
+ $X2=3.05 $Y2=0.805
r77 13 16 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.05 $Y=0.88 $X2=3.05
+ $Y2=1.18
r78 10 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.05 $Y=0.73
+ $X2=3.05 $Y2=0.805
r79 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.05 $Y=0.73 $X2=3.05
+ $Y2=0.445
r80 8 18 172.675 $w=2.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.06 $Y=2.545
+ $X2=3.06 $Y2=1.85
r81 4 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.975 $Y=0.805
+ $X2=3.05 $Y2=0.805
r82 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.975 $Y=0.805
+ $X2=2.765 $Y2=0.805
r83 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.69 $Y=0.73
+ $X2=2.765 $Y2=0.805
r84 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.69 $Y=0.73 $X2=2.69
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_LP%D1 1 3 8 10 12 16 19 20 21 22 23 27
c48 22 0 9.59571e-20 $X=3.6 $Y=1.295
r49 22 23 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.66 $Y=1.295
+ $X2=3.66 $Y2=1.665
r50 22 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.67
+ $Y=1.34 $X2=3.67 $Y2=1.34
r51 20 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.67 $Y=1.68
+ $X2=3.67 $Y2=1.34
r52 20 21 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.68
+ $X2=3.67 $Y2=1.845
r53 19 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.175
+ $X2=3.67 $Y2=1.34
r54 15 16 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.58 $Y=0.805
+ $X2=3.84 $Y2=0.805
r55 13 15 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=3.48 $Y=0.805 $X2=3.58
+ $Y2=0.805
r56 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=0.73
+ $X2=3.84 $Y2=0.805
r57 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.84 $Y=0.73 $X2=3.84
+ $Y2=0.445
r58 8 21 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.63 $Y=2.545 $X2=3.63
+ $Y2=1.845
r59 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.58 $Y=0.88 $X2=3.58
+ $Y2=0.805
r60 4 19 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=3.58 $Y=0.88
+ $X2=3.58 $Y2=1.175
r61 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.48 $Y=0.73 $X2=3.48
+ $Y2=0.805
r62 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.48 $Y=0.73 $X2=3.48
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_LP%VPWR 1 2 7 9 13 17 19 26 27 33
r38 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r39 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r42 24 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r43 23 26 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=4.08 $Y2=3.33
r44 23 24 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 21 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=3.33
+ $X2=1.325 $Y2=3.33
r46 21 23 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.49 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 19 27 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 19 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 15 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=3.245
+ $X2=1.325 $Y2=3.33
r50 15 17 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.325 $Y=3.245
+ $X2=1.325 $Y2=2.54
r51 14 30 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=3.33
+ $X2=0.215 $Y2=3.33
r52 13 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=1.325 $Y2=3.33
r53 13 14 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=0.43 $Y2=3.33
r54 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.265 $Y=2.19
+ $X2=0.265 $Y2=2.9
r55 7 30 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.265 $Y=3.245
+ $X2=0.215 $Y2=3.33
r56 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.265 $Y=3.245
+ $X2=0.265 $Y2=2.9
r57 2 17 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=1.185
+ $Y=2.045 $X2=1.325 $Y2=2.54
r58 1 12 400 $w=1.7e-07 $l=9.17701e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.265 $Y2=2.9
r59 1 9 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.265 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_LP%A_131_409# 1 2 7 9 11 13 15
r34 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=2.195
+ $X2=2.305 $Y2=2.11
r35 13 15 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=2.305 $Y=2.195
+ $X2=2.305 $Y2=2.9
r36 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=2.11
+ $X2=0.795 $Y2=2.11
r37 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=2.11
+ $X2=2.305 $Y2=2.11
r38 11 12 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=2.14 $Y=2.11
+ $X2=0.96 $Y2=2.11
r39 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=2.195
+ $X2=0.795 $Y2=2.11
r40 7 9 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.795 $Y=2.195
+ $X2=0.795 $Y2=2.9
r41 2 20 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.16
+ $Y=2.045 $X2=2.305 $Y2=2.19
r42 2 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.16
+ $Y=2.045 $X2=2.305 $Y2=2.9
r43 1 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=2.045 $X2=0.795 $Y2=2.19
r44 1 9 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=2.045 $X2=0.795 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_LP%Y 1 2 3 4 15 17 18 21 23 25 29 33 35 37
+ 38 39 42
c89 23 0 1.26081e-19 $X=3.005 $Y=0.91
r90 39 42 2.30489 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=3.217 $Y=0.555
+ $X2=3.217 $Y2=0.47
r91 37 38 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.957 $Y=2.19
+ $X2=3.957 $Y2=2.025
r92 34 39 7.3214 $w=4.23e-07 $l=2.7e-07 $layer=LI1_cond $X=3.217 $Y=0.825
+ $X2=3.217 $Y2=0.555
r93 34 35 1.63918 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.217 $Y=0.825
+ $X2=3.217 $Y2=0.91
r94 31 38 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=4.1 $Y=0.995
+ $X2=4.1 $Y2=2.025
r95 27 37 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=3.957 $Y=2.252
+ $X2=3.957 $Y2=2.19
r96 27 29 17.0343 $w=4.53e-07 $l=6.48e-07 $layer=LI1_cond $X=3.957 $Y=2.252
+ $X2=3.957 $Y2=2.9
r97 26 35 10.2049 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=3.43 $Y=0.91
+ $X2=3.217 $Y2=0.91
r98 25 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=0.91
+ $X2=4.1 $Y2=0.995
r99 25 26 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.015 $Y=0.91
+ $X2=3.43 $Y2=0.91
r100 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=0.91
+ $X2=1.945 $Y2=0.91
r101 23 35 10.2049 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.005 $Y=0.91
+ $X2=3.217 $Y2=0.91
r102 23 24 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.005 $Y=0.91
+ $X2=2.11 $Y2=0.91
r103 19 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=0.825
+ $X2=1.945 $Y2=0.91
r104 19 21 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.945 $Y=0.825
+ $X2=1.945 $Y2=0.495
r105 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0.91
+ $X2=1.945 $Y2=0.91
r106 17 18 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=1.78 $Y=0.91
+ $X2=0.5 $Y2=0.91
r107 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.335 $Y=0.825
+ $X2=0.5 $Y2=0.91
r108 13 15 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.335 $Y=0.825
+ $X2=0.335 $Y2=0.495
r109 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=2.045 $X2=3.895 $Y2=2.19
r110 4 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=2.045 $X2=3.895 $Y2=2.9
r111 3 42 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.125
+ $Y=0.235 $X2=3.265 $Y2=0.47
r112 2 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.285 $X2=1.945 $Y2=0.495
r113 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.285 $X2=0.335 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_LP%VGND 1 2 3 12 16 18 20 23 24 25 27 36 44
+ 48
r61 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r62 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r63 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r64 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r65 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r66 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r67 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 36 47 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.105
+ $Y2=0
r69 36 41 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=3.6
+ $Y2=0
r70 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.155
+ $Y2=0
r71 32 34 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=2.16
+ $Y2=0
r72 30 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r73 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r74 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.155
+ $Y2=0
r75 27 29 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r76 25 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r77 25 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r78 25 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r79 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.64
+ $Y2=0
r80 23 34 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.16
+ $Y2=0
r81 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.475
+ $Y2=0
r82 18 47 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.105 $Y2=0
r83 18 20 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.055 $Y2=0.43
r84 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0
r85 14 16 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0.43
r86 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r87 10 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.455
r88 3 20 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.235 $X2=4.055 $Y2=0.43
r89 2 16 182 $w=1.7e-07 $l=2.51744e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.235 $X2=2.475 $Y2=0.43
r90 1 12 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.285 $X2=1.155 $Y2=0.455
.ends

