# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 1.515000 2.545000 1.840000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.130000 1.845000 10.475000 3.075000 ;
        RECT 10.205000 0.365000 10.475000 1.845000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.585000 2.475000 4.915000 2.635000 ;
        RECT 4.585000 2.635000 5.935000 2.805000 ;
        RECT 4.585000 2.805000 4.915000 2.985000 ;
        RECT 5.765000 2.805000 5.935000 2.905000 ;
        RECT 5.765000 2.905000 7.395000 3.075000 ;
        RECT 7.225000 1.555000 8.145000 1.885000 ;
        RECT 7.225000 1.885000 7.395000 2.905000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.450000 0.470000 2.130000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.245000 10.560000 3.415000 ;
      RECT 0.095000  0.620000  0.425000 1.100000 ;
      RECT 0.095000  1.100000  1.125000 1.280000 ;
      RECT 0.095000  2.300000  0.835000 2.470000 ;
      RECT 0.095000  2.470000  0.355000 2.970000 ;
      RECT 0.525000  2.640000  0.855000 3.245000 ;
      RECT 0.595000  0.085000  0.785000 0.930000 ;
      RECT 0.665000  1.280000  1.125000 1.770000 ;
      RECT 0.665000  1.770000  0.835000 2.300000 ;
      RECT 0.955000  0.280000  1.825000 0.450000 ;
      RECT 0.955000  0.450000  1.125000 1.100000 ;
      RECT 1.025000  1.940000  1.485000 2.135000 ;
      RECT 1.025000  2.135000  2.905000 2.335000 ;
      RECT 1.025000  2.335000  1.285000 2.960000 ;
      RECT 1.295000  0.620000  1.485000 1.940000 ;
      RECT 1.480000  2.505000  3.245000 2.675000 ;
      RECT 1.480000  2.675000  1.740000 3.035000 ;
      RECT 1.655000  0.450000  1.825000 1.175000 ;
      RECT 1.655000  1.175000  2.685000 1.345000 ;
      RECT 1.910000  2.845000  2.240000 3.245000 ;
      RECT 2.005000  0.085000  2.335000 1.005000 ;
      RECT 2.410000  2.675000  2.640000 3.035000 ;
      RECT 2.515000  0.470000  4.835000 0.525000 ;
      RECT 2.515000  0.525000  6.345000 0.640000 ;
      RECT 2.515000  0.640000  2.685000 1.175000 ;
      RECT 2.810000  2.845000  3.585000 3.075000 ;
      RECT 2.855000  0.810000  3.055000 1.785000 ;
      RECT 2.855000  1.785000  3.245000 1.955000 ;
      RECT 3.075000  1.955000  3.245000 2.505000 ;
      RECT 3.225000  0.640000  3.395000 1.605000 ;
      RECT 3.415000  2.445000  4.415000 2.615000 ;
      RECT 3.415000  2.615000  3.585000 2.845000 ;
      RECT 3.455000  1.875000  4.015000 2.180000 ;
      RECT 3.565000  0.810000  4.145000 0.930000 ;
      RECT 3.565000  0.930000  5.485000 1.140000 ;
      RECT 3.685000  1.310000  4.015000 1.875000 ;
      RECT 3.755000  2.795000  3.975000 3.245000 ;
      RECT 4.145000  2.615000  4.415000 3.035000 ;
      RECT 4.195000  2.125000  5.485000 2.295000 ;
      RECT 4.195000  2.295000  4.415000 2.445000 ;
      RECT 4.225000  1.355000  4.555000 1.495000 ;
      RECT 4.225000  1.495000  5.935000 1.665000 ;
      RECT 4.225000  1.665000  4.555000 1.955000 ;
      RECT 4.470000  0.640000  6.345000 0.705000 ;
      RECT 5.005000  0.085000  5.335000 0.355000 ;
      RECT 5.155000  1.140000  5.485000 1.315000 ;
      RECT 5.155000  1.845000  5.485000 2.125000 ;
      RECT 5.255000  2.975000  5.585000 3.245000 ;
      RECT 5.505000  0.255000  7.175000 0.525000 ;
      RECT 5.665000  0.875000  5.995000 1.065000 ;
      RECT 5.665000  1.065000  5.935000 1.495000 ;
      RECT 5.765000  1.665000  5.935000 2.265000 ;
      RECT 5.765000  2.265000  6.200000 2.465000 ;
      RECT 6.105000  1.755000  6.345000 2.085000 ;
      RECT 6.175000  0.705000  6.345000 1.755000 ;
      RECT 6.370000  2.265000  6.695000 2.735000 ;
      RECT 6.515000  0.695000  6.775000 1.195000 ;
      RECT 6.515000  1.195000  8.655000 1.365000 ;
      RECT 6.515000  1.365000  6.695000 2.265000 ;
      RECT 6.865000  1.545000  7.055000 2.215000 ;
      RECT 7.510000  0.085000  7.840000 1.025000 ;
      RECT 7.565000  2.095000  8.995000 2.265000 ;
      RECT 7.565000  2.265000  8.465000 2.425000 ;
      RECT 7.565000  2.630000  7.905000 3.245000 ;
      RECT 8.160000  2.425000  8.465000 2.960000 ;
      RECT 8.300000  0.695000  8.995000 1.025000 ;
      RECT 8.395000  1.365000  8.655000 1.865000 ;
      RECT 8.635000  2.630000  8.920000 3.245000 ;
      RECT 8.825000  1.025000  8.995000 2.095000 ;
      RECT 9.165000  0.430000  9.525000 1.335000 ;
      RECT 9.165000  1.335000 10.035000 1.665000 ;
      RECT 9.165000  1.665000  9.390000 2.490000 ;
      RECT 9.585000  1.845000  9.960000 3.245000 ;
      RECT 9.695000  0.085000 10.035000 1.165000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.950000  1.285000 2.120000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  1.950000  3.685000 2.120000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  1.950000  7.045000 2.120000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
    LAYER met1 ;
      RECT 1.055000 1.920000 1.345000 1.965000 ;
      RECT 1.055000 1.965000 7.105000 2.105000 ;
      RECT 1.055000 2.105000 1.345000 2.150000 ;
      RECT 3.455000 1.920000 3.745000 1.965000 ;
      RECT 3.455000 2.105000 3.745000 2.150000 ;
      RECT 6.815000 1.920000 7.105000 1.965000 ;
      RECT 6.815000 2.105000 7.105000 2.150000 ;
  END
END sky130_fd_sc_lp__dfrtp_1
