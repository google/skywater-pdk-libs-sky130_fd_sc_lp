# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__and4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__and4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.690000 1.425000 6.140000 1.760000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.470000 0.855000 2.120000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.480000 1.210000 3.900000 1.790000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 1.210000 3.310000 1.795000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 1.075000 2.515000 1.245000 ;
        RECT 1.115000 1.245000 1.295000 1.815000 ;
        RECT 1.115000 1.815000 2.505000 2.145000 ;
        RECT 1.425000 0.255000 1.655000 1.075000 ;
        RECT 2.325000 0.255000 2.515000 1.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.205000  0.700000 0.455000 2.465000 ;
      RECT 0.205000  2.465000 4.960000 2.645000 ;
      RECT 0.965000  2.815000 1.295000 3.245000 ;
      RECT 1.025000  0.085000 1.255000 0.905000 ;
      RECT 1.465000  1.415000 2.855000 1.645000 ;
      RECT 1.825000  0.085000 2.155000 0.905000 ;
      RECT 1.825000  2.815000 2.155000 3.245000 ;
      RECT 2.685000  0.870000 5.100000 0.905000 ;
      RECT 2.685000  0.905000 4.405000 1.040000 ;
      RECT 2.685000  1.040000 2.855000 1.415000 ;
      RECT 2.685000  1.645000 2.855000 1.965000 ;
      RECT 2.685000  1.965000 4.610000 2.295000 ;
      RECT 2.765000  2.815000 3.095000 3.245000 ;
      RECT 2.790000  0.085000 3.120000 0.700000 ;
      RECT 3.460000  0.255000 5.100000 0.870000 ;
      RECT 3.750000  2.815000 4.080000 3.245000 ;
      RECT 4.105000  1.345000 4.445000 1.615000 ;
      RECT 4.105000  1.615000 4.960000 1.785000 ;
      RECT 4.645000  1.075000 6.145000 1.245000 ;
      RECT 4.645000  1.245000 4.975000 1.445000 ;
      RECT 4.770000  2.815000 5.100000 3.245000 ;
      RECT 4.790000  1.785000 4.960000 2.465000 ;
      RECT 5.340000  1.245000 5.510000 1.930000 ;
      RECT 5.340000  1.930000 5.640000 2.260000 ;
      RECT 5.385000  0.085000 5.715000 0.905000 ;
      RECT 5.885000  0.695000 6.145000 1.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__and4bb_4
END LIBRARY
