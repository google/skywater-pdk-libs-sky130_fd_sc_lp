* File: sky130_fd_sc_lp__clkbuf_16.spice
* Created: Wed Sep  2 09:38:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkbuf_16.pex.spice"
.subckt sky130_fd_sc_lp__clkbuf_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1011 N_A_116_47#_M1011_d N_A_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1239 PD=0.7 PS=1.43 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75008.8
+ A=0.063 P=1.14 MULT=1
MM1026 N_A_116_47#_M1011_d N_A_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75008.3
+ A=0.063 P=1.14 MULT=1
MM1029 N_A_116_47#_M1029_d N_A_M1029_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75007.9
+ A=0.063 P=1.14 MULT=1
MM1030 N_A_116_47#_M1029_d N_A_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1407 PD=0.7 PS=1.09 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75007.5
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1030_s N_A_116_47#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1407 AS=0.0588 PD=1.09 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.3 SB=75006.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_116_47#_M1003_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.8 SB=75006.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1003_d N_A_116_47#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.2 SB=75005.8
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_116_47#_M1006_g N_X_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.6 SB=75005.3
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1006_d N_A_116_47#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.1 SB=75004.9
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_116_47#_M1008_g N_X_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.5 SB=75004.5
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1008_d N_A_116_47#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.9 SB=75004.1
+ A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_116_47#_M1012_g N_X_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.3 SB=75003.6
+ A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1012_d N_A_116_47#_M1018_g N_X_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.8 SB=75003.2
+ A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_116_47#_M1020_g N_X_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.2 SB=75002.8
+ A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1020_d N_A_116_47#_M1023_g N_X_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006.6 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_116_47#_M1024_g N_X_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.1 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1024_d N_A_116_47#_M1027_g N_X_M1027_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.5 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_A_116_47#_M1031_g N_X_M1027_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.9 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1031_d N_A_116_47#_M1033_g N_X_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75008.4 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_A_116_47#_M1036_g N_X_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75008.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_116_47#_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3717 AS=0.1764 PD=3.11 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75008.8 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1021_d N_A_M1021_g N_A_116_47#_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75008.3 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1021_d N_A_M1025_g N_A_116_47#_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75007.9 A=0.189 P=2.82 MULT=1
MM1035 N_VPWR_M1035_d N_A_M1035_g N_A_116_47#_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4221 AS=0.1764 PD=1.93 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75007.5 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1035_d N_A_116_47#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4221 AS=0.1764 PD=1.93 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75006.6 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A_116_47#_M1002_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75006.2 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1002_d N_A_116_47#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75005.8 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A_116_47#_M1013_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75005.3 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1013_d N_A_116_47#_M1014_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1015 N_VPWR_M1015_d N_A_116_47#_M1015_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1015_d N_A_116_47#_M1016_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.9
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_A_116_47#_M1017_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.3
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1017_d N_A_116_47#_M1019_g N_X_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.8
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_A_116_47#_M1022_g N_X_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.2
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1028 N_VPWR_M1022_d N_A_116_47#_M1028_g N_X_M1028_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.6
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1032 N_VPWR_M1032_d N_A_116_47#_M1032_g N_X_M1028_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.1
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1034 N_VPWR_M1032_d N_A_116_47#_M1034_g N_X_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.5
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1037_d N_A_116_47#_M1037_g N_X_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.9
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1038 N_VPWR_M1037_d N_A_116_47#_M1038_g N_X_M1038_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1039 N_VPWR_M1039_d N_A_116_47#_M1039_g N_X_M1038_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75008.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=18.6127 P=23.69
*
.include "sky130_fd_sc_lp__clkbuf_16.pxi.spice"
*
.ends
*
*
