* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_2 A0 A1 S VGND VNB VPB VPWR X
X0 VGND S a_284_279# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_319_48# A0 a_86_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR S a_284_279# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_508_449# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_86_21# A0 a_508_449# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_350_449# A1 a_86_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_86_21# A1 a_499_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_86_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR a_86_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND a_284_279# a_319_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR a_284_279# a_350_449# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 X a_86_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 X a_86_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_499_48# S VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
