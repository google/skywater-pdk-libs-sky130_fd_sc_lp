* File: sky130_fd_sc_lp__o31ai_1.spice
* Created: Wed Sep  2 10:25:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o31ai_1.pex.spice"
.subckt sky130_fd_sc_lp__o31ai_1  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_A_110_47#_M1004_d N_A1_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_110_47#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1003 N_A_110_47#_M1003_d N_A3_M1003_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.2604 PD=1.19 PS=1.46 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_110_47#_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.147 PD=2.21 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1007 A_110_367# N_A1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1006 A_182_367# N_A2_M1006_g A_110_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_A3_M1002_g A_182_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.40005
+ AS=0.2457 PD=1.895 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4 SA=75001.1 SB=75001
+ A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.40005 PD=3.05 PS=1.895 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__o31ai_1.pxi.spice"
*
.ends
*
*
