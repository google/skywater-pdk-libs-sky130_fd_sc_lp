* File: sky130_fd_sc_lp__lsbuf_lp.pex.spice
* Created: Fri Aug 28 10:42:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%VGND 1 2 3 26 42 46 52 64 65 71 83 87
c95 46 0 1.8723e-19 $X=1.88 $Y=3.715
r96 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r97 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r98 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r99 78 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r101 75 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r102 75 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r104 72 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=3.33
+ $X2=3.27 $Y2=3.33
r105 72 74 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.435 $Y=3.33
+ $X2=4.08 $Y2=3.33
r106 71 86 3.44808 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.41 $Y=3.33
+ $X2=4.605 $Y2=3.33
r107 71 74 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.41 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 70 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 67 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r111 67 69 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 65 84 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r113 65 70 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r114 64 69 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.68 $Y2=3.33
r115 59 86 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=4.56 $Y=3.415
+ $X2=4.605 $Y2=3.33
r116 54 86 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=4.56 $Y=3.245
+ $X2=4.605 $Y2=3.33
r117 50 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=3.415
+ $X2=3.27 $Y2=3.33
r118 50 52 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.27 $Y=3.415
+ $X2=3.27 $Y2=3.715
r119 44 64 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.855 $Y=3.415
+ $X2=1.715 $Y2=3.33
r120 44 46 12.3476 $w=2.78e-07 $l=3e-07 $layer=LI1_cond $X=1.855 $Y=3.415
+ $X2=1.855 $Y2=3.715
r121 40 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=3.33
r122 40 42 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=2.44
r123 39 77 3.44808 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r124 38 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r125 38 39 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.39 $Y2=3.33
r126 33 77 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.24 $Y=3.415
+ $X2=0.195 $Y2=3.33
r127 28 77 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.195 $Y2=3.33
r128 26 59 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=4.56 $Y=3.855
+ $X2=4.56 $Y2=3.415
r129 26 54 32.8446 $w=2.98e-07 $l=8.55e-07 $layer=LI1_cond $X=4.56 $Y=2.39
+ $X2=4.56 $Y2=3.245
r130 26 33 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=0.24 $Y=3.855
+ $X2=0.24 $Y2=3.415
r131 26 28 32.8446 $w=2.98e-07 $l=8.55e-07 $layer=LI1_cond $X=0.24 $Y=2.39
+ $X2=0.24 $Y2=3.245
r132 3 52 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.125
+ $Y=3.59 $X2=3.27 $Y2=3.715
r133 2 46 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.74
+ $Y=3.59 $X2=1.88 $Y2=3.715
r134 1 42 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=2.23 $X2=0.74 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%VPB 7 9 10 11 12 13 14
r19 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=4.56 $Y=0.925
+ $X2=4.56 $Y2=1.295
r20 12 13 15.3659 $w=2.98e-07 $l=4e-07 $layer=LI1_cond $X=4.56 $Y=0.525 $X2=4.56
+ $Y2=0.925
r21 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.295
r22 9 10 15.3659 $w=2.98e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=0.525 $X2=0.24
+ $Y2=0.925
r23 7 12 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=4.475 $Y=0.32 $X2=4.56 $Y2=0.525
r24 7 9 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0.155
+ $Y=0.32 $X2=0.24 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%DESTVPB 7 9 10 11 12 13 14
r44 13 14 15.558 $w=2.98e-07 $l=4.05e-07 $layer=LI1_cond $X=4.56 $Y=5.7 $X2=4.56
+ $Y2=6.105
r45 12 13 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=4.56 $Y=5.365
+ $X2=4.56 $Y2=5.7
r46 10 11 15.558 $w=2.98e-07 $l=4.05e-07 $layer=LI1_cond $X=0.24 $Y=5.7 $X2=0.24
+ $Y2=6.105
r47 9 10 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=5.365
+ $X2=0.24 $Y2=5.7
r48 7 13 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=4.475 $Y=5.495 $X2=4.56 $Y2=5.7
r49 7 10 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=0.155 $Y=5.495 $X2=0.24 $Y2=5.7
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%A_246_987# 1 2 9 13 15 17 19 24 26 28 30 34
+ 44
c83 15 0 1.01247e-19 $X=2.505 $Y=5.44
r84 34 36 11.5428 $w=4.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.72 $Y=3.715
+ $X2=2.72 $Y2=4.14
r85 31 44 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.515 $Y=5.1
+ $X2=1.665 $Y2=5.1
r86 31 41 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.515 $Y=5.1
+ $X2=1.305 $Y2=5.1
r87 30 32 16.4603 $w=2.52e-07 $l=3.4e-07 $layer=LI1_cond $X=1.515 $Y=5.1
+ $X2=1.515 $Y2=5.44
r88 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.515
+ $Y=5.1 $X2=1.515 $Y2=5.1
r89 27 28 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.075 $Y=4.57
+ $X2=3.075 $Y2=5.16
r90 26 36 4.04103 $w=3.83e-07 $l=1.35e-07 $layer=LI1_cond $X=2.742 $Y=4.275
+ $X2=2.742 $Y2=4.14
r91 24 27 32.7629 $w=1.24e-07 $l=3.73087e-07 $layer=LI1_cond $X=2.742 $Y=4.4
+ $X2=3.075 $Y2=4.485
r92 24 26 3.7417 $w=3.83e-07 $l=1.25e-07 $layer=LI1_cond $X=2.742 $Y=4.4
+ $X2=2.742 $Y2=4.275
r93 19 21 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.67 $Y=5.55
+ $X2=2.67 $Y2=6.3
r94 17 28 22.4591 $w=2.2e-07 $l=4.87581e-07 $layer=LI1_cond $X=2.67 $Y=5.342
+ $X2=3.075 $Y2=5.16
r95 17 19 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.67 $Y=5.525
+ $X2=2.67 $Y2=5.55
r96 16 32 3.04159 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=5.44
+ $X2=1.515 $Y2=5.44
r97 15 17 9.81194 $w=2.2e-07 $l=2.08315e-07 $layer=LI1_cond $X=2.505 $Y=5.44
+ $X2=2.67 $Y2=5.342
r98 15 16 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.505 $Y=5.44
+ $X2=1.68 $Y2=5.44
r99 11 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=5.265
+ $X2=1.665 $Y2=5.1
r100 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.665 $Y=5.265
+ $X2=1.665 $Y2=5.925
r101 7 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.305 $Y=5.265
+ $X2=1.305 $Y2=5.1
r102 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.305 $Y=5.265
+ $X2=1.305 $Y2=5.925
r103 2 21 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=5.425 $X2=2.67 $Y2=6.3
r104 2 19 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=5.425 $X2=2.67 $Y2=5.55
r105 1 34 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=3.59 $X2=2.67 $Y2=3.715
r106 1 26 182 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=3.59 $X2=2.67 $Y2=4.275
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%A 3 5 7 10 14 19 22 25 26 28 31 38 42 48
r64 41 42 51.7485 $w=3.26e-07 $l=3.5e-07 $layer=POLY_cond $X=1.315 $Y=2.925
+ $X2=1.665 $Y2=2.925
r65 40 41 1.47853 $w=3.26e-07 $l=1e-08 $layer=POLY_cond $X=1.305 $Y=2.925
+ $X2=1.315 $Y2=2.925
r66 37 48 1.38389 $w=6.03e-07 $l=7e-08 $layer=LI1_cond $X=1.09 $Y=1.832 $X2=1.16
+ $Y2=1.832
r67 36 38 38.1866 $w=3.4e-07 $l=2.25e-07 $layer=POLY_cond $X=1.09 $Y=1.96
+ $X2=1.315 $Y2=1.96
r68 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.09
+ $Y=1.955 $X2=1.09 $Y2=1.955
r69 33 36 22.912 $w=3.4e-07 $l=1.35e-07 $layer=POLY_cond $X=0.955 $Y=1.96
+ $X2=1.09 $Y2=1.96
r70 31 37 7.21601 $w=6.03e-07 $l=3.65e-07 $layer=LI1_cond $X=0.725 $Y=1.832
+ $X2=1.09 $Y2=1.832
r71 29 42 11.8282 $w=3.26e-07 $l=8e-08 $layer=POLY_cond $X=1.745 $Y=2.925
+ $X2=1.665 $Y2=2.925
r72 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.745
+ $Y=2.925 $X2=1.745 $Y2=2.925
r73 26 28 19.2074 $w=2.98e-07 $l=5e-07 $layer=LI1_cond $X=1.245 $Y=2.925
+ $X2=1.745 $Y2=2.925
r74 25 26 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.16 $Y=2.775
+ $X2=1.245 $Y2=2.925
r75 24 48 8.37032 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=1.16 $Y=2.135
+ $X2=1.16 $Y2=1.832
r76 24 25 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.16 $Y=2.135
+ $X2=1.16 $Y2=2.775
r77 20 42 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=3.09
+ $X2=1.665 $Y2=2.925
r78 20 22 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=1.665 $Y=3.09
+ $X2=1.665 $Y2=4.01
r79 17 41 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.315 $Y=2.76
+ $X2=1.315 $Y2=2.925
r80 17 19 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.315 $Y=2.76
+ $X2=1.315 $Y2=2.44
r81 16 38 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.315 $Y=2.13
+ $X2=1.315 $Y2=1.96
r82 16 19 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.315 $Y=2.13
+ $X2=1.315 $Y2=2.44
r83 12 38 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.315 $Y=1.79
+ $X2=1.315 $Y2=1.96
r84 12 14 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=1.315 $Y=1.79
+ $X2=1.315 $Y2=0.735
r85 8 40 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.305 $Y=3.09
+ $X2=1.305 $Y2=2.925
r86 8 10 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=1.305 $Y=3.09
+ $X2=1.305 $Y2=4.01
r87 5 33 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.955 $Y=2.13
+ $X2=0.955 $Y2=1.96
r88 5 7 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.955 $Y=2.13
+ $X2=0.955 $Y2=2.44
r89 1 33 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.955 $Y=1.79
+ $X2=0.955 $Y2=1.96
r90 1 3 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=0.955 $Y=1.79
+ $X2=0.955 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%A_278_47# 1 2 7 9 10 11 12 14 17 22 23 26
+ 27 33
c67 33 0 1.01247e-19 $X=2.6 $Y=4.615
c68 26 0 2.4388e-19 $X=2.25 $Y=4.31
c69 10 0 6.03389e-20 $X=2.38 $Y=4.615
r70 32 33 31.8302 $w=3.18e-07 $l=2.1e-07 $layer=POLY_cond $X=2.6 $Y=4.825
+ $X2=2.6 $Y2=4.615
r71 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.655
+ $Y=4.825 $X2=2.655 $Y2=4.825
r72 26 31 21.8592 $w=3.31e-07 $l=6.24384e-07 $layer=LI1_cond $X=2.25 $Y=4.31
+ $X2=2.492 $Y2=4.825
r73 25 26 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=2.25 $Y=2.605
+ $X2=2.25 $Y2=4.31
r74 24 29 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.715 $Y=2.52
+ $X2=1.565 $Y2=2.52
r75 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.165 $Y=2.52
+ $X2=2.25 $Y2=2.605
r76 23 24 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.165 $Y=2.52
+ $X2=1.715 $Y2=2.52
r77 22 29 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=2.435
+ $X2=1.565 $Y2=2.52
r78 22 27 41.2959 $w=2.98e-07 $l=1.075e-06 $layer=LI1_cond $X=1.565 $Y=2.435
+ $X2=1.565 $Y2=1.36
r79 17 20 23.3781 $w=3.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.54 $Y=0.38
+ $X2=1.54 $Y2=1.09
r80 15 27 6.02978 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=1.54 $Y=1.185
+ $X2=1.54 $Y2=1.36
r81 15 20 3.12806 $w=3.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.54 $Y=1.185
+ $X2=1.54 $Y2=1.09
r82 12 33 24.9017 $w=3.18e-07 $l=1.78606e-07 $layer=POLY_cond $X=2.455 $Y=4.54
+ $X2=2.6 $Y2=4.615
r83 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.455 $Y=4.54
+ $X2=2.455 $Y2=4.01
r84 10 33 20.3436 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.38 $Y=4.615
+ $X2=2.6 $Y2=4.615
r85 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.38 $Y=4.615
+ $X2=2.17 $Y2=4.615
r86 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.095 $Y=4.54
+ $X2=2.17 $Y2=4.615
r87 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.095 $Y=4.54
+ $X2=2.095 $Y2=4.01
r88 2 20 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.39
+ $Y=0.235 $X2=1.53 $Y2=1.09
r89 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.39
+ $Y=0.235 $X2=1.53 $Y2=0.38
r90 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.39
+ $Y=2.23 $X2=1.53 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%A_193_718# 1 2 7 9 10 12 13 14 15 19 23 25
+ 29 33 35 39 40 43 49 51 54 55 57 58 62
c116 62 0 6.03389e-20 $X=2.115 $Y=5.1
c117 35 0 6.27731e-20 $X=3.105 $Y=5.01
c118 14 0 1.8723e-19 $X=2.53 $Y=5.275
c119 13 0 1.81107e-19 $X=3.03 $Y=5.275
r120 63 65 3.32414 $w=2.9e-07 $l=2e-08 $layer=POLY_cond $X=2.115 $Y=5.142
+ $X2=2.095 $Y2=5.142
r121 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=5.1 $X2=2.115 $Y2=5.1
r122 57 58 5.31505 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=1.1 $Y=5.57
+ $X2=1.1 $Y2=5.435
r123 54 62 10.1403 $w=1.73e-07 $l=1.6e-07 $layer=LI1_cond $X=1.955 $Y=5.097
+ $X2=2.115 $Y2=5.097
r124 53 54 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.955 $Y=4.82
+ $X2=1.955 $Y2=5.01
r125 52 55 3.01551 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.205 $Y=4.735
+ $X2=1.065 $Y2=4.735
r126 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.87 $Y=4.735
+ $X2=1.955 $Y2=4.82
r127 51 52 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.87 $Y=4.735
+ $X2=1.205 $Y2=4.735
r128 47 57 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=1.1 $Y=5.61 $X2=1.1
+ $Y2=5.57
r129 47 49 22.0611 $w=3.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.1 $Y=5.61 $X2=1.1
+ $Y2=6.28
r130 45 55 3.49088 $w=2.67e-07 $l=9.12688e-08 $layer=LI1_cond $X=1.052 $Y=4.82
+ $X2=1.065 $Y2=4.735
r131 45 58 27.7942 $w=2.53e-07 $l=6.15e-07 $layer=LI1_cond $X=1.052 $Y=4.82
+ $X2=1.052 $Y2=5.435
r132 41 55 3.49088 $w=2.67e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=4.65
+ $X2=1.065 $Y2=4.735
r133 41 43 37.0428 $w=2.78e-07 $l=9e-07 $layer=LI1_cond $X=1.065 $Y=4.65
+ $X2=1.065 $Y2=3.75
r134 35 37 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.105 $Y=5.01
+ $X2=3.105 $Y2=5.275
r135 31 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.845 $Y=5.085
+ $X2=3.845 $Y2=5.01
r136 31 33 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.845 $Y=5.085
+ $X2=3.845 $Y2=5.925
r137 27 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.845 $Y=4.935
+ $X2=3.845 $Y2=5.01
r138 27 29 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.845 $Y=4.935
+ $X2=3.845 $Y2=4.01
r139 26 39 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=5.01 $X2=3.485
+ $Y2=5.01
r140 25 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=5.01
+ $X2=3.845 $Y2=5.01
r141 25 26 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.77 $Y=5.01
+ $X2=3.56 $Y2=5.01
r142 21 39 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=5.085
+ $X2=3.485 $Y2=5.01
r143 21 23 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.485 $Y=5.085
+ $X2=3.485 $Y2=5.925
r144 17 39 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.485 $Y=4.935
+ $X2=3.485 $Y2=5.01
r145 17 19 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.485 $Y=4.935
+ $X2=3.485 $Y2=4.01
r146 16 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.18 $Y=5.01
+ $X2=3.105 $Y2=5.01
r147 15 39 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=5.01 $X2=3.485
+ $Y2=5.01
r148 15 16 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.41 $Y=5.01
+ $X2=3.18 $Y2=5.01
r149 13 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.03 $Y=5.275
+ $X2=3.105 $Y2=5.275
r150 13 14 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.03 $Y=5.275
+ $X2=2.53 $Y2=5.275
r151 10 14 23.6571 $w=2.9e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.455 $Y=5.35
+ $X2=2.53 $Y2=5.275
r152 10 63 56.5103 $w=2.9e-07 $l=4.31648e-07 $layer=POLY_cond $X=2.455 $Y=5.35
+ $X2=2.115 $Y2=5.142
r153 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.455 $Y=5.35
+ $X2=2.455 $Y2=5.925
r154 7 65 18.1727 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=2.095 $Y=5.35
+ $X2=2.095 $Y2=5.142
r155 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.095 $Y=5.35
+ $X2=2.095 $Y2=5.925
r156 2 57 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=5.425 $X2=1.09 $Y2=5.57
r157 2 49 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.965
+ $Y=5.425 $X2=1.09 $Y2=6.28
r158 1 43 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=0.965
+ $Y=3.59 $X2=1.09 $Y2=3.75
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%VPWR 1 6 10 12 22 23 26
r24 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r25 22 23 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r26 20 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r27 19 22 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r28 19 20 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r29 17 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.74
+ $Y2=0
r30 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.2
+ $Y2=0
r31 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r32 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 12 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.74
+ $Y2=0
r34 12 14 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.24
+ $Y2=0
r35 10 23 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=4.56
+ $Y2=0
r36 10 20 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r37 6 8 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.74 $Y=0.38 $X2=0.74
+ $Y2=1.09
r38 4 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0
r39 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.38
r40 1 8 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.74 $Y2=1.09
r41 1 6 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.74 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%DESTPWR 1 2 9 13 18 19 20 29 38 39 42
r53 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=6.66
+ $X2=3.12 $Y2=6.66
r54 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=6.66
+ $X2=4.56 $Y2=6.66
r55 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=6.66
+ $X2=4.56 $Y2=6.66
r56 36 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=6.66
+ $X2=3.12 $Y2=6.66
r57 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=6.66 $X2=4.56
+ $Y2=6.66
r58 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=6.66 $X2=3.6
+ $Y2=6.66
r59 33 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=6.66
+ $X2=3.27 $Y2=6.66
r60 33 35 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=6.66
+ $X2=3.6 $Y2=6.66
r61 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=6.66
+ $X2=2.16 $Y2=6.66
r62 29 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=6.66
+ $X2=3.27 $Y2=6.66
r63 29 31 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.105 $Y=6.66
+ $X2=2.16 $Y2=6.66
r64 28 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=6.66
+ $X2=2.16 $Y2=6.66
r65 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=6.66
+ $X2=1.68 $Y2=6.66
r66 24 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=6.66
+ $X2=1.68 $Y2=6.66
r67 23 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=6.66
+ $X2=1.68 $Y2=6.66
r68 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=6.66
+ $X2=0.24 $Y2=6.66
r69 20 43 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=6.66
+ $X2=3.12 $Y2=6.66
r70 20 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=6.66
+ $X2=2.16 $Y2=6.66
r71 18 27 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.715 $Y=6.66
+ $X2=1.68 $Y2=6.66
r72 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=6.66
+ $X2=1.88 $Y2=6.66
r73 17 31 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.045 $Y=6.66
+ $X2=2.16 $Y2=6.66
r74 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=6.66
+ $X2=1.88 $Y2=6.66
r75 13 16 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=3.27 $Y=5.585
+ $X2=3.27 $Y2=6.3
r76 11 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=6.575
+ $X2=3.27 $Y2=6.66
r77 11 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.27 $Y=6.575
+ $X2=3.27 $Y2=6.3
r78 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=6.575 $X2=1.88
+ $Y2=6.66
r79 7 9 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=1.88 $Y=6.575
+ $X2=1.88 $Y2=5.78
r80 2 16 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=5.425 $X2=3.27 $Y2=6.3
r81 2 13 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=5.425 $X2=3.27 $Y2=5.585
r82 1 9 300 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=2 $X=1.74
+ $Y=5.425 $X2=1.88 $Y2=5.78
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUF_LP%X 1 2 7 8 9 10 11 12 20
r15 12 37 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=4.06 $Y=5.735
+ $X2=4.06 $Y2=6.28
r16 12 33 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=5.735
+ $X2=4.06 $Y2=5.57
r17 11 33 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.06 $Y=5.365
+ $X2=4.06 $Y2=5.57
r18 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.06 $Y=4.995
+ $X2=4.06 $Y2=5.365
r19 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.06 $Y=4.625
+ $X2=4.06 $Y2=4.995
r20 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.06 $Y=4.255 $X2=4.06
+ $Y2=4.625
r21 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.06 $Y=3.885 $X2=4.06
+ $Y2=4.255
r22 7 20 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.06 $Y=3.885
+ $X2=4.06 $Y2=3.735
r23 2 37 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=5.425 $X2=4.06 $Y2=6.28
r24 2 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=5.425 $X2=4.06 $Y2=5.57
r25 1 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.92
+ $Y=3.59 $X2=4.06 $Y2=3.735
.ends

