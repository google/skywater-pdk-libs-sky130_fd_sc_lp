* File: sky130_fd_sc_lp__nand3b_lp.pxi.spice
* Created: Wed Sep  2 10:05:06 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3B_LP%A_90_247# N_A_90_247#_M1004_d
+ N_A_90_247#_M1008_d N_A_90_247#_M1007_g N_A_90_247#_M1000_g N_A_90_247#_c_55_n
+ N_A_90_247#_c_56_n N_A_90_247#_c_65_n N_A_90_247#_c_66_n N_A_90_247#_c_57_n
+ N_A_90_247#_c_58_n N_A_90_247#_c_59_n N_A_90_247#_c_60_n N_A_90_247#_c_67_n
+ N_A_90_247#_c_61_n N_A_90_247#_c_62_n PM_SKY130_FD_SC_LP__NAND3B_LP%A_90_247#
x_PM_SKY130_FD_SC_LP__NAND3B_LP%B N_B_M1005_g N_B_M1003_g B N_B_c_124_n
+ PM_SKY130_FD_SC_LP__NAND3B_LP%B
x_PM_SKY130_FD_SC_LP__NAND3B_LP%C N_C_c_158_n N_C_M1002_g N_C_M1001_g
+ N_C_c_159_n C C N_C_c_161_n N_C_c_162_n PM_SKY130_FD_SC_LP__NAND3B_LP%C
x_PM_SKY130_FD_SC_LP__NAND3B_LP%A_N N_A_N_c_201_n N_A_N_M1006_g N_A_N_M1008_g
+ N_A_N_M1004_g N_A_N_c_204_n A_N A_N N_A_N_c_206_n
+ PM_SKY130_FD_SC_LP__NAND3B_LP%A_N
x_PM_SKY130_FD_SC_LP__NAND3B_LP%Y N_Y_M1000_s N_Y_M1007_s N_Y_M1003_d
+ N_Y_c_238_n N_Y_c_239_n N_Y_c_248_n N_Y_c_242_n N_Y_c_252_n Y Y Y
+ PM_SKY130_FD_SC_LP__NAND3B_LP%Y
x_PM_SKY130_FD_SC_LP__NAND3B_LP%VPWR N_VPWR_M1007_d N_VPWR_M1001_d
+ N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n
+ N_VPWR_c_288_n VPWR N_VPWR_c_289_n N_VPWR_c_282_n
+ PM_SKY130_FD_SC_LP__NAND3B_LP%VPWR
x_PM_SKY130_FD_SC_LP__NAND3B_LP%VGND N_VGND_M1002_d N_VGND_c_321_n VGND
+ N_VGND_c_322_n N_VGND_c_323_n N_VGND_c_324_n N_VGND_c_325_n
+ PM_SKY130_FD_SC_LP__NAND3B_LP%VGND
cc_1 VNB N_A_90_247#_c_55_n 0.0178627f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.235
cc_2 VNB N_A_90_247#_c_56_n 0.0195434f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.74
cc_3 VNB N_A_90_247#_c_57_n 0.0176104f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.4
cc_4 VNB N_A_90_247#_c_58_n 0.0354428f $X=-0.19 $Y=-0.245 $X2=2.435 $Y2=1.285
cc_5 VNB N_A_90_247#_c_59_n 0.00334294f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.285
cc_6 VNB N_A_90_247#_c_60_n 0.0138158f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=0.955
cc_7 VNB N_A_90_247#_c_61_n 0.0135364f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.06
cc_8 VNB N_A_90_247#_c_62_n 0.0130312f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.285
cc_9 VNB N_B_M1005_g 0.0318398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB B 0.00218746f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.58
cc_11 VNB N_B_c_124_n 0.0094845f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.915
cc_12 VNB N_C_c_158_n 0.0155405f $X=-0.19 $Y=-0.245 $X2=2.46 $Y2=0.705
cc_13 VNB N_C_c_159_n 0.0174687f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.915
cc_14 VNB C 0.00260783f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.235
cc_15 VNB N_C_c_161_n 0.0108875f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.4
cc_16 VNB N_C_c_162_n 0.0129954f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.4
cc_17 VNB N_A_N_c_201_n 0.0157664f $X=-0.19 $Y=-0.245 $X2=2.46 $Y2=0.705
cc_18 VNB N_A_N_M1008_g 5.60619e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_N_M1004_g 0.0313869f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.235
cc_20 VNB N_A_N_c_204_n 0.0183516f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.915
cc_21 VNB A_N 0.0263767f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.235
cc_22 VNB N_A_N_c_206_n 0.049481f $X=-0.19 $Y=-0.245 $X2=2.435 $Y2=1.285
cc_23 VNB N_Y_c_238_n 0.0289631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_239_n 0.0305506f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.235
cc_25 VNB Y 0.0179284f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.285
cc_26 VNB N_VPWR_c_282_n 0.123877f $X=-0.19 $Y=-0.245 $X2=2.52 $Y2=2.225
cc_27 VNB N_VGND_c_321_n 0.0214469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_322_n 0.0430497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_323_n 0.0279052f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.4
cc_30 VNB N_VGND_c_324_n 0.197499f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.4
cc_31 VNB N_VGND_c_325_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.285
cc_32 VPB N_A_90_247#_M1007_g 0.0302088f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.58
cc_33 VPB N_A_90_247#_c_56_n 0.00637818f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.74
cc_34 VPB N_A_90_247#_c_65_n 0.0147548f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.905
cc_35 VPB N_A_90_247#_c_66_n 7.54448e-19 $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.4
cc_36 VPB N_A_90_247#_c_67_n 0.0495349f $X=-0.19 $Y=1.655 $X2=2.52 $Y2=2.225
cc_37 VPB N_A_90_247#_c_61_n 0.0197033f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.06
cc_38 VPB N_B_M1003_g 0.0257346f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.905
cc_39 VPB B 7.38391e-19 $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.58
cc_40 VPB N_B_c_124_n 0.020666f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.915
cc_41 VPB N_C_M1001_g 0.0286488f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.58
cc_42 VPB C 0.00430931f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.235
cc_43 VPB N_C_c_161_n 0.0150198f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.4
cc_44 VPB N_A_N_M1008_g 0.0481122f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_Y_c_239_n 0.0206871f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=1.235
cc_46 VPB N_Y_c_242_n 0.0430018f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.4
cc_47 VPB N_VPWR_c_283_n 8.75318e-19 $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.58
cc_48 VPB N_VPWR_c_284_n 0.00609586f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.915
cc_49 VPB N_VPWR_c_285_n 0.0203637f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.37
cc_50 VPB N_VPWR_c_286_n 0.00455177f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.4
cc_51 VPB N_VPWR_c_287_n 0.0182443f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.4
cc_52 VPB N_VPWR_c_288_n 0.00522215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_289_n 0.022723f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.225
cc_54 VPB N_VPWR_c_282_n 0.053496f $X=-0.19 $Y=1.655 $X2=2.52 $Y2=2.225
cc_55 N_A_90_247#_c_55_n N_B_M1005_g 0.0561901f $X=0.615 $Y=1.235 $X2=0 $Y2=0
cc_56 N_A_90_247#_c_66_n N_B_M1005_g 0.00120662f $X=0.615 $Y=1.4 $X2=0 $Y2=0
cc_57 N_A_90_247#_c_58_n N_B_M1005_g 0.0101086f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_58 N_A_90_247#_M1007_g N_B_M1003_g 0.0424582f $X=0.625 $Y=2.58 $X2=0 $Y2=0
cc_59 N_A_90_247#_c_56_n B 0.00133772f $X=0.615 $Y=1.74 $X2=0 $Y2=0
cc_60 N_A_90_247#_c_66_n B 0.0226338f $X=0.615 $Y=1.4 $X2=0 $Y2=0
cc_61 N_A_90_247#_c_58_n B 0.0241149f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_62 N_A_90_247#_M1007_g N_B_c_124_n 8.41017e-19 $X=0.625 $Y=2.58 $X2=0 $Y2=0
cc_63 N_A_90_247#_c_56_n N_B_c_124_n 0.0191658f $X=0.615 $Y=1.74 $X2=0 $Y2=0
cc_64 N_A_90_247#_c_66_n N_B_c_124_n 0.00109648f $X=0.615 $Y=1.4 $X2=0 $Y2=0
cc_65 N_A_90_247#_c_58_n N_B_c_124_n 0.00110374f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_66 N_A_90_247#_c_67_n N_C_M1001_g 2.81111e-19 $X=2.52 $Y=2.225 $X2=0 $Y2=0
cc_67 N_A_90_247#_c_58_n N_C_c_159_n 0.0167459f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_68 N_A_90_247#_c_58_n C 0.0519034f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_69 N_A_90_247#_c_61_n C 0.0163183f $X=2.56 $Y=2.06 $X2=0 $Y2=0
cc_70 N_A_90_247#_c_58_n N_C_c_161_n 0.00439954f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_71 N_A_90_247#_c_58_n N_C_c_162_n 0.00298719f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_72 N_A_90_247#_c_58_n N_A_N_c_201_n 0.00988853f $X=2.435 $Y=1.285 $X2=-0.19
+ $Y2=-0.245
cc_73 N_A_90_247#_c_60_n N_A_N_c_201_n 0.00139038f $X=2.6 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_74 N_A_90_247#_c_67_n N_A_N_M1008_g 0.022155f $X=2.52 $Y=2.225 $X2=0 $Y2=0
cc_75 N_A_90_247#_c_61_n N_A_N_M1008_g 0.00957836f $X=2.56 $Y=2.06 $X2=0 $Y2=0
cc_76 N_A_90_247#_c_58_n N_A_N_M1004_g 0.0130701f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_77 N_A_90_247#_c_60_n N_A_N_M1004_g 0.0079225f $X=2.6 $Y=0.955 $X2=0 $Y2=0
cc_78 N_A_90_247#_c_61_n N_A_N_M1004_g 0.00719872f $X=2.56 $Y=2.06 $X2=0 $Y2=0
cc_79 N_A_90_247#_c_62_n N_A_N_M1004_g 0.00492103f $X=2.6 $Y=1.285 $X2=0 $Y2=0
cc_80 N_A_90_247#_c_58_n N_A_N_c_204_n 0.00557189f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_81 N_A_90_247#_c_67_n N_A_N_c_204_n 0.00298743f $X=2.52 $Y=2.225 $X2=0 $Y2=0
cc_82 N_A_90_247#_c_58_n A_N 0.0128377f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_83 N_A_90_247#_c_60_n A_N 0.0235024f $X=2.6 $Y=0.955 $X2=0 $Y2=0
cc_84 N_A_90_247#_M1007_g N_Y_c_239_n 0.00600702f $X=0.625 $Y=2.58 $X2=0 $Y2=0
cc_85 N_A_90_247#_c_55_n N_Y_c_239_n 0.00483579f $X=0.615 $Y=1.235 $X2=0 $Y2=0
cc_86 N_A_90_247#_c_66_n N_Y_c_239_n 0.0384063f $X=0.615 $Y=1.4 $X2=0 $Y2=0
cc_87 N_A_90_247#_c_57_n N_Y_c_239_n 0.0128179f $X=0.615 $Y=1.4 $X2=0 $Y2=0
cc_88 N_A_90_247#_c_59_n N_Y_c_239_n 0.0131681f $X=0.78 $Y=1.285 $X2=0 $Y2=0
cc_89 N_A_90_247#_M1007_g N_Y_c_248_n 0.0179867f $X=0.625 $Y=2.58 $X2=0 $Y2=0
cc_90 N_A_90_247#_c_66_n N_Y_c_248_n 0.0164626f $X=0.615 $Y=1.4 $X2=0 $Y2=0
cc_91 N_A_90_247#_M1007_g N_Y_c_242_n 0.0209867f $X=0.625 $Y=2.58 $X2=0 $Y2=0
cc_92 N_A_90_247#_c_66_n N_Y_c_242_n 0.00397635f $X=0.615 $Y=1.4 $X2=0 $Y2=0
cc_93 N_A_90_247#_M1007_g N_Y_c_252_n 0.00100717f $X=0.625 $Y=2.58 $X2=0 $Y2=0
cc_94 N_A_90_247#_c_55_n Y 0.0184607f $X=0.615 $Y=1.235 $X2=0 $Y2=0
cc_95 N_A_90_247#_c_57_n Y 0.00108959f $X=0.615 $Y=1.4 $X2=0 $Y2=0
cc_96 N_A_90_247#_c_58_n Y 0.0335495f $X=2.435 $Y=1.285 $X2=0 $Y2=0
cc_97 N_A_90_247#_c_59_n Y 0.025185f $X=0.78 $Y=1.285 $X2=0 $Y2=0
cc_98 N_A_90_247#_M1007_g N_VPWR_c_283_n 0.0197097f $X=0.625 $Y=2.58 $X2=0 $Y2=0
cc_99 N_A_90_247#_c_67_n N_VPWR_c_284_n 0.0301865f $X=2.52 $Y=2.225 $X2=0 $Y2=0
cc_100 N_A_90_247#_M1007_g N_VPWR_c_285_n 0.00818185f $X=0.625 $Y=2.58 $X2=0
+ $Y2=0
cc_101 N_A_90_247#_c_67_n N_VPWR_c_289_n 0.025152f $X=2.52 $Y=2.225 $X2=0 $Y2=0
cc_102 N_A_90_247#_M1007_g N_VPWR_c_282_n 0.0145557f $X=0.625 $Y=2.58 $X2=0
+ $Y2=0
cc_103 N_A_90_247#_c_67_n N_VPWR_c_282_n 0.015666f $X=2.52 $Y=2.225 $X2=0 $Y2=0
cc_104 N_A_90_247#_c_58_n N_VGND_c_321_n 0.0227959f $X=2.435 $Y=1.285 $X2=0
+ $Y2=0
cc_105 N_A_90_247#_c_60_n N_VGND_c_321_n 0.00510094f $X=2.6 $Y=0.955 $X2=0 $Y2=0
cc_106 N_A_90_247#_c_55_n N_VGND_c_322_n 5.6543e-19 $X=0.615 $Y=1.235 $X2=0
+ $Y2=0
cc_107 N_A_90_247#_c_60_n N_VGND_c_324_n 9.36254e-19 $X=2.6 $Y=0.955 $X2=0 $Y2=0
cc_108 N_B_M1005_g N_C_c_158_n 0.0405804f $X=1.095 $Y=0.915 $X2=-0.19 $Y2=-0.245
cc_109 N_B_M1003_g N_C_M1001_g 0.0263669f $X=1.155 $Y=2.58 $X2=0 $Y2=0
cc_110 B C 0.0200938f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_111 N_B_c_124_n C 0.00106198f $X=1.155 $Y=1.755 $X2=0 $Y2=0
cc_112 B N_C_c_161_n 8.02603e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_113 N_B_c_124_n N_C_c_161_n 0.0177681f $X=1.155 $Y=1.755 $X2=0 $Y2=0
cc_114 N_B_M1005_g N_C_c_162_n 0.00847105f $X=1.095 $Y=0.915 $X2=0 $Y2=0
cc_115 N_B_M1003_g N_Y_c_248_n 0.0178513f $X=1.155 $Y=2.58 $X2=0 $Y2=0
cc_116 B N_Y_c_248_n 0.016964f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_117 N_B_M1003_g N_Y_c_242_n 0.00100361f $X=1.155 $Y=2.58 $X2=0 $Y2=0
cc_118 N_B_M1003_g N_Y_c_252_n 0.0177728f $X=1.155 $Y=2.58 $X2=0 $Y2=0
cc_119 B N_Y_c_252_n 0.00332706f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_120 N_B_M1005_g Y 0.0183811f $X=1.095 $Y=0.915 $X2=0 $Y2=0
cc_121 N_B_M1003_g N_VPWR_c_283_n 0.0187576f $X=1.155 $Y=2.58 $X2=0 $Y2=0
cc_122 N_B_M1003_g N_VPWR_c_284_n 0.00132364f $X=1.155 $Y=2.58 $X2=0 $Y2=0
cc_123 N_B_M1003_g N_VPWR_c_287_n 0.00818185f $X=1.155 $Y=2.58 $X2=0 $Y2=0
cc_124 N_B_M1003_g N_VPWR_c_282_n 0.0136091f $X=1.155 $Y=2.58 $X2=0 $Y2=0
cc_125 N_B_M1005_g N_VGND_c_321_n 3.72866e-19 $X=1.095 $Y=0.915 $X2=0 $Y2=0
cc_126 N_B_M1005_g N_VGND_c_322_n 5.6543e-19 $X=1.095 $Y=0.915 $X2=0 $Y2=0
cc_127 N_C_c_159_n N_A_N_c_201_n 0.00301839f $X=1.635 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_128 C N_A_N_c_201_n 8.2243e-19 $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_129 N_C_M1001_g N_A_N_M1008_g 0.0147288f $X=1.685 $Y=2.58 $X2=0 $Y2=0
cc_130 C N_A_N_M1008_g 0.0152463f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_131 N_C_c_159_n N_A_N_M1004_g 0.00470697f $X=1.635 $Y=1.275 $X2=0 $Y2=0
cc_132 C N_A_N_c_204_n 0.00452923f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_133 N_C_c_161_n N_A_N_c_204_n 0.0181257f $X=1.725 $Y=1.715 $X2=0 $Y2=0
cc_134 N_C_c_162_n N_A_N_c_204_n 0.00203968f $X=1.725 $Y=1.55 $X2=0 $Y2=0
cc_135 N_C_c_158_n N_A_N_c_206_n 0.0129651f $X=1.485 $Y=1.2 $X2=0 $Y2=0
cc_136 N_C_M1001_g N_Y_c_252_n 0.0198306f $X=1.685 $Y=2.58 $X2=0 $Y2=0
cc_137 C N_Y_c_252_n 0.00158785f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_138 N_C_c_158_n Y 0.00349806f $X=1.485 $Y=1.2 $X2=0 $Y2=0
cc_139 N_C_M1001_g N_VPWR_c_283_n 0.0011034f $X=1.685 $Y=2.58 $X2=0 $Y2=0
cc_140 N_C_M1001_g N_VPWR_c_284_n 0.022734f $X=1.685 $Y=2.58 $X2=0 $Y2=0
cc_141 C N_VPWR_c_284_n 0.0273201f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_142 N_C_c_161_n N_VPWR_c_284_n 0.00185447f $X=1.725 $Y=1.715 $X2=0 $Y2=0
cc_143 N_C_M1001_g N_VPWR_c_287_n 0.00818185f $X=1.685 $Y=2.58 $X2=0 $Y2=0
cc_144 N_C_M1001_g N_VPWR_c_282_n 0.0136091f $X=1.685 $Y=2.58 $X2=0 $Y2=0
cc_145 N_C_c_158_n N_VGND_c_321_n 0.00752086f $X=1.485 $Y=1.2 $X2=0 $Y2=0
cc_146 N_C_c_159_n N_VGND_c_321_n 0.00388286f $X=1.635 $Y=1.275 $X2=0 $Y2=0
cc_147 N_C_c_158_n N_VGND_c_322_n 0.0031218f $X=1.485 $Y=1.2 $X2=0 $Y2=0
cc_148 N_C_c_158_n N_VGND_c_324_n 0.00376215f $X=1.485 $Y=1.2 $X2=0 $Y2=0
cc_149 N_A_N_M1008_g N_VPWR_c_284_n 0.00336873f $X=2.255 $Y=2.58 $X2=0 $Y2=0
cc_150 N_A_N_M1008_g N_VPWR_c_289_n 0.00914935f $X=2.255 $Y=2.58 $X2=0 $Y2=0
cc_151 N_A_N_M1008_g N_VPWR_c_282_n 0.0169826f $X=2.255 $Y=2.58 $X2=0 $Y2=0
cc_152 A_N N_VGND_c_321_n 0.0324453f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_153 N_A_N_c_206_n N_VGND_c_321_n 0.0167463f $X=2.385 $Y=0.43 $X2=0 $Y2=0
cc_154 A_N N_VGND_c_323_n 0.0444402f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_155 N_A_N_c_206_n N_VGND_c_323_n 0.0140846f $X=2.385 $Y=0.43 $X2=0 $Y2=0
cc_156 A_N N_VGND_c_324_n 0.0268292f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A_N_c_206_n N_VGND_c_324_n 0.018165f $X=2.385 $Y=0.43 $X2=0 $Y2=0
cc_158 N_Y_c_248_n N_VPWR_M1007_d 0.00814128f $X=1.255 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_159 N_Y_c_248_n N_VPWR_c_283_n 0.0164319f $X=1.255 $Y=2.185 $X2=0 $Y2=0
cc_160 N_Y_c_242_n N_VPWR_c_283_n 0.0413224f $X=0.36 $Y=2.25 $X2=0 $Y2=0
cc_161 N_Y_c_252_n N_VPWR_c_283_n 0.0405228f $X=1.42 $Y=2.265 $X2=0 $Y2=0
cc_162 N_Y_c_252_n N_VPWR_c_284_n 0.0642563f $X=1.42 $Y=2.265 $X2=0 $Y2=0
cc_163 N_Y_c_242_n N_VPWR_c_285_n 0.0261633f $X=0.36 $Y=2.25 $X2=0 $Y2=0
cc_164 N_Y_c_252_n N_VPWR_c_287_n 0.0177952f $X=1.42 $Y=2.265 $X2=0 $Y2=0
cc_165 N_Y_c_242_n N_VPWR_c_282_n 0.0162464f $X=0.36 $Y=2.25 $X2=0 $Y2=0
cc_166 N_Y_c_252_n N_VPWR_c_282_n 0.0124497f $X=1.42 $Y=2.265 $X2=0 $Y2=0
cc_167 Y A_156_141# 0.0014282f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_168 Y A_234_141# 0.00386746f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_169 Y N_VGND_c_321_n 0.0401799f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_170 N_Y_c_238_n N_VGND_c_322_n 0.00555891f $X=0.185 $Y=1.02 $X2=0 $Y2=0
cc_171 Y N_VGND_c_322_n 0.0336569f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_172 N_Y_c_238_n N_VGND_c_324_n 0.00592732f $X=0.185 $Y=1.02 $X2=0 $Y2=0
cc_173 Y N_VGND_c_324_n 0.0361737f $X=1.115 $Y=0.47 $X2=0 $Y2=0
