* File: sky130_fd_sc_lp__clkinvlp_2.spice
* Created: Wed Sep  2 09:41:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkinvlp_2.pex.spice"
.subckt sky130_fd_sc_lp__clkinvlp_2  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 A_185_67# N_A_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.55 AD=0.066
+ AS=0.15675 PD=0.79 PS=1.67 NRD=14.172 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_185_67# VNB NSHORT L=0.15 W=0.55 AD=0.15675
+ AS=0.066 PD=1.67 PS=0.79 NRD=0 NRS=14.172 M=1 R=3.66667 SA=75000.6 SB=75000.2
+ A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000 A=0.25 P=2.5
+ MULT=1
DX4_noxref VNB VPB NWDIODE A=4.2895 P=8.33
*
.include "sky130_fd_sc_lp__clkinvlp_2.pxi.spice"
*
.ends
*
*
