* File: sky130_fd_sc_lp__inv_1.pex.spice
* Created: Fri Aug 28 10:38:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INV_1%A 3 6 8 9 13 15
r18 13 16 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.372 $Y=1.375
+ $X2=0.372 $Y2=1.54
r19 13 15 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.372 $Y=1.375
+ $X2=0.372 $Y2=1.21
r20 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.375 $X2=0.35 $Y2=1.375
r21 9 14 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=1.375
r22 8 14 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=0.26 $Y=1.295 $X2=0.26
+ $Y2=1.375
r23 6 16 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.485 $Y=2.465
+ $X2=0.485 $Y2=1.54
r24 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.485 $Y=0.68
+ $X2=0.485 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__INV_1%VPWR 1 4 6 10 14 15
r13 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r14 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r15 12 18 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r16 12 14 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r17 10 15 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=3.33
+ $X2=0.72 $Y2=3.33
r18 10 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=3.33
+ $X2=0.24 $Y2=3.33
r19 6 9 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.27 $Y=2.005
+ $X2=0.27 $Y2=2.95
r20 4 18 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r21 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.95
r22 1 9 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.95
r23 1 6 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__INV_1%Y 1 2 7 8 9 10 11 12 13 22
r10 13 40 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.74 $Y=2.775
+ $X2=0.74 $Y2=2.91
r11 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=2.405
+ $X2=0.74 $Y2=2.775
r12 11 12 16.6464 $w=2.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.74 $Y=2.015
+ $X2=0.74 $Y2=2.405
r13 10 11 14.9391 $w=2.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.74 $Y=1.665
+ $X2=0.74 $Y2=2.015
r14 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=1.295
+ $X2=0.74 $Y2=1.665
r15 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=0.925 $X2=0.74
+ $Y2=1.295
r16 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=0.555 $X2=0.74
+ $Y2=0.925
r17 7 22 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.74 $Y=0.555
+ $X2=0.74 $Y2=0.42
r18 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=2.91
r19 2 11 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=0.56 $Y=1.835
+ $X2=0.7 $Y2=2.015
r20 1 22 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.26 $X2=0.7 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__INV_1%VGND 1 4 6 8 12 13
r12 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r13 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r14 10 16 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r15 10 12 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.72
+ $Y2=0
r16 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r17 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r18 4 16 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.217 $Y2=0
r19 4 6 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.27 $Y=0.085 $X2=0.27
+ $Y2=0.405
r20 1 6 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.26 $X2=0.27 $Y2=0.405
.ends

