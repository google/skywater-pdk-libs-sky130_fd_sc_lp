* File: sky130_fd_sc_lp__o221ai_0.pxi.spice
* Created: Wed Sep  2 10:18:55 2020
* 
x_PM_SKY130_FD_SC_LP__O221AI_0%C1 N_C1_M1002_g N_C1_M1001_g C1 N_C1_c_76_n
+ N_C1_c_77_n PM_SKY130_FD_SC_LP__O221AI_0%C1
x_PM_SKY130_FD_SC_LP__O221AI_0%B1 N_B1_M1006_g N_B1_M1003_g B1 B1 B1
+ N_B1_c_110_n N_B1_c_111_n N_B1_c_112_n PM_SKY130_FD_SC_LP__O221AI_0%B1
x_PM_SKY130_FD_SC_LP__O221AI_0%B2 N_B2_M1005_g N_B2_M1007_g N_B2_c_158_n B2 B2
+ B2 B2 B2 B2 B2 N_B2_c_162_n N_B2_c_163_n N_B2_c_159_n N_B2_c_165_n
+ N_B2_c_166_n PM_SKY130_FD_SC_LP__O221AI_0%B2
x_PM_SKY130_FD_SC_LP__O221AI_0%A2 N_A2_c_215_n N_A2_M1009_g N_A2_c_216_n
+ N_A2_M1008_g N_A2_c_218_n A2 A2 N_A2_c_220_n PM_SKY130_FD_SC_LP__O221AI_0%A2
x_PM_SKY130_FD_SC_LP__O221AI_0%A1 N_A1_c_264_n N_A1_c_265_n N_A1_M1000_g
+ N_A1_M1004_g A1 A1 N_A1_c_268_n PM_SKY130_FD_SC_LP__O221AI_0%A1
x_PM_SKY130_FD_SC_LP__O221AI_0%Y N_Y_M1002_s N_Y_M1001_s N_Y_M1005_d N_Y_c_306_n
+ N_Y_c_307_n N_Y_c_308_n N_Y_c_311_n N_Y_c_312_n N_Y_c_313_n N_Y_c_339_n Y Y Y
+ N_Y_c_316_n PM_SKY130_FD_SC_LP__O221AI_0%Y
x_PM_SKY130_FD_SC_LP__O221AI_0%VPWR N_VPWR_M1001_d N_VPWR_M1000_d N_VPWR_c_373_n
+ N_VPWR_c_374_n N_VPWR_c_375_n N_VPWR_c_376_n VPWR N_VPWR_c_377_n
+ N_VPWR_c_378_n N_VPWR_c_372_n N_VPWR_c_380_n PM_SKY130_FD_SC_LP__O221AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O221AI_0%A_110_47# N_A_110_47#_M1002_d N_A_110_47#_M1007_d
+ N_A_110_47#_c_416_n N_A_110_47#_c_417_n N_A_110_47#_c_418_n
+ N_A_110_47#_c_419_n N_A_110_47#_c_424_n N_A_110_47#_c_420_n
+ N_A_110_47#_c_421_n PM_SKY130_FD_SC_LP__O221AI_0%A_110_47#
x_PM_SKY130_FD_SC_LP__O221AI_0%A_196_47# N_A_196_47#_M1006_d N_A_196_47#_M1004_d
+ N_A_196_47#_c_460_n N_A_196_47#_c_461_n N_A_196_47#_c_462_n
+ PM_SKY130_FD_SC_LP__O221AI_0%A_196_47#
x_PM_SKY130_FD_SC_LP__O221AI_0%VGND N_VGND_M1009_d VGND N_VGND_c_487_n
+ N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n PM_SKY130_FD_SC_LP__O221AI_0%VGND
cc_1 VNB N_C1_M1002_g 0.0669274f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_2 VNB N_B1_M1006_g 0.0354996f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_3 VNB N_B1_M1003_g 0.0105208f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.66
cc_4 VNB B1 0.00298006f $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=2.015
cc_5 VNB N_B1_c_110_n 0.0306622f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.035
cc_6 VNB N_B1_c_111_n 0.00495294f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.035
cc_7 VNB N_B1_c_112_n 0.00277472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B2_M1007_g 0.0366287f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.66
cc_9 VNB N_B2_c_158_n 0.0314944f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.015
cc_10 VNB N_B2_c_159_n 0.0320192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_c_215_n 0.0220083f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.85
cc_12 VNB N_A2_c_216_n 0.0239831f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.18
cc_13 VNB N_A2_M1008_g 7.66603e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_218_n 0.0168826f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.015
cc_15 VNB A2 0.002421f $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=2.18
cc_16 VNB N_A2_c_220_n 0.0514733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_264_n 0.00559992f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.85
cc_18 VNB N_A1_c_265_n 0.0156622f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_19 VNB N_A1_M1004_g 0.0411954f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_20 VNB A1 0.018763f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.015
cc_21 VNB N_A1_c_268_n 0.0273022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_306_n 0.0629768f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.015
cc_23 VNB N_Y_c_307_n 0.00430949f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.035
cc_24 VNB N_Y_c_308_n 0.00340131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_372_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_110_47#_c_416_n 0.00187888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_110_47#_c_417_n 0.00154943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_110_47#_c_418_n 0.0278676f $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=2.015
cc_29 VNB N_A_110_47#_c_419_n 0.0259787f $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=2.18
cc_30 VNB N_A_110_47#_c_420_n 0.0101998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_110_47#_c_421_n 0.00189664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_196_47#_c_460_n 0.00671863f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.66
cc_33 VNB N_A_196_47#_c_461_n 0.00240564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_196_47#_c_462_n 0.00281026f $X=-0.19 $Y=-0.245 $X2=0.447 $Y2=2.18
cc_35 VNB N_VGND_c_487_n 0.0348703f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=2.035
cc_36 VNB N_VGND_c_488_n 0.196384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_489_n 0.0402677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_490_n 0.0180777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_C1_M1002_g 0.0142341f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_40 VPB N_C1_M1001_g 0.0264848f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.66
cc_41 VPB N_C1_c_76_n 0.0431145f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.015
cc_42 VPB N_C1_c_77_n 0.0149865f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.015
cc_43 VPB N_B1_M1003_g 0.0456465f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.66
cc_44 VPB B1 0.00362337f $X=-0.19 $Y=1.655 $X2=0.447 $Y2=2.015
cc_45 VPB N_B2_M1005_g 0.0205255f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_46 VPB B2 0.0473548f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B2_c_162_n 0.032857f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_B2_c_163_n 0.0455465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B2_c_159_n 0.0141126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B2_c_165_n 0.0365685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B2_c_166_n 0.00894607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A2_M1008_g 0.0472716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB A2 0.00553239f $X=-0.19 $Y=1.655 $X2=0.447 $Y2=2.18
cc_54 VPB N_A1_M1000_g 0.0456714f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.18
cc_55 VPB A1 0.00967846f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.015
cc_56 VPB N_A1_c_268_n 0.0176014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_307_n 0.00257612f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.035
cc_58 VPB N_Y_c_308_n 0.00642699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_Y_c_311_n 0.001961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_Y_c_312_n 0.00459857f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_Y_c_313_n 0.0305535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB Y 0.00269486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB Y 0.00304467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_Y_c_316_n 0.003013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_373_n 0.00344978f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_66 VPB N_VPWR_c_374_n 0.0239291f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=2.015
cc_67 VPB N_VPWR_c_375_n 0.0422209f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.035
cc_68 VPB N_VPWR_c_376_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_377_n 0.0193281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_378_n 0.0209635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_372_n 0.0798338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_380_n 0.00577233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 N_C1_M1002_g N_B1_M1006_g 0.0437518f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_74 N_C1_M1002_g N_B1_M1003_g 0.011483f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_75 N_C1_c_76_n N_B1_M1003_g 0.0379567f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_76 N_C1_c_77_n N_B1_M1003_g 2.08226e-19 $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_77 N_C1_M1002_g B1 2.0569e-19 $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_78 N_C1_M1002_g N_B1_c_111_n 0.00436131f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_79 N_C1_M1002_g N_Y_c_306_n 0.0280011f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_80 N_C1_M1002_g N_Y_c_307_n 0.0167374f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_81 N_C1_c_76_n N_Y_c_307_n 0.00367942f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_82 N_C1_c_77_n N_Y_c_307_n 0.0154903f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_83 N_C1_c_76_n N_Y_c_308_n 0.00278981f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_84 N_C1_c_77_n N_Y_c_308_n 0.0228504f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_85 N_C1_M1001_g N_Y_c_311_n 0.0105124f $X=0.565 $Y=2.66 $X2=0 $Y2=0
cc_86 N_C1_c_76_n N_Y_c_311_n 0.00122594f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_87 N_C1_c_77_n N_Y_c_311_n 0.00984566f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_88 N_C1_M1002_g N_Y_c_312_n 0.00202314f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_89 N_C1_c_76_n N_Y_c_312_n 0.00696309f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_90 N_C1_c_77_n N_Y_c_312_n 0.0170248f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_91 N_C1_M1001_g N_Y_c_313_n 4.46816e-19 $X=0.565 $Y=2.66 $X2=0 $Y2=0
cc_92 N_C1_c_76_n N_Y_c_313_n 0.00476468f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_93 N_C1_c_77_n N_Y_c_313_n 0.0216736f $X=0.42 $Y=2.015 $X2=0 $Y2=0
cc_94 N_C1_M1001_g N_VPWR_c_373_n 0.0101777f $X=0.565 $Y=2.66 $X2=0 $Y2=0
cc_95 N_C1_M1001_g N_VPWR_c_377_n 0.00396895f $X=0.565 $Y=2.66 $X2=0 $Y2=0
cc_96 N_C1_M1001_g N_VPWR_c_372_n 0.00417037f $X=0.565 $Y=2.66 $X2=0 $Y2=0
cc_97 N_C1_M1002_g N_A_110_47#_c_416_n 0.00420848f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_98 N_C1_M1002_g N_A_110_47#_c_417_n 0.00369885f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_99 N_C1_M1002_g N_A_110_47#_c_424_n 0.00319146f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_100 N_C1_M1002_g N_VGND_c_488_n 0.0118279f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_101 N_C1_M1002_g N_VGND_c_489_n 0.0057945f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_102 N_B1_M1003_g N_B2_c_162_n 0.0765402f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_103 B1 N_B2_c_162_n 2.67885e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B1_M1003_g N_B2_c_165_n 0.00154505f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_105 B1 N_B2_c_165_n 0.0153789f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_106 N_B1_c_110_n N_B2_c_165_n 2.02426e-19 $X=0.995 $Y=1.3 $X2=0 $Y2=0
cc_107 N_B1_M1006_g N_A2_c_215_n 0.0202874f $X=0.905 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_108 N_B1_M1006_g N_A2_c_216_n 0.00685452f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_109 N_B1_c_110_n N_A2_c_216_n 0.0211028f $X=0.995 $Y=1.3 $X2=0 $Y2=0
cc_110 N_B1_c_112_n N_A2_c_216_n 0.00378617f $X=1.197 $Y=1.41 $X2=0 $Y2=0
cc_111 B1 N_A2_M1008_g 3.97202e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_112 B1 A2 0.0285615f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_113 N_B1_c_112_n A2 0.00882527f $X=1.197 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B1_M1003_g N_A2_c_220_n 0.00617591f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_115 B1 N_A2_c_220_n 0.00186509f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_116 N_B1_c_111_n N_Y_c_306_n 0.0156699f $X=1.105 $Y=1.31 $X2=0 $Y2=0
cc_117 N_B1_M1003_g N_Y_c_307_n 0.00436839f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_118 B1 N_Y_c_307_n 0.0136669f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_119 N_B1_c_110_n N_Y_c_307_n 0.00261783f $X=0.995 $Y=1.3 $X2=0 $Y2=0
cc_120 N_B1_c_111_n N_Y_c_307_n 0.0307431f $X=1.105 $Y=1.31 $X2=0 $Y2=0
cc_121 N_B1_M1003_g N_Y_c_312_n 0.0140897f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_122 B1 N_Y_c_312_n 6.86112e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_123 N_B1_M1003_g N_Y_c_339_n 0.00243966f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_124 N_B1_M1003_g N_Y_c_316_n 0.0125795f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_125 N_B1_M1003_g N_VPWR_c_373_n 0.0100983f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_126 N_B1_M1003_g N_VPWR_c_375_n 0.00396895f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_127 N_B1_M1003_g N_VPWR_c_372_n 0.00394667f $X=0.995 $Y=2.66 $X2=0 $Y2=0
cc_128 N_B1_M1006_g N_A_110_47#_c_416_n 0.00430038f $X=0.905 $Y=0.445 $X2=0
+ $Y2=0
cc_129 N_B1_c_111_n N_A_110_47#_c_417_n 0.0144772f $X=1.105 $Y=1.31 $X2=0 $Y2=0
cc_130 N_B1_M1006_g N_A_110_47#_c_424_n 0.0029226f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_131 N_B1_M1006_g N_A_110_47#_c_420_n 0.0151882f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_132 N_B1_c_110_n N_A_110_47#_c_420_n 0.00479399f $X=0.995 $Y=1.3 $X2=0 $Y2=0
cc_133 N_B1_c_111_n N_A_110_47#_c_420_n 0.0280382f $X=1.105 $Y=1.31 $X2=0 $Y2=0
cc_134 N_B1_c_112_n N_A_110_47#_c_420_n 0.0151134f $X=1.197 $Y=1.41 $X2=0 $Y2=0
cc_135 N_B1_M1006_g N_A_196_47#_c_461_n 5.04263e-19 $X=0.905 $Y=0.445 $X2=0
+ $Y2=0
cc_136 N_B1_M1006_g N_VGND_c_488_n 0.0108508f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_137 N_B1_M1006_g N_VGND_c_489_n 0.0057945f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_138 N_B2_M1005_g N_A2_M1008_g 0.0177735f $X=1.355 $Y=2.66 $X2=0 $Y2=0
cc_139 N_B2_c_162_n N_A2_M1008_g 0.0219978f $X=1.445 $Y=2.015 $X2=0 $Y2=0
cc_140 N_B2_c_165_n N_A2_M1008_g 0.0155352f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_141 N_B2_c_162_n A2 0.0010273f $X=1.445 $Y=2.015 $X2=0 $Y2=0
cc_142 N_B2_c_159_n A2 6.44287e-19 $X=3.085 $Y=1.85 $X2=0 $Y2=0
cc_143 N_B2_c_165_n A2 0.0650349f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_144 N_B2_c_162_n N_A2_c_220_n 0.0160999f $X=1.445 $Y=2.015 $X2=0 $Y2=0
cc_145 N_B2_c_165_n N_A2_c_220_n 0.00182325f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_146 N_B2_c_158_n N_A1_c_264_n 0.0171913f $X=2.995 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_147 N_B2_c_159_n N_A1_c_265_n 0.00494747f $X=3.085 $Y=1.85 $X2=0 $Y2=0
cc_148 B2 N_A1_M1000_g 0.00467259f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_149 N_B2_c_159_n N_A1_M1000_g 0.00854828f $X=3.085 $Y=1.85 $X2=0 $Y2=0
cc_150 N_B2_c_165_n N_A1_M1000_g 0.0192331f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_151 N_B2_M1007_g N_A1_M1004_g 0.0171913f $X=2.695 $Y=0.445 $X2=0 $Y2=0
cc_152 N_B2_c_158_n A1 0.00522893f $X=2.995 $Y=1.135 $X2=0 $Y2=0
cc_153 N_B2_c_163_n A1 0.00449931f $X=3.085 $Y=2.015 $X2=0 $Y2=0
cc_154 N_B2_c_159_n A1 0.0186294f $X=3.085 $Y=1.85 $X2=0 $Y2=0
cc_155 N_B2_c_165_n A1 0.0387743f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_156 N_B2_c_166_n A1 0.0255035f $X=3.115 $Y=2.14 $X2=0 $Y2=0
cc_157 N_B2_c_158_n N_A1_c_268_n 0.00599726f $X=2.995 $Y=1.135 $X2=0 $Y2=0
cc_158 N_B2_c_159_n N_A1_c_268_n 0.0213844f $X=3.085 $Y=1.85 $X2=0 $Y2=0
cc_159 N_B2_c_165_n N_A1_c_268_n 0.00673801f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_160 N_B2_c_162_n N_Y_c_312_n 0.00149502f $X=1.445 $Y=2.015 $X2=0 $Y2=0
cc_161 N_B2_c_165_n N_Y_c_312_n 0.0167794f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_162 N_B2_c_162_n Y 0.0035198f $X=1.445 $Y=2.015 $X2=0 $Y2=0
cc_163 N_B2_c_165_n Y 0.0265538f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_164 N_B2_M1005_g Y 0.0029938f $X=1.355 $Y=2.66 $X2=0 $Y2=0
cc_165 N_B2_M1005_g N_Y_c_316_n 0.011743f $X=1.355 $Y=2.66 $X2=0 $Y2=0
cc_166 N_B2_c_162_n N_Y_c_316_n 8.14816e-19 $X=1.445 $Y=2.015 $X2=0 $Y2=0
cc_167 N_B2_c_165_n N_Y_c_316_n 0.0250978f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_168 N_B2_M1005_g N_VPWR_c_373_n 0.00161585f $X=1.355 $Y=2.66 $X2=0 $Y2=0
cc_169 B2 N_VPWR_c_374_n 0.0380147f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_170 N_B2_c_165_n N_VPWR_c_374_n 0.0259803f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_171 N_B2_M1005_g N_VPWR_c_375_n 0.00478016f $X=1.355 $Y=2.66 $X2=0 $Y2=0
cc_172 B2 N_VPWR_c_378_n 0.0124374f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_173 N_B2_M1005_g N_VPWR_c_372_n 0.0050291f $X=1.355 $Y=2.66 $X2=0 $Y2=0
cc_174 B2 N_VPWR_c_372_n 0.0114937f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_175 N_B2_M1007_g N_A_110_47#_c_418_n 0.0163562f $X=2.695 $Y=0.445 $X2=0 $Y2=0
cc_176 N_B2_c_158_n N_A_110_47#_c_418_n 0.00983882f $X=2.995 $Y=1.135 $X2=0
+ $Y2=0
cc_177 N_B2_M1007_g N_A_110_47#_c_419_n 0.00909898f $X=2.695 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_B2_M1007_g N_A_196_47#_c_462_n 4.20102e-19 $X=2.695 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_B2_M1007_g N_VGND_c_487_n 0.00585385f $X=2.695 $Y=0.445 $X2=0 $Y2=0
cc_180 N_B2_M1007_g N_VGND_c_488_n 0.0121599f $X=2.695 $Y=0.445 $X2=0 $Y2=0
cc_181 N_A2_c_216_n N_A1_c_264_n 0.00482804f $X=1.445 $Y=1.31 $X2=-0.19
+ $Y2=-0.245
cc_182 A2 N_A1_c_265_n 0.00600357f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_183 N_A2_c_220_n N_A1_c_265_n 0.0560509f $X=1.895 $Y=1.475 $X2=0 $Y2=0
cc_184 A2 N_A1_M1000_g 0.00167915f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A2_c_218_n N_A1_M1004_g 0.00539762f $X=1.445 $Y=0.85 $X2=0 $Y2=0
cc_186 A2 A1 0.0268889f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A2_M1008_g N_A1_c_268_n 0.0560509f $X=1.895 $Y=2.66 $X2=0 $Y2=0
cc_188 A2 N_A1_c_268_n 0.0108798f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A2_M1008_g Y 5.06755e-19 $X=1.895 $Y=2.66 $X2=0 $Y2=0
cc_190 N_A2_M1008_g N_VPWR_c_375_n 0.00478016f $X=1.895 $Y=2.66 $X2=0 $Y2=0
cc_191 N_A2_M1008_g N_VPWR_c_372_n 0.0094764f $X=1.895 $Y=2.66 $X2=0 $Y2=0
cc_192 N_A2_c_216_n N_A_110_47#_c_420_n 0.00652148f $X=1.445 $Y=1.31 $X2=0 $Y2=0
cc_193 N_A2_c_218_n N_A_110_47#_c_420_n 0.00594902f $X=1.445 $Y=0.85 $X2=0 $Y2=0
cc_194 A2 N_A_110_47#_c_420_n 2.29607e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A2_c_216_n N_A_110_47#_c_421_n 0.00396217f $X=1.445 $Y=1.31 $X2=0 $Y2=0
cc_196 N_A2_c_218_n N_A_110_47#_c_421_n 0.0018086f $X=1.445 $Y=0.85 $X2=0 $Y2=0
cc_197 A2 N_A_110_47#_c_421_n 0.04538f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A2_c_220_n N_A_110_47#_c_421_n 0.00998607f $X=1.895 $Y=1.475 $X2=0
+ $Y2=0
cc_199 N_A2_c_215_n N_A_196_47#_c_460_n 0.0106758f $X=1.335 $Y=0.775 $X2=0 $Y2=0
cc_200 N_A2_c_218_n N_A_196_47#_c_460_n 0.00324108f $X=1.445 $Y=0.85 $X2=0 $Y2=0
cc_201 N_A2_c_215_n N_A_196_47#_c_461_n 0.010222f $X=1.335 $Y=0.775 $X2=0 $Y2=0
cc_202 N_A2_c_215_n N_VGND_c_488_n 0.00701853f $X=1.335 $Y=0.775 $X2=0 $Y2=0
cc_203 N_A2_c_215_n N_VGND_c_489_n 0.00402633f $X=1.335 $Y=0.775 $X2=0 $Y2=0
cc_204 N_A2_c_215_n N_VGND_c_490_n 0.00716575f $X=1.335 $Y=0.775 $X2=0 $Y2=0
cc_205 N_A1_M1000_g N_VPWR_c_374_n 0.018075f $X=2.255 $Y=2.66 $X2=0 $Y2=0
cc_206 N_A1_M1000_g N_VPWR_c_375_n 0.00478016f $X=2.255 $Y=2.66 $X2=0 $Y2=0
cc_207 N_A1_M1000_g N_VPWR_c_372_n 0.00960321f $X=2.255 $Y=2.66 $X2=0 $Y2=0
cc_208 N_A1_c_264_n N_A_110_47#_c_418_n 3.15372e-19 $X=2.26 $Y=1.18 $X2=0 $Y2=0
cc_209 N_A1_M1004_g N_A_110_47#_c_418_n 0.0140282f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_210 A1 N_A_110_47#_c_418_n 0.0274915f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_211 N_A1_c_268_n N_A_110_47#_c_418_n 0.00696474f $X=2.545 $Y=1.585 $X2=0
+ $Y2=0
cc_212 N_A1_M1004_g N_A_196_47#_c_460_n 0.0107014f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_213 N_A1_M1004_g N_A_196_47#_c_462_n 0.0102469f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A1_M1004_g N_VGND_c_487_n 0.00402633f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A1_M1004_g N_VGND_c_488_n 0.00701853f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_216 N_A1_M1004_g N_VGND_c_490_n 0.00716575f $X=2.265 $Y=0.445 $X2=0 $Y2=0
cc_217 N_Y_c_311_n N_VPWR_M1001_d 7.02569e-19 $X=0.765 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_218 N_Y_c_339_n N_VPWR_M1001_d 0.00106976f $X=0.85 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_219 N_Y_c_311_n N_VPWR_c_373_n 0.00712262f $X=0.765 $Y=2.405 $X2=0 $Y2=0
cc_220 N_Y_c_313_n N_VPWR_c_373_n 0.0135201f $X=0.35 $Y=2.485 $X2=0 $Y2=0
cc_221 N_Y_c_339_n N_VPWR_c_373_n 0.00981978f $X=0.85 $Y=2.405 $X2=0 $Y2=0
cc_222 Y N_VPWR_c_373_n 0.00513141f $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_223 N_Y_c_316_n N_VPWR_c_373_n 6.38214e-19 $X=1.465 $Y=2.405 $X2=0 $Y2=0
cc_224 Y N_VPWR_c_374_n 3.37782e-19 $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_225 Y N_VPWR_c_374_n 3.18865e-19 $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_226 Y N_VPWR_c_375_n 0.0152302f $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_227 N_Y_c_313_n N_VPWR_c_377_n 0.0125145f $X=0.35 $Y=2.485 $X2=0 $Y2=0
cc_228 N_Y_c_311_n N_VPWR_c_372_n 0.00543208f $X=0.765 $Y=2.405 $X2=0 $Y2=0
cc_229 N_Y_c_313_n N_VPWR_c_372_n 0.00964185f $X=0.35 $Y=2.485 $X2=0 $Y2=0
cc_230 N_Y_c_339_n N_VPWR_c_372_n 6.13426e-19 $X=0.85 $Y=2.405 $X2=0 $Y2=0
cc_231 Y N_VPWR_c_372_n 0.0121804f $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_232 N_Y_c_316_n N_VPWR_c_372_n 0.0160356f $X=1.465 $Y=2.405 $X2=0 $Y2=0
cc_233 N_Y_c_316_n A_214_468# 0.00193007f $X=1.465 $Y=2.405 $X2=-0.19 $Y2=-0.245
cc_234 N_Y_c_306_n N_A_110_47#_c_417_n 0.013454f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_235 N_Y_c_306_n N_A_110_47#_c_424_n 0.0282568f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_236 N_Y_M1002_s N_VGND_c_488_n 0.00342001f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_237 N_Y_c_306_n N_VGND_c_488_n 0.0102927f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_238 N_Y_c_306_n N_VGND_c_489_n 0.0156583f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_239 N_A_110_47#_c_418_n N_A_196_47#_c_460_n 0.0491867f $X=2.77 $Y=0.96 $X2=0
+ $Y2=0
cc_240 N_A_110_47#_c_420_n N_A_196_47#_c_460_n 0.0249924f $X=1.465 $Y=0.957
+ $X2=0 $Y2=0
cc_241 N_A_110_47#_c_416_n N_A_196_47#_c_461_n 0.00335327f $X=0.63 $Y=0.87 $X2=0
+ $Y2=0
cc_242 N_A_110_47#_c_420_n N_A_196_47#_c_461_n 0.0223813f $X=1.465 $Y=0.957
+ $X2=0 $Y2=0
cc_243 N_A_110_47#_c_418_n N_A_196_47#_c_462_n 0.0223185f $X=2.77 $Y=0.96 $X2=0
+ $Y2=0
cc_244 N_A_110_47#_c_419_n N_A_196_47#_c_462_n 0.0183993f $X=2.91 $Y=0.445 $X2=0
+ $Y2=0
cc_245 N_A_110_47#_c_419_n N_VGND_c_487_n 0.0167415f $X=2.91 $Y=0.445 $X2=0
+ $Y2=0
cc_246 N_A_110_47#_M1002_d N_VGND_c_488_n 0.00226149f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_247 N_A_110_47#_M1007_d N_VGND_c_488_n 0.00216084f $X=2.77 $Y=0.235 $X2=0
+ $Y2=0
cc_248 N_A_110_47#_c_419_n N_VGND_c_488_n 0.0116369f $X=2.91 $Y=0.445 $X2=0
+ $Y2=0
cc_249 N_A_110_47#_c_424_n N_VGND_c_488_n 0.0109167f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_250 N_A_110_47#_c_424_n N_VGND_c_489_n 0.0138131f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_251 N_A_196_47#_c_460_n N_VGND_M1009_d 0.00954051f $X=2.315 $Y=0.615
+ $X2=-0.19 $Y2=-0.245
cc_252 N_A_196_47#_c_460_n N_VGND_c_487_n 0.00334901f $X=2.315 $Y=0.615 $X2=0
+ $Y2=0
cc_253 N_A_196_47#_c_462_n N_VGND_c_487_n 0.0139227f $X=2.48 $Y=0.445 $X2=0
+ $Y2=0
cc_254 N_A_196_47#_M1006_d N_VGND_c_488_n 0.00316506f $X=0.98 $Y=0.235 $X2=0
+ $Y2=0
cc_255 N_A_196_47#_M1004_d N_VGND_c_488_n 0.00299129f $X=2.34 $Y=0.235 $X2=0
+ $Y2=0
cc_256 N_A_196_47#_c_460_n N_VGND_c_488_n 0.0135672f $X=2.315 $Y=0.615 $X2=0
+ $Y2=0
cc_257 N_A_196_47#_c_461_n N_VGND_c_488_n 0.0104144f $X=1.12 $Y=0.445 $X2=0
+ $Y2=0
cc_258 N_A_196_47#_c_462_n N_VGND_c_488_n 0.0106039f $X=2.48 $Y=0.445 $X2=0
+ $Y2=0
cc_259 N_A_196_47#_c_460_n N_VGND_c_489_n 0.00334901f $X=2.315 $Y=0.615 $X2=0
+ $Y2=0
cc_260 N_A_196_47#_c_461_n N_VGND_c_489_n 0.013768f $X=1.12 $Y=0.445 $X2=0 $Y2=0
cc_261 N_A_196_47#_c_460_n N_VGND_c_490_n 0.0486499f $X=2.315 $Y=0.615 $X2=0
+ $Y2=0
