* File: sky130_fd_sc_lp__o221a_0.pex.spice
* Created: Wed Sep  2 10:18:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221A_0%C1 3 7 11 12 13 14 15 20
c39 20 0 1.77549e-19 $X=0.55 $Y=1.615
c40 7 0 1.3453e-19 $X=0.56 $Y=0.74
c41 3 0 7.20622e-20 $X=0.5 $Y=2.74
r42 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.55
+ $Y=1.615 $X2=0.55 $Y2=1.615
r43 14 15 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.665 $Y=1.665
+ $X2=0.665 $Y2=2.035
r44 14 21 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=0.665 $Y=1.665
+ $X2=0.665 $Y2=1.615
r45 13 21 9.21954 $w=3.98e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=1.295
+ $X2=0.665 $Y2=1.615
r46 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.55 $Y=1.955
+ $X2=0.55 $Y2=1.615
r47 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.955
+ $X2=0.55 $Y2=2.12
r48 10 20 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.45
+ $X2=0.55 $Y2=1.615
r49 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.56 $Y=0.74 $X2=0.56
+ $Y2=1.45
r50 3 12 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.5 $Y=2.74 $X2=0.5
+ $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%B1 3 7 10 12 13 14 15 16 20 22
c46 22 0 2.3898e-20 $X=1.15 $Y=1.545
c47 15 0 7.20622e-20 $X=1.2 $Y=1.665
c48 13 0 1.12826e-19 $X=1.01 $Y=1.21
r49 20 22 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.71
+ $X2=1.15 $Y2=1.545
r50 15 16 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=1.187 $Y=1.665
+ $X2=1.187 $Y2=2.035
r51 15 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.12
+ $Y=1.71 $X2=1.12 $Y2=1.71
r52 13 22 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.03 $Y=1.21
+ $X2=1.03 $Y2=1.545
r53 12 13 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.01 $Y=1.06
+ $X2=1.01 $Y2=1.21
r54 10 14 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=1.27 $Y=2.74
+ $X2=1.27 $Y2=2.215
r55 7 14 49.7341 $w=3.9e-07 $l=1.95e-07 $layer=POLY_cond $X=1.15 $Y=2.02
+ $X2=1.15 $Y2=2.215
r56 6 20 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=1.15 $Y=1.74 $X2=1.15
+ $Y2=1.71
r57 6 7 39.929 $w=3.9e-07 $l=2.8e-07 $layer=POLY_cond $X=1.15 $Y=1.74 $X2=1.15
+ $Y2=2.02
r58 3 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.99 $Y=0.74 $X2=0.99
+ $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%B2 1 3 8 12 15 16 17 18 20 27
c51 20 0 2.3898e-20 $X=2.16 $Y=2.035
c52 17 0 1.82648e-19 $X=1.72 $Y=2.17
r53 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.72
+ $Y=1.665 $X2=1.72 $Y2=1.665
r54 20 28 7.73933 $w=6.78e-07 $l=4.4e-07 $layer=LI1_cond $X=2.16 $Y=1.875
+ $X2=1.72 $Y2=1.875
r55 18 28 0.703576 $w=6.78e-07 $l=4e-08 $layer=LI1_cond $X=1.68 $Y=1.875
+ $X2=1.72 $Y2=1.875
r56 16 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.72 $Y=2.005
+ $X2=1.72 $Y2=1.665
r57 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.72 $Y=2.005
+ $X2=1.72 $Y2=2.17
r58 15 27 43.2685 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.72 $Y=1.5
+ $X2=1.72 $Y2=1.665
r59 10 12 111.27 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=1.42 $Y=1.135
+ $X2=1.637 $Y2=1.135
r60 8 17 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.63 $Y=2.74 $X2=1.63
+ $Y2=2.17
r61 4 12 0.660903 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.637 $Y=1.21
+ $X2=1.637 $Y2=1.135
r62 4 15 126.33 $w=1.65e-07 $l=2.9e-07 $layer=POLY_cond $X=1.637 $Y=1.21
+ $X2=1.637 $Y2=1.5
r63 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.42 $Y=1.06 $X2=1.42
+ $Y2=1.135
r64 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.42 $Y=1.06 $X2=1.42
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%A2 3 5 7 8 13
c45 13 0 1.2307e-19 $X=2.17 $Y=0.93
r46 11 13 14.0661 $w=2.57e-07 $l=7.5e-08 $layer=POLY_cond $X=2.095 $Y=0.93
+ $X2=2.17 $Y2=0.93
r47 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.095
+ $Y=0.93 $X2=2.095 $Y2=0.93
r48 5 13 45.0117 $w=2.57e-07 $l=3.11769e-07 $layer=POLY_cond $X=2.41 $Y=0.765
+ $X2=2.17 $Y2=0.93
r49 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.41 $Y=0.765 $X2=2.41
+ $Y2=0.445
r50 1 13 15.359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.095
+ $X2=2.17 $Y2=0.93
r51 1 3 843.5 $w=1.5e-07 $l=1.645e-06 $layer=POLY_cond $X=2.17 $Y=1.095 $X2=2.17
+ $Y2=2.74
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%A1 1 3 6 9 13 14 15 20
c47 13 0 1.2307e-19 $X=3.12 $Y=0.925
c48 1 0 9.54985e-20 $X=2.53 $Y=1.69
r49 20 22 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=2.867 $Y=1.035
+ $X2=2.867 $Y2=0.87
r50 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.875
+ $Y=1.035 $X2=2.875 $Y2=1.035
r51 14 15 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.027 $Y=1.295
+ $X2=3.027 $Y2=1.665
r52 14 21 6.54696 $w=4.73e-07 $l=2.6e-07 $layer=LI1_cond $X=3.027 $Y=1.295
+ $X2=3.027 $Y2=1.035
r53 13 21 2.76987 $w=4.73e-07 $l=1.1e-07 $layer=LI1_cond $X=3.027 $Y=0.925
+ $X2=3.027 $Y2=1.035
r54 9 22 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.84 $Y=0.445
+ $X2=2.84 $Y2=0.87
r55 5 20 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=2.867 $Y=1.042
+ $X2=2.867 $Y2=1.035
r56 5 6 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=2.867 $Y=1.042
+ $X2=2.867 $Y2=1.368
r57 1 6 80.8129 $w=2.01e-07 $l=4.09666e-07 $layer=POLY_cond $X=2.53 $Y=1.69
+ $X2=2.867 $Y2=1.529
r58 1 3 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.53 $Y=1.69 $X2=2.53
+ $Y2=2.74
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%A_32_484# 1 2 3 12 16 19 22 24 28 30 34 40
+ 42 43 47
c76 34 0 9.54985e-20 $X=3.1 $Y=2.095
c77 24 0 1.82648e-19 $X=1.735 $Y=2.47
r78 46 47 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.3 $Y=2.095
+ $X2=3.355 $Y2=2.095
r79 37 40 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.205 $Y=0.74
+ $X2=0.345 $Y2=0.74
r80 35 46 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=3.1 $Y=2.095 $X2=3.3
+ $Y2=2.095
r81 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.1
+ $Y=2.095 $X2=3.1 $Y2=2.095
r82 32 34 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.1 $Y=2.385 $X2=3.1
+ $Y2=2.095
r83 31 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=2.47
+ $X2=1.9 $Y2=2.47
r84 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.935 $Y=2.47
+ $X2=3.1 $Y2=2.385
r85 30 31 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.935 $Y=2.47
+ $X2=2.065 $Y2=2.47
r86 26 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.9 $Y=2.555 $X2=1.9
+ $Y2=2.47
r87 26 28 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.9 $Y=2.555 $X2=1.9
+ $Y2=2.56
r88 25 42 2.32734 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=0.38 $Y=2.47
+ $X2=0.247 $Y2=2.47
r89 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=2.47
+ $X2=1.9 $Y2=2.47
r90 24 25 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=1.735 $Y=2.47
+ $X2=0.38 $Y2=2.47
r91 20 42 4.10697 $w=2.22e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=2.555
+ $X2=0.247 $Y2=2.47
r92 20 22 0.434884 $w=2.63e-07 $l=1e-08 $layer=LI1_cond $X=0.247 $Y=2.555
+ $X2=0.247 $Y2=2.565
r93 19 42 4.10697 $w=2.22e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.205 $Y=2.385
+ $X2=0.247 $Y2=2.47
r94 18 37 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.205 $Y=0.905
+ $X2=0.205 $Y2=0.74
r95 18 19 91.1919 $w=1.78e-07 $l=1.48e-06 $layer=LI1_cond $X=0.205 $Y=0.905
+ $X2=0.205 $Y2=2.385
r96 14 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.93
+ $X2=3.355 $Y2=2.095
r97 14 16 761.457 $w=1.5e-07 $l=1.485e-06 $layer=POLY_cond $X=3.355 $Y=1.93
+ $X2=3.355 $Y2=0.445
r98 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=2.26 $X2=3.3
+ $Y2=2.095
r99 10 12 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.3 $Y=2.26 $X2=3.3
+ $Y2=2.74
r100 3 28 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=1.705
+ $Y=2.42 $X2=1.9 $Y2=2.56
r101 2 22 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=2.42 $X2=0.285 $Y2=2.565
r102 1 40 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.22
+ $Y=0.53 $X2=0.345 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%VPWR 1 2 9 18 19 24 30 34 40
r41 38 40 10.1341 $w=6.88e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=3.07
+ $X2=3.25 $Y2=3.07
r42 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 36 38 0.606706 $w=6.88e-07 $l=3.5e-08 $layer=LI1_cond $X=3.085 $Y=3.07
+ $X2=3.12 $Y2=3.07
r44 33 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 32 36 7.71384 $w=6.88e-07 $l=4.45e-07 $layer=LI1_cond $X=2.64 $Y=3.07
+ $X2=3.085 $Y2=3.07
r46 32 34 8.92072 $w=6.88e-07 $l=6e-08 $layer=LI1_cond $X=2.64 $Y=3.07 $X2=2.58
+ $Y2=3.07
r47 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 30 34 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.22 $Y=3.33
+ $X2=2.58 $Y2=3.33
r49 28 30 8.22735 $w=6.88e-07 $l=2e-08 $layer=LI1_cond $X=1.2 $Y=3.07 $X2=1.22
+ $Y2=3.07
r50 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 26 28 2.5135 $w=6.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.07
+ $X2=1.2 $Y2=3.07
r52 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 22 26 5.80705 $w=6.88e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=3.07
+ $X2=1.055 $Y2=3.07
r54 22 24 10.8275 $w=6.88e-07 $l=1.7e-07 $layer=LI1_cond $X=0.72 $Y=3.07
+ $X2=0.55 $Y2=3.07
r55 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 19 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 18 40 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=3.25
+ $Y2=3.33
r58 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r59 14 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 13 24 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=0.55 $Y2=3.33
r61 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 9 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 9 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33 $X2=1.2
+ $Y2=3.33
r64 2 36 300 $w=1.7e-07 $l=6.60908e-07 $layer=licon1_PDIFF $count=2 $X=2.605
+ $Y=2.42 $X2=3.085 $Y2=2.85
r65 1 26 300 $w=1.7e-07 $l=6.60908e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=2.42 $X2=1.055 $Y2=2.85
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%X 1 2 7 8 9 10 11 12 21
r13 12 34 4.98819 $w=3.33e-07 $l=1.45e-07 $layer=LI1_cond $X=3.587 $Y=2.775
+ $X2=3.587 $Y2=2.63
r14 11 34 8.10312 $w=3.18e-07 $l=2.25e-07 $layer=LI1_cond $X=3.595 $Y=2.405
+ $X2=3.595 $Y2=2.63
r15 10 11 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.595 $Y=2.035
+ $X2=3.595 $Y2=2.405
r16 9 10 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.595 $Y=1.665
+ $X2=3.595 $Y2=2.035
r17 8 9 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.595 $Y=1.295
+ $X2=3.595 $Y2=1.665
r18 7 8 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.595 $Y=0.925
+ $X2=3.595 $Y2=1.295
r19 7 21 17.2866 $w=3.18e-07 $l=4.8e-07 $layer=LI1_cond $X=3.595 $Y=0.925
+ $X2=3.595 $Y2=0.445
r20 2 12 600 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=2.42 $X2=3.515 $Y2=2.795
r21 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.235 $X2=3.57 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%A_127_106# 1 2 9 11 12 15
c24 11 0 1.12826e-19 $X=1.54 $Y=0.347
c25 9 0 1.77549e-19 $X=0.775 $Y=0.74
r26 13 15 16.6364 $w=1.98e-07 $l=3e-07 $layer=LI1_cond $X=1.64 $Y=0.44 $X2=1.64
+ $Y2=0.74
r27 11 13 6.82996 $w=1.85e-07 $l=1.38924e-07 $layer=LI1_cond $X=1.54 $Y=0.347
+ $X2=1.64 $Y2=0.44
r28 11 12 40.1671 $w=1.83e-07 $l=6.7e-07 $layer=LI1_cond $X=1.54 $Y=0.347
+ $X2=0.87 $Y2=0.347
r29 7 12 6.88292 $w=1.85e-07 $l=1.49432e-07 $layer=LI1_cond $X=0.76 $Y=0.44
+ $X2=0.87 $Y2=0.347
r30 7 9 15.7151 $w=2.18e-07 $l=3e-07 $layer=LI1_cond $X=0.76 $Y=0.44 $X2=0.76
+ $Y2=0.74
r31 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.53 $X2=1.635 $Y2=0.74
r32 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.635
+ $Y=0.53 $X2=0.775 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%A_213_106# 1 2 9 11 12 14 18
c42 12 0 1.3453e-19 $X=1.37 $Y=1.28
r43 15 18 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.535 $Y=0.445
+ $X2=2.625 $Y2=0.445
r44 13 15 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=0.61
+ $X2=2.535 $Y2=0.445
r45 13 14 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.535 $Y=0.61
+ $X2=2.535 $Y2=1.195
r46 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.45 $Y=1.28
+ $X2=2.535 $Y2=1.195
r47 11 12 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=2.45 $Y=1.28
+ $X2=1.37 $Y2=1.28
r48 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.205 $Y=1.195
+ $X2=1.37 $Y2=1.28
r49 7 9 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.205 $Y=1.195
+ $X2=1.205 $Y2=0.74
r50 2 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.625 $Y2=0.445
r51 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.53 $X2=1.205 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_0%VGND 1 2 9 13 15 17 25 32 33 36 39
r46 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r49 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.1
+ $Y2=0
r51 30 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.6
+ $Y2=0
r52 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r53 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r54 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r55 26 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.155
+ $Y2=0
r56 26 28 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.64
+ $Y2=0
r57 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=3.1
+ $Y2=0
r58 25 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=2.64
+ $Y2=0
r59 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 20 24 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r61 19 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r62 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 17 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.155
+ $Y2=0
r64 17 23 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=1.68
+ $Y2=0
r65 15 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r66 15 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r67 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0
r68 11 13 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0.445
r69 7 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.155 $Y2=0
r70 7 9 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.155 $Y2=0.43
r71 2 13 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.445
r72 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.235 $X2=2.195 $Y2=0.43
.ends

