* File: sky130_fd_sc_lp__o2111ai_m.pex.spice
* Created: Wed Sep  2 10:13:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111AI_M%D1 2 3 4 7 9 11 14 17 19 20 21 22 28
c48 7 0 1.8461e-19 $X=0.85 $Y=2.885
r49 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=0.945 $X2=0.58 $Y2=0.945
r50 21 22 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.65 $Y=1.665
+ $X2=0.65 $Y2=2.035
r51 20 21 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.65 $Y=1.295
+ $X2=0.65 $Y2=1.665
r52 20 29 13.0115 $w=3.08e-07 $l=3.5e-07 $layer=LI1_cond $X=0.65 $Y=1.295
+ $X2=0.65 $Y2=0.945
r53 19 29 0.743512 $w=3.08e-07 $l=2e-08 $layer=LI1_cond $X=0.65 $Y=0.925
+ $X2=0.65 $Y2=0.945
r54 15 17 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.67 $Y=2.155
+ $X2=0.85 $Y2=2.155
r55 13 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.58 $Y=1.285
+ $X2=0.58 $Y2=0.945
r56 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.285
+ $X2=0.58 $Y2=1.45
r57 12 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.58 $Y=0.93
+ $X2=0.58 $Y2=0.945
r58 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.99 $Y=0.78 $X2=0.99
+ $Y2=0.46
r59 5 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.85 $Y=2.23 $X2=0.85
+ $Y2=2.155
r60 5 7 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.85 $Y=2.23 $X2=0.85
+ $Y2=2.885
r61 4 12 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.745 $Y=0.855
+ $X2=0.58 $Y2=0.93
r62 3 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.915 $Y=0.855
+ $X2=0.99 $Y2=0.78
r63 3 4 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.915 $Y=0.855
+ $X2=0.745 $Y2=0.855
r64 2 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.67 $Y=2.08 $X2=0.67
+ $Y2=2.155
r65 2 14 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.67 $Y=2.08 $X2=0.67
+ $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_M%C1 5 8 12 14 15 16 17 18 19 20 21 28
c57 16 0 2.18351e-19 $X=1.245 $Y=2.56
r58 20 21 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.665
+ $X2=1.175 $Y2=2.035
r59 19 20 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.295
+ $X2=1.175 $Y2=1.665
r60 19 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.335 $X2=1.15 $Y2=1.335
r61 18 19 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=0.925
+ $X2=1.175 $Y2=1.295
r62 17 18 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=0.555
+ $X2=1.175 $Y2=0.925
r63 15 16 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.245 $Y=2.41
+ $X2=1.245 $Y2=2.56
r64 14 15 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.21 $Y=1.84
+ $X2=1.21 $Y2=2.41
r65 13 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.15 $Y=1.675
+ $X2=1.15 $Y2=1.335
r66 13 14 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.675
+ $X2=1.15 $Y2=1.84
r67 12 28 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=1.15 $Y=1.29
+ $X2=1.15 $Y2=1.335
r68 11 12 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.205 $Y=1.14
+ $X2=1.205 $Y2=1.29
r69 8 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.35 $Y=0.46 $X2=1.35
+ $Y2=1.14
r70 5 16 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.28 $Y=2.885
+ $X2=1.28 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_M%B1 3 7 11 12 13 14 15 20
c44 20 0 1.36011e-19 $X=1.69 $Y=1.695
c45 7 0 1.01012e-19 $X=1.71 $Y=2.885
r46 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=1.665
+ $X2=1.69 $Y2=2.035
r47 14 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.695 $X2=1.69 $Y2=1.695
r48 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=1.295
+ $X2=1.69 $Y2=1.665
r49 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.69 $Y=2.035
+ $X2=1.69 $Y2=1.695
r50 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=2.035
+ $X2=1.69 $Y2=2.2
r51 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.53
+ $X2=1.69 $Y2=1.695
r52 7 12 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=1.71 $Y=2.885
+ $X2=1.71 $Y2=2.2
r53 3 10 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.71 $Y=0.46 $X2=1.71
+ $Y2=1.53
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_M%A2 3 7 11 12 13 14 15 20
c42 12 0 1.32761e-19 $X=2.23 $Y=1.88
r43 14 15 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=2.035
r44 13 14 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=1.295
+ $X2=2.195 $Y2=1.665
r45 13 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23
+ $Y=1.375 $X2=2.23 $Y2=1.375
r46 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.23 $Y=1.715
+ $X2=2.23 $Y2=1.375
r47 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.715
+ $X2=2.23 $Y2=1.88
r48 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.21
+ $X2=2.23 $Y2=1.375
r49 7 12 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=2.14 $Y=2.885
+ $X2=2.14 $Y2=1.88
r50 3 10 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.14 $Y=0.46 $X2=2.14
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_M%A1 3 7 14 18 21 22 23 24 25 31
c36 18 0 2.58839e-20 $X=2.71 $Y=0.895
r37 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.8
+ $Y=1.765 $X2=2.8 $Y2=1.765
r38 24 25 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.72 $Y=2.035
+ $X2=2.72 $Y2=2.405
r39 24 32 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.72 $Y=2.035
+ $X2=2.72 $Y2=1.765
r40 23 32 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.72 $Y=1.665 $X2=2.72
+ $Y2=1.765
r41 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.72 $Y=1.295
+ $X2=2.72 $Y2=1.665
r42 21 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.8 $Y=1.6 $X2=2.8
+ $Y2=1.765
r43 16 18 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.57 $Y=0.895
+ $X2=2.71 $Y2=0.895
r44 14 31 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.8 $Y=2.12 $X2=2.8
+ $Y2=1.765
r45 11 14 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.5 $Y=2.195 $X2=2.8
+ $Y2=2.195
r46 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.71 $Y=0.97 $X2=2.71
+ $Y2=0.895
r47 9 21 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.71 $Y=0.97 $X2=2.71
+ $Y2=1.6
r48 5 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.57 $Y=0.82 $X2=2.57
+ $Y2=0.895
r49 5 7 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.57 $Y=0.82 $X2=2.57
+ $Y2=0.46
r50 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.5 $Y=2.27 $X2=2.5
+ $Y2=2.195
r51 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.5 $Y=2.27 $X2=2.5
+ $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_M%VPWR 1 2 3 10 12 16 20 23 24 25 31 37 38
+ 44
c44 38 0 2.66457e-20 $X=3.12 $Y=3.33
c45 23 0 1.91706e-19 $X=1.39 $Y=3.33
r46 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 38 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 35 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=2.715 $Y2=3.33
r51 35 37 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 34 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=3.33
+ $X2=2.715 $Y2=3.33
r55 31 33 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.55 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 30 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 27 41 3.49867 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r59 27 29 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 25 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 25 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 23 29 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.39 $Y=3.33 $X2=1.2
+ $Y2=3.33
r63 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.495 $Y2=3.33
r64 22 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.6 $Y=3.33 $X2=2.16
+ $Y2=3.33
r65 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.6 $Y=3.33
+ $X2=1.495 $Y2=3.33
r66 18 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=3.245
+ $X2=2.715 $Y2=3.33
r67 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.715 $Y=3.245
+ $X2=2.715 $Y2=2.95
r68 14 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.495 $Y=3.245
+ $X2=1.495 $Y2=3.33
r69 14 16 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.495 $Y=3.245
+ $X2=1.495 $Y2=2.97
r70 10 41 3.34522 $w=1.9e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.227 $Y2=3.33
r71 10 12 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.36 $Y2=2.95
r72 3 20 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=2.675 $X2=2.715 $Y2=2.95
r73 2 16 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.355
+ $Y=2.675 $X2=1.495 $Y2=2.97
r74 1 12 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=2.675 $X2=0.37 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_M%Y 1 2 3 11 15 17 18 20 21 28 31
c54 28 0 1.8461e-19 $X=1.82 $Y=2.472
c55 21 0 1.32761e-19 $X=2.16 $Y=2.405
c56 18 0 1.01012e-19 $X=0.72 $Y=2.405
r57 39 41 7.7801 $w=5.33e-07 $l=3.48e-07 $layer=LI1_cond $X=0.902 $Y=2.472
+ $X2=0.902 $Y2=2.82
r58 29 39 4.03697 $w=3.05e-07 $l=2.68e-07 $layer=LI1_cond $X=1.17 $Y=2.472
+ $X2=0.902 $Y2=2.472
r59 29 31 1.13355 $w=3.03e-07 $l=3e-08 $layer=LI1_cond $X=1.17 $Y=2.472 $X2=1.2
+ $Y2=2.472
r60 28 48 8.89415 $w=4.23e-07 $l=3.28e-07 $layer=LI1_cond $X=2.032 $Y=2.472
+ $X2=2.032 $Y2=2.8
r61 21 28 1.81679 $w=4.23e-07 $l=6.7e-08 $layer=LI1_cond $X=2.032 $Y=2.405
+ $X2=2.032 $Y2=2.472
r62 20 28 5.2899 $w=3.03e-07 $l=1.4e-07 $layer=LI1_cond $X=1.68 $Y=2.472
+ $X2=1.82 $Y2=2.472
r63 18 39 1.49789 $w=5.33e-07 $l=6.7e-08 $layer=LI1_cond $X=0.902 $Y=2.405
+ $X2=0.902 $Y2=2.472
r64 18 20 17.1166 $w=3.03e-07 $l=4.53e-07 $layer=LI1_cond $X=1.227 $Y=2.472
+ $X2=1.68 $Y2=2.472
r65 18 31 1.0202 $w=3.03e-07 $l=2.7e-08 $layer=LI1_cond $X=1.227 $Y=2.472
+ $X2=1.2 $Y2=2.472
r66 17 18 12.2861 $w=3.38e-07 $l=3.2e-07 $layer=LI1_cond $X=0.315 $Y=2.405
+ $X2=0.635 $Y2=2.405
r67 12 15 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.23 $Y=0.435
+ $X2=0.64 $Y2=0.435
r68 11 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.23 $Y=2.32
+ $X2=0.315 $Y2=2.405
r69 10 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.23 $Y=0.6 $X2=0.23
+ $Y2=0.435
r70 10 11 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=0.23 $Y=0.6
+ $X2=0.23 $Y2=2.32
r71 3 48 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.785
+ $Y=2.675 $X2=1.925 $Y2=2.8
r72 2 41 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.925
+ $Y=2.675 $X2=1.065 $Y2=2.82
r73 1 15 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.515
+ $Y=0.25 $X2=0.64 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_M%A_357_50# 1 2 9 11 12 15
c26 12 0 1.36011e-19 $X=2.03 $Y=0.825
r27 13 15 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.785 $Y=0.74
+ $X2=2.785 $Y2=0.525
r28 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.68 $Y=0.825
+ $X2=2.785 $Y2=0.74
r29 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.68 $Y=0.825
+ $X2=2.03 $Y2=0.825
r30 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.925 $Y=0.74
+ $X2=2.03 $Y2=0.825
r31 7 9 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.925 $Y=0.74
+ $X2=1.925 $Y2=0.525
r32 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.25 $X2=2.785 $Y2=0.525
r33 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.785
+ $Y=0.25 $X2=1.925 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__O2111AI_M%VGND 1 6 9 10 11 21 22
c32 22 0 2.58839e-20 $X=3.12 $Y=0
r33 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r34 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r35 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r36 14 18 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r37 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r38 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r39 11 15 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r40 9 18 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.16
+ $Y2=0
r41 9 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.355
+ $Y2=0
r42 8 21 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=3.12
+ $Y2=0
r43 8 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.355
+ $Y2=0
r44 4 10 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=0.085
+ $X2=2.355 $Y2=0
r45 4 6 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=2.355 $Y=0.085
+ $X2=2.355 $Y2=0.395
r46 1 6 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.25 $X2=2.355 $Y2=0.395
.ends

