* NGSPICE file created from sky130_fd_sc_lp__o31a_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 VGND A2 a_275_49# VNB nshort w=840000u l=150000u
+  ad=8.82e+11p pd=5.46e+06u as=4.914e+11p ps=4.53e+06u
M1001 a_86_23# A3 a_367_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.914e+11p pd=3.3e+06u as=3.654e+11p ps=3.1e+06u
M1002 a_275_49# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_86_23# X VPB phighvt w=1.26e+06u l=150000u
+  ad=1.1466e+12p pd=6.86e+06u as=3.339e+11p ps=3.05e+06u
M1004 a_275_49# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_86_23# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1006 VPWR B1 a_86_23# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_275_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.906e+11p pd=3.14e+06u as=0p ps=0u
M1008 a_86_23# B1 a_275_49# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1009 a_367_367# A2 a_275_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

