* File: sky130_fd_sc_lp__a221o_4.pex.spice
* Created: Wed Sep  2 09:21:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221O_4%A_83_21# 1 2 3 4 5 18 22 26 30 34 38 42 46
+ 48 56 58 60 63 64 66 70 72 76 78 82 90 99
c169 99 0 9.42274e-20 $X=1.78 $Y=1.49
c170 56 0 1.79433e-19 $X=4.125 $Y=1.782
r171 96 97 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.92 $Y=1.49
+ $X2=1.35 $Y2=1.49
r172 82 85 6.12235 $w=3.18e-07 $l=1.7e-07 $layer=LI1_cond $X=3.37 $Y=0.34
+ $X2=3.37 $Y2=0.51
r173 78 80 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.935 $Y=1.492
+ $X2=1.935 $Y2=1.782
r174 74 92 3.47416 $w=2.6e-07 $l=1.35e-07 $layer=LI1_cond $X=5.235 $Y=0.385
+ $X2=5.1 $Y2=0.385
r175 74 76 31.9138 $w=2.58e-07 $l=7.2e-07 $layer=LI1_cond $X=5.235 $Y=0.385
+ $X2=5.955 $Y2=0.385
r176 72 92 3.34549 $w=2.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.1 $Y=0.515 $X2=5.1
+ $Y2=0.385
r177 72 73 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.1 $Y=0.515
+ $X2=5.1 $Y2=0.855
r178 68 70 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.665 $Y=1.875
+ $X2=4.665 $Y2=2.14
r179 67 89 2.0246 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.365 $Y=0.94
+ $X2=4.245 $Y2=0.94
r180 66 73 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.965 $Y=0.94
+ $X2=5.1 $Y2=0.855
r181 66 67 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.965 $Y=0.94
+ $X2=4.365 $Y2=0.94
r182 65 90 4.98297 $w=1.77e-07 $l=8.89101e-08 $layer=LI1_cond $X=4.295 $Y=1.79
+ $X2=4.21 $Y2=1.782
r183 64 68 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.5 $Y=1.79
+ $X2=4.665 $Y2=1.875
r184 64 65 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.5 $Y=1.79
+ $X2=4.295 $Y2=1.79
r185 63 90 1.49848 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=4.21 $Y=1.69
+ $X2=4.21 $Y2=1.782
r186 62 89 4.40882 $w=2.05e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.21 $Y=1.025
+ $X2=4.245 $Y2=0.94
r187 62 63 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.21 $Y=1.025
+ $X2=4.21 $Y2=1.69
r188 61 89 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=0.855
+ $X2=4.245 $Y2=0.94
r189 60 88 2.93484 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=0.425
+ $X2=4.245 $Y2=0.34
r190 60 61 20.6479 $w=2.38e-07 $l=4.3e-07 $layer=LI1_cond $X=4.245 $Y=0.425
+ $X2=4.245 $Y2=0.855
r191 59 82 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.53 $Y=0.34
+ $X2=3.37 $Y2=0.34
r192 58 88 4.1433 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.125 $Y=0.34
+ $X2=4.245 $Y2=0.34
r193 58 59 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.125 $Y=0.34
+ $X2=3.53 $Y2=0.34
r194 57 80 0.22998 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=1.782
+ $X2=1.935 $Y2=1.782
r195 56 90 4.98297 $w=1.77e-07 $l=8.5e-08 $layer=LI1_cond $X=4.125 $Y=1.782
+ $X2=4.21 $Y2=1.782
r196 56 57 126.197 $w=1.83e-07 $l=2.105e-06 $layer=LI1_cond $X=4.125 $Y=1.782
+ $X2=2.02 $Y2=1.782
r197 55 99 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.69 $Y=1.49 $X2=1.78
+ $Y2=1.49
r198 55 97 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.69 $Y=1.49
+ $X2=1.35 $Y2=1.49
r199 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.49 $X2=1.69 $Y2=1.49
r200 51 96 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.67 $Y=1.49
+ $X2=0.92 $Y2=1.49
r201 51 93 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.67 $Y=1.49
+ $X2=0.49 $Y2=1.49
r202 50 54 61.1499 $w=1.83e-07 $l=1.02e-06 $layer=LI1_cond $X=0.67 $Y=1.492
+ $X2=1.69 $Y2=1.492
r203 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.67
+ $Y=1.49 $X2=0.67 $Y2=1.49
r204 48 78 0.22998 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.85 $Y=1.492
+ $X2=1.935 $Y2=1.492
r205 48 54 9.59214 $w=1.83e-07 $l=1.6e-07 $layer=LI1_cond $X=1.85 $Y=1.492
+ $X2=1.69 $Y2=1.492
r206 44 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.655
+ $X2=1.78 $Y2=1.49
r207 44 46 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.78 $Y=1.655
+ $X2=1.78 $Y2=2.465
r208 40 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=1.49
r209 40 42 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=0.655
r210 36 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.655
+ $X2=1.35 $Y2=1.49
r211 36 38 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.35 $Y=1.655
+ $X2=1.35 $Y2=2.465
r212 32 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=1.49
r213 32 34 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=0.655
r214 28 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.655
+ $X2=0.92 $Y2=1.49
r215 28 30 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.92 $Y=1.655
+ $X2=0.92 $Y2=2.465
r216 24 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.325
+ $X2=0.92 $Y2=1.49
r217 24 26 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.92 $Y=1.325
+ $X2=0.92 $Y2=0.655
r218 20 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.655
+ $X2=0.49 $Y2=1.49
r219 20 22 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.49 $Y=1.655
+ $X2=0.49 $Y2=2.465
r220 16 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.49
r221 16 18 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=0.655
r222 5 70 600 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=4.525
+ $Y=1.835 $X2=4.665 $Y2=2.14
r223 4 76 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.235 $X2=5.955 $Y2=0.4
r224 3 92 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.955
+ $Y=0.235 $X2=5.095 $Y2=0.42
r225 2 88 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.095
+ $Y=0.235 $X2=4.235 $Y2=0.42
r226 1 85 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.235 $X2=3.375 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%A2 1 3 6 8 10 13 15 16 23
c47 23 0 1.27343e-19 $X=2.64 $Y=1.352
c48 16 0 9.42274e-20 $X=3.12 $Y=1.295
r49 21 23 2.91239 $w=3.31e-07 $l=2e-08 $layer=POLY_cond $X=2.62 $Y=1.352
+ $X2=2.64 $Y2=1.352
r50 15 16 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.62 $Y=1.35 $X2=3.12
+ $Y2=1.35
r51 15 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.62
+ $Y=1.35 $X2=2.62 $Y2=1.35
r52 11 23 21.295 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=2.64 $Y=1.52
+ $X2=2.64 $Y2=1.352
r53 11 13 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=2.64 $Y=1.52
+ $X2=2.64 $Y2=2.465
r54 8 23 21.295 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=2.64 $Y=1.185
+ $X2=2.64 $Y2=1.352
r55 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.64 $Y=1.185
+ $X2=2.64 $Y2=0.655
r56 4 21 59.7039 $w=3.31e-07 $l=4.1e-07 $layer=POLY_cond $X=2.21 $Y=1.352
+ $X2=2.62 $Y2=1.352
r57 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.21 $Y=1.515 $X2=2.21
+ $Y2=2.465
r58 1 4 21.295 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=2.21 $Y=1.185 $X2=2.21
+ $Y2=1.352
r59 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.21 $Y=1.185 $X2=2.21
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%A1 3 7 9 11 12 14 15 23 24
c46 23 0 1.27343e-19 $X=3.835 $Y=1.35
r47 22 24 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.835 $Y=1.35
+ $X2=4.02 $Y2=1.35
r48 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.835
+ $Y=1.35 $X2=3.835 $Y2=1.35
r49 20 22 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=3.59 $Y=1.35
+ $X2=3.835 $Y2=1.35
r50 19 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.5 $Y=1.35 $X2=3.59
+ $Y2=1.35
r51 17 19 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.07 $Y=1.35 $X2=3.5
+ $Y2=1.35
r52 15 23 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=3.6 $Y=1.35
+ $X2=3.835 $Y2=1.35
r53 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.02 $Y=1.185
+ $X2=4.02 $Y2=1.35
r54 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.02 $Y=1.185
+ $X2=4.02 $Y2=0.655
r55 9 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.59 $Y=1.185
+ $X2=3.59 $Y2=1.35
r56 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.59 $Y=1.185
+ $X2=3.59 $Y2=0.655
r57 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.5 $Y=1.515 $X2=3.5
+ $Y2=1.35
r58 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.5 $Y=1.515 $X2=3.5
+ $Y2=2.465
r59 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.515
+ $X2=3.07 $Y2=1.35
r60 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.07 $Y=1.515 $X2=3.07
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%C1 1 3 6 8 10 13 15 16 24
r48 22 24 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=4.72 $Y=1.36
+ $X2=4.88 $Y2=1.36
r49 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.72
+ $Y=1.36 $X2=4.72 $Y2=1.36
r50 19 22 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=4.45 $Y=1.36
+ $X2=4.72 $Y2=1.36
r51 16 23 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=5.04 $Y=1.36
+ $X2=4.72 $Y2=1.36
r52 15 23 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.56 $Y=1.36 $X2=4.72
+ $Y2=1.36
r53 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.88 $Y=1.525
+ $X2=4.88 $Y2=1.36
r54 11 13 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.88 $Y=1.525 $X2=4.88
+ $Y2=2.465
r55 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.88 $Y=1.195
+ $X2=4.88 $Y2=1.36
r56 8 10 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=4.88 $Y=1.195 $X2=4.88
+ $Y2=0.655
r57 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.45 $Y=1.525
+ $X2=4.45 $Y2=1.36
r58 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.45 $Y=1.525 $X2=4.45
+ $Y2=2.465
r59 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.45 $Y=1.195
+ $X2=4.45 $Y2=1.36
r60 1 3 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=4.45 $Y=1.195 $X2=4.45
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%B1 1 3 6 8 10 13 15 16 24
c50 24 0 1.79196e-19 $X=5.74 $Y=1.36
r51 22 24 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.72 $Y=1.36 $X2=5.74
+ $Y2=1.36
r52 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.72
+ $Y=1.36 $X2=5.72 $Y2=1.36
r53 19 22 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=5.31 $Y=1.36
+ $X2=5.72 $Y2=1.36
r54 16 23 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6 $Y=1.36 $X2=5.72
+ $Y2=1.36
r55 15 23 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=5.52 $Y=1.36 $X2=5.72
+ $Y2=1.36
r56 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.74 $Y=1.525
+ $X2=5.74 $Y2=1.36
r57 11 13 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=5.74 $Y=1.525 $X2=5.74
+ $Y2=2.465
r58 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.74 $Y=1.195
+ $X2=5.74 $Y2=1.36
r59 8 10 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.74 $Y=1.195 $X2=5.74
+ $Y2=0.655
r60 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.525
+ $X2=5.31 $Y2=1.36
r61 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=5.31 $Y=1.525 $X2=5.31
+ $Y2=2.465
r62 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.195
+ $X2=5.31 $Y2=1.36
r63 1 3 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=5.31 $Y=1.195 $X2=5.31
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%B2 3 7 11 15 17 18 25 29 37
r46 29 37 0.884058 $w=3.45e-07 $l=2.5e-08 $layer=LI1_cond $X=6.985 $Y=1.577
+ $X2=6.96 $Y2=1.577
r47 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.135
+ $Y=1.49 $X2=7.135 $Y2=1.49
r48 25 27 2.12023 $w=3.41e-07 $l=1.5e-08 $layer=POLY_cond $X=7.12 $Y=1.5
+ $X2=7.135 $Y2=1.5
r49 24 25 60.7801 $w=3.41e-07 $l=4.3e-07 $layer=POLY_cond $X=6.69 $Y=1.5
+ $X2=7.12 $Y2=1.5
r50 23 24 12.7214 $w=3.41e-07 $l=9e-08 $layer=POLY_cond $X=6.6 $Y=1.5 $X2=6.69
+ $Y2=1.5
r51 22 23 60.7801 $w=3.41e-07 $l=4.3e-07 $layer=POLY_cond $X=6.17 $Y=1.5 $X2=6.6
+ $Y2=1.5
r52 18 28 10.1883 $w=3.43e-07 $l=3.05e-07 $layer=LI1_cond $X=7.44 $Y=1.577
+ $X2=7.135 $Y2=1.577
r53 17 37 1.07331 $w=3.41e-07 $l=3e-08 $layer=LI1_cond $X=6.93 $Y=1.577 $X2=6.96
+ $Y2=1.577
r54 17 28 4.0085 $w=3.43e-07 $l=1.2e-07 $layer=LI1_cond $X=7.015 $Y=1.577
+ $X2=7.135 $Y2=1.577
r55 17 29 1.00212 $w=3.43e-07 $l=3e-08 $layer=LI1_cond $X=7.015 $Y=1.577
+ $X2=6.985 $Y2=1.577
r56 13 25 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=7.12 $Y=1.325
+ $X2=7.12 $Y2=1.5
r57 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.12 $Y=1.325
+ $X2=7.12 $Y2=0.665
r58 9 24 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.69 $Y=1.325
+ $X2=6.69 $Y2=1.5
r59 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.69 $Y=1.325
+ $X2=6.69 $Y2=0.665
r60 5 23 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.6 $Y=1.675 $X2=6.6
+ $Y2=1.5
r61 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.6 $Y=1.675 $X2=6.6
+ $Y2=2.465
r62 1 22 22.0049 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.17 $Y=1.675
+ $X2=6.17 $Y2=1.5
r63 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.17 $Y=1.675 $X2=6.17
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%VPWR 1 2 3 4 5 16 18 24 30 36 38 42 45 46 47
+ 48 49 51 68 69 75 78
r109 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r110 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r111 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r112 68 69 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r113 66 69 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 65 68 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=7.44 $Y2=3.33
r115 65 66 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r116 63 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=3.33
+ $X2=3.715 $Y2=3.33
r117 63 65 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.88 $Y=3.33 $X2=4.08
+ $Y2=3.33
r118 62 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r119 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r121 59 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 56 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.135 $Y2=3.33
r124 56 58 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.68 $Y2=3.33
r125 55 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 55 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r127 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r128 52 72 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r129 52 54 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 51 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.135 $Y2=3.33
r131 51 54 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.72 $Y2=3.33
r132 49 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 49 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r134 47 61 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=3.33 $X2=2.64
+ $Y2=3.33
r135 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=2.855 $Y2=3.33
r136 45 58 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=1.68 $Y2=3.33
r137 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=1.995 $Y2=3.33
r138 44 61 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r139 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=1.995 $Y2=3.33
r140 40 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=3.245
+ $X2=3.715 $Y2=3.33
r141 40 42 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=3.715 $Y=3.245
+ $X2=3.715 $Y2=2.47
r142 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=2.855 $Y2=3.33
r143 38 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=3.33
+ $X2=3.715 $Y2=3.33
r144 38 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.55 $Y=3.33
+ $X2=3.02 $Y2=3.33
r145 34 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=3.245
+ $X2=2.855 $Y2=3.33
r146 34 36 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=2.855 $Y=3.245
+ $X2=2.855 $Y2=2.48
r147 30 33 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=1.995 $Y=2.13
+ $X2=1.995 $Y2=2.95
r148 28 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=3.245
+ $X2=1.995 $Y2=3.33
r149 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.995 $Y=3.245
+ $X2=1.995 $Y2=2.95
r150 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=2.18
+ $X2=1.135 $Y2=2.95
r151 22 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=3.33
r152 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=2.95
r153 18 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.275 $Y=2.18
+ $X2=0.275 $Y2=2.95
r154 16 72 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r155 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.95
r156 5 42 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=3.575
+ $Y=1.835 $X2=3.715 $Y2=2.47
r157 4 36 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=2.715
+ $Y=1.835 $X2=2.855 $Y2=2.48
r158 3 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=1.995 $Y2=2.95
r159 3 30 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=1.995 $Y2=2.13
r160 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.95
r161 2 24 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.18
r162 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.95
r163 1 18 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%X 1 2 3 4 13 15 16 19 23 27 29 33 37 42 43
+ 44 45 49 51
r56 49 51 3.32928 $w=2.23e-07 $l=6.5e-08 $layer=LI1_cond $X=0.222 $Y=1.23
+ $X2=0.222 $Y2=1.295
r57 44 49 3.00067 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.222 $Y=1.145
+ $X2=0.222 $Y2=1.23
r58 44 45 18.4391 $w=2.23e-07 $l=3.6e-07 $layer=LI1_cond $X=0.222 $Y=1.305
+ $X2=0.222 $Y2=1.665
r59 44 51 0.512197 $w=2.23e-07 $l=1e-08 $layer=LI1_cond $X=0.222 $Y=1.305
+ $X2=0.222 $Y2=1.295
r60 41 45 4.60977 $w=2.23e-07 $l=9e-08 $layer=LI1_cond $X=0.222 $Y=1.755
+ $X2=0.222 $Y2=1.665
r61 37 39 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.565 $Y=1.98
+ $X2=1.565 $Y2=2.91
r62 35 37 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.565 $Y=1.925
+ $X2=1.565 $Y2=1.98
r63 31 33 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=1.565 $Y=1.045
+ $X2=1.565 $Y2=0.42
r64 30 42 5.465 $w=1.77e-07 $l=9.5e-08 $layer=LI1_cond $X=0.8 $Y=1.137 $X2=0.705
+ $Y2=1.137
r65 29 31 6.81807 $w=1.85e-07 $l=1.33285e-07 $layer=LI1_cond $X=1.47 $Y=1.137
+ $X2=1.565 $Y2=1.045
r66 29 30 40.1671 $w=1.83e-07 $l=6.7e-07 $layer=LI1_cond $X=1.47 $Y=1.137
+ $X2=0.8 $Y2=1.137
r67 28 43 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.79 $Y=1.84 $X2=0.7
+ $Y2=1.84
r68 27 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.47 $Y=1.84
+ $X2=1.565 $Y2=1.925
r69 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.47 $Y=1.84
+ $X2=0.79 $Y2=1.84
r70 23 25 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=0.7 $Y=1.98 $X2=0.7
+ $Y2=2.91
r71 21 43 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=1.925 $X2=0.7
+ $Y2=1.84
r72 21 23 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=0.7 $Y=1.925 $X2=0.7
+ $Y2=1.98
r73 17 42 1.09868 $w=1.9e-07 $l=9.2e-08 $layer=LI1_cond $X=0.705 $Y=1.045
+ $X2=0.705 $Y2=1.137
r74 17 19 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=0.705 $Y=1.045
+ $X2=0.705 $Y2=0.42
r75 16 41 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.335 $Y=1.84
+ $X2=0.222 $Y2=1.755
r76 15 43 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.61 $Y=1.84 $X2=0.7
+ $Y2=1.84
r77 15 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.61 $Y=1.84
+ $X2=0.335 $Y2=1.84
r78 14 44 3.98913 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.335 $Y=1.145
+ $X2=0.222 $Y2=1.145
r79 13 42 5.465 $w=1.77e-07 $l=9.89192e-08 $layer=LI1_cond $X=0.61 $Y=1.145
+ $X2=0.705 $Y2=1.137
r80 13 14 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.61 $Y=1.145
+ $X2=0.335 $Y2=1.145
r81 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=2.91
r82 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=1.98
r83 3 25 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.91
r84 3 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=1.98
r85 2 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.425
+ $Y=0.235 $X2=1.565 $Y2=0.42
r86 1 19 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.705 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%A_457_367# 1 2 3 4 13 15 17 21 23 26 27 28
+ 32 33 34 37 42
r68 35 37 6.4697 $w=1.78e-07 $l=1.05e-07 $layer=LI1_cond $X=6.38 $Y=1.875
+ $X2=6.38 $Y2=1.98
r69 33 35 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.29 $Y=1.79
+ $X2=6.38 $Y2=1.875
r70 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.29 $Y=1.79
+ $X2=5.62 $Y2=1.79
r71 30 32 20.611 $w=2.58e-07 $l=4.65e-07 $layer=LI1_cond $X=5.49 $Y=2.445
+ $X2=5.49 $Y2=1.98
r72 29 34 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.49 $Y=1.875
+ $X2=5.62 $Y2=1.79
r73 29 32 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=5.49 $Y=1.875
+ $X2=5.49 $Y2=1.98
r74 27 30 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.36 $Y=2.53
+ $X2=5.49 $Y2=2.445
r75 27 28 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=5.36 $Y=2.53
+ $X2=4.315 $Y2=2.53
r76 26 28 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=4.192 $Y=2.445
+ $X2=4.315 $Y2=2.53
r77 25 26 10.8189 $w=2.43e-07 $l=2.3e-07 $layer=LI1_cond $X=4.192 $Y=2.215
+ $X2=4.192 $Y2=2.445
r78 24 42 5.52892 $w=1.75e-07 $l=9.74679e-08 $layer=LI1_cond $X=3.38 $Y=2.13
+ $X2=3.285 $Y2=2.135
r79 23 25 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=4.07 $Y=2.13
+ $X2=4.192 $Y2=2.215
r80 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.07 $Y=2.13 $X2=3.38
+ $Y2=2.13
r81 19 42 1.04816 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=3.285 $Y=2.225
+ $X2=3.285 $Y2=2.135
r82 19 21 39.4019 $w=1.88e-07 $l=6.75e-07 $layer=LI1_cond $X=3.285 $Y=2.225
+ $X2=3.285 $Y2=2.9
r83 18 40 3.50369 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.52 $Y=2.135
+ $X2=2.425 $Y2=2.135
r84 17 42 5.52892 $w=1.75e-07 $l=9.5e-08 $layer=LI1_cond $X=3.19 $Y=2.135
+ $X2=3.285 $Y2=2.135
r85 17 18 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.19 $Y=2.135
+ $X2=2.52 $Y2=2.135
r86 13 40 3.31928 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=2.425 $Y=2.225
+ $X2=2.425 $Y2=2.135
r87 13 15 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=2.425 $Y=2.225
+ $X2=2.425 $Y2=2.91
r88 4 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.245
+ $Y=1.835 $X2=6.385 $Y2=1.98
r89 3 32 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=5.385
+ $Y=1.835 $X2=5.525 $Y2=1.98
r90 2 42 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=1.835 $X2=3.285 $Y2=2.21
r91 2 21 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=1.835 $X2=3.285 $Y2=2.9
r92 1 40 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.835 $X2=2.425 $Y2=2.21
r93 1 15 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.835 $X2=2.425 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%A_822_367# 1 2 3 4 13 21 23 25 27 30
c48 1 0 1.79433e-19 $X=4.11 $Y=1.835
r49 25 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=2.895
+ $X2=6.815 $Y2=2.98
r50 25 27 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=6.815 $Y=2.895
+ $X2=6.815 $Y2=2.005
r51 24 30 7.01393 $w=2.25e-07 $l=1.90526e-07 $layer=LI1_cond $X=6.12 $Y=2.98
+ $X2=5.955 $Y2=2.925
r52 23 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.65 $Y=2.98
+ $X2=6.815 $Y2=2.98
r53 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.65 $Y=2.98
+ $X2=6.12 $Y2=2.98
r54 19 30 0.00725833 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=5.955 $Y=2.785
+ $X2=5.955 $Y2=2.925
r55 19 21 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=5.955 $Y=2.785
+ $X2=5.955 $Y2=2.145
r56 15 18 35.3965 $w=2.78e-07 $l=8.6e-07 $layer=LI1_cond $X=4.235 $Y=2.925
+ $X2=5.095 $Y2=2.925
r57 13 30 7.01393 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=5.79 $Y=2.925
+ $X2=5.955 $Y2=2.925
r58 13 18 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=5.79 $Y=2.925
+ $X2=5.095 $Y2=2.925
r59 4 32 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=6.675
+ $Y=1.835 $X2=6.815 $Y2=2.9
r60 4 27 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=6.675
+ $Y=1.835 $X2=6.815 $Y2=2.005
r61 3 30 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=5.815
+ $Y=1.835 $X2=5.955 $Y2=2.9
r62 3 21 400 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_PDIFF $count=1 $X=5.815
+ $Y=1.835 $X2=5.955 $Y2=2.145
r63 2 18 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=4.955
+ $Y=1.835 $X2=5.095 $Y2=2.9
r64 1 15 600 $w=1.7e-07 $l=1.12577e-06 $layer=licon1_PDIFF $count=1 $X=4.11
+ $Y=1.835 $X2=4.235 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 47 48 49 51 63 67 77 78 84 87 90
r115 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r116 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r117 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r118 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r119 78 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r120 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r121 75 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.07 $Y=0 $X2=6.905
+ $Y2=0
r122 75 77 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.07 $Y=0 $X2=7.44
+ $Y2=0
r123 74 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r124 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r125 71 74 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r126 71 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r127 70 73 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.48
+ $Y2=0
r128 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r129 68 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.665
+ $Y2=0
r130 68 70 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=5.04
+ $Y2=0
r131 67 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.74 $Y=0 $X2=6.905
+ $Y2=0
r132 67 73 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.74 $Y=0 $X2=6.48
+ $Y2=0
r133 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r134 63 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.535 $Y=0 $X2=4.665
+ $Y2=0
r135 63 65 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=4.535 $Y=0
+ $X2=3.12 $Y2=0
r136 62 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r137 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r138 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r139 59 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r140 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r141 56 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.135
+ $Y2=0
r142 56 58 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.68
+ $Y2=0
r143 55 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r144 55 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r145 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r146 52 81 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r147 52 54 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.72
+ $Y2=0
r148 51 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.135
+ $Y2=0
r149 51 54 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.72
+ $Y2=0
r150 49 88 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=4.56
+ $Y2=0
r151 49 66 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.12
+ $Y2=0
r152 47 61 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.64
+ $Y2=0
r153 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.855
+ $Y2=0
r154 46 65 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=3.12
+ $Y2=0
r155 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=2.855
+ $Y2=0
r156 44 58 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.68
+ $Y2=0
r157 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.995
+ $Y2=0
r158 43 61 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r159 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.995
+ $Y2=0
r160 39 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0
r161 39 41 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0.39
r162 35 87 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=0.085
+ $X2=4.665 $Y2=0
r163 35 37 19.2813 $w=2.58e-07 $l=4.35e-07 $layer=LI1_cond $X=4.665 $Y=0.085
+ $X2=4.665 $Y2=0.52
r164 31 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0
r165 31 33 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0.51
r166 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0
r167 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0.38
r168 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0
r169 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0.36
r170 19 81 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r171 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.38
r172 6 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.765
+ $Y=0.245 $X2=6.905 $Y2=0.39
r173 5 37 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.235 $X2=4.665 $Y2=0.52
r174 4 33 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.855 $Y2=0.51
r175 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.855
+ $Y=0.235 $X2=1.995 $Y2=0.38
r176 2 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.995
+ $Y=0.235 $X2=1.135 $Y2=0.36
r177 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%A_457_47# 1 2 9 11 12 14
r25 11 14 7.68295 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=3.827 $Y=0.93
+ $X2=3.827 $Y2=0.76
r26 11 12 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=3.7 $Y=0.93 $X2=2.52
+ $Y2=0.93
r27 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.425 $Y=0.845
+ $X2=2.52 $Y2=0.93
r28 7 9 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=2.425 $Y=0.845
+ $X2=2.425 $Y2=0.42
r29 2 14 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.235 $X2=3.805 $Y2=0.76
r30 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.285
+ $Y=0.235 $X2=2.425 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A221O_4%A_1077_47# 1 2 3 10 16 18 22 24
c34 24 0 1.79196e-19 $X=6.31 $Y=0.685
r35 20 22 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=7.37 $Y=1.065
+ $X2=7.37 $Y2=0.42
r36 19 24 5.33677 $w=2.5e-07 $l=5.80625e-07 $layer=LI1_cond $X=6.57 $Y=1.15
+ $X2=6.31 $Y2=0.685
r37 18 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.24 $Y=1.15
+ $X2=7.37 $Y2=1.065
r38 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.24 $Y=1.15
+ $X2=6.57 $Y2=1.15
r39 14 24 1.20171 $w=2.6e-07 $l=1.3e-07 $layer=LI1_cond $X=6.44 $Y=0.685
+ $X2=6.31 $Y2=0.685
r40 14 16 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=6.44 $Y=0.685
+ $X2=6.44 $Y2=0.42
r41 10 24 5.33677 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=6.31 $Y=0.85
+ $X2=6.31 $Y2=0.685
r42 10 12 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=6.31 $Y=0.85
+ $X2=5.525 $Y2=0.85
r43 3 22 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=7.195
+ $Y=0.245 $X2=7.335 $Y2=0.42
r44 2 16 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=6.35
+ $Y=0.245 $X2=6.475 $Y2=0.42
r45 1 12 182 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_NDIFF $count=1 $X=5.385
+ $Y=0.235 $X2=5.525 $Y2=0.85
.ends

