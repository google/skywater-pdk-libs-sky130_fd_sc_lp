* NGSPICE file created from sky130_fd_sc_lp__dlclkp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
M1000 a_80_269# a_315_382# a_273_480# VPB phighvt w=640000u l=150000u
+  ad=2.221e+11p pd=2.06e+06u as=1.344e+11p ps=1.7e+06u
M1001 VPWR a_27_367# a_453_480# VPB phighvt w=420000u l=150000u
+  ad=2.04465e+12p pd=1.399e+07u as=8.82e+10p ps=1.26e+06u
M1002 a_279_81# GATE VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.07688e+12p ps=9.44e+06u
M1003 a_315_382# a_321_55# VPWR VPB phighvt w=640000u l=150000u
+  ad=2.752e+11p pd=2.14e+06u as=0p ps=0u
M1004 VGND a_27_367# a_437_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1005 a_1046_367# a_27_367# a_1002_79# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1006 a_1046_367# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1007 a_1002_79# CLK VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_80_269# a_27_367# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1009 a_453_480# a_321_55# a_80_269# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_437_81# a_315_382# a_80_269# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1011 VPWR CLK a_321_55# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.464e+11p ps=2.05e+06u
M1012 a_315_382# a_321_55# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1013 VGND CLK a_321_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1014 GCLK a_1046_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1015 GCLK a_1046_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1016 a_80_269# a_321_55# a_279_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_27_367# a_1046_367# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_273_480# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_80_269# a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

