* NGSPICE file created from sky130_fd_sc_lp__and3b_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and3b_lp A_N B C VGND VNB VPB VPWR X
M1000 a_666_57# a_248_409# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.066e+11p ps=3.14e+06u
M1001 a_391_57# a_137_408# a_248_409# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1002 X a_248_409# a_666_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1003 a_248_409# B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.65e+11p pd=5.13e+06u as=9.5e+11p ps=7.9e+06u
M1004 X a_248_409# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1005 a_114_57# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1006 a_469_57# B a_391_57# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 VGND C a_469_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_137_408# a_248_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_137_408# A_N VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1010 VPWR C a_248_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_137_408# A_N a_114_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends

