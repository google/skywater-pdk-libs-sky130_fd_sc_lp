* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2i_lp A0 A1 S VGND VNB VPB VPWR Y
X0 VGND S a_114_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR S a_125_527# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_324_49# a_365_255# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_289_527# a_365_255# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_509_49# S a_365_255# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y A0 a_324_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_125_527# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 Y A1 a_289_527# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND S a_509_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR S a_510_527# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_510_527# S a_365_255# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_114_49# A1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
