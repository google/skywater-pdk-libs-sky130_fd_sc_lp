# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__and4bb_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__and4bb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.670000 0.690000 1.785000 ;
        RECT 0.440000 1.785000 0.880000 2.530000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.785000 1.080000 1.115000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 0.750000 3.265000 1.515000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.985000 2.625000 3.345000 3.075000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.925000 0.255000 4.235000 1.095000 ;
        RECT 3.925000 2.035000 4.235000 3.075000 ;
        RECT 4.025000 1.095000 4.235000 2.035000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.090000  0.285000 0.390000 1.330000 ;
      RECT 0.090000  1.330000 1.095000 1.425000 ;
      RECT 0.090000  1.425000 1.590000 1.500000 ;
      RECT 0.090000  1.500000 0.260000 2.700000 ;
      RECT 0.090000  2.700000 0.455000 3.030000 ;
      RECT 0.560000  0.085000 0.820000 0.615000 ;
      RECT 0.625000  2.700000 0.955000 3.245000 ;
      RECT 0.925000  1.500000 1.590000 1.615000 ;
      RECT 0.990000  0.255000 2.675000 0.505000 ;
      RECT 0.990000  0.505000 1.500000 0.615000 ;
      RECT 1.125000  1.785000 1.940000 1.955000 ;
      RECT 1.125000  1.955000 1.385000 3.030000 ;
      RECT 1.330000  0.615000 1.500000 1.085000 ;
      RECT 1.330000  1.085000 1.940000 1.255000 ;
      RECT 1.610000  2.125000 1.940000 3.245000 ;
      RECT 1.680000  0.675000 2.310000 0.915000 ;
      RECT 1.770000  1.255000 1.940000 1.785000 ;
      RECT 2.110000  0.915000 2.310000 1.705000 ;
      RECT 2.110000  1.705000 3.855000 1.875000 ;
      RECT 2.110000  1.875000 2.315000 2.340000 ;
      RECT 2.485000  2.045000 2.815000 3.245000 ;
      RECT 2.985000  1.875000 3.240000 2.340000 ;
      RECT 3.410000  2.045000 3.755000 2.375000 ;
      RECT 3.435000  0.085000 3.755000 1.095000 ;
      RECT 3.515000  2.375000 3.755000 3.245000 ;
      RECT 3.605000  1.345000 3.855000 1.705000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__and4bb_1
END LIBRARY
