* File: sky130_fd_sc_lp__lsbufiso0p_lp.pxi.spice
* Created: Wed Sep  2 09:59:04 2020
* 
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%VGND N_VGND_M1017_s N_VGND_M1022_d
+ N_VGND_M1018_s N_VGND_M1014_d N_VGND_M1017_b N_VGND_c_12_p N_VGND_c_7_p
+ N_VGND_c_97_p N_VGND_c_76_p N_VGND_c_101_p VGND N_VGND_c_13_p N_VGND_c_102_p
+ N_VGND_c_77_p N_VGND_c_18_p N_VGND_c_8_p
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%VGND
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%VPB N_VPB_M1013_b VPB VPB VPB VPB VPB VPB
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%VPB
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%DESTVPB N_DESTVPB_M1020_b DESTVPB DESTVPB
+ DESTVPB DESTVPB DESTVPB DESTVPB PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%DESTVPB
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_176_987# N_A_176_987#_M1021_d
+ N_A_176_987#_M1010_d N_A_176_987#_M1020_g N_A_176_987#_M1019_g
+ N_A_176_987#_c_265_n N_A_176_987#_c_258_n N_A_176_987#_c_267_n
+ N_A_176_987#_c_268_n N_A_176_987#_c_259_n N_A_176_987#_c_269_n
+ N_A_176_987#_c_262_n PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_176_987#
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A N_A_M1013_g N_A_c_334_n N_A_M1017_g
+ N_A_M1008_g N_A_c_343_n N_A_c_346_n N_A_M1006_g N_A_M1012_g N_A_c_352_n
+ N_A_M1001_g N_A_c_360_n N_A_c_362_n A N_A_c_366_n N_A_c_368_n
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_278_47# N_A_278_47#_M1012_d
+ N_A_278_47#_M1006_d N_A_278_47#_c_405_n N_A_278_47#_M1003_g
+ N_A_278_47#_c_407_n N_A_278_47#_c_410_n N_A_278_47#_c_413_n
+ N_A_278_47#_c_416_n N_A_278_47#_M1021_g N_A_278_47#_c_419_n
+ N_A_278_47#_c_432_n N_A_278_47#_c_422_n N_A_278_47#_c_425_n
+ N_A_278_47#_c_428_n N_A_278_47#_c_433_n N_A_278_47#_c_431_n
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_278_47#
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_123_718# N_A_123_718#_M1008_s
+ N_A_123_718#_M1020_s N_A_123_718#_c_498_n N_A_123_718#_M1009_g
+ N_A_123_718#_c_499_n N_A_123_718#_M1010_g N_A_123_718#_c_500_n
+ N_A_123_718#_c_476_n N_A_123_718#_M1011_g N_A_123_718#_M1004_g
+ N_A_123_718#_M1023_g N_A_123_718#_c_485_n N_A_123_718#_c_504_n
+ N_A_123_718#_c_488_n N_A_123_718#_c_489_n N_A_123_718#_c_506_n
+ N_A_123_718#_c_490_n N_A_123_718#_c_508_n N_A_123_718#_c_509_n
+ N_A_123_718#_c_576_p N_A_123_718#_c_510_n N_A_123_718#_c_491_n
+ N_A_123_718#_c_492_n N_A_123_718#_c_493_n N_A_123_718#_c_512_n
+ N_A_123_718#_c_494_n N_A_123_718#_c_515_n N_A_123_718#_c_495_n
+ N_A_123_718#_c_497_n PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_123_718#
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_517_420# N_A_517_420#_M1016_d
+ N_A_517_420#_M1015_d N_A_517_420#_c_633_n N_A_517_420#_M1022_g
+ N_A_517_420#_c_636_n N_A_517_420#_c_641_n N_A_517_420#_c_645_n
+ N_A_517_420#_c_649_n N_A_517_420#_c_650_n N_A_517_420#_c_651_n
+ N_A_517_420#_c_652_n N_A_517_420#_c_653_n N_A_517_420#_c_656_n
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_517_420#
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%SLEEP N_SLEEP_c_707_n N_SLEEP_M1018_g
+ N_SLEEP_c_711_n N_SLEEP_M1016_g N_SLEEP_M1002_g N_SLEEP_c_716_n
+ N_SLEEP_M1005_g N_SLEEP_c_718_n N_SLEEP_c_719_n N_SLEEP_c_739_n
+ N_SLEEP_M1015_g N_SLEEP_c_720_n N_SLEEP_c_740_n N_SLEEP_c_721_n
+ N_SLEEP_M1007_g N_SLEEP_c_725_n N_SLEEP_c_726_n N_SLEEP_M1014_g
+ N_SLEEP_c_741_n N_SLEEP_M1000_g N_SLEEP_c_730_n N_SLEEP_c_731_n
+ N_SLEEP_c_742_n N_SLEEP_c_732_n SLEEP N_SLEEP_c_733_n N_SLEEP_c_735_n
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%SLEEP
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%VPWR N_VPWR_M1013_s N_VPWR_c_823_n VPWR
+ N_VPWR_c_825_n N_VPWR_c_827_n N_VPWR_c_822_n N_VPWR_c_832_n
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%VPWR
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_278_1085# N_A_278_1085#_M1019_d
+ N_A_278_1085#_M1002_s N_A_278_1085#_c_853_n N_A_278_1085#_c_849_n
+ N_A_278_1085#_c_859_n N_A_278_1085#_c_850_n N_A_278_1085#_c_851_n
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_278_1085#
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%DESTPWR N_DESTPWR_M1002_d N_DESTPWR_M1000_s
+ N_DESTPWR_c_886_n N_DESTPWR_c_887_n DESTPWR N_DESTPWR_c_888_n
+ N_DESTPWR_c_890_n N_DESTPWR_c_891_n N_DESTPWR_c_885_n N_DESTPWR_c_896_n
+ N_DESTPWR_c_897_n PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%DESTPWR
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%X N_X_M1007_s N_X_M1004_d N_X_M1023_d
+ N_X_c_954_n N_X_c_958_n N_X_c_961_n X X X X X X N_X_c_964_n X
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%X
x_PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_278_718# N_A_278_718#_M1001_d
+ N_A_278_718#_M1022_s N_A_278_718#_c_1002_n N_A_278_718#_c_1006_n
+ N_A_278_718#_c_1007_n N_A_278_718#_c_1013_n N_A_278_718#_c_1016_n
+ PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_278_718#
cc_1 N_VGND_M1017_b VPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_2 N_VGND_M1017_b VPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=6.395 $Y2=0.47
cc_3 N_VGND_M1017_b DESTVPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_4 N_VGND_M1017_b DESTVPB 0.0141757f $X=-0.025 $Y=-0.245 $X2=6.395 $Y2=0.47
cc_5 N_VGND_M1017_b N_A_176_987#_c_258_n 0.016137f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_6 N_VGND_M1017_b N_A_176_987#_c_259_n 0.00431945f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_7 N_VGND_c_7_p N_A_176_987#_c_259_n 0.0120094f $X=2.865 $Y=4.155 $X2=0 $Y2=0
cc_8 N_VGND_c_8_p N_A_176_987#_c_259_n 0.00149965f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_9 N_VGND_M1017_b N_A_176_987#_c_262_n 0.0169579f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_10 N_VGND_M1017_b N_A_M1013_g 0.00622578f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_11 N_VGND_M1017_b N_A_c_334_n 0.0206818f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_12 N_VGND_c_12_p N_A_c_334_n 0.00818476f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_13 N_VGND_c_13_p N_A_c_334_n 9.22492e-19 $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_14 N_VGND_c_8_p N_A_c_334_n 7.18026e-19 $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_15 N_VGND_M1017_b N_A_M1008_g 0.0399099f $X=-0.025 $Y=-0.245 $X2=0.155
+ $Y2=0.84
cc_16 N_VGND_c_12_p N_A_M1008_g 0.00429861f $X=0.74 $Y=2.44 $X2=0.155 $Y2=0.84
cc_17 N_VGND_c_13_p N_A_M1008_g 0.00909137f $X=1.68 $Y=3.33 $X2=0.155 $Y2=0.84
cc_18 N_VGND_c_18_p N_A_M1008_g 0.00506743f $X=0.72 $Y=3.33 $X2=0.155 $Y2=0.84
cc_19 N_VGND_c_8_p N_A_M1008_g 0.0108583f $X=6.48 $Y=3.33 $X2=0.155 $Y2=0.84
cc_20 N_VGND_M1017_b N_A_c_343_n 0.0114117f $X=-0.025 $Y=-0.245 $X2=6.395
+ $Y2=0.47
cc_21 N_VGND_c_13_p N_A_c_343_n 5.14398e-19 $X=1.68 $Y=3.33 $X2=6.395 $Y2=0.47
cc_22 N_VGND_c_8_p N_A_c_343_n 0.00400159f $X=6.48 $Y=3.33 $X2=6.395 $Y2=0.47
cc_23 N_VGND_M1017_b N_A_c_346_n 0.00960464f $X=-0.025 $Y=-0.245 $X2=6.395
+ $Y2=0.84
cc_24 N_VGND_c_12_p N_A_c_346_n 0.00626201f $X=0.74 $Y=2.44 $X2=6.395 $Y2=0.84
cc_25 N_VGND_c_8_p N_A_c_346_n 0.00228999f $X=6.48 $Y=3.33 $X2=6.395 $Y2=0.84
cc_26 N_VGND_M1017_b N_A_M1006_g 0.00537455f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_27 N_VGND_M1017_b N_A_M1012_g 0.0097482f $X=-0.025 $Y=-0.245 $X2=0.24
+ $Y2=0.525
cc_28 N_VGND_c_12_p N_A_M1012_g 3.60856e-19 $X=0.74 $Y=2.44 $X2=0.24 $Y2=0.525
cc_29 N_VGND_M1017_b N_A_c_352_n 0.032122f $X=-0.025 $Y=-0.245 $X2=0.24
+ $Y2=0.525
cc_30 N_VGND_c_12_p N_A_c_352_n 5.98673e-19 $X=0.74 $Y=2.44 $X2=0.24 $Y2=0.525
cc_31 N_VGND_c_13_p N_A_c_352_n 0.0030635f $X=1.68 $Y=3.33 $X2=0.24 $Y2=0.525
cc_32 N_VGND_c_8_p N_A_c_352_n 0.00643718f $X=6.48 $Y=3.33 $X2=0.24 $Y2=0.525
cc_33 N_VGND_M1017_b N_A_M1001_g 0.029645f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_34 N_VGND_c_12_p N_A_M1001_g 8.81789e-19 $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_35 N_VGND_c_13_p N_A_M1001_g 0.0110813f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_36 N_VGND_c_8_p N_A_M1001_g 0.00964689f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_37 N_VGND_M1017_b N_A_c_360_n 0.00229529f $X=-0.025 $Y=-0.245 $X2=0.24
+ $Y2=1.295
cc_38 N_VGND_c_12_p N_A_c_360_n 0.0223008f $X=0.74 $Y=2.44 $X2=0.24 $Y2=1.295
cc_39 N_VGND_M1017_b N_A_c_362_n 0.00551809f $X=-0.025 $Y=-0.245 $X2=6.48
+ $Y2=0.525
cc_40 N_VGND_c_12_p N_A_c_362_n 0.0252639f $X=0.74 $Y=2.44 $X2=6.48 $Y2=0.525
cc_41 N_VGND_c_13_p N_A_c_362_n 0.0362016f $X=1.68 $Y=3.33 $X2=6.48 $Y2=0.525
cc_42 N_VGND_c_8_p N_A_c_362_n 0.0196655f $X=6.48 $Y=3.33 $X2=6.48 $Y2=0.525
cc_43 N_VGND_M1017_b N_A_c_366_n 0.0674831f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_44 N_VGND_c_12_p N_A_c_366_n 0.00213349f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_45 N_VGND_M1017_b N_A_c_368_n 0.0344278f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_46 N_VGND_c_12_p N_A_c_368_n 0.0262117f $X=0.74 $Y=2.44 $X2=0 $Y2=0
cc_47 N_VGND_M1017_b N_A_278_47#_c_405_n 0.012966f $X=-0.025 $Y=-0.245
+ $X2=-0.025 $Y2=-0.19
cc_48 N_VGND_c_8_p N_A_278_47#_c_405_n 0.00222998f $X=6.48 $Y=3.33 $X2=-0.025
+ $Y2=-0.19
cc_49 N_VGND_M1017_b N_A_278_47#_c_407_n 0.00602992f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=0.84
cc_50 N_VGND_c_13_p N_A_278_47#_c_407_n 0.00312162f $X=1.68 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_51 N_VGND_c_8_p N_A_278_47#_c_407_n 2.63629e-19 $X=6.48 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_52 N_VGND_M1017_b N_A_278_47#_c_410_n 0.00857286f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=1.21
cc_53 N_VGND_c_13_p N_A_278_47#_c_410_n 0.00482701f $X=1.68 $Y=3.33 $X2=0.155
+ $Y2=1.21
cc_54 N_VGND_c_8_p N_A_278_47#_c_410_n 6.46318e-19 $X=6.48 $Y=3.33 $X2=0.155
+ $Y2=1.21
cc_55 N_VGND_M1017_b N_A_278_47#_c_413_n 0.0164815f $X=-0.025 $Y=-0.245
+ $X2=6.395 $Y2=0.84
cc_56 N_VGND_c_13_p N_A_278_47#_c_413_n 0.00507498f $X=1.68 $Y=3.33 $X2=6.395
+ $Y2=0.84
cc_57 N_VGND_c_8_p N_A_278_47#_c_413_n 0.00497945f $X=6.48 $Y=3.33 $X2=6.395
+ $Y2=0.84
cc_58 N_VGND_M1017_b N_A_278_47#_c_416_n 0.0162397f $X=-0.025 $Y=-0.245
+ $X2=6.395 $Y2=1.21
cc_59 N_VGND_c_7_p N_A_278_47#_c_416_n 0.00860948f $X=2.865 $Y=4.155 $X2=6.395
+ $Y2=1.21
cc_60 N_VGND_c_8_p N_A_278_47#_c_416_n 0.00271031f $X=6.48 $Y=3.33 $X2=6.395
+ $Y2=1.21
cc_61 N_VGND_M1017_b N_A_278_47#_c_419_n 0.00923091f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_62 N_VGND_c_13_p N_A_278_47#_c_419_n 0.00190461f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_63 N_VGND_c_8_p N_A_278_47#_c_419_n 0.00291644f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_64 N_VGND_M1017_b N_A_278_47#_c_422_n 0.0216596f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_65 N_VGND_c_13_p N_A_278_47#_c_422_n 0.00259986f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_66 N_VGND_c_8_p N_A_278_47#_c_422_n 0.00569686f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_67 N_VGND_M1017_b N_A_278_47#_c_425_n 0.00372993f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_68 N_VGND_c_13_p N_A_278_47#_c_425_n 0.0220216f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_69 N_VGND_c_8_p N_A_278_47#_c_425_n 0.012589f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_70 N_VGND_M1017_b N_A_278_47#_c_428_n 0.0371605f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_71 N_VGND_c_13_p N_A_278_47#_c_428_n 8.65569e-19 $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_72 N_VGND_c_8_p N_A_278_47#_c_428_n 0.00157003f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_73 N_VGND_M1017_b N_A_278_47#_c_431_n 0.0355797f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_74 N_VGND_M1017_b N_A_123_718#_c_476_n 0.0149084f $X=-0.025 $Y=-0.245
+ $X2=6.395 $Y2=1.21
cc_75 N_VGND_M1017_b N_A_123_718#_M1011_g 0.0207676f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_76 N_VGND_c_76_p N_A_123_718#_M1011_g 0.00982261f $X=5.19 $Y=3.715 $X2=0
+ $Y2=0
cc_77 N_VGND_c_77_p N_A_123_718#_M1011_g 0.00465098f $X=6.33 $Y=3.33 $X2=0 $Y2=0
cc_78 N_VGND_c_8_p N_A_123_718#_M1011_g 0.00800632f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_79 N_VGND_M1017_b N_A_123_718#_M1004_g 0.0309972f $X=-0.025 $Y=-0.245
+ $X2=0.24 $Y2=0.525
cc_80 N_VGND_c_76_p N_A_123_718#_M1004_g 0.00178951f $X=5.19 $Y=3.715 $X2=0.24
+ $Y2=0.525
cc_81 N_VGND_c_77_p N_A_123_718#_M1004_g 0.00525141f $X=6.33 $Y=3.33 $X2=0.24
+ $Y2=0.525
cc_82 N_VGND_c_8_p N_A_123_718#_M1004_g 0.01053f $X=6.48 $Y=3.33 $X2=0.24
+ $Y2=0.525
cc_83 N_VGND_M1017_b N_A_123_718#_c_485_n 0.101989f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_84 N_VGND_c_18_p N_A_123_718#_c_485_n 0.0205041f $X=0.72 $Y=3.33 $X2=0 $Y2=0
cc_85 N_VGND_c_8_p N_A_123_718#_c_485_n 0.0106717f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_86 N_VGND_M1017_b N_A_123_718#_c_488_n 0.0267048f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_87 N_VGND_M1017_b N_A_123_718#_c_489_n 0.00597888f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_88 N_VGND_M1017_b N_A_123_718#_c_490_n 0.00640786f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_89 N_VGND_M1017_b N_A_123_718#_c_491_n 0.00794591f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_90 N_VGND_M1017_b N_A_123_718#_c_492_n 0.00690568f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_91 N_VGND_M1017_b N_A_123_718#_c_493_n 0.0152338f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_92 N_VGND_M1017_b N_A_123_718#_c_494_n 0.0119951f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_93 N_VGND_M1017_b N_A_123_718#_c_495_n 0.0155539f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_94 N_VGND_c_7_p N_A_123_718#_c_495_n 0.00116779f $X=2.865 $Y=4.155 $X2=0
+ $Y2=0
cc_95 N_VGND_M1017_b N_A_123_718#_c_497_n 0.036852f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_96 N_VGND_M1017_b N_A_517_420#_c_633_n 0.0273206f $X=-0.025 $Y=-0.245
+ $X2=-0.025 $Y2=-0.19
cc_97 N_VGND_c_97_p N_A_517_420#_c_633_n 0.0108288f $X=2.875 $Y=2.515 $X2=-0.025
+ $Y2=-0.19
cc_98 N_VGND_c_8_p N_A_517_420#_c_633_n 0.00642949f $X=6.48 $Y=3.33 $X2=-0.025
+ $Y2=-0.19
cc_99 N_VGND_M1017_b N_A_517_420#_c_636_n 0.0943772f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=0.84
cc_100 N_VGND_c_97_p N_A_517_420#_c_636_n 0.012424f $X=2.875 $Y=2.515 $X2=0.155
+ $Y2=0.84
cc_101 N_VGND_c_101_p N_A_517_420#_c_636_n 0.00850832f $X=2.87 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_102 N_VGND_c_102_p N_A_517_420#_c_636_n 0.0351019f $X=5.025 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_103 N_VGND_c_8_p N_A_517_420#_c_636_n 0.0103238f $X=6.48 $Y=3.33 $X2=0.155
+ $Y2=0.84
cc_104 N_VGND_M1017_b N_A_517_420#_c_641_n 0.0101923f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=1.21
cc_105 N_VGND_c_97_p N_A_517_420#_c_641_n 7.79356e-19 $X=2.875 $Y=2.515
+ $X2=0.155 $Y2=1.21
cc_106 N_VGND_c_101_p N_A_517_420#_c_641_n 0.00153142f $X=2.87 $Y=3.33 $X2=0.155
+ $Y2=1.21
cc_107 N_VGND_c_8_p N_A_517_420#_c_641_n 0.00282686f $X=6.48 $Y=3.33 $X2=0.155
+ $Y2=1.21
cc_108 N_VGND_M1017_b N_A_517_420#_c_645_n 0.0159984f $X=-0.025 $Y=-0.245
+ $X2=6.395 $Y2=1.21
cc_109 N_VGND_c_7_p N_A_517_420#_c_645_n 0.025063f $X=2.865 $Y=4.155 $X2=6.395
+ $Y2=1.21
cc_110 N_VGND_c_102_p N_A_517_420#_c_645_n 0.0400923f $X=5.025 $Y=3.33 $X2=6.395
+ $Y2=1.21
cc_111 N_VGND_c_8_p N_A_517_420#_c_645_n 0.0217427f $X=6.48 $Y=3.33 $X2=6.395
+ $Y2=1.21
cc_112 N_VGND_M1017_b N_A_517_420#_c_649_n 0.00529491f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_113 N_VGND_M1017_b N_A_517_420#_c_650_n 0.0120215f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_114 N_VGND_M1017_b N_A_517_420#_c_651_n 0.00296389f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_115 N_VGND_M1017_b N_A_517_420#_c_652_n 0.00148259f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_116 N_VGND_M1017_b N_A_517_420#_c_653_n 0.0406717f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_117 N_VGND_c_102_p N_A_517_420#_c_653_n 0.00336816f $X=5.025 $Y=3.33 $X2=0
+ $Y2=0
cc_118 N_VGND_c_8_p N_A_517_420#_c_653_n 0.00254324f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_119 N_VGND_M1017_b N_A_517_420#_c_656_n 0.0217853f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_120 N_VGND_c_102_p N_A_517_420#_c_656_n 0.00847838f $X=5.025 $Y=3.33 $X2=0
+ $Y2=0
cc_121 N_VGND_c_8_p N_A_517_420#_c_656_n 0.00581174f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_122 N_VGND_M1017_b N_SLEEP_c_707_n 0.0164714f $X=-0.025 $Y=-0.245 $X2=0.155
+ $Y2=0.32
cc_123 N_VGND_c_7_p N_SLEEP_c_707_n 0.00923491f $X=2.865 $Y=4.155 $X2=0.155
+ $Y2=0.32
cc_124 N_VGND_c_102_p N_SLEEP_c_707_n 0.00153691f $X=5.025 $Y=3.33 $X2=0.155
+ $Y2=0.32
cc_125 N_VGND_c_8_p N_SLEEP_c_707_n 0.00245232f $X=6.48 $Y=3.33 $X2=0.155
+ $Y2=0.32
cc_126 N_VGND_M1017_b N_SLEEP_c_711_n 0.0152475f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_127 N_VGND_c_7_p N_SLEEP_c_711_n 9.79299e-19 $X=2.865 $Y=4.155 $X2=0 $Y2=0
cc_128 N_VGND_c_102_p N_SLEEP_c_711_n 0.00171734f $X=5.025 $Y=3.33 $X2=0 $Y2=0
cc_129 N_VGND_c_8_p N_SLEEP_c_711_n 0.00243285f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_130 N_VGND_M1017_b N_SLEEP_M1002_g 0.00758372f $X=-0.025 $Y=-0.245 $X2=0.155
+ $Y2=0.47
cc_131 N_VGND_M1017_b N_SLEEP_c_716_n 0.0126934f $X=-0.025 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_132 N_VGND_M1017_b N_SLEEP_M1005_g 0.0138913f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_133 N_VGND_M1017_b N_SLEEP_c_718_n 0.0101995f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_134 N_VGND_M1017_b N_SLEEP_c_719_n 0.0154757f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_135 N_VGND_M1017_b N_SLEEP_c_720_n 0.0127025f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_136 N_VGND_M1017_b N_SLEEP_c_721_n 0.0158388f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_137 N_VGND_c_76_p N_SLEEP_c_721_n 0.00180098f $X=5.19 $Y=3.715 $X2=0 $Y2=0
cc_138 N_VGND_c_102_p N_SLEEP_c_721_n 0.00525297f $X=5.025 $Y=3.33 $X2=0 $Y2=0
cc_139 N_VGND_c_8_p N_SLEEP_c_721_n 0.0099313f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_140 N_VGND_M1017_b N_SLEEP_c_725_n 0.0184474f $X=-0.025 $Y=-0.245 $X2=6.48
+ $Y2=0.525
cc_141 N_VGND_M1017_b N_SLEEP_c_726_n 0.0131929f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_142 N_VGND_c_76_p N_SLEEP_c_726_n 0.00982947f $X=5.19 $Y=3.715 $X2=0 $Y2=0
cc_143 N_VGND_c_102_p N_SLEEP_c_726_n 0.00465098f $X=5.025 $Y=3.33 $X2=0 $Y2=0
cc_144 N_VGND_c_8_p N_SLEEP_c_726_n 0.00800632f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_145 N_VGND_M1017_b N_SLEEP_c_730_n 0.00688864f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_146 N_VGND_M1017_b N_SLEEP_c_731_n 0.00994534f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_147 N_VGND_M1017_b N_SLEEP_c_732_n 0.00639424f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_148 N_VGND_M1017_b N_SLEEP_c_733_n 0.0126999f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_149 N_VGND_c_7_p N_SLEEP_c_733_n 0.010359f $X=2.865 $Y=4.155 $X2=0 $Y2=0
cc_150 N_VGND_M1017_b N_SLEEP_c_735_n 0.0456607f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_151 N_VGND_M1017_b N_VPWR_c_822_n 0.283096f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_152 N_VGND_M1017_b N_DESTPWR_c_885_n 0.283096f $X=-0.025 $Y=-0.245 $X2=0
+ $Y2=0
cc_153 N_VGND_M1017_b N_X_c_954_n 0.00144788f $X=-0.025 $Y=-0.245 $X2=6.395
+ $Y2=0.47
cc_154 N_VGND_c_76_p N_X_c_954_n 0.00958206f $X=5.19 $Y=3.715 $X2=6.395 $Y2=0.47
cc_155 N_VGND_c_102_p N_X_c_954_n 0.0169429f $X=5.025 $Y=3.33 $X2=6.395 $Y2=0.47
cc_156 N_VGND_c_8_p N_X_c_954_n 0.0105342f $X=6.48 $Y=3.33 $X2=6.395 $Y2=0.47
cc_157 N_VGND_M1014_d N_X_c_958_n 0.00279751f $X=5.05 $Y=3.59 $X2=6.395 $Y2=1.21
cc_158 N_VGND_M1017_b N_X_c_958_n 0.00881818f $X=-0.025 $Y=-0.245 $X2=6.395
+ $Y2=1.21
cc_159 N_VGND_c_76_p N_X_c_958_n 0.00828326f $X=5.19 $Y=3.715 $X2=6.395 $Y2=1.21
cc_160 N_VGND_M1017_b N_X_c_961_n 0.00340813f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_161 N_VGND_M1017_b X 0.0161518f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_162 N_VGND_M1017_b X 0.0347182f $X=-0.025 $Y=-0.245 $X2=0 $Y2=0
cc_163 N_VGND_M1017_b N_X_c_964_n 0.0675226f $X=-0.025 $Y=-0.245 $X2=6.48
+ $Y2=0.525
cc_164 N_VGND_c_76_p N_X_c_964_n 0.00986992f $X=5.19 $Y=3.715 $X2=6.48 $Y2=0.525
cc_165 N_VGND_c_77_p N_X_c_964_n 0.0234355f $X=6.33 $Y=3.33 $X2=6.48 $Y2=0.525
cc_166 N_VGND_c_8_p N_X_c_964_n 0.0124904f $X=6.48 $Y=3.33 $X2=6.48 $Y2=0.525
cc_167 N_VGND_M1017_b N_A_278_718#_c_1002_n 0.00481358f $X=-0.025 $Y=-0.245
+ $X2=0.155 $Y2=0.47
cc_168 N_VGND_c_7_p N_A_278_718#_c_1002_n 0.0127465f $X=2.865 $Y=4.155 $X2=0.155
+ $Y2=0.47
cc_169 N_VGND_c_13_p N_A_278_718#_c_1002_n 0.03008f $X=1.68 $Y=3.33 $X2=0.155
+ $Y2=0.47
cc_170 N_VGND_c_8_p N_A_278_718#_c_1002_n 0.0273016f $X=6.48 $Y=3.33 $X2=0.155
+ $Y2=0.47
cc_171 N_VGND_M1017_b N_A_278_718#_c_1006_n 0.00602893f $X=-0.025 $Y=-0.245
+ $X2=6.395 $Y2=0.84
cc_172 N_VGND_M1017_b N_A_278_718#_c_1007_n 0.00954178f $X=-0.025 $Y=-0.245
+ $X2=0 $Y2=0
cc_173 N_VGND_c_7_p N_A_278_718#_c_1007_n 0.00977302f $X=2.865 $Y=4.155 $X2=0
+ $Y2=0
cc_174 N_VGND_c_97_p N_A_278_718#_c_1007_n 0.00780714f $X=2.875 $Y=2.515 $X2=0
+ $Y2=0
cc_175 N_VGND_c_101_p N_A_278_718#_c_1007_n 0.009578f $X=2.87 $Y=3.33 $X2=0
+ $Y2=0
cc_176 N_VGND_c_13_p N_A_278_718#_c_1007_n 0.0115155f $X=1.68 $Y=3.33 $X2=0
+ $Y2=0
cc_177 N_VGND_c_8_p N_A_278_718#_c_1007_n 0.0299959f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_178 N_VGND_M1017_b N_A_278_718#_c_1013_n 0.00440914f $X=-0.025 $Y=-0.245
+ $X2=0 $Y2=0
cc_179 N_VGND_c_13_p N_A_278_718#_c_1013_n 0.0199194f $X=1.68 $Y=3.33 $X2=0
+ $Y2=0
cc_180 N_VGND_c_8_p N_A_278_718#_c_1013_n 0.0106419f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_181 N_VGND_M1017_b N_A_278_718#_c_1016_n 0.00150928f $X=-0.025 $Y=-0.245
+ $X2=0 $Y2=0
cc_182 N_VGND_c_97_p N_A_278_718#_c_1016_n 0.0242302f $X=2.875 $Y=2.515 $X2=0
+ $Y2=0
cc_183 N_VGND_c_8_p N_A_278_718#_c_1016_n 0.0150209f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPB_M1013_b N_A_M1013_g 0.0389027f $X=-0.025 $Y=-0.19 $X2=2.74 $Y2=4.01
cc_185 VPB N_A_M1013_g 0.00621856f $X=0.155 $Y=0.47 $X2=2.74 $Y2=4.01
cc_186 N_VPB_M1013_b N_A_M1006_g 0.0358449f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_187 N_VPB_M1013_b N_A_c_368_n 0.0183257f $X=-0.025 $Y=-0.19 $X2=2.875
+ $Y2=3.245
cc_188 N_VPB_M1013_b N_A_278_47#_c_432_n 0.0369401f $X=-0.025 $Y=-0.19 $X2=0
+ $Y2=0
cc_189 N_VPB_M1013_b N_A_278_47#_c_433_n 0.00836222f $X=-0.025 $Y=-0.19 $X2=0.24
+ $Y2=3.245
cc_190 N_VPB_M1013_b N_A_278_47#_c_431_n 0.0164461f $X=-0.025 $Y=-0.19 $X2=0
+ $Y2=0
cc_191 N_VPB_M1013_b N_VPWR_c_823_n 0.0144492f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_823_n 0.0708842f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_193 N_VPB_M1013_b N_VPWR_c_825_n 0.0176917f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_825_n 0.0200925f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_195 N_VPB_M1013_b N_VPWR_c_827_n 0.180182f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_827_n 0.0200925f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_197 N_VPB_M1013_b N_VPWR_c_822_n 0.2494f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_822_n 0.0115306f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_822_n 0.0115306f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_200 N_VPB_M1013_b N_VPWR_c_832_n 0.00513431f $X=-0.025 $Y=-0.19 $X2=0 $Y2=0
cc_201 N_DESTVPB_M1020_b N_A_176_987#_M1020_g 0.0210833f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_202 N_DESTVPB_M1020_b N_A_176_987#_M1019_g 0.0170453f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_203 N_DESTVPB_M1020_b N_A_176_987#_c_265_n 0.00720677f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_204 N_DESTVPB_M1020_b N_A_176_987#_c_258_n 0.00300406f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_205 N_DESTVPB_M1020_b N_A_176_987#_c_267_n 0.0088759f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_206 N_DESTVPB_M1020_b N_A_176_987#_c_268_n 0.00229064f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_207 N_DESTVPB_M1020_b N_A_176_987#_c_269_n 0.00401794f $X=-0.025 $Y=4.985
+ $X2=0.24 $Y2=3.245
cc_208 N_DESTVPB_M1020_b N_A_176_987#_c_262_n 0.0274464f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_209 N_DESTVPB_M1020_b N_A_123_718#_c_498_n 0.0130622f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_210 N_DESTVPB_M1020_b N_A_123_718#_c_499_n 0.0167244f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_211 N_DESTVPB_M1020_b N_A_123_718#_c_500_n 0.0141652f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_212 N_DESTVPB_M1020_b N_A_123_718#_c_476_n 0.0331088f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_213 N_DESTVPB_M1020_b N_A_123_718#_M1023_g 0.0458036f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_214 DESTVPB N_A_123_718#_M1023_g 0.00224388f $X=6.395 $Y=5.28 $X2=0 $Y2=0
cc_215 N_DESTVPB_M1020_b N_A_123_718#_c_504_n 0.00931091f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_216 N_DESTVPB_M1020_b N_A_123_718#_c_489_n 3.94425e-19 $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_217 N_DESTVPB_M1020_b N_A_123_718#_c_506_n 0.0353002f $X=-0.025 $Y=4.985
+ $X2=0.575 $Y2=3.33
cc_218 N_DESTVPB_M1020_b N_A_123_718#_c_490_n 6.71603e-19 $X=-0.025 $Y=4.985
+ $X2=0.39 $Y2=3.33
cc_219 N_DESTVPB_M1020_b N_A_123_718#_c_508_n 0.00153126f $X=-0.025 $Y=4.985
+ $X2=0.74 $Y2=2.44
cc_220 N_DESTVPB_M1020_b N_A_123_718#_c_509_n 0.00872435f $X=-0.025 $Y=4.985
+ $X2=0.74 $Y2=2.44
cc_221 N_DESTVPB_M1020_b N_A_123_718#_c_510_n 0.0263702f $X=-0.025 $Y=4.985
+ $X2=2.865 $Y2=4.155
cc_222 N_DESTVPB_M1020_b N_A_123_718#_c_492_n 0.00435325f $X=-0.025 $Y=4.985
+ $X2=2.875 $Y2=3.245
cc_223 N_DESTVPB_M1020_b N_A_123_718#_c_512_n 0.00192794f $X=-0.025 $Y=4.985
+ $X2=5.19 $Y2=3.715
cc_224 N_DESTVPB_M1020_b N_A_123_718#_c_494_n 0.0165636f $X=-0.025 $Y=4.985
+ $X2=5.19 $Y2=3.715
cc_225 DESTVPB N_A_123_718#_c_494_n 0.0914628f $X=0.155 $Y=5.28 $X2=5.19
+ $Y2=3.715
cc_226 N_DESTVPB_M1020_b N_A_123_718#_c_515_n 0.00338836f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_227 N_DESTVPB_M1020_b N_A_123_718#_c_495_n 0.0426489f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_228 N_DESTVPB_M1020_b N_A_123_718#_c_497_n 0.0144582f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_229 N_DESTVPB_M1020_b N_A_517_420#_c_652_n 0.0047836f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_230 N_DESTVPB_M1020_b N_SLEEP_M1002_g 0.0403619f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_231 N_DESTVPB_M1020_b N_SLEEP_M1005_g 0.0298061f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_232 N_DESTVPB_M1020_b N_SLEEP_c_719_n 0.00862085f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_233 N_DESTVPB_M1020_b N_SLEEP_c_739_n 0.0163404f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_234 N_DESTVPB_M1020_b N_SLEEP_c_740_n 0.0772177f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_235 N_DESTVPB_M1020_b N_SLEEP_c_741_n 0.016382f $X=-0.025 $Y=4.985 $X2=0.24
+ $Y2=3.415
cc_236 N_DESTVPB_M1020_b N_SLEEP_c_742_n 0.00388587f $X=-0.025 $Y=4.985
+ $X2=0.575 $Y2=3.33
cc_237 N_DESTVPB_M1020_b N_A_278_1085#_c_849_n 0.0278512f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_238 N_DESTVPB_M1020_b N_A_278_1085#_c_850_n 4.74859e-19 $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_239 N_DESTVPB_M1020_b N_A_278_1085#_c_851_n 0.0172271f $X=-0.025 $Y=4.985
+ $X2=0 $Y2=0
cc_240 N_DESTVPB_M1020_b N_DESTPWR_c_886_n 0.0062934f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_241 N_DESTVPB_M1020_b N_DESTPWR_c_887_n 0.0154453f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_242 N_DESTVPB_M1020_b N_DESTPWR_c_888_n 0.0900644f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_243 DESTVPB N_DESTPWR_c_888_n 0.0200925f $X=0.155 $Y=5.28 $X2=0 $Y2=0
cc_244 N_DESTVPB_M1020_b N_DESTPWR_c_890_n 0.0328717f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_245 N_DESTVPB_M1020_b N_DESTPWR_c_891_n 0.0385711f $X=-0.025 $Y=4.985
+ $X2=0.24 $Y2=3.415
cc_246 DESTVPB N_DESTPWR_c_891_n 0.0200925f $X=6.395 $Y=5.28 $X2=0.24 $Y2=3.415
cc_247 N_DESTVPB_M1020_b N_DESTPWR_c_885_n 0.0806078f $X=-0.025 $Y=4.985
+ $X2=0.24 $Y2=3.855
cc_248 DESTVPB N_DESTPWR_c_885_n 0.0115306f $X=0.155 $Y=5.28 $X2=0.24 $Y2=3.855
cc_249 DESTVPB N_DESTPWR_c_885_n 0.0115306f $X=6.395 $Y=5.28 $X2=0.24 $Y2=3.855
cc_250 N_DESTVPB_M1020_b N_DESTPWR_c_896_n 0.00324402f $X=-0.025 $Y=4.985 $X2=0
+ $Y2=0
cc_251 N_DESTVPB_M1020_b N_DESTPWR_c_897_n 0.00481989f $X=-0.025 $Y=4.985
+ $X2=0.74 $Y2=3.245
cc_252 N_DESTVPB_M1020_b X 0.0240847f $X=-0.025 $Y=4.985 $X2=0 $Y2=0
cc_253 DESTVPB X 0.0915263f $X=6.395 $Y=5.28 $X2=0 $Y2=0
cc_254 N_A_176_987#_c_262_n N_A_M1008_g 0.00436304f $X=1.315 $Y=5.1 $X2=0 $Y2=0
cc_255 N_A_176_987#_c_262_n N_A_M1001_g 0.00436304f $X=1.315 $Y=5.1 $X2=0 $Y2=0
cc_256 N_A_176_987#_c_259_n N_A_278_47#_c_405_n 0.00155306f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_257 N_A_176_987#_c_258_n N_A_278_47#_c_416_n 0.00534252f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_258 N_A_176_987#_c_259_n N_A_278_47#_c_416_n 0.00599326f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_259 N_A_176_987#_c_265_n N_A_123_718#_c_498_n 0.0137915f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_260 N_A_176_987#_c_267_n N_A_123_718#_c_498_n 0.00182938f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_261 N_A_176_987#_c_265_n N_A_123_718#_c_499_n 0.0137481f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_262 N_A_176_987#_c_267_n N_A_123_718#_c_499_n 0.00899114f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_263 N_A_176_987#_c_269_n N_A_123_718#_c_499_n 0.0015814f $X=2.155 $Y=5.355
+ $X2=0 $Y2=0
cc_264 N_A_176_987#_c_258_n N_A_123_718#_c_500_n 0.0124296f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_265 N_A_176_987#_c_269_n N_A_123_718#_c_500_n 0.00779865f $X=2.155 $Y=5.355
+ $X2=0 $Y2=0
cc_266 N_A_176_987#_M1019_g N_A_123_718#_c_476_n 0.0275551f $X=1.315 $Y=5.925
+ $X2=0 $Y2=0
cc_267 N_A_176_987#_c_265_n N_A_123_718#_c_476_n 0.00279508f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_268 N_A_176_987#_c_258_n N_A_123_718#_c_476_n 0.00893677f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_269 N_A_176_987#_c_268_n N_A_123_718#_c_476_n 0.00130944f $X=1.165 $Y=5.1
+ $X2=0 $Y2=0
cc_270 N_A_176_987#_c_262_n N_A_123_718#_c_476_n 0.0219836f $X=1.315 $Y=5.1
+ $X2=0 $Y2=0
cc_271 N_A_176_987#_M1020_g N_A_123_718#_c_504_n 0.0139667f $X=0.955 $Y=5.925
+ $X2=0 $Y2=0
cc_272 N_A_176_987#_c_265_n N_A_123_718#_c_488_n 0.00619807f $X=2.155 $Y=5.44
+ $X2=0.24 $Y2=3.855
cc_273 N_A_176_987#_c_258_n N_A_123_718#_c_488_n 0.00714341f $X=2.24 $Y=5.355
+ $X2=0.24 $Y2=3.855
cc_274 N_A_176_987#_c_268_n N_A_123_718#_c_488_n 0.0252464f $X=1.165 $Y=5.1
+ $X2=0.24 $Y2=3.855
cc_275 N_A_176_987#_c_262_n N_A_123_718#_c_488_n 0.0102483f $X=1.315 $Y=5.1
+ $X2=0.24 $Y2=3.855
cc_276 N_A_176_987#_c_258_n N_A_123_718#_c_489_n 0.00682589f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_277 N_A_176_987#_c_268_n N_A_123_718#_c_489_n 0.00138846f $X=1.165 $Y=5.1
+ $X2=0 $Y2=0
cc_278 N_A_176_987#_c_262_n N_A_123_718#_c_489_n 0.00132465f $X=1.315 $Y=5.1
+ $X2=0 $Y2=0
cc_279 N_A_176_987#_c_258_n N_A_123_718#_c_490_n 0.0269829f $X=2.24 $Y=5.355
+ $X2=0.39 $Y2=3.33
cc_280 N_A_176_987#_M1020_g N_A_123_718#_c_512_n 0.00381798f $X=0.955 $Y=5.925
+ $X2=5.19 $Y2=3.715
cc_281 N_A_176_987#_M1019_g N_A_123_718#_c_512_n 0.00296352f $X=1.315 $Y=5.925
+ $X2=5.19 $Y2=3.715
cc_282 N_A_176_987#_c_268_n N_A_123_718#_c_512_n 0.00581585f $X=1.165 $Y=5.1
+ $X2=5.19 $Y2=3.715
cc_283 N_A_176_987#_c_268_n N_A_123_718#_c_494_n 0.0299155f $X=1.165 $Y=5.1
+ $X2=5.19 $Y2=3.715
cc_284 N_A_176_987#_c_262_n N_A_123_718#_c_494_n 0.0143834f $X=1.315 $Y=5.1
+ $X2=5.19 $Y2=3.715
cc_285 N_A_176_987#_c_265_n N_A_123_718#_c_515_n 0.0290917f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_286 N_A_176_987#_c_258_n N_A_123_718#_c_515_n 0.0107546f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_287 N_A_176_987#_c_268_n N_A_123_718#_c_515_n 0.0129286f $X=1.165 $Y=5.1
+ $X2=0 $Y2=0
cc_288 N_A_176_987#_c_262_n N_A_123_718#_c_515_n 0.00119275f $X=1.315 $Y=5.1
+ $X2=0 $Y2=0
cc_289 N_A_176_987#_c_258_n N_A_123_718#_c_495_n 0.00266191f $X=2.24 $Y=5.355
+ $X2=0 $Y2=0
cc_290 N_A_176_987#_c_259_n N_A_123_718#_c_495_n 0.00195932f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_291 N_A_176_987#_c_258_n N_SLEEP_c_707_n 0.00213092f $X=2.24 $Y=5.355
+ $X2=0.615 $Y2=2.23
cc_292 N_A_176_987#_c_259_n N_SLEEP_c_707_n 0.00282641f $X=2.32 $Y=4.235
+ $X2=0.615 $Y2=2.23
cc_293 N_A_176_987#_c_258_n N_SLEEP_c_733_n 0.0156707f $X=2.24 $Y=5.355
+ $X2=2.865 $Y2=4.155
cc_294 N_A_176_987#_c_258_n N_SLEEP_c_735_n 0.00148894f $X=2.24 $Y=5.355
+ $X2=2.875 $Y2=3.245
cc_295 N_A_176_987#_c_268_n A_206_1085# 0.00200208f $X=1.165 $Y=5.1 $X2=0.615
+ $Y2=2.23
cc_296 N_A_176_987#_c_265_n N_A_278_1085#_M1019_d 0.00176461f $X=2.155 $Y=5.44
+ $X2=0.615 $Y2=2.23
cc_297 N_A_176_987#_M1020_g N_A_278_1085#_c_853_n 0.00145208f $X=0.955 $Y=5.925
+ $X2=0 $Y2=0
cc_298 N_A_176_987#_M1019_g N_A_278_1085#_c_853_n 0.0102531f $X=1.315 $Y=5.925
+ $X2=0 $Y2=0
cc_299 N_A_176_987#_c_265_n N_A_278_1085#_c_853_n 0.0171383f $X=2.155 $Y=5.44
+ $X2=0 $Y2=0
cc_300 N_A_176_987#_c_267_n N_A_278_1085#_c_853_n 0.0120446f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_301 N_A_176_987#_M1010_d N_A_278_1085#_c_849_n 0.00559995f $X=2.18 $Y=5.425
+ $X2=0 $Y2=0
cc_302 N_A_176_987#_c_267_n N_A_278_1085#_c_849_n 0.019416f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_303 N_A_176_987#_M1020_g N_A_278_1085#_c_859_n 4.5542e-19 $X=0.955 $Y=5.925
+ $X2=0 $Y2=0
cc_304 N_A_176_987#_M1019_g N_A_278_1085#_c_859_n 0.00285177f $X=1.315 $Y=5.925
+ $X2=0 $Y2=0
cc_305 N_A_176_987#_c_267_n N_A_278_1085#_c_851_n 0.0189219f $X=2.32 $Y=5.55
+ $X2=0 $Y2=0
cc_306 N_A_176_987#_c_269_n N_A_278_1085#_c_851_n 0.00227118f $X=2.155 $Y=5.355
+ $X2=0 $Y2=0
cc_307 N_A_176_987#_c_265_n A_364_1085# 0.00366293f $X=2.155 $Y=5.44 $X2=0.615
+ $Y2=2.23
cc_308 N_A_176_987#_M1020_g N_DESTPWR_c_888_n 0.00518588f $X=0.955 $Y=5.925
+ $X2=0 $Y2=0
cc_309 N_A_176_987#_M1019_g N_DESTPWR_c_888_n 0.00547432f $X=1.315 $Y=5.925
+ $X2=0 $Y2=0
cc_310 N_A_176_987#_M1010_d N_DESTPWR_c_885_n 0.00232737f $X=2.18 $Y=5.425
+ $X2=0.24 $Y2=3.855
cc_311 N_A_176_987#_M1020_g N_DESTPWR_c_885_n 0.0103683f $X=0.955 $Y=5.925
+ $X2=0.24 $Y2=3.855
cc_312 N_A_176_987#_M1019_g N_DESTPWR_c_885_n 0.00979813f $X=1.315 $Y=5.925
+ $X2=0.24 $Y2=3.855
cc_313 N_A_176_987#_M1021_d N_A_278_718#_c_1002_n 0.00426626f $X=2.18 $Y=3.59
+ $X2=0 $Y2=0
cc_314 N_A_176_987#_c_259_n N_A_278_718#_c_1002_n 0.0126536f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_315 N_A_176_987#_c_259_n N_A_278_718#_c_1013_n 0.00705761f $X=2.32 $Y=4.235
+ $X2=0 $Y2=0
cc_316 N_A_M1001_g N_A_278_47#_c_410_n 0.0237825f $X=1.315 $Y=4.01 $X2=0 $Y2=0
cc_317 N_A_c_352_n N_A_278_47#_c_413_n 0.00454236f $X=1.315 $Y=3.14 $X2=0 $Y2=0
cc_318 N_A_M1013_g N_A_278_47#_c_432_n 0.00339963f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_319 N_A_M1006_g N_A_278_47#_c_432_n 0.0148505f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_320 N_A_c_352_n N_A_278_47#_c_422_n 0.00346449f $X=1.315 $Y=3.14 $X2=0 $Y2=0
cc_321 N_A_c_362_n N_A_278_47#_c_422_n 0.0154334f $X=1.405 $Y=2.925 $X2=0 $Y2=0
cc_322 N_A_M1012_g N_A_278_47#_c_425_n 0.00232378f $X=1.315 $Y=2.44 $X2=0 $Y2=0
cc_323 N_A_c_352_n N_A_278_47#_c_425_n 3.97765e-19 $X=1.315 $Y=3.14 $X2=0 $Y2=0
cc_324 N_A_c_360_n N_A_278_47#_c_425_n 0.00510196f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_325 N_A_c_362_n N_A_278_47#_c_425_n 0.0247675f $X=1.405 $Y=2.925 $X2=0 $Y2=0
cc_326 N_A_c_352_n N_A_278_47#_c_428_n 0.0171629f $X=1.315 $Y=3.14 $X2=-0.025
+ $Y2=-0.245
cc_327 N_A_c_362_n N_A_278_47#_c_428_n 0.00191938f $X=1.405 $Y=2.925 $X2=-0.025
+ $Y2=-0.245
cc_328 N_A_M1006_g N_A_278_47#_c_433_n 0.00684213f $X=1.315 $Y=0.735 $X2=0.24
+ $Y2=3.245
cc_329 N_A_M1006_g N_A_278_47#_c_431_n 0.0272488f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_330 N_A_c_360_n N_A_278_47#_c_431_n 0.0140219f $X=1.16 $Y=2.775 $X2=0 $Y2=0
cc_331 N_A_c_368_n N_A_278_47#_c_431_n 0.0500336f $X=1.16 $Y=1.832 $X2=0 $Y2=0
cc_332 N_A_M1008_g N_A_123_718#_c_485_n 0.00781951f $X=0.955 $Y=4.01 $X2=-0.025
+ $Y2=-0.245
cc_333 N_A_M1008_g N_A_123_718#_c_488_n 0.00392017f $X=0.955 $Y=4.01 $X2=0.24
+ $Y2=3.855
cc_334 N_A_M1001_g N_A_123_718#_c_488_n 0.00352781f $X=1.315 $Y=4.01 $X2=0.24
+ $Y2=3.855
cc_335 N_A_M1013_g N_VPWR_c_823_n 0.0213886f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_336 N_A_M1006_g N_VPWR_c_823_n 0.00375886f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_337 N_A_c_366_n N_VPWR_c_823_n 0.00119966f $X=1.315 $Y=1.96 $X2=0 $Y2=0
cc_338 N_A_c_368_n N_VPWR_c_823_n 0.0154497f $X=1.16 $Y=1.832 $X2=0 $Y2=0
cc_339 N_A_M1013_g N_VPWR_c_827_n 0.00486043f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_340 N_A_M1006_g N_VPWR_c_827_n 0.00549284f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_341 N_A_M1013_g N_VPWR_c_822_n 0.00814425f $X=0.955 $Y=0.735 $X2=0 $Y2=0
cc_342 N_A_M1006_g N_VPWR_c_822_n 0.0111098f $X=1.315 $Y=0.735 $X2=0 $Y2=0
cc_343 N_A_M1008_g N_A_278_718#_c_1013_n 0.00250397f $X=0.955 $Y=4.01 $X2=0
+ $Y2=0
cc_344 N_A_M1001_g N_A_278_718#_c_1013_n 0.0175796f $X=1.315 $Y=4.01 $X2=0 $Y2=0
cc_345 N_A_278_47#_c_405_n N_A_123_718#_c_476_n 0.006115f $X=1.745 $Y=3.515
+ $X2=0 $Y2=0
cc_346 N_A_278_47#_c_416_n N_A_123_718#_c_476_n 0.00407187f $X=2.105 $Y=3.515
+ $X2=0 $Y2=0
cc_347 N_A_278_47#_c_405_n N_A_123_718#_c_488_n 5.99168e-19 $X=1.745 $Y=3.515
+ $X2=0.24 $Y2=3.855
cc_348 N_A_278_47#_c_405_n N_A_123_718#_c_515_n 8.15435e-19 $X=1.745 $Y=3.515
+ $X2=0 $Y2=0
cc_349 N_A_278_47#_c_428_n N_A_517_420#_c_633_n 0.00490025f $X=1.98 $Y=2.925
+ $X2=0 $Y2=0
cc_350 N_A_278_47#_c_413_n N_A_517_420#_c_641_n 0.00490025f $X=2.07 $Y=3.365
+ $X2=0 $Y2=0
cc_351 N_A_278_47#_c_416_n N_SLEEP_c_733_n 2.77866e-19 $X=2.105 $Y=3.515
+ $X2=2.865 $Y2=4.155
cc_352 N_A_278_47#_c_432_n N_VPWR_c_823_n 0.0305839f $X=1.53 $Y=0.38 $X2=0 $Y2=0
cc_353 N_A_278_47#_c_432_n N_VPWR_c_827_n 0.0211337f $X=1.53 $Y=0.38 $X2=0 $Y2=0
cc_354 N_A_278_47#_M1006_d N_VPWR_c_822_n 0.00215406f $X=1.39 $Y=0.235 $X2=0
+ $Y2=0
cc_355 N_A_278_47#_c_432_n N_VPWR_c_822_n 0.0132819f $X=1.53 $Y=0.38 $X2=0 $Y2=0
cc_356 N_A_278_47#_c_405_n N_A_278_718#_c_1002_n 0.012303f $X=1.745 $Y=3.515
+ $X2=0 $Y2=0
cc_357 N_A_278_47#_c_407_n N_A_278_718#_c_1002_n 5.62214e-19 $X=1.995 $Y=3.44
+ $X2=0 $Y2=0
cc_358 N_A_278_47#_c_416_n N_A_278_718#_c_1002_n 0.0151615f $X=2.105 $Y=3.515
+ $X2=0 $Y2=0
cc_359 N_A_278_47#_c_422_n N_A_278_718#_c_1006_n 0.0144198f $X=1.98 $Y=2.605
+ $X2=0 $Y2=0
cc_360 N_A_278_47#_c_425_n N_A_278_718#_c_1006_n 0.036567f $X=1.98 $Y=2.925
+ $X2=0 $Y2=0
cc_361 N_A_278_47#_c_428_n N_A_278_718#_c_1006_n 0.00279589f $X=1.98 $Y=2.925
+ $X2=0 $Y2=0
cc_362 N_A_278_47#_c_431_n N_A_278_718#_c_1006_n 0.00349796f $X=1.53 $Y=2.44
+ $X2=0 $Y2=0
cc_363 N_A_278_47#_c_413_n N_A_278_718#_c_1007_n 6.18037e-19 $X=2.07 $Y=3.365
+ $X2=0 $Y2=0
cc_364 N_A_278_47#_c_419_n N_A_278_718#_c_1007_n 0.00617354f $X=2.087 $Y=3.44
+ $X2=0 $Y2=0
cc_365 N_A_278_47#_c_405_n N_A_278_718#_c_1013_n 0.00138154f $X=1.745 $Y=3.515
+ $X2=0 $Y2=0
cc_366 N_A_278_47#_c_413_n N_A_278_718#_c_1016_n 0.00279589f $X=2.07 $Y=3.365
+ $X2=0 $Y2=0
cc_367 N_A_123_718#_c_509_n N_A_517_420#_M1015_d 0.00726325f $X=4.7 $Y=6.32
+ $X2=2.735 $Y2=2.23
cc_368 N_A_123_718#_c_506_n N_A_517_420#_c_650_n 0.0264452f $X=3.99 $Y=5.165
+ $X2=0 $Y2=0
cc_369 N_A_123_718#_c_491_n N_A_517_420#_c_650_n 0.0159282f $X=4.87 $Y=4.825
+ $X2=0 $Y2=0
cc_370 N_A_123_718#_c_506_n N_A_517_420#_c_651_n 0.0187956f $X=3.99 $Y=5.165
+ $X2=0 $Y2=0
cc_371 N_A_123_718#_c_506_n N_A_517_420#_c_652_n 0.013514f $X=3.99 $Y=5.165
+ $X2=0 $Y2=0
cc_372 N_A_123_718#_c_508_n N_A_517_420#_c_652_n 0.0335424f $X=4.075 $Y=6.235
+ $X2=0 $Y2=0
cc_373 N_A_123_718#_c_509_n N_A_517_420#_c_652_n 0.0121011f $X=4.7 $Y=6.32 $X2=0
+ $Y2=0
cc_374 N_A_123_718#_c_510_n N_A_517_420#_c_652_n 0.0791492f $X=4.785 $Y=6.235
+ $X2=0 $Y2=0
cc_375 N_A_123_718#_c_491_n N_A_517_420#_c_652_n 0.00679352f $X=4.87 $Y=4.825
+ $X2=0 $Y2=0
cc_376 N_A_123_718#_c_506_n N_SLEEP_M1002_g 0.0185729f $X=3.99 $Y=5.165 $X2=0
+ $Y2=0
cc_377 N_A_123_718#_c_490_n N_SLEEP_M1002_g 8.56956e-19 $X=2.745 $Y=5.165 $X2=0
+ $Y2=0
cc_378 N_A_123_718#_c_495_n N_SLEEP_M1002_g 0.00742904f $X=2.58 $Y=5.1 $X2=0
+ $Y2=0
cc_379 N_A_123_718#_c_506_n N_SLEEP_c_716_n 4.01661e-19 $X=3.99 $Y=5.165 $X2=0
+ $Y2=0
cc_380 N_A_123_718#_c_506_n N_SLEEP_M1005_g 0.0145847f $X=3.99 $Y=5.165 $X2=0
+ $Y2=0
cc_381 N_A_123_718#_c_508_n N_SLEEP_M1005_g 0.00664656f $X=4.075 $Y=6.235 $X2=0
+ $Y2=0
cc_382 N_A_123_718#_c_506_n N_SLEEP_c_719_n 0.0027719f $X=3.99 $Y=5.165 $X2=0
+ $Y2=0
cc_383 N_A_123_718#_c_491_n N_SLEEP_c_719_n 9.63508e-19 $X=4.87 $Y=4.825 $X2=0
+ $Y2=0
cc_384 N_A_123_718#_c_508_n N_SLEEP_c_739_n 0.0151466f $X=4.075 $Y=6.235 $X2=0
+ $Y2=0
cc_385 N_A_123_718#_c_509_n N_SLEEP_c_739_n 0.0137572f $X=4.7 $Y=6.32 $X2=0
+ $Y2=0
cc_386 N_A_123_718#_c_576_p N_SLEEP_c_739_n 0.00110234f $X=4.16 $Y=6.32 $X2=0
+ $Y2=0
cc_387 N_A_123_718#_c_510_n N_SLEEP_c_739_n 0.00372942f $X=4.785 $Y=6.235 $X2=0
+ $Y2=0
cc_388 N_A_123_718#_M1023_g N_SLEEP_c_740_n 0.0806592f $X=5.765 $Y=5.925 $X2=0
+ $Y2=0
cc_389 N_A_123_718#_c_510_n N_SLEEP_c_740_n 0.0178671f $X=4.785 $Y=6.235 $X2=0
+ $Y2=0
cc_390 N_A_123_718#_c_492_n N_SLEEP_c_740_n 0.0120446f $X=5.495 $Y=4.825 $X2=0
+ $Y2=0
cc_391 N_A_123_718#_c_497_n N_SLEEP_c_740_n 0.0112999f $X=5.765 $Y=4.825 $X2=0
+ $Y2=0
cc_392 N_A_123_718#_c_491_n N_SLEEP_c_725_n 0.00259927f $X=4.87 $Y=4.825
+ $X2=0.24 $Y2=3.245
cc_393 N_A_123_718#_c_492_n N_SLEEP_c_725_n 0.00271874f $X=5.495 $Y=4.825
+ $X2=0.24 $Y2=3.245
cc_394 N_A_123_718#_M1011_g N_SLEEP_c_726_n 0.0437228f $X=5.405 $Y=4.01 $X2=0
+ $Y2=0
cc_395 N_A_123_718#_c_510_n N_SLEEP_c_741_n 0.00280665f $X=4.785 $Y=6.235
+ $X2=0.24 $Y2=3.415
cc_396 N_A_123_718#_c_506_n N_SLEEP_c_742_n 0.0012043f $X=3.99 $Y=5.165
+ $X2=0.575 $Y2=3.33
cc_397 N_A_123_718#_c_508_n N_SLEEP_c_742_n 0.00198545f $X=4.075 $Y=6.235
+ $X2=0.575 $Y2=3.33
cc_398 N_A_123_718#_c_506_n N_SLEEP_c_733_n 0.0467041f $X=3.99 $Y=5.165
+ $X2=2.865 $Y2=4.155
cc_399 N_A_123_718#_c_506_n N_SLEEP_c_735_n 0.00224573f $X=3.99 $Y=5.165
+ $X2=2.875 $Y2=3.245
cc_400 N_A_123_718#_c_498_n N_A_278_1085#_c_853_n 0.0106887f $X=1.745 $Y=5.35
+ $X2=0 $Y2=0
cc_401 N_A_123_718#_c_499_n N_A_278_1085#_c_853_n 0.00187953f $X=2.105 $Y=5.35
+ $X2=0 $Y2=0
cc_402 N_A_123_718#_c_504_n N_A_278_1085#_c_853_n 0.0188335f $X=0.74 $Y=6.28
+ $X2=0 $Y2=0
cc_403 N_A_123_718#_c_498_n N_A_278_1085#_c_849_n 0.010046f $X=1.745 $Y=5.35
+ $X2=0 $Y2=0
cc_404 N_A_123_718#_c_499_n N_A_278_1085#_c_849_n 0.0151541f $X=2.105 $Y=5.35
+ $X2=0 $Y2=0
cc_405 N_A_123_718#_c_498_n N_A_278_1085#_c_859_n 5.81207e-19 $X=1.745 $Y=5.35
+ $X2=0 $Y2=0
cc_406 N_A_123_718#_c_504_n N_A_278_1085#_c_859_n 0.00629328f $X=0.74 $Y=6.28
+ $X2=0 $Y2=0
cc_407 N_A_123_718#_c_506_n N_A_278_1085#_c_851_n 0.0205931f $X=3.99 $Y=5.165
+ $X2=0 $Y2=0
cc_408 N_A_123_718#_c_506_n N_DESTPWR_c_886_n 0.0141894f $X=3.99 $Y=5.165 $X2=0
+ $Y2=0
cc_409 N_A_123_718#_c_508_n N_DESTPWR_c_886_n 2.29837e-19 $X=4.075 $Y=6.235
+ $X2=0 $Y2=0
cc_410 N_A_123_718#_M1023_g N_DESTPWR_c_887_n 0.00390966f $X=5.765 $Y=5.925
+ $X2=0 $Y2=0
cc_411 N_A_123_718#_c_509_n N_DESTPWR_c_887_n 0.0149884f $X=4.7 $Y=6.32 $X2=0
+ $Y2=0
cc_412 N_A_123_718#_c_510_n N_DESTPWR_c_887_n 0.0643412f $X=4.785 $Y=6.235 $X2=0
+ $Y2=0
cc_413 N_A_123_718#_c_492_n N_DESTPWR_c_887_n 0.0142746f $X=5.495 $Y=4.825 $X2=0
+ $Y2=0
cc_414 N_A_123_718#_c_498_n N_DESTPWR_c_888_n 0.00357842f $X=1.745 $Y=5.35 $X2=0
+ $Y2=0
cc_415 N_A_123_718#_c_499_n N_DESTPWR_c_888_n 0.00357877f $X=2.105 $Y=5.35 $X2=0
+ $Y2=0
cc_416 N_A_123_718#_c_504_n N_DESTPWR_c_888_n 0.0224101f $X=0.74 $Y=6.28 $X2=0
+ $Y2=0
cc_417 N_A_123_718#_c_509_n N_DESTPWR_c_890_n 0.0445984f $X=4.7 $Y=6.32 $X2=0
+ $Y2=0
cc_418 N_A_123_718#_c_576_p N_DESTPWR_c_890_n 0.00950638f $X=4.16 $Y=6.32 $X2=0
+ $Y2=0
cc_419 N_A_123_718#_M1023_g N_DESTPWR_c_891_n 0.0054895f $X=5.765 $Y=5.925
+ $X2=0.24 $Y2=3.415
cc_420 N_A_123_718#_M1020_s N_DESTPWR_c_885_n 0.00215158f $X=0.615 $Y=5.425
+ $X2=0.24 $Y2=3.855
cc_421 N_A_123_718#_c_498_n N_DESTPWR_c_885_n 0.00516571f $X=1.745 $Y=5.35
+ $X2=0.24 $Y2=3.855
cc_422 N_A_123_718#_c_499_n N_DESTPWR_c_885_n 0.0066108f $X=2.105 $Y=5.35
+ $X2=0.24 $Y2=3.855
cc_423 N_A_123_718#_M1023_g N_DESTPWR_c_885_n 0.0111524f $X=5.765 $Y=5.925
+ $X2=0.24 $Y2=3.855
cc_424 N_A_123_718#_c_504_n N_DESTPWR_c_885_n 0.0132444f $X=0.74 $Y=6.28
+ $X2=0.24 $Y2=3.855
cc_425 N_A_123_718#_c_509_n N_DESTPWR_c_885_n 0.0262447f $X=4.7 $Y=6.32 $X2=0.24
+ $Y2=3.855
cc_426 N_A_123_718#_c_576_p N_DESTPWR_c_885_n 0.00657636f $X=4.16 $Y=6.32
+ $X2=0.24 $Y2=3.855
cc_427 N_A_123_718#_c_576_p A_789_1085# 9.38685e-19 $X=4.16 $Y=6.32 $X2=0.615
+ $Y2=2.23
cc_428 N_A_123_718#_M1011_g N_X_c_958_n 0.0140172f $X=5.405 $Y=4.01 $X2=0 $Y2=0
cc_429 N_A_123_718#_M1004_g N_X_c_958_n 0.0144626f $X=5.765 $Y=4.01 $X2=0 $Y2=0
cc_430 N_A_123_718#_c_491_n N_X_c_958_n 0.0143516f $X=4.87 $Y=4.825 $X2=0 $Y2=0
cc_431 N_A_123_718#_c_492_n N_X_c_958_n 0.0540891f $X=5.495 $Y=4.825 $X2=0 $Y2=0
cc_432 N_A_123_718#_c_497_n N_X_c_958_n 9.75531e-19 $X=5.765 $Y=4.825 $X2=0
+ $Y2=0
cc_433 N_A_123_718#_M1004_g X 0.00158184f $X=5.765 $Y=4.01 $X2=0 $Y2=0
cc_434 N_A_123_718#_M1011_g X 8.44505e-19 $X=5.405 $Y=4.01 $X2=0 $Y2=0
cc_435 N_A_123_718#_M1004_g X 0.00631209f $X=5.765 $Y=4.01 $X2=0 $Y2=0
cc_436 N_A_123_718#_M1023_g X 0.0375216f $X=5.765 $Y=5.925 $X2=0 $Y2=0
cc_437 N_A_123_718#_c_492_n X 0.0201866f $X=5.495 $Y=4.825 $X2=0 $Y2=0
cc_438 N_A_123_718#_c_497_n X 0.0128845f $X=5.765 $Y=4.825 $X2=0 $Y2=0
cc_439 N_A_123_718#_M1011_g N_X_c_964_n 0.00300668f $X=5.405 $Y=4.01 $X2=0.24
+ $Y2=3.245
cc_440 N_A_123_718#_M1004_g N_X_c_964_n 0.0157235f $X=5.765 $Y=4.01 $X2=0.24
+ $Y2=3.245
cc_441 N_A_123_718#_c_485_n N_A_278_718#_c_1013_n 0.0147015f $X=0.74 $Y=3.75
+ $X2=0 $Y2=0
cc_442 N_A_123_718#_c_488_n N_A_278_718#_c_1013_n 0.0239528f $X=1.52 $Y=4.735
+ $X2=0 $Y2=0
cc_443 N_A_517_420#_c_636_n N_SLEEP_c_707_n 0.0024026f $X=3.83 $Y=3.22 $X2=0.615
+ $Y2=2.23
cc_444 N_A_517_420#_c_645_n N_SLEEP_c_707_n 9.80946e-19 $X=3.702 $Y=4.24
+ $X2=0.615 $Y2=2.23
cc_445 N_A_517_420#_c_636_n N_SLEEP_c_711_n 0.00239275f $X=3.83 $Y=3.22 $X2=5.05
+ $Y2=3.59
cc_446 N_A_517_420#_c_645_n N_SLEEP_c_711_n 0.00974027f $X=3.702 $Y=4.24
+ $X2=5.05 $Y2=3.59
cc_447 N_A_517_420#_c_649_n N_SLEEP_c_711_n 0.00830112f $X=3.702 $Y=4.74
+ $X2=5.05 $Y2=3.59
cc_448 N_A_517_420#_c_653_n N_SLEEP_c_711_n 0.00135899f $X=3.995 $Y=3.75
+ $X2=5.05 $Y2=3.59
cc_449 N_A_517_420#_c_649_n N_SLEEP_c_716_n 0.011511f $X=3.702 $Y=4.74 $X2=0
+ $Y2=0
cc_450 N_A_517_420#_c_649_n N_SLEEP_M1005_g 0.00207384f $X=3.702 $Y=4.74 $X2=0
+ $Y2=0
cc_451 N_A_517_420#_c_650_n N_SLEEP_M1005_g 0.0102332f $X=4.33 $Y=4.825 $X2=0
+ $Y2=0
cc_452 N_A_517_420#_c_651_n N_SLEEP_M1005_g 0.00206052f $X=3.815 $Y=4.825 $X2=0
+ $Y2=0
cc_453 N_A_517_420#_c_652_n N_SLEEP_M1005_g 2.44465e-19 $X=4.445 $Y=5.55 $X2=0
+ $Y2=0
cc_454 N_A_517_420#_c_650_n N_SLEEP_c_718_n 0.00112662f $X=4.33 $Y=4.825 $X2=0
+ $Y2=0
cc_455 N_A_517_420#_c_649_n N_SLEEP_c_719_n 4.83723e-19 $X=3.702 $Y=4.74 $X2=0
+ $Y2=0
cc_456 N_A_517_420#_c_650_n N_SLEEP_c_719_n 0.0187948f $X=4.33 $Y=4.825 $X2=0
+ $Y2=0
cc_457 N_A_517_420#_c_652_n N_SLEEP_c_719_n 0.00761657f $X=4.445 $Y=5.55 $X2=0
+ $Y2=0
cc_458 N_A_517_420#_c_652_n N_SLEEP_c_739_n 0.00169277f $X=4.445 $Y=5.55 $X2=0
+ $Y2=0
cc_459 N_A_517_420#_c_650_n N_SLEEP_c_720_n 0.00290535f $X=4.33 $Y=4.825 $X2=0
+ $Y2=0
cc_460 N_A_517_420#_c_650_n N_SLEEP_c_740_n 5.28578e-19 $X=4.33 $Y=4.825 $X2=0
+ $Y2=0
cc_461 N_A_517_420#_c_652_n N_SLEEP_c_740_n 0.013374f $X=4.445 $Y=5.55 $X2=0
+ $Y2=0
cc_462 N_A_517_420#_c_653_n N_SLEEP_c_721_n 0.00431241f $X=3.995 $Y=3.75 $X2=0
+ $Y2=0
cc_463 N_A_517_420#_c_656_n N_SLEEP_c_721_n 0.00277014f $X=3.995 $Y=3.585 $X2=0
+ $Y2=0
cc_464 N_A_517_420#_c_645_n N_SLEEP_c_730_n 0.00197198f $X=3.702 $Y=4.24 $X2=0
+ $Y2=0
cc_465 N_A_517_420#_c_649_n N_SLEEP_c_730_n 0.00759926f $X=3.702 $Y=4.74 $X2=0
+ $Y2=0
cc_466 N_A_517_420#_c_653_n N_SLEEP_c_730_n 0.00660115f $X=3.995 $Y=3.75 $X2=0
+ $Y2=0
cc_467 N_A_517_420#_c_649_n N_SLEEP_c_733_n 0.0182428f $X=3.702 $Y=4.74
+ $X2=2.865 $Y2=4.155
cc_468 N_A_517_420#_c_651_n N_SLEEP_c_733_n 0.014862f $X=3.815 $Y=4.825
+ $X2=2.865 $Y2=4.155
cc_469 N_A_517_420#_c_649_n N_SLEEP_c_735_n 6.91261e-19 $X=3.702 $Y=4.74
+ $X2=2.875 $Y2=3.245
cc_470 N_A_517_420#_c_651_n N_SLEEP_c_735_n 0.00150219f $X=3.815 $Y=4.825
+ $X2=2.875 $Y2=3.245
cc_471 N_A_517_420#_M1015_d N_DESTPWR_c_885_n 0.00232737f $X=4.305 $Y=5.425
+ $X2=0.24 $Y2=3.855
cc_472 N_A_517_420#_c_645_n N_X_c_954_n 0.0354593f $X=3.702 $Y=4.24 $X2=0 $Y2=0
cc_473 N_A_517_420#_c_649_n N_X_c_954_n 0.00299499f $X=3.702 $Y=4.74 $X2=0 $Y2=0
cc_474 N_A_517_420#_c_653_n N_X_c_954_n 0.00288777f $X=3.995 $Y=3.75 $X2=0 $Y2=0
cc_475 N_A_517_420#_c_649_n N_X_c_961_n 0.00701637f $X=3.702 $Y=4.74 $X2=0 $Y2=0
cc_476 N_A_517_420#_c_650_n N_X_c_961_n 0.0170557f $X=4.33 $Y=4.825 $X2=0 $Y2=0
cc_477 N_A_517_420#_c_633_n N_A_278_718#_c_1007_n 0.00165736f $X=2.66 $Y=3.145
+ $X2=0 $Y2=0
cc_478 N_A_517_420#_c_633_n N_A_278_718#_c_1016_n 9.27717e-19 $X=2.66 $Y=3.145
+ $X2=0 $Y2=0
cc_479 N_SLEEP_M1002_g N_A_278_1085#_c_850_n 0.00197018f $X=3.44 $Y=5.925 $X2=0
+ $Y2=0
cc_480 N_SLEEP_M1002_g N_A_278_1085#_c_851_n 0.00832486f $X=3.44 $Y=5.925 $X2=0
+ $Y2=0
cc_481 N_SLEEP_M1002_g N_DESTPWR_c_886_n 0.00281775f $X=3.44 $Y=5.925 $X2=0
+ $Y2=0
cc_482 N_SLEEP_M1005_g N_DESTPWR_c_886_n 0.00275486f $X=3.87 $Y=5.925 $X2=0
+ $Y2=0
cc_483 N_SLEEP_c_740_n N_DESTPWR_c_887_n 0.00543646f $X=5.33 $Y=5.275 $X2=0
+ $Y2=0
cc_484 N_SLEEP_c_741_n N_DESTPWR_c_887_n 0.0222504f $X=5.405 $Y=5.35 $X2=0 $Y2=0
cc_485 N_SLEEP_M1002_g N_DESTPWR_c_888_n 0.00547432f $X=3.44 $Y=5.925 $X2=0
+ $Y2=0
cc_486 N_SLEEP_M1005_g N_DESTPWR_c_890_n 0.00585385f $X=3.87 $Y=5.925 $X2=0
+ $Y2=0
cc_487 N_SLEEP_c_739_n N_DESTPWR_c_890_n 0.0035787f $X=4.23 $Y=5.35 $X2=0 $Y2=0
cc_488 N_SLEEP_c_741_n N_DESTPWR_c_891_n 0.00486043f $X=5.405 $Y=5.35 $X2=0.24
+ $Y2=3.415
cc_489 N_SLEEP_M1002_g N_DESTPWR_c_885_n 0.0110556f $X=3.44 $Y=5.925 $X2=0.24
+ $Y2=3.855
cc_490 N_SLEEP_M1005_g N_DESTPWR_c_885_n 0.0105424f $X=3.87 $Y=5.925 $X2=0.24
+ $Y2=3.855
cc_491 N_SLEEP_c_739_n N_DESTPWR_c_885_n 0.00661079f $X=4.23 $Y=5.35 $X2=0.24
+ $Y2=3.855
cc_492 N_SLEEP_c_741_n N_DESTPWR_c_885_n 0.00818711f $X=5.405 $Y=5.35 $X2=0.24
+ $Y2=3.855
cc_493 N_SLEEP_c_721_n N_X_c_954_n 0.0130481f $X=4.615 $Y=4.505 $X2=0 $Y2=0
cc_494 N_SLEEP_c_726_n N_X_c_954_n 0.0029998f $X=4.975 $Y=4.505 $X2=0 $Y2=0
cc_495 N_SLEEP_c_721_n N_X_c_958_n 0.0137628f $X=4.615 $Y=4.505 $X2=0 $Y2=0
cc_496 N_SLEEP_c_725_n N_X_c_958_n 6.90929e-19 $X=4.9 $Y=4.58 $X2=0 $Y2=0
cc_497 N_SLEEP_c_726_n N_X_c_958_n 0.0133831f $X=4.975 $Y=4.505 $X2=0 $Y2=0
cc_498 N_SLEEP_c_721_n N_X_c_961_n 0.00366132f $X=4.615 $Y=4.505 $X2=0 $Y2=0
cc_499 N_SLEEP_c_731_n N_X_c_961_n 0.00443951f $X=4.23 $Y=4.58 $X2=0 $Y2=0
cc_500 N_SLEEP_c_740_n X 0.00390383f $X=5.33 $Y=5.275 $X2=0 $Y2=0
cc_501 N_VPWR_c_822_n A_206_47# 0.00899413f $X=6.48 $Y=0 $X2=0.615 $Y2=2.23
cc_502 A_206_1085# N_DESTPWR_c_885_n 0.00899413f $X=1.03 $Y=5.425 $X2=0 $Y2=0
cc_503 N_A_278_1085#_c_849_n A_364_1085# 0.00456442f $X=3.06 $Y=6.32 $X2=0.155
+ $Y2=5.495
cc_504 N_A_278_1085#_c_849_n N_DESTPWR_c_888_n 0.0817564f $X=3.06 $Y=6.32
+ $X2=0.24 $Y2=5.365
cc_505 N_A_278_1085#_c_859_n N_DESTPWR_c_888_n 0.019107f $X=1.695 $Y=6.32
+ $X2=0.24 $Y2=5.365
cc_506 N_A_278_1085#_c_850_n N_DESTPWR_c_888_n 0.0211797f $X=3.225 $Y=6.235
+ $X2=0.24 $Y2=5.365
cc_507 N_A_278_1085#_M1019_d N_DESTPWR_c_885_n 0.00223559f $X=1.39 $Y=5.425
+ $X2=0 $Y2=0
cc_508 N_A_278_1085#_M1002_s N_DESTPWR_c_885_n 0.00219347f $X=3.095 $Y=5.425
+ $X2=0 $Y2=0
cc_509 N_A_278_1085#_c_849_n N_DESTPWR_c_885_n 0.0500621f $X=3.06 $Y=6.32 $X2=0
+ $Y2=0
cc_510 N_A_278_1085#_c_859_n N_DESTPWR_c_885_n 0.0124689f $X=1.695 $Y=6.32 $X2=0
+ $Y2=0
cc_511 N_A_278_1085#_c_850_n N_DESTPWR_c_885_n 0.0126421f $X=3.225 $Y=6.235
+ $X2=0 $Y2=0
cc_512 A_364_1085# N_DESTPWR_c_885_n 0.00168889f $X=1.82 $Y=5.425 $X2=0 $Y2=0
cc_513 N_DESTPWR_c_885_n A_789_1085# 0.00325419f $X=6.48 $Y=6.66 $X2=0.615
+ $Y2=2.23
cc_514 N_DESTPWR_c_885_n A_1096_1085# 0.00899413f $X=6.48 $Y=6.66 $X2=0.615
+ $Y2=2.23
cc_515 N_DESTPWR_c_885_n N_X_M1023_d 0.00215158f $X=6.48 $Y=6.66 $X2=2.74
+ $Y2=4.01
cc_516 N_DESTPWR_c_887_n X 0.0328385f $X=5.19 $Y=5.585 $X2=0 $Y2=0
cc_517 N_DESTPWR_c_891_n X 0.0210467f $X=6.48 $Y=6.66 $X2=0 $Y2=0
cc_518 N_DESTPWR_c_885_n X 0.0125689f $X=6.48 $Y=6.66 $X2=0 $Y2=0
cc_519 N_X_c_958_n A_938_718# 0.00366293f $X=5.815 $Y=4.405 $X2=0.615 $Y2=2.23
cc_520 N_X_c_958_n A_1096_718# 0.00366293f $X=5.815 $Y=4.405 $X2=0.615 $Y2=2.23
cc_521 N_A_278_718#_c_1002_n A_364_718# 0.00366293f $X=2.315 $Y=3.67 $X2=0.615
+ $Y2=2.23
