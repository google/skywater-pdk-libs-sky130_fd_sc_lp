# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o41a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o41a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.395000 1.210000 7.595000 1.435000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.345000 1.210000 6.225000 1.435000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985000 1.210000 5.175000 1.435000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.455000 1.210000 3.815000 1.435000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.690000 1.210000 3.285000 1.435000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 1.660000 1.225000 ;
        RECT 0.085000 1.225000 0.335000 1.755000 ;
        RECT 0.085000 1.755000 1.660000 1.925000 ;
        RECT 0.610000 0.255000 0.800000 1.055000 ;
        RECT 0.610000 1.925000 0.800000 3.075000 ;
        RECT 1.470000 0.255000 1.660000 1.055000 ;
        RECT 1.470000 1.925000 1.660000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.110000  0.085000 0.440000 0.885000 ;
      RECT 0.110000  2.095000 0.440000 3.245000 ;
      RECT 0.505000  1.395000 2.510000 1.585000 ;
      RECT 0.970000  0.085000 1.300000 0.885000 ;
      RECT 0.970000  2.105000 1.300000 3.245000 ;
      RECT 1.830000  0.085000 2.150000 1.105000 ;
      RECT 1.830000  1.815000 2.160000 3.245000 ;
      RECT 2.320000  0.860000 3.120000 1.040000 ;
      RECT 2.320000  1.040000 2.510000 1.395000 ;
      RECT 2.330000  1.585000 2.510000 1.605000 ;
      RECT 2.330000  1.605000 3.910000 1.815000 ;
      RECT 2.330000  1.815000 2.520000 3.075000 ;
      RECT 2.360000  0.255000 3.515000 0.425000 ;
      RECT 2.360000  0.425000 2.620000 0.690000 ;
      RECT 2.690000  1.985000 3.020000 3.245000 ;
      RECT 2.790000  0.595000 3.120000 0.860000 ;
      RECT 3.220000  1.985000 3.550000 2.905000 ;
      RECT 3.220000  2.905000 4.410000 3.075000 ;
      RECT 3.290000  0.425000 3.515000 0.870000 ;
      RECT 3.290000  0.870000 7.500000 1.040000 ;
      RECT 3.685000  0.085000 3.945000 0.700000 ;
      RECT 3.720000  1.815000 3.910000 2.735000 ;
      RECT 4.080000  1.605000 5.270000 1.775000 ;
      RECT 4.080000  1.775000 4.410000 2.905000 ;
      RECT 4.115000  0.255000 4.375000 0.870000 ;
      RECT 4.545000  0.085000 4.800000 0.700000 ;
      RECT 4.580000  1.945000 4.770000 2.895000 ;
      RECT 4.580000  2.895000 6.260000 3.075000 ;
      RECT 4.940000  1.775000 5.270000 2.725000 ;
      RECT 4.970000  0.255000 5.235000 0.870000 ;
      RECT 5.405000  0.085000 6.150000 0.700000 ;
      RECT 5.500000  1.705000 7.490000 1.875000 ;
      RECT 5.500000  1.875000 5.760000 2.725000 ;
      RECT 5.930000  2.055000 6.260000 2.895000 ;
      RECT 6.320000  0.255000 6.585000 0.870000 ;
      RECT 6.430000  1.875000 6.620000 3.075000 ;
      RECT 6.755000  0.085000 7.015000 0.700000 ;
      RECT 6.790000  2.105000 7.120000 3.245000 ;
      RECT 7.185000  0.265000 7.500000 0.870000 ;
      RECT 7.290000  1.875000 7.490000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__o41a_4
