* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_27_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_726_47# A2 a_919_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_27_367# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_110_47# B1 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND B1 a_110_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_27_367# B1 a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_919_67# A1 a_110_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_110_47# A1 a_919_67# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_919_67# A2 a_726_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VGND A3 a_726_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_726_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VPWR A1 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_27_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR A2 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_110_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 VPWR A3 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
