* File: sky130_fd_sc_lp__a311oi_lp.pxi.spice
* Created: Wed Sep  2 09:25:59 2020
* 
x_PM_SKY130_FD_SC_LP__A311OI_LP%A1 N_A1_c_78_n N_A1_M1001_g N_A1_M1006_g
+ N_A1_c_75_n A1 N_A1_c_76_n N_A1_c_77_n PM_SKY130_FD_SC_LP__A311OI_LP%A1
x_PM_SKY130_FD_SC_LP__A311OI_LP%A2 N_A2_M1003_g N_A2_M1005_g A2 A2 N_A2_c_109_n
+ N_A2_c_110_n PM_SKY130_FD_SC_LP__A311OI_LP%A2
x_PM_SKY130_FD_SC_LP__A311OI_LP%A3 N_A3_M1002_g N_A3_M1000_g N_A3_c_157_n
+ N_A3_c_161_n A3 A3 N_A3_c_159_n PM_SKY130_FD_SC_LP__A311OI_LP%A3
x_PM_SKY130_FD_SC_LP__A311OI_LP%B1 N_B1_c_200_n N_B1_M1009_g N_B1_c_201_n
+ N_B1_c_202_n N_B1_c_203_n N_B1_M1007_g N_B1_c_209_n N_B1_M1008_g N_B1_c_204_n
+ N_B1_c_205_n N_B1_c_206_n B1 B1 N_B1_c_208_n PM_SKY130_FD_SC_LP__A311OI_LP%B1
x_PM_SKY130_FD_SC_LP__A311OI_LP%C1 N_C1_c_265_n N_C1_M1010_g N_C1_c_271_n
+ N_C1_M1004_g N_C1_c_266_n N_C1_M1011_g N_C1_c_267_n N_C1_c_272_n C1
+ N_C1_c_268_n N_C1_c_269_n N_C1_c_270_n PM_SKY130_FD_SC_LP__A311OI_LP%C1
x_PM_SKY130_FD_SC_LP__A311OI_LP%VPWR N_VPWR_M1001_s N_VPWR_M1005_d
+ N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n VPWR
+ N_VPWR_c_323_n N_VPWR_c_318_n N_VPWR_c_325_n
+ PM_SKY130_FD_SC_LP__A311OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A311OI_LP%A_134_409# N_A_134_409#_M1001_d
+ N_A_134_409#_M1000_d N_A_134_409#_c_355_n N_A_134_409#_c_356_n
+ N_A_134_409#_c_357_n N_A_134_409#_c_358_n
+ PM_SKY130_FD_SC_LP__A311OI_LP%A_134_409#
x_PM_SKY130_FD_SC_LP__A311OI_LP%Y N_Y_M1006_s N_Y_M1007_d N_Y_M1004_d
+ N_Y_c_401_n N_Y_c_390_n N_Y_c_391_n N_Y_c_392_n N_Y_c_428_n N_Y_c_398_n
+ N_Y_c_393_n N_Y_c_394_n N_Y_c_399_n N_Y_c_395_n Y N_Y_c_396_n N_Y_c_397_n
+ PM_SKY130_FD_SC_LP__A311OI_LP%Y
x_PM_SKY130_FD_SC_LP__A311OI_LP%VGND N_VGND_M1002_d N_VGND_M1011_d
+ N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n
+ VGND N_VGND_c_486_n N_VGND_c_487_n PM_SKY130_FD_SC_LP__A311OI_LP%VGND
cc_1 VNB N_A1_M1006_g 0.0255309f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.445
cc_2 VNB N_A1_c_75_n 0.038127f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.9
cc_3 VNB N_A1_c_76_n 0.0341614f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.975
cc_4 VNB N_A1_c_77_n 0.0182528f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.975
cc_5 VNB N_A2_M1003_g 0.0527739f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.025
cc_6 VNB N_A2_c_109_n 0.0172404f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.975
cc_7 VNB N_A2_c_110_n 0.018242f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.81
cc_8 VNB N_A3_M1002_g 0.0352083f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.025
cc_9 VNB N_A3_c_157_n 0.0334708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A3 0.00341007f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.81
cc_11 VNB N_A3_c_159_n 0.0264118f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.975
cc_12 VNB N_B1_c_200_n 0.0137255f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.14
cc_13 VNB N_B1_c_201_n 0.00994843f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_14 VNB N_B1_c_202_n 0.00739473f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_15 VNB N_B1_c_203_n 0.0135266f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.81
cc_16 VNB N_B1_c_204_n 0.0178702f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.81
cc_17 VNB N_B1_c_205_n 0.0225419f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.14
cc_18 VNB N_B1_c_206_n 0.00437176f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.975
cc_19 VNB B1 0.00167457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_208_n 0.0166342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C1_c_265_n 0.0157123f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.14
cc_22 VNB N_C1_c_266_n 0.0216315f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_23 VNB N_C1_c_267_n 0.0245474f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.14
cc_24 VNB N_C1_c_268_n 0.0252146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C1_c_269_n 0.00395983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C1_c_270_n 0.025537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_318_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_390_n 0.00155664f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.975
cc_29 VNB N_Y_c_391_n 0.0189612f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.975
cc_30 VNB N_Y_c_392_n 0.00197331f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.975
cc_31 VNB N_Y_c_393_n 0.0141788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_394_n 0.00659774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_395_n 0.0306421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_396_n 0.00888417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_397_n 0.0155399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_481_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_482_n 0.0109794f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_38 VNB N_VGND_c_483_n 0.0177348f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.975
cc_39 VNB N_VGND_c_484_n 0.0375543f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=0.81
cc_40 VNB N_VGND_c_485_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.14
cc_41 VNB N_VGND_c_486_n 0.0345943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_487_n 0.189739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A1_c_78_n 0.0330309f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.025
cc_44 VPB N_A1_c_75_n 0.0159859f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.9
cc_45 VPB N_A2_M1005_g 0.0288608f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.445
cc_46 VPB N_A2_c_109_n 0.0148386f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.975
cc_47 VPB N_A2_c_110_n 0.0151982f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.81
cc_48 VPB N_A3_M1000_g 0.0286439f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.445
cc_49 VPB N_A3_c_161_n 0.0126695f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.975
cc_50 VPB A3 0.00236586f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.81
cc_51 VPB N_A3_c_159_n 0.0012012f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.975
cc_52 VPB N_B1_c_209_n 0.0138955f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_53 VPB N_B1_M1008_g 0.029037f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.975
cc_54 VPB N_B1_c_205_n 0.00134252f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.14
cc_55 VPB B1 0.00195814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_C1_c_271_n 0.0291324f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.445
cc_57 VPB N_C1_c_272_n 0.0138546f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_C1_c_268_n 0.00482861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_C1_c_269_n 0.00493212f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_319_n 0.0113568f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.445
cc_61 VPB N_VPWR_c_320_n 0.0473652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_321_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.975
cc_63 VPB N_VPWR_c_322_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.14
cc_64 VPB N_VPWR_c_323_n 0.0532502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_318_n 0.0640245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_325_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_134_409#_c_355_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_68 VPB N_A_134_409#_c_356_n 0.0164824f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.975
cc_69 VPB N_A_134_409#_c_357_n 0.00229072f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=0.975
cc_70 VPB N_A_134_409#_c_358_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_Y_c_398_n 0.0390561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_Y_c_399_n 0.0180592f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_Y_c_395_n 0.0184462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 N_A1_M1006_g N_A2_M1003_g 0.0555789f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A1_c_75_n N_A2_M1003_g 0.0285982f $X=0.545 $Y=1.9 $X2=0 $Y2=0
cc_76 N_A1_c_77_n N_A2_M1003_g 0.00116895f $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_77 N_A1_c_78_n N_A2_M1005_g 0.0141135f $X=0.545 $Y=2.025 $X2=0 $Y2=0
cc_78 N_A1_c_75_n N_A2_M1005_g 0.00236504f $X=0.545 $Y=1.9 $X2=0 $Y2=0
cc_79 N_A1_c_75_n N_A2_c_109_n 0.00714727f $X=0.545 $Y=1.9 $X2=0 $Y2=0
cc_80 N_A1_c_78_n N_A2_c_110_n 0.00451642f $X=0.545 $Y=2.025 $X2=0 $Y2=0
cc_81 N_A1_c_75_n N_A2_c_110_n 0.0246604f $X=0.545 $Y=1.9 $X2=0 $Y2=0
cc_82 N_A1_c_76_n N_A2_c_110_n 0.00361447f $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_83 N_A1_c_77_n N_A2_c_110_n 0.0200978f $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_84 N_A1_c_78_n N_VPWR_c_320_n 0.0236653f $X=0.545 $Y=2.025 $X2=0 $Y2=0
cc_85 N_A1_c_78_n N_VPWR_c_321_n 0.00769046f $X=0.545 $Y=2.025 $X2=0 $Y2=0
cc_86 N_A1_c_78_n N_VPWR_c_322_n 8.50498e-19 $X=0.545 $Y=2.025 $X2=0 $Y2=0
cc_87 N_A1_c_78_n N_VPWR_c_318_n 0.0134474f $X=0.545 $Y=2.025 $X2=0 $Y2=0
cc_88 N_A1_c_78_n N_A_134_409#_c_355_n 0.0157118f $X=0.545 $Y=2.025 $X2=0 $Y2=0
cc_89 N_A1_c_78_n N_A_134_409#_c_357_n 0.00367688f $X=0.545 $Y=2.025 $X2=0 $Y2=0
cc_90 N_A1_M1006_g N_Y_c_401_n 0.00811163f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A1_c_77_n N_Y_c_401_n 0.00823421f $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_92 N_A1_M1006_g N_Y_c_390_n 0.00360117f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A1_c_77_n N_Y_c_390_n 6.30874e-19 $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_94 N_A1_c_76_n N_Y_c_392_n 6.69696e-19 $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_95 N_A1_c_77_n N_Y_c_392_n 0.0141042f $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_96 N_A1_M1006_g N_Y_c_393_n 0.00486538f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A1_c_76_n N_Y_c_393_n 0.00397641f $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_98 N_A1_c_77_n N_Y_c_393_n 0.0220874f $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_99 N_A1_M1006_g N_VGND_c_484_n 0.00392332f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A1_M1006_g N_VGND_c_487_n 0.00654883f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A1_c_77_n N_VGND_c_487_n 7.52054e-19 $X=0.415 $Y=0.975 $X2=0 $Y2=0
cc_102 N_A2_M1003_g N_A3_M1002_g 0.0635831f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_103 N_A2_M1005_g N_A3_M1000_g 0.0280068f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_104 N_A2_M1003_g A3 0.00174528f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A2_c_109_n A3 4.12603e-19 $X=1.045 $Y=1.675 $X2=0 $Y2=0
cc_106 N_A2_c_110_n A3 0.0222637f $X=1.045 $Y=1.675 $X2=0 $Y2=0
cc_107 N_A2_M1003_g N_A3_c_159_n 0.00699895f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A2_c_109_n N_A3_c_159_n 0.0207596f $X=1.045 $Y=1.675 $X2=0 $Y2=0
cc_109 N_A2_c_110_n N_A3_c_159_n 0.00113718f $X=1.045 $Y=1.675 $X2=0 $Y2=0
cc_110 N_A2_M1005_g N_VPWR_c_320_n 9.44933e-19 $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_111 N_A2_c_110_n N_VPWR_c_320_n 0.0263685f $X=1.045 $Y=1.675 $X2=0 $Y2=0
cc_112 N_A2_M1005_g N_VPWR_c_321_n 0.00769046f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_113 N_A2_M1005_g N_VPWR_c_322_n 0.016528f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_114 N_A2_M1005_g N_VPWR_c_318_n 0.0134474f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_115 N_A2_M1005_g N_A_134_409#_c_355_n 0.0157714f $X=1.075 $Y=2.545 $X2=0
+ $Y2=0
cc_116 N_A2_M1005_g N_A_134_409#_c_356_n 0.0179769f $X=1.075 $Y=2.545 $X2=0
+ $Y2=0
cc_117 N_A2_c_109_n N_A_134_409#_c_356_n 2.22766e-19 $X=1.045 $Y=1.675 $X2=0
+ $Y2=0
cc_118 N_A2_c_110_n N_A_134_409#_c_356_n 0.0160355f $X=1.045 $Y=1.675 $X2=0
+ $Y2=0
cc_119 N_A2_M1005_g N_A_134_409#_c_357_n 0.00104211f $X=1.075 $Y=2.545 $X2=0
+ $Y2=0
cc_120 N_A2_c_109_n N_A_134_409#_c_357_n 0.0022054f $X=1.045 $Y=1.675 $X2=0
+ $Y2=0
cc_121 N_A2_c_110_n N_A_134_409#_c_357_n 0.0274076f $X=1.045 $Y=1.675 $X2=0
+ $Y2=0
cc_122 N_A2_M1005_g N_A_134_409#_c_358_n 8.9791e-19 $X=1.075 $Y=2.545 $X2=0
+ $Y2=0
cc_123 N_A2_M1003_g N_Y_c_401_n 0.00711998f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A2_M1003_g N_Y_c_390_n 0.00507444f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A2_M1003_g N_Y_c_391_n 0.00423625f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A2_c_109_n N_Y_c_391_n 0.00475432f $X=1.045 $Y=1.675 $X2=0 $Y2=0
cc_127 N_A2_c_110_n N_Y_c_391_n 0.00890453f $X=1.045 $Y=1.675 $X2=0 $Y2=0
cc_128 N_A2_M1003_g N_Y_c_392_n 0.0053571f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_129 N_A2_c_110_n N_Y_c_392_n 0.0058338f $X=1.045 $Y=1.675 $X2=0 $Y2=0
cc_130 N_A2_M1003_g N_Y_c_393_n 0.00104762f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A2_M1003_g N_VGND_c_481_n 0.00269023f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A2_M1003_g N_VGND_c_484_n 0.0044714f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_133 N_A2_M1003_g N_VGND_c_487_n 0.00570261f $X=0.895 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A3_M1002_g N_B1_c_200_n 0.0190653f $X=1.285 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A3_c_157_n N_B1_c_202_n 0.00612653f $X=1.585 $Y=1.27 $X2=0 $Y2=0
cc_136 A3 N_B1_c_202_n 3.60584e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_137 N_A3_c_161_n N_B1_c_209_n 0.0117887f $X=1.585 $Y=1.84 $X2=0 $Y2=0
cc_138 N_A3_M1000_g N_B1_M1008_g 0.0174701f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_139 N_A3_M1002_g N_B1_c_204_n 0.00437327f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A3_c_157_n N_B1_c_204_n 0.00308701f $X=1.585 $Y=1.27 $X2=0 $Y2=0
cc_141 N_A3_c_159_n N_B1_c_205_n 0.0117887f $X=1.585 $Y=1.335 $X2=0 $Y2=0
cc_142 N_A3_c_157_n B1 7.8095e-19 $X=1.585 $Y=1.27 $X2=0 $Y2=0
cc_143 A3 B1 0.04827f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A3_c_157_n N_B1_c_208_n 0.0117887f $X=1.585 $Y=1.27 $X2=0 $Y2=0
cc_145 A3 N_B1_c_208_n 0.00411717f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A3_M1000_g N_VPWR_c_322_n 0.0147848f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_147 N_A3_M1000_g N_VPWR_c_323_n 0.00840515f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_148 N_A3_M1000_g N_VPWR_c_318_n 0.0146909f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_149 N_A3_M1000_g N_A_134_409#_c_355_n 8.82255e-19 $X=1.625 $Y=2.545 $X2=0
+ $Y2=0
cc_150 N_A3_M1000_g N_A_134_409#_c_356_n 0.019556f $X=1.625 $Y=2.545 $X2=0 $Y2=0
cc_151 N_A3_c_161_n N_A_134_409#_c_356_n 5.42828e-19 $X=1.585 $Y=1.84 $X2=0
+ $Y2=0
cc_152 A3 N_A_134_409#_c_356_n 0.0283233f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_153 N_A3_M1000_g N_A_134_409#_c_358_n 0.0162817f $X=1.625 $Y=2.545 $X2=0
+ $Y2=0
cc_154 N_A3_M1002_g N_Y_c_401_n 5.51478e-19 $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_155 N_A3_M1002_g N_Y_c_390_n 0.00110316f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_156 N_A3_M1002_g N_Y_c_391_n 0.0162338f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A3_c_157_n N_Y_c_391_n 0.00903104f $X=1.585 $Y=1.27 $X2=0 $Y2=0
cc_158 A3 N_Y_c_391_n 0.0287058f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A3_M1002_g N_VGND_c_481_n 0.0120617f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A3_M1002_g N_VGND_c_484_n 0.00486043f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A3_M1002_g N_VGND_c_487_n 0.00449619f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_162 N_B1_c_203_n N_C1_c_265_n 0.0104623f $X=2.075 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_163 N_B1_c_206_n N_C1_c_267_n 0.0104623f $X=2.075 $Y=0.805 $X2=0 $Y2=0
cc_164 N_B1_c_209_n N_C1_c_272_n 0.0120211f $X=2.155 $Y=1.84 $X2=0 $Y2=0
cc_165 N_B1_M1008_g N_C1_c_272_n 0.0630873f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_166 B1 N_C1_c_272_n 3.88778e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_167 N_B1_c_205_n N_C1_c_268_n 0.0120211f $X=2.155 $Y=1.675 $X2=0 $Y2=0
cc_168 B1 N_C1_c_268_n 5.20067e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_169 N_B1_c_205_n N_C1_c_269_n 0.0026715f $X=2.155 $Y=1.675 $X2=0 $Y2=0
cc_170 B1 N_C1_c_269_n 0.0301371f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_171 N_B1_c_204_n N_C1_c_270_n 0.00804482f $X=2.155 $Y=1.17 $X2=0 $Y2=0
cc_172 B1 N_C1_c_270_n 0.00112745f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_B1_c_208_n N_C1_c_270_n 0.0120211f $X=2.155 $Y=1.335 $X2=0 $Y2=0
cc_174 N_B1_M1008_g N_VPWR_c_322_n 8.33168e-19 $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_175 N_B1_M1008_g N_VPWR_c_323_n 0.0086001f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_176 N_B1_M1008_g N_VPWR_c_318_n 0.0157977f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_177 N_B1_c_209_n N_A_134_409#_c_356_n 3.02892e-19 $X=2.155 $Y=1.84 $X2=0
+ $Y2=0
cc_178 N_B1_M1008_g N_A_134_409#_c_356_n 0.00438558f $X=2.155 $Y=2.545 $X2=0
+ $Y2=0
cc_179 B1 N_A_134_409#_c_356_n 0.00534367f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_180 N_B1_M1008_g N_A_134_409#_c_358_n 0.0181312f $X=2.155 $Y=2.545 $X2=0
+ $Y2=0
cc_181 N_B1_c_201_n N_Y_c_391_n 0.00924795f $X=2 $Y=0.805 $X2=0 $Y2=0
cc_182 N_B1_c_202_n N_Y_c_391_n 0.0061019f $X=1.79 $Y=0.805 $X2=0 $Y2=0
cc_183 N_B1_c_204_n N_Y_c_391_n 0.00515277f $X=2.155 $Y=1.17 $X2=0 $Y2=0
cc_184 N_B1_c_206_n N_Y_c_391_n 0.0036223f $X=2.075 $Y=0.805 $X2=0 $Y2=0
cc_185 B1 N_Y_c_391_n 0.0097368f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_186 N_B1_c_200_n N_Y_c_428_n 0.00146708f $X=1.715 $Y=0.73 $X2=0 $Y2=0
cc_187 N_B1_c_203_n N_Y_c_428_n 0.00870123f $X=2.075 $Y=0.73 $X2=0 $Y2=0
cc_188 N_B1_c_206_n N_Y_c_428_n 0.00525299f $X=2.075 $Y=0.805 $X2=0 $Y2=0
cc_189 N_B1_c_204_n N_Y_c_394_n 0.00213381f $X=2.155 $Y=1.17 $X2=0 $Y2=0
cc_190 N_B1_c_206_n N_Y_c_394_n 8.54856e-19 $X=2.075 $Y=0.805 $X2=0 $Y2=0
cc_191 B1 N_Y_c_394_n 0.016429f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_192 N_B1_c_208_n N_Y_c_394_n 0.00131253f $X=2.155 $Y=1.335 $X2=0 $Y2=0
cc_193 N_B1_M1008_g N_Y_c_399_n 0.00445114f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_194 N_B1_c_200_n N_VGND_c_481_n 0.0118476f $X=1.715 $Y=0.73 $X2=0 $Y2=0
cc_195 N_B1_c_203_n N_VGND_c_481_n 0.00230268f $X=2.075 $Y=0.73 $X2=0 $Y2=0
cc_196 N_B1_c_200_n N_VGND_c_486_n 0.00486043f $X=1.715 $Y=0.73 $X2=0 $Y2=0
cc_197 N_B1_c_201_n N_VGND_c_486_n 4.87571e-19 $X=2 $Y=0.805 $X2=0 $Y2=0
cc_198 N_B1_c_203_n N_VGND_c_486_n 0.00549284f $X=2.075 $Y=0.73 $X2=0 $Y2=0
cc_199 N_B1_c_200_n N_VGND_c_487_n 0.00436662f $X=1.715 $Y=0.73 $X2=0 $Y2=0
cc_200 N_B1_c_201_n N_VGND_c_487_n 6.51792e-19 $X=2 $Y=0.805 $X2=0 $Y2=0
cc_201 N_B1_c_203_n N_VGND_c_487_n 0.00611432f $X=2.075 $Y=0.73 $X2=0 $Y2=0
cc_202 N_C1_c_271_n N_VPWR_c_323_n 0.0086001f $X=2.685 $Y=2.04 $X2=0 $Y2=0
cc_203 N_C1_c_271_n N_VPWR_c_318_n 0.0165018f $X=2.685 $Y=2.04 $X2=0 $Y2=0
cc_204 N_C1_c_271_n N_A_134_409#_c_356_n 7.23126e-19 $X=2.685 $Y=2.04 $X2=0
+ $Y2=0
cc_205 N_C1_c_271_n N_A_134_409#_c_358_n 0.00376238f $X=2.685 $Y=2.04 $X2=0
+ $Y2=0
cc_206 N_C1_c_265_n N_Y_c_428_n 0.0101675f $X=2.505 $Y=0.78 $X2=0 $Y2=0
cc_207 N_C1_c_266_n N_Y_c_428_n 0.0017408f $X=2.865 $Y=0.78 $X2=0 $Y2=0
cc_208 N_C1_c_267_n N_Y_c_428_n 0.00213085f $X=2.865 $Y=0.855 $X2=0 $Y2=0
cc_209 N_C1_c_271_n N_Y_c_398_n 0.0176224f $X=2.685 $Y=2.04 $X2=0 $Y2=0
cc_210 N_C1_c_267_n N_Y_c_394_n 0.00194918f $X=2.865 $Y=0.855 $X2=0 $Y2=0
cc_211 N_C1_c_271_n N_Y_c_399_n 0.00528392f $X=2.685 $Y=2.04 $X2=0 $Y2=0
cc_212 N_C1_c_268_n N_Y_c_399_n 5.00779e-19 $X=2.725 $Y=1.51 $X2=0 $Y2=0
cc_213 N_C1_c_269_n N_Y_c_399_n 0.00710328f $X=2.725 $Y=1.51 $X2=0 $Y2=0
cc_214 N_C1_c_271_n N_Y_c_395_n 0.00361244f $X=2.685 $Y=2.04 $X2=0 $Y2=0
cc_215 N_C1_c_272_n N_Y_c_395_n 0.00424773f $X=2.685 $Y=1.915 $X2=0 $Y2=0
cc_216 N_C1_c_268_n N_Y_c_395_n 0.00735127f $X=2.725 $Y=1.51 $X2=0 $Y2=0
cc_217 N_C1_c_269_n N_Y_c_395_n 0.0320005f $X=2.725 $Y=1.51 $X2=0 $Y2=0
cc_218 N_C1_c_270_n N_Y_c_395_n 0.00851932f $X=2.725 $Y=1.345 $X2=0 $Y2=0
cc_219 N_C1_c_267_n N_Y_c_396_n 0.0219871f $X=2.865 $Y=0.855 $X2=0 $Y2=0
cc_220 N_C1_c_268_n N_Y_c_396_n 6.68119e-19 $X=2.725 $Y=1.51 $X2=0 $Y2=0
cc_221 N_C1_c_269_n N_Y_c_396_n 0.0156911f $X=2.725 $Y=1.51 $X2=0 $Y2=0
cc_222 N_C1_c_270_n N_Y_c_396_n 0.00610749f $X=2.725 $Y=1.345 $X2=0 $Y2=0
cc_223 N_C1_c_267_n N_Y_c_397_n 2.98157e-19 $X=2.865 $Y=0.855 $X2=0 $Y2=0
cc_224 N_C1_c_270_n N_Y_c_397_n 0.00152854f $X=2.725 $Y=1.345 $X2=0 $Y2=0
cc_225 N_C1_c_265_n N_VGND_c_483_n 0.00227546f $X=2.505 $Y=0.78 $X2=0 $Y2=0
cc_226 N_C1_c_266_n N_VGND_c_483_n 0.0128863f $X=2.865 $Y=0.78 $X2=0 $Y2=0
cc_227 N_C1_c_265_n N_VGND_c_486_n 0.00549284f $X=2.505 $Y=0.78 $X2=0 $Y2=0
cc_228 N_C1_c_266_n N_VGND_c_486_n 0.00486043f $X=2.865 $Y=0.78 $X2=0 $Y2=0
cc_229 N_C1_c_267_n N_VGND_c_486_n 5.84996e-19 $X=2.865 $Y=0.855 $X2=0 $Y2=0
cc_230 N_C1_c_265_n N_VGND_c_487_n 0.00611432f $X=2.505 $Y=0.78 $X2=0 $Y2=0
cc_231 N_C1_c_266_n N_VGND_c_487_n 0.00436662f $X=2.865 $Y=0.78 $X2=0 $Y2=0
cc_232 N_C1_c_267_n N_VGND_c_487_n 7.94744e-19 $X=2.865 $Y=0.855 $X2=0 $Y2=0
cc_233 N_VPWR_c_320_n N_A_134_409#_c_355_n 0.0576214f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_321_n N_A_134_409#_c_355_n 0.021949f $X=1.175 $Y=3.33 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_322_n N_A_134_409#_c_355_n 0.045794f $X=1.34 $Y=2.535 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_318_n N_A_134_409#_c_355_n 0.0124703f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_237 N_VPWR_M1005_d N_A_134_409#_c_356_n 0.00202522f $X=1.2 $Y=2.045 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_322_n N_A_134_409#_c_356_n 0.0164557f $X=1.34 $Y=2.535 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_320_n N_A_134_409#_c_357_n 0.0114859f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_322_n N_A_134_409#_c_358_n 0.0424406f $X=1.34 $Y=2.535 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_323_n N_A_134_409#_c_358_n 0.021949f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_242 N_VPWR_c_318_n N_A_134_409#_c_358_n 0.0124703f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_323_n N_Y_c_398_n 0.0304602f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_318_n N_Y_c_398_n 0.0174175f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_245 N_Y_c_401_n A_116_47# 0.00632947f $X=0.76 $Y=0.545 $X2=-0.19 $Y2=-0.245
cc_246 N_Y_c_390_n A_116_47# 2.80249e-19 $X=0.845 $Y=0.82 $X2=-0.19 $Y2=-0.245
cc_247 N_Y_c_401_n N_VGND_c_481_n 0.00653474f $X=0.76 $Y=0.545 $X2=0 $Y2=0
cc_248 N_Y_c_390_n N_VGND_c_481_n 3.37807e-19 $X=0.845 $Y=0.82 $X2=0 $Y2=0
cc_249 N_Y_c_391_n N_VGND_c_481_n 0.0200683f $X=2.125 $Y=0.905 $X2=0 $Y2=0
cc_250 N_Y_c_428_n N_VGND_c_481_n 0.0125465f $X=2.29 $Y=0.47 $X2=0 $Y2=0
cc_251 N_Y_c_428_n N_VGND_c_483_n 0.0122119f $X=2.29 $Y=0.47 $X2=0 $Y2=0
cc_252 N_Y_c_396_n N_VGND_c_483_n 0.00403394f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_253 N_Y_c_397_n N_VGND_c_483_n 0.0185669f $X=3.155 $Y=0.925 $X2=0 $Y2=0
cc_254 N_Y_c_401_n N_VGND_c_484_n 0.0115084f $X=0.76 $Y=0.545 $X2=0 $Y2=0
cc_255 N_Y_c_393_n N_VGND_c_484_n 0.0189827f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_256 N_Y_c_428_n N_VGND_c_486_n 0.0178561f $X=2.29 $Y=0.47 $X2=0 $Y2=0
cc_257 N_Y_M1006_s N_VGND_c_487_n 0.00232985f $X=0.145 $Y=0.235 $X2=0 $Y2=0
cc_258 N_Y_M1007_d N_VGND_c_487_n 0.0022543f $X=2.15 $Y=0.235 $X2=0 $Y2=0
cc_259 N_Y_c_401_n N_VGND_c_487_n 0.0145831f $X=0.76 $Y=0.545 $X2=0 $Y2=0
cc_260 N_Y_c_391_n N_VGND_c_487_n 0.0278189f $X=2.125 $Y=0.905 $X2=0 $Y2=0
cc_261 N_Y_c_428_n N_VGND_c_487_n 0.0124703f $X=2.29 $Y=0.47 $X2=0 $Y2=0
cc_262 N_Y_c_393_n N_VGND_c_487_n 0.0123683f $X=0.29 $Y=0.445 $X2=0 $Y2=0
cc_263 N_Y_c_396_n N_VGND_c_487_n 0.0139776f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_264 N_Y_c_397_n N_VGND_c_487_n 8.29304e-19 $X=3.155 $Y=0.925 $X2=0 $Y2=0
cc_265 A_116_47# N_VGND_c_487_n 0.00224316f $X=0.58 $Y=0.235 $X2=3.012 $Y2=2.025
cc_266 A_194_47# N_VGND_c_487_n 0.00345006f $X=0.97 $Y=0.235 $X2=3.12 $Y2=0
cc_267 N_VGND_c_487_n A_358_47# 0.00301881f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_268 N_VGND_c_487_n A_516_47# 0.00301881f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
