# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__sdfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__sdfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.510000 0.470000 1.775000 2.130000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.305000 0.255000 10.535000 0.945000 ;
        RECT 10.305000 0.945000 11.910000 1.115000 ;
        RECT 10.310000 1.655000 11.910000 1.825000 ;
        RECT 10.310000 1.825000 10.535000 3.075000 ;
        RECT 11.195000 1.115000 11.910000 1.655000 ;
        RECT 11.205000 0.255000 11.395000 0.945000 ;
        RECT 11.205000 1.825000 11.910000 1.925000 ;
        RECT 11.205000 1.925000 11.395000 3.075000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.395000 2.725000 1.795000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.480000 1.145000 1.340000 1.475000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.255000 1.190000 3.695000 2.120000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 12.000000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 12.190000 3.520000 ;
        RECT  8.735000 1.515000  9.795000 1.655000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.130000  0.635000  0.675000 0.965000 ;
      RECT  0.130000  0.965000  0.310000 1.655000 ;
      RECT  0.130000  1.655000  1.270000 2.300000 ;
      RECT  0.130000  2.300000  2.310000 2.470000 ;
      RECT  0.130000  2.470000  0.855000 2.945000 ;
      RECT  0.845000  0.085000  1.175000 0.975000 ;
      RECT  1.025000  2.640000  1.355000 3.245000 ;
      RECT  1.815000  2.640000  2.650000 2.970000 ;
      RECT  1.945000  0.725000  2.135000 1.045000 ;
      RECT  1.945000  1.045000  3.075000 1.215000 ;
      RECT  2.050000  1.965000  2.310000 2.300000 ;
      RECT  2.480000  2.155000  3.075000 2.335000 ;
      RECT  2.480000  2.335000  3.010000 2.490000 ;
      RECT  2.480000  2.490000  2.650000 2.640000 ;
      RECT  2.750000  0.085000  3.080000 0.875000 ;
      RECT  2.820000  2.660000  3.010000 3.245000 ;
      RECT  2.905000  1.215000  3.075000 2.155000 ;
      RECT  3.180000  2.505000  3.510000 3.075000 ;
      RECT  3.275000  0.785000  4.300000 1.020000 ;
      RECT  3.340000  2.300000  4.300000 2.470000 ;
      RECT  3.340000  2.470000  3.510000 2.505000 ;
      RECT  3.700000  2.640000  3.960000 3.245000 ;
      RECT  3.795000  0.085000  4.125000 0.615000 ;
      RECT  3.865000  1.020000  4.300000 2.300000 ;
      RECT  4.130000  2.470000  4.300000 2.895000 ;
      RECT  4.130000  2.895000  6.045000 3.065000 ;
      RECT  4.295000  0.255000  5.890000 0.495000 ;
      RECT  4.295000  0.495000  4.665000 0.595000 ;
      RECT  4.470000  0.595000  4.665000 1.235000 ;
      RECT  4.470000  1.235000  4.750000 2.725000 ;
      RECT  4.835000  0.665000  5.150000 0.995000 ;
      RECT  4.920000  0.995000  5.150000 2.295000 ;
      RECT  4.920000  2.295000  5.190000 2.625000 ;
      RECT  5.320000  0.665000  5.550000 1.055000 ;
      RECT  5.320000  1.055000  7.095000 1.120000 ;
      RECT  5.360000  1.120000  7.095000 1.305000 ;
      RECT  5.360000  1.305000  5.540000 2.225000 ;
      RECT  5.360000  2.225000  5.705000 2.725000 ;
      RECT  5.710000  1.515000  6.045000 1.845000 ;
      RECT  5.720000  0.495000  5.890000 0.555000 ;
      RECT  5.720000  0.555000  6.935000 0.725000 ;
      RECT  5.875000  1.845000  6.045000 2.635000 ;
      RECT  5.875000  2.635000  7.600000 2.805000 ;
      RECT  5.875000  2.805000  6.045000 2.895000 ;
      RECT  6.225000  1.475000  7.445000 1.655000 ;
      RECT  6.225000  1.655000  7.090000 2.075000 ;
      RECT  6.255000  0.085000  6.585000 0.385000 ;
      RECT  6.410000  2.975000  6.740000 3.245000 ;
      RECT  6.765000  0.255000  7.795000 0.425000 ;
      RECT  6.765000  0.425000  6.935000 0.555000 ;
      RECT  6.920000  2.075000  7.090000 2.205000 ;
      RECT  6.920000  2.205000  7.250000 2.465000 ;
      RECT  7.115000  0.595000  7.445000 0.885000 ;
      RECT  7.270000  1.825000  7.975000 2.005000 ;
      RECT  7.270000  2.005000  7.600000 2.035000 ;
      RECT  7.275000  0.885000  7.445000 1.475000 ;
      RECT  7.430000  2.035000  7.600000 2.635000 ;
      RECT  7.615000  0.425000  7.795000 1.165000 ;
      RECT  7.770000  2.580000  8.325000 2.910000 ;
      RECT  7.805000  1.345000  8.335000 1.515000 ;
      RECT  7.805000  1.515000  7.975000 1.825000 ;
      RECT  7.965000  0.345000  8.685000 0.675000 ;
      RECT  7.975000  0.855000  8.335000 1.345000 ;
      RECT  8.155000  1.695000  8.685000 1.865000 ;
      RECT  8.155000  1.865000  8.325000 2.580000 ;
      RECT  8.495000  2.045000  9.595000 2.215000 ;
      RECT  8.495000  2.215000  8.725000 2.375000 ;
      RECT  8.495000  2.580000  9.225000 3.245000 ;
      RECT  8.515000  0.675000  8.685000 1.185000 ;
      RECT  8.515000  1.185000  9.235000 1.515000 ;
      RECT  8.515000  1.515000  8.685000 1.695000 ;
      RECT  8.855000  0.085000  9.175000 1.015000 ;
      RECT  8.895000  2.405000  9.225000 2.580000 ;
      RECT  9.345000  0.255000  9.605000 1.005000 ;
      RECT  9.395000  2.215000  9.595000 2.975000 ;
      RECT  9.405000  1.005000  9.605000 1.285000 ;
      RECT  9.405000  1.285000 11.015000 1.485000 ;
      RECT  9.405000  1.485000  9.595000 2.045000 ;
      RECT  9.845000  0.085000 10.135000 1.115000 ;
      RECT  9.845000  1.815000 10.140000 3.245000 ;
      RECT 10.705000  0.085000 11.035000 0.775000 ;
      RECT 10.705000  1.995000 11.035000 3.245000 ;
      RECT 11.565000  0.085000 11.895000 0.775000 ;
      RECT 11.565000  2.095000 11.895000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  2.320000  2.725000 2.490000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  2.320000  5.125000 2.490000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
    LAYER met1 ;
      RECT 2.495000 2.290000 2.785000 2.335000 ;
      RECT 2.495000 2.335000 5.185000 2.475000 ;
      RECT 2.495000 2.475000 2.785000 2.520000 ;
      RECT 4.895000 2.290000 5.185000 2.335000 ;
      RECT 4.895000 2.475000 5.185000 2.520000 ;
  END
END sky130_fd_sc_lp__sdfxtp_4
END LIBRARY
