* File: sky130_fd_sc_lp__inputiso0p_lp.pxi.spice
* Created: Fri Aug 28 10:37:09 2020
* 
x_PM_SKY130_FD_SC_LP__INPUTISO0P_LP%SLEEP N_SLEEP_M1012_g N_SLEEP_M1005_g
+ N_SLEEP_M1006_g N_SLEEP_M1002_g SLEEP SLEEP N_SLEEP_c_65_n
+ PM_SKY130_FD_SC_LP__INPUTISO0P_LP%SLEEP
x_PM_SKY130_FD_SC_LP__INPUTISO0P_LP%A_27_93# N_A_27_93#_M1012_s
+ N_A_27_93#_M1005_s N_A_27_93#_M1011_g N_A_27_93#_M1007_g N_A_27_93#_M1013_g
+ N_A_27_93#_c_97_n N_A_27_93#_c_102_n N_A_27_93#_c_103_n N_A_27_93#_c_116_n
+ N_A_27_93#_c_98_n N_A_27_93#_c_105_n
+ PM_SKY130_FD_SC_LP__INPUTISO0P_LP%A_27_93#
x_PM_SKY130_FD_SC_LP__INPUTISO0P_LP%A N_A_M1001_g N_A_c_151_n N_A_M1000_g
+ N_A_M1010_g N_A_c_154_n N_A_c_155_n A N_A_c_156_n N_A_c_159_n
+ PM_SKY130_FD_SC_LP__INPUTISO0P_LP%A
x_PM_SKY130_FD_SC_LP__INPUTISO0P_LP%A_342_489# N_A_342_489#_M1001_d
+ N_A_342_489#_M1013_d N_A_342_489#_c_197_n N_A_342_489#_M1003_g
+ N_A_342_489#_M1008_g N_A_342_489#_c_198_n N_A_342_489#_M1004_g
+ N_A_342_489#_M1009_g N_A_342_489#_c_207_n N_A_342_489#_c_208_n
+ N_A_342_489#_c_209_n N_A_342_489#_c_199_n N_A_342_489#_c_200_n
+ N_A_342_489#_c_201_n N_A_342_489#_c_202_n N_A_342_489#_c_203_n
+ N_A_342_489#_c_204_n PM_SKY130_FD_SC_LP__INPUTISO0P_LP%A_342_489#
x_PM_SKY130_FD_SC_LP__INPUTISO0P_LP%VPWR N_VPWR_M1002_d N_VPWR_M1010_d
+ N_VPWR_c_266_n N_VPWR_c_267_n VPWR N_VPWR_c_268_n N_VPWR_c_269_n
+ N_VPWR_c_270_n N_VPWR_c_265_n N_VPWR_c_272_n N_VPWR_c_273_n
+ PM_SKY130_FD_SC_LP__INPUTISO0P_LP%VPWR
x_PM_SKY130_FD_SC_LP__INPUTISO0P_LP%X N_X_M1004_d N_X_M1009_d X X X X X
+ N_X_c_311_n PM_SKY130_FD_SC_LP__INPUTISO0P_LP%X
x_PM_SKY130_FD_SC_LP__INPUTISO0P_LP%VGND N_VGND_M1006_d N_VGND_M1003_s
+ N_VGND_c_321_n N_VGND_c_322_n VGND N_VGND_c_323_n N_VGND_c_324_n
+ N_VGND_c_325_n N_VGND_c_326_n N_VGND_c_327_n N_VGND_c_328_n
+ PM_SKY130_FD_SC_LP__INPUTISO0P_LP%VGND
cc_1 VNB N_SLEEP_M1012_g 0.0340203f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.675
cc_2 VNB N_SLEEP_M1006_g 0.035339f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=0.675
cc_3 VNB SLEEP 0.00855277f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_SLEEP_c_65_n 0.0357139f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.465
cc_5 VNB N_A_27_93#_M1007_g 0.0380418f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.985
cc_6 VNB N_A_27_93#_c_97_n 0.0426945f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.465
cc_7 VNB N_A_27_93#_c_98_n 0.0440266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_c_151_n 0.0109922f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.985
cc_9 VNB N_A_M1000_g 3.61206e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_M1010_g 3.74535e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_154_n 0.017557f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.655
cc_12 VNB N_A_c_155_n 0.0170764f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.655
cc_13 VNB N_A_c_156_n 0.0536741f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.465
cc_14 VNB N_A_342_489#_c_197_n 0.0188631f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.655
cc_15 VNB N_A_342_489#_c_198_n 0.020326f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.655
cc_16 VNB N_A_342_489#_c_199_n 0.00555058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_342_489#_c_200_n 0.0220155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_342_489#_c_201_n 0.0010417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_342_489#_c_202_n 0.0015967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_342_489#_c_203_n 0.00393769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_342_489#_c_204_n 0.0639765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_265_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_311_n 0.0647669f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_24 VNB N_VGND_c_321_n 0.0162715f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.3
cc_25 VNB N_VGND_c_322_n 0.0186777f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.985
cc_26 VNB N_VGND_c_323_n 0.0291685f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_27 VNB N_VGND_c_324_n 0.0295741f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.465
cc_28 VNB N_VGND_c_325_n 0.0303334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_326_n 0.271448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_327_n 0.0130796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_328_n 0.00644364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_SLEEP_M1005_g 0.038312f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.655
cc_33 VPB N_SLEEP_M1002_g 0.0307205f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.655
cc_34 VPB N_SLEEP_c_65_n 0.0330344f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.465
cc_35 VPB N_A_27_93#_M1011_g 0.0304093f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.3
cc_36 VPB N_A_27_93#_M1013_g 0.0324565f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_37 VPB N_A_27_93#_c_97_n 0.0197538f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.465
cc_38 VPB N_A_27_93#_c_102_n 0.0100893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_93#_c_103_n 0.0322681f $X=-0.19 $Y=1.655 $X2=0.732 $Y2=1.465
cc_40 VPB N_A_27_93#_c_98_n 0.0320078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_27_93#_c_105_n 0.00739525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_M1000_g 0.0475243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_M1010_g 0.0488228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_c_159_n 0.00506862f $X=-0.19 $Y=1.655 $X2=0.732 $Y2=1.295
cc_45 VPB N_A_342_489#_M1008_g 0.0180556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_342_489#_M1009_g 0.0199177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_342_489#_c_207_n 0.00687382f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.465
cc_48 VPB N_A_342_489#_c_208_n 0.0120722f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_342_489#_c_209_n 0.00990386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_342_489#_c_203_n 0.00161812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_342_489#_c_204_n 0.00366798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_266_n 0.0133194f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.3
cc_53 VPB N_VPWR_c_267_n 0.0106604f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.985
cc_54 VPB N_VPWR_c_268_n 0.0292919f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_55 VPB N_VPWR_c_269_n 0.0399828f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.465
cc_56 VPB N_VPWR_c_270_n 0.02737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_265_n 0.0972216f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_272_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_273_n 0.00601838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_X_c_311_n 0.0630605f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_61 N_SLEEP_M1002_g N_A_27_93#_M1011_g 0.0312625f $X=0.845 $Y=2.655 $X2=0
+ $Y2=0
cc_62 N_SLEEP_M1006_g N_A_27_93#_M1007_g 0.0116365f $X=0.845 $Y=0.675 $X2=0
+ $Y2=0
cc_63 SLEEP N_A_27_93#_M1007_g 7.25913e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_64 N_SLEEP_M1012_g N_A_27_93#_c_97_n 0.0412295f $X=0.485 $Y=0.675 $X2=0 $Y2=0
cc_65 SLEEP N_A_27_93#_c_97_n 0.0568433f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_66 N_SLEEP_M1005_g N_A_27_93#_c_102_n 0.00952698f $X=0.485 $Y=2.655 $X2=0
+ $Y2=0
cc_67 N_SLEEP_M1005_g N_A_27_93#_c_103_n 0.0200033f $X=0.485 $Y=2.655 $X2=0
+ $Y2=0
cc_68 N_SLEEP_M1002_g N_A_27_93#_c_103_n 0.0138102f $X=0.845 $Y=2.655 $X2=0
+ $Y2=0
cc_69 SLEEP N_A_27_93#_c_103_n 0.0292015f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_SLEEP_c_65_n N_A_27_93#_c_103_n 8.69237e-19 $X=0.71 $Y=1.465 $X2=0 $Y2=0
cc_71 SLEEP N_A_27_93#_c_116_n 0.0260401f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_SLEEP_c_65_n N_A_27_93#_c_116_n 0.0032643f $X=0.71 $Y=1.465 $X2=0 $Y2=0
cc_73 SLEEP N_A_27_93#_c_98_n 0.00270332f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_SLEEP_c_65_n N_A_27_93#_c_98_n 0.0312625f $X=0.71 $Y=1.465 $X2=0 $Y2=0
cc_75 N_SLEEP_M1005_g N_VPWR_c_266_n 0.00185559f $X=0.485 $Y=2.655 $X2=0 $Y2=0
cc_76 N_SLEEP_M1002_g N_VPWR_c_266_n 0.0124876f $X=0.845 $Y=2.655 $X2=0 $Y2=0
cc_77 N_SLEEP_M1005_g N_VPWR_c_268_n 0.00510437f $X=0.485 $Y=2.655 $X2=0 $Y2=0
cc_78 N_SLEEP_M1002_g N_VPWR_c_268_n 0.00424179f $X=0.845 $Y=2.655 $X2=0 $Y2=0
cc_79 N_SLEEP_M1005_g N_VPWR_c_265_n 0.00515964f $X=0.485 $Y=2.655 $X2=0 $Y2=0
cc_80 N_SLEEP_M1002_g N_VPWR_c_265_n 0.0043341f $X=0.845 $Y=2.655 $X2=0 $Y2=0
cc_81 N_SLEEP_M1012_g N_VGND_c_321_n 0.00161762f $X=0.485 $Y=0.675 $X2=0 $Y2=0
cc_82 N_SLEEP_M1006_g N_VGND_c_321_n 0.0125781f $X=0.845 $Y=0.675 $X2=0 $Y2=0
cc_83 SLEEP N_VGND_c_321_n 0.00116827f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_84 N_SLEEP_M1012_g N_VGND_c_323_n 0.00510437f $X=0.485 $Y=0.675 $X2=0 $Y2=0
cc_85 N_SLEEP_M1006_g N_VGND_c_323_n 0.00424179f $X=0.845 $Y=0.675 $X2=0 $Y2=0
cc_86 N_SLEEP_M1012_g N_VGND_c_326_n 0.00515964f $X=0.485 $Y=0.675 $X2=0 $Y2=0
cc_87 N_SLEEP_M1006_g N_VGND_c_326_n 0.0043341f $X=0.845 $Y=0.675 $X2=0 $Y2=0
cc_88 N_A_27_93#_M1007_g N_A_c_151_n 0.00439272f $X=1.625 $Y=0.675 $X2=0 $Y2=0
cc_89 N_A_27_93#_c_116_n N_A_M1000_g 0.0011996f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_90 N_A_27_93#_c_98_n N_A_M1000_g 0.0386444f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_91 N_A_27_93#_M1007_g N_A_c_154_n 0.0484202f $X=1.625 $Y=0.675 $X2=0 $Y2=0
cc_92 N_A_27_93#_c_116_n N_A_c_156_n 9.47243e-19 $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_93 N_A_27_93#_c_98_n N_A_c_156_n 0.021439f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_94 N_A_27_93#_c_116_n N_A_c_159_n 0.0152671f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_95 N_A_27_93#_c_98_n N_A_c_159_n 0.0020496f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_96 N_A_27_93#_M1013_g N_A_342_489#_c_207_n 0.00628397f $X=1.635 $Y=2.655
+ $X2=0 $Y2=0
cc_97 N_A_27_93#_c_103_n N_A_342_489#_c_207_n 0.00888624f $X=1.2 $Y=2.15 $X2=0
+ $Y2=0
cc_98 N_A_27_93#_c_103_n N_A_342_489#_c_209_n 0.00534853f $X=1.2 $Y=2.15 $X2=0
+ $Y2=0
cc_99 N_A_27_93#_c_116_n N_A_342_489#_c_209_n 0.00931347f $X=1.43 $Y=1.475 $X2=0
+ $Y2=0
cc_100 N_A_27_93#_c_98_n N_A_342_489#_c_209_n 0.0014554f $X=1.43 $Y=1.475 $X2=0
+ $Y2=0
cc_101 N_A_27_93#_M1007_g N_A_342_489#_c_201_n 0.00100859f $X=1.625 $Y=0.675
+ $X2=0 $Y2=0
cc_102 N_A_27_93#_M1011_g N_VPWR_c_266_n 0.0126163f $X=1.275 $Y=2.655 $X2=0
+ $Y2=0
cc_103 N_A_27_93#_M1013_g N_VPWR_c_266_n 0.00186774f $X=1.635 $Y=2.655 $X2=0
+ $Y2=0
cc_104 N_A_27_93#_c_103_n N_VPWR_c_266_n 0.0186033f $X=1.2 $Y=2.15 $X2=0 $Y2=0
cc_105 N_A_27_93#_c_102_n N_VPWR_c_268_n 0.00593896f $X=0.27 $Y=2.61 $X2=0 $Y2=0
cc_106 N_A_27_93#_M1011_g N_VPWR_c_269_n 0.00424179f $X=1.275 $Y=2.655 $X2=0
+ $Y2=0
cc_107 N_A_27_93#_M1013_g N_VPWR_c_269_n 0.00510437f $X=1.635 $Y=2.655 $X2=0
+ $Y2=0
cc_108 N_A_27_93#_M1011_g N_VPWR_c_265_n 0.0043341f $X=1.275 $Y=2.655 $X2=0
+ $Y2=0
cc_109 N_A_27_93#_M1013_g N_VPWR_c_265_n 0.00515964f $X=1.635 $Y=2.655 $X2=0
+ $Y2=0
cc_110 N_A_27_93#_c_102_n N_VPWR_c_265_n 0.00742155f $X=0.27 $Y=2.61 $X2=0 $Y2=0
cc_111 N_A_27_93#_M1007_g N_VGND_c_321_n 0.0127454f $X=1.625 $Y=0.675 $X2=0
+ $Y2=0
cc_112 N_A_27_93#_c_97_n N_VGND_c_321_n 0.00748999f $X=0.27 $Y=0.72 $X2=0 $Y2=0
cc_113 N_A_27_93#_c_116_n N_VGND_c_321_n 0.0118129f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_114 N_A_27_93#_c_98_n N_VGND_c_321_n 0.00765182f $X=1.43 $Y=1.475 $X2=0 $Y2=0
cc_115 N_A_27_93#_c_97_n N_VGND_c_323_n 0.00734893f $X=0.27 $Y=0.72 $X2=0 $Y2=0
cc_116 N_A_27_93#_M1007_g N_VGND_c_324_n 0.00424179f $X=1.625 $Y=0.675 $X2=0
+ $Y2=0
cc_117 N_A_27_93#_M1007_g N_VGND_c_326_n 0.0043341f $X=1.625 $Y=0.675 $X2=0
+ $Y2=0
cc_118 N_A_27_93#_c_97_n N_VGND_c_326_n 0.00765198f $X=0.27 $Y=0.72 $X2=0 $Y2=0
cc_119 N_A_M1000_g N_A_342_489#_c_207_n 0.00652706f $X=2.085 $Y=2.655 $X2=0
+ $Y2=0
cc_120 N_A_M1000_g N_A_342_489#_c_208_n 0.0144643f $X=2.085 $Y=2.655 $X2=0 $Y2=0
cc_121 N_A_M1010_g N_A_342_489#_c_208_n 0.01506f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_122 N_A_c_156_n N_A_342_489#_c_208_n 9.9437e-19 $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_123 N_A_c_159_n N_A_342_489#_c_208_n 0.0443923f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_124 N_A_c_154_n N_A_342_489#_c_199_n 0.00656473f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_155_n N_A_342_489#_c_199_n 0.00111161f $X=2.02 $Y=1.145 $X2=0 $Y2=0
cc_126 N_A_c_156_n N_A_342_489#_c_200_n 0.00949144f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_127 N_A_c_159_n N_A_342_489#_c_200_n 0.0266037f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_128 N_A_c_151_n N_A_342_489#_c_201_n 0.00403612f $X=2.055 $Y=1.315 $X2=0
+ $Y2=0
cc_129 N_A_c_155_n N_A_342_489#_c_201_n 0.00634201f $X=2.02 $Y=1.145 $X2=0 $Y2=0
cc_130 N_A_c_156_n N_A_342_489#_c_201_n 0.00511378f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_131 N_A_c_159_n N_A_342_489#_c_201_n 0.0177261f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_132 N_A_c_151_n N_A_342_489#_c_203_n 0.00198796f $X=2.055 $Y=1.315 $X2=0
+ $Y2=0
cc_133 N_A_M1010_g N_A_342_489#_c_203_n 0.00248423f $X=2.445 $Y=2.655 $X2=0
+ $Y2=0
cc_134 N_A_c_156_n N_A_342_489#_c_203_n 0.00356425f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_135 N_A_c_159_n N_A_342_489#_c_203_n 0.0305846f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_136 N_A_M1010_g N_A_342_489#_c_204_n 0.0310943f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_137 N_A_c_156_n N_A_342_489#_c_204_n 0.0217991f $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_138 N_A_c_159_n N_A_342_489#_c_204_n 6.78031e-19 $X=2.485 $Y=1.48 $X2=0 $Y2=0
cc_139 N_A_M1010_g N_VPWR_c_267_n 0.00861135f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_140 N_A_M1000_g N_VPWR_c_269_n 0.00510437f $X=2.085 $Y=2.655 $X2=0 $Y2=0
cc_141 N_A_M1010_g N_VPWR_c_269_n 0.00510437f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_142 N_A_M1000_g N_VPWR_c_265_n 0.00515964f $X=2.085 $Y=2.655 $X2=0 $Y2=0
cc_143 N_A_M1010_g N_VPWR_c_265_n 0.00515964f $X=2.445 $Y=2.655 $X2=0 $Y2=0
cc_144 N_A_c_154_n N_VGND_c_321_n 0.00161762f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_154_n N_VGND_c_322_n 0.00333051f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_154_n N_VGND_c_324_n 0.00510437f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_154_n N_VGND_c_326_n 0.00515964f $X=2.02 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_342_489#_c_208_n N_VPWR_M1010_d 0.00859922f $X=2.82 $Y=2.04 $X2=0
+ $Y2=0
cc_149 N_A_342_489#_M1008_g N_VPWR_c_267_n 0.0241518f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_342_489#_M1009_g N_VPWR_c_267_n 0.00358702f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_342_489#_c_207_n N_VPWR_c_267_n 0.00530717f $X=1.87 $Y=2.61 $X2=0
+ $Y2=0
cc_152 N_A_342_489#_c_208_n N_VPWR_c_267_n 0.0268559f $X=2.82 $Y=2.04 $X2=0
+ $Y2=0
cc_153 N_A_342_489#_c_207_n N_VPWR_c_269_n 0.00564047f $X=1.87 $Y=2.61 $X2=0
+ $Y2=0
cc_154 N_A_342_489#_M1008_g N_VPWR_c_270_n 0.00388479f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_342_489#_M1009_g N_VPWR_c_270_n 0.00585385f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_342_489#_M1008_g N_VPWR_c_265_n 0.006597f $X=2.935 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_342_489#_M1009_g N_VPWR_c_265_n 0.0116546f $X=3.295 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A_342_489#_c_207_n N_VPWR_c_265_n 0.00707389f $X=1.87 $Y=2.61 $X2=0
+ $Y2=0
cc_159 N_A_342_489#_c_208_n A_602_367# 0.00433061f $X=2.82 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_342_489#_c_198_n N_X_c_311_n 0.032245f $X=3.295 $Y=1.005 $X2=0 $Y2=0
cc_161 N_A_342_489#_c_202_n N_X_c_311_n 0.0185607f $X=3.025 $Y=1.225 $X2=0 $Y2=0
cc_162 N_A_342_489#_c_203_n N_X_c_311_n 0.0538185f $X=3.025 $Y=1.955 $X2=0 $Y2=0
cc_163 N_A_342_489#_c_199_n N_VGND_c_321_n 0.00748572f $X=2.2 $Y=0.72 $X2=0
+ $Y2=0
cc_164 N_A_342_489#_c_197_n N_VGND_c_322_n 0.0132046f $X=2.935 $Y=1.17 $X2=0
+ $Y2=0
cc_165 N_A_342_489#_c_198_n N_VGND_c_322_n 0.00168986f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_166 N_A_342_489#_c_199_n N_VGND_c_322_n 0.0247472f $X=2.2 $Y=0.72 $X2=0 $Y2=0
cc_167 N_A_342_489#_c_200_n N_VGND_c_322_n 0.0219254f $X=2.82 $Y=1.115 $X2=0
+ $Y2=0
cc_168 N_A_342_489#_c_202_n N_VGND_c_322_n 0.00386325f $X=3.025 $Y=1.225 $X2=0
+ $Y2=0
cc_169 N_A_342_489#_c_199_n N_VGND_c_324_n 0.00701182f $X=2.2 $Y=0.72 $X2=0
+ $Y2=0
cc_170 N_A_342_489#_c_197_n N_VGND_c_325_n 0.00424179f $X=2.935 $Y=1.17 $X2=0
+ $Y2=0
cc_171 N_A_342_489#_c_198_n N_VGND_c_325_n 0.00510437f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_172 N_A_342_489#_c_197_n N_VGND_c_326_n 0.0043341f $X=2.935 $Y=1.17 $X2=0
+ $Y2=0
cc_173 N_A_342_489#_c_198_n N_VGND_c_326_n 0.00515964f $X=3.295 $Y=1.005 $X2=0
+ $Y2=0
cc_174 N_A_342_489#_c_199_n N_VGND_c_326_n 0.00730097f $X=2.2 $Y=0.72 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_265_n A_602_367# 0.00899413f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_176 N_VPWR_c_265_n N_X_M1009_d 0.00319521f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_177 N_VPWR_c_270_n N_X_c_311_n 0.0240782f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_178 N_VPWR_c_265_n N_X_c_311_n 0.0137238f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_179 N_X_c_311_n N_VGND_c_325_n 0.0101312f $X=3.51 $Y=0.72 $X2=0 $Y2=0
cc_180 N_X_c_311_n N_VGND_c_326_n 0.0121005f $X=3.51 $Y=0.72 $X2=0 $Y2=0
