# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfrtp_ov2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfrtp_ov2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.565000 2.255000 1.805000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.085000 0.255000 13.355000 3.075000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.800000 1.940000 6.130000 2.320000 ;
        RECT 5.800000 2.320000 6.950000 2.490000 ;
        RECT 5.800000 2.490000 6.130000 2.545000 ;
        RECT 6.770000 2.490000 6.950000 2.905000 ;
        RECT 6.770000 2.905000 8.285000 3.075000 ;
        RECT 8.035000 2.475000 9.270000 2.570000 ;
        RECT 8.035000 2.570000 9.215000 2.645000 ;
        RECT 8.035000 2.645000 8.285000 2.905000 ;
        RECT 8.940000 2.255000 9.270000 2.475000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 1.175000 3.310000 2.145000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.285000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.200000 2.795000 1.395000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 11.550000 1.425000 11.880000 2.500000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.440000 0.085000 ;
      RECT  0.000000  3.245000 13.440000 3.415000 ;
      RECT  0.090000  0.415000  0.430000 0.860000 ;
      RECT  0.090000  0.860000  1.510000 1.030000 ;
      RECT  0.090000  1.030000  0.370000 1.975000 ;
      RECT  0.090000  1.975000  2.675000 2.145000 ;
      RECT  0.090000  2.145000  1.140000 2.965000 ;
      RECT  0.600000  0.085000  0.895000 0.690000 ;
      RECT  1.145000  0.265000  3.225000 0.435000 ;
      RECT  1.145000  0.435000  1.355000 0.595000 ;
      RECT  1.320000  2.390000  1.650000 3.245000 ;
      RECT  1.990000  0.615000  2.320000 0.815000 ;
      RECT  1.990000  0.815000  4.215000 0.985000 ;
      RECT  2.110000  2.315000  3.885000 2.485000 ;
      RECT  2.110000  2.485000  2.440000 2.680000 ;
      RECT  2.425000  1.815000  2.675000 1.975000 ;
      RECT  2.895000  0.435000  3.225000 0.635000 ;
      RECT  3.070000  2.655000  3.400000 3.245000 ;
      RECT  3.405000  0.085000  3.735000 0.635000 ;
      RECT  3.480000  0.985000  3.685000 2.295000 ;
      RECT  3.480000  2.295000  3.885000 2.315000 ;
      RECT  3.590000  2.485000  3.885000 2.625000 ;
      RECT  3.855000  1.155000  4.215000 1.915000 ;
      RECT  4.015000  0.655000  4.215000 0.815000 ;
      RECT  4.065000  2.085000  4.555000 2.165000 ;
      RECT  4.065000  2.165000  5.630000 2.335000 ;
      RECT  4.065000  2.335000  4.385000 2.690000 ;
      RECT  4.385000  0.785000  5.670000 0.995000 ;
      RECT  4.385000  0.995000  4.555000 2.085000 ;
      RECT  4.725000  1.600000  6.835000 1.770000 ;
      RECT  4.725000  1.770000  5.015000 1.995000 ;
      RECT  4.735000  1.165000  5.125000 1.430000 ;
      RECT  4.865000  2.505000  5.195000 3.245000 ;
      RECT  5.365000  2.335000  5.630000 2.690000 ;
      RECT  5.465000  0.995000  5.670000 1.170000 ;
      RECT  5.465000  1.170000  6.475000 1.430000 ;
      RECT  6.145000  0.085000  6.475000 0.940000 ;
      RECT  6.270000  2.660000  6.600000 3.245000 ;
      RECT  6.645000  0.630000  6.835000 1.600000 ;
      RECT  6.655000  1.770000  6.835000 1.960000 ;
      RECT  6.655000  1.960000  7.145000 2.150000 ;
      RECT  7.005000  0.745000  8.320000 0.915000 ;
      RECT  7.005000  0.915000  7.175000 1.620000 ;
      RECT  7.005000  1.620000  7.575000 1.790000 ;
      RECT  7.200000  0.625000  7.870000 0.745000 ;
      RECT  7.315000  1.790000  7.575000 2.735000 ;
      RECT  7.345000  1.095000  7.940000 1.425000 ;
      RECT  7.770000  1.425000  7.940000 2.055000 ;
      RECT  7.770000  2.055000  8.120000 2.305000 ;
      RECT  8.110000  0.915000  8.320000 1.135000 ;
      RECT  8.110000  1.135000 10.045000 1.305000 ;
      RECT  8.110000  1.485000  8.370000 1.555000 ;
      RECT  8.110000  1.555000 10.045000 1.725000 ;
      RECT  8.110000  1.725000  8.370000 1.815000 ;
      RECT  8.400000  2.055000  9.620000 2.075000 ;
      RECT  8.400000  2.075000  8.730000 2.305000 ;
      RECT  8.455000  2.855000  9.190000 3.245000 ;
      RECT  8.490000  0.085000  8.820000 0.965000 ;
      RECT  8.560000  1.905000  9.620000 2.055000 ;
      RECT  9.360000  2.745000  9.620000 3.075000 ;
      RECT  9.425000  0.255000 10.155000 0.475000 ;
      RECT  9.425000  0.475000  9.705000 0.965000 ;
      RECT  9.450000  2.075000  9.620000 2.745000 ;
      RECT  9.480000  1.305000 10.045000 1.385000 ;
      RECT  9.790000  2.710000 10.050000 3.245000 ;
      RECT  9.800000  1.725000 10.045000 2.370000 ;
      RECT  9.800000  2.370000 11.380000 2.540000 ;
      RECT  9.875000  0.645000 11.980000 0.815000 ;
      RECT  9.875000  0.815000 10.045000 1.135000 ;
      RECT 10.215000  0.985000 10.575000 1.165000 ;
      RECT 10.215000  1.165000 10.545000 2.200000 ;
      RECT 10.715000  1.345000 11.380000 2.370000 ;
      RECT 10.755000  0.085000 11.085000 0.475000 ;
      RECT 10.755000  2.710000 11.040000 3.245000 ;
      RECT 11.200000  0.985000 11.630000 1.185000 ;
      RECT 11.200000  1.185000 11.380000 1.345000 ;
      RECT 11.210000  2.540000 11.380000 2.715000 ;
      RECT 11.210000  2.715000 11.630000 3.045000 ;
      RECT 11.810000  0.815000 11.980000 0.985000 ;
      RECT 11.810000  0.985000 12.455000 1.165000 ;
      RECT 12.050000  1.675000 12.915000 1.845000 ;
      RECT 12.050000  1.845000 12.260000 2.495000 ;
      RECT 12.125000  1.165000 12.455000 1.505000 ;
      RECT 12.150000  0.275000 12.405000 0.645000 ;
      RECT 12.150000  0.645000 12.915000 0.815000 ;
      RECT 12.430000  2.015000 12.915000 3.245000 ;
      RECT 12.575000  0.085000 12.915000 0.475000 ;
      RECT 12.665000  0.815000 12.915000 1.675000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  1.210000  4.165000 1.380000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.210000  5.125000 1.380000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.210000  7.525000 1.380000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  1.210000 10.405000 1.380000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
    LAYER met1 ;
      RECT  3.935000 1.180000  4.225000 1.225000 ;
      RECT  3.935000 1.225000 10.465000 1.365000 ;
      RECT  3.935000 1.365000  4.225000 1.410000 ;
      RECT  4.895000 1.180000  5.185000 1.225000 ;
      RECT  4.895000 1.365000  5.185000 1.410000 ;
      RECT  7.295000 1.180000  7.585000 1.225000 ;
      RECT  7.295000 1.365000  7.585000 1.410000 ;
      RECT 10.175000 1.180000 10.465000 1.225000 ;
      RECT 10.175000 1.365000 10.465000 1.410000 ;
  END
END sky130_fd_sc_lp__sdfrtp_ov2
