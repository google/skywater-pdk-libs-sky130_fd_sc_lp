* File: sky130_fd_sc_lp__einvn_1.pex.spice
* Created: Wed Sep  2 09:51:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVN_1%A 3 6 8 9 13 15
c29 15 0 1.09601e-19 $X=0.665 $Y=1.315
r30 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.48
+ $X2=0.665 $Y2=1.645
r31 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.48
+ $X2=0.665 $Y2=1.315
r32 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.665
+ $Y=1.48 $X2=0.665 $Y2=1.48
r33 9 14 5.33005 $w=3.98e-07 $l=1.85e-07 $layer=LI1_cond $X=0.7 $Y=1.665 $X2=0.7
+ $Y2=1.48
r34 8 14 5.33005 $w=3.98e-07 $l=1.85e-07 $layer=LI1_cond $X=0.7 $Y=1.295 $X2=0.7
+ $Y2=1.48
r35 6 16 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.755 $Y=2.465
+ $X2=0.755 $Y2=1.645
r36 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.755 $Y=0.785
+ $X2=0.755 $Y2=1.315
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_1%A_214_21# 1 2 7 9 10 11 13 17 22 23 26 28
r46 26 27 8.11215 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=1.105
+ $X2=2.115 $Y2=1.27
r47 23 27 38.9681 $w=1.83e-07 $l=6.5e-07 $layer=LI1_cond $X=2.222 $Y=1.92
+ $X2=2.222 $Y2=1.27
r48 22 23 8.2055 $w=5.13e-07 $l=1.3e-07 $layer=LI1_cond $X=2.057 $Y=2.05
+ $X2=2.057 $Y2=1.92
r49 18 28 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.945 $Y=0.38
+ $X2=1.945 $Y2=0.18
r50 17 20 6.37706 $w=5.33e-07 $l=2.5e-07 $layer=LI1_cond $X=2.047 $Y=0.38
+ $X2=2.047 $Y2=0.63
r51 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.945
+ $Y=0.38 $X2=1.945 $Y2=0.38
r52 13 26 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=2.115 $Y=1.07
+ $X2=2.115 $Y2=1.105
r53 13 20 12.6769 $w=3.98e-07 $l=4.4e-07 $layer=LI1_cond $X=2.115 $Y=1.07
+ $X2=2.115 $Y2=0.63
r54 10 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=0.18
+ $X2=1.945 $Y2=0.18
r55 10 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.78 $Y=0.18
+ $X2=1.22 $Y2=0.18
r56 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.145 $Y=0.255
+ $X2=1.22 $Y2=0.18
r57 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.145 $Y=0.255
+ $X2=1.145 $Y2=0.785
r58 2 22 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=1.905 $X2=1.965 $Y2=2.05
r59 1 26 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.885 $X2=2.045 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_1%TE_B 1 3 4 5 8 12 13 14 18 19 20
c45 5 0 2.61772e-20 $X=1.22 $Y=1.635
r46 21 22 36.5941 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.795 $Y=1.635
+ $X2=1.795 $Y2=1.745
r47 18 21 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.795 $Y=1.58
+ $X2=1.795 $Y2=1.635
r48 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.58
+ $X2=1.795 $Y2=1.415
r49 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.795
+ $Y=1.58 $X2=1.795 $Y2=1.58
r50 14 19 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.622
+ $X2=1.795 $Y2=1.622
r51 13 14 21.693 $w=2.53e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.622 $X2=1.68
+ $Y2=1.622
r52 12 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.83 $Y=1.095
+ $X2=1.83 $Y2=1.415
r53 8 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.75 $Y=2.225
+ $X2=1.75 $Y2=1.745
r54 4 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.635
+ $X2=1.795 $Y2=1.635
r55 4 5 159.371 $w=1.8e-07 $l=4.1e-07 $layer=POLY_cond $X=1.63 $Y=1.635 $X2=1.22
+ $Y2=1.635
r56 1 5 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.145 $Y=1.725
+ $X2=1.22 $Y2=1.635
r57 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.145 $Y=1.725
+ $X2=1.145 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_1%Z 1 2 7 9 16 17 18
r26 18 43 2.56827 $w=8.13e-07 $l=1.75e-07 $layer=LI1_cond $X=0.492 $Y=2.775
+ $X2=0.492 $Y2=2.95
r27 17 18 5.43005 $w=8.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.492 $Y=2.405
+ $X2=0.492 $Y2=2.775
r28 16 17 5.43005 $w=8.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.492 $Y=2.035
+ $X2=0.492 $Y2=2.405
r29 12 16 26.4604 $w=4.13e-07 $l=9.1e-07 $layer=LI1_cond $X=0.207 $Y=1.04
+ $X2=0.207 $Y2=1.95
r30 11 12 2.58917 $w=2.45e-07 $l=1.68e-07 $layer=LI1_cond $X=0.207 $Y=0.872
+ $X2=0.207 $Y2=1.04
r31 7 11 11.4556 $w=3.33e-07 $l=3.33e-07 $layer=LI1_cond $X=0.54 $Y=0.872
+ $X2=0.207 $Y2=0.872
r32 7 9 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.54 $Y=0.705
+ $X2=0.54 $Y2=0.51
r33 2 43 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.415
+ $Y=1.835 $X2=0.54 $Y2=2.95
r34 2 16 400 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.415
+ $Y=1.835 $X2=0.54 $Y2=2.035
r35 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.415
+ $Y=0.365 $X2=0.54 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_1%VPWR 1 6 10 12 19 20 23
r24 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r25 17 23 10.3577 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=1.63 $Y=3.33
+ $X2=1.412 $Y2=3.33
r26 17 19 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.63 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 12 23 10.3577 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.412 $Y2=3.33
r29 12 14 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 10 20 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 10 15 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 10 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 6 9 12.4517 $w=4.33e-07 $l=4.7e-07 $layer=LI1_cond $X=1.412 $Y=2.085
+ $X2=1.412 $Y2=2.555
r34 4 23 1.70358 $w=4.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.412 $Y=3.245
+ $X2=1.412 $Y2=3.33
r35 4 9 18.2801 $w=4.33e-07 $l=6.9e-07 $layer=LI1_cond $X=1.412 $Y=3.245
+ $X2=1.412 $Y2=2.555
r36 1 9 300 $w=1.7e-07 $l=8.22679e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=1.835 $X2=1.44 $Y2=2.555
r37 1 6 600 $w=1.7e-07 $l=4.21871e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=1.835 $X2=1.535 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_1%VGND 1 7 9 12 14 21 22 25
c37 9 0 1.35778e-19 $X=1.615 $Y=1.16
r38 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 19 25 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.402
+ $Y2=0
r40 19 21 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.16
+ $Y2=0
r41 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r42 14 25 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.402
+ $Y2=0
r43 14 16 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=0.24
+ $Y2=0
r44 12 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r45 12 17 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r46 12 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 9 10 4.33665 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=1.16
+ $X2=1.47 $Y2=0.995
r48 7 10 14.0237 $w=4.13e-07 $l=5.05e-07 $layer=LI1_cond $X=1.402 $Y=0.49
+ $X2=1.402 $Y2=0.995
r49 4 25 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.402 $Y=0.085
+ $X2=1.402 $Y2=0
r50 4 7 11.2467 $w=4.13e-07 $l=4.05e-07 $layer=LI1_cond $X=1.402 $Y=0.085
+ $X2=1.402 $Y2=0.49
r51 1 9 182 $w=1.7e-07 $l=9.72651e-07 $layer=licon1_NDIFF $count=1 $X=1.22
+ $Y=0.365 $X2=1.615 $Y2=1.16
r52 1 7 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.22
+ $Y=0.365 $X2=1.36 $Y2=0.49
.ends

