* File: sky130_fd_sc_lp__o2bb2ai_0.pxi.spice
* Created: Fri Aug 28 11:12:26 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2AI_0%A1_N N_A1_N_c_84_n N_A1_N_M1003_g N_A1_N_c_91_n
+ N_A1_N_c_92_n N_A1_N_M1005_g N_A1_N_c_86_n N_A1_N_c_87_n A1_N A1_N A1_N A1_N
+ A1_N A1_N N_A1_N_c_89_n PM_SKY130_FD_SC_LP__O2BB2AI_0%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_0%A2_N N_A2_N_M1000_g N_A2_N_c_130_n
+ N_A2_N_c_131_n N_A2_N_M1001_g N_A2_N_c_127_n A2_N A2_N A2_N A2_N
+ N_A2_N_c_129_n PM_SKY130_FD_SC_LP__O2BB2AI_0%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_0%A_195_56# N_A_195_56#_M1000_d
+ N_A_195_56#_M1005_d N_A_195_56#_c_178_n N_A_195_56#_c_179_n
+ N_A_195_56#_M1009_g N_A_195_56#_M1006_g N_A_195_56#_c_182_n
+ N_A_195_56#_c_191_n N_A_195_56#_c_192_n N_A_195_56#_c_183_n
+ N_A_195_56#_c_184_n N_A_195_56#_c_185_n N_A_195_56#_c_186_n
+ N_A_195_56#_c_187_n N_A_195_56#_c_188_n N_A_195_56#_c_189_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_0%A_195_56#
x_PM_SKY130_FD_SC_LP__O2BB2AI_0%B2 N_B2_M1004_g N_B2_M1007_g N_B2_c_253_n
+ N_B2_c_257_n B2 B2 N_B2_c_255_n PM_SKY130_FD_SC_LP__O2BB2AI_0%B2
x_PM_SKY130_FD_SC_LP__O2BB2AI_0%B1 N_B1_M1008_g N_B1_M1002_g N_B1_c_301_n
+ N_B1_c_302_n N_B1_c_294_n N_B1_c_295_n N_B1_c_296_n N_B1_c_297_n N_B1_c_304_n
+ B1 B1 B1 N_B1_c_299_n PM_SKY130_FD_SC_LP__O2BB2AI_0%B1
x_PM_SKY130_FD_SC_LP__O2BB2AI_0%VPWR N_VPWR_M1005_s N_VPWR_M1001_d
+ N_VPWR_M1008_d N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n N_VPWR_c_341_n
+ VPWR N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n N_VPWR_c_345_n
+ N_VPWR_c_337_n PM_SKY130_FD_SC_LP__O2BB2AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2AI_0%Y N_Y_M1009_s N_Y_M1006_d N_Y_c_384_n
+ N_Y_c_385_n N_Y_c_381_n Y Y N_Y_c_383_n Y PM_SKY130_FD_SC_LP__O2BB2AI_0%Y
x_PM_SKY130_FD_SC_LP__O2BB2AI_0%VGND N_VGND_M1003_s N_VGND_M1007_d
+ N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n VGND N_VGND_c_435_n
+ N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_0%VGND
x_PM_SKY130_FD_SC_LP__O2BB2AI_0%A_400_47# N_A_400_47#_M1009_d
+ N_A_400_47#_M1002_d N_A_400_47#_c_473_n N_A_400_47#_c_474_n
+ N_A_400_47#_c_475_n N_A_400_47#_c_476_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_0%A_400_47#
cc_1 VNB N_A1_N_c_84_n 0.00891946f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.11
cc_2 VNB N_A1_N_M1003_g 0.0232274f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.49
cc_3 VNB N_A1_N_c_86_n 0.0310338f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.99
cc_4 VNB N_A1_N_c_87_n 0.0185667f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_5 VNB A1_N 0.0339238f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A1_N_c_89_n 0.0299899f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_7 VNB N_A2_N_M1000_g 0.0379586f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.84
cc_8 VNB N_A2_N_c_127_n 0.0177479f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_9 VNB A2_N 0.0118135f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.84
cc_10 VNB N_A2_N_c_129_n 0.015539f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.69
cc_11 VNB N_A_195_56#_c_178_n 0.0164807f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.185
cc_12 VNB N_A_195_56#_c_179_n 0.0163515f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=2.185
cc_13 VNB N_A_195_56#_M1009_g 0.0235042f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.735
cc_14 VNB N_A_195_56#_M1006_g 0.036117f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.99
cc_15 VNB N_A_195_56#_c_182_n 0.00556614f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_16 VNB N_A_195_56#_c_183_n 0.00150898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_195_56#_c_184_n 0.00514819f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_18 VNB N_A_195_56#_c_185_n 0.00300654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_195_56#_c_186_n 0.00469837f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.295
cc_20 VNB N_A_195_56#_c_187_n 0.0385445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_195_56#_c_188_n 0.0028439f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=1.665
cc_22 VNB N_A_195_56#_c_189_n 0.00111214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B2_M1007_g 0.0368634f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.185
cc_24 VNB N_B2_c_253_n 0.0215498f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.735
cc_25 VNB B2 0.00602684f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_26 VNB N_B2_c_255_n 0.015621f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_27 VNB N_B1_c_294_n 0.0194855f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_28 VNB N_B1_c_295_n 0.0131616f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_29 VNB N_B1_c_296_n 0.0220493f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_B1_c_297_n 0.0227414f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_31 VNB B1 0.0254248f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_32 VNB N_B1_c_299_n 0.018587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_337_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.237 $Y2=2.775
cc_34 VNB N_Y_c_381_n 0.00403391f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_35 VNB Y 0.00510342f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_36 VNB N_Y_c_383_n 0.00630729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_432_n 0.0118233f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.185
cc_38 VNB N_VGND_c_433_n 0.019822f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.26
cc_39 VNB N_VGND_c_434_n 0.00522139f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_40 VNB N_VGND_c_435_n 0.0545876f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_41 VNB N_VGND_c_436_n 0.0193622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_437_n 0.19969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_438_n 0.00497572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_400_47#_c_473_n 0.00201706f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.26
cc_45 VNB N_A_400_47#_c_474_n 0.0211366f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.735
cc_46 VNB N_A_400_47#_c_475_n 0.00345143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_400_47#_c_476_n 0.020394f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.99
cc_48 VPB N_A1_N_c_84_n 0.0290741f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.11
cc_49 VPB N_A1_N_c_91_n 0.0478784f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.185
cc_50 VPB N_A1_N_c_92_n 0.0121793f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.185
cc_51 VPB N_A1_N_M1005_g 0.0229564f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.735
cc_52 VPB A1_N 0.0644339f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_53 VPB N_A2_N_c_130_n 0.0376814f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.49
cc_54 VPB N_A2_N_c_131_n 0.0102888f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A2_N_M1001_g 0.0371795f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.26
cc_56 VPB N_A2_N_c_127_n 0.00668111f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_57 VPB A2_N 0.00432183f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=0.84
cc_58 VPB N_A_195_56#_M1006_g 0.0488343f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=0.99
cc_59 VPB N_A_195_56#_c_191_n 0.001049f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_60 VPB N_A_195_56#_c_192_n 0.00190422f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_61 VPB N_A_195_56#_c_185_n 0.0113312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_B2_M1004_g 0.0405852f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.84
cc_63 VPB N_B2_c_257_n 0.0179157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB B2 0.00546551f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_65 VPB N_B1_M1008_g 0.0280681f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.84
cc_66 VPB N_B1_c_301_n 0.012313f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.735
cc_67 VPB N_B1_c_302_n 0.0233146f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=0.84
cc_68 VPB N_B1_c_297_n 0.00480911f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_69 VPB N_B1_c_304_n 0.0188836f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_70 VPB B1 0.0291139f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_71 VPB N_VPWR_c_338_n 0.0198391f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=0.84
cc_72 VPB N_VPWR_c_339_n 0.00414834f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_73 VPB N_VPWR_c_340_n 0.0151088f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_74 VPB N_VPWR_c_341_n 0.0329212f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_75 VPB N_VPWR_c_342_n 0.015301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_343_n 0.0254914f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_77 VPB N_VPWR_c_344_n 0.0273137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_345_n 0.00456098f $X=-0.19 $Y=1.655 $X2=0.237 $Y2=2.035
cc_79 VPB N_VPWR_c_337_n 0.0806516f $X=-0.19 $Y=1.655 $X2=0.237 $Y2=2.775
cc_80 VPB N_Y_c_384_n 0.00968624f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.26
cc_81 VPB N_Y_c_385_n 0.00486751f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.735
cc_82 VPB Y 0.00149747f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_83 N_A1_N_M1003_g N_A2_N_M1000_g 0.0444139f $X=0.51 $Y=0.49 $X2=0 $Y2=0
cc_84 A1_N N_A2_N_M1000_g 2.9992e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_85 N_A1_N_c_89_n N_A2_N_M1000_g 0.00638248f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_86 N_A1_N_c_84_n N_A2_N_c_131_n 0.0113237f $X=0.36 $Y=2.11 $X2=0 $Y2=0
cc_87 N_A1_N_c_91_n N_A2_N_c_131_n 0.031464f $X=0.99 $Y=2.185 $X2=0 $Y2=0
cc_88 N_A1_N_c_91_n N_A2_N_M1001_g 0.0175269f $X=0.99 $Y=2.185 $X2=0 $Y2=0
cc_89 N_A1_N_c_87_n N_A2_N_c_127_n 0.0113237f $X=0.27 $Y=1.51 $X2=0 $Y2=0
cc_90 N_A1_N_M1003_g A2_N 5.13607e-19 $X=0.51 $Y=0.49 $X2=0 $Y2=0
cc_91 N_A1_N_c_91_n A2_N 0.0189541f $X=0.99 $Y=2.185 $X2=0 $Y2=0
cc_92 N_A1_N_c_86_n A2_N 0.0041418f $X=0.345 $Y=0.99 $X2=0 $Y2=0
cc_93 A1_N A2_N 0.102177f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_94 N_A1_N_c_89_n A2_N 0.0107225f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_95 A1_N N_A2_N_c_129_n 6.56367e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_96 N_A1_N_c_89_n N_A2_N_c_129_n 0.0113237f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_97 N_A1_N_M1005_g N_A_195_56#_c_191_n 2.31079e-19 $X=1.065 $Y=2.735 $X2=0
+ $Y2=0
cc_98 N_A1_N_M1003_g N_A_195_56#_c_184_n 9.2831e-19 $X=0.51 $Y=0.49 $X2=0 $Y2=0
cc_99 N_A1_N_c_91_n N_A_195_56#_c_185_n 0.00574837f $X=0.99 $Y=2.185 $X2=0 $Y2=0
cc_100 N_A1_N_c_91_n N_VPWR_c_338_n 0.0062554f $X=0.99 $Y=2.185 $X2=0 $Y2=0
cc_101 N_A1_N_M1005_g N_VPWR_c_338_n 0.00388854f $X=1.065 $Y=2.735 $X2=0 $Y2=0
cc_102 A1_N N_VPWR_c_338_n 0.0316398f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_103 N_A1_N_M1005_g N_VPWR_c_339_n 5.73114e-19 $X=1.065 $Y=2.735 $X2=0 $Y2=0
cc_104 N_A1_N_M1005_g N_VPWR_c_342_n 0.00545548f $X=1.065 $Y=2.735 $X2=0 $Y2=0
cc_105 A1_N N_VPWR_c_344_n 0.0125142f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_106 N_A1_N_M1005_g N_VPWR_c_337_n 0.0113151f $X=1.065 $Y=2.735 $X2=0 $Y2=0
cc_107 A1_N N_VPWR_c_337_n 0.011055f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_108 N_A1_N_M1003_g N_VGND_c_433_n 0.0133924f $X=0.51 $Y=0.49 $X2=0 $Y2=0
cc_109 N_A1_N_c_86_n N_VGND_c_433_n 0.00190323f $X=0.345 $Y=0.99 $X2=0 $Y2=0
cc_110 A1_N N_VGND_c_433_n 0.0226729f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_111 N_A1_N_M1003_g N_VGND_c_435_n 0.00448994f $X=0.51 $Y=0.49 $X2=0 $Y2=0
cc_112 N_A1_N_M1003_g N_VGND_c_437_n 0.00779992f $X=0.51 $Y=0.49 $X2=0 $Y2=0
cc_113 A1_N N_VGND_c_437_n 0.00275806f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_114 N_A2_N_M1000_g N_A_195_56#_c_179_n 0.0229155f $X=0.9 $Y=0.49 $X2=0 $Y2=0
cc_115 A2_N N_A_195_56#_c_179_n 0.00141704f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_116 N_A2_N_c_130_n N_A_195_56#_M1006_g 0.0350663f $X=1.42 $Y=1.825 $X2=0
+ $Y2=0
cc_117 N_A2_N_c_130_n N_A_195_56#_c_191_n 0.00127379f $X=1.42 $Y=1.825 $X2=0
+ $Y2=0
cc_118 N_A2_N_M1000_g N_A_195_56#_c_184_n 0.00605075f $X=0.9 $Y=0.49 $X2=0 $Y2=0
cc_119 A2_N N_A_195_56#_c_184_n 0.00318588f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_120 N_A2_N_c_130_n N_A_195_56#_c_185_n 0.013693f $X=1.42 $Y=1.825 $X2=0 $Y2=0
cc_121 N_A2_N_M1001_g N_A_195_56#_c_185_n 0.00842698f $X=1.495 $Y=2.735 $X2=0
+ $Y2=0
cc_122 N_A2_N_c_127_n N_A_195_56#_c_185_n 0.00368369f $X=0.84 $Y=1.75 $X2=0
+ $Y2=0
cc_123 N_A2_N_M1000_g N_A_195_56#_c_186_n 0.00133103f $X=0.9 $Y=0.49 $X2=0 $Y2=0
cc_124 A2_N N_A_195_56#_c_186_n 0.101327f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_125 N_A2_N_c_130_n N_A_195_56#_c_187_n 0.0173335f $X=1.42 $Y=1.825 $X2=0
+ $Y2=0
cc_126 A2_N N_A_195_56#_c_187_n 3.03214e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_127 N_A2_N_c_129_n N_A_195_56#_c_187_n 0.0156447f $X=0.84 $Y=1.395 $X2=0
+ $Y2=0
cc_128 N_A2_N_M1000_g N_A_195_56#_c_188_n 0.00486252f $X=0.9 $Y=0.49 $X2=0 $Y2=0
cc_129 N_A2_N_c_130_n N_A_195_56#_c_189_n 9.64946e-19 $X=1.42 $Y=1.825 $X2=0
+ $Y2=0
cc_130 N_A2_N_c_129_n N_A_195_56#_c_189_n 0.00368369f $X=0.84 $Y=1.395 $X2=0
+ $Y2=0
cc_131 A2_N N_VPWR_c_338_n 0.0230936f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_132 N_A2_N_M1001_g N_VPWR_c_339_n 0.0101941f $X=1.495 $Y=2.735 $X2=0 $Y2=0
cc_133 N_A2_N_M1001_g N_VPWR_c_342_n 0.00489337f $X=1.495 $Y=2.735 $X2=0 $Y2=0
cc_134 N_A2_N_M1001_g N_VPWR_c_337_n 0.00879071f $X=1.495 $Y=2.735 $X2=0 $Y2=0
cc_135 N_A2_N_M1001_g N_Y_c_384_n 0.00388533f $X=1.495 $Y=2.735 $X2=0 $Y2=0
cc_136 N_A2_N_M1000_g N_Y_c_381_n 7.64997e-19 $X=0.9 $Y=0.49 $X2=0 $Y2=0
cc_137 N_A2_N_c_130_n Y 0.00435942f $X=1.42 $Y=1.825 $X2=0 $Y2=0
cc_138 N_A2_N_M1001_g Y 0.00230347f $X=1.495 $Y=2.735 $X2=0 $Y2=0
cc_139 N_A2_N_M1000_g N_VGND_c_433_n 0.0021062f $X=0.9 $Y=0.49 $X2=0 $Y2=0
cc_140 N_A2_N_M1000_g N_VGND_c_435_n 0.00507563f $X=0.9 $Y=0.49 $X2=0 $Y2=0
cc_141 N_A2_N_M1000_g N_VGND_c_437_n 0.00671799f $X=0.9 $Y=0.49 $X2=0 $Y2=0
cc_142 A2_N N_VGND_c_437_n 0.0139997f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_143 N_A_195_56#_M1006_g N_B2_M1004_g 0.031752f $X=1.925 $Y=2.735 $X2=0 $Y2=0
cc_144 N_A_195_56#_M1009_g N_B2_M1007_g 0.0244085f $X=1.925 $Y=0.445 $X2=0 $Y2=0
cc_145 N_A_195_56#_M1006_g B2 0.00493764f $X=1.925 $Y=2.735 $X2=0 $Y2=0
cc_146 N_A_195_56#_M1006_g N_B2_c_255_n 0.0329331f $X=1.925 $Y=2.735 $X2=0 $Y2=0
cc_147 N_A_195_56#_c_191_n N_VPWR_c_338_n 0.00225185f $X=1.267 $Y=2.512 $X2=0
+ $Y2=0
cc_148 N_A_195_56#_M1006_g N_VPWR_c_339_n 0.0109643f $X=1.925 $Y=2.735 $X2=0
+ $Y2=0
cc_149 N_A_195_56#_c_191_n N_VPWR_c_339_n 0.026007f $X=1.267 $Y=2.512 $X2=0
+ $Y2=0
cc_150 N_A_195_56#_c_192_n N_VPWR_c_342_n 0.0157066f $X=1.28 $Y=2.56 $X2=0 $Y2=0
cc_151 N_A_195_56#_M1006_g N_VPWR_c_343_n 0.00489337f $X=1.925 $Y=2.735 $X2=0
+ $Y2=0
cc_152 N_A_195_56#_M1006_g N_VPWR_c_337_n 0.00879071f $X=1.925 $Y=2.735 $X2=0
+ $Y2=0
cc_153 N_A_195_56#_c_192_n N_VPWR_c_337_n 0.00901482f $X=1.28 $Y=2.56 $X2=0
+ $Y2=0
cc_154 N_A_195_56#_M1006_g N_Y_c_384_n 0.0173543f $X=1.925 $Y=2.735 $X2=0 $Y2=0
cc_155 N_A_195_56#_c_185_n N_Y_c_384_n 0.0135323f $X=1.267 $Y=2.395 $X2=0 $Y2=0
cc_156 N_A_195_56#_M1006_g N_Y_c_385_n 0.0033809f $X=1.925 $Y=2.735 $X2=0 $Y2=0
cc_157 N_A_195_56#_c_185_n N_Y_c_385_n 0.00663916f $X=1.267 $Y=2.395 $X2=0 $Y2=0
cc_158 N_A_195_56#_c_178_n N_Y_c_381_n 0.00765056f $X=1.85 $Y=0.885 $X2=0 $Y2=0
cc_159 N_A_195_56#_M1009_g N_Y_c_381_n 0.00436063f $X=1.925 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_195_56#_c_184_n N_Y_c_381_n 0.0233358f $X=1.28 $Y=0.49 $X2=0 $Y2=0
cc_161 N_A_195_56#_c_178_n Y 0.0021943f $X=1.85 $Y=0.885 $X2=0 $Y2=0
cc_162 N_A_195_56#_M1006_g Y 0.0132025f $X=1.925 $Y=2.735 $X2=0 $Y2=0
cc_163 N_A_195_56#_c_185_n Y 0.0331423f $X=1.267 $Y=2.395 $X2=0 $Y2=0
cc_164 N_A_195_56#_c_178_n N_Y_c_383_n 0.0069321f $X=1.85 $Y=0.885 $X2=0 $Y2=0
cc_165 N_A_195_56#_M1009_g N_Y_c_383_n 0.00537096f $X=1.925 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A_195_56#_M1006_g N_Y_c_383_n 0.0135163f $X=1.925 $Y=2.735 $X2=0 $Y2=0
cc_167 N_A_195_56#_c_182_n N_Y_c_383_n 0.0018089f $X=1.925 $Y=0.885 $X2=0 $Y2=0
cc_168 N_A_195_56#_c_184_n N_Y_c_383_n 0.00205405f $X=1.28 $Y=0.49 $X2=0 $Y2=0
cc_169 N_A_195_56#_c_185_n N_Y_c_383_n 0.00763031f $X=1.267 $Y=2.395 $X2=0 $Y2=0
cc_170 N_A_195_56#_c_186_n N_Y_c_383_n 0.0419897f $X=1.38 $Y=0.975 $X2=0 $Y2=0
cc_171 N_A_195_56#_c_187_n N_Y_c_383_n 0.00351427f $X=1.38 $Y=0.975 $X2=0 $Y2=0
cc_172 N_A_195_56#_c_188_n N_Y_c_383_n 0.00692493f $X=1.37 $Y=0.81 $X2=0 $Y2=0
cc_173 N_A_195_56#_c_184_n N_VGND_c_433_n 0.0105995f $X=1.28 $Y=0.49 $X2=0 $Y2=0
cc_174 N_A_195_56#_M1009_g N_VGND_c_435_n 0.00518687f $X=1.925 $Y=0.445 $X2=0
+ $Y2=0
cc_175 N_A_195_56#_c_184_n N_VGND_c_435_n 0.017892f $X=1.28 $Y=0.49 $X2=0 $Y2=0
cc_176 N_A_195_56#_M1009_g N_VGND_c_437_n 0.0108337f $X=1.925 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_A_195_56#_c_184_n N_VGND_c_437_n 0.0150726f $X=1.28 $Y=0.49 $X2=0 $Y2=0
cc_178 N_A_195_56#_c_186_n N_VGND_c_437_n 0.00646009f $X=1.38 $Y=0.975 $X2=0
+ $Y2=0
cc_179 N_A_195_56#_M1009_g N_A_400_47#_c_473_n 0.00214944f $X=1.925 $Y=0.445
+ $X2=0 $Y2=0
cc_180 N_A_195_56#_M1009_g N_A_400_47#_c_475_n 0.00170671f $X=1.925 $Y=0.445
+ $X2=0 $Y2=0
cc_181 N_B2_M1004_g N_B1_c_302_n 0.0569463f $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_182 N_B2_M1007_g N_B1_c_294_n 0.0190622f $X=2.395 $Y=0.445 $X2=0 $Y2=0
cc_183 N_B2_M1007_g N_B1_c_296_n 0.00957013f $X=2.395 $Y=0.445 $X2=0 $Y2=0
cc_184 B2 N_B1_c_296_n 0.00249909f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_185 N_B2_c_255_n N_B1_c_296_n 0.0118636f $X=2.405 $Y=1.32 $X2=0 $Y2=0
cc_186 N_B2_c_257_n N_B1_c_297_n 0.0118636f $X=2.405 $Y=1.825 $X2=0 $Y2=0
cc_187 N_B2_M1004_g N_B1_c_304_n 0.0077026f $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_188 N_B2_M1004_g B1 0.00143082f $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_189 B2 B1 0.0274435f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_190 N_B2_c_255_n B1 0.00226679f $X=2.405 $Y=1.32 $X2=0 $Y2=0
cc_191 N_B2_c_253_n N_B1_c_299_n 0.0118636f $X=2.405 $Y=1.66 $X2=0 $Y2=0
cc_192 N_B2_M1004_g N_VPWR_c_339_n 0.00104684f $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_193 N_B2_M1004_g N_VPWR_c_341_n 0.00280799f $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_194 N_B2_M1004_g N_VPWR_c_343_n 0.00511657f $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_195 N_B2_M1004_g N_VPWR_c_337_n 0.00961146f $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_196 N_B2_M1004_g N_Y_c_384_n 0.00549575f $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_197 N_B2_c_257_n N_Y_c_384_n 2.75182e-19 $X=2.405 $Y=1.825 $X2=0 $Y2=0
cc_198 B2 N_Y_c_384_n 0.0190483f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_199 N_B2_M1004_g N_Y_c_385_n 0.0175754f $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_200 N_B2_M1004_g Y 9.08855e-19 $X=2.355 $Y=2.735 $X2=0 $Y2=0
cc_201 N_B2_M1007_g N_Y_c_383_n 0.00105411f $X=2.395 $Y=0.445 $X2=0 $Y2=0
cc_202 B2 N_Y_c_383_n 0.0552671f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_203 N_B2_M1007_g N_VGND_c_434_n 0.00319241f $X=2.395 $Y=0.445 $X2=0 $Y2=0
cc_204 N_B2_M1007_g N_VGND_c_435_n 0.00585385f $X=2.395 $Y=0.445 $X2=0 $Y2=0
cc_205 N_B2_M1007_g N_VGND_c_437_n 0.00628213f $X=2.395 $Y=0.445 $X2=0 $Y2=0
cc_206 N_B2_M1007_g N_A_400_47#_c_473_n 0.00188931f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_B2_M1007_g N_A_400_47#_c_474_n 0.0115421f $X=2.395 $Y=0.445 $X2=0 $Y2=0
cc_208 B2 N_A_400_47#_c_474_n 0.0143032f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_209 N_B2_c_255_n N_A_400_47#_c_474_n 0.00341934f $X=2.405 $Y=1.32 $X2=0 $Y2=0
cc_210 B2 N_A_400_47#_c_475_n 0.0224289f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_211 N_B2_c_255_n N_A_400_47#_c_475_n 4.59403e-19 $X=2.405 $Y=1.32 $X2=0 $Y2=0
cc_212 N_B1_M1008_g N_VPWR_c_341_n 0.0182446f $X=2.745 $Y=2.735 $X2=0 $Y2=0
cc_213 N_B1_c_302_n N_VPWR_c_341_n 0.00528274f $X=2.885 $Y=2.14 $X2=0 $Y2=0
cc_214 N_B1_c_304_n N_VPWR_c_341_n 6.58127e-19 $X=2.975 $Y=1.88 $X2=0 $Y2=0
cc_215 B1 N_VPWR_c_341_n 0.0194818f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_216 N_B1_M1008_g N_VPWR_c_343_n 0.00452967f $X=2.745 $Y=2.735 $X2=0 $Y2=0
cc_217 N_B1_M1008_g N_VPWR_c_337_n 0.00809218f $X=2.745 $Y=2.735 $X2=0 $Y2=0
cc_218 N_B1_c_302_n N_Y_c_384_n 3.56836e-19 $X=2.885 $Y=2.14 $X2=0 $Y2=0
cc_219 B1 N_Y_c_384_n 0.00485898f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_220 N_B1_c_302_n N_Y_c_385_n 0.00295391f $X=2.885 $Y=2.14 $X2=0 $Y2=0
cc_221 B1 N_Y_c_385_n 6.74009e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_222 N_B1_c_294_n N_VGND_c_434_n 0.00313081f $X=2.855 $Y=0.765 $X2=0 $Y2=0
cc_223 N_B1_c_294_n N_VGND_c_436_n 0.00585385f $X=2.855 $Y=0.765 $X2=0 $Y2=0
cc_224 N_B1_c_295_n N_VGND_c_436_n 2.3855e-19 $X=2.855 $Y=0.915 $X2=0 $Y2=0
cc_225 N_B1_c_294_n N_VGND_c_437_n 0.00724162f $X=2.855 $Y=0.765 $X2=0 $Y2=0
cc_226 N_B1_c_295_n N_A_400_47#_c_474_n 0.0110093f $X=2.855 $Y=0.915 $X2=0 $Y2=0
cc_227 N_B1_c_296_n N_A_400_47#_c_474_n 0.00611111f $X=2.975 $Y=1.21 $X2=0 $Y2=0
cc_228 B1 N_A_400_47#_c_474_n 0.0286117f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_229 N_B1_c_299_n N_A_400_47#_c_474_n 0.00111322f $X=2.975 $Y=1.375 $X2=0
+ $Y2=0
cc_230 N_B1_c_294_n N_A_400_47#_c_476_n 0.0036232f $X=2.855 $Y=0.765 $X2=0 $Y2=0
cc_231 N_B1_c_295_n N_A_400_47#_c_476_n 0.00178905f $X=2.855 $Y=0.915 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_339_n N_Y_c_384_n 0.0214598f $X=1.71 $Y=2.56 $X2=0 $Y2=0
cc_233 N_VPWR_c_339_n N_Y_c_385_n 0.0260305f $X=1.71 $Y=2.56 $X2=0 $Y2=0
cc_234 N_VPWR_c_341_n N_Y_c_385_n 0.0209047f $X=2.96 $Y=2.56 $X2=0 $Y2=0
cc_235 N_VPWR_c_343_n N_Y_c_385_n 0.0179866f $X=2.795 $Y=3.33 $X2=0 $Y2=0
cc_236 N_VPWR_c_337_n N_Y_c_385_n 0.0102592f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_237 N_Y_c_381_n N_VGND_c_435_n 0.0184511f $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_238 N_Y_M1009_s N_VGND_c_437_n 0.0021695f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_239 N_Y_c_381_n N_VGND_c_437_n 0.0129536f $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_240 N_Y_c_381_n N_A_400_47#_c_473_n 0.0250862f $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_241 N_Y_c_383_n N_A_400_47#_c_473_n 0.0123984f $X=1.725 $Y=1.57 $X2=0 $Y2=0
cc_242 N_Y_c_383_n N_A_400_47#_c_475_n 0.0136802f $X=1.725 $Y=1.57 $X2=0 $Y2=0
cc_243 N_VGND_c_437_n N_A_400_47#_M1009_d 0.00495563f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_244 N_VGND_c_437_n N_A_400_47#_M1002_d 0.00218933f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_245 N_VGND_c_435_n N_A_400_47#_c_473_n 0.0131849f $X=2.475 $Y=0 $X2=0 $Y2=0
cc_246 N_VGND_c_437_n N_A_400_47#_c_473_n 0.00913662f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_247 N_VGND_c_434_n N_A_400_47#_c_474_n 0.0166313f $X=2.61 $Y=0.445 $X2=0
+ $Y2=0
cc_248 N_VGND_c_437_n N_A_400_47#_c_474_n 0.0110596f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_249 N_VGND_c_436_n N_A_400_47#_c_476_n 0.0165706f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_250 N_VGND_c_437_n N_A_400_47#_c_476_n 0.01144f $X=3.12 $Y=0 $X2=0 $Y2=0
