* File: sky130_fd_sc_lp__mux2_lp2.spice
* Created: Wed Sep  2 10:00:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2_lp2.pex.spice"
.subckt sky130_fd_sc_lp__mux2_lp2  VNB VPB A1 A0 S X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* S	S
* A0	A0
* A1	A1
* VPB	VPB
* VNB	VNB
MM1001 A_115_57# N_A_84_259#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.9 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_84_259#_M1007_g A_115_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1386 AS=0.0441 PD=1.08 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1012 A_349_57# N_A_182_303#_M1012_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1386 PD=0.66 PS=1.08 NRD=18.564 NRS=108.564 M=1 R=2.8
+ SA=75001.4 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1006 N_A_84_259#_M1006_d N_A0_M1006_g A_349_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.13965 AS=0.0504 PD=1.085 PS=0.66 NRD=109.992 NRS=18.564 M=1 R=2.8
+ SA=75001.8 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1004 A_590_57# N_A1_M1004_g N_A_84_259#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.13965 PD=0.77 PS=1.085 NRD=34.284 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_S_M1002_g A_590_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=34.284 M=1 R=2.8 SA=75003.1 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1008 A_776_57# N_S_M1008_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.5 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_182_303#_M1009_d N_S_M1009_g A_776_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_84_259#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.25 W=1
+ AD=0.305 AS=0.285 PD=1.61 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1011 A_306_401# N_A_182_303#_M1011_g N_VPWR_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.305 PD=1.24 PS=1.61 NRD=12.7853 NRS=65.01 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1003 N_A_84_259#_M1003_d N_A1_M1003_g A_306_401# VPB PHIGHVT L=0.25 W=1
+ AD=0.16 AS=0.12 PD=1.32 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125002 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1000 A_518_401# N_A0_M1000_g N_A_84_259#_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.16 PD=1.24 PS=1.32 NRD=12.7853 NRS=7.8603 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_S_M1005_g A_518_401# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125003 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1013 N_A_182_303#_M1013_d N_S_M1013_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__mux2_lp2.pxi.spice"
*
.ends
*
*
