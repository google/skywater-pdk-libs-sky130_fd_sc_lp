* File: sky130_fd_sc_lp__mux4_4.spice
* Created: Fri Aug 28 10:46:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux4_4.pex.spice"
.subckt sky130_fd_sc_lp__mux4_4  VNB VPB S1 A1 A0 A3 A2 S0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S0	S0
* A2	A2
* A3	A3
* A0	A0
* A1	A1
* S1	S1
* VPB	VPB
* VNB	VNB
MM1008 N_A_114_119#_M1008_d N_S1_M1008_g N_A_27_119#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_200_119#_M1006_d N_A_84_277#_M1006_g N_A_114_119#_M1008_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_S1_M1007_g N_A_84_277#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1197 PD=0.913333 PS=1.41 NRD=60 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75006.4 A=0.063 P=1.14 MULT=1
MM1014 N_X_M1014_d N_A_114_119#_M1014_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=1.82667 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75004 A=0.126 P=1.98 MULT=1
MM1015 N_X_M1014_d N_A_114_119#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001 SB=75003.5
+ A=0.126 P=1.98 MULT=1
MM1024 N_X_M1024_d N_A_114_119#_M1024_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1027 N_X_M1024_d N_A_114_119#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1834 PD=1.12 PS=1.64 NRD=0 NRS=0 M=1 R=5.6 SA=75001.8
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1001 A_952_119# N_A1_M1001_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0917 PD=0.63 PS=0.82 NRD=14.28 NRS=31.428 M=1 R=2.8 SA=75002.6 SB=75004.6
+ A=0.063 P=1.14 MULT=1
MM1029 N_A_200_119#_M1029_d N_S0_M1029_g A_952_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003
+ SB=75004.3 A=0.063 P=1.14 MULT=1
MM1002 A_1110_119# N_A_1041_333#_M1002_g N_A_200_119#_M1029_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.4
+ SB=75003.8 A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_A0_M1030_g A_1110_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.177975 AS=0.0441 PD=1.3 PS=0.63 NRD=24.276 NRS=14.28 M=1 R=2.8 SA=75003.8
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1025 A_1367_119# N_A3_M1025_g N_VGND_M1030_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.177975 PD=0.63 PS=1.3 NRD=14.28 NRS=120 M=1 R=2.8 SA=75004.7
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1017 N_A_27_119#_M1017_d N_S0_M1017_g A_1367_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75005.1
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1023 A_1525_119# N_A_1041_333#_M1023_g N_A_27_119#_M1017_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75005.5
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_A2_M1028_g A_1525_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.19425 AS=0.0672 PD=1.345 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75006
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1021 N_A_1041_333#_M1021_d N_S0_M1021_g N_VGND_M1028_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.19425 PD=1.41 PS=1.345 NRD=5.712 NRS=184.284 M=1 R=2.8
+ SA=75007 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_A_114_119#_M1031_d N_A_84_277#_M1031_g N_A_27_119#_M1031_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=6.1464 M=1
+ R=4.26667 SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1009 N_A_200_119#_M1009_d N_S1_M1009_g N_A_114_119#_M1031_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_S1_M1016_g N_A_84_277#_M1016_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.144674 AS=0.24375 PD=1.11495 PS=2.28 NRD=52.6384 NRS=66.1723 M=1
+ R=4.26667 SA=75000.3 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1016_d N_A_114_119#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.284826 AS=0.1764 PD=2.19505 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75003.9 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_114_119#_M1011_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001 SB=75003.5
+ A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1011_d N_A_114_119#_M1018_g N_X_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.4
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_A_114_119#_M1022_g N_X_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.581788 AS=0.1764 PD=2.69905 PS=1.54 NRD=54.7069 NRS=0 M=1 R=8.4
+ SA=75001.8 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1004 A_999_431# N_A1_M1004_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.295512 PD=0.85 PS=1.37095 NRD=15.3857 NRS=45.3888 M=1 R=4.26667
+ SA=75002.6 SB=75003.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_200_119#_M1000_d N_A_1041_333#_M1000_g A_999_431# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75003 SB=75003.4 A=0.096 P=1.58 MULT=1
MM1020 A_1157_431# N_S0_M1020_g N_A_200_119#_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1194 AS=0.0896 PD=1.06 PS=0.92 NRD=40.4835 NRS=0 M=1 R=4.26667 SA=75003.4
+ SB=75003 A=0.096 P=1.58 MULT=1
MM1019 N_VPWR_M1019_d N_A0_M1019_g A_1157_431# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1194 PD=1.21 PS=1.06 NRD=0 NRS=40.4835 M=1 R=4.26667 SA=75003.6
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1012 A_1403_419# N_A3_M1012_g N_VPWR_M1019_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.21 NRD=15.3857 NRS=89.2607 M=1 R=4.26667
+ SA=75004.3 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1013 N_A_27_119#_M1013_d N_A_1041_333#_M1013_g A_1403_419# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.13785 AS=0.0672 PD=1.12 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75004.7 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1010 A_1589_431# N_S0_M1010_g N_A_27_119#_M1013_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1194 AS=0.13785 PD=1.06 PS=1.12 NRD=40.4835 NRS=43.0839 M=1 R=4.26667
+ SA=75005.1 SB=75001 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g A_1589_431# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1194 PD=0.92 PS=1.06 NRD=0 NRS=40.4835 M=1 R=4.26667 SA=75005.5
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1026 N_A_1041_333#_M1026_d N_S0_M1026_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75006
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX32_noxref VNB VPB NWDIODE A=19.1263 P=24.01
c_97 VNB 0 1.9535e-19 $X=0 $Y=0
c_1287 A_999_431# 0 8.77531e-20 $X=4.995 $Y=2.155
c_1415 A_1110_119# 0 4.44719e-20 $X=5.55 $Y=0.595
*
.include "sky130_fd_sc_lp__mux4_4.pxi.spice"
*
.ends
*
*
