* File: sky130_fd_sc_lp__dlclkp_lp.spice
* Created: Wed Sep  2 09:46:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlclkp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dlclkp_lp  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1013 A_110_47# N_A_80_21#_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_80_21#_M1000_g A_110_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0441 PD=0.78 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1009 A_284_47# N_GATE_M1009_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=22.848 M=1 R=2.8 SA=75001.1
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1010 N_A_352_419#_M1010_d N_A_80_21#_M1010_g A_284_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1022 A_448_47# N_A_27_47#_M1022_g N_A_352_419#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1428 AS=0.0588 PD=1.1 PS=0.7 NRD=81.42 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_584_21#_M1011_g A_448_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1428 PD=0.7 PS=1.1 NRD=0 NRS=81.42 M=1 R=2.8 SA=75002.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1019 A_700_47# N_A_352_419#_M1019_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75003.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1023 N_A_584_21#_M1023_d N_A_352_419#_M1023_g A_700_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 A_923_185# N_CLK_M1016_g N_A_80_21#_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.1197 PD=0.745 PS=1.41 NRD=30.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_CLK_M1014_g A_923_185# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.06825 PD=0.7 PS=0.745 NRD=0 NRS=30.708 M=1 R=2.8 SA=75000.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1017 A_1104_185# N_CLK_M1017_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_1147_419#_M1005_d N_A_584_21#_M1005_g A_1104_185# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_1284_47# N_A_1147_419#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_GCLK_M1006_d N_A_1147_419#_M1006_g A_1284_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_80_21#_M1003_g N_A_27_47#_M1003_s VPB PHIGHVT L=0.25
+ W=1 AD=0.16 AS=0.285 PD=1.32 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1007 A_254_419# N_GATE_M1007_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.16 PD=1.24 PS=1.32 NRD=12.7853 NRS=7.8603 M=1 R=4 SA=125001 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1018 N_A_352_419#_M1018_d N_A_27_47#_M1018_g A_254_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.31 AS=0.12 PD=1.62 PS=1.24 NRD=66.98 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1012 A_526_419# N_A_80_21#_M1012_g N_A_352_419#_M1018_d VPB PHIGHVT L=0.25 W=1
+ AD=0.16 AS=0.31 PD=1.32 PS=1.62 NRD=20.6653 NRS=0 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A_584_21#_M1001_g A_526_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.1775 AS=0.16 PD=1.355 PS=1.32 NRD=0.9653 NRS=20.6653 M=1 R=4 SA=125003
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1015 N_A_584_21#_M1015_d N_A_352_419#_M1015_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.1775 PD=2.57 PS=1.355 NRD=0 NRS=13.7703 M=1 R=4
+ SA=125003 SB=125000 A=0.25 P=2.5 MULT=1
MM1020 N_VPWR_M1020_d N_CLK_M1020_g N_A_80_21#_M1020_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1008 N_A_1147_419#_M1008_d N_CLK_M1008_g N_VPWR_M1020_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_584_21#_M1004_g N_A_1147_419#_M1008_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1021 N_GCLK_M1021_d N_A_1147_419#_M1021_g N_VPWR_M1004_d VPB PHIGHVT L=0.25
+ W=1 AD=0.27 AS=0.14 PD=2.54 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.7419 P=19.41
*
.include "sky130_fd_sc_lp__dlclkp_lp.pxi.spice"
*
.ends
*
*
