* File: sky130_fd_sc_lp__einvp_lp.pex.spice
* Created: Wed Sep  2 09:52:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVP_LP%A 1 3 8 10 11 15
r24 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=0.43
+ $X2=0.505 $Y2=0.595
r25 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.505
+ $Y=0.43 $X2=0.505 $Y2=0.43
r26 11 16 8.43408 $w=3.11e-07 $l=2.15e-07 $layer=LI1_cond $X=0.72 $Y=0.467
+ $X2=0.505 $Y2=0.467
r27 10 16 10.3955 $w=3.11e-07 $l=2.65e-07 $layer=LI1_cond $X=0.24 $Y=0.467
+ $X2=0.505 $Y2=0.467
r28 8 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.595 $Y=0.915
+ $X2=0.595 $Y2=1.235
r29 8 18 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.595 $Y=0.915
+ $X2=0.595 $Y2=0.595
r30 1 9 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.545 $Y=1.36
+ $X2=0.545 $Y2=1.235
r31 1 3 306.84 $w=2.5e-07 $l=1.235e-06 $layer=POLY_cond $X=0.545 $Y=1.36
+ $X2=0.545 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_LP%A_182_321# 1 2 9 11 15 19 21 25 27
r42 25 30 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.77
+ $X2=1.075 $Y2=1.935
r43 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.075
+ $Y=1.77 $X2=1.075 $Y2=1.77
r44 21 24 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.075 $Y=1.69 $X2=1.075
+ $Y2=1.77
r45 17 27 3.03453 $w=3.12e-07 $l=9.31128e-08 $layer=LI1_cond $X=2.132 $Y=1.605
+ $X2=2.115 $Y2=1.69
r46 17 19 34.7686 $w=2.93e-07 $l=8.9e-07 $layer=LI1_cond $X=2.132 $Y=1.605
+ $X2=2.132 $Y2=0.715
r47 13 27 3.03453 $w=3.12e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=1.775
+ $X2=2.115 $Y2=1.69
r48 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.115 $Y=1.775
+ $X2=2.115 $Y2=2.24
r49 12 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=1.69
+ $X2=1.075 $Y2=1.69
r50 11 27 3.60271 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=1.69
+ $X2=2.115 $Y2=1.69
r51 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.95 $Y=1.69
+ $X2=1.24 $Y2=1.69
r52 9 30 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.035 $Y=2.595
+ $X2=1.035 $Y2=1.935
r53 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.975
+ $Y=2.095 $X2=2.115 $Y2=2.24
r54 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.505 $X2=2.07 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_LP%TE 1 3 5 6 8 11 13 15 16 17 18 23 28
r42 27 28 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.85 $Y=1.2 $X2=1.855
+ $Y2=1.2
r43 25 27 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.63 $Y=1.2 $X2=1.85
+ $Y2=1.2
r44 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.2 $X2=1.63 $Y2=1.2
r45 22 25 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=1.495 $Y=1.2
+ $X2=1.63 $Y2=1.2
r46 22 23 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.495 $Y=1.2 $X2=1.42
+ $Y2=1.2
r47 18 26 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.63 $Y=1.295
+ $X2=1.63 $Y2=1.2
r48 17 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.63 $Y=0.925
+ $X2=1.63 $Y2=1.2
r49 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.63 $Y=0.555
+ $X2=1.63 $Y2=0.925
r50 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.035
+ $X2=1.855 $Y2=1.2
r51 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.855 $Y=1.035
+ $X2=1.855 $Y2=0.715
r52 9 27 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.365
+ $X2=1.85 $Y2=1.2
r53 9 11 305.598 $w=2.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.85 $Y=1.365
+ $X2=1.85 $Y2=2.595
r54 6 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.035
+ $X2=1.495 $Y2=1.2
r55 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.495 $Y=1.035
+ $X2=1.495 $Y2=0.715
r56 5 23 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.06 $Y=1.275
+ $X2=1.42 $Y2=1.275
r57 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.985 $Y=1.2
+ $X2=1.06 $Y2=1.275
r58 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.985 $Y=1.2 $X2=0.985
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_LP%Z 1 2 7 8 9 10 11 18
r15 10 11 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=2.405
+ $X2=0.29 $Y2=2.775
r16 10 27 5.43295 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.29 $Y=2.405
+ $X2=0.29 $Y2=2.24
r17 9 27 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.29 $Y=2.035
+ $X2=0.29 $Y2=2.24
r18 8 9 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=2.035
r19 7 8 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295 $X2=0.29
+ $Y2=1.665
r20 7 18 9.21954 $w=3.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.015
r21 2 27 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.24
r22 1 18 182 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.705 $X2=0.3 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_LP%VPWR 1 6 11 12 13 23 24
r23 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r24 16 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r25 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r26 13 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 13 17 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 13 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r29 11 20 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.42 $Y=3.33 $X2=1.2
+ $Y2=3.33
r30 11 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=3.33
+ $X2=1.585 $Y2=3.33
r31 10 23 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.75 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 10 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.75 $Y=3.33
+ $X2=1.585 $Y2=3.33
r33 6 9 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.585 $Y=2.24 $X2=1.585
+ $Y2=2.95
r34 4 12 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=3.245
+ $X2=1.585 $Y2=3.33
r35 4 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.585 $Y=3.245
+ $X2=1.585 $Y2=2.95
r36 1 9 400 $w=1.7e-07 $l=1.04614e-06 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=2.095 $X2=1.585 $Y2=2.95
r37 1 6 400 $w=1.7e-07 $l=4.92189e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=2.095 $X2=1.585 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_LP%VGND 1 6 8 10 17 18 21
r30 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r31 15 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.16
+ $Y2=0
r32 15 17 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=2.16
+ $Y2=0
r33 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r34 10 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.16
+ $Y2=0
r35 10 12 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.72
+ $Y2=0
r36 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r37 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r38 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r39 4 21 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0
r40 4 6 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.16 $Y=0.085 $X2=1.16
+ $Y2=0.915
r41 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.705 $X2=1.2 $Y2=0.915
.ends

