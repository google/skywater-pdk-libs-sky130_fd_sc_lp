* File: sky130_fd_sc_lp__mux2_2.spice
* Created: Fri Aug 28 10:43:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2_2.pex.spice"
.subckt sky130_fd_sc_lp__mux2_2  VNB VPB A0 A1 S VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1007 N_X_M1007_d N_A_86_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1007_d N_A_86_21#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2228 PD=1.12 PS=1.78 NRD=0 NRS=9.276 M=1 R=5.6 SA=75000.6
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1001 A_319_48# N_A_284_279#_M1001_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1114 PD=0.63 PS=0.89 NRD=14.28 NRS=28.56 M=1 R=2.8 SA=75001.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1013 N_A_86_21#_M1013_d N_A0_M1013_g A_319_48# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=2.856 NRS=14.28 M=1 R=2.8 SA=75001.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1005 A_499_48# N_A1_M1005_g N_A_86_21#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=28.56 M=1 R=2.8 SA=75002.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_S_M1003_g A_499_48# VNB NSHORT L=0.15 W=0.42 AD=0.08505
+ AS=0.0441 PD=0.825 PS=0.63 NRD=21.42 NRS=14.28 M=1 R=2.8 SA=75002.5 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_284_279#_M1009_d N_S_M1009_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.08505 PD=1.37 PS=0.825 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_86_21#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1011 N_X_M1006_d N_A_86_21#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.358536 PD=1.54 PS=2.45368 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1000 A_350_449# N_A_284_279#_M1000_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.182114 PD=0.85 PS=1.24632 NRD=15.3857 NRS=70.6442 M=1 R=4.26667
+ SA=75001.4 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1010 N_A_86_21#_M1010_d N_A1_M1010_g A_350_449# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.7
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1004 A_508_449# N_A0_M1004_g N_A_86_21#_M1010_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=32.308 NRS=0 M=1 R=4.26667 SA=75002.1
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_S_M1002_g A_508_449# VPB PHIGHVT L=0.15 W=0.64 AD=0.0896
+ AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=32.308 M=1 R=4.26667 SA=75002.6 SB=75000.6
+ A=0.096 P=1.58 MULT=1
MM1012 N_A_284_279#_M1012_d N_S_M1012_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__mux2_2.pxi.spice"
*
.ends
*
*
