* File: sky130_fd_sc_lp__sdfstp_lp.pxi.spice
* Created: Fri Aug 28 11:30:03 2020
* 
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%SCE N_SCE_M1006_g N_SCE_M1017_g N_SCE_M1004_g
+ N_SCE_M1044_g N_SCE_M1018_g N_SCE_c_320_n N_SCE_c_321_n N_SCE_c_322_n
+ N_SCE_c_323_n N_SCE_c_324_n N_SCE_c_332_n N_SCE_c_325_n SCE SCE N_SCE_c_326_n
+ N_SCE_c_327_n N_SCE_c_328_n PM_SKY130_FD_SC_LP__SDFSTP_LP%SCE
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_27_409# N_A_27_409#_M1017_s
+ N_A_27_409#_M1006_s N_A_27_409#_M1016_g N_A_27_409#_c_412_n
+ N_A_27_409#_c_413_n N_A_27_409#_M1022_g N_A_27_409#_c_414_n
+ N_A_27_409#_c_415_n N_A_27_409#_c_416_n N_A_27_409#_c_417_n
+ N_A_27_409#_c_424_n N_A_27_409#_c_418_n N_A_27_409#_c_419_n
+ N_A_27_409#_c_420_n PM_SKY130_FD_SC_LP__SDFSTP_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%D N_D_M1001_g N_D_M1023_g D D N_D_c_483_n
+ PM_SKY130_FD_SC_LP__SDFSTP_LP%D
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%SCD N_SCD_c_522_n N_SCD_M1024_g N_SCD_M1000_g
+ N_SCD_c_523_n SCD SCD N_SCD_c_525_n N_SCD_c_526_n
+ PM_SKY130_FD_SC_LP__SDFSTP_LP%SCD
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%CLK N_CLK_M1041_g N_CLK_c_573_n N_CLK_M1002_g
+ N_CLK_M1029_g N_CLK_c_575_n CLK N_CLK_c_577_n
+ PM_SKY130_FD_SC_LP__SDFSTP_LP%CLK
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_986_409# N_A_986_409#_M1030_d
+ N_A_986_409#_M1035_d N_A_986_409#_M1019_g N_A_986_409#_M1045_g
+ N_A_986_409#_M1042_g N_A_986_409#_M1013_g N_A_986_409#_c_640_n
+ N_A_986_409#_c_641_n N_A_986_409#_c_642_n N_A_986_409#_c_643_n
+ N_A_986_409#_c_627_n N_A_986_409#_c_628_n N_A_986_409#_c_654_p
+ N_A_986_409#_c_655_p N_A_986_409#_c_649_p N_A_986_409#_c_672_p
+ N_A_986_409#_c_629_n N_A_986_409#_c_630_n N_A_986_409#_c_631_n
+ N_A_986_409#_c_632_n N_A_986_409#_c_633_n N_A_986_409#_c_634_n
+ N_A_986_409#_c_661_p N_A_986_409#_c_635_n N_A_986_409#_c_636_n
+ N_A_986_409#_c_637_n PM_SKY130_FD_SC_LP__SDFSTP_LP%A_986_409#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_1425_99# N_A_1425_99#_M1025_s
+ N_A_1425_99#_M1036_d N_A_1425_99#_M1034_g N_A_1425_99#_c_832_n
+ N_A_1425_99#_M1009_g N_A_1425_99#_c_833_n N_A_1425_99#_c_839_n
+ N_A_1425_99#_c_834_n N_A_1425_99#_c_840_n N_A_1425_99#_c_841_n
+ N_A_1425_99#_c_835_n N_A_1425_99#_c_836_n
+ PM_SKY130_FD_SC_LP__SDFSTP_LP%A_1425_99#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_1199_419# N_A_1199_419#_M1020_d
+ N_A_1199_419#_M1019_d N_A_1199_419#_M1036_g N_A_1199_419#_c_907_n
+ N_A_1199_419#_c_908_n N_A_1199_419#_M1025_g N_A_1199_419#_M1043_g
+ N_A_1199_419#_M1008_g N_A_1199_419#_c_911_n N_A_1199_419#_c_931_n
+ N_A_1199_419#_c_947_n N_A_1199_419#_c_932_n N_A_1199_419#_c_933_n
+ N_A_1199_419#_c_912_n N_A_1199_419#_c_913_n N_A_1199_419#_c_914_n
+ N_A_1199_419#_c_915_n N_A_1199_419#_c_916_n N_A_1199_419#_c_917_n
+ N_A_1199_419#_c_918_n N_A_1199_419#_c_919_n N_A_1199_419#_c_920_n
+ N_A_1199_419#_c_921_n N_A_1199_419#_c_922_n N_A_1199_419#_c_923_n
+ N_A_1199_419#_c_924_n N_A_1199_419#_c_1014_n N_A_1199_419#_c_925_n
+ N_A_1199_419#_c_926_n N_A_1199_419#_c_927_n
+ PM_SKY130_FD_SC_LP__SDFSTP_LP%A_1199_419#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%SET_B N_SET_B_M1010_g N_SET_B_M1014_g
+ N_SET_B_c_1094_n N_SET_B_M1038_g N_SET_B_c_1095_n N_SET_B_c_1096_n
+ N_SET_B_M1021_g N_SET_B_c_1102_n N_SET_B_c_1103_n N_SET_B_c_1117_n SET_B
+ N_SET_B_c_1097_n N_SET_B_c_1106_n N_SET_B_c_1098_n N_SET_B_c_1099_n
+ PM_SKY130_FD_SC_LP__SDFSTP_LP%SET_B
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_750_108# N_A_750_108#_M1041_s
+ N_A_750_108#_M1002_s N_A_750_108#_M1035_g N_A_750_108#_M1031_g
+ N_A_750_108#_c_1220_n N_A_750_108#_c_1221_n N_A_750_108#_M1030_g
+ N_A_750_108#_c_1223_n N_A_750_108#_M1020_g N_A_750_108#_c_1225_n
+ N_A_750_108#_c_1226_n N_A_750_108#_c_1227_n N_A_750_108#_c_1240_n
+ N_A_750_108#_c_1241_n N_A_750_108#_c_1242_n N_A_750_108#_M1028_g
+ N_A_750_108#_c_1243_n N_A_750_108#_M1011_g N_A_750_108#_c_1244_n
+ N_A_750_108#_c_1245_n N_A_750_108#_c_1228_n N_A_750_108#_M1039_g
+ N_A_750_108#_c_1230_n N_A_750_108#_c_1231_n N_A_750_108#_c_1232_n
+ N_A_750_108#_c_1233_n N_A_750_108#_c_1247_n N_A_750_108#_c_1234_n
+ N_A_750_108#_c_1249_n N_A_750_108#_c_1235_n N_A_750_108#_c_1236_n
+ N_A_750_108#_c_1237_n N_A_750_108#_c_1252_n
+ PM_SKY130_FD_SC_LP__SDFSTP_LP%A_750_108#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_2172_40# N_A_2172_40#_M1005_s
+ N_A_2172_40#_M1015_s N_A_2172_40#_M1040_g N_A_2172_40#_c_1428_n
+ N_A_2172_40#_c_1429_n N_A_2172_40#_M1033_g N_A_2172_40#_c_1430_n
+ N_A_2172_40#_c_1431_n N_A_2172_40#_c_1432_n N_A_2172_40#_c_1433_n
+ N_A_2172_40#_c_1434_n N_A_2172_40#_c_1435_n N_A_2172_40#_c_1436_n
+ PM_SKY130_FD_SC_LP__SDFSTP_LP%A_2172_40#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_2006_125# N_A_2006_125#_M1042_d
+ N_A_2006_125#_M1011_d N_A_2006_125#_M1021_d N_A_2006_125#_c_1510_n
+ N_A_2006_125#_M1005_g N_A_2006_125#_c_1511_n N_A_2006_125#_c_1512_n
+ N_A_2006_125#_c_1513_n N_A_2006_125#_M1007_g N_A_2006_125#_M1015_g
+ N_A_2006_125#_c_1514_n N_A_2006_125#_M1027_g N_A_2006_125#_c_1516_n
+ N_A_2006_125#_M1003_g N_A_2006_125#_M1012_g N_A_2006_125#_c_1519_n
+ N_A_2006_125#_c_1520_n N_A_2006_125#_c_1521_n N_A_2006_125#_c_1522_n
+ N_A_2006_125#_c_1523_n N_A_2006_125#_c_1541_n N_A_2006_125#_c_1524_n
+ N_A_2006_125#_c_1525_n N_A_2006_125#_c_1548_n N_A_2006_125#_c_1526_n
+ N_A_2006_125#_c_1565_n N_A_2006_125#_c_1533_n N_A_2006_125#_c_1534_n
+ N_A_2006_125#_c_1535_n N_A_2006_125#_c_1536_n N_A_2006_125#_c_1606_n
+ N_A_2006_125#_c_1527_n N_A_2006_125#_c_1537_n N_A_2006_125#_c_1538_n
+ N_A_2006_125#_c_1611_n N_A_2006_125#_c_1539_n
+ PM_SKY130_FD_SC_LP__SDFSTP_LP%A_2006_125#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_2767_57# N_A_2767_57#_M1027_s
+ N_A_2767_57#_M1003_s N_A_2767_57#_M1032_g N_A_2767_57#_M1037_g
+ N_A_2767_57#_M1026_g N_A_2767_57#_c_1693_n N_A_2767_57#_c_1694_n
+ N_A_2767_57#_c_1695_n N_A_2767_57#_c_1696_n N_A_2767_57#_c_1697_n
+ N_A_2767_57#_c_1698_n N_A_2767_57#_c_1699_n N_A_2767_57#_c_1700_n
+ N_A_2767_57#_c_1701_n PM_SKY130_FD_SC_LP__SDFSTP_LP%A_2767_57#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%VPWR N_VPWR_M1006_d N_VPWR_M1018_d
+ N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_M1010_d N_VPWR_M1033_d N_VPWR_M1015_d
+ N_VPWR_M1003_d N_VPWR_c_1766_n N_VPWR_c_1767_n N_VPWR_c_1768_n N_VPWR_c_1769_n
+ N_VPWR_c_1770_n N_VPWR_c_1771_n N_VPWR_c_1772_n N_VPWR_c_1773_n
+ N_VPWR_c_1774_n N_VPWR_c_1775_n N_VPWR_c_1776_n N_VPWR_c_1777_n VPWR
+ N_VPWR_c_1778_n N_VPWR_c_1779_n N_VPWR_c_1780_n N_VPWR_c_1781_n
+ N_VPWR_c_1782_n N_VPWR_c_1783_n N_VPWR_c_1765_n N_VPWR_c_1785_n
+ N_VPWR_c_1786_n N_VPWR_c_1787_n N_VPWR_c_1788_n N_VPWR_c_1789_n
+ N_VPWR_c_1790_n PM_SKY130_FD_SC_LP__SDFSTP_LP%VPWR
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_245_406# N_A_245_406#_M1016_s
+ N_A_245_406#_M1000_d N_A_245_406#_c_1931_n N_A_245_406#_c_1932_n
+ N_A_245_406#_c_1933_n N_A_245_406#_c_1940_n N_A_245_406#_c_1941_n
+ N_A_245_406#_c_1951_n N_A_245_406#_c_1934_n N_A_245_406#_c_1935_n
+ N_A_245_406#_c_1936_n PM_SKY130_FD_SC_LP__SDFSTP_LP%A_245_406#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%A_352_406# N_A_352_406#_M1023_d
+ N_A_352_406#_M1020_s N_A_352_406#_M1016_d N_A_352_406#_M1019_s
+ N_A_352_406#_c_2012_n N_A_352_406#_c_2006_n N_A_352_406#_c_2007_n
+ N_A_352_406#_c_1991_n N_A_352_406#_c_1992_n N_A_352_406#_c_1993_n
+ N_A_352_406#_c_1994_n N_A_352_406#_c_1995_n N_A_352_406#_c_1996_n
+ N_A_352_406#_c_1997_n N_A_352_406#_c_1998_n N_A_352_406#_c_2062_n
+ N_A_352_406#_c_1999_n N_A_352_406#_c_2000_n N_A_352_406#_c_2001_n
+ N_A_352_406#_c_2009_n N_A_352_406#_c_2002_n N_A_352_406#_c_2003_n
+ N_A_352_406#_c_2051_n N_A_352_406#_c_2004_n N_A_352_406#_c_2005_n
+ N_A_352_406#_c_2011_n PM_SKY130_FD_SC_LP__SDFSTP_LP%A_352_406#
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%Q N_Q_M1026_d N_Q_M1037_d N_Q_c_2181_n Q Q Q Q Q
+ N_Q_c_2185_n Q PM_SKY130_FD_SC_LP__SDFSTP_LP%Q
x_PM_SKY130_FD_SC_LP__SDFSTP_LP%VGND N_VGND_M1004_d N_VGND_M1024_d
+ N_VGND_M1029_d N_VGND_M1034_d N_VGND_M1014_d N_VGND_M1038_d N_VGND_M1007_d
+ N_VGND_M1012_d N_VGND_c_2203_n N_VGND_c_2204_n N_VGND_c_2205_n N_VGND_c_2206_n
+ N_VGND_c_2207_n N_VGND_c_2208_n N_VGND_c_2209_n N_VGND_c_2210_n
+ N_VGND_c_2211_n N_VGND_c_2212_n N_VGND_c_2213_n N_VGND_c_2214_n
+ N_VGND_c_2215_n N_VGND_c_2216_n VGND N_VGND_c_2217_n N_VGND_c_2218_n
+ N_VGND_c_2219_n N_VGND_c_2220_n N_VGND_c_2221_n N_VGND_c_2222_n
+ N_VGND_c_2223_n N_VGND_c_2224_n N_VGND_c_2225_n N_VGND_c_2226_n
+ N_VGND_c_2227_n N_VGND_c_2228_n PM_SKY130_FD_SC_LP__SDFSTP_LP%VGND
cc_1 VNB N_SCE_M1006_g 0.0427438f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_2 VNB N_SCE_M1017_g 0.0233828f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.445
cc_3 VNB N_SCE_M1004_g 0.0226883f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_4 VNB N_SCE_M1044_g 0.0335591f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.445
cc_5 VNB N_SCE_c_320_n 0.0236987f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.625
cc_6 VNB N_SCE_c_321_n 0.00205846f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.79
cc_7 VNB N_SCE_c_322_n 0.00582476f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.045
cc_8 VNB N_SCE_c_323_n 0.00600931f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.045
cc_9 VNB N_SCE_c_324_n 0.0121024f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.195
cc_10 VNB N_SCE_c_325_n 0.0159395f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_11 VNB N_SCE_c_326_n 0.0557461f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.02
cc_12 VNB N_SCE_c_327_n 0.0125325f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.045
cc_13 VNB N_SCE_c_328_n 0.0046114f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=1.045
cc_14 VNB N_A_27_409#_c_412_n 0.0363763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_409#_c_413_n 0.0164534f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.12
cc_16 VNB N_A_27_409#_c_414_n 0.0243003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_409#_c_415_n 0.00987081f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_18 VNB N_A_27_409#_c_416_n 0.0147561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_409#_c_417_n 0.034586f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.625
cc_20 VNB N_A_27_409#_c_418_n 0.00338121f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.195
cc_21 VNB N_A_27_409#_c_419_n 0.0212352f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_22 VNB N_A_27_409#_c_420_n 0.0088434f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.84
cc_23 VNB N_D_M1023_g 0.0491821f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.445
cc_24 VNB D 0.00314213f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_25 VNB N_D_c_483_n 0.0153543f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.445
cc_26 VNB N_SCD_c_522_n 0.0167014f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.185
cc_27 VNB N_SCD_c_523_n 0.0196493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB SCD 0.00511008f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.445
cc_29 VNB N_SCD_c_525_n 0.0629181f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=2.53
cc_30 VNB N_SCD_c_526_n 0.0175307f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_31 VNB N_CLK_M1041_g 0.0224242f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_32 VNB N_CLK_c_573_n 0.026721f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.445
cc_33 VNB N_CLK_M1029_g 0.0210687f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.12
cc_34 VNB N_CLK_c_575_n 0.0185747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB CLK 0.00236067f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_36 VNB N_CLK_c_577_n 0.00249638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_986_409#_M1045_g 0.0239136f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.12
cc_38 VNB N_A_986_409#_M1042_g 0.0244773f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_39 VNB N_A_986_409#_c_627_n 0.0126921f $X=-0.19 $Y=-0.245 $X2=2.672 $Y2=1.285
cc_40 VNB N_A_986_409#_c_628_n 0.032059f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_41 VNB N_A_986_409#_c_629_n 4.47893e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_986_409#_c_630_n 0.0134463f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.02
cc_43 VNB N_A_986_409#_c_631_n 0.0087483f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.045
cc_44 VNB N_A_986_409#_c_632_n 0.00644975f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.045
cc_45 VNB N_A_986_409#_c_633_n 0.0035526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_986_409#_c_634_n 0.0135028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_986_409#_c_635_n 0.0302581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_986_409#_c_636_n 0.00388401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_986_409#_c_637_n 0.00912808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1425_99#_M1034_g 0.0220336f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.855
cc_51 VNB N_A_1425_99#_c_832_n 0.0571353f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.445
cc_52 VNB N_A_1425_99#_c_833_n 0.00315975f $X=-0.19 $Y=-0.245 $X2=2.585
+ $Y2=0.445
cc_53 VNB N_A_1425_99#_c_834_n 0.0173161f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_54 VNB N_A_1425_99#_c_835_n 0.00695255f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.79
cc_55 VNB N_A_1425_99#_c_836_n 0.0126091f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.045
cc_56 VNB N_A_1199_419#_c_907_n 0.0194217f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.12
cc_57 VNB N_A_1199_419#_c_908_n 0.00919322f $X=-0.19 $Y=-0.245 $X2=2.585
+ $Y2=0.445
cc_58 VNB N_A_1199_419#_M1025_g 0.0206249f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_59 VNB N_A_1199_419#_M1008_g 0.0215614f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.02
cc_60 VNB N_A_1199_419#_c_911_n 0.0169652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1199_419#_c_912_n 0.00588726f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_62 VNB N_A_1199_419#_c_913_n 0.00513605f $X=-0.19 $Y=-0.245 $X2=2.075
+ $Y2=0.84
cc_63 VNB N_A_1199_419#_c_914_n 0.00714464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1199_419#_c_915_n 0.0124553f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.02
cc_65 VNB N_A_1199_419#_c_916_n 0.025629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1199_419#_c_917_n 0.00348498f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.02
cc_67 VNB N_A_1199_419#_c_918_n 0.00220516f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.02
cc_68 VNB N_A_1199_419#_c_919_n 0.0102835f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.045
cc_69 VNB N_A_1199_419#_c_920_n 0.00329787f $X=-0.19 $Y=-0.245 $X2=2.16
+ $Y2=1.045
cc_70 VNB N_A_1199_419#_c_921_n 0.00947584f $X=-0.19 $Y=-0.245 $X2=2.275
+ $Y2=1.045
cc_71 VNB N_A_1199_419#_c_922_n 0.00684256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1199_419#_c_923_n 0.00535137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1199_419#_c_924_n 0.00671756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1199_419#_c_925_n 0.00546133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1199_419#_c_926_n 0.0145769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1199_419#_c_927_n 0.0132055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_SET_B_M1014_g 0.0402952f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.445
cc_78 VNB N_SET_B_c_1094_n 0.0187067f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.855
cc_79 VNB N_SET_B_c_1095_n 0.0666229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_SET_B_c_1096_n 0.0064741f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.12
cc_81 VNB N_SET_B_c_1097_n 0.0573702f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.045
cc_82 VNB N_SET_B_c_1098_n 0.00148747f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_83 VNB N_SET_B_c_1099_n 0.0134554f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_84 VNB N_A_750_108#_M1031_g 0.0173002f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=1.12
cc_85 VNB N_A_750_108#_c_1220_n 0.0177294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_750_108#_c_1221_n 0.00711524f $X=-0.19 $Y=-0.245 $X2=2.655
+ $Y2=1.79
cc_87 VNB N_A_750_108#_M1030_g 0.0205832f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_88 VNB N_A_750_108#_c_1223_n 0.0499981f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.625
cc_89 VNB N_A_750_108#_M1020_g 0.0292054f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.02
cc_90 VNB N_A_750_108#_c_1225_n 0.0197077f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.045
cc_91 VNB N_A_750_108#_c_1226_n 0.313104f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.045
cc_92 VNB N_A_750_108#_c_1227_n 0.012806f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.195
cc_93 VNB N_A_750_108#_c_1228_n 0.0214876f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.02
cc_94 VNB N_A_750_108#_M1039_g 0.0239767f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.02
cc_95 VNB N_A_750_108#_c_1230_n 0.00458405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_750_108#_c_1231_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=1.68
+ $Y2=1.045
cc_97 VNB N_A_750_108#_c_1232_n 0.00611956f $X=-0.19 $Y=-0.245 $X2=1.565
+ $Y2=1.045
cc_98 VNB N_A_750_108#_c_1233_n 0.0137937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_750_108#_c_1234_n 0.0133243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_750_108#_c_1235_n 0.00127691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_750_108#_c_1236_n 0.016939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_750_108#_c_1237_n 0.00232128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2172_40#_M1040_g 0.0354732f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.855
cc_104 VNB N_A_2172_40#_c_1428_n 0.0202272f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.445
cc_105 VNB N_A_2172_40#_c_1429_n 0.00815301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2172_40#_c_1430_n 0.00235378f $X=-0.19 $Y=-0.245 $X2=2.655
+ $Y2=2.53
cc_107 VNB N_A_2172_40#_c_1431_n 0.00951594f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.12
cc_108 VNB N_A_2172_40#_c_1432_n 8.40012e-19 $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.625
cc_109 VNB N_A_2172_40#_c_1433_n 0.025401f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.02
cc_110 VNB N_A_2172_40#_c_1434_n 0.0166951f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.02
cc_111 VNB N_A_2172_40#_c_1435_n 0.0121871f $X=-0.19 $Y=-0.245 $X2=2.04
+ $Y2=1.045
cc_112 VNB N_A_2172_40#_c_1436_n 0.0492363f $X=-0.19 $Y=-0.245 $X2=2.672
+ $Y2=1.285
cc_113 VNB N_A_2006_125#_c_1510_n 0.020185f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.445
cc_114 VNB N_A_2006_125#_c_1511_n 0.0103315f $X=-0.19 $Y=-0.245 $X2=2.585
+ $Y2=1.12
cc_115 VNB N_A_2006_125#_c_1512_n 0.00898983f $X=-0.19 $Y=-0.245 $X2=2.585
+ $Y2=0.445
cc_116 VNB N_A_2006_125#_c_1513_n 0.0209802f $X=-0.19 $Y=-0.245 $X2=2.585
+ $Y2=0.445
cc_117 VNB N_A_2006_125#_c_1514_n 0.0223269f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.12
cc_118 VNB N_A_2006_125#_M1027_g 0.047819f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.02
cc_119 VNB N_A_2006_125#_c_1516_n 0.00622978f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.02
cc_120 VNB N_A_2006_125#_M1003_g 0.0056572f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.195
cc_121 VNB N_A_2006_125#_M1012_g 0.0437846f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_122 VNB N_A_2006_125#_c_1519_n 0.025162f $X=-0.19 $Y=-0.245 $X2=1.595
+ $Y2=0.84
cc_123 VNB N_A_2006_125#_c_1520_n 0.00952398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_2006_125#_c_1521_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2006_125#_c_1522_n 0.00847484f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_126 VNB N_A_2006_125#_c_1523_n 0.00697891f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.02
cc_127 VNB N_A_2006_125#_c_1524_n 0.0221473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_2006_125#_c_1525_n 0.0046914f $X=-0.19 $Y=-0.245 $X2=2.16
+ $Y2=1.045
cc_129 VNB N_A_2006_125#_c_1526_n 0.00519088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_2006_125#_c_1527_n 0.0431905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_2767_57#_M1032_g 0.0241349f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=0.855
cc_132 VNB N_A_2767_57#_M1026_g 0.0279877f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=1.79
cc_133 VNB N_A_2767_57#_c_1693_n 0.0245459f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.625
cc_134 VNB N_A_2767_57#_c_1694_n 0.0123324f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.02
cc_135 VNB N_A_2767_57#_c_1695_n 0.00531848f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.02
cc_136 VNB N_A_2767_57#_c_1696_n 0.00550225f $X=-0.19 $Y=-0.245 $X2=1.8
+ $Y2=1.045
cc_137 VNB N_A_2767_57#_c_1697_n 0.0109226f $X=-0.19 $Y=-0.245 $X2=2.672
+ $Y2=1.285
cc_138 VNB N_A_2767_57#_c_1698_n 0.0174539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_2767_57#_c_1699_n 0.0100926f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=1.02
cc_140 VNB N_A_2767_57#_c_1700_n 0.00142388f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.02
cc_141 VNB N_A_2767_57#_c_1701_n 0.0279586f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.02
cc_142 VNB N_VPWR_c_1765_n 0.661241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_352_406#_c_1991_n 0.010657f $X=-0.19 $Y=-0.245 $X2=2.655 $Y2=2.53
cc_144 VNB N_A_352_406#_c_1992_n 0.00535067f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.12
cc_145 VNB N_A_352_406#_c_1993_n 0.00924181f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.625
cc_146 VNB N_A_352_406#_c_1994_n 0.00784801f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.02
cc_147 VNB N_A_352_406#_c_1995_n 0.019365f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.02
cc_148 VNB N_A_352_406#_c_1996_n 0.00353386f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=1.02
cc_149 VNB N_A_352_406#_c_1997_n 0.00454056f $X=-0.19 $Y=-0.245 $X2=2.04
+ $Y2=1.045
cc_150 VNB N_A_352_406#_c_1998_n 0.0103953f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.045
cc_151 VNB N_A_352_406#_c_1999_n 0.00220255f $X=-0.19 $Y=-0.245 $X2=2.672
+ $Y2=1.28
cc_152 VNB N_A_352_406#_c_2000_n 0.020878f $X=-0.19 $Y=-0.245 $X2=2.672
+ $Y2=1.285
cc_153 VNB N_A_352_406#_c_2001_n 0.00267466f $X=-0.19 $Y=-0.245 $X2=2.675
+ $Y2=1.285
cc_154 VNB N_A_352_406#_c_2002_n 0.00703304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_A_352_406#_c_2003_n 0.0029333f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.02
cc_156 VNB N_A_352_406#_c_2004_n 0.00729677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_A_352_406#_c_2005_n 0.00712722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_Q_c_2181_n 0.0223955f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.855
cc_159 VNB Q 0.0478482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2203_n 0.00608103f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.02
cc_161 VNB N_VGND_c_2204_n 0.00240024f $X=-0.19 $Y=-0.245 $X2=1.8 $Y2=1.045
cc_162 VNB N_VGND_c_2205_n 0.0144133f $X=-0.19 $Y=-0.245 $X2=2.672 $Y2=1.285
cc_163 VNB N_VGND_c_2206_n 0.0119842f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=0.84
cc_164 VNB N_VGND_c_2207_n 0.015886f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=1.285
cc_165 VNB N_VGND_c_2208_n 0.0232945f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.02
cc_166 VNB N_VGND_c_2209_n 0.0102818f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.045
cc_167 VNB N_VGND_c_2210_n 0.00475893f $X=-0.19 $Y=-0.245 $X2=2.275 $Y2=1.045
cc_168 VNB N_VGND_c_2211_n 0.0336361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2212_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2213_n 0.0570966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2214_n 0.00585462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2215_n 0.0455168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2216_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2217_n 0.0302588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2218_n 0.0458216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2219_n 0.066685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2220_n 0.0355252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2221_n 0.0275301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2222_n 0.0271986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2223_n 0.816082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2224_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2225_n 0.00356907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2226_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2227_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2228_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VPB N_SCE_M1006_g 0.0557053f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_187 VPB N_SCE_M1018_g 0.0298127f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=2.53
cc_188 VPB N_SCE_c_321_n 0.0114869f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.79
cc_189 VPB N_SCE_c_332_n 6.99016e-19 $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_190 VPB N_A_27_409#_M1016_g 0.0398327f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.855
cc_191 VPB N_A_27_409#_c_414_n 0.024046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_27_409#_c_415_n 0.0049422f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=1.79
cc_193 VPB N_A_27_409#_c_424_n 0.0516919f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.02
cc_194 VPB N_A_27_409#_c_418_n 0.00631498f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.195
cc_195 VPB N_A_27_409#_c_420_n 0.00612236f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.84
cc_196 VPB N_D_M1001_g 0.0299465f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_197 VPB D 0.00288225f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.445
cc_198 VPB N_D_c_483_n 0.0093985f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=0.445
cc_199 VPB N_SCD_M1000_g 0.031816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB SCD 0.00521534f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=0.445
cc_201 VPB N_SCD_c_525_n 0.0287329f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=2.53
cc_202 VPB N_CLK_M1002_g 0.0319121f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.855
cc_203 VPB CLK 0.00275386f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=1.79
cc_204 VPB N_CLK_c_577_n 0.0193092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_986_409#_M1019_g 0.0364776f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.855
cc_206 VPB N_A_986_409#_M1013_g 0.026613f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_207 VPB N_A_986_409#_c_640_n 0.00722948f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.02
cc_208 VPB N_A_986_409#_c_641_n 0.010463f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.02
cc_209 VPB N_A_986_409#_c_642_n 0.00253984f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.02
cc_210 VPB N_A_986_409#_c_643_n 0.00248188f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.195
cc_211 VPB N_A_986_409#_c_629_n 0.00629199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_986_409#_c_630_n 5.13679e-19 $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.02
cc_213 VPB N_A_986_409#_c_632_n 0.00439862f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.045
cc_214 VPB N_A_986_409#_c_634_n 0.0145452f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_986_409#_c_637_n 0.0217237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_1425_99#_c_832_n 0.0364729f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.445
cc_217 VPB N_A_1425_99#_M1009_g 0.0312251f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=1.12
cc_218 VPB N_A_1425_99#_c_839_n 0.00332961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1425_99#_c_840_n 3.51419e-19 $X=-0.19 $Y=1.655 $X2=2.655 $Y2=2.53
cc_220 VPB N_A_1425_99#_c_841_n 0.0114339f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_221 VPB N_A_1199_419#_M1036_g 0.0316409f $X=-0.19 $Y=1.655 $X2=1.005
+ $Y2=0.855
cc_222 VPB N_A_1199_419#_M1043_g 0.0277925f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.285
cc_223 VPB N_A_1199_419#_c_911_n 0.00718046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_1199_419#_c_931_n 0.0145467f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=1.045
cc_225 VPB N_A_1199_419#_c_932_n 0.00614413f $X=-0.19 $Y=1.655 $X2=2.672
+ $Y2=1.285
cc_226 VPB N_A_1199_419#_c_933_n 0.00276195f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.285
cc_227 VPB N_A_1199_419#_c_913_n 0.00941752f $X=-0.19 $Y=1.655 $X2=2.075
+ $Y2=0.84
cc_228 VPB N_A_1199_419#_c_918_n 0.0039712f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.02
cc_229 VPB N_A_1199_419#_c_919_n 0.0160659f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.045
cc_230 VPB N_A_1199_419#_c_925_n 9.02542e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_SET_B_M1010_g 0.0270064f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_232 VPB N_SET_B_M1021_g 0.031323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_SET_B_c_1102_n 0.0161347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_SET_B_c_1103_n 0.0254179f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_235 VPB SET_B 9.33844e-19 $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.02
cc_236 VPB N_SET_B_c_1097_n 0.00926324f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=1.045
cc_237 VPB N_SET_B_c_1106_n 0.00224522f $X=-0.19 $Y=1.655 $X2=1.8 $Y2=1.045
cc_238 VPB N_SET_B_c_1098_n 0.00201299f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_239 VPB N_SET_B_c_1099_n 0.0323657f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_240 VPB N_A_750_108#_M1035_g 0.0296819f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.855
cc_241 VPB N_A_750_108#_c_1225_n 0.0128181f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=1.045
cc_242 VPB N_A_750_108#_c_1240_n 0.0262822f $X=-0.19 $Y=1.655 $X2=2.275
+ $Y2=1.195
cc_243 VPB N_A_750_108#_c_1241_n 0.0115398f $X=-0.19 $Y=1.655 $X2=2.672 $Y2=1.28
cc_244 VPB N_A_750_108#_c_1242_n 0.0220437f $X=-0.19 $Y=1.655 $X2=2.672
+ $Y2=1.285
cc_245 VPB N_A_750_108#_c_1243_n 0.0212961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_750_108#_c_1244_n 0.0283613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_750_108#_c_1245_n 0.00935016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_750_108#_c_1228_n 0.0123727f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.02
cc_249 VPB N_A_750_108#_c_1247_n 0.0101373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_750_108#_c_1234_n 0.00814918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_750_108#_c_1249_n 0.00346979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_750_108#_c_1235_n 0.00105063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_750_108#_c_1236_n 0.0268152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_750_108#_c_1252_n 0.00375396f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_2172_40#_M1033_g 0.0296154f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=0.445
cc_256 VPB N_A_2172_40#_c_1430_n 0.00313155f $X=-0.19 $Y=1.655 $X2=2.655
+ $Y2=2.53
cc_257 VPB N_A_2172_40#_c_1435_n 0.0150564f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=1.045
cc_258 VPB N_A_2172_40#_c_1436_n 0.029609f $X=-0.19 $Y=1.655 $X2=2.672 $Y2=1.285
cc_259 VPB N_A_2006_125#_M1015_g 0.0300241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_2006_125#_c_1514_n 0.0157925f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.12
cc_261 VPB N_A_2006_125#_M1003_g 0.0317764f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.195
cc_262 VPB N_A_2006_125#_c_1520_n 0.00471867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_2006_125#_c_1526_n 0.003589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_2006_125#_c_1533_n 0.00234021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_2006_125#_c_1534_n 0.00411508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_2006_125#_c_1535_n 0.024152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_2006_125#_c_1536_n 2.73935e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_2006_125#_c_1537_n 0.00440917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_2006_125#_c_1538_n 0.00293285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_2006_125#_c_1539_n 0.00463457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_2767_57#_M1037_g 0.0327251f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=1.12
cc_272 VPB N_A_2767_57#_c_1694_n 0.00261142f $X=-0.19 $Y=1.655 $X2=0.915
+ $Y2=1.02
cc_273 VPB N_A_2767_57#_c_1696_n 0.0172535f $X=-0.19 $Y=1.655 $X2=1.8 $Y2=1.045
cc_274 VPB N_A_2767_57#_c_1700_n 7.59613e-19 $X=-0.19 $Y=1.655 $X2=0.645
+ $Y2=1.02
cc_275 VPB N_VPWR_c_1766_n 0.0166114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1767_n 0.00216255f $X=-0.19 $Y=1.655 $X2=2.672 $Y2=1.285
cc_277 VPB N_VPWR_c_1768_n 0.00177638f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=0.84
cc_278 VPB N_VPWR_c_1769_n 0.00487982f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.285
cc_279 VPB N_VPWR_c_1770_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.02
cc_280 VPB N_VPWR_c_1771_n 0.00284591f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=1.045
cc_281 VPB N_VPWR_c_1772_n 0.0261478f $X=-0.19 $Y=1.655 $X2=2.275 $Y2=1.045
cc_282 VPB N_VPWR_c_1773_n 0.0202407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1774_n 0.0448104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1775_n 0.00516205f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1776_n 0.0216466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_1777_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_1778_n 0.0344024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_1779_n 0.0651706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_1780_n 0.0270015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_1781_n 0.069175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1782_n 0.0462043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_1783_n 0.0253236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_1765_n 0.122913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_1785_n 0.0243996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_1786_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_1787_n 0.00631504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_1788_n 0.00510188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_1789_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_1790_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_300 VPB N_A_245_406#_c_1931_n 0.010689f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=0.855
cc_301 VPB N_A_245_406#_c_1932_n 0.003222f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=1.12
cc_302 VPB N_A_245_406#_c_1933_n 0.00392134f $X=-0.19 $Y=1.655 $X2=2.585
+ $Y2=0.445
cc_303 VPB N_A_245_406#_c_1934_n 0.00455709f $X=-0.19 $Y=1.655 $X2=2.675
+ $Y2=1.285
cc_304 VPB N_A_245_406#_c_1935_n 0.00710892f $X=-0.19 $Y=1.655 $X2=1.565
+ $Y2=1.02
cc_305 VPB N_A_245_406#_c_1936_n 0.00152567f $X=-0.19 $Y=1.655 $X2=0.915
+ $Y2=1.02
cc_306 VPB N_A_352_406#_c_2006_n 0.0137929f $X=-0.19 $Y=1.655 $X2=2.655 $Y2=1.79
cc_307 VPB N_A_352_406#_c_2007_n 0.00245018f $X=-0.19 $Y=1.655 $X2=2.655
+ $Y2=2.53
cc_308 VPB N_A_352_406#_c_1992_n 0.0026312f $X=-0.19 $Y=1.655 $X2=2.675 $Y2=1.12
cc_309 VPB N_A_352_406#_c_2009_n 0.0059824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_310 VPB N_A_352_406#_c_2005_n 0.00741352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_311 VPB N_A_352_406#_c_2011_n 0.0173087f $X=-0.19 $Y=1.655 $X2=2.275
+ $Y2=1.045
cc_312 VPB Q 0.0107174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_313 VPB Q 0.0417159f $X=-0.19 $Y=1.655 $X2=2.585 $Y2=0.445
cc_314 VPB N_Q_c_2185_n 0.0224082f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_315 N_SCE_c_323_n N_A_27_409#_c_412_n 0.0199245f $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_316 N_SCE_c_326_n N_A_27_409#_c_412_n 0.00444069f $X=1.005 $Y=1.02 $X2=0
+ $Y2=0
cc_317 N_SCE_M1004_g N_A_27_409#_c_413_n 0.00639606f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_318 N_SCE_M1006_g N_A_27_409#_c_414_n 0.00979362f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_319 N_SCE_c_326_n N_A_27_409#_c_414_n 0.00116338f $X=1.005 $Y=1.02 $X2=0
+ $Y2=0
cc_320 N_SCE_c_327_n N_A_27_409#_c_414_n 0.013257f $X=1.565 $Y=1.045 $X2=0 $Y2=0
cc_321 N_SCE_c_323_n N_A_27_409#_c_415_n 0.0012047f $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_322 N_SCE_M1004_g N_A_27_409#_c_416_n 0.00444069f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_323 N_SCE_c_322_n N_A_27_409#_c_416_n 0.00282681f $X=2.04 $Y=1.045 $X2=0
+ $Y2=0
cc_324 N_SCE_c_323_n N_A_27_409#_c_416_n 0.00764278f $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_325 N_SCE_M1006_g N_A_27_409#_c_417_n 0.0177015f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_326 N_SCE_M1017_g N_A_27_409#_c_417_n 0.00697224f $X=0.645 $Y=0.445 $X2=0
+ $Y2=0
cc_327 N_SCE_c_326_n N_A_27_409#_c_417_n 0.0143008f $X=1.005 $Y=1.02 $X2=0 $Y2=0
cc_328 N_SCE_c_327_n N_A_27_409#_c_417_n 0.0163704f $X=1.565 $Y=1.045 $X2=0
+ $Y2=0
cc_329 N_SCE_M1006_g N_A_27_409#_c_424_n 0.0343357f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_330 N_SCE_M1006_g N_A_27_409#_c_418_n 0.0322447f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_331 N_SCE_c_326_n N_A_27_409#_c_418_n 0.0107525f $X=1.005 $Y=1.02 $X2=0 $Y2=0
cc_332 N_SCE_c_327_n N_A_27_409#_c_418_n 0.035032f $X=1.565 $Y=1.045 $X2=0 $Y2=0
cc_333 N_SCE_M1017_g N_A_27_409#_c_419_n 0.00856247f $X=0.645 $Y=0.445 $X2=0
+ $Y2=0
cc_334 N_SCE_M1004_g N_A_27_409#_c_419_n 0.00111271f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_335 N_SCE_c_326_n N_A_27_409#_c_419_n 0.0056226f $X=1.005 $Y=1.02 $X2=0 $Y2=0
cc_336 N_SCE_M1006_g N_A_27_409#_c_420_n 0.00744399f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_337 N_SCE_M1018_g N_D_M1001_g 0.0756772f $X=2.655 $Y=2.53 $X2=0 $Y2=0
cc_338 N_SCE_M1044_g N_D_M1023_g 0.0432552f $X=2.585 $Y=0.445 $X2=0 $Y2=0
cc_339 N_SCE_c_332_n N_D_M1023_g 0.00111852f $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_340 N_SCE_c_328_n N_D_M1023_g 0.0216649f $X=2.275 $Y=1.045 $X2=0 $Y2=0
cc_341 N_SCE_c_320_n D 0.00113718f $X=2.675 $Y=1.625 $X2=0 $Y2=0
cc_342 N_SCE_c_323_n D 0.0566405f $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_343 N_SCE_c_332_n D 0.0220339f $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_344 N_SCE_c_320_n N_D_c_483_n 0.0207503f $X=2.675 $Y=1.625 $X2=0 $Y2=0
cc_345 N_SCE_c_322_n N_D_c_483_n 0.00266912f $X=2.04 $Y=1.045 $X2=0 $Y2=0
cc_346 N_SCE_c_332_n N_D_c_483_n 4.1374e-19 $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_347 N_SCE_c_328_n N_D_c_483_n 0.00181781f $X=2.275 $Y=1.045 $X2=0 $Y2=0
cc_348 N_SCE_M1044_g N_SCD_c_522_n 0.0404789f $X=2.585 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_349 N_SCE_M1018_g N_SCD_c_525_n 0.046459f $X=2.655 $Y=2.53 $X2=0 $Y2=0
cc_350 N_SCE_c_320_n N_SCD_c_525_n 0.0197677f $X=2.675 $Y=1.625 $X2=0 $Y2=0
cc_351 N_SCE_c_332_n N_SCD_c_525_n 5.76655e-19 $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_352 N_SCE_M1044_g N_SCD_c_526_n 0.00628173f $X=2.585 $Y=0.445 $X2=0 $Y2=0
cc_353 N_SCE_c_324_n N_SCD_c_526_n 2.19935e-19 $X=2.51 $Y=1.195 $X2=0 $Y2=0
cc_354 N_SCE_c_325_n N_SCD_c_526_n 0.0197677f $X=2.675 $Y=1.285 $X2=0 $Y2=0
cc_355 N_SCE_M1006_g N_VPWR_c_1766_n 0.025033f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_356 N_SCE_M1018_g N_VPWR_c_1767_n 0.0108277f $X=2.655 $Y=2.53 $X2=0 $Y2=0
cc_357 N_SCE_M1018_g N_VPWR_c_1774_n 0.00781473f $X=2.655 $Y=2.53 $X2=0 $Y2=0
cc_358 N_SCE_M1006_g N_VPWR_c_1765_n 0.014085f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_359 N_SCE_M1018_g N_VPWR_c_1765_n 0.00750628f $X=2.655 $Y=2.53 $X2=0 $Y2=0
cc_360 N_SCE_M1006_g N_VPWR_c_1785_n 0.00769046f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_361 N_SCE_M1006_g N_A_245_406#_c_1931_n 0.00195302f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_362 N_SCE_M1018_g N_A_245_406#_c_1932_n 0.00169926f $X=2.655 $Y=2.53 $X2=0
+ $Y2=0
cc_363 N_SCE_M1006_g N_A_245_406#_c_1933_n 3.95513e-19 $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_364 N_SCE_M1018_g N_A_245_406#_c_1940_n 0.00579089f $X=2.655 $Y=2.53 $X2=0
+ $Y2=0
cc_365 N_SCE_M1018_g N_A_245_406#_c_1941_n 0.0167879f $X=2.655 $Y=2.53 $X2=0
+ $Y2=0
cc_366 N_SCE_M1018_g N_A_352_406#_c_2012_n 9.35961e-19 $X=2.655 $Y=2.53 $X2=0
+ $Y2=0
cc_367 N_SCE_M1018_g N_A_352_406#_c_2006_n 0.0146929f $X=2.655 $Y=2.53 $X2=0
+ $Y2=0
cc_368 N_SCE_c_321_n N_A_352_406#_c_2006_n 7.46077e-19 $X=2.675 $Y=1.79 $X2=0
+ $Y2=0
cc_369 N_SCE_c_332_n N_A_352_406#_c_2006_n 0.0237712f $X=2.675 $Y=1.285 $X2=0
+ $Y2=0
cc_370 N_SCE_M1044_g N_A_352_406#_c_1991_n 0.00386743f $X=2.585 $Y=0.445 $X2=0
+ $Y2=0
cc_371 N_SCE_c_324_n N_A_352_406#_c_1991_n 0.0167042f $X=2.51 $Y=1.195 $X2=0
+ $Y2=0
cc_372 N_SCE_c_325_n N_A_352_406#_c_1991_n 0.00137074f $X=2.675 $Y=1.285 $X2=0
+ $Y2=0
cc_373 N_SCE_M1044_g N_A_352_406#_c_1992_n 0.00315661f $X=2.585 $Y=0.445 $X2=0
+ $Y2=0
cc_374 N_SCE_M1018_g N_A_352_406#_c_1992_n 0.00348712f $X=2.655 $Y=2.53 $X2=0
+ $Y2=0
cc_375 N_SCE_c_324_n N_A_352_406#_c_1992_n 0.0130532f $X=2.51 $Y=1.195 $X2=0
+ $Y2=0
cc_376 N_SCE_c_332_n N_A_352_406#_c_1992_n 0.0365638f $X=2.675 $Y=1.285 $X2=0
+ $Y2=0
cc_377 N_SCE_c_325_n N_A_352_406#_c_1992_n 0.00365786f $X=2.675 $Y=1.285 $X2=0
+ $Y2=0
cc_378 N_SCE_M1044_g N_A_352_406#_c_2003_n 0.0168833f $X=2.585 $Y=0.445 $X2=0
+ $Y2=0
cc_379 N_SCE_c_324_n N_A_352_406#_c_2003_n 0.0201314f $X=2.51 $Y=1.195 $X2=0
+ $Y2=0
cc_380 N_SCE_c_328_n N_A_352_406#_c_2003_n 0.0142643f $X=2.275 $Y=1.045 $X2=0
+ $Y2=0
cc_381 N_SCE_M1017_g N_VGND_c_2203_n 0.00239794f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_382 N_SCE_M1004_g N_VGND_c_2203_n 0.0135711f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_383 N_SCE_c_327_n N_VGND_c_2203_n 0.0269388f $X=1.565 $Y=1.045 $X2=0 $Y2=0
cc_384 N_SCE_M1044_g N_VGND_c_2204_n 0.00206514f $X=2.585 $Y=0.445 $X2=0 $Y2=0
cc_385 N_SCE_M1017_g N_VGND_c_2217_n 0.00549284f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_386 N_SCE_M1004_g N_VGND_c_2217_n 0.00486043f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_387 N_SCE_M1044_g N_VGND_c_2218_n 0.00379072f $X=2.585 $Y=0.445 $X2=0 $Y2=0
cc_388 N_SCE_M1017_g N_VGND_c_2223_n 0.0110208f $X=0.645 $Y=0.445 $X2=0 $Y2=0
cc_389 N_SCE_M1004_g N_VGND_c_2223_n 0.00443987f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_390 N_SCE_M1044_g N_VGND_c_2223_n 0.00558182f $X=2.585 $Y=0.445 $X2=0 $Y2=0
cc_391 N_SCE_c_323_n N_VGND_c_2223_n 0.0226439f $X=1.8 $Y=1.045 $X2=0 $Y2=0
cc_392 N_SCE_c_326_n N_VGND_c_2223_n 6.74651e-19 $X=1.005 $Y=1.02 $X2=0 $Y2=0
cc_393 N_SCE_c_327_n N_VGND_c_2223_n 0.0171553f $X=1.565 $Y=1.045 $X2=0 $Y2=0
cc_394 N_A_27_409#_M1016_g N_D_M1001_g 0.0320039f $X=1.635 $Y=2.53 $X2=0 $Y2=0
cc_395 N_A_27_409#_c_412_n N_D_M1023_g 0.0231976f $X=1.685 $Y=1.46 $X2=0 $Y2=0
cc_396 N_A_27_409#_c_413_n N_D_M1023_g 0.0420076f $X=1.765 $Y=0.73 $X2=0 $Y2=0
cc_397 N_A_27_409#_c_415_n D 0.0247986f $X=1.635 $Y=1.625 $X2=0 $Y2=0
cc_398 N_A_27_409#_c_416_n D 2.72519e-19 $X=1.765 $Y=0.805 $X2=0 $Y2=0
cc_399 N_A_27_409#_c_418_n D 0.0265069f $X=1.22 $Y=1.625 $X2=0 $Y2=0
cc_400 N_A_27_409#_c_415_n N_D_c_483_n 0.0215238f $X=1.635 $Y=1.625 $X2=0 $Y2=0
cc_401 N_A_27_409#_M1016_g N_VPWR_c_1766_n 0.00357456f $X=1.635 $Y=2.53 $X2=0
+ $Y2=0
cc_402 N_A_27_409#_c_424_n N_VPWR_c_1766_n 0.0685263f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_403 N_A_27_409#_c_418_n N_VPWR_c_1766_n 0.0229033f $X=1.22 $Y=1.625 $X2=0
+ $Y2=0
cc_404 N_A_27_409#_M1016_g N_VPWR_c_1774_n 0.00531075f $X=1.635 $Y=2.53 $X2=0
+ $Y2=0
cc_405 N_A_27_409#_M1016_g N_VPWR_c_1765_n 0.0080075f $X=1.635 $Y=2.53 $X2=0
+ $Y2=0
cc_406 N_A_27_409#_c_424_n N_VPWR_c_1765_n 0.0125808f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_407 N_A_27_409#_c_424_n N_VPWR_c_1785_n 0.0220321f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_408 N_A_27_409#_M1016_g N_A_245_406#_c_1931_n 0.0169147f $X=1.635 $Y=2.53
+ $X2=0 $Y2=0
cc_409 N_A_27_409#_c_414_n N_A_245_406#_c_1931_n 0.00930681f $X=1.51 $Y=1.625
+ $X2=0 $Y2=0
cc_410 N_A_27_409#_c_418_n N_A_245_406#_c_1931_n 0.0124468f $X=1.22 $Y=1.625
+ $X2=0 $Y2=0
cc_411 N_A_27_409#_M1016_g N_A_245_406#_c_1932_n 0.016384f $X=1.635 $Y=2.53
+ $X2=0 $Y2=0
cc_412 N_A_27_409#_M1016_g N_A_245_406#_c_1933_n 0.00126082f $X=1.635 $Y=2.53
+ $X2=0 $Y2=0
cc_413 N_A_27_409#_M1016_g N_A_245_406#_c_1940_n 7.43022e-19 $X=1.635 $Y=2.53
+ $X2=0 $Y2=0
cc_414 N_A_27_409#_M1016_g N_A_352_406#_c_2012_n 0.0103858f $X=1.635 $Y=2.53
+ $X2=0 $Y2=0
cc_415 N_A_27_409#_M1016_g N_A_352_406#_c_2007_n 0.00535365f $X=1.635 $Y=2.53
+ $X2=0 $Y2=0
cc_416 N_A_27_409#_c_413_n N_A_352_406#_c_2003_n 0.00180619f $X=1.765 $Y=0.73
+ $X2=0 $Y2=0
cc_417 N_A_27_409#_c_413_n N_VGND_c_2203_n 0.0118404f $X=1.765 $Y=0.73 $X2=0
+ $Y2=0
cc_418 N_A_27_409#_c_419_n N_VGND_c_2203_n 0.0141221f $X=0.43 $Y=0.47 $X2=0
+ $Y2=0
cc_419 N_A_27_409#_c_419_n N_VGND_c_2217_n 0.0296879f $X=0.43 $Y=0.47 $X2=0
+ $Y2=0
cc_420 N_A_27_409#_c_413_n N_VGND_c_2218_n 0.00585385f $X=1.765 $Y=0.73 $X2=0
+ $Y2=0
cc_421 N_A_27_409#_c_416_n N_VGND_c_2218_n 0.0016562f $X=1.765 $Y=0.805 $X2=0
+ $Y2=0
cc_422 N_A_27_409#_M1017_s N_VGND_c_2223_n 0.00232985f $X=0.285 $Y=0.235 $X2=0
+ $Y2=0
cc_423 N_A_27_409#_c_413_n N_VGND_c_2223_n 0.00705373f $X=1.765 $Y=0.73 $X2=0
+ $Y2=0
cc_424 N_A_27_409#_c_416_n N_VGND_c_2223_n 0.00218182f $X=1.765 $Y=0.805 $X2=0
+ $Y2=0
cc_425 N_A_27_409#_c_419_n N_VGND_c_2223_n 0.0183089f $X=0.43 $Y=0.47 $X2=0
+ $Y2=0
cc_426 N_D_M1001_g N_VPWR_c_1767_n 9.0827e-19 $X=2.165 $Y=2.53 $X2=0 $Y2=0
cc_427 N_D_M1001_g N_VPWR_c_1774_n 0.00531052f $X=2.165 $Y=2.53 $X2=0 $Y2=0
cc_428 N_D_M1001_g N_VPWR_c_1765_n 0.00720256f $X=2.165 $Y=2.53 $X2=0 $Y2=0
cc_429 N_D_M1001_g N_A_245_406#_c_1931_n 8.97374e-19 $X=2.165 $Y=2.53 $X2=0
+ $Y2=0
cc_430 N_D_M1001_g N_A_245_406#_c_1932_n 0.0170768f $X=2.165 $Y=2.53 $X2=0 $Y2=0
cc_431 N_D_M1001_g N_A_245_406#_c_1940_n 0.00993317f $X=2.165 $Y=2.53 $X2=0
+ $Y2=0
cc_432 N_D_M1001_g N_A_245_406#_c_1951_n 0.00554657f $X=2.165 $Y=2.53 $X2=0
+ $Y2=0
cc_433 N_D_M1001_g N_A_352_406#_c_2012_n 0.0100996f $X=2.165 $Y=2.53 $X2=0 $Y2=0
cc_434 N_D_M1001_g N_A_352_406#_c_2006_n 0.0169748f $X=2.165 $Y=2.53 $X2=0 $Y2=0
cc_435 D N_A_352_406#_c_2006_n 0.0160355f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_436 N_D_c_483_n N_A_352_406#_c_2006_n 2.22766e-19 $X=2.135 $Y=1.625 $X2=0
+ $Y2=0
cc_437 N_D_M1001_g N_A_352_406#_c_2007_n 0.00145704f $X=2.165 $Y=2.53 $X2=0
+ $Y2=0
cc_438 D N_A_352_406#_c_2007_n 0.027305f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_439 N_D_c_483_n N_A_352_406#_c_2007_n 0.00162266f $X=2.135 $Y=1.625 $X2=0
+ $Y2=0
cc_440 N_D_M1023_g N_A_352_406#_c_2003_n 0.0110385f $X=2.155 $Y=0.445 $X2=0
+ $Y2=0
cc_441 N_D_M1023_g N_VGND_c_2218_n 0.0054778f $X=2.155 $Y=0.445 $X2=0 $Y2=0
cc_442 N_D_M1023_g N_VGND_c_2223_n 0.00623217f $X=2.155 $Y=0.445 $X2=0 $Y2=0
cc_443 N_SCD_c_525_n N_CLK_M1041_g 0.0212414f $X=3.525 $Y=1.325 $X2=0 $Y2=0
cc_444 N_SCD_M1000_g N_A_750_108#_c_1247_n 0.00137517f $X=3.185 $Y=2.53 $X2=0
+ $Y2=0
cc_445 N_SCD_M1000_g N_A_750_108#_c_1234_n 0.0043777f $X=3.185 $Y=2.53 $X2=0
+ $Y2=0
cc_446 SCD N_A_750_108#_c_1234_n 0.048119f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_447 N_SCD_c_525_n N_A_750_108#_c_1234_n 0.00523056f $X=3.525 $Y=1.325 $X2=0
+ $Y2=0
cc_448 N_SCD_c_526_n N_A_750_108#_c_1234_n 0.00371494f $X=3.375 $Y=1.16 $X2=0
+ $Y2=0
cc_449 N_SCD_c_523_n N_A_750_108#_c_1237_n 5.73316e-19 $X=3.135 $Y=0.805 $X2=0
+ $Y2=0
cc_450 N_SCD_c_526_n N_A_750_108#_c_1237_n 7.30551e-19 $X=3.375 $Y=1.16 $X2=0
+ $Y2=0
cc_451 N_SCD_M1000_g N_VPWR_c_1767_n 0.0116112f $X=3.185 $Y=2.53 $X2=0 $Y2=0
cc_452 N_SCD_M1000_g N_VPWR_c_1778_n 0.00781473f $X=3.185 $Y=2.53 $X2=0 $Y2=0
cc_453 N_SCD_M1000_g N_VPWR_c_1765_n 0.00831119f $X=3.185 $Y=2.53 $X2=0 $Y2=0
cc_454 N_SCD_M1000_g N_A_245_406#_c_1941_n 0.0187281f $X=3.185 $Y=2.53 $X2=0
+ $Y2=0
cc_455 N_SCD_M1000_g N_A_245_406#_c_1934_n 4.90931e-19 $X=3.185 $Y=2.53 $X2=0
+ $Y2=0
cc_456 SCD N_A_245_406#_c_1934_n 0.0211474f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_457 N_SCD_c_525_n N_A_245_406#_c_1934_n 0.00192767f $X=3.525 $Y=1.325 $X2=0
+ $Y2=0
cc_458 N_SCD_M1000_g N_A_245_406#_c_1935_n 5.20695e-19 $X=3.185 $Y=2.53 $X2=0
+ $Y2=0
cc_459 N_SCD_M1000_g N_A_352_406#_c_2006_n 0.00877477f $X=3.185 $Y=2.53 $X2=0
+ $Y2=0
cc_460 N_SCD_c_523_n N_A_352_406#_c_1991_n 0.00719882f $X=3.135 $Y=0.805 $X2=0
+ $Y2=0
cc_461 N_SCD_M1000_g N_A_352_406#_c_1992_n 0.0074731f $X=3.185 $Y=2.53 $X2=0
+ $Y2=0
cc_462 SCD N_A_352_406#_c_1992_n 0.0455899f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_463 N_SCD_c_525_n N_A_352_406#_c_1992_n 0.0192636f $X=3.525 $Y=1.325 $X2=0
+ $Y2=0
cc_464 N_SCD_c_526_n N_A_352_406#_c_1992_n 0.0114716f $X=3.375 $Y=1.16 $X2=0
+ $Y2=0
cc_465 N_SCD_c_523_n N_A_352_406#_c_1993_n 0.00299032f $X=3.135 $Y=0.805 $X2=0
+ $Y2=0
cc_466 SCD N_A_352_406#_c_1993_n 0.0176552f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_467 N_SCD_c_525_n N_A_352_406#_c_1993_n 0.00790305f $X=3.525 $Y=1.325 $X2=0
+ $Y2=0
cc_468 N_SCD_c_526_n N_A_352_406#_c_1993_n 0.00220996f $X=3.375 $Y=1.16 $X2=0
+ $Y2=0
cc_469 N_SCD_c_522_n N_A_352_406#_c_1994_n 0.0038599f $X=2.975 $Y=0.73 $X2=0
+ $Y2=0
cc_470 N_SCD_c_523_n N_A_352_406#_c_1994_n 0.00101587f $X=3.135 $Y=0.805 $X2=0
+ $Y2=0
cc_471 N_SCD_c_522_n N_A_352_406#_c_2003_n 0.00212691f $X=2.975 $Y=0.73 $X2=0
+ $Y2=0
cc_472 N_SCD_c_523_n N_A_352_406#_c_2051_n 0.00445598f $X=3.135 $Y=0.805 $X2=0
+ $Y2=0
cc_473 N_SCD_c_526_n N_A_352_406#_c_2051_n 0.0013265f $X=3.375 $Y=1.16 $X2=0
+ $Y2=0
cc_474 N_SCD_c_522_n N_VGND_c_2204_n 0.0112713f $X=2.975 $Y=0.73 $X2=0 $Y2=0
cc_475 N_SCD_c_523_n N_VGND_c_2204_n 0.00421813f $X=3.135 $Y=0.805 $X2=0 $Y2=0
cc_476 N_SCD_c_522_n N_VGND_c_2218_n 0.00367946f $X=2.975 $Y=0.73 $X2=0 $Y2=0
cc_477 N_SCD_c_522_n N_VGND_c_2223_n 0.00436992f $X=2.975 $Y=0.73 $X2=0 $Y2=0
cc_478 N_CLK_M1029_g N_A_750_108#_M1031_g 0.0104419f $X=4.5 $Y=0.75 $X2=0 $Y2=0
cc_479 N_CLK_c_573_n N_A_750_108#_c_1220_n 0.00908215f $X=4.252 $Y=1.623 $X2=0
+ $Y2=0
cc_480 CLK N_A_750_108#_c_1220_n 5.22851e-19 $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_481 N_CLK_c_575_n N_A_750_108#_c_1230_n 0.0104419f $X=4.305 $Y=1.315 $X2=0
+ $Y2=0
cc_482 N_CLK_M1002_g N_A_750_108#_c_1247_n 0.0157596f $X=4.275 $Y=2.545 $X2=0
+ $Y2=0
cc_483 N_CLK_M1041_g N_A_750_108#_c_1234_n 0.0149469f $X=4.11 $Y=0.75 $X2=0
+ $Y2=0
cc_484 N_CLK_M1002_g N_A_750_108#_c_1234_n 0.00690216f $X=4.275 $Y=2.545 $X2=0
+ $Y2=0
cc_485 CLK N_A_750_108#_c_1234_n 0.0241661f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_486 N_CLK_M1002_g N_A_750_108#_c_1249_n 0.0190356f $X=4.275 $Y=2.545 $X2=0
+ $Y2=0
cc_487 CLK N_A_750_108#_c_1249_n 0.0309857f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_488 N_CLK_c_577_n N_A_750_108#_c_1249_n 0.00183219f $X=4.305 $Y=1.675 $X2=0
+ $Y2=0
cc_489 N_CLK_c_573_n N_A_750_108#_c_1235_n 2.07603e-19 $X=4.252 $Y=1.623 $X2=0
+ $Y2=0
cc_490 N_CLK_M1002_g N_A_750_108#_c_1235_n 8.86822e-19 $X=4.275 $Y=2.545 $X2=0
+ $Y2=0
cc_491 CLK N_A_750_108#_c_1235_n 0.021809f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_492 N_CLK_c_573_n N_A_750_108#_c_1236_n 0.0179676f $X=4.252 $Y=1.623 $X2=0
+ $Y2=0
cc_493 N_CLK_M1002_g N_A_750_108#_c_1236_n 0.0294821f $X=4.275 $Y=2.545 $X2=0
+ $Y2=0
cc_494 CLK N_A_750_108#_c_1236_n 0.00230926f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_495 N_CLK_M1041_g N_A_750_108#_c_1237_n 0.00559423f $X=4.11 $Y=0.75 $X2=0
+ $Y2=0
cc_496 N_CLK_M1002_g N_A_750_108#_c_1252_n 0.00216931f $X=4.275 $Y=2.545 $X2=0
+ $Y2=0
cc_497 N_CLK_c_577_n N_A_750_108#_c_1252_n 0.00550457f $X=4.305 $Y=1.675 $X2=0
+ $Y2=0
cc_498 N_CLK_M1002_g N_VPWR_c_1768_n 0.0174514f $X=4.275 $Y=2.545 $X2=0 $Y2=0
cc_499 N_CLK_M1002_g N_VPWR_c_1778_n 0.00769046f $X=4.275 $Y=2.545 $X2=0 $Y2=0
cc_500 N_CLK_M1002_g N_VPWR_c_1765_n 0.0143431f $X=4.275 $Y=2.545 $X2=0 $Y2=0
cc_501 N_CLK_M1002_g N_A_245_406#_c_1934_n 5.39842e-19 $X=4.275 $Y=2.545 $X2=0
+ $Y2=0
cc_502 N_CLK_M1002_g N_A_245_406#_c_1935_n 9.21169e-19 $X=4.275 $Y=2.545 $X2=0
+ $Y2=0
cc_503 N_CLK_M1041_g N_A_352_406#_c_1994_n 0.00294561f $X=4.11 $Y=0.75 $X2=0
+ $Y2=0
cc_504 N_CLK_M1041_g N_A_352_406#_c_1995_n 0.00958377f $X=4.11 $Y=0.75 $X2=0
+ $Y2=0
cc_505 N_CLK_M1029_g N_A_352_406#_c_1995_n 2.32904e-19 $X=4.5 $Y=0.75 $X2=0
+ $Y2=0
cc_506 N_CLK_M1041_g N_A_352_406#_c_1997_n 0.00415822f $X=4.11 $Y=0.75 $X2=0
+ $Y2=0
cc_507 N_CLK_M1029_g N_A_352_406#_c_1997_n 0.00489413f $X=4.5 $Y=0.75 $X2=0
+ $Y2=0
cc_508 N_CLK_c_573_n N_A_352_406#_c_1998_n 0.00110106f $X=4.252 $Y=1.623 $X2=0
+ $Y2=0
cc_509 N_CLK_M1029_g N_A_352_406#_c_1998_n 0.0066768f $X=4.5 $Y=0.75 $X2=0 $Y2=0
cc_510 N_CLK_c_575_n N_A_352_406#_c_1998_n 0.00558211f $X=4.305 $Y=1.315 $X2=0
+ $Y2=0
cc_511 CLK N_A_352_406#_c_1998_n 0.0173858f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_512 N_CLK_c_573_n N_A_352_406#_c_2062_n 0.00291278f $X=4.252 $Y=1.623 $X2=0
+ $Y2=0
cc_513 N_CLK_c_575_n N_A_352_406#_c_2062_n 0.00551859f $X=4.305 $Y=1.315 $X2=0
+ $Y2=0
cc_514 CLK N_A_352_406#_c_2062_n 0.0129587f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_515 N_CLK_M1029_g N_A_352_406#_c_1999_n 7.00847e-19 $X=4.5 $Y=0.75 $X2=0
+ $Y2=0
cc_516 CLK N_A_352_406#_c_2005_n 0.0014091f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_517 N_CLK_M1029_g N_VGND_c_2205_n 0.00127668f $X=4.5 $Y=0.75 $X2=0 $Y2=0
cc_518 N_CLK_M1041_g N_VGND_c_2211_n 6.5362e-19 $X=4.11 $Y=0.75 $X2=0 $Y2=0
cc_519 N_CLK_M1029_g N_VGND_c_2211_n 0.00463045f $X=4.5 $Y=0.75 $X2=0 $Y2=0
cc_520 N_CLK_M1029_g N_VGND_c_2223_n 0.00493565f $X=4.5 $Y=0.75 $X2=0 $Y2=0
cc_521 N_A_986_409#_c_649_p N_A_1425_99#_M1036_d 0.0047688f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_522 N_A_986_409#_M1045_g N_A_1425_99#_M1034_g 0.0266791f $X=6.84 $Y=0.835
+ $X2=0 $Y2=0
cc_523 N_A_986_409#_c_627_n N_A_1425_99#_c_832_n 3.5911e-19 $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_524 N_A_986_409#_c_628_n N_A_1425_99#_c_832_n 0.0416558f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_525 N_A_986_409#_c_649_p N_A_1425_99#_c_832_n 9.21303e-19 $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_526 N_A_986_409#_c_654_p N_A_1425_99#_M1009_g 0.00194618f $X=6.81 $Y=2.98
+ $X2=0 $Y2=0
cc_527 N_A_986_409#_c_655_p N_A_1425_99#_M1009_g 0.00421674f $X=6.895 $Y=2.895
+ $X2=0 $Y2=0
cc_528 N_A_986_409#_c_649_p N_A_1425_99#_M1009_g 0.0232454f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_529 N_A_986_409#_c_649_p N_A_1425_99#_c_840_n 0.0243994f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_530 N_A_986_409#_c_649_p N_A_1425_99#_c_841_n 0.0461265f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_531 N_A_986_409#_c_643_n N_A_1199_419#_M1019_d 0.0086935f $X=6.035 $Y=2.895
+ $X2=0 $Y2=0
cc_532 N_A_986_409#_c_654_p N_A_1199_419#_M1019_d 0.0159428f $X=6.81 $Y=2.98
+ $X2=0 $Y2=0
cc_533 N_A_986_409#_c_661_p N_A_1199_419#_M1019_d 6.69812e-19 $X=6.035 $Y=2.98
+ $X2=0 $Y2=0
cc_534 N_A_986_409#_c_649_p N_A_1199_419#_M1036_g 0.0187081f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_535 N_A_986_409#_c_649_p N_A_1199_419#_M1043_g 0.0211617f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_536 N_A_986_409#_M1042_g N_A_1199_419#_M1008_g 0.041776f $X=9.955 $Y=0.835
+ $X2=0 $Y2=0
cc_537 N_A_986_409#_c_629_n N_A_1199_419#_c_911_n 0.00968448f $X=9.935 $Y=2.505
+ $X2=0 $Y2=0
cc_538 N_A_986_409#_c_636_n N_A_1199_419#_c_911_n 7.44355e-19 $X=10.18 $Y=1.465
+ $X2=0 $Y2=0
cc_539 N_A_986_409#_c_649_p N_A_1199_419#_c_931_n 2.21279e-19 $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_540 N_A_986_409#_M1019_g N_A_1199_419#_c_947_n 0.00152258f $X=5.87 $Y=2.595
+ $X2=0 $Y2=0
cc_541 N_A_986_409#_c_643_n N_A_1199_419#_c_947_n 0.0343853f $X=6.035 $Y=2.895
+ $X2=0 $Y2=0
cc_542 N_A_986_409#_c_654_p N_A_1199_419#_c_947_n 0.0194739f $X=6.81 $Y=2.98
+ $X2=0 $Y2=0
cc_543 N_A_986_409#_c_655_p N_A_1199_419#_c_947_n 0.00269616f $X=6.895 $Y=2.895
+ $X2=0 $Y2=0
cc_544 N_A_986_409#_c_672_p N_A_1199_419#_c_947_n 0.0129587f $X=6.98 $Y=2.59
+ $X2=0 $Y2=0
cc_545 N_A_986_409#_c_627_n N_A_1199_419#_c_932_n 0.00881594f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_546 N_A_986_409#_c_628_n N_A_1199_419#_c_932_n 0.00201348f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_547 N_A_986_409#_c_654_p N_A_1199_419#_c_932_n 0.00396791f $X=6.81 $Y=2.98
+ $X2=0 $Y2=0
cc_548 N_A_986_409#_c_649_p N_A_1199_419#_c_932_n 0.0110988f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_549 N_A_986_409#_c_672_p N_A_1199_419#_c_932_n 0.00637416f $X=6.98 $Y=2.59
+ $X2=0 $Y2=0
cc_550 N_A_986_409#_M1019_g N_A_1199_419#_c_933_n 6.20042e-19 $X=5.87 $Y=2.595
+ $X2=0 $Y2=0
cc_551 N_A_986_409#_c_643_n N_A_1199_419#_c_933_n 0.0133149f $X=6.035 $Y=2.895
+ $X2=0 $Y2=0
cc_552 N_A_986_409#_c_627_n N_A_1199_419#_c_933_n 0.0142118f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_553 N_A_986_409#_M1045_g N_A_1199_419#_c_912_n 0.0117957f $X=6.84 $Y=0.835
+ $X2=0 $Y2=0
cc_554 N_A_986_409#_c_627_n N_A_1199_419#_c_912_n 0.0096427f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_555 N_A_986_409#_c_628_n N_A_1199_419#_c_912_n 8.62438e-19 $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_556 N_A_986_409#_M1045_g N_A_1199_419#_c_913_n 0.00557216f $X=6.84 $Y=0.835
+ $X2=0 $Y2=0
cc_557 N_A_986_409#_c_627_n N_A_1199_419#_c_913_n 0.0250966f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_558 N_A_986_409#_c_628_n N_A_1199_419#_c_913_n 5.47377e-19 $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_559 N_A_986_409#_c_649_p N_A_1199_419#_c_918_n 6.40744e-19 $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_560 N_A_986_409#_M1045_g N_A_1199_419#_c_924_n 0.00238746f $X=6.84 $Y=0.835
+ $X2=0 $Y2=0
cc_561 N_A_986_409#_c_627_n N_A_1199_419#_c_924_n 0.0217436f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_562 N_A_986_409#_c_628_n N_A_1199_419#_c_924_n 0.00352136f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_563 N_A_986_409#_M1042_g N_A_1199_419#_c_925_n 3.5045e-19 $X=9.955 $Y=0.835
+ $X2=0 $Y2=0
cc_564 N_A_986_409#_c_649_p N_A_1199_419#_c_925_n 0.00337217f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_565 N_A_986_409#_c_629_n N_A_1199_419#_c_925_n 0.0182476f $X=9.935 $Y=2.505
+ $X2=0 $Y2=0
cc_566 N_A_986_409#_c_635_n N_A_1199_419#_c_925_n 2.69668e-19 $X=10.015 $Y=1.465
+ $X2=0 $Y2=0
cc_567 N_A_986_409#_c_636_n N_A_1199_419#_c_925_n 0.0218887f $X=10.18 $Y=1.465
+ $X2=0 $Y2=0
cc_568 N_A_986_409#_c_635_n N_A_1199_419#_c_926_n 0.0209697f $X=10.015 $Y=1.465
+ $X2=0 $Y2=0
cc_569 N_A_986_409#_c_649_p N_SET_B_M1010_g 0.0226293f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_570 N_A_986_409#_M1013_g N_SET_B_c_1103_n 0.00795378f $X=10.905 $Y=2.595
+ $X2=0 $Y2=0
cc_571 N_A_986_409#_c_649_p N_SET_B_c_1103_n 0.0224065f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_572 N_A_986_409#_c_629_n N_SET_B_c_1103_n 0.0220497f $X=9.935 $Y=2.505 $X2=0
+ $Y2=0
cc_573 N_A_986_409#_c_630_n N_SET_B_c_1103_n 0.00950669f $X=10.75 $Y=1.545 $X2=0
+ $Y2=0
cc_574 N_A_986_409#_c_635_n N_SET_B_c_1103_n 8.24116e-19 $X=10.015 $Y=1.465
+ $X2=0 $Y2=0
cc_575 N_A_986_409#_c_636_n N_SET_B_c_1103_n 0.021763f $X=10.18 $Y=1.465 $X2=0
+ $Y2=0
cc_576 N_A_986_409#_c_637_n N_SET_B_c_1103_n 7.08039e-19 $X=10.915 $Y=1.77 $X2=0
+ $Y2=0
cc_577 N_A_986_409#_c_649_p N_SET_B_c_1117_n 0.00355211f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_578 N_A_986_409#_c_649_p N_SET_B_c_1098_n 0.0084572f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_579 N_A_986_409#_c_649_p N_SET_B_c_1099_n 0.00104218f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_580 N_A_986_409#_c_640_n N_A_750_108#_M1035_g 0.00911739f $X=5.07 $Y=2.535
+ $X2=0 $Y2=0
cc_581 N_A_986_409#_c_642_n N_A_750_108#_M1035_g 0.00358952f $X=5.235 $Y=2.98
+ $X2=0 $Y2=0
cc_582 N_A_986_409#_c_631_n N_A_750_108#_M1031_g 2.85022e-19 $X=5.715 $Y=0.797
+ $X2=0 $Y2=0
cc_583 N_A_986_409#_c_632_n N_A_750_108#_c_1220_n 3.17403e-19 $X=5.875 $Y=1.465
+ $X2=0 $Y2=0
cc_584 N_A_986_409#_c_634_n N_A_750_108#_c_1220_n 4.73556e-19 $X=5.83 $Y=1.675
+ $X2=0 $Y2=0
cc_585 N_A_986_409#_c_631_n N_A_750_108#_M1030_g 0.00482427f $X=5.715 $Y=0.797
+ $X2=0 $Y2=0
cc_586 N_A_986_409#_c_633_n N_A_750_108#_M1030_g 0.00275279f $X=5.875 $Y=1.3
+ $X2=0 $Y2=0
cc_587 N_A_986_409#_c_631_n N_A_750_108#_c_1223_n 0.00776483f $X=5.715 $Y=0.797
+ $X2=0 $Y2=0
cc_588 N_A_986_409#_c_632_n N_A_750_108#_c_1223_n 0.0086844f $X=5.875 $Y=1.465
+ $X2=0 $Y2=0
cc_589 N_A_986_409#_c_633_n N_A_750_108#_c_1223_n 0.0162166f $X=5.875 $Y=1.3
+ $X2=0 $Y2=0
cc_590 N_A_986_409#_c_634_n N_A_750_108#_c_1223_n 0.0170355f $X=5.83 $Y=1.675
+ $X2=0 $Y2=0
cc_591 N_A_986_409#_M1045_g N_A_750_108#_M1020_g 0.0223259f $X=6.84 $Y=0.835
+ $X2=0 $Y2=0
cc_592 N_A_986_409#_c_633_n N_A_750_108#_M1020_g 0.00158157f $X=5.875 $Y=1.3
+ $X2=0 $Y2=0
cc_593 N_A_986_409#_c_627_n N_A_750_108#_c_1225_n 0.0238185f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_594 N_A_986_409#_c_628_n N_A_750_108#_c_1225_n 0.0213403f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_595 N_A_986_409#_c_632_n N_A_750_108#_c_1225_n 0.00666406f $X=5.875 $Y=1.465
+ $X2=0 $Y2=0
cc_596 N_A_986_409#_c_633_n N_A_750_108#_c_1225_n 7.7427e-19 $X=5.875 $Y=1.3
+ $X2=0 $Y2=0
cc_597 N_A_986_409#_c_634_n N_A_750_108#_c_1225_n 0.0160542f $X=5.83 $Y=1.675
+ $X2=0 $Y2=0
cc_598 N_A_986_409#_M1045_g N_A_750_108#_c_1226_n 0.00865213f $X=6.84 $Y=0.835
+ $X2=0 $Y2=0
cc_599 N_A_986_409#_M1042_g N_A_750_108#_c_1226_n 0.00907339f $X=9.955 $Y=0.835
+ $X2=0 $Y2=0
cc_600 N_A_986_409#_c_627_n N_A_750_108#_c_1240_n 0.0057037f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_601 N_A_986_409#_c_628_n N_A_750_108#_c_1240_n 0.016667f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_602 N_A_986_409#_M1019_g N_A_750_108#_c_1241_n 0.0160542f $X=5.87 $Y=2.595
+ $X2=0 $Y2=0
cc_603 N_A_986_409#_c_643_n N_A_750_108#_c_1241_n 0.00500669f $X=6.035 $Y=2.895
+ $X2=0 $Y2=0
cc_604 N_A_986_409#_M1019_g N_A_750_108#_c_1242_n 0.0145942f $X=5.87 $Y=2.595
+ $X2=0 $Y2=0
cc_605 N_A_986_409#_c_643_n N_A_750_108#_c_1242_n 0.00490093f $X=6.035 $Y=2.895
+ $X2=0 $Y2=0
cc_606 N_A_986_409#_c_654_p N_A_750_108#_c_1242_n 0.0160827f $X=6.81 $Y=2.98
+ $X2=0 $Y2=0
cc_607 N_A_986_409#_c_655_p N_A_750_108#_c_1242_n 0.00991566f $X=6.895 $Y=2.895
+ $X2=0 $Y2=0
cc_608 N_A_986_409#_c_672_p N_A_750_108#_c_1242_n 0.0060717f $X=6.98 $Y=2.59
+ $X2=0 $Y2=0
cc_609 N_A_986_409#_M1013_g N_A_750_108#_c_1243_n 0.0144374f $X=10.905 $Y=2.595
+ $X2=0 $Y2=0
cc_610 N_A_986_409#_c_649_p N_A_750_108#_c_1243_n 0.00882806f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_611 N_A_986_409#_c_629_n N_A_750_108#_c_1243_n 0.0126461f $X=9.935 $Y=2.505
+ $X2=0 $Y2=0
cc_612 N_A_986_409#_M1013_g N_A_750_108#_c_1244_n 0.00530853f $X=10.905 $Y=2.595
+ $X2=0 $Y2=0
cc_613 N_A_986_409#_c_630_n N_A_750_108#_c_1244_n 0.00491141f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_614 N_A_986_409#_c_629_n N_A_750_108#_c_1245_n 0.00909518f $X=9.935 $Y=2.505
+ $X2=0 $Y2=0
cc_615 N_A_986_409#_c_635_n N_A_750_108#_c_1245_n 0.0171208f $X=10.015 $Y=1.465
+ $X2=0 $Y2=0
cc_616 N_A_986_409#_c_636_n N_A_750_108#_c_1245_n 0.00124929f $X=10.18 $Y=1.465
+ $X2=0 $Y2=0
cc_617 N_A_986_409#_c_629_n N_A_750_108#_c_1228_n 0.00663125f $X=9.935 $Y=2.505
+ $X2=0 $Y2=0
cc_618 N_A_986_409#_c_630_n N_A_750_108#_c_1228_n 0.0153262f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_619 N_A_986_409#_c_635_n N_A_750_108#_c_1228_n 0.0205198f $X=10.015 $Y=1.465
+ $X2=0 $Y2=0
cc_620 N_A_986_409#_c_636_n N_A_750_108#_c_1228_n 0.00106267f $X=10.18 $Y=1.465
+ $X2=0 $Y2=0
cc_621 N_A_986_409#_c_637_n N_A_750_108#_c_1228_n 0.0216102f $X=10.915 $Y=1.77
+ $X2=0 $Y2=0
cc_622 N_A_986_409#_M1042_g N_A_750_108#_M1039_g 0.0134082f $X=9.955 $Y=0.835
+ $X2=0 $Y2=0
cc_623 N_A_986_409#_M1042_g N_A_750_108#_c_1233_n 0.00744792f $X=9.955 $Y=0.835
+ $X2=0 $Y2=0
cc_624 N_A_986_409#_c_630_n N_A_750_108#_c_1233_n 0.00223464f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_625 N_A_986_409#_M1035_d N_A_750_108#_c_1249_n 0.00278829f $X=4.93 $Y=2.045
+ $X2=0 $Y2=0
cc_626 N_A_986_409#_M1019_g N_A_750_108#_c_1249_n 5.41252e-19 $X=5.87 $Y=2.595
+ $X2=0 $Y2=0
cc_627 N_A_986_409#_c_640_n N_A_750_108#_c_1249_n 0.0116184f $X=5.07 $Y=2.535
+ $X2=0 $Y2=0
cc_628 N_A_986_409#_M1019_g N_A_750_108#_c_1236_n 5.48299e-19 $X=5.87 $Y=2.595
+ $X2=0 $Y2=0
cc_629 N_A_986_409#_c_640_n N_A_750_108#_c_1236_n 0.00140188f $X=5.07 $Y=2.535
+ $X2=0 $Y2=0
cc_630 N_A_986_409#_c_634_n N_A_750_108#_c_1236_n 0.0046034f $X=5.83 $Y=1.675
+ $X2=0 $Y2=0
cc_631 N_A_986_409#_c_630_n N_A_2172_40#_c_1429_n 0.0021382f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_632 N_A_986_409#_c_637_n N_A_2172_40#_c_1429_n 0.0119535f $X=10.915 $Y=1.77
+ $X2=0 $Y2=0
cc_633 N_A_986_409#_M1013_g N_A_2172_40#_M1033_g 0.0602571f $X=10.905 $Y=2.595
+ $X2=0 $Y2=0
cc_634 N_A_986_409#_c_630_n N_A_2172_40#_c_1436_n 0.00118771f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_635 N_A_986_409#_c_637_n N_A_2172_40#_c_1436_n 0.0173564f $X=10.915 $Y=1.77
+ $X2=0 $Y2=0
cc_636 N_A_986_409#_M1042_g N_A_2006_125#_c_1523_n 0.00401673f $X=9.955 $Y=0.835
+ $X2=0 $Y2=0
cc_637 N_A_986_409#_c_649_p N_A_2006_125#_c_1541_n 0.0114736f $X=9.85 $Y=2.59
+ $X2=0 $Y2=0
cc_638 N_A_986_409#_c_630_n N_A_2006_125#_c_1524_n 0.0229278f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_639 N_A_986_409#_c_637_n N_A_2006_125#_c_1524_n 6.04575e-19 $X=10.915 $Y=1.77
+ $X2=0 $Y2=0
cc_640 N_A_986_409#_M1042_g N_A_2006_125#_c_1525_n 0.00183568f $X=9.955 $Y=0.835
+ $X2=0 $Y2=0
cc_641 N_A_986_409#_c_630_n N_A_2006_125#_c_1525_n 0.0162186f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_642 N_A_986_409#_c_635_n N_A_2006_125#_c_1525_n 0.00216175f $X=10.015
+ $Y=1.465 $X2=0 $Y2=0
cc_643 N_A_986_409#_c_636_n N_A_2006_125#_c_1525_n 0.00671973f $X=10.18 $Y=1.465
+ $X2=0 $Y2=0
cc_644 N_A_986_409#_M1013_g N_A_2006_125#_c_1548_n 0.0195375f $X=10.905 $Y=2.595
+ $X2=0 $Y2=0
cc_645 N_A_986_409#_c_630_n N_A_2006_125#_c_1548_n 0.00524002f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_646 N_A_986_409#_M1013_g N_A_2006_125#_c_1526_n 0.00484557f $X=10.905
+ $Y=2.595 $X2=0 $Y2=0
cc_647 N_A_986_409#_c_630_n N_A_2006_125#_c_1526_n 0.0345858f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_648 N_A_986_409#_c_637_n N_A_2006_125#_c_1526_n 0.00196901f $X=10.915 $Y=1.77
+ $X2=0 $Y2=0
cc_649 N_A_986_409#_M1013_g N_A_2006_125#_c_1538_n 0.0188768f $X=10.905 $Y=2.595
+ $X2=0 $Y2=0
cc_650 N_A_986_409#_c_629_n N_A_2006_125#_c_1538_n 0.0257837f $X=9.935 $Y=2.505
+ $X2=0 $Y2=0
cc_651 N_A_986_409#_c_630_n N_A_2006_125#_c_1538_n 0.00766198f $X=10.75 $Y=1.545
+ $X2=0 $Y2=0
cc_652 N_A_986_409#_c_649_p N_VPWR_M1009_d 0.0153853f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_653 N_A_986_409#_c_649_p N_VPWR_M1010_d 0.0150829f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_654 N_A_986_409#_c_640_n N_VPWR_c_1768_n 0.0345597f $X=5.07 $Y=2.535 $X2=0
+ $Y2=0
cc_655 N_A_986_409#_c_642_n N_VPWR_c_1768_n 0.0119061f $X=5.235 $Y=2.98 $X2=0
+ $Y2=0
cc_656 N_A_986_409#_c_649_p N_VPWR_c_1769_n 0.0238466f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_657 N_A_986_409#_c_649_p N_VPWR_c_1770_n 0.0196062f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_658 N_A_986_409#_M1013_g N_VPWR_c_1771_n 0.00263095f $X=10.905 $Y=2.595 $X2=0
+ $Y2=0
cc_659 N_A_986_409#_M1019_g N_VPWR_c_1779_n 0.00599878f $X=5.87 $Y=2.595 $X2=0
+ $Y2=0
cc_660 N_A_986_409#_c_641_n N_VPWR_c_1779_n 0.040934f $X=5.95 $Y=2.98 $X2=0
+ $Y2=0
cc_661 N_A_986_409#_c_642_n N_VPWR_c_1779_n 0.0221998f $X=5.235 $Y=2.98 $X2=0
+ $Y2=0
cc_662 N_A_986_409#_c_654_p N_VPWR_c_1779_n 0.0483813f $X=6.81 $Y=2.98 $X2=0
+ $Y2=0
cc_663 N_A_986_409#_c_649_p N_VPWR_c_1779_n 0.00656068f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_664 N_A_986_409#_c_661_p N_VPWR_c_1779_n 0.0092477f $X=6.035 $Y=2.98 $X2=0
+ $Y2=0
cc_665 N_A_986_409#_c_649_p N_VPWR_c_1780_n 0.01523f $X=9.85 $Y=2.59 $X2=0 $Y2=0
cc_666 N_A_986_409#_M1013_g N_VPWR_c_1781_n 0.00975641f $X=10.905 $Y=2.595 $X2=0
+ $Y2=0
cc_667 N_A_986_409#_c_649_p N_VPWR_c_1781_n 0.0135362f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_668 N_A_986_409#_M1019_g N_VPWR_c_1765_n 0.0100086f $X=5.87 $Y=2.595 $X2=0
+ $Y2=0
cc_669 N_A_986_409#_M1013_g N_VPWR_c_1765_n 0.0105056f $X=10.905 $Y=2.595 $X2=0
+ $Y2=0
cc_670 N_A_986_409#_c_641_n N_VPWR_c_1765_n 0.0257755f $X=5.95 $Y=2.98 $X2=0
+ $Y2=0
cc_671 N_A_986_409#_c_642_n N_VPWR_c_1765_n 0.0126612f $X=5.235 $Y=2.98 $X2=0
+ $Y2=0
cc_672 N_A_986_409#_c_654_p N_VPWR_c_1765_n 0.0311775f $X=6.81 $Y=2.98 $X2=0
+ $Y2=0
cc_673 N_A_986_409#_c_649_p N_VPWR_c_1765_n 0.0646345f $X=9.85 $Y=2.59 $X2=0
+ $Y2=0
cc_674 N_A_986_409#_c_661_p N_VPWR_c_1765_n 0.00636511f $X=6.035 $Y=2.98 $X2=0
+ $Y2=0
cc_675 N_A_986_409#_c_641_n N_A_352_406#_M1019_s 0.00534965f $X=5.95 $Y=2.98
+ $X2=0 $Y2=0
cc_676 N_A_986_409#_c_631_n N_A_352_406#_c_1999_n 0.0144118f $X=5.715 $Y=0.797
+ $X2=0 $Y2=0
cc_677 N_A_986_409#_c_633_n N_A_352_406#_c_1999_n 0.0063732f $X=5.875 $Y=1.3
+ $X2=0 $Y2=0
cc_678 N_A_986_409#_c_631_n N_A_352_406#_c_2000_n 0.0304199f $X=5.715 $Y=0.797
+ $X2=0 $Y2=0
cc_679 N_A_986_409#_M1019_g N_A_352_406#_c_2009_n 0.01181f $X=5.87 $Y=2.595
+ $X2=0 $Y2=0
cc_680 N_A_986_409#_c_640_n N_A_352_406#_c_2009_n 0.0251928f $X=5.07 $Y=2.535
+ $X2=0 $Y2=0
cc_681 N_A_986_409#_c_641_n N_A_352_406#_c_2009_n 0.0196819f $X=5.95 $Y=2.98
+ $X2=0 $Y2=0
cc_682 N_A_986_409#_c_627_n N_A_352_406#_c_2002_n 0.00204395f $X=6.73 $Y=1.465
+ $X2=0 $Y2=0
cc_683 N_A_986_409#_c_631_n N_A_352_406#_c_2002_n 0.0280321f $X=5.715 $Y=0.797
+ $X2=0 $Y2=0
cc_684 N_A_986_409#_c_632_n N_A_352_406#_c_2002_n 0.0102745f $X=5.875 $Y=1.465
+ $X2=0 $Y2=0
cc_685 N_A_986_409#_c_633_n N_A_352_406#_c_2002_n 0.00605939f $X=5.875 $Y=1.3
+ $X2=0 $Y2=0
cc_686 N_A_986_409#_c_631_n N_A_352_406#_c_2004_n 0.00788995f $X=5.715 $Y=0.797
+ $X2=0 $Y2=0
cc_687 N_A_986_409#_c_633_n N_A_352_406#_c_2004_n 0.0128609f $X=5.875 $Y=1.3
+ $X2=0 $Y2=0
cc_688 N_A_986_409#_M1019_g N_A_352_406#_c_2005_n 0.00330551f $X=5.87 $Y=2.595
+ $X2=0 $Y2=0
cc_689 N_A_986_409#_c_643_n N_A_352_406#_c_2005_n 0.00569922f $X=6.035 $Y=2.895
+ $X2=0 $Y2=0
cc_690 N_A_986_409#_c_632_n N_A_352_406#_c_2005_n 0.0400899f $X=5.875 $Y=1.465
+ $X2=0 $Y2=0
cc_691 N_A_986_409#_c_634_n N_A_352_406#_c_2005_n 0.00117547f $X=5.83 $Y=1.675
+ $X2=0 $Y2=0
cc_692 N_A_986_409#_M1019_g N_A_352_406#_c_2011_n 0.00702305f $X=5.87 $Y=2.595
+ $X2=0 $Y2=0
cc_693 N_A_986_409#_c_643_n N_A_352_406#_c_2011_n 0.0477521f $X=6.035 $Y=2.895
+ $X2=0 $Y2=0
cc_694 N_A_986_409#_c_632_n N_A_352_406#_c_2011_n 0.011847f $X=5.875 $Y=1.465
+ $X2=0 $Y2=0
cc_695 N_A_986_409#_c_634_n N_A_352_406#_c_2011_n 6.26457e-19 $X=5.83 $Y=1.675
+ $X2=0 $Y2=0
cc_696 N_A_986_409#_c_654_p A_1371_419# 0.00292004f $X=6.81 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_697 N_A_986_409#_c_655_p A_1371_419# 0.00254812f $X=6.895 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_698 N_A_986_409#_c_649_p A_1371_419# 0.00294021f $X=9.85 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_699 N_A_986_409#_c_672_p A_1371_419# 9.0912e-19 $X=6.98 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_700 N_A_986_409#_c_649_p A_1928_419# 0.00434279f $X=9.85 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_701 N_A_986_409#_M1045_g N_VGND_c_2223_n 9.49986e-19 $X=6.84 $Y=0.835 $X2=0
+ $Y2=0
cc_702 N_A_986_409#_M1042_g N_VGND_c_2223_n 9.49986e-19 $X=9.955 $Y=0.835 $X2=0
+ $Y2=0
cc_703 N_A_1425_99#_M1009_g N_A_1199_419#_M1036_g 0.0204793f $X=7.26 $Y=2.595
+ $X2=0 $Y2=0
cc_704 N_A_1425_99#_c_839_n N_A_1199_419#_M1036_g 0.00433088f $X=7.59 $Y=2.075
+ $X2=0 $Y2=0
cc_705 N_A_1425_99#_c_841_n N_A_1199_419#_M1036_g 0.0180572f $X=8.425 $Y=2.24
+ $X2=0 $Y2=0
cc_706 N_A_1425_99#_c_832_n N_A_1199_419#_c_908_n 0.00949949f $X=7.26 $Y=1.885
+ $X2=0 $Y2=0
cc_707 N_A_1425_99#_c_834_n N_A_1199_419#_c_908_n 0.007556f $X=8.095 $Y=1.3
+ $X2=0 $Y2=0
cc_708 N_A_1425_99#_c_836_n N_A_1199_419#_c_908_n 0.00701034f $X=8.39 $Y=0.84
+ $X2=0 $Y2=0
cc_709 N_A_1425_99#_c_835_n N_A_1199_419#_M1025_g 0.002946f $X=8.18 $Y=1.215
+ $X2=0 $Y2=0
cc_710 N_A_1425_99#_c_836_n N_A_1199_419#_M1025_g 0.0064556f $X=8.39 $Y=0.84
+ $X2=0 $Y2=0
cc_711 N_A_1425_99#_M1009_g N_A_1199_419#_c_947_n 0.00122719f $X=7.26 $Y=2.595
+ $X2=0 $Y2=0
cc_712 N_A_1425_99#_M1009_g N_A_1199_419#_c_932_n 0.00728523f $X=7.26 $Y=2.595
+ $X2=0 $Y2=0
cc_713 N_A_1425_99#_c_840_n N_A_1199_419#_c_932_n 0.00772304f $X=7.755 $Y=2.2
+ $X2=0 $Y2=0
cc_714 N_A_1425_99#_M1034_g N_A_1199_419#_c_913_n 0.00752601f $X=7.2 $Y=0.835
+ $X2=0 $Y2=0
cc_715 N_A_1425_99#_c_832_n N_A_1199_419#_c_913_n 0.0218441f $X=7.26 $Y=1.885
+ $X2=0 $Y2=0
cc_716 N_A_1425_99#_M1009_g N_A_1199_419#_c_913_n 0.00455902f $X=7.26 $Y=2.595
+ $X2=0 $Y2=0
cc_717 N_A_1425_99#_c_833_n N_A_1199_419#_c_913_n 0.0123662f $X=7.59 $Y=1.385
+ $X2=0 $Y2=0
cc_718 N_A_1425_99#_c_839_n N_A_1199_419#_c_913_n 0.0477088f $X=7.59 $Y=2.075
+ $X2=0 $Y2=0
cc_719 N_A_1425_99#_M1034_g N_A_1199_419#_c_914_n 0.00623975f $X=7.2 $Y=0.835
+ $X2=0 $Y2=0
cc_720 N_A_1425_99#_c_832_n N_A_1199_419#_c_914_n 0.00744269f $X=7.26 $Y=1.885
+ $X2=0 $Y2=0
cc_721 N_A_1425_99#_c_833_n N_A_1199_419#_c_914_n 0.025034f $X=7.59 $Y=1.385
+ $X2=0 $Y2=0
cc_722 N_A_1425_99#_c_834_n N_A_1199_419#_c_914_n 0.0129405f $X=8.095 $Y=1.3
+ $X2=0 $Y2=0
cc_723 N_A_1425_99#_c_836_n N_A_1199_419#_c_914_n 0.0148555f $X=8.39 $Y=0.84
+ $X2=0 $Y2=0
cc_724 N_A_1425_99#_M1034_g N_A_1199_419#_c_915_n 0.00473436f $X=7.2 $Y=0.835
+ $X2=0 $Y2=0
cc_725 N_A_1425_99#_c_836_n N_A_1199_419#_c_915_n 0.0195222f $X=8.39 $Y=0.84
+ $X2=0 $Y2=0
cc_726 N_A_1425_99#_c_836_n N_A_1199_419#_c_916_n 0.0334088f $X=8.39 $Y=0.84
+ $X2=0 $Y2=0
cc_727 N_A_1425_99#_c_832_n N_A_1199_419#_c_918_n 0.00132319f $X=7.26 $Y=1.885
+ $X2=0 $Y2=0
cc_728 N_A_1425_99#_c_839_n N_A_1199_419#_c_918_n 0.0197405f $X=7.59 $Y=2.075
+ $X2=0 $Y2=0
cc_729 N_A_1425_99#_c_834_n N_A_1199_419#_c_918_n 0.0197186f $X=8.095 $Y=1.3
+ $X2=0 $Y2=0
cc_730 N_A_1425_99#_c_841_n N_A_1199_419#_c_918_n 0.0443808f $X=8.425 $Y=2.24
+ $X2=0 $Y2=0
cc_731 N_A_1425_99#_c_836_n N_A_1199_419#_c_918_n 0.0070016f $X=8.39 $Y=0.84
+ $X2=0 $Y2=0
cc_732 N_A_1425_99#_c_832_n N_A_1199_419#_c_919_n 0.0179213f $X=7.26 $Y=1.885
+ $X2=0 $Y2=0
cc_733 N_A_1425_99#_c_839_n N_A_1199_419#_c_919_n 4.48216e-19 $X=7.59 $Y=2.075
+ $X2=0 $Y2=0
cc_734 N_A_1425_99#_c_834_n N_A_1199_419#_c_919_n 0.00458383f $X=8.095 $Y=1.3
+ $X2=0 $Y2=0
cc_735 N_A_1425_99#_c_841_n N_A_1199_419#_c_919_n 0.00194249f $X=8.425 $Y=2.24
+ $X2=0 $Y2=0
cc_736 N_A_1425_99#_c_834_n N_A_1199_419#_c_921_n 0.00110685f $X=8.095 $Y=1.3
+ $X2=0 $Y2=0
cc_737 N_A_1425_99#_c_835_n N_A_1199_419#_c_921_n 0.00553806f $X=8.18 $Y=1.215
+ $X2=0 $Y2=0
cc_738 N_A_1425_99#_c_836_n N_A_1199_419#_c_921_n 0.0179238f $X=8.39 $Y=0.84
+ $X2=0 $Y2=0
cc_739 N_A_1425_99#_c_834_n N_A_1199_419#_c_923_n 0.0112835f $X=8.095 $Y=1.3
+ $X2=0 $Y2=0
cc_740 N_A_1425_99#_c_836_n N_A_1199_419#_c_923_n 0.00802851f $X=8.39 $Y=0.84
+ $X2=0 $Y2=0
cc_741 N_A_1425_99#_M1034_g N_A_1199_419#_c_1014_n 0.00673013f $X=7.2 $Y=0.835
+ $X2=0 $Y2=0
cc_742 N_A_1425_99#_c_839_n N_A_1199_419#_c_927_n 0.00101368f $X=7.59 $Y=2.075
+ $X2=0 $Y2=0
cc_743 N_A_1425_99#_c_834_n N_A_1199_419#_c_927_n 0.00187457f $X=8.095 $Y=1.3
+ $X2=0 $Y2=0
cc_744 N_A_1425_99#_c_841_n N_SET_B_M1010_g 0.010625f $X=8.425 $Y=2.24 $X2=0
+ $Y2=0
cc_745 N_A_1425_99#_c_841_n N_SET_B_c_1117_n 0.0021036f $X=8.425 $Y=2.24 $X2=0
+ $Y2=0
cc_746 N_A_1425_99#_c_841_n N_SET_B_c_1098_n 0.00395695f $X=8.425 $Y=2.24 $X2=0
+ $Y2=0
cc_747 N_A_1425_99#_M1034_g N_A_750_108#_c_1226_n 0.00865126f $X=7.2 $Y=0.835
+ $X2=0 $Y2=0
cc_748 N_A_1425_99#_c_832_n N_A_750_108#_c_1240_n 0.0309379f $X=7.26 $Y=1.885
+ $X2=0 $Y2=0
cc_749 N_A_1425_99#_M1009_g N_A_750_108#_c_1242_n 0.0309379f $X=7.26 $Y=2.595
+ $X2=0 $Y2=0
cc_750 N_A_1425_99#_c_840_n N_VPWR_M1009_d 0.00754175f $X=7.755 $Y=2.2 $X2=0
+ $Y2=0
cc_751 N_A_1425_99#_c_841_n N_VPWR_M1009_d 0.00370683f $X=8.425 $Y=2.24 $X2=0
+ $Y2=0
cc_752 N_A_1425_99#_M1009_g N_VPWR_c_1769_n 0.00568281f $X=7.26 $Y=2.595 $X2=0
+ $Y2=0
cc_753 N_A_1425_99#_M1009_g N_VPWR_c_1779_n 0.00713369f $X=7.26 $Y=2.595 $X2=0
+ $Y2=0
cc_754 N_A_1425_99#_M1036_d N_VPWR_c_1765_n 0.00333718f $X=8.285 $Y=2.095 $X2=0
+ $Y2=0
cc_755 N_A_1425_99#_M1009_g N_VPWR_c_1765_n 0.00963348f $X=7.26 $Y=2.595 $X2=0
+ $Y2=0
cc_756 N_A_1425_99#_M1034_g N_VGND_c_2206_n 0.00627416f $X=7.2 $Y=0.835 $X2=0
+ $Y2=0
cc_757 N_A_1425_99#_M1034_g N_VGND_c_2223_n 9.49986e-19 $X=7.2 $Y=0.835 $X2=0
+ $Y2=0
cc_758 N_A_1199_419#_M1043_g N_SET_B_M1010_g 0.0238257f $X=9.515 $Y=2.595 $X2=0
+ $Y2=0
cc_759 N_A_1199_419#_M1025_g N_SET_B_M1014_g 0.0391973f $X=8.605 $Y=0.835 $X2=0
+ $Y2=0
cc_760 N_A_1199_419#_M1008_g N_SET_B_M1014_g 0.0125976f $X=9.565 $Y=0.835 $X2=0
+ $Y2=0
cc_761 N_A_1199_419#_c_918_n N_SET_B_M1014_g 0.00100389f $X=8.445 $Y=1.73 $X2=0
+ $Y2=0
cc_762 N_A_1199_419#_c_920_n N_SET_B_M1014_g 0.00297973f $X=8.53 $Y=1.565 $X2=0
+ $Y2=0
cc_763 N_A_1199_419#_c_921_n N_SET_B_M1014_g 0.00716454f $X=8.82 $Y=1.245 $X2=0
+ $Y2=0
cc_764 N_A_1199_419#_c_922_n N_SET_B_M1014_g 0.0149663f $X=9.31 $Y=1.33 $X2=0
+ $Y2=0
cc_765 N_A_1199_419#_c_925_n N_SET_B_M1014_g 0.00122465f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_766 N_A_1199_419#_c_926_n N_SET_B_M1014_g 0.0194015f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_767 N_A_1199_419#_c_927_n N_SET_B_M1014_g 0.00289763f $X=8.16 $Y=1.565 $X2=0
+ $Y2=0
cc_768 N_A_1199_419#_M1043_g N_SET_B_c_1103_n 0.00882558f $X=9.515 $Y=2.595
+ $X2=0 $Y2=0
cc_769 N_A_1199_419#_c_922_n N_SET_B_c_1103_n 0.00692633f $X=9.31 $Y=1.33 $X2=0
+ $Y2=0
cc_770 N_A_1199_419#_c_925_n N_SET_B_c_1103_n 0.0114042f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_771 N_A_1199_419#_M1036_g N_SET_B_c_1117_n 7.27401e-19 $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_772 N_A_1199_419#_c_923_n N_SET_B_c_1117_n 0.00276155f $X=8.905 $Y=1.33 $X2=0
+ $Y2=0
cc_773 N_A_1199_419#_M1036_g N_SET_B_c_1098_n 0.00127749f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_774 N_A_1199_419#_M1043_g N_SET_B_c_1098_n 0.00405655f $X=9.515 $Y=2.595
+ $X2=0 $Y2=0
cc_775 N_A_1199_419#_c_911_n N_SET_B_c_1098_n 0.00107725f $X=9.475 $Y=1.75 $X2=0
+ $Y2=0
cc_776 N_A_1199_419#_c_918_n N_SET_B_c_1098_n 0.0218185f $X=8.445 $Y=1.73 $X2=0
+ $Y2=0
cc_777 N_A_1199_419#_c_923_n N_SET_B_c_1098_n 0.0203881f $X=8.905 $Y=1.33 $X2=0
+ $Y2=0
cc_778 N_A_1199_419#_c_925_n N_SET_B_c_1098_n 0.0194963f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_779 N_A_1199_419#_M1036_g N_SET_B_c_1099_n 0.0502033f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_780 N_A_1199_419#_c_907_n N_SET_B_c_1099_n 0.00643005f $X=8.53 $Y=1.29 $X2=0
+ $Y2=0
cc_781 N_A_1199_419#_M1043_g N_SET_B_c_1099_n 9.70237e-19 $X=9.515 $Y=2.595
+ $X2=0 $Y2=0
cc_782 N_A_1199_419#_c_911_n N_SET_B_c_1099_n 0.0195771f $X=9.475 $Y=1.75 $X2=0
+ $Y2=0
cc_783 N_A_1199_419#_c_918_n N_SET_B_c_1099_n 0.00999645f $X=8.445 $Y=1.73 $X2=0
+ $Y2=0
cc_784 N_A_1199_419#_c_919_n N_SET_B_c_1099_n 0.0159962f $X=8.16 $Y=1.73 $X2=0
+ $Y2=0
cc_785 N_A_1199_419#_c_923_n N_SET_B_c_1099_n 0.00697957f $X=8.905 $Y=1.33 $X2=0
+ $Y2=0
cc_786 N_A_1199_419#_c_925_n N_SET_B_c_1099_n 0.00118191f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_787 N_A_1199_419#_c_924_n N_A_750_108#_M1020_g 0.00294311f $X=6.56 $Y=0.835
+ $X2=0 $Y2=0
cc_788 N_A_1199_419#_M1025_g N_A_750_108#_c_1226_n 0.00737233f $X=8.605 $Y=0.835
+ $X2=0 $Y2=0
cc_789 N_A_1199_419#_M1008_g N_A_750_108#_c_1226_n 0.00907339f $X=9.565 $Y=0.835
+ $X2=0 $Y2=0
cc_790 N_A_1199_419#_c_912_n N_A_750_108#_c_1226_n 0.003295f $X=7.075 $Y=0.965
+ $X2=0 $Y2=0
cc_791 N_A_1199_419#_c_914_n N_A_750_108#_c_1226_n 0.00473275f $X=7.745 $Y=0.95
+ $X2=0 $Y2=0
cc_792 N_A_1199_419#_c_916_n N_A_750_108#_c_1226_n 0.0209179f $X=8.735 $Y=0.35
+ $X2=0 $Y2=0
cc_793 N_A_1199_419#_c_917_n N_A_750_108#_c_1226_n 0.00418768f $X=7.915 $Y=0.35
+ $X2=0 $Y2=0
cc_794 N_A_1199_419#_c_924_n N_A_750_108#_c_1226_n 0.00537854f $X=6.56 $Y=0.835
+ $X2=0 $Y2=0
cc_795 N_A_1199_419#_c_1014_n N_A_750_108#_c_1226_n 3.82766e-19 $X=7.16 $Y=0.965
+ $X2=0 $Y2=0
cc_796 N_A_1199_419#_c_913_n N_A_750_108#_c_1240_n 0.00417154f $X=7.16 $Y=2.075
+ $X2=0 $Y2=0
cc_797 N_A_1199_419#_c_933_n N_A_750_108#_c_1241_n 0.00892503f $X=6.63 $Y=2.16
+ $X2=0 $Y2=0
cc_798 N_A_1199_419#_c_947_n N_A_750_108#_c_1242_n 0.0109411f $X=6.465 $Y=2.395
+ $X2=0 $Y2=0
cc_799 N_A_1199_419#_c_932_n N_A_750_108#_c_1242_n 0.0148744f $X=7.075 $Y=2.16
+ $X2=0 $Y2=0
cc_800 N_A_1199_419#_c_933_n N_A_750_108#_c_1242_n 0.00277341f $X=6.63 $Y=2.16
+ $X2=0 $Y2=0
cc_801 N_A_1199_419#_M1043_g N_A_750_108#_c_1243_n 0.0381472f $X=9.515 $Y=2.595
+ $X2=0 $Y2=0
cc_802 N_A_1199_419#_c_931_n N_A_750_108#_c_1245_n 0.0381472f $X=9.475 $Y=1.915
+ $X2=0 $Y2=0
cc_803 N_A_1199_419#_M1036_g N_VPWR_c_1769_n 0.0080577f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_804 N_A_1199_419#_M1036_g N_VPWR_c_1770_n 0.00189234f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_805 N_A_1199_419#_M1043_g N_VPWR_c_1770_n 0.00780519f $X=9.515 $Y=2.595 $X2=0
+ $Y2=0
cc_806 N_A_1199_419#_M1036_g N_VPWR_c_1780_n 0.00713369f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_807 N_A_1199_419#_M1043_g N_VPWR_c_1781_n 0.00713369f $X=9.515 $Y=2.595 $X2=0
+ $Y2=0
cc_808 N_A_1199_419#_M1019_d N_VPWR_c_1765_n 0.00499582f $X=5.995 $Y=2.095 $X2=0
+ $Y2=0
cc_809 N_A_1199_419#_M1036_g N_VPWR_c_1765_n 0.00975378f $X=8.16 $Y=2.595 $X2=0
+ $Y2=0
cc_810 N_A_1199_419#_M1043_g N_VPWR_c_1765_n 0.00953645f $X=9.515 $Y=2.595 $X2=0
+ $Y2=0
cc_811 N_A_1199_419#_c_924_n N_A_352_406#_c_2002_n 0.00233138f $X=6.56 $Y=0.835
+ $X2=0 $Y2=0
cc_812 N_A_1199_419#_c_932_n A_1371_419# 0.00208762f $X=7.075 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_813 N_A_1199_419#_c_914_n N_VGND_M1034_d 0.00772331f $X=7.745 $Y=0.95 $X2=0
+ $Y2=0
cc_814 N_A_1199_419#_c_914_n N_VGND_c_2206_n 0.0180852f $X=7.745 $Y=0.95 $X2=0
+ $Y2=0
cc_815 N_A_1199_419#_c_915_n N_VGND_c_2206_n 0.0182235f $X=7.83 $Y=0.865 $X2=0
+ $Y2=0
cc_816 N_A_1199_419#_c_917_n N_VGND_c_2206_n 0.0140721f $X=7.915 $Y=0.35 $X2=0
+ $Y2=0
cc_817 N_A_1199_419#_c_924_n N_VGND_c_2206_n 6.42296e-19 $X=6.56 $Y=0.835 $X2=0
+ $Y2=0
cc_818 N_A_1199_419#_M1008_g N_VGND_c_2207_n 0.00889597f $X=9.565 $Y=0.835 $X2=0
+ $Y2=0
cc_819 N_A_1199_419#_c_916_n N_VGND_c_2207_n 0.0144411f $X=8.735 $Y=0.35 $X2=0
+ $Y2=0
cc_820 N_A_1199_419#_c_921_n N_VGND_c_2207_n 0.0157946f $X=8.82 $Y=1.245 $X2=0
+ $Y2=0
cc_821 N_A_1199_419#_c_922_n N_VGND_c_2207_n 0.0181313f $X=9.31 $Y=1.33 $X2=0
+ $Y2=0
cc_822 N_A_1199_419#_c_925_n N_VGND_c_2207_n 0.00886836f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_823 N_A_1199_419#_c_926_n N_VGND_c_2207_n 8.08179e-19 $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_824 N_A_1199_419#_c_924_n N_VGND_c_2219_n 0.0068634f $X=6.56 $Y=0.835 $X2=0
+ $Y2=0
cc_825 N_A_1199_419#_c_916_n N_VGND_c_2220_n 0.0611043f $X=8.735 $Y=0.35 $X2=0
+ $Y2=0
cc_826 N_A_1199_419#_c_917_n N_VGND_c_2220_n 0.0114574f $X=7.915 $Y=0.35 $X2=0
+ $Y2=0
cc_827 N_A_1199_419#_M1008_g N_VGND_c_2223_n 9.49986e-19 $X=9.565 $Y=0.835 $X2=0
+ $Y2=0
cc_828 N_A_1199_419#_c_916_n N_VGND_c_2223_n 0.0332665f $X=8.735 $Y=0.35 $X2=0
+ $Y2=0
cc_829 N_A_1199_419#_c_917_n N_VGND_c_2223_n 0.00589978f $X=7.915 $Y=0.35 $X2=0
+ $Y2=0
cc_830 N_A_1199_419#_c_924_n N_VGND_c_2223_n 0.00870304f $X=6.56 $Y=0.835 $X2=0
+ $Y2=0
cc_831 N_A_1199_419#_c_1014_n N_VGND_c_2223_n 0.00545057f $X=7.16 $Y=0.965 $X2=0
+ $Y2=0
cc_832 N_A_1199_419#_c_912_n A_1383_125# 0.00165482f $X=7.075 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_833 N_A_1199_419#_c_921_n A_1736_125# 0.00292914f $X=8.82 $Y=1.245 $X2=-0.19
+ $Y2=-0.245
cc_834 N_SET_B_M1014_g N_A_750_108#_c_1226_n 0.00907339f $X=8.995 $Y=0.835 $X2=0
+ $Y2=0
cc_835 N_SET_B_c_1103_n N_A_750_108#_c_1243_n 0.00556136f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_836 N_SET_B_c_1103_n N_A_750_108#_c_1244_n 0.00845492f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_837 N_SET_B_c_1103_n N_A_750_108#_c_1245_n 0.00107753f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_838 N_SET_B_c_1094_n N_A_2172_40#_M1040_g 0.0433565f $X=11.325 $Y=0.825 $X2=0
+ $Y2=0
cc_839 N_SET_B_c_1096_n N_A_2172_40#_c_1428_n 0.0181626f $X=11.4 $Y=0.9 $X2=0
+ $Y2=0
cc_840 N_SET_B_c_1103_n N_A_2172_40#_c_1428_n 0.00259692f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_841 N_SET_B_c_1102_n N_A_2172_40#_M1033_g 0.0251384f $X=12.265 $Y=1.935 $X2=0
+ $Y2=0
cc_842 N_SET_B_c_1103_n N_A_2172_40#_M1033_g 0.010222f $X=12.095 $Y=2.035 $X2=0
+ $Y2=0
cc_843 SET_B N_A_2172_40#_M1033_g 0.00120324f $X=12.155 $Y=1.95 $X2=0 $Y2=0
cc_844 N_SET_B_c_1106_n N_A_2172_40#_M1033_g 0.00194194f $X=12.265 $Y=1.43 $X2=0
+ $Y2=0
cc_845 N_SET_B_c_1103_n N_A_2172_40#_c_1430_n 0.0102464f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_846 N_SET_B_c_1097_n N_A_2172_40#_c_1430_n 0.00748419f $X=12.265 $Y=1.43
+ $X2=0 $Y2=0
cc_847 N_SET_B_c_1106_n N_A_2172_40#_c_1430_n 0.0390243f $X=12.265 $Y=1.43 $X2=0
+ $Y2=0
cc_848 N_SET_B_c_1095_n N_A_2172_40#_c_1431_n 0.0274962f $X=12.1 $Y=0.9 $X2=0
+ $Y2=0
cc_849 N_SET_B_c_1097_n N_A_2172_40#_c_1431_n 0.0129849f $X=12.265 $Y=1.43 $X2=0
+ $Y2=0
cc_850 N_SET_B_c_1106_n N_A_2172_40#_c_1431_n 0.0238596f $X=12.265 $Y=1.43 $X2=0
+ $Y2=0
cc_851 N_SET_B_c_1095_n N_A_2172_40#_c_1432_n 0.0148381f $X=12.1 $Y=0.9 $X2=0
+ $Y2=0
cc_852 N_SET_B_c_1095_n N_A_2172_40#_c_1433_n 0.00277498f $X=12.1 $Y=0.9 $X2=0
+ $Y2=0
cc_853 N_SET_B_M1021_g N_A_2172_40#_c_1435_n 0.00604253f $X=12.225 $Y=2.595
+ $X2=0 $Y2=0
cc_854 SET_B N_A_2172_40#_c_1435_n 0.00147374f $X=12.155 $Y=1.95 $X2=0 $Y2=0
cc_855 N_SET_B_c_1097_n N_A_2172_40#_c_1435_n 0.0175512f $X=12.265 $Y=1.43 $X2=0
+ $Y2=0
cc_856 N_SET_B_c_1106_n N_A_2172_40#_c_1435_n 0.0319036f $X=12.265 $Y=1.43 $X2=0
+ $Y2=0
cc_857 N_SET_B_c_1095_n N_A_2172_40#_c_1436_n 0.0181626f $X=12.1 $Y=0.9 $X2=0
+ $Y2=0
cc_858 N_SET_B_c_1103_n N_A_2172_40#_c_1436_n 4.92627e-19 $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_859 N_SET_B_c_1097_n N_A_2172_40#_c_1436_n 0.0431131f $X=12.265 $Y=1.43 $X2=0
+ $Y2=0
cc_860 N_SET_B_c_1106_n N_A_2172_40#_c_1436_n 0.00241081f $X=12.265 $Y=1.43
+ $X2=0 $Y2=0
cc_861 N_SET_B_c_1103_n N_A_2006_125#_M1011_d 0.00598621f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_862 N_SET_B_c_1106_n N_A_2006_125#_M1021_d 0.00121553f $X=12.265 $Y=1.43
+ $X2=0 $Y2=0
cc_863 N_SET_B_c_1095_n N_A_2006_125#_c_1512_n 0.00523856f $X=12.1 $Y=0.9 $X2=0
+ $Y2=0
cc_864 N_SET_B_c_1095_n N_A_2006_125#_c_1524_n 8.93333e-19 $X=12.1 $Y=0.9 $X2=0
+ $Y2=0
cc_865 N_SET_B_c_1096_n N_A_2006_125#_c_1524_n 0.00993687f $X=11.4 $Y=0.9 $X2=0
+ $Y2=0
cc_866 N_SET_B_c_1097_n N_A_2006_125#_c_1524_n 3.1732e-19 $X=12.265 $Y=1.43
+ $X2=0 $Y2=0
cc_867 N_SET_B_c_1103_n N_A_2006_125#_c_1548_n 0.0224831f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_868 N_SET_B_c_1102_n N_A_2006_125#_c_1526_n 0.00200526f $X=12.265 $Y=1.935
+ $X2=0 $Y2=0
cc_869 N_SET_B_c_1103_n N_A_2006_125#_c_1526_n 0.0259073f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_870 N_SET_B_M1021_g N_A_2006_125#_c_1565_n 0.0149523f $X=12.225 $Y=2.595
+ $X2=0 $Y2=0
cc_871 N_SET_B_c_1103_n N_A_2006_125#_c_1565_n 0.0236569f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_872 SET_B N_A_2006_125#_c_1565_n 0.00179801f $X=12.155 $Y=1.95 $X2=0 $Y2=0
cc_873 N_SET_B_c_1106_n N_A_2006_125#_c_1565_n 0.0127306f $X=12.265 $Y=1.43
+ $X2=0 $Y2=0
cc_874 N_SET_B_M1021_g N_A_2006_125#_c_1533_n 7.27872e-19 $X=12.225 $Y=2.595
+ $X2=0 $Y2=0
cc_875 N_SET_B_c_1102_n N_A_2006_125#_c_1533_n 2.60945e-19 $X=12.265 $Y=1.935
+ $X2=0 $Y2=0
cc_876 SET_B N_A_2006_125#_c_1533_n 4.90986e-19 $X=12.155 $Y=1.95 $X2=0 $Y2=0
cc_877 N_SET_B_c_1106_n N_A_2006_125#_c_1533_n 0.004071f $X=12.265 $Y=1.43 $X2=0
+ $Y2=0
cc_878 N_SET_B_M1021_g N_A_2006_125#_c_1534_n 0.0125354f $X=12.225 $Y=2.595
+ $X2=0 $Y2=0
cc_879 N_SET_B_M1021_g N_A_2006_125#_c_1536_n 0.0036057f $X=12.225 $Y=2.595
+ $X2=0 $Y2=0
cc_880 N_SET_B_c_1103_n N_A_2006_125#_c_1538_n 0.0236052f $X=12.095 $Y=2.035
+ $X2=0 $Y2=0
cc_881 N_SET_B_c_1103_n N_VPWR_M1010_d 0.00304251f $X=12.095 $Y=2.035 $X2=0
+ $Y2=0
cc_882 N_SET_B_c_1117_n N_VPWR_M1010_d 0.00158531f $X=9.025 $Y=2.035 $X2=0 $Y2=0
cc_883 N_SET_B_c_1098_n N_VPWR_M1010_d 0.00352445f $X=8.935 $Y=1.77 $X2=0 $Y2=0
cc_884 N_SET_B_c_1103_n N_VPWR_M1033_d 0.00448682f $X=12.095 $Y=2.035 $X2=0
+ $Y2=0
cc_885 SET_B N_VPWR_M1033_d 8.48526e-19 $X=12.155 $Y=1.95 $X2=0 $Y2=0
cc_886 N_SET_B_M1010_g N_VPWR_c_1770_n 0.0106736f $X=8.69 $Y=2.595 $X2=0 $Y2=0
cc_887 N_SET_B_M1021_g N_VPWR_c_1771_n 0.00732292f $X=12.225 $Y=2.595 $X2=0
+ $Y2=0
cc_888 N_SET_B_M1010_g N_VPWR_c_1780_n 0.00641304f $X=8.69 $Y=2.595 $X2=0 $Y2=0
cc_889 N_SET_B_M1021_g N_VPWR_c_1782_n 0.00938036f $X=12.225 $Y=2.595 $X2=0
+ $Y2=0
cc_890 N_SET_B_M1010_g N_VPWR_c_1765_n 0.00717129f $X=8.69 $Y=2.595 $X2=0 $Y2=0
cc_891 N_SET_B_M1021_g N_VPWR_c_1765_n 0.0113389f $X=12.225 $Y=2.595 $X2=0 $Y2=0
cc_892 N_SET_B_c_1103_n A_1928_419# 0.00218517f $X=12.095 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_893 N_SET_B_c_1103_n A_2206_419# 0.00172233f $X=12.095 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_894 N_SET_B_M1014_g N_VGND_c_2207_n 0.00171181f $X=8.995 $Y=0.835 $X2=0 $Y2=0
cc_895 N_SET_B_c_1094_n N_VGND_c_2208_n 0.0134773f $X=11.325 $Y=0.825 $X2=0
+ $Y2=0
cc_896 N_SET_B_c_1095_n N_VGND_c_2208_n 0.00941714f $X=12.1 $Y=0.9 $X2=0 $Y2=0
cc_897 N_SET_B_c_1094_n N_VGND_c_2213_n 0.00411131f $X=11.325 $Y=0.825 $X2=0
+ $Y2=0
cc_898 N_SET_B_M1014_g N_VGND_c_2223_n 9.49986e-19 $X=8.995 $Y=0.835 $X2=0 $Y2=0
cc_899 N_SET_B_c_1094_n N_VGND_c_2223_n 0.00781653f $X=11.325 $Y=0.825 $X2=0
+ $Y2=0
cc_900 N_SET_B_c_1095_n N_VGND_c_2223_n 0.0166505f $X=12.1 $Y=0.9 $X2=0 $Y2=0
cc_901 N_A_750_108#_c_1226_n N_A_2172_40#_M1040_g 0.0294613f $X=10.47 $Y=0.18
+ $X2=0 $Y2=0
cc_902 N_A_750_108#_c_1228_n N_A_2172_40#_c_1429_n 0.00424283f $X=10.465 $Y=1.87
+ $X2=0 $Y2=0
cc_903 N_A_750_108#_M1039_g N_A_2172_40#_c_1429_n 0.0294613f $X=10.545 $Y=0.54
+ $X2=0 $Y2=0
cc_904 N_A_750_108#_c_1226_n N_A_2006_125#_c_1523_n 0.00710251f $X=10.47 $Y=0.18
+ $X2=0 $Y2=0
cc_905 N_A_750_108#_M1039_g N_A_2006_125#_c_1523_n 0.0234574f $X=10.545 $Y=0.54
+ $X2=0 $Y2=0
cc_906 N_A_750_108#_M1039_g N_A_2006_125#_c_1524_n 0.00845566f $X=10.545 $Y=0.54
+ $X2=0 $Y2=0
cc_907 N_A_750_108#_M1039_g N_A_2006_125#_c_1525_n 0.00482363f $X=10.545 $Y=0.54
+ $X2=0 $Y2=0
cc_908 N_A_750_108#_c_1233_n N_A_2006_125#_c_1525_n 0.00289117f $X=10.545
+ $Y=1.195 $X2=0 $Y2=0
cc_909 N_A_750_108#_c_1228_n N_A_2006_125#_c_1526_n 0.00220964f $X=10.465
+ $Y=1.87 $X2=0 $Y2=0
cc_910 N_A_750_108#_c_1243_n N_A_2006_125#_c_1538_n 0.018917f $X=10.005 $Y=2.02
+ $X2=0 $Y2=0
cc_911 N_A_750_108#_c_1244_n N_A_2006_125#_c_1538_n 0.0074013f $X=10.39 $Y=1.945
+ $X2=0 $Y2=0
cc_912 N_A_750_108#_c_1249_n N_VPWR_M1002_d 0.00180746f $X=4.825 $Y=2.105 $X2=0
+ $Y2=0
cc_913 N_A_750_108#_M1035_g N_VPWR_c_1768_n 0.0174444f $X=4.805 $Y=2.545 $X2=0
+ $Y2=0
cc_914 N_A_750_108#_c_1247_n N_VPWR_c_1768_n 0.045794f $X=4.01 $Y=2.9 $X2=0
+ $Y2=0
cc_915 N_A_750_108#_c_1249_n N_VPWR_c_1768_n 0.0163515f $X=4.825 $Y=2.105 $X2=0
+ $Y2=0
cc_916 N_A_750_108#_c_1247_n N_VPWR_c_1778_n 0.0220321f $X=4.01 $Y=2.9 $X2=0
+ $Y2=0
cc_917 N_A_750_108#_M1035_g N_VPWR_c_1779_n 0.00767656f $X=4.805 $Y=2.545 $X2=0
+ $Y2=0
cc_918 N_A_750_108#_c_1242_n N_VPWR_c_1779_n 0.00599878f $X=6.73 $Y=2.02 $X2=0
+ $Y2=0
cc_919 N_A_750_108#_c_1243_n N_VPWR_c_1781_n 0.00828633f $X=10.005 $Y=2.02 $X2=0
+ $Y2=0
cc_920 N_A_750_108#_M1035_g N_VPWR_c_1765_n 0.014306f $X=4.805 $Y=2.545 $X2=0
+ $Y2=0
cc_921 N_A_750_108#_c_1242_n N_VPWR_c_1765_n 0.00861531f $X=6.73 $Y=2.02 $X2=0
+ $Y2=0
cc_922 N_A_750_108#_c_1243_n N_VPWR_c_1765_n 0.0132413f $X=10.005 $Y=2.02 $X2=0
+ $Y2=0
cc_923 N_A_750_108#_c_1247_n N_VPWR_c_1765_n 0.0125808f $X=4.01 $Y=2.9 $X2=0
+ $Y2=0
cc_924 N_A_750_108#_c_1247_n N_A_245_406#_c_1934_n 0.00851797f $X=4.01 $Y=2.9
+ $X2=0 $Y2=0
cc_925 N_A_750_108#_c_1234_n N_A_245_406#_c_1934_n 5.64154e-19 $X=3.95 $Y=2.02
+ $X2=0 $Y2=0
cc_926 N_A_750_108#_c_1252_n N_A_245_406#_c_1934_n 0.011925f $X=4.01 $Y=2.105
+ $X2=0 $Y2=0
cc_927 N_A_750_108#_c_1247_n N_A_245_406#_c_1935_n 0.0369449f $X=4.01 $Y=2.9
+ $X2=0 $Y2=0
cc_928 N_A_750_108#_c_1247_n N_A_245_406#_c_1936_n 0.0121616f $X=4.01 $Y=2.9
+ $X2=0 $Y2=0
cc_929 N_A_750_108#_c_1237_n N_A_352_406#_c_1992_n 0.00132047f $X=3.895 $Y=0.795
+ $X2=0 $Y2=0
cc_930 N_A_750_108#_c_1237_n N_A_352_406#_c_1993_n 0.0136369f $X=3.895 $Y=0.795
+ $X2=0 $Y2=0
cc_931 N_A_750_108#_c_1237_n N_A_352_406#_c_1994_n 0.0103474f $X=3.895 $Y=0.795
+ $X2=0 $Y2=0
cc_932 N_A_750_108#_c_1237_n N_A_352_406#_c_1995_n 0.0157629f $X=3.895 $Y=0.795
+ $X2=0 $Y2=0
cc_933 N_A_750_108#_c_1234_n N_A_352_406#_c_1997_n 0.0118074f $X=3.95 $Y=2.02
+ $X2=0 $Y2=0
cc_934 N_A_750_108#_c_1237_n N_A_352_406#_c_1997_n 0.0132237f $X=3.895 $Y=0.795
+ $X2=0 $Y2=0
cc_935 N_A_750_108#_c_1220_n N_A_352_406#_c_1998_n 0.00357582f $X=4.93 $Y=1.555
+ $X2=0 $Y2=0
cc_936 N_A_750_108#_c_1230_n N_A_352_406#_c_1998_n 0.00855772f $X=4.93 $Y=1.195
+ $X2=0 $Y2=0
cc_937 N_A_750_108#_c_1235_n N_A_352_406#_c_1998_n 0.0169523f $X=4.96 $Y=1.72
+ $X2=0 $Y2=0
cc_938 N_A_750_108#_c_1236_n N_A_352_406#_c_1998_n 0.00590221f $X=4.96 $Y=1.72
+ $X2=0 $Y2=0
cc_939 N_A_750_108#_c_1234_n N_A_352_406#_c_2062_n 0.0117724f $X=3.95 $Y=2.02
+ $X2=0 $Y2=0
cc_940 N_A_750_108#_M1031_g N_A_352_406#_c_1999_n 0.0118036f $X=4.93 $Y=0.75
+ $X2=0 $Y2=0
cc_941 N_A_750_108#_c_1221_n N_A_352_406#_c_1999_n 0.00272233f $X=5.215 $Y=1.195
+ $X2=0 $Y2=0
cc_942 N_A_750_108#_M1030_g N_A_352_406#_c_1999_n 0.00526182f $X=5.29 $Y=0.75
+ $X2=0 $Y2=0
cc_943 N_A_750_108#_c_1230_n N_A_352_406#_c_1999_n 7.50555e-19 $X=4.93 $Y=1.195
+ $X2=0 $Y2=0
cc_944 N_A_750_108#_M1030_g N_A_352_406#_c_2000_n 0.00960218f $X=5.29 $Y=0.75
+ $X2=0 $Y2=0
cc_945 N_A_750_108#_c_1223_n N_A_352_406#_c_2000_n 0.00362861f $X=6.205 $Y=1.195
+ $X2=0 $Y2=0
cc_946 N_A_750_108#_M1020_g N_A_352_406#_c_2000_n 0.00858239f $X=6.28 $Y=0.835
+ $X2=0 $Y2=0
cc_947 N_A_750_108#_M1031_g N_A_352_406#_c_2001_n 7.3726e-19 $X=4.93 $Y=0.75
+ $X2=0 $Y2=0
cc_948 N_A_750_108#_M1035_g N_A_352_406#_c_2009_n 0.00452671f $X=4.805 $Y=2.545
+ $X2=0 $Y2=0
cc_949 N_A_750_108#_M1030_g N_A_352_406#_c_2002_n 0.00424696f $X=5.29 $Y=0.75
+ $X2=0 $Y2=0
cc_950 N_A_750_108#_c_1223_n N_A_352_406#_c_2002_n 0.00326111f $X=6.205 $Y=1.195
+ $X2=0 $Y2=0
cc_951 N_A_750_108#_M1020_g N_A_352_406#_c_2002_n 0.00806602f $X=6.28 $Y=0.835
+ $X2=0 $Y2=0
cc_952 N_A_750_108#_c_1220_n N_A_352_406#_c_2004_n 0.00159507f $X=4.93 $Y=1.555
+ $X2=0 $Y2=0
cc_953 N_A_750_108#_c_1221_n N_A_352_406#_c_2004_n 0.00655679f $X=5.215 $Y=1.195
+ $X2=0 $Y2=0
cc_954 N_A_750_108#_c_1223_n N_A_352_406#_c_2004_n 0.00493994f $X=6.205 $Y=1.195
+ $X2=0 $Y2=0
cc_955 N_A_750_108#_c_1231_n N_A_352_406#_c_2004_n 0.00970865f $X=5.29 $Y=1.195
+ $X2=0 $Y2=0
cc_956 N_A_750_108#_c_1236_n N_A_352_406#_c_2004_n 0.00113113f $X=4.96 $Y=1.72
+ $X2=0 $Y2=0
cc_957 N_A_750_108#_M1035_g N_A_352_406#_c_2005_n 0.00151603f $X=4.805 $Y=2.545
+ $X2=0 $Y2=0
cc_958 N_A_750_108#_c_1220_n N_A_352_406#_c_2005_n 0.00602087f $X=4.93 $Y=1.555
+ $X2=0 $Y2=0
cc_959 N_A_750_108#_c_1231_n N_A_352_406#_c_2005_n 0.00139177f $X=5.29 $Y=1.195
+ $X2=0 $Y2=0
cc_960 N_A_750_108#_c_1235_n N_A_352_406#_c_2005_n 0.0334879f $X=4.96 $Y=1.72
+ $X2=0 $Y2=0
cc_961 N_A_750_108#_c_1236_n N_A_352_406#_c_2005_n 0.00336924f $X=4.96 $Y=1.72
+ $X2=0 $Y2=0
cc_962 N_A_750_108#_c_1249_n N_A_352_406#_c_2011_n 0.0146f $X=4.825 $Y=2.105
+ $X2=0 $Y2=0
cc_963 N_A_750_108#_M1031_g N_VGND_c_2205_n 0.0012123f $X=4.93 $Y=0.75 $X2=0
+ $Y2=0
cc_964 N_A_750_108#_c_1226_n N_VGND_c_2206_n 0.0210695f $X=10.47 $Y=0.18 $X2=0
+ $Y2=0
cc_965 N_A_750_108#_c_1226_n N_VGND_c_2207_n 0.0261591f $X=10.47 $Y=0.18 $X2=0
+ $Y2=0
cc_966 N_A_750_108#_c_1226_n N_VGND_c_2213_n 0.0369976f $X=10.47 $Y=0.18 $X2=0
+ $Y2=0
cc_967 N_A_750_108#_M1031_g N_VGND_c_2219_n 0.00423267f $X=4.93 $Y=0.75 $X2=0
+ $Y2=0
cc_968 N_A_750_108#_M1030_g N_VGND_c_2219_n 6.5362e-19 $X=5.29 $Y=0.75 $X2=0
+ $Y2=0
cc_969 N_A_750_108#_c_1227_n N_VGND_c_2219_n 0.0364304f $X=6.355 $Y=0.18 $X2=0
+ $Y2=0
cc_970 N_A_750_108#_c_1226_n N_VGND_c_2220_n 0.0361813f $X=10.47 $Y=0.18 $X2=0
+ $Y2=0
cc_971 N_A_750_108#_M1031_g N_VGND_c_2223_n 0.00444208f $X=4.93 $Y=0.75 $X2=0
+ $Y2=0
cc_972 N_A_750_108#_c_1226_n N_VGND_c_2223_n 0.12596f $X=10.47 $Y=0.18 $X2=0
+ $Y2=0
cc_973 N_A_750_108#_c_1227_n N_VGND_c_2223_n 0.0116041f $X=6.355 $Y=0.18 $X2=0
+ $Y2=0
cc_974 N_A_2172_40#_c_1433_n N_A_2006_125#_c_1510_n 0.0126504f $X=12.63 $Y=0.495
+ $X2=0 $Y2=0
cc_975 N_A_2172_40#_c_1434_n N_A_2006_125#_c_1511_n 0.0135802f $X=13.01 $Y=1.085
+ $X2=0 $Y2=0
cc_976 N_A_2172_40#_c_1433_n N_A_2006_125#_c_1512_n 0.005422f $X=12.63 $Y=0.495
+ $X2=0 $Y2=0
cc_977 N_A_2172_40#_c_1434_n N_A_2006_125#_c_1512_n 0.0097739f $X=13.01 $Y=1.085
+ $X2=0 $Y2=0
cc_978 N_A_2172_40#_c_1435_n N_A_2006_125#_c_1512_n 0.00151451f $X=13.05 $Y=1.88
+ $X2=0 $Y2=0
cc_979 N_A_2172_40#_c_1433_n N_A_2006_125#_c_1513_n 0.00174859f $X=12.63
+ $Y=0.495 $X2=0 $Y2=0
cc_980 N_A_2172_40#_c_1434_n N_A_2006_125#_c_1519_n 0.00112993f $X=13.01
+ $Y=1.085 $X2=0 $Y2=0
cc_981 N_A_2172_40#_M1040_g N_A_2006_125#_c_1523_n 0.0031992f $X=10.935 $Y=0.54
+ $X2=0 $Y2=0
cc_982 N_A_2172_40#_M1040_g N_A_2006_125#_c_1524_n 0.0160271f $X=10.935 $Y=0.54
+ $X2=0 $Y2=0
cc_983 N_A_2172_40#_c_1428_n N_A_2006_125#_c_1524_n 0.00742319f $X=11.32 $Y=1.29
+ $X2=0 $Y2=0
cc_984 N_A_2172_40#_c_1432_n N_A_2006_125#_c_1524_n 0.0147436f $X=11.89 $Y=1
+ $X2=0 $Y2=0
cc_985 N_A_2172_40#_M1040_g N_A_2006_125#_c_1526_n 0.00416286f $X=10.935 $Y=0.54
+ $X2=0 $Y2=0
cc_986 N_A_2172_40#_c_1428_n N_A_2006_125#_c_1526_n 0.0071263f $X=11.32 $Y=1.29
+ $X2=0 $Y2=0
cc_987 N_A_2172_40#_M1033_g N_A_2006_125#_c_1526_n 0.014639f $X=11.445 $Y=2.595
+ $X2=0 $Y2=0
cc_988 N_A_2172_40#_c_1430_n N_A_2006_125#_c_1526_n 0.0551777f $X=11.725 $Y=1.38
+ $X2=0 $Y2=0
cc_989 N_A_2172_40#_c_1436_n N_A_2006_125#_c_1526_n 0.0204573f $X=11.605 $Y=1.29
+ $X2=0 $Y2=0
cc_990 N_A_2172_40#_M1033_g N_A_2006_125#_c_1565_n 0.0120516f $X=11.445 $Y=2.595
+ $X2=0 $Y2=0
cc_991 N_A_2172_40#_c_1430_n N_A_2006_125#_c_1565_n 0.00493162f $X=11.725
+ $Y=1.38 $X2=0 $Y2=0
cc_992 N_A_2172_40#_c_1436_n N_A_2006_125#_c_1565_n 0.00157019f $X=11.605
+ $Y=1.29 $X2=0 $Y2=0
cc_993 N_A_2172_40#_c_1435_n N_A_2006_125#_c_1533_n 0.011925f $X=13.05 $Y=1.88
+ $X2=0 $Y2=0
cc_994 N_A_2172_40#_c_1435_n N_A_2006_125#_c_1534_n 0.0141629f $X=13.05 $Y=1.88
+ $X2=0 $Y2=0
cc_995 N_A_2172_40#_c_1435_n N_A_2006_125#_c_1535_n 0.0183398f $X=13.05 $Y=1.88
+ $X2=0 $Y2=0
cc_996 N_A_2172_40#_c_1433_n N_A_2006_125#_c_1606_n 3.00845e-19 $X=12.63
+ $Y=0.495 $X2=0 $Y2=0
cc_997 N_A_2172_40#_c_1434_n N_A_2006_125#_c_1606_n 0.0132649f $X=13.01 $Y=1.085
+ $X2=0 $Y2=0
cc_998 N_A_2172_40#_c_1435_n N_A_2006_125#_c_1606_n 0.0792281f $X=13.05 $Y=1.88
+ $X2=0 $Y2=0
cc_999 N_A_2172_40#_c_1434_n N_A_2006_125#_c_1527_n 0.00311101f $X=13.01
+ $Y=1.085 $X2=0 $Y2=0
cc_1000 N_A_2172_40#_c_1435_n N_A_2006_125#_c_1527_n 0.0239983f $X=13.05 $Y=1.88
+ $X2=0 $Y2=0
cc_1001 N_A_2172_40#_M1033_g N_A_2006_125#_c_1611_n 0.00577012f $X=11.445
+ $Y=2.595 $X2=0 $Y2=0
cc_1002 N_A_2172_40#_M1033_g N_VPWR_c_1771_n 0.0146179f $X=11.445 $Y=2.595 $X2=0
+ $Y2=0
cc_1003 N_A_2172_40#_M1033_g N_VPWR_c_1781_n 0.008763f $X=11.445 $Y=2.595 $X2=0
+ $Y2=0
cc_1004 N_A_2172_40#_M1033_g N_VPWR_c_1765_n 0.00785204f $X=11.445 $Y=2.595
+ $X2=0 $Y2=0
cc_1005 N_A_2172_40#_M1040_g N_VGND_c_2208_n 0.00279447f $X=10.935 $Y=0.54 $X2=0
+ $Y2=0
cc_1006 N_A_2172_40#_c_1432_n N_VGND_c_2208_n 0.00998028f $X=11.89 $Y=1 $X2=0
+ $Y2=0
cc_1007 N_A_2172_40#_c_1433_n N_VGND_c_2209_n 0.0153904f $X=12.63 $Y=0.495 $X2=0
+ $Y2=0
cc_1008 N_A_2172_40#_M1040_g N_VGND_c_2213_n 0.00495161f $X=10.935 $Y=0.54 $X2=0
+ $Y2=0
cc_1009 N_A_2172_40#_c_1433_n N_VGND_c_2215_n 0.0219574f $X=12.63 $Y=0.495 $X2=0
+ $Y2=0
cc_1010 N_A_2172_40#_M1040_g N_VGND_c_2223_n 0.0097634f $X=10.935 $Y=0.54 $X2=0
+ $Y2=0
cc_1011 N_A_2172_40#_c_1433_n N_VGND_c_2223_n 0.0125652f $X=12.63 $Y=0.495 $X2=0
+ $Y2=0
cc_1012 N_A_2006_125#_M1012_g N_A_2767_57#_M1032_g 0.0395279f $X=14.555 $Y=0.495
+ $X2=0 $Y2=0
cc_1013 N_A_2006_125#_M1003_g N_A_2767_57#_M1037_g 0.0163172f $X=14.575 $Y=2.37
+ $X2=0 $Y2=0
cc_1014 N_A_2006_125#_M1003_g N_A_2767_57#_c_1694_n 0.00766063f $X=14.575
+ $Y=2.37 $X2=0 $Y2=0
cc_1015 N_A_2006_125#_M1027_g N_A_2767_57#_c_1695_n 0.010329f $X=14.195 $Y=0.495
+ $X2=0 $Y2=0
cc_1016 N_A_2006_125#_M1012_g N_A_2767_57#_c_1695_n 0.00175877f $X=14.555
+ $Y=0.495 $X2=0 $Y2=0
cc_1017 N_A_2006_125#_c_1519_n N_A_2767_57#_c_1695_n 0.00204063f $X=13.387
+ $Y=0.9 $X2=0 $Y2=0
cc_1018 N_A_2006_125#_c_1606_n N_A_2767_57#_c_1695_n 0.00304483f $X=13.48
+ $Y=1.07 $X2=0 $Y2=0
cc_1019 N_A_2006_125#_M1015_g N_A_2767_57#_c_1696_n 0.00225207f $X=13.315
+ $Y=2.235 $X2=0 $Y2=0
cc_1020 N_A_2006_125#_c_1514_n N_A_2767_57#_c_1696_n 0.00453915f $X=14.12 $Y=1.5
+ $X2=0 $Y2=0
cc_1021 N_A_2006_125#_M1027_g N_A_2767_57#_c_1696_n 0.00748594f $X=14.195
+ $Y=0.495 $X2=0 $Y2=0
cc_1022 N_A_2006_125#_c_1516_n N_A_2767_57#_c_1696_n 0.00540806f $X=14.45 $Y=1.5
+ $X2=0 $Y2=0
cc_1023 N_A_2006_125#_M1003_g N_A_2767_57#_c_1696_n 0.0297615f $X=14.575 $Y=2.37
+ $X2=0 $Y2=0
cc_1024 N_A_2006_125#_M1012_g N_A_2767_57#_c_1696_n 0.00317353f $X=14.555
+ $Y=0.495 $X2=0 $Y2=0
cc_1025 N_A_2006_125#_c_1521_n N_A_2767_57#_c_1696_n 0.00588934f $X=14.195
+ $Y=1.5 $X2=0 $Y2=0
cc_1026 N_A_2006_125#_c_1522_n N_A_2767_57#_c_1696_n 0.00269777f $X=14.575
+ $Y=1.5 $X2=0 $Y2=0
cc_1027 N_A_2006_125#_c_1606_n N_A_2767_57#_c_1696_n 0.0153809f $X=13.48 $Y=1.07
+ $X2=0 $Y2=0
cc_1028 N_A_2006_125#_c_1527_n N_A_2767_57#_c_1696_n 0.00208619f $X=13.48
+ $Y=1.07 $X2=0 $Y2=0
cc_1029 N_A_2006_125#_c_1537_n N_A_2767_57#_c_1696_n 0.00559149f $X=13.4
+ $Y=2.895 $X2=0 $Y2=0
cc_1030 N_A_2006_125#_M1012_g N_A_2767_57#_c_1697_n 0.0184611f $X=14.555
+ $Y=0.495 $X2=0 $Y2=0
cc_1031 N_A_2006_125#_c_1522_n N_A_2767_57#_c_1697_n 0.00262418f $X=14.575
+ $Y=1.5 $X2=0 $Y2=0
cc_1032 N_A_2006_125#_c_1513_n N_A_2767_57#_c_1698_n 0.00100153f $X=13.205
+ $Y=0.825 $X2=0 $Y2=0
cc_1033 N_A_2006_125#_M1027_g N_A_2767_57#_c_1698_n 0.0128629f $X=14.195
+ $Y=0.495 $X2=0 $Y2=0
cc_1034 N_A_2006_125#_M1012_g N_A_2767_57#_c_1698_n 0.00151759f $X=14.555
+ $Y=0.495 $X2=0 $Y2=0
cc_1035 N_A_2006_125#_M1027_g N_A_2767_57#_c_1699_n 0.005487f $X=14.195 $Y=0.495
+ $X2=0 $Y2=0
cc_1036 N_A_2006_125#_c_1606_n N_A_2767_57#_c_1699_n 0.00693741f $X=13.48
+ $Y=1.07 $X2=0 $Y2=0
cc_1037 N_A_2006_125#_c_1527_n N_A_2767_57#_c_1699_n 0.00144622f $X=13.48
+ $Y=1.07 $X2=0 $Y2=0
cc_1038 N_A_2006_125#_M1012_g N_A_2767_57#_c_1700_n 9.65688e-19 $X=14.555
+ $Y=0.495 $X2=0 $Y2=0
cc_1039 N_A_2006_125#_c_1522_n N_A_2767_57#_c_1700_n 0.00101735f $X=14.575
+ $Y=1.5 $X2=0 $Y2=0
cc_1040 N_A_2006_125#_c_1522_n N_A_2767_57#_c_1701_n 0.00766063f $X=14.575
+ $Y=1.5 $X2=0 $Y2=0
cc_1041 N_A_2006_125#_c_1565_n N_VPWR_M1033_d 0.0129524f $X=12.325 $Y=2.415
+ $X2=0 $Y2=0
cc_1042 N_A_2006_125#_c_1565_n N_VPWR_c_1771_n 0.0197154f $X=12.325 $Y=2.415
+ $X2=0 $Y2=0
cc_1043 N_A_2006_125#_c_1534_n N_VPWR_c_1771_n 0.00784614f $X=12.49 $Y=2.895
+ $X2=0 $Y2=0
cc_1044 N_A_2006_125#_c_1536_n N_VPWR_c_1771_n 0.00656934f $X=12.655 $Y=2.98
+ $X2=0 $Y2=0
cc_1045 N_A_2006_125#_M1015_g N_VPWR_c_1772_n 0.00710853f $X=13.315 $Y=2.235
+ $X2=0 $Y2=0
cc_1046 N_A_2006_125#_c_1514_n N_VPWR_c_1772_n 0.0105821f $X=14.12 $Y=1.5 $X2=0
+ $Y2=0
cc_1047 N_A_2006_125#_M1003_g N_VPWR_c_1772_n 0.00461224f $X=14.575 $Y=2.37
+ $X2=0 $Y2=0
cc_1048 N_A_2006_125#_c_1535_n N_VPWR_c_1772_n 0.0141601f $X=13.315 $Y=2.98
+ $X2=0 $Y2=0
cc_1049 N_A_2006_125#_c_1537_n N_VPWR_c_1772_n 0.0479842f $X=13.4 $Y=2.895 $X2=0
+ $Y2=0
cc_1050 N_A_2006_125#_M1003_g N_VPWR_c_1773_n 0.0265364f $X=14.575 $Y=2.37 $X2=0
+ $Y2=0
cc_1051 N_A_2006_125#_M1003_g N_VPWR_c_1776_n 0.00747382f $X=14.575 $Y=2.37
+ $X2=0 $Y2=0
cc_1052 N_A_2006_125#_c_1541_n N_VPWR_c_1781_n 0.0216692f $X=10.405 $Y=2.9 $X2=0
+ $Y2=0
cc_1053 N_A_2006_125#_M1015_g N_VPWR_c_1782_n 6.29517e-19 $X=13.315 $Y=2.235
+ $X2=0 $Y2=0
cc_1054 N_A_2006_125#_c_1535_n N_VPWR_c_1782_n 0.0514264f $X=13.315 $Y=2.98
+ $X2=0 $Y2=0
cc_1055 N_A_2006_125#_c_1536_n N_VPWR_c_1782_n 0.0198894f $X=12.655 $Y=2.98
+ $X2=0 $Y2=0
cc_1056 N_A_2006_125#_M1011_d N_VPWR_c_1765_n 0.0105425f $X=10.13 $Y=2.095 $X2=0
+ $Y2=0
cc_1057 N_A_2006_125#_M1021_d N_VPWR_c_1765_n 0.0023218f $X=12.35 $Y=2.095 $X2=0
+ $Y2=0
cc_1058 N_A_2006_125#_M1003_g N_VPWR_c_1765_n 0.00779694f $X=14.575 $Y=2.37
+ $X2=0 $Y2=0
cc_1059 N_A_2006_125#_c_1541_n N_VPWR_c_1765_n 0.0126914f $X=10.405 $Y=2.9 $X2=0
+ $Y2=0
cc_1060 N_A_2006_125#_c_1548_n N_VPWR_c_1765_n 0.0213707f $X=11.235 $Y=2.415
+ $X2=0 $Y2=0
cc_1061 N_A_2006_125#_c_1565_n N_VPWR_c_1765_n 0.0190568f $X=12.325 $Y=2.415
+ $X2=0 $Y2=0
cc_1062 N_A_2006_125#_c_1535_n N_VPWR_c_1765_n 0.0312358f $X=13.315 $Y=2.98
+ $X2=0 $Y2=0
cc_1063 N_A_2006_125#_c_1536_n N_VPWR_c_1765_n 0.0125808f $X=12.655 $Y=2.98
+ $X2=0 $Y2=0
cc_1064 N_A_2006_125#_c_1611_n N_VPWR_c_1765_n 0.00606883f $X=11.32 $Y=2.415
+ $X2=0 $Y2=0
cc_1065 N_A_2006_125#_c_1548_n A_2206_419# 0.00494602f $X=11.235 $Y=2.415
+ $X2=-0.19 $Y2=-0.245
cc_1066 N_A_2006_125#_c_1526_n A_2206_419# 0.00331016f $X=11.32 $Y=2.33
+ $X2=-0.19 $Y2=-0.245
cc_1067 N_A_2006_125#_c_1611_n A_2206_419# 6.35756e-19 $X=11.32 $Y=2.415
+ $X2=-0.19 $Y2=-0.245
cc_1068 N_A_2006_125#_M1003_g N_Q_c_2185_n 2.75707e-19 $X=14.575 $Y=2.37 $X2=0
+ $Y2=0
cc_1069 N_A_2006_125#_c_1523_n N_VGND_c_2207_n 0.014278f $X=10.25 $Y=0.475 $X2=0
+ $Y2=0
cc_1070 N_A_2006_125#_c_1525_n N_VGND_c_2207_n 0.0024802f $X=10.53 $Y=1 $X2=0
+ $Y2=0
cc_1071 N_A_2006_125#_c_1524_n N_VGND_c_2208_n 0.00210116f $X=11.235 $Y=1 $X2=0
+ $Y2=0
cc_1072 N_A_2006_125#_c_1510_n N_VGND_c_2209_n 0.002112f $X=12.845 $Y=0.825
+ $X2=0 $Y2=0
cc_1073 N_A_2006_125#_c_1513_n N_VGND_c_2209_n 0.0149349f $X=13.205 $Y=0.825
+ $X2=0 $Y2=0
cc_1074 N_A_2006_125#_M1027_g N_VGND_c_2209_n 0.00281003f $X=14.195 $Y=0.495
+ $X2=0 $Y2=0
cc_1075 N_A_2006_125#_c_1519_n N_VGND_c_2209_n 0.00986306f $X=13.387 $Y=0.9
+ $X2=0 $Y2=0
cc_1076 N_A_2006_125#_c_1606_n N_VGND_c_2209_n 0.0228655f $X=13.48 $Y=1.07 $X2=0
+ $Y2=0
cc_1077 N_A_2006_125#_M1027_g N_VGND_c_2210_n 0.00202687f $X=14.195 $Y=0.495
+ $X2=0 $Y2=0
cc_1078 N_A_2006_125#_M1012_g N_VGND_c_2210_n 0.0115615f $X=14.555 $Y=0.495
+ $X2=0 $Y2=0
cc_1079 N_A_2006_125#_c_1523_n N_VGND_c_2213_n 0.0233299f $X=10.25 $Y=0.475
+ $X2=0 $Y2=0
cc_1080 N_A_2006_125#_c_1510_n N_VGND_c_2215_n 0.00502664f $X=12.845 $Y=0.825
+ $X2=0 $Y2=0
cc_1081 N_A_2006_125#_c_1513_n N_VGND_c_2215_n 0.00445056f $X=13.205 $Y=0.825
+ $X2=0 $Y2=0
cc_1082 N_A_2006_125#_M1027_g N_VGND_c_2221_n 0.00334669f $X=14.195 $Y=0.495
+ $X2=0 $Y2=0
cc_1083 N_A_2006_125#_M1012_g N_VGND_c_2221_n 0.00445056f $X=14.555 $Y=0.495
+ $X2=0 $Y2=0
cc_1084 N_A_2006_125#_c_1510_n N_VGND_c_2223_n 0.010303f $X=12.845 $Y=0.825
+ $X2=0 $Y2=0
cc_1085 N_A_2006_125#_c_1511_n N_VGND_c_2223_n 6.16811e-19 $X=13.13 $Y=0.9 $X2=0
+ $Y2=0
cc_1086 N_A_2006_125#_c_1513_n N_VGND_c_2223_n 0.00796275f $X=13.205 $Y=0.825
+ $X2=0 $Y2=0
cc_1087 N_A_2006_125#_M1027_g N_VGND_c_2223_n 0.00581109f $X=14.195 $Y=0.495
+ $X2=0 $Y2=0
cc_1088 N_A_2006_125#_M1012_g N_VGND_c_2223_n 0.00796275f $X=14.555 $Y=0.495
+ $X2=0 $Y2=0
cc_1089 N_A_2006_125#_c_1519_n N_VGND_c_2223_n 0.00157435f $X=13.387 $Y=0.9
+ $X2=0 $Y2=0
cc_1090 N_A_2006_125#_c_1523_n N_VGND_c_2223_n 0.0149002f $X=10.25 $Y=0.475
+ $X2=0 $Y2=0
cc_1091 N_A_2767_57#_c_1696_n N_VPWR_c_1772_n 0.0898892f $X=14.31 $Y=2.015 $X2=0
+ $Y2=0
cc_1092 N_A_2767_57#_M1037_g N_VPWR_c_1773_n 0.0257478f $X=15.105 $Y=2.37 $X2=0
+ $Y2=0
cc_1093 N_A_2767_57#_c_1694_n N_VPWR_c_1773_n 5.32278e-19 $X=15.075 $Y=1.66
+ $X2=0 $Y2=0
cc_1094 N_A_2767_57#_c_1696_n N_VPWR_c_1773_n 0.0692741f $X=14.31 $Y=2.015 $X2=0
+ $Y2=0
cc_1095 N_A_2767_57#_c_1700_n N_VPWR_c_1773_n 0.00750214f $X=15.075 $Y=1.155
+ $X2=0 $Y2=0
cc_1096 N_A_2767_57#_c_1696_n N_VPWR_c_1776_n 0.0122968f $X=14.31 $Y=2.015 $X2=0
+ $Y2=0
cc_1097 N_A_2767_57#_M1037_g N_VPWR_c_1783_n 0.00747382f $X=15.105 $Y=2.37 $X2=0
+ $Y2=0
cc_1098 N_A_2767_57#_M1037_g N_VPWR_c_1765_n 0.00779694f $X=15.105 $Y=2.37 $X2=0
+ $Y2=0
cc_1099 N_A_2767_57#_c_1696_n N_VPWR_c_1765_n 0.0131561f $X=14.31 $Y=2.015 $X2=0
+ $Y2=0
cc_1100 N_A_2767_57#_M1032_g N_Q_c_2181_n 0.00125204f $X=14.985 $Y=0.495 $X2=0
+ $Y2=0
cc_1101 N_A_2767_57#_M1026_g N_Q_c_2181_n 0.0100348f $X=15.345 $Y=0.495 $X2=0
+ $Y2=0
cc_1102 N_A_2767_57#_M1037_g Q 0.00651453f $X=15.105 $Y=2.37 $X2=0 $Y2=0
cc_1103 N_A_2767_57#_M1026_g Q 0.014928f $X=15.345 $Y=0.495 $X2=0 $Y2=0
cc_1104 N_A_2767_57#_c_1700_n Q 0.0398637f $X=15.075 $Y=1.155 $X2=0 $Y2=0
cc_1105 N_A_2767_57#_c_1701_n Q 0.0108771f $X=15.075 $Y=1.155 $X2=0 $Y2=0
cc_1106 N_A_2767_57#_M1037_g Q 0.0139894f $X=15.105 $Y=2.37 $X2=0 $Y2=0
cc_1107 N_A_2767_57#_M1037_g N_Q_c_2185_n 0.00522616f $X=15.105 $Y=2.37 $X2=0
+ $Y2=0
cc_1108 N_A_2767_57#_c_1700_n N_Q_c_2185_n 0.00259106f $X=15.075 $Y=1.155 $X2=0
+ $Y2=0
cc_1109 N_A_2767_57#_c_1698_n N_VGND_c_2209_n 0.0317249f $X=14.18 $Y=0.495 $X2=0
+ $Y2=0
cc_1110 N_A_2767_57#_M1032_g N_VGND_c_2210_n 0.012605f $X=14.985 $Y=0.495 $X2=0
+ $Y2=0
cc_1111 N_A_2767_57#_M1026_g N_VGND_c_2210_n 0.002112f $X=15.345 $Y=0.495 $X2=0
+ $Y2=0
cc_1112 N_A_2767_57#_c_1697_n N_VGND_c_2210_n 0.0185923f $X=14.91 $Y=1.075 $X2=0
+ $Y2=0
cc_1113 N_A_2767_57#_c_1698_n N_VGND_c_2210_n 0.0202525f $X=14.18 $Y=0.495 $X2=0
+ $Y2=0
cc_1114 N_A_2767_57#_c_1700_n N_VGND_c_2210_n 0.00141855f $X=15.075 $Y=1.155
+ $X2=0 $Y2=0
cc_1115 N_A_2767_57#_c_1698_n N_VGND_c_2221_n 0.0288109f $X=14.18 $Y=0.495 $X2=0
+ $Y2=0
cc_1116 N_A_2767_57#_M1032_g N_VGND_c_2222_n 0.00445056f $X=14.985 $Y=0.495
+ $X2=0 $Y2=0
cc_1117 N_A_2767_57#_M1026_g N_VGND_c_2222_n 0.00502664f $X=15.345 $Y=0.495
+ $X2=0 $Y2=0
cc_1118 N_A_2767_57#_M1032_g N_VGND_c_2223_n 0.00796275f $X=14.985 $Y=0.495
+ $X2=0 $Y2=0
cc_1119 N_A_2767_57#_M1026_g N_VGND_c_2223_n 0.0100616f $X=15.345 $Y=0.495 $X2=0
+ $Y2=0
cc_1120 N_A_2767_57#_c_1698_n N_VGND_c_2223_n 0.016554f $X=14.18 $Y=0.495 $X2=0
+ $Y2=0
cc_1121 N_VPWR_c_1766_n N_A_245_406#_c_1931_n 0.0586203f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_1122 N_VPWR_c_1767_n N_A_245_406#_c_1932_n 0.00830303f $X=2.92 $Y=2.86 $X2=0
+ $Y2=0
cc_1123 N_VPWR_c_1774_n N_A_245_406#_c_1932_n 0.0530763f $X=2.755 $Y=3.33 $X2=0
+ $Y2=0
cc_1124 N_VPWR_c_1765_n N_A_245_406#_c_1932_n 0.0309297f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1125 N_VPWR_c_1766_n N_A_245_406#_c_1933_n 0.0121616f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_1126 N_VPWR_c_1774_n N_A_245_406#_c_1933_n 0.0221635f $X=2.755 $Y=3.33 $X2=0
+ $Y2=0
cc_1127 N_VPWR_c_1765_n N_A_245_406#_c_1933_n 0.0126536f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1128 N_VPWR_c_1767_n N_A_245_406#_c_1940_n 0.00972699f $X=2.92 $Y=2.86 $X2=0
+ $Y2=0
cc_1129 N_VPWR_M1018_d N_A_245_406#_c_1941_n 0.00356107f $X=2.78 $Y=2.03 $X2=0
+ $Y2=0
cc_1130 N_VPWR_c_1767_n N_A_245_406#_c_1941_n 0.0159264f $X=2.92 $Y=2.86 $X2=0
+ $Y2=0
cc_1131 N_VPWR_c_1765_n N_A_245_406#_c_1941_n 0.0192581f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1132 N_VPWR_c_1767_n N_A_245_406#_c_1935_n 0.0101047f $X=2.92 $Y=2.86 $X2=0
+ $Y2=0
cc_1133 N_VPWR_c_1778_n N_A_245_406#_c_1935_n 0.0153477f $X=4.375 $Y=3.33 $X2=0
+ $Y2=0
cc_1134 N_VPWR_c_1765_n N_A_245_406#_c_1935_n 0.00952457f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1135 N_VPWR_c_1765_n N_A_352_406#_M1019_s 0.00224633f $X=15.6 $Y=3.33 $X2=0
+ $Y2=0
cc_1136 N_VPWR_M1018_d N_A_352_406#_c_2006_n 0.00181172f $X=2.78 $Y=2.03 $X2=0
+ $Y2=0
cc_1137 N_VPWR_c_1765_n A_1371_419# 0.00285375f $X=15.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1138 N_VPWR_c_1765_n A_1928_419# 0.00286f $X=15.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1139 N_VPWR_c_1765_n A_2206_419# 0.00421098f $X=15.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1140 N_VPWR_c_1783_n Q 0.0168747f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1141 N_VPWR_c_1765_n Q 0.0180375f $X=15.6 $Y=3.33 $X2=0 $Y2=0
cc_1142 N_VPWR_c_1773_n N_Q_c_2185_n 0.0709584f $X=14.84 $Y=2.015 $X2=0 $Y2=0
cc_1143 N_A_245_406#_c_1932_n N_A_352_406#_M1016_d 0.00180746f $X=2.245 $Y=2.98
+ $X2=0 $Y2=0
cc_1144 N_A_245_406#_c_1931_n N_A_352_406#_c_2012_n 0.0378542f $X=1.37 $Y=2.175
+ $X2=0 $Y2=0
cc_1145 N_A_245_406#_c_1932_n N_A_352_406#_c_2012_n 0.015238f $X=2.245 $Y=2.98
+ $X2=0 $Y2=0
cc_1146 N_A_245_406#_c_1940_n N_A_352_406#_c_2012_n 0.0153156f $X=2.33 $Y=2.895
+ $X2=0 $Y2=0
cc_1147 N_A_245_406#_c_1951_n N_A_352_406#_c_2012_n 0.0129587f $X=2.415 $Y=2.405
+ $X2=0 $Y2=0
cc_1148 N_A_245_406#_c_1941_n N_A_352_406#_c_2006_n 0.0407967f $X=3.365 $Y=2.405
+ $X2=0 $Y2=0
cc_1149 N_A_245_406#_c_1951_n N_A_352_406#_c_2006_n 0.00857425f $X=2.415
+ $Y=2.405 $X2=0 $Y2=0
cc_1150 N_A_245_406#_c_1934_n N_A_352_406#_c_2006_n 0.0059602f $X=3.45 $Y=2.175
+ $X2=0 $Y2=0
cc_1151 N_A_245_406#_c_1931_n N_A_352_406#_c_2007_n 0.0091047f $X=1.37 $Y=2.175
+ $X2=0 $Y2=0
cc_1152 N_A_245_406#_c_1932_n A_458_406# 0.00154159f $X=2.245 $Y=2.98 $X2=-0.19
+ $Y2=1.655
cc_1153 N_A_245_406#_c_1940_n A_458_406# 0.00445973f $X=2.33 $Y=2.895 $X2=-0.19
+ $Y2=1.655
cc_1154 N_A_245_406#_c_1941_n A_458_406# 0.00176808f $X=3.365 $Y=2.405 $X2=-0.19
+ $Y2=1.655
cc_1155 N_A_245_406#_c_1951_n A_458_406# 7.72785e-19 $X=2.415 $Y=2.405 $X2=-0.19
+ $Y2=1.655
cc_1156 N_A_352_406#_c_2006_n A_458_406# 0.00137342f $X=3.015 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_1157 N_A_352_406#_c_1993_n N_VGND_c_2204_n 0.00668062f $X=3.455 $Y=0.845
+ $X2=0 $Y2=0
cc_1158 N_A_352_406#_c_1994_n N_VGND_c_2204_n 0.0105542f $X=3.54 $Y=0.76 $X2=0
+ $Y2=0
cc_1159 N_A_352_406#_c_1996_n N_VGND_c_2204_n 0.0139102f $X=3.625 $Y=0.35 $X2=0
+ $Y2=0
cc_1160 N_A_352_406#_c_2003_n N_VGND_c_2204_n 0.0118667f $X=2.37 $Y=0.445 $X2=0
+ $Y2=0
cc_1161 N_A_352_406#_c_2051_n N_VGND_c_2204_n 0.0102206f $X=3.1 $Y=0.845 $X2=0
+ $Y2=0
cc_1162 N_A_352_406#_c_1995_n N_VGND_c_2205_n 0.0119743f $X=4.24 $Y=0.35 $X2=0
+ $Y2=0
cc_1163 N_A_352_406#_c_1997_n N_VGND_c_2205_n 0.00769201f $X=4.325 $Y=1.16 $X2=0
+ $Y2=0
cc_1164 N_A_352_406#_c_1998_n N_VGND_c_2205_n 0.0136256f $X=4.99 $Y=1.245 $X2=0
+ $Y2=0
cc_1165 N_A_352_406#_c_1999_n N_VGND_c_2205_n 0.0211433f $X=5.075 $Y=1.16 $X2=0
+ $Y2=0
cc_1166 N_A_352_406#_c_2001_n N_VGND_c_2205_n 0.0131556f $X=5.16 $Y=0.35 $X2=0
+ $Y2=0
cc_1167 N_A_352_406#_c_1993_n N_VGND_c_2211_n 0.00254764f $X=3.455 $Y=0.845
+ $X2=0 $Y2=0
cc_1168 N_A_352_406#_c_1995_n N_VGND_c_2211_n 0.0486978f $X=4.24 $Y=0.35 $X2=0
+ $Y2=0
cc_1169 N_A_352_406#_c_1996_n N_VGND_c_2211_n 0.0114429f $X=3.625 $Y=0.35 $X2=0
+ $Y2=0
cc_1170 N_A_352_406#_c_1991_n N_VGND_c_2218_n 0.0052665f $X=3.015 $Y=0.845 $X2=0
+ $Y2=0
cc_1171 N_A_352_406#_c_2003_n N_VGND_c_2218_n 0.0231253f $X=2.37 $Y=0.445 $X2=0
+ $Y2=0
cc_1172 N_A_352_406#_c_2000_n N_VGND_c_2219_n 0.0611279f $X=5.98 $Y=0.35 $X2=0
+ $Y2=0
cc_1173 N_A_352_406#_c_2001_n N_VGND_c_2219_n 0.0114622f $X=5.16 $Y=0.35 $X2=0
+ $Y2=0
cc_1174 N_A_352_406#_M1023_d N_VGND_c_2223_n 0.0022543f $X=2.23 $Y=0.235 $X2=0
+ $Y2=0
cc_1175 N_A_352_406#_c_1991_n N_VGND_c_2223_n 0.00935798f $X=3.015 $Y=0.845
+ $X2=0 $Y2=0
cc_1176 N_A_352_406#_c_1993_n N_VGND_c_2223_n 0.00501995f $X=3.455 $Y=0.845
+ $X2=0 $Y2=0
cc_1177 N_A_352_406#_c_1995_n N_VGND_c_2223_n 0.029554f $X=4.24 $Y=0.35 $X2=0
+ $Y2=0
cc_1178 N_A_352_406#_c_1996_n N_VGND_c_2223_n 0.00657383f $X=3.625 $Y=0.35 $X2=0
+ $Y2=0
cc_1179 N_A_352_406#_c_2000_n N_VGND_c_2223_n 0.0372155f $X=5.98 $Y=0.35 $X2=0
+ $Y2=0
cc_1180 N_A_352_406#_c_2001_n N_VGND_c_2223_n 0.00657784f $X=5.16 $Y=0.35 $X2=0
+ $Y2=0
cc_1181 N_A_352_406#_c_2003_n N_VGND_c_2223_n 0.015428f $X=2.37 $Y=0.445 $X2=0
+ $Y2=0
cc_1182 N_A_352_406#_c_2051_n N_VGND_c_2223_n 8.68625e-19 $X=3.1 $Y=0.845 $X2=0
+ $Y2=0
cc_1183 N_A_352_406#_c_1997_n A_837_108# 0.00242534f $X=4.325 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_1184 N_Q_c_2181_n N_VGND_c_2210_n 0.0153904f $X=15.56 $Y=0.495 $X2=0 $Y2=0
cc_1185 N_Q_c_2181_n N_VGND_c_2222_n 0.0218641f $X=15.56 $Y=0.495 $X2=0 $Y2=0
cc_1186 N_Q_c_2181_n N_VGND_c_2223_n 0.0125454f $X=15.56 $Y=0.495 $X2=0 $Y2=0
cc_1187 A_144_47# N_VGND_c_2223_n 0.00396664f $X=0.72 $Y=0.235 $X2=15.6 $Y2=0
cc_1188 N_VGND_c_2223_n A_368_47# 0.0034141f $X=15.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1189 N_VGND_c_2223_n A_532_47# 0.00323414f $X=15.6 $Y=0 $X2=-0.19 $Y2=-0.245
