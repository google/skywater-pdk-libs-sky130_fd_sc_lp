* File: sky130_fd_sc_lp__a21boi_4.spice
* Created: Fri Aug 28 09:50:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21boi_4.pex.spice"
.subckt sky130_fd_sc_lp__a21boi_4  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_B1_N_M1014_g N_A_33_367#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.2226 PD=1.14 PS=2.21 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75005.7 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1014_d N_A_33_367#_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.126 AS=0.1176 PD=1.14 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6 SB=75005.3
+ A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A_33_367#_M1005_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.8 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1005_d N_A_33_367#_M1017_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75004.4 A=0.126 P=1.98 MULT=1
MM1018 N_VGND_M1018_d N_A_33_367#_M1018_g N_Y_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9 SB=75004
+ A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1018_d N_A2_M1004_g N_A_658_47#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.7
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1003 N_A_658_47#_M1004_s N_A1_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.1
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1008 N_A_658_47#_M1008_d N_A1_M1008_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1020 N_A_658_47#_M1008_d N_A1_M1020_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004 SB=75001.9
+ A=0.126 P=1.98 MULT=1
MM1021 N_A_658_47#_M1021_d N_A1_M1021_g N_Y_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.4
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_658_47#_M1021_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.9
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1010_d N_A2_M1015_g N_A_658_47#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.3
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1023 N_VGND_M1023_d N_A2_M1023_g N_A_658_47#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_B1_N_M1007_g N_A_33_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_A_223_367#_M1002_d N_A_33_367#_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005 A=0.189 P=2.82 MULT=1
MM1009 N_A_223_367#_M1009_d N_A_33_367#_M1009_g N_Y_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1016 N_A_223_367#_M1009_d N_A_33_367#_M1016_g N_Y_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1022 N_A_223_367#_M1022_d N_A_33_367#_M1022_g N_Y_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1953 AS=0.1764 PD=1.57 PS=1.54 NRD=4.6886 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75003.7 A=0.189 P=2.82 MULT=1
MM1001 N_A_223_367#_M1022_d N_A2_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1953 AS=0.1827 PD=1.57 PS=1.55 NRD=0 NRS=1.5563 M=1 R=8.4
+ SA=75001.9 SB=75003.2 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1001_s N_A1_M1006_g N_A_223_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1827 AS=0.1764 PD=1.55 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g N_A_223_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1012_d N_A1_M1019_g N_A_223_367#_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1024 N_VPWR_M1024_d N_A1_M1024_g N_A_223_367#_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_A_223_367#_M1011_d N_A2_M1011_g N_VPWR_M1024_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1013 N_A_223_367#_M1011_d N_A2_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_A_223_367#_M1025_d N_A2_M1025_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=13.2415 P=17.93
*
.include "sky130_fd_sc_lp__a21boi_4.pxi.spice"
*
.ends
*
*
