* NGSPICE file created from sky130_fd_sc_lp__a31oi_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a31oi_lp A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 VPWR A2 a_139_409# VPB phighvt w=1e+06u l=250000u
+  ad=6.05e+11p pd=5.21e+06u as=5.6e+11p ps=5.12e+06u
M1001 a_139_409# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_175_47# A3 VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.394e+11p ps=2.82e+06u
M1003 a_253_47# A2 a_175_47# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1004 Y A1 a_253_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1005 a_417_47# B1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1006 VGND B1 a_417_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_139_409# A3 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y B1 a_139_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends

