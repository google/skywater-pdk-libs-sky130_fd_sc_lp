* File: sky130_fd_sc_lp__a21o_2.spice
* Created: Wed Sep  2 09:20:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21o_2.pex.spice"
.subckt sky130_fd_sc_lp__a21o_2  VNB VPB B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_X_M1001_d N_A_86_269#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1009 N_X_M1001_d N_A_86_269#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1428 PD=1.12 PS=1.18 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1003 N_A_86_269#_M1003_d N_B1_M1003_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.21 AS=0.1428 PD=1.34 PS=1.18 NRD=0 NRS=8.568 M=1 R=5.6 SA=75001.1
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1005 A_464_47# N_A1_M1005_g N_A_86_269#_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.21 PD=1.23 PS=1.34 NRD=19.992 NRS=31.428 M=1 R=5.6 SA=75001.8
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g A_464_47# VNB NSHORT L=0.15 W=0.84 AD=0.231
+ AS=0.1638 PD=2.23 PS=1.23 NRD=1.428 NRS=19.992 M=1 R=5.6 SA=75002.3 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1002 N_X_M1002_d N_A_86_269#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_X_M1002_d N_A_86_269#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_A_392_367#_M1000_d N_B1_M1000_g N_A_86_269#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_392_367#_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1004 N_A_392_367#_M1004_d N_A2_M1004_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2016 PD=3.05 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a21o_2.pxi.spice"
*
.ends
*
*
