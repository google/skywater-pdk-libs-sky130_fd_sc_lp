* NGSPICE file created from sky130_fd_sc_lp__einvp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__einvp_2 A TE VGND VNB VPB VPWR Z
M1000 VGND TE a_30_131# VNB nshort w=420000u l=150000u
+  ad=4.914e+11p pd=4.64e+06u as=1.113e+11p ps=1.37e+06u
M1001 Z A a_249_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.0206e+12p ps=9.18e+06u
M1002 a_218_47# A Z VNB nshort w=840000u l=150000u
+  ad=6.804e+11p pd=6.66e+06u as=2.352e+11p ps=2.24e+06u
M1003 VPWR a_30_131# a_249_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=5.224e+11p pd=4.89e+06u as=0p ps=0u
M1004 a_218_47# TE VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_249_367# a_30_131# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR TE a_30_131# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1007 a_249_367# A Z VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND TE a_218_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z A a_218_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

