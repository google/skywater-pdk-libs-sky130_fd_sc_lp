* File: sky130_fd_sc_lp__o211a_4.pex.spice
* Created: Fri Aug 28 11:02:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211A_4%A_80_21# 1 2 3 4 15 19 23 27 31 35 39 43 45
+ 54 56 57 58 59 60 63 67 71 73 75 77 82 93
c149 2 0 1.61007e-19 $X=2.66 $Y=1.835
r150 90 91 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.725 $Y=1.48
+ $X2=1.765 $Y2=1.48
r151 89 90 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=1.335 $Y=1.48
+ $X2=1.725 $Y2=1.48
r152 88 89 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.295 $Y=1.48
+ $X2=1.335 $Y2=1.48
r153 87 88 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=0.905 $Y=1.48
+ $X2=1.295 $Y2=1.48
r154 86 87 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.865 $Y=1.48
+ $X2=0.905 $Y2=1.48
r155 77 79 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.535 $Y=1.07
+ $X2=3.535 $Y2=1.15
r156 69 71 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=5.5 $Y=2.27
+ $X2=5.5 $Y2=2.035
r157 68 82 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=4.3 $Y=2.355
+ $X2=4.132 $Y2=2.355
r158 67 69 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.335 $Y=2.355
+ $X2=5.5 $Y2=2.27
r159 67 68 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=5.335 $Y=2.355
+ $X2=4.3 $Y2=2.355
r160 64 75 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.295 $Y=2.355
+ $X2=3 $Y2=2.355
r161 63 82 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=3.965 $Y=2.355
+ $X2=4.132 $Y2=2.355
r162 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.965 $Y=2.355
+ $X2=3.295 $Y2=2.355
r163 59 75 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.705 $Y=2.355
+ $X2=3 $Y2=2.355
r164 59 60 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.705 $Y=2.355
+ $X2=2.375 $Y2=2.355
r165 57 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.37 $Y=1.15
+ $X2=3.535 $Y2=1.15
r166 57 58 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=3.37 $Y=1.15
+ $X2=2.375 $Y2=1.15
r167 56 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.29 $Y=2.27
+ $X2=2.375 $Y2=2.355
r168 55 73 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.29 $Y=1.585 $X2=2.29
+ $Y2=1.485
r169 55 56 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.29 $Y=1.585
+ $X2=2.29 $Y2=2.27
r170 54 73 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.29 $Y=1.385 $X2=2.29
+ $Y2=1.485
r171 53 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.29 $Y=1.235
+ $X2=2.375 $Y2=1.15
r172 53 54 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.29 $Y=1.235
+ $X2=2.29 $Y2=1.385
r173 52 93 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.065 $Y=1.48
+ $X2=2.155 $Y2=1.48
r174 52 91 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.065 $Y=1.48
+ $X2=1.765 $Y2=1.48
r175 51 52 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.065
+ $Y=1.48 $X2=2.065 $Y2=1.48
r176 48 86 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.705 $Y=1.48
+ $X2=0.865 $Y2=1.48
r177 48 83 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=0.705 $Y=1.48
+ $X2=0.475 $Y2=1.48
r178 47 51 75.4182 $w=1.98e-07 $l=1.36e-06 $layer=LI1_cond $X=0.705 $Y=1.485
+ $X2=2.065 $Y2=1.485
r179 47 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.705
+ $Y=1.48 $X2=0.705 $Y2=1.48
r180 45 73 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=1.485
+ $X2=2.29 $Y2=1.485
r181 45 51 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=2.205 $Y=1.485
+ $X2=2.065 $Y2=1.485
r182 41 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.645
+ $X2=2.155 $Y2=1.48
r183 41 43 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.155 $Y=1.645
+ $X2=2.155 $Y2=2.465
r184 37 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.315
+ $X2=1.765 $Y2=1.48
r185 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.765 $Y=1.315
+ $X2=1.765 $Y2=0.655
r186 33 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.645
+ $X2=1.725 $Y2=1.48
r187 33 35 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.725 $Y=1.645
+ $X2=1.725 $Y2=2.465
r188 29 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.315
+ $X2=1.335 $Y2=1.48
r189 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.315
+ $X2=1.335 $Y2=0.655
r190 25 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.295 $Y=1.645
+ $X2=1.295 $Y2=1.48
r191 25 27 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.295 $Y=1.645
+ $X2=1.295 $Y2=2.465
r192 21 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.315
+ $X2=0.905 $Y2=1.48
r193 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.315
+ $X2=0.905 $Y2=0.655
r194 17 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.865 $Y=1.645
+ $X2=0.865 $Y2=1.48
r195 17 19 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.865 $Y=1.645
+ $X2=0.865 $Y2=2.465
r196 13 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.315
+ $X2=0.475 $Y2=1.48
r197 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.315
+ $X2=0.475 $Y2=0.655
r198 4 71 300 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=2 $X=5.36
+ $Y=1.835 $X2=5.5 $Y2=2.035
r199 3 82 300 $w=1.7e-07 $l=6.97137e-07 $layer=licon1_PDIFF $count=2 $X=3.92
+ $Y=1.835 $X2=4.13 $Y2=2.435
r200 2 75 150 $w=1.7e-07 $l=8.27043e-07 $layer=licon1_PDIFF $count=4 $X=2.66
+ $Y=1.835 $X2=3.2 $Y2=2.435
r201 1 77 182 $w=1.7e-07 $l=9.35147e-07 $layer=licon1_NDIFF $count=1 $X=3.3
+ $Y=0.245 $X2=3.535 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%B1 3 7 11 15 17 21 22 24 25 33 44
c85 33 0 1.27614e-19 $X=2.795 $Y=1.51
c86 22 0 1.84755e-19 $X=4.295 $Y=1.51
c87 17 0 1.61007e-19 $X=4.13 $Y=2.015
c88 15 0 8.24151e-20 $X=4.385 $Y=2.465
r89 31 33 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=2.71 $Y=1.51
+ $X2=2.795 $Y2=1.51
r90 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.51 $X2=2.71 $Y2=1.51
r91 28 31 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.585 $Y=1.51
+ $X2=2.71 $Y2=1.51
r92 25 44 10.6009 $w=6.93e-07 $l=1.55e-07 $layer=LI1_cond $X=3.12 $Y=1.752
+ $X2=3.275 $Y2=1.752
r93 25 32 7.056 $w=6.93e-07 $l=4.1e-07 $layer=LI1_cond $X=3.12 $Y=1.752 $X2=2.71
+ $Y2=1.752
r94 24 32 1.20468 $w=6.93e-07 $l=7e-08 $layer=LI1_cond $X=2.64 $Y=1.752 $X2=2.71
+ $Y2=1.752
r95 22 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.295 $Y=1.51
+ $X2=4.295 $Y2=1.675
r96 22 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.295 $Y=1.51
+ $X2=4.295 $Y2=1.345
r97 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.51 $X2=4.295 $Y2=1.51
r98 19 21 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.295 $Y=1.93
+ $X2=4.295 $Y2=1.51
r99 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.13 $Y=2.015
+ $X2=4.295 $Y2=1.93
r100 17 44 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.13 $Y=2.015
+ $X2=3.275 $Y2=2.015
r101 15 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.385 $Y=2.465
+ $X2=4.385 $Y2=1.675
r102 11 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.275 $Y=0.665
+ $X2=4.275 $Y2=1.345
r103 5 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.345
+ $X2=2.795 $Y2=1.51
r104 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.795 $Y=1.345
+ $X2=2.795 $Y2=0.665
r105 1 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.585 $Y=1.675
+ $X2=2.585 $Y2=1.51
r106 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.585 $Y=1.675
+ $X2=2.585 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%C1 3 7 11 15 17 24 25
c48 24 0 2.10029e-19 $X=3.755 $Y=1.51
r49 23 25 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.755 $Y=1.51
+ $X2=3.845 $Y2=1.51
r50 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.755
+ $Y=1.51 $X2=3.755 $Y2=1.51
r51 21 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.415 $Y=1.51
+ $X2=3.755 $Y2=1.51
r52 19 21 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.225 $Y=1.51
+ $X2=3.415 $Y2=1.51
r53 17 24 5.03179 $w=3.53e-07 $l=1.55e-07 $layer=LI1_cond $X=3.6 $Y=1.582
+ $X2=3.755 $Y2=1.582
r54 13 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.675
+ $X2=3.845 $Y2=1.51
r55 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.845 $Y=1.675
+ $X2=3.845 $Y2=2.465
r56 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.345
+ $X2=3.845 $Y2=1.51
r57 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.845 $Y=1.345
+ $X2=3.845 $Y2=0.665
r58 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=1.675
+ $X2=3.415 $Y2=1.51
r59 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.415 $Y=1.675
+ $X2=3.415 $Y2=2.465
r60 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.225 $Y=1.345
+ $X2=3.225 $Y2=1.51
r61 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.225 $Y=1.345
+ $X2=3.225 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%A1 3 6 8 10 13 15 17 20 21 22 27 32 35 37
c71 37 0 5.26839e-20 $X=6.48 $Y=1.295
c72 20 0 1.24029e-19 $X=4.835 $Y=1.36
c73 17 0 1.24362e-19 $X=4.835 $Y=1.17
r74 35 37 1.44055 $w=3.18e-07 $l=4e-08 $layer=LI1_cond $X=6.475 $Y=1.255
+ $X2=6.475 $Y2=1.295
r75 29 32 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=6.145 $Y=1.36
+ $X2=6.45 $Y2=1.36
r76 21 35 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.475 $Y=1.17
+ $X2=6.475 $Y2=1.255
r77 21 22 12.5328 $w=3.18e-07 $l=3.48e-07 $layer=LI1_cond $X=6.475 $Y=1.317
+ $X2=6.475 $Y2=1.665
r78 21 37 0.792305 $w=3.18e-07 $l=2.2e-08 $layer=LI1_cond $X=6.475 $Y=1.317
+ $X2=6.475 $Y2=1.295
r79 21 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.36 $X2=6.45 $Y2=1.36
r80 20 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.36
+ $X2=4.835 $Y2=1.525
r81 20 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.36
+ $X2=4.835 $Y2=1.195
r82 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.835
+ $Y=1.36 $X2=4.835 $Y2=1.36
r83 17 19 7.9931 $w=2.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.835 $Y=1.17
+ $X2=4.835 $Y2=1.36
r84 16 17 3.86198 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5 $Y=1.17 $X2=4.835
+ $Y2=1.17
r85 15 21 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.315 $Y=1.17
+ $X2=6.475 $Y2=1.17
r86 15 16 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=6.315 $Y=1.17
+ $X2=5 $Y2=1.17
r87 11 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.145 $Y=1.525
+ $X2=6.145 $Y2=1.36
r88 11 13 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=6.145 $Y=1.525 $X2=6.145
+ $Y2=2.465
r89 8 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.145 $Y=1.195
+ $X2=6.145 $Y2=1.36
r90 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.145 $Y=1.195
+ $X2=6.145 $Y2=0.665
r91 6 28 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.855 $Y=2.465 $X2=4.855
+ $Y2=1.525
r92 3 27 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.745 $Y=0.665
+ $X2=4.745 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%A2 3 7 11 15 17 18 26
c53 26 0 1.77046e-19 $X=5.715 $Y=1.51
c54 18 0 1.24029e-19 $X=6 $Y=1.665
r55 24 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.375 $Y=1.51
+ $X2=5.715 $Y2=1.51
r56 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.375
+ $Y=1.51 $X2=5.375 $Y2=1.51
r57 21 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.285 $Y=1.51
+ $X2=5.375 $Y2=1.51
r58 17 18 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.592 $X2=6
+ $Y2=1.592
r59 17 25 4.98819 $w=3.33e-07 $l=1.45e-07 $layer=LI1_cond $X=5.52 $Y=1.592
+ $X2=5.375 $Y2=1.592
r60 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.675
+ $X2=5.715 $Y2=1.51
r61 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.715 $Y=1.675
+ $X2=5.715 $Y2=2.465
r62 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.345
+ $X2=5.715 $Y2=1.51
r63 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.715 $Y=1.345
+ $X2=5.715 $Y2=0.665
r64 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.675
+ $X2=5.285 $Y2=1.51
r65 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.285 $Y=1.675
+ $X2=5.285 $Y2=2.465
r66 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.345
+ $X2=5.285 $Y2=1.51
r67 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.285 $Y=1.345
+ $X2=5.285 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%VPWR 1 2 3 4 5 6 21 27 33 37 41 43 45 50 51
+ 53 54 55 57 69 73 78 87 90 93 97
r96 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r97 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r98 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r99 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 85 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r101 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r102 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r103 82 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r104 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r105 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 79 93 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.735 $Y=3.33
+ $X2=4.602 $Y2=3.33
r107 79 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.735 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 78 96 4.58274 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=6.457 $Y2=3.33
r109 78 84 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=6 $Y2=3.33
r110 77 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r111 77 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r112 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r113 74 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.63 $Y2=3.33
r114 74 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=4.08 $Y2=3.33
r115 73 93 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.47 $Y=3.33
+ $X2=4.602 $Y2=3.33
r116 73 76 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.47 $Y=3.33
+ $X2=4.08 $Y2=3.33
r117 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r118 69 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.63 $Y2=3.33
r119 69 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.12 $Y2=3.33
r120 68 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r121 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r122 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r123 65 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r125 62 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.65 $Y2=3.33
r126 62 64 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 60 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r128 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r129 57 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.65 $Y2=3.33
r130 57 59 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.24 $Y2=3.33
r131 55 91 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r132 55 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r133 53 67 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.205 $Y=3.33
+ $X2=2.16 $Y2=3.33
r134 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=3.33
+ $X2=2.37 $Y2=3.33
r135 52 71 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=3.12 $Y2=3.33
r136 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=2.37 $Y2=3.33
r137 50 64 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.51 $Y2=3.33
r139 49 67 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=2.16 $Y2=3.33
r140 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=3.33
+ $X2=1.51 $Y2=3.33
r141 45 48 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=6.36 $Y=2.015
+ $X2=6.36 $Y2=2.95
r142 43 96 3.18343 $w=3.3e-07 $l=1.32868e-07 $layer=LI1_cond $X=6.36 $Y=3.245
+ $X2=6.457 $Y2=3.33
r143 43 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.36 $Y=3.245
+ $X2=6.36 $Y2=2.95
r144 39 93 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.602 $Y=3.245
+ $X2=4.602 $Y2=3.33
r145 39 41 20.4396 $w=2.63e-07 $l=4.7e-07 $layer=LI1_cond $X=4.602 $Y=3.245
+ $X2=4.602 $Y2=2.775
r146 35 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=3.245
+ $X2=3.63 $Y2=3.33
r147 35 37 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=3.63 $Y=3.245
+ $X2=3.63 $Y2=2.775
r148 31 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=3.245
+ $X2=2.37 $Y2=3.33
r149 31 33 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=2.37 $Y=3.245
+ $X2=2.37 $Y2=2.73
r150 27 30 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.51 $Y=2.18
+ $X2=1.51 $Y2=2.95
r151 25 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=3.245
+ $X2=1.51 $Y2=3.33
r152 25 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.51 $Y=3.245
+ $X2=1.51 $Y2=2.95
r153 21 24 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.65 $Y=2.18
+ $X2=0.65 $Y2=2.95
r154 19 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=3.245
+ $X2=0.65 $Y2=3.33
r155 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.65 $Y=3.245
+ $X2=0.65 $Y2=2.95
r156 6 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.22
+ $Y=1.835 $X2=6.36 $Y2=2.95
r157 6 45 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=6.22
+ $Y=1.835 $X2=6.36 $Y2=2.015
r158 5 41 600 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=1.835 $X2=4.6 $Y2=2.775
r159 4 37 600 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=1.835 $X2=3.63 $Y2=2.775
r160 3 33 600 $w=1.7e-07 $l=9.62458e-07 $layer=licon1_PDIFF $count=1 $X=2.23
+ $Y=1.835 $X2=2.37 $Y2=2.73
r161 2 30 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.37
+ $Y=1.835 $X2=1.51 $Y2=2.95
r162 2 27 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.37
+ $Y=1.835 $X2=1.51 $Y2=2.18
r163 1 24 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.525
+ $Y=1.835 $X2=0.65 $Y2=2.95
r164 1 21 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.525
+ $Y=1.835 $X2=0.65 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%X 1 2 3 4 13 15 16 19 21 25 29 33 37 42 43
+ 44 45 49 51
r55 49 51 3.23493 $w=2.83e-07 $l=8e-08 $layer=LI1_cond $X=0.227 $Y=1.215
+ $X2=0.227 $Y2=1.295
r56 44 49 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.227 $Y=1.13
+ $X2=0.227 $Y2=1.215
r57 44 45 14.8807 $w=2.83e-07 $l=3.68e-07 $layer=LI1_cond $X=0.227 $Y=1.297
+ $X2=0.227 $Y2=1.665
r58 44 51 0.0808732 $w=2.83e-07 $l=2e-09 $layer=LI1_cond $X=0.227 $Y=1.297
+ $X2=0.227 $Y2=1.295
r59 41 45 3.63929 $w=2.83e-07 $l=9e-08 $layer=LI1_cond $X=0.227 $Y=1.755
+ $X2=0.227 $Y2=1.665
r60 37 39 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.94 $Y=1.98
+ $X2=1.94 $Y2=2.91
r61 35 37 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.94 $Y=1.925
+ $X2=1.94 $Y2=1.98
r62 31 33 34.6591 $w=1.98e-07 $l=6.25e-07 $layer=LI1_cond $X=1.555 $Y=1.045
+ $X2=1.555 $Y2=0.42
r63 30 43 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.165 $Y=1.84 $X2=1.075
+ $Y2=1.84
r64 29 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.845 $Y=1.84
+ $X2=1.94 $Y2=1.925
r65 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.845 $Y=1.84
+ $X2=1.165 $Y2=1.84
r66 25 27 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=1.075 $Y=1.98
+ $X2=1.075 $Y2=2.91
r67 23 43 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.075 $Y=1.925
+ $X2=1.075 $Y2=1.84
r68 23 25 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=1.075 $Y=1.925
+ $X2=1.075 $Y2=1.98
r69 22 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.785 $Y=1.13
+ $X2=0.69 $Y2=1.13
r70 21 31 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.455 $Y=1.13
+ $X2=1.555 $Y2=1.045
r71 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.455 $Y=1.13
+ $X2=0.785 $Y2=1.13
r72 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.045
+ $X2=0.69 $Y2=1.13
r73 17 19 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=0.69 $Y=1.045
+ $X2=0.69 $Y2=0.42
r74 16 41 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.37 $Y=1.84
+ $X2=0.227 $Y2=1.755
r75 15 43 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.985 $Y=1.84 $X2=1.075
+ $Y2=1.84
r76 15 16 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.985 $Y=1.84
+ $X2=0.37 $Y2=1.84
r77 14 44 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=0.37 $Y=1.13
+ $X2=0.227 $Y2=1.13
r78 13 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.595 $Y=1.13
+ $X2=0.69 $Y2=1.13
r79 13 14 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.595 $Y=1.13
+ $X2=0.37 $Y2=1.13
r80 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.8
+ $Y=1.835 $X2=1.94 $Y2=2.91
r81 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.8
+ $Y=1.835 $X2=1.94 $Y2=1.98
r82 3 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.94
+ $Y=1.835 $X2=1.08 $Y2=2.91
r83 3 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.94
+ $Y=1.835 $X2=1.08 $Y2=1.98
r84 2 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.42
r85 1 19 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%A_986_367# 1 2 7 11 13
r13 11 16 4.39812 $w=1.9e-07 $l=1.47e-07 $layer=LI1_cond $X=5.93 $Y=2.78
+ $X2=5.93 $Y2=2.927
r14 11 13 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=5.93 $Y=2.78
+ $X2=5.93 $Y2=2.095
r15 7 16 2.84233 $w=2.95e-07 $l=9.5e-08 $layer=LI1_cond $X=5.835 $Y=2.927
+ $X2=5.93 $Y2=2.927
r16 7 9 29.8854 $w=2.93e-07 $l=7.65e-07 $layer=LI1_cond $X=5.835 $Y=2.927
+ $X2=5.07 $Y2=2.927
r17 2 16 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.835 $X2=5.93 $Y2=2.91
r18 2 13 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=5.79
+ $Y=1.835 $X2=5.93 $Y2=2.095
r19 1 9 600 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=4.93
+ $Y=1.835 $X2=5.07 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 42 44 53 65 66 72 75
r98 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r99 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r100 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r101 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r102 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r103 63 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r104 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r105 60 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5
+ $Y2=0
r106 60 62 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.52 $Y2=0
r107 59 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r108 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r109 55 58 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r110 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r111 53 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5
+ $Y2=0
r112 53 58 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.56 $Y2=0
r113 52 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r114 52 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r115 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r116 49 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r117 49 51 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.68 $Y2=0
r118 48 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r119 48 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r120 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 45 69 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r122 45 47 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r123 44 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r124 44 47 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=0
+ $X2=0.72 $Y2=0
r125 42 59 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.56
+ $Y2=0
r126 42 56 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.16
+ $Y2=0
r127 40 62 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.835 $Y=0
+ $X2=5.52 $Y2=0
r128 40 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.835 $Y=0 $X2=5.93
+ $Y2=0
r129 39 65 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.025 $Y=0
+ $X2=6.48 $Y2=0
r130 39 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.025 $Y=0 $X2=5.93
+ $Y2=0
r131 37 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.68
+ $Y2=0
r132 37 38 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.967
+ $Y2=0
r133 36 55 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.16
+ $Y2=0
r134 36 38 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=2.085 $Y=0
+ $X2=1.967 $Y2=0
r135 32 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=0.085
+ $X2=5.93 $Y2=0
r136 32 34 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=5.93 $Y=0.085
+ $X2=5.93 $Y2=0.41
r137 28 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r138 28 30 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.44
r139 24 38 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.967 $Y=0.085
+ $X2=1.967 $Y2=0
r140 24 26 14.4668 $w=2.33e-07 $l=2.95e-07 $layer=LI1_cond $X=1.967 $Y=0.085
+ $X2=1.967 $Y2=0.38
r141 20 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r142 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.36
r143 16 69 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r144 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r145 5 34 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.79
+ $Y=0.245 $X2=5.93 $Y2=0.41
r146 4 30 182 $w=1.7e-07 $l=2.70416e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.245 $X2=5 $Y2=0.44
r147 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.38
r148 2 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.36
r149 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%A_475_49# 1 2 3 4 13 15 17 21 23 27 29 33 38
+ 41
c68 17 0 1.84755e-19 $X=4.365 $Y=0.72
r69 38 40 1.22819 $w=2.98e-07 $l=3e-08 $layer=LI1_cond $X=4.515 $Y=0.83
+ $X2=4.515 $Y2=0.86
r70 37 38 4.50336 $w=2.98e-07 $l=1.1e-07 $layer=LI1_cond $X=4.515 $Y=0.72
+ $X2=4.515 $Y2=0.83
r71 31 33 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.36 $Y=0.745
+ $X2=6.36 $Y2=0.42
r72 30 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=0.83
+ $X2=5.5 $Y2=0.83
r73 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.195 $Y=0.83
+ $X2=6.36 $Y2=0.745
r74 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.195 $Y=0.83
+ $X2=5.665 $Y2=0.83
r75 25 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=0.745 $X2=5.5
+ $Y2=0.83
r76 25 27 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.5 $Y=0.745
+ $X2=5.5 $Y2=0.42
r77 24 38 4.02169 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.665 $Y=0.83
+ $X2=4.515 $Y2=0.83
r78 23 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0.83
+ $X2=5.5 $Y2=0.83
r79 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.335 $Y=0.83
+ $X2=4.665 $Y2=0.83
r80 19 37 3.61266 $w=2.98e-07 $l=9.21954e-08 $layer=LI1_cond $X=4.53 $Y=0.635
+ $X2=4.515 $Y2=0.72
r81 19 21 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.53 $Y=0.635
+ $X2=4.53 $Y2=0.43
r82 18 36 4.79676 $w=1.7e-07 $l=1.86145e-07 $layer=LI1_cond $X=2.665 $Y=0.72
+ $X2=2.5 $Y2=0.765
r83 17 37 4.02169 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.365 $Y=0.72
+ $X2=4.515 $Y2=0.72
r84 17 18 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=4.365 $Y=0.72
+ $X2=2.665 $Y2=0.72
r85 13 36 2.96942 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=2.5 $Y=0.635 $X2=2.5
+ $Y2=0.765
r86 13 15 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.5 $Y=0.635
+ $X2=2.5 $Y2=0.39
r87 4 33 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=6.22
+ $Y=0.245 $X2=6.36 $Y2=0.42
r88 3 27 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.245 $X2=5.5 $Y2=0.42
r89 2 40 182 $w=1.7e-07 $l=6.99232e-07 $layer=licon1_NDIFF $count=1 $X=4.35
+ $Y=0.245 $X2=4.53 $Y2=0.86
r90 2 21 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=4.35
+ $Y=0.245 $X2=4.53 $Y2=0.43
r91 1 36 182 $w=1.7e-07 $l=5.94222e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.245 $X2=2.5 $Y2=0.78
r92 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.245 $X2=2.5 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_4%A_574_49# 1 2 11
r13 8 11 55.4545 $w=2.08e-07 $l=1.05e-06 $layer=LI1_cond $X=3.01 $Y=0.36
+ $X2=4.06 $Y2=0.36
r14 2 11 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.245 $X2=4.06 $Y2=0.37
r15 1 8 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.87
+ $Y=0.245 $X2=3.01 $Y2=0.37
.ends

