* File: sky130_fd_sc_lp__or2b_4.pex.spice
* Created: Fri Aug 28 11:22:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2B_4%B_N 3 5 6 7 9 12 13 14 15 16 17 24
r35 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=0.93 $X2=0.385 $Y2=0.93
r36 16 17 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=2.035
r37 15 16 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.315 $Y=1.295
+ $X2=0.315 $Y2=1.665
r38 15 25 9.49062 $w=4.58e-07 $l=3.65e-07 $layer=LI1_cond $X=0.315 $Y=1.295
+ $X2=0.315 $Y2=0.93
r39 14 25 0.130009 $w=4.58e-07 $l=5e-09 $layer=LI1_cond $X=0.315 $Y=0.925
+ $X2=0.315 $Y2=0.93
r40 13 14 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.315 $Y=0.555
+ $X2=0.315 $Y2=0.925
r41 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.27
+ $X2=0.385 $Y2=0.93
r42 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.27
+ $X2=0.385 $Y2=1.435
r43 10 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.385 $Y=0.915
+ $X2=0.385 $Y2=0.93
r44 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.095 $Y=0.765
+ $X2=1.095 $Y2=0.445
r45 6 10 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.55 $Y=0.84
+ $X2=0.385 $Y2=0.915
r46 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.02 $Y=0.84
+ $X2=1.095 $Y2=0.765
r47 5 6 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.02 $Y=0.84 $X2=0.55
+ $Y2=0.84
r48 3 12 643.521 $w=1.5e-07 $l=1.255e-06 $layer=POLY_cond $X=0.475 $Y=2.69
+ $X2=0.475 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_4%A_27_496# 1 2 7 8 9 11 14 17 20 22 23 26 30
r58 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=1.35 $X2=0.955 $Y2=1.35
r59 26 29 31.7795 $w=3.28e-07 $l=9.1e-07 $layer=LI1_cond $X=0.88 $Y=0.44
+ $X2=0.88 $Y2=1.35
r60 24 29 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=0.88 $Y=2.3 $X2=0.88
+ $Y2=1.35
r61 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.715 $Y=2.385
+ $X2=0.88 $Y2=2.3
r62 22 23 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.715 $Y=2.385
+ $X2=0.355 $Y2=2.385
r63 18 23 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=2.47
+ $X2=0.355 $Y2=2.385
r64 18 20 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=0.225 $Y=2.47
+ $X2=0.225 $Y2=2.69
r65 16 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.955 $Y=1.335
+ $X2=0.955 $Y2=1.35
r66 12 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.62 $Y=1.335
+ $X2=1.62 $Y2=1.26
r67 12 14 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=1.62 $Y=1.335
+ $X2=1.62 $Y2=2.465
r68 9 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.62 $Y=1.185
+ $X2=1.62 $Y2=1.26
r69 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.62 $Y=1.185
+ $X2=1.62 $Y2=0.655
r70 8 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.12 $Y=1.26
+ $X2=0.955 $Y2=1.335
r71 7 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.545 $Y=1.26
+ $X2=1.62 $Y2=1.26
r72 7 8 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=1.545 $Y=1.26
+ $X2=1.12 $Y2=1.26
r73 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.48 $X2=0.26 $Y2=2.69
r74 1 26 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.755
+ $Y=0.235 $X2=0.88 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_4%A 3 7 9 10 14
r32 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.51
+ $X2=2.07 $Y2=1.675
r33 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.51
+ $X2=2.07 $Y2=1.345
r34 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=1.51 $X2=2.07 $Y2=1.51
r35 10 15 3.09612 $w=3.33e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=1.592 $X2=2.07
+ $Y2=1.592
r36 9 15 13.4165 $w=3.33e-07 $l=3.9e-07 $layer=LI1_cond $X=1.68 $Y=1.592
+ $X2=2.07 $Y2=1.592
r37 7 16 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.05 $Y=0.655
+ $X2=2.05 $Y2=1.345
r38 3 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.98 $Y=2.465
+ $X2=1.98 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_4%A_256_367# 1 2 9 13 17 21 25 29 33 37 43 45
+ 46 49 51 58 62 63 64 77
r116 69 71 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.61 $Y=1.5 $X2=2.52
+ $Y2=1.5
r117 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.5 $X2=2.61 $Y2=1.5
r118 62 63 6.71914 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.405 $Y=2.05
+ $X2=1.405 $Y2=1.93
r119 59 77 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.63 $Y=1.5 $X2=3.81
+ $Y2=1.5
r120 59 75 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.63 $Y=1.5
+ $X2=3.38 $Y2=1.5
r121 58 59 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.63
+ $Y=1.5 $X2=3.63 $Y2=1.5
r122 56 75 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.95 $Y=1.5
+ $X2=3.38 $Y2=1.5
r123 56 69 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.95 $Y=1.5
+ $X2=2.61 $Y2=1.5
r124 55 58 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.95 $Y=1.5
+ $X2=3.63 $Y2=1.5
r125 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.5 $X2=2.95 $Y2=1.5
r126 53 68 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.79 $Y=1.5
+ $X2=2.617 $Y2=1.5
r127 53 55 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.79 $Y=1.5
+ $X2=2.95 $Y2=1.5
r128 52 64 6.19399 $w=1.8e-07 $l=1.13e-07 $layer=LI1_cond $X=1.965 $Y=1.165
+ $X2=1.852 $Y2=1.165
r129 51 68 11.1904 $w=3.43e-07 $l=3.35e-07 $layer=LI1_cond $X=2.617 $Y=1.165
+ $X2=2.617 $Y2=1.5
r130 51 52 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=2.445 $Y=1.165
+ $X2=1.965 $Y2=1.165
r131 47 64 0.552779 $w=2.25e-07 $l=9e-08 $layer=LI1_cond $X=1.852 $Y=1.075
+ $X2=1.852 $Y2=1.165
r132 47 49 33.5489 $w=2.23e-07 $l=6.55e-07 $layer=LI1_cond $X=1.852 $Y=1.075
+ $X2=1.852 $Y2=0.42
r133 45 64 6.19399 $w=1.8e-07 $l=1.12e-07 $layer=LI1_cond $X=1.74 $Y=1.165
+ $X2=1.852 $Y2=1.165
r134 45 46 20.0253 $w=1.78e-07 $l=3.25e-07 $layer=LI1_cond $X=1.74 $Y=1.165
+ $X2=1.415 $Y2=1.165
r135 41 62 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.405 $Y=2.095
+ $X2=1.405 $Y2=2.05
r136 41 43 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.405 $Y=2.095
+ $X2=1.405 $Y2=2.95
r137 39 46 6.81825 $w=1.8e-07 $l=1.2657e-07 $layer=LI1_cond $X=1.327 $Y=1.255
+ $X2=1.415 $Y2=1.165
r138 39 63 42.7792 $w=1.73e-07 $l=6.75e-07 $layer=LI1_cond $X=1.327 $Y=1.255
+ $X2=1.327 $Y2=1.93
r139 35 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.665
+ $X2=3.81 $Y2=1.5
r140 35 37 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.81 $Y=1.665
+ $X2=3.81 $Y2=2.465
r141 31 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.335
+ $X2=3.81 $Y2=1.5
r142 31 33 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.81 $Y=1.335
+ $X2=3.81 $Y2=0.655
r143 27 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.665
+ $X2=3.38 $Y2=1.5
r144 27 29 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.38 $Y=1.665
+ $X2=3.38 $Y2=2.465
r145 23 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.335
+ $X2=3.38 $Y2=1.5
r146 23 25 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.38 $Y=1.335
+ $X2=3.38 $Y2=0.655
r147 19 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.665
+ $X2=2.95 $Y2=1.5
r148 19 21 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.95 $Y=1.665
+ $X2=2.95 $Y2=2.465
r149 15 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.335
+ $X2=2.95 $Y2=1.5
r150 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.95 $Y=1.335
+ $X2=2.95 $Y2=0.655
r151 11 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.52 $Y=1.665
+ $X2=2.52 $Y2=1.5
r152 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.52 $Y=1.665
+ $X2=2.52 $Y2=2.465
r153 7 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.52 $Y=1.335
+ $X2=2.52 $Y2=1.5
r154 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.52 $Y=1.335
+ $X2=2.52 $Y2=0.655
r155 2 62 400 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=1.28
+ $Y=1.835 $X2=1.405 $Y2=2.05
r156 2 43 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=1.28
+ $Y=1.835 $X2=1.405 $Y2=2.95
r157 1 49 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.695
+ $Y=0.235 $X2=1.835 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_4%VPWR 1 2 3 4 15 19 25 29 31 35 37 42 47 52 58
+ 61 64 68
r61 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 56 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 56 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r67 53 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=3.33
+ $X2=3.165 $Y2=3.33
r68 53 55 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.33 $Y=3.33 $X2=3.6
+ $Y2=3.33
r69 52 67 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.86 $Y=3.33 $X2=4.09
+ $Y2=3.33
r70 52 55 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.86 $Y=3.33 $X2=3.6
+ $Y2=3.33
r71 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r73 48 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.245 $Y2=3.33
r74 48 50 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.64 $Y2=3.33
r75 47 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3 $Y=3.33 $X2=3.165
+ $Y2=3.33
r76 47 50 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3 $Y=3.33 $X2=2.64
+ $Y2=3.33
r77 46 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r79 43 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r80 43 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r81 42 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.08 $Y=3.33
+ $X2=2.245 $Y2=3.33
r82 42 45 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=2.08 $Y=3.33 $X2=1.2
+ $Y2=3.33
r83 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r84 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r85 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r86 37 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 35 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r89 35 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r90 31 34 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=4.025 $Y=2.2
+ $X2=4.025 $Y2=2.97
r91 29 67 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.025 $Y=3.245
+ $X2=4.09 $Y2=3.33
r92 29 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.025 $Y=3.245
+ $X2=4.025 $Y2=2.97
r93 25 28 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.165 $Y=2.2
+ $X2=3.165 $Y2=2.97
r94 23 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=3.245
+ $X2=3.165 $Y2=3.33
r95 23 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.165 $Y=3.245
+ $X2=3.165 $Y2=2.97
r96 19 22 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=2.245 $Y=2.015
+ $X2=2.245 $Y2=2.95
r97 17 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=3.245
+ $X2=2.245 $Y2=3.33
r98 17 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.245 $Y=3.245
+ $X2=2.245 $Y2=2.95
r99 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r100 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.745
r101 4 34 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.835 $X2=4.025 $Y2=2.97
r102 4 31 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.835 $X2=4.025 $Y2=2.2
r103 3 28 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.025
+ $Y=1.835 $X2=3.165 $Y2=2.97
r104 3 25 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=3.025
+ $Y=1.835 $X2=3.165 $Y2=2.2
r105 2 22 400 $w=1.7e-07 $l=1.20626e-06 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.835 $X2=2.245 $Y2=2.95
r106 2 19 400 $w=1.7e-07 $l=2.65141e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.835 $X2=2.245 $Y2=2.015
r107 1 15 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.48 $X2=0.69 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 44 45
+ 47 48 52 54
r68 52 54 2.13415 $w=2.68e-07 $l=5e-08 $layer=LI1_cond $X=4.1 $Y=1.245 $X2=4.1
+ $Y2=1.295
r69 47 52 2.87089 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=4.1 $Y=1.155 $X2=4.1
+ $Y2=1.245
r70 47 48 15.0671 $w=2.68e-07 $l=3.53e-07 $layer=LI1_cond $X=4.1 $Y=1.312
+ $X2=4.1 $Y2=1.665
r71 47 54 0.725612 $w=2.68e-07 $l=1.7e-08 $layer=LI1_cond $X=4.1 $Y=1.312
+ $X2=4.1 $Y2=1.295
r72 46 48 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=4.1 $Y=1.755 $X2=4.1
+ $Y2=1.665
r73 40 45 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.69 $Y=1.85
+ $X2=3.595 $Y2=1.85
r74 39 46 7.08811 $w=1.9e-07 $l=1.7621e-07 $layer=LI1_cond $X=3.965 $Y=1.85
+ $X2=4.1 $Y2=1.755
r75 39 40 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=3.965 $Y=1.85
+ $X2=3.69 $Y2=1.85
r76 38 44 3.06858 $w=3.45e-07 $l=2.07123e-07 $layer=LI1_cond $X=3.69 $Y=1.155
+ $X2=3.595 $Y2=0.99
r77 37 47 4.30634 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=3.965 $Y=1.155
+ $X2=4.1 $Y2=1.155
r78 37 38 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=3.965 $Y=1.155
+ $X2=3.69 $Y2=1.155
r79 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.595 $Y=1.98
+ $X2=3.595 $Y2=2.91
r80 31 45 1.34256 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.595 $Y=1.945
+ $X2=3.595 $Y2=1.85
r81 31 33 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=3.595 $Y=1.945
+ $X2=3.595 $Y2=1.98
r82 27 44 3.55614 $w=1.9e-07 $l=2.55e-07 $layer=LI1_cond $X=3.595 $Y=0.735
+ $X2=3.595 $Y2=0.99
r83 27 29 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=3.595 $Y=0.735
+ $X2=3.595 $Y2=0.42
r84 25 44 3.06858 $w=3.45e-07 $l=9.5e-08 $layer=LI1_cond $X=3.5 $Y=0.99
+ $X2=3.595 $Y2=0.99
r85 25 26 6.68397 $w=5.08e-07 $l=2.85e-07 $layer=LI1_cond $X=3.5 $Y=0.99
+ $X2=3.215 $Y2=0.99
r86 23 45 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.5 $Y=1.85 $X2=3.595
+ $Y2=1.85
r87 23 24 39.11 $w=1.88e-07 $l=6.7e-07 $layer=LI1_cond $X=3.5 $Y=1.85 $X2=2.83
+ $Y2=1.85
r88 19 21 42.8709 $w=2.48e-07 $l=9.3e-07 $layer=LI1_cond $X=2.705 $Y=1.98
+ $X2=2.705 $Y2=2.91
r89 17 24 6.98266 $w=1.9e-07 $l=1.65831e-07 $layer=LI1_cond $X=2.705 $Y=1.945
+ $X2=2.83 $Y2=1.85
r90 17 19 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=2.705 $Y=1.945
+ $X2=2.705 $Y2=1.98
r91 13 26 14.2942 $w=5.1e-07 $l=6.29722e-07 $layer=LI1_cond $X=2.7 $Y=0.735
+ $X2=3.215 $Y2=0.99
r92 13 15 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.7 $Y=0.735
+ $X2=2.7 $Y2=0.42
r93 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.835 $X2=3.595 $Y2=2.91
r94 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.835 $X2=3.595 $Y2=1.98
r95 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.595
+ $Y=1.835 $X2=2.735 $Y2=2.91
r96 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.595
+ $Y=1.835 $X2=2.735 $Y2=1.98
r97 2 44 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.235 $X2=3.595 $Y2=0.93
r98 2 29 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.235 $X2=3.595 $Y2=0.42
r99 1 13 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.235 $X2=2.735 $Y2=0.82
r100 1 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.235 $X2=2.735 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR2B_4%VGND 1 2 3 4 15 17 21 25 27 29 31 32 33 42 47
+ 53 56 60
r73 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r74 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r75 51 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r76 51 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r77 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r78 48 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.165
+ $Y2=0
r79 48 50 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.6
+ $Y2=0
r80 47 59 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.86 $Y=0 $X2=4.09
+ $Y2=0
r81 47 50 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.86 $Y=0 $X2=3.6
+ $Y2=0
r82 46 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r83 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r84 43 53 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.267
+ $Y2=0
r85 43 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r86 42 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3 $Y=0 $X2=3.165
+ $Y2=0
r87 42 45 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3 $Y=0 $X2=2.64
+ $Y2=0
r88 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r89 37 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r90 36 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r91 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r92 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r93 33 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r94 33 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r95 31 40 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.2
+ $Y2=0
r96 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=0 $X2=1.405
+ $Y2=0
r97 27 59 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.025 $Y=0.085
+ $X2=4.09 $Y2=0
r98 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.025 $Y=0.085
+ $X2=4.025 $Y2=0.38
r99 23 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=0.085
+ $X2=3.165 $Y2=0
r100 23 25 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.165 $Y=0.085
+ $X2=3.165 $Y2=0.445
r101 19 53 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.267 $Y=0.085
+ $X2=2.267 $Y2=0
r102 19 21 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=2.267 $Y=0.085
+ $X2=2.267 $Y2=0.38
r103 18 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.405
+ $Y2=0
r104 17 53 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.135 $Y=0
+ $X2=2.267 $Y2=0
r105 17 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.135 $Y=0 $X2=1.57
+ $Y2=0
r106 13 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.405 $Y=0.085
+ $X2=1.405 $Y2=0
r107 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.405 $Y=0.085
+ $X2=1.405 $Y2=0.38
r108 4 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.235 $X2=4.025 $Y2=0.38
r109 3 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.235 $X2=3.165 $Y2=0.445
r110 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.125
+ $Y=0.235 $X2=2.265 $Y2=0.38
r111 1 15 91 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=2 $X=1.17
+ $Y=0.235 $X2=1.405 $Y2=0.38
.ends

