* File: sky130_fd_sc_lp__nand3_2.pex.spice
* Created: Fri Aug 28 10:49:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3_2%A 1 3 6 8 10 12 15 17 18 19 27
c45 10 0 5.42978e-20 $X=0.985 $Y=1.275
r46 26 27 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.555 $Y=1.44
+ $X2=0.63 $Y2=1.44
r47 23 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.34 $Y=1.44
+ $X2=0.555 $Y2=1.44
r48 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.44 $X2=0.34 $Y2=1.44
r49 19 24 6.1738 $w=4.18e-07 $l=2.25e-07 $layer=LI1_cond $X=0.295 $Y=1.665
+ $X2=0.295 $Y2=1.44
r50 18 24 3.97867 $w=4.18e-07 $l=1.45e-07 $layer=LI1_cond $X=0.295 $Y=1.295
+ $X2=0.295 $Y2=1.44
r51 13 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.985 $Y=1.425
+ $X2=0.985 $Y2=1.35
r52 13 15 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=0.985 $Y=1.425
+ $X2=0.985 $Y2=2.465
r53 10 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.985 $Y=1.275
+ $X2=0.985 $Y2=1.35
r54 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.985 $Y=1.275
+ $X2=0.985 $Y2=0.745
r55 8 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.91 $Y=1.35
+ $X2=0.985 $Y2=1.35
r56 8 27 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.91 $Y=1.35 $X2=0.63
+ $Y2=1.35
r57 4 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.605
+ $X2=0.555 $Y2=1.44
r58 4 6 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.555 $Y=1.605
+ $X2=0.555 $Y2=2.465
r59 1 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.275
+ $X2=0.555 $Y2=1.44
r60 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.555 $Y=1.275
+ $X2=0.555 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_2%B 3 7 11 15 18 19 21 22 24 26 27 34 35 41 44
c84 34 0 9.92477e-20 $X=1.435 $Y=1.51
c85 18 0 5.23255e-20 $X=2.617 $Y=1.92
c86 7 0 8.37963e-20 $X=1.455 $Y=2.465
r87 42 50 6.0869 $w=2e-07 $l=2.48e-07 $layer=LI1_cond $X=1.6 $Y=2.02 $X2=1.352
+ $Y2=2.02
r88 42 44 4.43636 $w=1.98e-07 $l=8e-08 $layer=LI1_cond $X=1.6 $Y=2.02 $X2=1.68
+ $Y2=2.02
r89 35 50 12.3232 $w=4.93e-07 $l=5.1e-07 $layer=LI1_cond $X=1.352 $Y=1.51
+ $X2=1.352 $Y2=2.02
r90 34 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.51
+ $X2=1.435 $Y2=1.675
r91 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.51
+ $X2=1.435 $Y2=1.345
r92 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.435
+ $Y=1.51 $X2=1.435 $Y2=1.51
r93 27 41 3.88656 $w=2e-07 $l=1.27e-07 $layer=LI1_cond $X=2.617 $Y=2.02 $X2=2.49
+ $Y2=2.02
r94 26 41 18.3 $w=1.98e-07 $l=3.3e-07 $layer=LI1_cond $X=2.16 $Y=2.02 $X2=2.49
+ $Y2=2.02
r95 24 50 0.362448 $w=4.93e-07 $l=1.5e-08 $layer=LI1_cond $X=1.352 $Y=2.035
+ $X2=1.352 $Y2=2.02
r96 24 26 26.5073 $w=1.98e-07 $l=4.78e-07 $layer=LI1_cond $X=1.682 $Y=2.02
+ $X2=2.16 $Y2=2.02
r97 24 44 0.110909 $w=1.98e-07 $l=2e-09 $layer=LI1_cond $X=1.682 $Y=2.02
+ $X2=1.68 $Y2=2.02
r98 22 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.51
+ $X2=2.885 $Y2=1.675
r99 22 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.51
+ $X2=2.885 $Y2=1.345
r100 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.885
+ $Y=1.51 $X2=2.885 $Y2=1.51
r101 19 21 7.33373 $w=2.18e-07 $l=1.4e-07 $layer=LI1_cond $X=2.745 $Y=1.535
+ $X2=2.885 $Y2=1.535
r102 18 27 3.06028 $w=2.55e-07 $l=1e-07 $layer=LI1_cond $X=2.617 $Y=1.92
+ $X2=2.617 $Y2=2.02
r103 17 19 6.86474 $w=2.2e-07 $l=1.74539e-07 $layer=LI1_cond $X=2.617 $Y=1.645
+ $X2=2.745 $Y2=1.535
r104 17 18 12.4283 $w=2.53e-07 $l=2.75e-07 $layer=LI1_cond $X=2.617 $Y=1.645
+ $X2=2.617 $Y2=1.92
r105 15 39 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.865 $Y=0.745
+ $X2=2.865 $Y2=1.345
r106 11 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.795 $Y=2.465
+ $X2=2.795 $Y2=1.675
r107 7 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.455 $Y=2.465
+ $X2=1.455 $Y2=1.675
r108 3 36 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.415 $Y=0.745
+ $X2=1.415 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_2%C 3 7 11 15 17 23
c52 17 0 8.37963e-20 $X=2.16 $Y=1.665
c53 3 0 6.40318e-20 $X=1.885 $Y=0.745
r54 23 24 10.8141 $w=3.12e-07 $l=7e-08 $layer=POLY_cond $X=2.365 $Y=1.51
+ $X2=2.435 $Y2=1.51
r55 21 23 60.25 $w=3.12e-07 $l=3.9e-07 $layer=POLY_cond $X=1.975 $Y=1.51
+ $X2=2.365 $Y2=1.51
r56 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.975
+ $Y=1.51 $X2=1.975 $Y2=1.51
r57 19 21 13.9038 $w=3.12e-07 $l=9e-08 $layer=POLY_cond $X=1.885 $Y=1.51
+ $X2=1.975 $Y2=1.51
r58 17 22 6.56006 $w=3.23e-07 $l=1.85e-07 $layer=LI1_cond $X=2.16 $Y=1.587
+ $X2=1.975 $Y2=1.587
r59 13 24 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.345
+ $X2=2.435 $Y2=1.51
r60 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.435 $Y=1.345
+ $X2=2.435 $Y2=0.745
r61 9 23 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.675
+ $X2=2.365 $Y2=1.51
r62 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.365 $Y=1.675
+ $X2=2.365 $Y2=2.465
r63 5 19 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.675
+ $X2=1.885 $Y2=1.51
r64 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.885 $Y=1.675
+ $X2=1.885 $Y2=2.465
r65 1 19 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.345
+ $X2=1.885 $Y2=1.51
r66 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.885 $Y=1.345 $X2=1.885
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_2%VPWR 1 2 3 4 13 15 21 25 27 29 33 35 40 45
+ 54 57 61
r57 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 49 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 49 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 46 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.12 $Y2=3.33
r65 46 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 45 60 4.01281 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r67 45 48 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 41 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.22 $Y2=3.33
r69 41 43 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 40 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=2.12 $Y2=3.33
r71 40 43 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 39 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 36 51 4.61231 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.252 $Y2=3.33
r76 36 38 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.505 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 35 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.22 $Y2=3.33
r78 35 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 33 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r80 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r81 33 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r82 29 32 42.995 $w=2.58e-07 $l=9.7e-07 $layer=LI1_cond $X=3.045 $Y=1.98
+ $X2=3.045 $Y2=2.95
r83 27 60 3.19941 $w=2.6e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.045 $Y=3.245
+ $X2=3.137 $Y2=3.33
r84 27 32 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.045 $Y=3.245
+ $X2=3.045 $Y2=2.95
r85 23 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=3.33
r86 23 25 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.785
r87 19 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r88 19 21 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.755
r89 15 18 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.34 $Y=2.005
+ $X2=0.34 $Y2=2.95
r90 13 51 3.15387 $w=3.3e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.252 $Y2=3.33
r91 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.34 $Y=3.245
+ $X2=0.34 $Y2=2.95
r92 4 32 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.835 $X2=3.01 $Y2=2.95
r93 4 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=1.835 $X2=3.01 $Y2=1.98
r94 3 25 600 $w=1.7e-07 $l=1.02689e-06 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.835 $X2=2.12 $Y2=2.785
r95 2 21 600 $w=1.7e-07 $l=9.96795e-07 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.835 $X2=1.22 $Y2=2.755
r96 1 18 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.95
r97 1 15 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.835 $X2=0.34 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_2%Y 1 2 3 4 16 19 23 25 27 30 36 39 40 43
c48 39 0 9.92477e-20 $X=1.67 $Y=2.375
r49 40 43 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=2.455 $Y=2.39
+ $X2=2.16 $Y2=2.39
r50 40 42 4.21383 $w=2e-07 $l=1.45e-07 $layer=LI1_cond $X=2.455 $Y=2.39 $X2=2.6
+ $Y2=2.39
r51 37 43 20.7955 $w=1.98e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=2.39
+ $X2=2.16 $Y2=2.39
r52 37 39 6.1674 $w=1.85e-07 $l=1.15e-07 $layer=LI1_cond $X=1.785 $Y=2.39
+ $X2=1.67 $Y2=2.39
r53 33 34 1.59825 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.77 $Y=1.04 $X2=0.77
+ $Y2=1.07
r54 30 33 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.77 $Y=0.68
+ $X2=0.77 $Y2=1.04
r55 25 42 2.90609 $w=2.9e-07 $l=1e-07 $layer=LI1_cond $X=2.6 $Y=2.49 $X2=2.6
+ $Y2=2.39
r56 25 27 16.6906 $w=2.88e-07 $l=4.2e-07 $layer=LI1_cond $X=2.6 $Y=2.49 $X2=2.6
+ $Y2=2.91
r57 21 39 0.571601 $w=2.3e-07 $l=1e-07 $layer=LI1_cond $X=1.67 $Y=2.49 $X2=1.67
+ $Y2=2.39
r58 21 23 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.67 $Y=2.49
+ $X2=1.67 $Y2=2.91
r59 20 36 2.53056 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.935 $Y=2.375
+ $X2=0.805 $Y2=2.375
r60 19 39 6.1674 $w=1.85e-07 $l=1.2227e-07 $layer=LI1_cond $X=1.555 $Y=2.375
+ $X2=1.67 $Y2=2.39
r61 19 20 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.555 $Y=2.375
+ $X2=0.935 $Y2=2.375
r62 16 34 39.449 $w=2.58e-07 $l=8.9e-07 $layer=LI1_cond $X=0.805 $Y=1.96
+ $X2=0.805 $Y2=1.07
r63 14 36 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=2.29
+ $X2=0.805 $Y2=2.375
r64 14 16 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=0.805 $Y=2.29
+ $X2=0.805 $Y2=1.96
r65 4 42 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.835 $X2=2.58 $Y2=2.375
r66 4 27 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.44
+ $Y=1.835 $X2=2.58 $Y2=2.91
r67 3 39 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.835 $X2=1.67 $Y2=2.375
r68 3 23 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.835 $X2=1.67 $Y2=2.91
r69 2 36 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=2.44
r70 2 16 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=1.96
r71 1 33 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.325 $X2=0.77 $Y2=1.04
r72 1 30 182 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.325 $X2=0.77 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_2%A_43_65# 1 2 3 12 14 15 20 21 24
r45 22 24 27.2597 $w=2.58e-07 $l=6.15e-07 $layer=LI1_cond $X=3.115 $Y=1.085
+ $X2=3.115 $Y2=0.47
r46 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.985 $Y=1.17
+ $X2=3.115 $Y2=1.085
r47 20 21 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=2.985 $Y=1.17
+ $X2=1.315 $Y2=1.17
r48 17 21 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.21 $Y=1.085
+ $X2=1.315 $Y2=1.17
r49 17 19 32.4805 $w=2.08e-07 $l=6.15e-07 $layer=LI1_cond $X=1.21 $Y=1.085
+ $X2=1.21 $Y2=0.47
r50 16 19 2.37662 $w=2.08e-07 $l=4.5e-08 $layer=LI1_cond $X=1.21 $Y=0.425
+ $X2=1.21 $Y2=0.47
r51 14 16 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.105 $Y=0.34
+ $X2=1.21 $Y2=0.425
r52 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.105 $Y=0.34
+ $X2=0.435 $Y2=0.34
r53 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.305 $Y=0.425
+ $X2=0.435 $Y2=0.34
r54 10 12 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=0.305 $Y=0.425
+ $X2=0.305 $Y2=0.47
r55 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.325 $X2=3.08 $Y2=0.47
r56 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.06
+ $Y=0.325 $X2=1.2 $Y2=0.47
r57 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.215
+ $Y=0.325 $X2=0.34 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_2%A_298_65# 1 2 9 11 12 15
c29 12 0 6.40318e-20 $X=1.815 $Y=0.83
c30 9 0 5.42978e-20 $X=1.65 $Y=0.45
r31 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.65 $Y=0.745
+ $X2=2.65 $Y2=0.45
r32 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.485 $Y=0.83
+ $X2=2.65 $Y2=0.745
r33 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.485 $Y=0.83
+ $X2=1.815 $Y2=0.83
r34 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.65 $Y=0.745
+ $X2=1.815 $Y2=0.83
r35 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.65 $Y=0.745
+ $X2=1.65 $Y2=0.45
r36 2 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.51
+ $Y=0.325 $X2=2.65 $Y2=0.45
r37 1 9 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=1.49
+ $Y=0.325 $X2=1.65 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_2%VGND 1 6 8 10 20 21 24
r38 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r39 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r40 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.15
+ $Y2=0
r42 18 20 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=3.12
+ $Y2=0
r43 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r44 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r45 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.15
+ $Y2=0
r46 10 16 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=1.68
+ $Y2=0
r47 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r48 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r49 8 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r50 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0.085 $X2=2.15
+ $Y2=0
r51 4 6 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0.45
r52 1 6 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.325 $X2=2.15 $Y2=0.45
.ends

