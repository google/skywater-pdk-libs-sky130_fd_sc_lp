* NGSPICE file created from sky130_fd_sc_lp__sleep_sergate_plv_14.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sleep_sergate_plv_14 VIRTPWR VPWR SLEEP VPB
M1000 VIRTPWR SLEEP VPWR VPB phighvt w=7e+06u l=150000u
+  ad=3.71e+12p pd=2.906e+07u as=1.96e+12p ps=1.456e+07u
M1001 VPWR SLEEP VIRTPWR VPB phighvt w=7e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

