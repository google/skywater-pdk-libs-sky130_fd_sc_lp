* File: sky130_fd_sc_lp__nand2_8.pxi.spice
* Created: Wed Sep  2 10:02:57 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2_8%B N_B_M1001_g N_B_M1000_g N_B_M1008_g N_B_M1004_g
+ N_B_M1012_g N_B_M1010_g N_B_M1014_g N_B_M1015_g N_B_M1019_g N_B_M1021_g
+ N_B_M1024_g N_B_M1022_g N_B_M1029_g N_B_M1028_g N_B_M1031_g N_B_M1030_g
+ N_B_c_153_p B B N_B_c_138_n N_B_c_148_n B B N_B_c_190_p N_B_c_150_n
+ PM_SKY130_FD_SC_LP__NAND2_8%B
x_PM_SKY130_FD_SC_LP__NAND2_8%A N_A_M1003_g N_A_M1002_g N_A_M1006_g N_A_M1005_g
+ N_A_M1009_g N_A_M1007_g N_A_c_280_n N_A_M1013_g N_A_M1011_g N_A_M1020_g
+ N_A_M1016_g N_A_M1023_g N_A_M1017_g N_A_M1026_g N_A_M1018_g N_A_M1027_g
+ N_A_M1025_g N_A_c_286_n N_A_c_287_n N_A_c_288_n N_A_c_289_n N_A_c_290_n A A A
+ N_A_c_306_n N_A_c_291_n PM_SKY130_FD_SC_LP__NAND2_8%A
x_PM_SKY130_FD_SC_LP__NAND2_8%VPWR N_VPWR_M1000_s N_VPWR_M1004_s N_VPWR_M1015_s
+ N_VPWR_M1022_s N_VPWR_M1030_s N_VPWR_M1005_d N_VPWR_M1011_d N_VPWR_M1017_d
+ N_VPWR_M1025_d N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n
+ N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n
+ N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n
+ N_VPWR_c_439_n N_VPWR_c_440_n VPWR N_VPWR_c_441_n N_VPWR_c_442_n
+ N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n
+ N_VPWR_c_448_n N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_424_n
+ PM_SKY130_FD_SC_LP__NAND2_8%VPWR
x_PM_SKY130_FD_SC_LP__NAND2_8%Y N_Y_M1003_d N_Y_M1009_d N_Y_M1020_d N_Y_M1026_d
+ N_Y_M1000_d N_Y_M1010_d N_Y_M1021_d N_Y_M1028_d N_Y_M1002_s N_Y_M1007_s
+ N_Y_M1016_s N_Y_M1018_s N_Y_c_656_n N_Y_c_560_n N_Y_c_561_n N_Y_c_562_n
+ N_Y_c_661_n N_Y_c_578_n N_Y_c_665_n N_Y_c_583_n N_Y_c_669_n N_Y_c_563_n
+ N_Y_c_564_n N_Y_c_673_n N_Y_c_601_n N_Y_c_555_n N_Y_c_677_n N_Y_c_609_n
+ N_Y_c_611_n N_Y_c_556_n N_Y_c_681_n N_Y_c_704_p N_Y_c_619_n N_Y_c_683_n
+ N_Y_c_590_n N_Y_c_565_n N_Y_c_622_n N_Y_c_557_n N_Y_c_558_n Y Y Y N_Y_c_639_n
+ Y PM_SKY130_FD_SC_LP__NAND2_8%Y
x_PM_SKY130_FD_SC_LP__NAND2_8%A_27_65# N_A_27_65#_M1001_d N_A_27_65#_M1008_d
+ N_A_27_65#_M1014_d N_A_27_65#_M1024_d N_A_27_65#_M1031_d N_A_27_65#_M1006_s
+ N_A_27_65#_M1013_s N_A_27_65#_M1023_s N_A_27_65#_M1027_s N_A_27_65#_c_709_n
+ N_A_27_65#_c_710_n N_A_27_65#_c_711_n N_A_27_65#_c_712_n N_A_27_65#_c_713_n
+ N_A_27_65#_c_714_n N_A_27_65#_c_715_n N_A_27_65#_c_716_n N_A_27_65#_c_717_n
+ N_A_27_65#_c_718_n N_A_27_65#_c_719_n N_A_27_65#_c_763_n N_A_27_65#_c_720_n
+ N_A_27_65#_c_767_n N_A_27_65#_c_721_n N_A_27_65#_c_771_n N_A_27_65#_c_722_n
+ N_A_27_65#_c_723_n N_A_27_65#_c_724_n N_A_27_65#_c_725_n N_A_27_65#_c_726_n
+ N_A_27_65#_c_727_n N_A_27_65#_c_728_n N_A_27_65#_c_729_n
+ PM_SKY130_FD_SC_LP__NAND2_8%A_27_65#
x_PM_SKY130_FD_SC_LP__NAND2_8%VGND N_VGND_M1001_s N_VGND_M1012_s N_VGND_M1019_s
+ N_VGND_M1029_s N_VGND_c_841_n N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n
+ N_VGND_c_845_n N_VGND_c_846_n N_VGND_c_847_n N_VGND_c_848_n N_VGND_c_849_n
+ VGND N_VGND_c_850_n N_VGND_c_851_n N_VGND_c_852_n N_VGND_c_853_n
+ N_VGND_c_854_n PM_SKY130_FD_SC_LP__NAND2_8%VGND
cc_1 VNB N_B_M1001_g 0.0262168f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.745
cc_2 VNB N_B_M1008_g 0.0191761f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.745
cc_3 VNB N_B_M1012_g 0.0191762f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.745
cc_4 VNB N_B_M1014_g 0.0191761f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.745
cc_5 VNB N_B_M1019_g 0.0191761f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.745
cc_6 VNB N_B_M1024_g 0.0191761f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.745
cc_7 VNB N_B_M1029_g 0.0191761f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=0.745
cc_8 VNB N_B_M1031_g 0.0194864f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=0.745
cc_9 VNB N_B_c_138_n 0.143645f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=1.51
cc_10 VNB N_A_M1003_g 0.019335f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.745
cc_11 VNB N_A_M1006_g 0.0198055f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.745
cc_12 VNB N_A_M1009_g 0.0206404f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.745
cc_13 VNB N_A_c_280_n 0.0154066f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.345
cc_14 VNB N_A_M1013_g 0.0206642f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.675
cc_15 VNB N_A_M1020_g 0.0201905f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.675
cc_16 VNB N_A_M1023_g 0.0186252f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.675
cc_17 VNB N_A_M1026_g 0.018254f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=1.675
cc_18 VNB N_A_M1027_g 0.0260721f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=1.675
cc_19 VNB N_A_c_286_n 0.0281326f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_20 VNB N_A_c_287_n 0.015408f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=1.51
cc_21 VNB N_A_c_288_n 0.004935f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=1.51
cc_22 VNB N_A_c_289_n 0.015408f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=1.51
cc_23 VNB N_A_c_290_n 0.0749315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_c_291_n 0.004935f $X=-0.19 $Y=-0.245 $X2=1.98 $Y2=1.51
cc_25 VNB N_VPWR_c_424_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_555_n 0.00311043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_556_n 0.00309095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_557_n 0.00227088f $X=-0.19 $Y=-0.245 $X2=2.66 $Y2=1.587
cc_29 VNB N_Y_c_558_n 4.39188e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB Y 8.58945e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_65#_c_709_n 0.0312591f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=2.465
cc_32 VNB N_A_27_65#_c_710_n 0.00332611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_65#_c_711_n 0.0115731f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.345
cc_34 VNB N_A_27_65#_c_712_n 0.00176121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_65#_c_713_n 0.00313892f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=2.465
cc_36 VNB N_A_27_65#_c_714_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.745
cc_37 VNB N_A_27_65#_c_715_n 0.00304705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_65#_c_716_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_65#_c_717_n 0.00680897f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=0.745
cc_40 VNB N_A_27_65#_c_718_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_65#_c_719_n 0.00190976f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=1.345
cc_42 VNB N_A_27_65#_c_720_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=2.465
cc_43 VNB N_A_27_65#_c_721_n 0.00227356f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_44 VNB N_A_27_65#_c_722_n 0.0122515f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=1.51
cc_45 VNB N_A_27_65#_c_723_n 0.0339267f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_46 VNB N_A_27_65#_c_724_n 0.00134924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_65#_c_725_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_65#_c_726_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_65#_c_727_n 0.00221189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_65#_c_728_n 0.00221131f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_51 VNB N_A_27_65#_c_729_n 0.00163793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_841_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_53 VNB N_VGND_c_842_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.745
cc_54 VNB N_VGND_c_843_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_55 VNB N_VGND_c_844_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.345
cc_56 VNB N_VGND_c_845_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=1.675
cc_57 VNB N_VGND_c_846_n 0.0143749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_847_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=1.345
cc_59 VNB N_VGND_c_848_n 0.0142895f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.745
cc_60 VNB N_VGND_c_849_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=0.745
cc_61 VNB N_VGND_c_850_n 0.0161944f $X=-0.19 $Y=-0.245 $X2=2.195 $Y2=2.465
cc_62 VNB N_VGND_c_851_n 0.098614f $X=-0.19 $Y=-0.245 $X2=3.055 $Y2=2.465
cc_63 VNB N_VGND_c_852_n 0.409365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_853_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=0.745
cc_65 VNB N_VGND_c_854_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=2.465
cc_66 VPB N_B_M1000_g 0.0249083f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_67 VPB N_B_M1004_g 0.0179297f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_68 VPB N_B_M1010_g 0.0179236f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_69 VPB N_B_M1015_g 0.01818f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.465
cc_70 VPB N_B_M1021_g 0.0178521f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=2.465
cc_71 VPB N_B_M1022_g 0.0178338f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=2.465
cc_72 VPB N_B_M1028_g 0.01825f $X=-0.19 $Y=1.655 $X2=3.055 $Y2=2.465
cc_73 VPB N_B_M1030_g 0.018168f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=2.465
cc_74 VPB N_B_c_138_n 0.025911f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=1.51
cc_75 VPB N_B_c_148_n 0.00260038f $X=-0.19 $Y=1.655 $X2=2.653 $Y2=1.587
cc_76 VPB B 0.00260385f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.665
cc_77 VPB N_B_c_150_n 0.00210831f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=1.587
cc_78 VPB N_A_M1002_g 0.0177655f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_79 VPB N_A_M1005_g 0.0194465f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_80 VPB N_A_M1007_g 0.0196195f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_81 VPB N_A_c_280_n 0.00559875f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.345
cc_82 VPB N_A_M1011_g 0.0196201f $X=-0.19 $Y=1.655 $X2=2.195 $Y2=1.345
cc_83 VPB N_A_M1016_g 0.0194742f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=1.345
cc_84 VPB N_A_M1017_g 0.0175255f $X=-0.19 $Y=1.655 $X2=3.055 $Y2=1.345
cc_85 VPB N_A_M1018_g 0.0171771f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=1.345
cc_86 VPB N_A_M1025_g 0.0255361f $X=-0.19 $Y=1.655 $X2=1.815 $Y2=1.505
cc_87 VPB N_A_c_286_n 0.00449101f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.51
cc_88 VPB N_A_c_287_n 0.00559875f $X=-0.19 $Y=1.655 $X2=1.64 $Y2=1.51
cc_89 VPB N_A_c_288_n 3.18387e-19 $X=-0.19 $Y=1.655 $X2=1.64 $Y2=1.51
cc_90 VPB N_A_c_289_n 0.00559875f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=1.51
cc_91 VPB N_A_c_290_n 0.0136599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_c_306_n 0.010146f $X=-0.19 $Y=1.655 $X2=1.98 $Y2=1.51
cc_93 VPB N_A_c_291_n 3.18387e-19 $X=-0.19 $Y=1.655 $X2=1.98 $Y2=1.51
cc_94 VPB N_VPWR_c_425_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_426_n 0.0567831f $X=-0.19 $Y=1.655 $X2=1.765 $Y2=2.465
cc_96 VPB N_VPWR_c_427_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_428_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=2.625 $Y2=0.745
cc_98 VPB N_VPWR_c_429_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=2.625 $Y2=2.465
cc_99 VPB N_VPWR_c_430_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_431_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_432_n 0.00443131f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=0.745
cc_102 VPB N_VPWR_c_433_n 0.00446949f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=2.465
cc_103 VPB N_VPWR_c_434_n 3.30321e-19 $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.505
cc_104 VPB N_VPWR_c_435_n 0.0124346f $X=-0.19 $Y=1.655 $X2=1.64 $Y2=1.505
cc_105 VPB N_VPWR_c_436_n 0.00903456f $X=-0.19 $Y=1.655 $X2=1.64 $Y2=1.51
cc_106 VPB N_VPWR_c_437_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_438_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.58
cc_108 VPB N_VPWR_c_439_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.58
cc_109 VPB N_VPWR_c_440_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_441_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_442_n 0.0147711f $X=-0.19 $Y=1.655 $X2=2.32 $Y2=1.51
cc_112 VPB N_VPWR_c_443_n 0.0181714f $X=-0.19 $Y=1.655 $X2=2.66 $Y2=1.51
cc_113 VPB N_VPWR_c_444_n 0.0156317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_445_n 0.0158018f $X=-0.19 $Y=1.655 $X2=2.202 $Y2=1.587
cc_115 VPB N_VPWR_c_446_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_447_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=1.587
cc_117 VPB N_VPWR_c_448_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_449_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_450_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_424_n 0.0473597f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_Y_c_560_n 0.00304538f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=0.745
cc_122 VPB N_Y_c_561_n 0.00221851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_Y_c_562_n 0.00209027f $X=-0.19 $Y=1.655 $X2=2.625 $Y2=1.675
cc_124 VPB N_Y_c_563_n 0.00557861f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=1.675
cc_125 VPB N_Y_c_564_n 6.30836e-19 $X=-0.19 $Y=1.655 $X2=3.485 $Y2=2.465
cc_126 VPB N_Y_c_565_n 0.00195933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_Y_c_558_n 0.00292033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB Y 6.3246e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 N_B_M1031_g N_A_M1003_g 0.0196923f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_130 N_B_M1030_g N_A_M1002_g 0.0196923f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_131 N_B_c_153_p N_A_c_286_n 8.15032e-19 $X=3.34 $Y=1.51 $X2=0 $Y2=0
cc_132 N_B_c_138_n N_A_c_286_n 0.0196923f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_133 N_B_M1000_g N_VPWR_c_426_n 0.0224359f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B_M1004_g N_VPWR_c_426_n 8.11603e-19 $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_135 N_B_M1000_g N_VPWR_c_427_n 7.24342e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_136 N_B_M1004_g N_VPWR_c_427_n 0.0141179f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_137 N_B_M1010_g N_VPWR_c_427_n 0.0141179f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_138 N_B_M1015_g N_VPWR_c_427_n 7.24342e-19 $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_139 N_B_M1010_g N_VPWR_c_428_n 6.77662e-19 $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_140 N_B_M1015_g N_VPWR_c_428_n 0.0149184f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_141 N_B_M1021_g N_VPWR_c_428_n 0.0149184f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_142 N_B_M1022_g N_VPWR_c_428_n 6.77662e-19 $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_143 N_B_M1021_g N_VPWR_c_429_n 6.77662e-19 $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_144 N_B_M1022_g N_VPWR_c_429_n 0.0149184f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_145 N_B_M1028_g N_VPWR_c_429_n 0.0149184f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_146 N_B_M1030_g N_VPWR_c_429_n 6.77662e-19 $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B_M1028_g N_VPWR_c_430_n 0.00486043f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_148 N_B_M1030_g N_VPWR_c_430_n 0.00486043f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_149 N_B_M1028_g N_VPWR_c_431_n 7.21513e-19 $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_150 N_B_M1030_g N_VPWR_c_431_n 0.0144515f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_151 N_B_M1010_g N_VPWR_c_437_n 0.00486043f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_152 N_B_M1015_g N_VPWR_c_437_n 0.00486043f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_153 N_B_M1021_g N_VPWR_c_439_n 0.00486043f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_154 N_B_M1022_g N_VPWR_c_439_n 0.00486043f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_155 N_B_M1000_g N_VPWR_c_441_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_156 N_B_M1004_g N_VPWR_c_441_n 0.00486043f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_157 N_B_M1000_g N_VPWR_c_424_n 0.00824727f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B_M1004_g N_VPWR_c_424_n 0.00824727f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B_M1010_g N_VPWR_c_424_n 0.00824727f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_160 N_B_M1015_g N_VPWR_c_424_n 0.00824727f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_161 N_B_M1021_g N_VPWR_c_424_n 0.00824727f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_162 N_B_M1022_g N_VPWR_c_424_n 0.00824727f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_163 N_B_M1028_g N_VPWR_c_424_n 0.00824727f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_164 N_B_M1030_g N_VPWR_c_424_n 0.00824727f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_165 N_B_M1004_g N_Y_c_560_n 0.0128166f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_166 N_B_M1010_g N_Y_c_560_n 0.0128501f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_167 N_B_c_138_n N_Y_c_560_n 0.00246472f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_168 N_B_c_190_p N_Y_c_560_n 0.0469271f $X=1.815 $Y=1.587 $X2=0 $Y2=0
cc_169 N_B_M1000_g N_Y_c_561_n 0.00188176f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_170 N_B_c_138_n N_Y_c_561_n 0.00256759f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_171 N_B_c_190_p N_Y_c_561_n 0.015388f $X=1.815 $Y=1.587 $X2=0 $Y2=0
cc_172 N_B_M1015_g N_Y_c_562_n 0.00218762f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_173 N_B_c_138_n N_Y_c_562_n 0.00256759f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_174 N_B_c_190_p N_Y_c_562_n 0.0145779f $X=1.815 $Y=1.587 $X2=0 $Y2=0
cc_175 N_B_M1015_g N_Y_c_578_n 0.0129743f $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_176 N_B_M1021_g N_Y_c_578_n 0.0121662f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_177 N_B_c_138_n N_Y_c_578_n 5.64665e-19 $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_178 B N_Y_c_578_n 0.0321215f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_179 N_B_c_190_p N_Y_c_578_n 0.00579577f $X=1.815 $Y=1.587 $X2=0 $Y2=0
cc_180 N_B_M1022_g N_Y_c_583_n 0.0122595f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B_M1028_g N_Y_c_583_n 0.0137383f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B_c_153_p N_Y_c_583_n 0.01127f $X=3.34 $Y=1.51 $X2=0 $Y2=0
cc_183 N_B_c_138_n N_Y_c_583_n 0.00161526f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_184 N_B_c_148_n N_Y_c_583_n 0.0202738f $X=2.653 $Y=1.587 $X2=0 $Y2=0
cc_185 N_B_M1030_g N_Y_c_563_n 0.0131405f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B_c_153_p N_Y_c_563_n 0.00974037f $X=3.34 $Y=1.51 $X2=0 $Y2=0
cc_187 N_B_c_138_n N_Y_c_590_n 6.37898e-19 $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_188 N_B_c_148_n N_Y_c_590_n 0.0154476f $X=2.653 $Y=1.587 $X2=0 $Y2=0
cc_189 N_B_M1022_g N_Y_c_565_n 8.08979e-19 $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_190 N_B_M1028_g N_Y_c_565_n 0.00362228f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B_c_153_p N_Y_c_565_n 0.019088f $X=3.34 $Y=1.51 $X2=0 $Y2=0
cc_192 N_B_c_138_n N_Y_c_565_n 0.00253619f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_193 N_B_M1031_g Y 0.00244993f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_194 N_B_c_153_p Y 0.0066183f $X=3.34 $Y=1.51 $X2=0 $Y2=0
cc_195 N_B_M1001_g N_A_27_65#_c_709_n 0.00354556f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_196 N_B_M1001_g N_A_27_65#_c_710_n 0.0151147f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_197 N_B_M1008_g N_A_27_65#_c_710_n 0.0132122f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_198 N_B_c_138_n N_A_27_65#_c_710_n 0.00243542f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_199 N_B_c_190_p N_A_27_65#_c_710_n 0.0399877f $X=1.815 $Y=1.587 $X2=0 $Y2=0
cc_200 N_B_M1008_g N_A_27_65#_c_712_n 8.2809e-19 $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_201 N_B_M1012_g N_A_27_65#_c_712_n 8.13915e-19 $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_202 N_B_M1012_g N_A_27_65#_c_713_n 0.0132122f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_203 N_B_M1014_g N_A_27_65#_c_713_n 0.0132122f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_204 N_B_c_138_n N_A_27_65#_c_713_n 0.00243542f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_205 N_B_c_190_p N_A_27_65#_c_713_n 0.0478626f $X=1.815 $Y=1.587 $X2=0 $Y2=0
cc_206 N_B_M1014_g N_A_27_65#_c_714_n 8.28776e-19 $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_207 N_B_M1019_g N_A_27_65#_c_714_n 8.28776e-19 $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_208 N_B_M1019_g N_A_27_65#_c_715_n 0.0132122f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_209 N_B_M1024_g N_A_27_65#_c_715_n 0.0132122f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_210 N_B_c_138_n N_A_27_65#_c_715_n 0.00243542f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_211 B N_A_27_65#_c_715_n 0.0492562f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_212 N_B_M1024_g N_A_27_65#_c_716_n 8.28776e-19 $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_213 N_B_M1029_g N_A_27_65#_c_716_n 8.28776e-19 $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_214 N_B_M1029_g N_A_27_65#_c_717_n 0.0131109f $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_215 N_B_M1031_g N_A_27_65#_c_717_n 0.0136563f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_216 N_B_c_153_p N_A_27_65#_c_717_n 0.0401504f $X=3.34 $Y=1.51 $X2=0 $Y2=0
cc_217 N_B_c_138_n N_A_27_65#_c_717_n 0.00243542f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_218 N_B_M1031_g N_A_27_65#_c_719_n 5.73473e-19 $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_219 N_B_c_138_n N_A_27_65#_c_724_n 0.00253619f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_220 N_B_c_190_p N_A_27_65#_c_724_n 0.014578f $X=1.815 $Y=1.587 $X2=0 $Y2=0
cc_221 N_B_c_138_n N_A_27_65#_c_725_n 0.00253619f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_222 B N_A_27_65#_c_725_n 0.0160732f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_223 N_B_c_138_n N_A_27_65#_c_726_n 0.00253619f $X=3.485 $Y=1.51 $X2=0 $Y2=0
cc_224 N_B_c_150_n N_A_27_65#_c_726_n 0.0156735f $X=2.825 $Y=1.587 $X2=0 $Y2=0
cc_225 N_B_M1001_g N_VGND_c_841_n 0.0124264f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_226 N_B_M1008_g N_VGND_c_841_n 0.0101212f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_227 N_B_M1012_g N_VGND_c_841_n 5.09471e-19 $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_228 N_B_M1008_g N_VGND_c_842_n 5.18777e-19 $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_229 N_B_M1012_g N_VGND_c_842_n 0.010259f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_230 N_B_M1014_g N_VGND_c_842_n 0.0101212f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_231 N_B_M1019_g N_VGND_c_842_n 5.09471e-19 $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_232 N_B_M1014_g N_VGND_c_843_n 5.09471e-19 $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_233 N_B_M1019_g N_VGND_c_843_n 0.0101212f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_234 N_B_M1024_g N_VGND_c_843_n 0.0101212f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_235 N_B_M1029_g N_VGND_c_843_n 5.09471e-19 $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_236 N_B_M1024_g N_VGND_c_844_n 0.00414769f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_237 N_B_M1029_g N_VGND_c_844_n 0.00414769f $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_238 N_B_M1024_g N_VGND_c_845_n 5.09471e-19 $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_239 N_B_M1029_g N_VGND_c_845_n 0.0101212f $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_240 N_B_M1031_g N_VGND_c_845_n 0.0101655f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_241 N_B_M1008_g N_VGND_c_846_n 0.00414769f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_242 N_B_M1012_g N_VGND_c_846_n 0.00414769f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_243 N_B_M1014_g N_VGND_c_848_n 0.00414769f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_244 N_B_M1019_g N_VGND_c_848_n 0.00414769f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_245 N_B_M1001_g N_VGND_c_850_n 0.00414769f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_246 N_B_M1031_g N_VGND_c_851_n 0.00414769f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_247 N_B_M1001_g N_VGND_c_852_n 0.00823375f $X=0.475 $Y=0.745 $X2=0 $Y2=0
cc_248 N_B_M1008_g N_VGND_c_852_n 0.00787505f $X=0.905 $Y=0.745 $X2=0 $Y2=0
cc_249 N_B_M1012_g N_VGND_c_852_n 0.00787505f $X=1.335 $Y=0.745 $X2=0 $Y2=0
cc_250 N_B_M1014_g N_VGND_c_852_n 0.00787505f $X=1.765 $Y=0.745 $X2=0 $Y2=0
cc_251 N_B_M1019_g N_VGND_c_852_n 0.00787505f $X=2.195 $Y=0.745 $X2=0 $Y2=0
cc_252 N_B_M1024_g N_VGND_c_852_n 0.00787505f $X=2.625 $Y=0.745 $X2=0 $Y2=0
cc_253 N_B_M1029_g N_VGND_c_852_n 0.00787505f $X=3.055 $Y=0.745 $X2=0 $Y2=0
cc_254 N_B_M1031_g N_VGND_c_852_n 0.0078848f $X=3.485 $Y=0.745 $X2=0 $Y2=0
cc_255 N_A_M1002_g N_VPWR_c_431_n 0.0145321f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_256 N_A_M1005_g N_VPWR_c_431_n 7.35732e-19 $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A_M1005_g N_VPWR_c_432_n 0.00287895f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A_M1007_g N_VPWR_c_432_n 0.00302413f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A_M1011_g N_VPWR_c_433_n 0.00302413f $X=5.345 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A_M1016_g N_VPWR_c_433_n 0.00292189f $X=5.845 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A_M1016_g N_VPWR_c_434_n 7.14262e-19 $X=5.845 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A_M1017_g N_VPWR_c_434_n 0.0147378f $X=6.305 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A_M1018_g N_VPWR_c_434_n 0.0147154f $X=6.735 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A_M1025_g N_VPWR_c_434_n 7.51354e-19 $X=7.165 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A_c_290_n N_VPWR_c_434_n 4.53654e-19 $X=7.165 $Y=1.51 $X2=0 $Y2=0
cc_266 N_A_M1025_g N_VPWR_c_436_n 0.00739609f $X=7.165 $Y=2.465 $X2=0 $Y2=0
cc_267 N_A_M1002_g N_VPWR_c_442_n 0.00486043f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A_M1005_g N_VPWR_c_442_n 0.00585385f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A_M1007_g N_VPWR_c_443_n 0.00585385f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_270 N_A_M1011_g N_VPWR_c_443_n 0.00585385f $X=5.345 $Y=2.465 $X2=0 $Y2=0
cc_271 N_A_M1016_g N_VPWR_c_444_n 0.00585385f $X=5.845 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A_M1017_g N_VPWR_c_444_n 0.00486043f $X=6.305 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A_M1018_g N_VPWR_c_445_n 0.00486043f $X=6.735 $Y=2.465 $X2=0 $Y2=0
cc_274 N_A_M1025_g N_VPWR_c_445_n 0.00585385f $X=7.165 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A_M1002_g N_VPWR_c_424_n 0.00824727f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A_M1005_g N_VPWR_c_424_n 0.0106935f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A_M1007_g N_VPWR_c_424_n 0.0108646f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_278 N_A_M1011_g N_VPWR_c_424_n 0.0108646f $X=5.345 $Y=2.465 $X2=0 $Y2=0
cc_279 N_A_M1016_g N_VPWR_c_424_n 0.0107697f $X=5.845 $Y=2.465 $X2=0 $Y2=0
cc_280 N_A_M1017_g N_VPWR_c_424_n 0.00832343f $X=6.305 $Y=2.465 $X2=0 $Y2=0
cc_281 N_A_M1018_g N_VPWR_c_424_n 0.00824727f $X=6.735 $Y=2.465 $X2=0 $Y2=0
cc_282 N_A_M1025_g N_VPWR_c_424_n 0.011559f $X=7.165 $Y=2.465 $X2=0 $Y2=0
cc_283 N_A_M1002_g N_Y_c_563_n 0.0141566f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_284 N_A_M1002_g N_Y_c_564_n 0.00216819f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_285 N_A_M1005_g N_Y_c_564_n 0.00197868f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A_M1005_g N_Y_c_601_n 0.0156001f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A_M1007_g N_Y_c_601_n 0.0133867f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_288 N_A_c_287_n N_Y_c_601_n 9.5993e-19 $X=4.77 $Y=1.51 $X2=0 $Y2=0
cc_289 N_A_c_306_n N_Y_c_601_n 0.033867f $X=5.615 $Y=1.51 $X2=0 $Y2=0
cc_290 N_A_M1006_g N_Y_c_555_n 0.0114552f $X=4.345 $Y=0.745 $X2=0 $Y2=0
cc_291 N_A_M1009_g N_Y_c_555_n 0.013136f $X=4.845 $Y=0.745 $X2=0 $Y2=0
cc_292 N_A_c_287_n N_Y_c_555_n 0.00419003f $X=4.77 $Y=1.51 $X2=0 $Y2=0
cc_293 N_A_c_306_n N_Y_c_555_n 0.0395828f $X=5.615 $Y=1.51 $X2=0 $Y2=0
cc_294 N_A_M1013_g N_Y_c_609_n 0.00687129f $X=5.345 $Y=0.745 $X2=0 $Y2=0
cc_295 N_A_M1020_g N_Y_c_609_n 2.75259e-19 $X=5.845 $Y=0.745 $X2=0 $Y2=0
cc_296 N_A_M1011_g N_Y_c_611_n 0.0133867f $X=5.345 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A_M1016_g N_Y_c_611_n 0.0154521f $X=5.845 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A_c_289_n N_Y_c_611_n 9.5993e-19 $X=5.77 $Y=1.51 $X2=0 $Y2=0
cc_299 N_A_c_306_n N_Y_c_611_n 0.0349993f $X=5.615 $Y=1.51 $X2=0 $Y2=0
cc_300 N_A_M1013_g N_Y_c_556_n 0.00985868f $X=5.345 $Y=0.745 $X2=0 $Y2=0
cc_301 N_A_M1020_g N_Y_c_556_n 0.0152187f $X=5.845 $Y=0.745 $X2=0 $Y2=0
cc_302 N_A_c_289_n N_Y_c_556_n 0.00419585f $X=5.77 $Y=1.51 $X2=0 $Y2=0
cc_303 N_A_c_306_n N_Y_c_556_n 0.0360351f $X=5.615 $Y=1.51 $X2=0 $Y2=0
cc_304 N_A_M1023_g N_Y_c_619_n 5.49489e-19 $X=6.305 $Y=0.745 $X2=0 $Y2=0
cc_305 N_A_M1026_g N_Y_c_619_n 0.0072112f $X=6.735 $Y=0.745 $X2=0 $Y2=0
cc_306 N_A_M1027_g N_Y_c_619_n 0.00617693f $X=7.165 $Y=0.745 $X2=0 $Y2=0
cc_307 N_A_c_280_n N_Y_c_622_n 0.00108443f $X=5.27 $Y=1.51 $X2=0 $Y2=0
cc_308 N_A_c_306_n N_Y_c_622_n 0.0244204f $X=5.615 $Y=1.51 $X2=0 $Y2=0
cc_309 N_A_c_280_n N_Y_c_557_n 0.00435292f $X=5.27 $Y=1.51 $X2=0 $Y2=0
cc_310 N_A_M1013_g N_Y_c_557_n 0.00203406f $X=5.345 $Y=0.745 $X2=0 $Y2=0
cc_311 N_A_c_306_n N_Y_c_557_n 0.0276412f $X=5.615 $Y=1.51 $X2=0 $Y2=0
cc_312 N_A_M1020_g N_Y_c_558_n 0.00135012f $X=5.845 $Y=0.745 $X2=0 $Y2=0
cc_313 N_A_M1016_g N_Y_c_558_n 0.00322662f $X=5.845 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A_M1023_g N_Y_c_558_n 0.015082f $X=6.305 $Y=0.745 $X2=0 $Y2=0
cc_315 N_A_M1017_g N_Y_c_558_n 0.0147427f $X=6.305 $Y=2.465 $X2=0 $Y2=0
cc_316 N_A_M1026_g N_Y_c_558_n 0.0135304f $X=6.735 $Y=0.745 $X2=0 $Y2=0
cc_317 N_A_M1018_g N_Y_c_558_n 0.0146004f $X=6.735 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A_M1027_g N_Y_c_558_n 0.00976683f $X=7.165 $Y=0.745 $X2=0 $Y2=0
cc_319 N_A_M1025_g N_Y_c_558_n 0.0047211f $X=7.165 $Y=2.465 $X2=0 $Y2=0
cc_320 N_A_c_290_n N_Y_c_558_n 0.0761296f $X=7.165 $Y=1.51 $X2=0 $Y2=0
cc_321 N_A_c_306_n N_Y_c_558_n 0.0285236f $X=5.615 $Y=1.51 $X2=0 $Y2=0
cc_322 N_A_M1003_g Y 0.00288173f $X=3.915 $Y=0.745 $X2=0 $Y2=0
cc_323 N_A_M1006_g Y 0.00214025f $X=4.345 $Y=0.745 $X2=0 $Y2=0
cc_324 N_A_M1003_g N_Y_c_639_n 0.00526144f $X=3.915 $Y=0.745 $X2=0 $Y2=0
cc_325 N_A_M1006_g N_Y_c_639_n 0.00697334f $X=4.345 $Y=0.745 $X2=0 $Y2=0
cc_326 N_A_M1009_g N_Y_c_639_n 2.7525e-19 $X=4.845 $Y=0.745 $X2=0 $Y2=0
cc_327 N_A_M1003_g Y 0.0024675f $X=3.915 $Y=0.745 $X2=0 $Y2=0
cc_328 N_A_M1002_g Y 0.0027479f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_329 N_A_M1006_g Y 0.00249892f $X=4.345 $Y=0.745 $X2=0 $Y2=0
cc_330 N_A_M1005_g Y 0.00109995f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_331 N_A_c_286_n Y 0.0262248f $X=4.42 $Y=1.51 $X2=0 $Y2=0
cc_332 N_A_c_306_n Y 0.0270828f $X=5.615 $Y=1.51 $X2=0 $Y2=0
cc_333 N_A_M1003_g N_A_27_65#_c_717_n 6.54275e-19 $X=3.915 $Y=0.745 $X2=0 $Y2=0
cc_334 N_A_M1003_g N_A_27_65#_c_718_n 0.0118056f $X=3.915 $Y=0.745 $X2=0 $Y2=0
cc_335 N_A_M1006_g N_A_27_65#_c_718_n 0.0115919f $X=4.345 $Y=0.745 $X2=0 $Y2=0
cc_336 N_A_M1009_g N_A_27_65#_c_763_n 0.00697842f $X=4.845 $Y=0.745 $X2=0 $Y2=0
cc_337 N_A_M1013_g N_A_27_65#_c_763_n 3.22114e-19 $X=5.345 $Y=0.745 $X2=0 $Y2=0
cc_338 N_A_M1009_g N_A_27_65#_c_720_n 0.00869988f $X=4.845 $Y=0.745 $X2=0 $Y2=0
cc_339 N_A_M1013_g N_A_27_65#_c_720_n 0.0120041f $X=5.345 $Y=0.745 $X2=0 $Y2=0
cc_340 N_A_M1020_g N_A_27_65#_c_767_n 0.00652982f $X=5.845 $Y=0.745 $X2=0 $Y2=0
cc_341 N_A_M1023_g N_A_27_65#_c_767_n 5.95627e-19 $X=6.305 $Y=0.745 $X2=0 $Y2=0
cc_342 N_A_M1020_g N_A_27_65#_c_721_n 0.00868531f $X=5.845 $Y=0.745 $X2=0 $Y2=0
cc_343 N_A_M1023_g N_A_27_65#_c_721_n 0.0132133f $X=6.305 $Y=0.745 $X2=0 $Y2=0
cc_344 N_A_c_290_n N_A_27_65#_c_771_n 5.08933e-19 $X=7.165 $Y=1.51 $X2=0 $Y2=0
cc_345 N_A_M1026_g N_A_27_65#_c_722_n 0.0122849f $X=6.735 $Y=0.745 $X2=0 $Y2=0
cc_346 N_A_M1027_g N_A_27_65#_c_722_n 0.0128465f $X=7.165 $Y=0.745 $X2=0 $Y2=0
cc_347 N_A_M1027_g N_A_27_65#_c_723_n 0.00365765f $X=7.165 $Y=0.745 $X2=0 $Y2=0
cc_348 N_A_M1009_g N_A_27_65#_c_727_n 0.00152703f $X=4.845 $Y=0.745 $X2=0 $Y2=0
cc_349 N_A_M1020_g N_A_27_65#_c_728_n 0.00154963f $X=5.845 $Y=0.745 $X2=0 $Y2=0
cc_350 N_A_M1003_g N_VGND_c_845_n 5.15399e-19 $X=3.915 $Y=0.745 $X2=0 $Y2=0
cc_351 N_A_M1003_g N_VGND_c_851_n 0.00302501f $X=3.915 $Y=0.745 $X2=0 $Y2=0
cc_352 N_A_M1006_g N_VGND_c_851_n 0.00302501f $X=4.345 $Y=0.745 $X2=0 $Y2=0
cc_353 N_A_M1009_g N_VGND_c_851_n 0.00302473f $X=4.845 $Y=0.745 $X2=0 $Y2=0
cc_354 N_A_M1013_g N_VGND_c_851_n 0.00302501f $X=5.345 $Y=0.745 $X2=0 $Y2=0
cc_355 N_A_M1020_g N_VGND_c_851_n 0.00302473f $X=5.845 $Y=0.745 $X2=0 $Y2=0
cc_356 N_A_M1023_g N_VGND_c_851_n 0.00302501f $X=6.305 $Y=0.745 $X2=0 $Y2=0
cc_357 N_A_M1026_g N_VGND_c_851_n 0.00302501f $X=6.735 $Y=0.745 $X2=0 $Y2=0
cc_358 N_A_M1027_g N_VGND_c_851_n 0.00302501f $X=7.165 $Y=0.745 $X2=0 $Y2=0
cc_359 N_A_M1003_g N_VGND_c_852_n 0.00435646f $X=3.915 $Y=0.745 $X2=0 $Y2=0
cc_360 N_A_M1006_g N_VGND_c_852_n 0.00441253f $X=4.345 $Y=0.745 $X2=0 $Y2=0
cc_361 N_A_M1009_g N_VGND_c_852_n 0.00447833f $X=4.845 $Y=0.745 $X2=0 $Y2=0
cc_362 N_A_M1013_g N_VGND_c_852_n 0.00447835f $X=5.345 $Y=0.745 $X2=0 $Y2=0
cc_363 N_A_M1020_g N_VGND_c_852_n 0.00444181f $X=5.845 $Y=0.745 $X2=0 $Y2=0
cc_364 N_A_M1023_g N_VGND_c_852_n 0.00437601f $X=6.305 $Y=0.745 $X2=0 $Y2=0
cc_365 N_A_M1026_g N_VGND_c_852_n 0.00434671f $X=6.735 $Y=0.745 $X2=0 $Y2=0
cc_366 N_A_M1027_g N_VGND_c_852_n 0.00471914f $X=7.165 $Y=0.745 $X2=0 $Y2=0
cc_367 N_VPWR_c_424_n N_Y_M1000_d 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_368 N_VPWR_c_424_n N_Y_M1010_d 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_369 N_VPWR_c_424_n N_Y_M1021_d 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_370 N_VPWR_c_424_n N_Y_M1028_d 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_371 N_VPWR_c_424_n N_Y_M1002_s 0.0041489f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_372 N_VPWR_c_424_n N_Y_M1007_s 0.00349426f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_373 N_VPWR_c_424_n N_Y_M1016_s 0.0050859f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_374 N_VPWR_c_424_n N_Y_M1018_s 0.00501859f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_375 N_VPWR_c_441_n N_Y_c_656_n 0.0124525f $X=0.955 $Y=3.33 $X2=0 $Y2=0
cc_376 N_VPWR_c_424_n N_Y_c_656_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_377 N_VPWR_M1004_s N_Y_c_560_n 0.00176461f $X=0.98 $Y=1.835 $X2=0 $Y2=0
cc_378 N_VPWR_c_427_n N_Y_c_560_n 0.0170777f $X=1.12 $Y=2.19 $X2=0 $Y2=0
cc_379 N_VPWR_c_426_n N_Y_c_561_n 0.00498824f $X=0.26 $Y=1.985 $X2=0 $Y2=0
cc_380 N_VPWR_c_437_n N_Y_c_661_n 0.0124525f $X=1.815 $Y=3.33 $X2=0 $Y2=0
cc_381 N_VPWR_c_424_n N_Y_c_661_n 0.00729316f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_382 N_VPWR_M1015_s N_Y_c_578_n 0.00333177f $X=1.84 $Y=1.835 $X2=0 $Y2=0
cc_383 N_VPWR_c_428_n N_Y_c_578_n 0.0170777f $X=1.98 $Y=2.355 $X2=0 $Y2=0
cc_384 N_VPWR_c_439_n N_Y_c_665_n 0.0124525f $X=2.675 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_c_424_n N_Y_c_665_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_M1022_s N_Y_c_583_n 0.00362809f $X=2.7 $Y=1.835 $X2=0 $Y2=0
cc_387 N_VPWR_c_429_n N_Y_c_583_n 0.0170777f $X=2.84 $Y=2.355 $X2=0 $Y2=0
cc_388 N_VPWR_c_430_n N_Y_c_669_n 0.0124525f $X=3.535 $Y=3.33 $X2=0 $Y2=0
cc_389 N_VPWR_c_424_n N_Y_c_669_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_390 N_VPWR_M1030_s N_Y_c_563_n 0.00176461f $X=3.56 $Y=1.835 $X2=0 $Y2=0
cc_391 N_VPWR_c_431_n N_Y_c_563_n 0.0170777f $X=3.7 $Y=2.2 $X2=0 $Y2=0
cc_392 N_VPWR_c_442_n N_Y_c_673_n 0.0136943f $X=4.43 $Y=3.33 $X2=0 $Y2=0
cc_393 N_VPWR_c_424_n N_Y_c_673_n 0.00866972f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_394 N_VPWR_M1005_d N_Y_c_601_n 0.00468059f $X=4.42 $Y=1.835 $X2=0 $Y2=0
cc_395 N_VPWR_c_432_n N_Y_c_601_n 0.0192006f $X=4.595 $Y=2.355 $X2=0 $Y2=0
cc_396 N_VPWR_c_443_n N_Y_c_677_n 0.019858f $X=5.43 $Y=3.33 $X2=0 $Y2=0
cc_397 N_VPWR_c_424_n N_Y_c_677_n 0.0127519f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_398 N_VPWR_M1011_d N_Y_c_611_n 0.00468059f $X=5.42 $Y=1.835 $X2=0 $Y2=0
cc_399 N_VPWR_c_433_n N_Y_c_611_n 0.0192006f $X=5.595 $Y=2.355 $X2=0 $Y2=0
cc_400 N_VPWR_c_444_n N_Y_c_681_n 0.0150941f $X=6.355 $Y=3.33 $X2=0 $Y2=0
cc_401 N_VPWR_c_424_n N_Y_c_681_n 0.0090585f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_402 N_VPWR_c_445_n N_Y_c_683_n 0.0128073f $X=7.275 $Y=3.33 $X2=0 $Y2=0
cc_403 N_VPWR_c_424_n N_Y_c_683_n 0.00769778f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_404 N_VPWR_M1017_d N_Y_c_558_n 0.001837f $X=6.38 $Y=1.835 $X2=0 $Y2=0
cc_405 N_VPWR_c_434_n N_Y_c_558_n 0.0189454f $X=6.52 $Y=2.18 $X2=0 $Y2=0
cc_406 N_VPWR_c_436_n N_Y_c_558_n 0.00135635f $X=7.38 $Y=1.98 $X2=0 $Y2=0
cc_407 N_VPWR_c_426_n N_A_27_65#_c_710_n 0.00227786f $X=0.26 $Y=1.985 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_426_n N_A_27_65#_c_711_n 0.0103538f $X=0.26 $Y=1.985 $X2=0 $Y2=0
cc_409 N_VPWR_c_436_n N_A_27_65#_c_723_n 0.00744828f $X=7.38 $Y=1.98 $X2=0 $Y2=0
cc_410 N_Y_c_555_n N_A_27_65#_M1006_s 0.00250873f $X=4.965 $Y=1.17 $X2=0 $Y2=0
cc_411 N_Y_c_556_n N_A_27_65#_M1013_s 0.00251316f $X=5.95 $Y=1.165 $X2=0 $Y2=0
cc_412 N_Y_c_558_n N_A_27_65#_M1023_s 0.001837f $X=6.95 $Y=1.587 $X2=0 $Y2=0
cc_413 N_Y_c_563_n N_A_27_65#_c_717_n 0.0102738f $X=3.965 $Y=1.86 $X2=0 $Y2=0
cc_414 Y N_A_27_65#_c_717_n 0.0104705f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_415 N_Y_M1003_d N_A_27_65#_c_718_n 0.00176461f $X=3.99 $Y=0.325 $X2=0 $Y2=0
cc_416 N_Y_c_555_n N_A_27_65#_c_718_n 0.00272017f $X=4.965 $Y=1.17 $X2=0 $Y2=0
cc_417 N_Y_c_639_n N_A_27_65#_c_718_n 0.0159766f $X=4.13 $Y=0.7 $X2=0 $Y2=0
cc_418 N_Y_c_555_n N_A_27_65#_c_763_n 0.0209355f $X=4.965 $Y=1.17 $X2=0 $Y2=0
cc_419 N_Y_M1009_d N_A_27_65#_c_720_n 0.00250873f $X=4.92 $Y=0.325 $X2=0 $Y2=0
cc_420 N_Y_c_555_n N_A_27_65#_c_720_n 0.00272017f $X=4.965 $Y=1.17 $X2=0 $Y2=0
cc_421 N_Y_c_609_n N_A_27_65#_c_720_n 0.0195903f $X=5.13 $Y=0.7 $X2=0 $Y2=0
cc_422 N_Y_c_556_n N_A_27_65#_c_720_n 0.00277195f $X=5.95 $Y=1.165 $X2=0 $Y2=0
cc_423 N_Y_c_556_n N_A_27_65#_c_767_n 0.0209908f $X=5.95 $Y=1.165 $X2=0 $Y2=0
cc_424 N_Y_M1020_d N_A_27_65#_c_721_n 0.0020872f $X=5.92 $Y=0.325 $X2=0 $Y2=0
cc_425 N_Y_c_556_n N_A_27_65#_c_721_n 0.00282518f $X=5.95 $Y=1.165 $X2=0 $Y2=0
cc_426 N_Y_c_704_p N_A_27_65#_c_721_n 0.0150119f $X=6.09 $Y=0.805 $X2=0 $Y2=0
cc_427 N_Y_c_558_n N_A_27_65#_c_771_n 0.0149668f $X=6.95 $Y=1.587 $X2=0 $Y2=0
cc_428 N_Y_M1026_d N_A_27_65#_c_722_n 0.00176773f $X=6.81 $Y=0.325 $X2=0 $Y2=0
cc_429 N_Y_c_619_n N_A_27_65#_c_722_n 0.0160814f $X=6.95 $Y=0.7 $X2=0 $Y2=0
cc_430 N_Y_c_558_n N_A_27_65#_c_723_n 0.00244151f $X=6.95 $Y=1.587 $X2=0 $Y2=0
cc_431 N_A_27_65#_c_710_n N_VGND_M1001_s 0.00176461f $X=1.025 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_432 N_A_27_65#_c_713_n N_VGND_M1012_s 0.00176461f $X=1.885 $Y=1.16 $X2=0
+ $Y2=0
cc_433 N_A_27_65#_c_715_n N_VGND_M1019_s 0.00176461f $X=2.745 $Y=1.16 $X2=0
+ $Y2=0
cc_434 N_A_27_65#_c_717_n N_VGND_M1029_s 0.00176461f $X=3.605 $Y=1.16 $X2=0
+ $Y2=0
cc_435 N_A_27_65#_c_709_n N_VGND_c_841_n 0.0232759f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_436 N_A_27_65#_c_710_n N_VGND_c_841_n 0.0170777f $X=1.025 $Y=1.16 $X2=0 $Y2=0
cc_437 N_A_27_65#_c_712_n N_VGND_c_841_n 0.0232345f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_438 N_A_27_65#_c_712_n N_VGND_c_842_n 0.0221973f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_439 N_A_27_65#_c_713_n N_VGND_c_842_n 0.0170777f $X=1.885 $Y=1.16 $X2=0 $Y2=0
cc_440 N_A_27_65#_c_714_n N_VGND_c_842_n 0.0232405f $X=1.98 $Y=0.47 $X2=0 $Y2=0
cc_441 N_A_27_65#_c_714_n N_VGND_c_843_n 0.0232405f $X=1.98 $Y=0.47 $X2=0 $Y2=0
cc_442 N_A_27_65#_c_715_n N_VGND_c_843_n 0.0170777f $X=2.745 $Y=1.16 $X2=0 $Y2=0
cc_443 N_A_27_65#_c_716_n N_VGND_c_843_n 0.0232405f $X=2.84 $Y=0.47 $X2=0 $Y2=0
cc_444 N_A_27_65#_c_716_n N_VGND_c_844_n 0.0102275f $X=2.84 $Y=0.47 $X2=0 $Y2=0
cc_445 N_A_27_65#_c_716_n N_VGND_c_845_n 0.0232405f $X=2.84 $Y=0.47 $X2=0 $Y2=0
cc_446 N_A_27_65#_c_717_n N_VGND_c_845_n 0.0170777f $X=3.605 $Y=1.16 $X2=0 $Y2=0
cc_447 N_A_27_65#_c_719_n N_VGND_c_845_n 0.00962585f $X=3.795 $Y=0.34 $X2=0
+ $Y2=0
cc_448 N_A_27_65#_c_712_n N_VGND_c_846_n 0.0096835f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_449 N_A_27_65#_c_714_n N_VGND_c_848_n 0.0102275f $X=1.98 $Y=0.47 $X2=0 $Y2=0
cc_450 N_A_27_65#_c_709_n N_VGND_c_850_n 0.0140356f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_451 N_A_27_65#_c_718_n N_VGND_c_851_n 0.0422287f $X=4.465 $Y=0.34 $X2=0 $Y2=0
cc_452 N_A_27_65#_c_719_n N_VGND_c_851_n 0.0136205f $X=3.795 $Y=0.34 $X2=0 $Y2=0
cc_453 N_A_27_65#_c_720_n N_VGND_c_851_n 0.0423044f $X=5.465 $Y=0.34 $X2=0 $Y2=0
cc_454 N_A_27_65#_c_721_n N_VGND_c_851_n 0.0376177f $X=6.39 $Y=0.345 $X2=0 $Y2=0
cc_455 N_A_27_65#_c_722_n N_VGND_c_851_n 0.0610304f $X=7.285 $Y=0.345 $X2=0
+ $Y2=0
cc_456 N_A_27_65#_c_727_n N_VGND_c_851_n 0.0235159f $X=4.63 $Y=0.34 $X2=0 $Y2=0
cc_457 N_A_27_65#_c_728_n N_VGND_c_851_n 0.023489f $X=5.63 $Y=0.345 $X2=0 $Y2=0
cc_458 N_A_27_65#_c_729_n N_VGND_c_851_n 0.0161295f $X=6.502 $Y=0.345 $X2=0
+ $Y2=0
cc_459 N_A_27_65#_c_709_n N_VGND_c_852_n 0.00977851f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_460 N_A_27_65#_c_712_n N_VGND_c_852_n 0.00674642f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_461 N_A_27_65#_c_714_n N_VGND_c_852_n 0.00712543f $X=1.98 $Y=0.47 $X2=0 $Y2=0
cc_462 N_A_27_65#_c_716_n N_VGND_c_852_n 0.00712543f $X=2.84 $Y=0.47 $X2=0 $Y2=0
cc_463 N_A_27_65#_c_718_n N_VGND_c_852_n 0.0238173f $X=4.465 $Y=0.34 $X2=0 $Y2=0
cc_464 N_A_27_65#_c_719_n N_VGND_c_852_n 0.00738676f $X=3.795 $Y=0.34 $X2=0
+ $Y2=0
cc_465 N_A_27_65#_c_720_n N_VGND_c_852_n 0.0239316f $X=5.465 $Y=0.34 $X2=0 $Y2=0
cc_466 N_A_27_65#_c_721_n N_VGND_c_852_n 0.0211384f $X=6.39 $Y=0.345 $X2=0 $Y2=0
cc_467 N_A_27_65#_c_722_n N_VGND_c_852_n 0.0339555f $X=7.285 $Y=0.345 $X2=0
+ $Y2=0
cc_468 N_A_27_65#_c_727_n N_VGND_c_852_n 0.0127052f $X=4.63 $Y=0.34 $X2=0 $Y2=0
cc_469 N_A_27_65#_c_728_n N_VGND_c_852_n 0.0127001f $X=5.63 $Y=0.345 $X2=0 $Y2=0
cc_470 N_A_27_65#_c_729_n N_VGND_c_852_n 0.00874748f $X=6.502 $Y=0.345 $X2=0
+ $Y2=0
