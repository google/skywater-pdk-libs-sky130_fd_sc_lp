* File: sky130_fd_sc_lp__dlxtp_1.spice
* Created: Wed Sep  2 09:48:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxtp_1.pex.spice"
.subckt sky130_fd_sc_lp__dlxtp_1  VNB VPB D GATE VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_D_M1008_g N_A_27_425#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_196_425#_M1009_d N_GATE_M1009_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_196_425#_M1001_g N_A_317_461#_M1001_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1003 A_530_125# N_A_27_425#_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1017 N_A_596_419#_M1017_d N_A_317_461#_M1017_g A_530_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.06195 AS=0.0441 PD=0.715 PS=0.63 NRD=4.284 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 A_691_125# N_A_196_425#_M1005_g N_A_596_419#_M1017_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.06195 PD=0.63 PS=0.715 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75001.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_733_99#_M1002_g A_691_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0917 AS=0.0441 PD=0.82 PS=0.63 NRD=46.656 NRS=14.28 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_A_733_99#_M1016_d N_A_596_419#_M1016_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1834 PD=2.21 PS=1.64 NRD=0 NRS=0 M=1 R=5.6 SA=75001.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1014 N_Q_M1014_d N_A_733_99#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_VPWR_M1007_d N_D_M1007_g N_A_27_425#_M1007_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1015 N_A_196_425#_M1015_d N_GATE_M1015_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_196_425#_M1000_g N_A_317_461#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.17665 AS=0.1696 PD=1.32 PS=1.81 NRD=29.2348 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1010 A_524_419# N_A_27_425#_M1010_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.17665 PD=0.85 PS=1.32 NRD=15.3857 NRS=30.7714 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1012 N_A_596_419#_M1012_d N_A_196_425#_M1012_g A_524_419# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.130294 AS=0.0672 PD=1.22566 PS=0.85 NRD=9.2196 NRS=15.3857 M=1
+ R=4.26667 SA=75001 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 A_701_419# N_A_317_461#_M1004_g N_A_596_419#_M1012_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0855057 PD=0.63 PS=0.80434 NRD=23.443 NRS=31.6579 M=1
+ R=2.8 SA=75001.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_733_99#_M1006_g A_701_419# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.101325 AS=0.0441 PD=0.8275 PS=0.63 NRD=56.2829 NRS=23.443 M=1 R=2.8
+ SA=75001.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_A_733_99#_M1013_d N_A_596_419#_M1013_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.303975 PD=3.05 PS=2.4825 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.9 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1011 N_Q_M1011_d N_A_733_99#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.6751 P=16.33
c_723 A_524_419# 0 1.64722e-19 $X=2.62 $Y=2.095
*
.include "sky130_fd_sc_lp__dlxtp_1.pxi.spice"
*
.ends
*
*
