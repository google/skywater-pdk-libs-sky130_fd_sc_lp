* File: sky130_fd_sc_lp__nor3b_m.spice
* Created: Fri Aug 28 10:56:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor3b_m.pex.spice"
.subckt sky130_fd_sc_lp__nor3b_m  VNB VPB C_N A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_C_N_M1003_g N_A_27_439#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.1 A=0.063
+ P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_27_439#_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_C_N_M1005_g N_A_27_439#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=32.8202 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1000 A_218_439# N_A_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=18.7544 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_290_439# N_B_M1001_g A_218_439# VPB PHIGHVT L=0.15 W=0.42 AD=0.0777
+ AS=0.0441 PD=0.79 PS=0.63 NRD=60.9715 NRS=23.443 M=1 R=2.8 SA=75001.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_A_27_439#_M1007_g A_290_439# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0777 PD=1.37 PS=0.79 NRD=0 NRS=60.9715 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
c_60 VPB 0 1.55344e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__nor3b_m.pxi.spice"
*
.ends
*
*
