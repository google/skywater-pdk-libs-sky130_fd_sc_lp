* File: sky130_fd_sc_lp__a221oi_2.pxi.spice
* Created: Wed Sep  2 09:21:55 2020
* 
x_PM_SKY130_FD_SC_LP__A221OI_2%C1 N_C1_M1005_g N_C1_M1003_g N_C1_M1018_g
+ N_C1_M1007_g C1 C1 N_C1_c_95_n PM_SKY130_FD_SC_LP__A221OI_2%C1
x_PM_SKY130_FD_SC_LP__A221OI_2%B2 N_B2_M1004_g N_B2_M1014_g N_B2_M1010_g
+ N_B2_M1017_g N_B2_c_133_n N_B2_c_134_n N_B2_c_135_n B2 B2 B2 N_B2_c_137_n
+ N_B2_c_138_n PM_SKY130_FD_SC_LP__A221OI_2%B2
x_PM_SKY130_FD_SC_LP__A221OI_2%B1 N_B1_c_213_n N_B1_M1002_g N_B1_M1000_g
+ N_B1_c_215_n N_B1_M1013_g N_B1_M1006_g B1 N_B1_c_218_n
+ PM_SKY130_FD_SC_LP__A221OI_2%B1
x_PM_SKY130_FD_SC_LP__A221OI_2%A2 N_A2_M1012_g N_A2_M1011_g N_A2_M1015_g
+ N_A2_M1016_g N_A2_c_268_n N_A2_c_269_n N_A2_c_270_n N_A2_c_271_n A2 A2
+ N_A2_c_273_n N_A2_c_274_n PM_SKY130_FD_SC_LP__A221OI_2%A2
x_PM_SKY130_FD_SC_LP__A221OI_2%A1 N_A1_c_342_n N_A1_M1001_g N_A1_M1009_g
+ N_A1_c_344_n N_A1_M1008_g N_A1_M1019_g A1 A1 A1 N_A1_c_347_n
+ PM_SKY130_FD_SC_LP__A221OI_2%A1
x_PM_SKY130_FD_SC_LP__A221OI_2%A_27_367# N_A_27_367#_M1005_d N_A_27_367#_M1018_d
+ N_A_27_367#_M1014_s N_A_27_367#_M1006_d N_A_27_367#_c_394_n
+ N_A_27_367#_c_395_n N_A_27_367#_c_401_n N_A_27_367#_c_396_n
+ N_A_27_367#_c_397_n N_A_27_367#_c_398_n N_A_27_367#_c_408_n
+ N_A_27_367#_c_409_n N_A_27_367#_c_412_n PM_SKY130_FD_SC_LP__A221OI_2%A_27_367#
x_PM_SKY130_FD_SC_LP__A221OI_2%Y N_Y_M1003_d N_Y_M1002_s N_Y_M1001_d N_Y_M1005_s
+ N_Y_c_469_n N_Y_c_446_n Y Y Y Y Y Y PM_SKY130_FD_SC_LP__A221OI_2%Y
x_PM_SKY130_FD_SC_LP__A221OI_2%A_303_367# N_A_303_367#_M1014_d
+ N_A_303_367#_M1000_s N_A_303_367#_M1017_d N_A_303_367#_M1009_s
+ N_A_303_367#_M1016_s N_A_303_367#_c_499_n N_A_303_367#_c_503_n
+ N_A_303_367#_c_500_n N_A_303_367#_c_535_n N_A_303_367#_c_504_n
+ N_A_303_367#_c_505_n N_A_303_367#_c_511_n N_A_303_367#_c_512_n
+ N_A_303_367#_c_516_n N_A_303_367#_c_517_n N_A_303_367#_c_501_n
+ N_A_303_367#_c_502_n N_A_303_367#_c_546_p N_A_303_367#_c_522_n
+ PM_SKY130_FD_SC_LP__A221OI_2%A_303_367#
x_PM_SKY130_FD_SC_LP__A221OI_2%VPWR N_VPWR_M1012_d N_VPWR_M1019_d N_VPWR_c_562_n
+ N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n
+ VPWR N_VPWR_c_568_n N_VPWR_c_561_n PM_SKY130_FD_SC_LP__A221OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A221OI_2%VGND N_VGND_M1003_s N_VGND_M1007_s N_VGND_M1010_s
+ N_VGND_M1015_s N_VGND_c_629_n N_VGND_c_630_n N_VGND_c_631_n N_VGND_c_632_n
+ N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n VGND
+ N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n N_VGND_c_640_n
+ PM_SKY130_FD_SC_LP__A221OI_2%VGND
x_PM_SKY130_FD_SC_LP__A221OI_2%A_384_47# N_A_384_47#_M1004_d N_A_384_47#_M1013_d
+ N_A_384_47#_c_696_n PM_SKY130_FD_SC_LP__A221OI_2%A_384_47#
x_PM_SKY130_FD_SC_LP__A221OI_2%A_760_47# N_A_760_47#_M1011_d N_A_760_47#_M1008_s
+ N_A_760_47#_c_707_n N_A_760_47#_c_708_n PM_SKY130_FD_SC_LP__A221OI_2%A_760_47#
cc_1 VNB N_C1_M1005_g 0.00703667f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB N_C1_M1003_g 0.023517f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.655
cc_3 VNB N_C1_M1018_g 0.00663591f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_4 VNB N_C1_M1007_g 0.0204108f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_5 VNB C1 0.0239943f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_C1_c_95_n 0.0741165f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.375
cc_7 VNB N_B2_M1004_g 0.0297723f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_8 VNB N_B2_M1010_g 0.024557f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_9 VNB N_B2_M1017_g 0.00128182f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_10 VNB N_B2_c_133_n 0.00582227f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_B2_c_134_n 2.57777e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B2_c_135_n 0.0324368f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_13 VNB B2 0.0141217f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.21
cc_14 VNB N_B2_c_137_n 0.0273161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_c_138_n 0.00162148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_213_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.54
cc_17 VNB N_B1_M1000_g 0.00596194f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.655
cc_18 VNB N_B1_c_215_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_M1006_g 0.00656831f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.21
cc_20 VNB B1 0.00279127f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_21 VNB N_B1_c_218_n 0.035642f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_22 VNB N_A2_M1011_g 0.0273283f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.655
cc_23 VNB N_A2_M1015_g 0.0243742f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_24 VNB N_A2_M1016_g 0.00662156f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_25 VNB N_A2_c_268_n 0.0102773f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_A2_c_269_n 0.0092694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A2_c_270_n 0.0012749f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_28 VNB N_A2_c_271_n 0.0260105f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_29 VNB A2 0.0276458f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.21
cc_30 VNB N_A2_c_273_n 0.0601928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_c_274_n 0.0016291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_c_342_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.54
cc_33 VNB N_A1_M1009_g 0.00650355f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.655
cc_34 VNB N_A1_c_344_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A1_M1019_g 0.00689546f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.21
cc_36 VNB A1 0.00948948f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_37 VNB N_A1_c_347_n 0.0345757f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.375
cc_38 VNB Y 0.00195071f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_39 VNB N_VPWR_c_561_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_629_n 0.0137379f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.21
cc_41 VNB N_VGND_c_630_n 0.034876f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.655
cc_42 VNB N_VGND_c_631_n 0.00561153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_632_n 0.0354775f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.375
cc_44 VNB N_VGND_c_633_n 0.0361336f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.375
cc_45 VNB N_VGND_c_634_n 0.00632255f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.21
cc_46 VNB N_VGND_c_635_n 0.0374415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_636_n 0.00499734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_637_n 0.0137583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_638_n 0.302923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_639_n 0.0154252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_640_n 0.0135337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_C1_M1005_g 0.0259883f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_53 VPB N_C1_M1018_g 0.0238463f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_54 VPB C1 0.00840075f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_55 VPB N_B2_M1014_g 0.0238089f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.655
cc_56 VPB N_B2_M1017_g 0.019473f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.655
cc_57 VPB N_B2_c_133_n 0.00473954f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_58 VPB N_B2_c_134_n 0.00406744f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB B2 0.0112491f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.21
cc_60 VPB N_B2_c_137_n 0.00652892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_B2_c_138_n 0.00125388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_B1_M1000_g 0.0188332f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.655
cc_63 VPB N_B1_M1006_g 0.0188867f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.21
cc_64 VPB N_A2_M1012_g 0.0202658f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_65 VPB N_A2_M1016_g 0.0247824f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.655
cc_66 VPB N_A2_c_269_n 0.0104001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A2_c_270_n 0.00114697f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.375
cc_68 VPB N_A2_c_271_n 0.00643251f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.375
cc_69 VPB N_A2_c_274_n 0.0177967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A1_M1009_g 0.019965f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.655
cc_71 VPB N_A1_M1019_g 0.0186439f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.21
cc_72 VPB N_A_27_367#_c_394_n 0.00746637f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.21
cc_73 VPB N_A_27_367#_c_395_n 0.0372165f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.655
cc_74 VPB N_A_27_367#_c_396_n 6.27129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_27_367#_c_397_n 0.00924297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_27_367#_c_398_n 0.0104114f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.375
cc_77 VPB Y 0.00136044f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.375
cc_78 VPB N_A_303_367#_c_499_n 0.00578576f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_79 VPB N_A_303_367#_c_500_n 0.00181169f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.375
cc_80 VPB N_A_303_367#_c_501_n 0.00745496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_303_367#_c_502_n 0.0358372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_562_n 0.00489487f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.54
cc_83 VPB N_VPWR_c_563_n 4.08532e-19 $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.21
cc_84 VPB N_VPWR_c_564_n 0.0889083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_565_n 0.00631455f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_86 VPB N_VPWR_c_566_n 0.0151943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_567_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_568_n 0.0240619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_561_n 0.0650598f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 N_C1_M1007_g N_B2_M1004_g 0.0140344f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_91 N_C1_c_95_n B2 0.00834781f $X=0.905 $Y=1.375 $X2=0 $Y2=0
cc_92 N_C1_c_95_n N_B2_c_137_n 0.00471508f $X=0.905 $Y=1.375 $X2=0 $Y2=0
cc_93 C1 N_A_27_367#_c_395_n 0.0223998f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_94 N_C1_c_95_n N_A_27_367#_c_395_n 7.07743e-19 $X=0.905 $Y=1.375 $X2=0 $Y2=0
cc_95 N_C1_M1005_g N_A_27_367#_c_401_n 0.0115031f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_96 N_C1_M1018_g N_A_27_367#_c_401_n 0.0115031f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_97 N_C1_M1007_g N_Y_c_446_n 0.0171244f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_98 N_C1_M1003_g Y 0.00621455f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_99 N_C1_M1003_g Y 0.00290792f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_100 N_C1_M1005_g Y 0.00515594f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_101 N_C1_M1003_g Y 0.00839382f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_102 N_C1_M1018_g Y 0.010675f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_103 N_C1_M1007_g Y 0.00407991f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_104 C1 Y 0.0405192f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_105 N_C1_c_95_n Y 0.0260106f $X=0.905 $Y=1.375 $X2=0 $Y2=0
cc_106 N_C1_M1005_g Y 0.0129453f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_107 N_C1_M1018_g Y 0.0127275f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_108 N_C1_M1005_g N_VPWR_c_564_n 0.00357877f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_109 N_C1_M1018_g N_VPWR_c_564_n 0.00357877f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_110 N_C1_M1005_g N_VPWR_c_561_n 0.00628381f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_111 N_C1_M1018_g N_VPWR_c_561_n 0.00665089f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_112 N_C1_M1003_g N_VGND_c_630_n 0.00521771f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_113 C1 N_VGND_c_630_n 0.0217463f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_114 N_C1_c_95_n N_VGND_c_630_n 0.00200262f $X=0.905 $Y=1.375 $X2=0 $Y2=0
cc_115 N_C1_M1003_g N_VGND_c_638_n 0.0108577f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_116 N_C1_M1007_g N_VGND_c_638_n 0.00448563f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_117 N_C1_M1003_g N_VGND_c_639_n 0.0054895f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_118 N_C1_M1007_g N_VGND_c_639_n 0.00486043f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_119 N_C1_M1003_g N_VGND_c_640_n 6.53151e-19 $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_120 N_C1_M1007_g N_VGND_c_640_n 0.0105049f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_121 N_B2_M1004_g N_B1_c_213_n 0.0419007f $X=1.845 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_122 N_B2_M1014_g N_B1_M1000_g 0.0355433f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B2_c_133_n N_B1_M1000_g 0.00780467f $X=3 $Y=1.7 $X2=0 $Y2=0
cc_124 N_B2_c_137_n N_B1_M1000_g 0.0097295f $X=1.825 $Y=1.51 $X2=0 $Y2=0
cc_125 N_B2_c_138_n N_B1_M1000_g 0.00622553f $X=2.255 $Y=1.605 $X2=0 $Y2=0
cc_126 N_B2_M1010_g N_B1_c_215_n 0.0383765f $X=3.135 $Y=0.655 $X2=0 $Y2=0
cc_127 N_B2_M1017_g N_B1_M1006_g 0.0377913f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_128 N_B2_c_133_n N_B1_M1006_g 0.00995412f $X=3 $Y=1.7 $X2=0 $Y2=0
cc_129 N_B2_c_138_n N_B1_M1006_g 4.96805e-19 $X=2.255 $Y=1.605 $X2=0 $Y2=0
cc_130 N_B2_M1004_g B1 5.47394e-19 $X=1.845 $Y=0.655 $X2=0 $Y2=0
cc_131 N_B2_M1010_g B1 0.00188886f $X=3.135 $Y=0.655 $X2=0 $Y2=0
cc_132 N_B2_c_133_n B1 0.0281021f $X=3 $Y=1.7 $X2=0 $Y2=0
cc_133 N_B2_c_134_n B1 0.00526935f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_134 N_B2_c_135_n B1 0.00230469f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_135 N_B2_c_137_n B1 3.70015e-19 $X=1.825 $Y=1.51 $X2=0 $Y2=0
cc_136 N_B2_c_138_n B1 0.00153522f $X=2.255 $Y=1.605 $X2=0 $Y2=0
cc_137 N_B2_c_133_n N_B1_c_218_n 0.00247657f $X=3 $Y=1.7 $X2=0 $Y2=0
cc_138 N_B2_c_134_n N_B1_c_218_n 0.00128179f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_139 N_B2_c_135_n N_B1_c_218_n 0.0211428f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_140 N_B2_c_137_n N_B1_c_218_n 0.0117496f $X=1.825 $Y=1.51 $X2=0 $Y2=0
cc_141 N_B2_c_138_n N_B1_c_218_n 0.00640124f $X=2.255 $Y=1.605 $X2=0 $Y2=0
cc_142 N_B2_M1010_g N_A2_M1011_g 0.0311051f $X=3.135 $Y=0.655 $X2=0 $Y2=0
cc_143 N_B2_c_135_n N_A2_M1011_g 0.00216033f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_144 N_B2_c_134_n N_A2_c_270_n 0.0260834f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_145 N_B2_c_135_n N_A2_c_270_n 0.00108681f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_146 N_B2_M1017_g N_A2_c_271_n 0.0188027f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B2_c_134_n N_A2_c_271_n 0.00191748f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_148 N_B2_c_135_n N_A2_c_271_n 0.0172639f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_149 B2 N_A_27_367#_c_396_n 0.0222158f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_150 N_B2_M1014_g N_A_27_367#_c_397_n 0.00329158f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_B2_M1014_g N_A_27_367#_c_398_n 0.0131906f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_152 B2 N_A_27_367#_c_398_n 0.0460137f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_153 N_B2_c_137_n N_A_27_367#_c_398_n 5.37952e-19 $X=1.825 $Y=1.51 $X2=0 $Y2=0
cc_154 N_B2_c_138_n N_A_27_367#_c_408_n 0.0334968f $X=2.255 $Y=1.605 $X2=0 $Y2=0
cc_155 N_B2_M1014_g N_A_27_367#_c_409_n 0.01171f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_156 B2 N_A_27_367#_c_409_n 0.0232019f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_157 N_B2_c_137_n N_A_27_367#_c_409_n 2.21398e-19 $X=1.825 $Y=1.51 $X2=0 $Y2=0
cc_158 N_B2_M1017_g N_A_27_367#_c_412_n 0.0109549f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B2_c_133_n N_A_27_367#_c_412_n 0.0166688f $X=3 $Y=1.7 $X2=0 $Y2=0
cc_160 N_B2_c_134_n N_A_27_367#_c_412_n 0.00553229f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_161 N_B2_c_135_n N_A_27_367#_c_412_n 2.45382e-19 $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_162 N_B2_M1004_g N_Y_c_446_n 0.0185192f $X=1.845 $Y=0.655 $X2=0 $Y2=0
cc_163 N_B2_M1010_g N_Y_c_446_n 0.0170169f $X=3.135 $Y=0.655 $X2=0 $Y2=0
cc_164 N_B2_c_133_n N_Y_c_446_n 0.00943636f $X=3 $Y=1.7 $X2=0 $Y2=0
cc_165 N_B2_c_134_n N_Y_c_446_n 0.0120643f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_166 N_B2_c_135_n N_Y_c_446_n 0.00363504f $X=3.165 $Y=1.46 $X2=0 $Y2=0
cc_167 B2 N_Y_c_446_n 0.048345f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_168 N_B2_c_137_n N_Y_c_446_n 0.00344256f $X=1.825 $Y=1.51 $X2=0 $Y2=0
cc_169 B2 Y 0.0293377f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_170 N_B2_M1014_g N_A_303_367#_c_503_n 0.0114565f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_B2_M1017_g N_A_303_367#_c_504_n 0.0114565f $X=3.145 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_B2_c_134_n N_A_303_367#_c_505_n 0.00512289f $X=3.165 $Y=1.46 $X2=0
+ $Y2=0
cc_173 N_B2_c_135_n N_A_303_367#_c_505_n 3.19279e-19 $X=3.165 $Y=1.46 $X2=0
+ $Y2=0
cc_174 N_B2_M1014_g N_VPWR_c_564_n 0.00357877f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_175 N_B2_M1017_g N_VPWR_c_564_n 0.00357877f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_176 N_B2_M1014_g N_VPWR_c_561_n 0.00667818f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_177 N_B2_M1017_g N_VPWR_c_561_n 0.00549753f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_178 N_B2_M1010_g N_VGND_c_631_n 0.00552762f $X=3.135 $Y=0.655 $X2=0 $Y2=0
cc_179 N_B2_M1004_g N_VGND_c_633_n 0.00564095f $X=1.845 $Y=0.655 $X2=0 $Y2=0
cc_180 N_B2_M1010_g N_VGND_c_633_n 0.00548501f $X=3.135 $Y=0.655 $X2=0 $Y2=0
cc_181 N_B2_M1004_g N_VGND_c_638_n 0.00513726f $X=1.845 $Y=0.655 $X2=0 $Y2=0
cc_182 N_B2_M1010_g N_VGND_c_638_n 0.00651887f $X=3.135 $Y=0.655 $X2=0 $Y2=0
cc_183 N_B2_M1004_g N_VGND_c_640_n 0.0104877f $X=1.845 $Y=0.655 $X2=0 $Y2=0
cc_184 N_B2_M1010_g N_A_384_47#_c_696_n 0.00402193f $X=3.135 $Y=0.655 $X2=0
+ $Y2=0
cc_185 N_B1_M1000_g N_A_27_367#_c_408_n 0.01115f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B1_M1006_g N_A_27_367#_c_408_n 0.01115f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_187 N_B1_M1000_g N_A_27_367#_c_409_n 0.0108074f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_188 N_B1_M1006_g N_A_27_367#_c_409_n 5.5933e-19 $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_189 N_B1_M1000_g N_A_27_367#_c_412_n 5.5933e-19 $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_190 N_B1_M1006_g N_A_27_367#_c_412_n 0.0108074f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B1_c_213_n N_Y_c_446_n 0.012325f $X=2.275 $Y=1.185 $X2=0 $Y2=0
cc_192 N_B1_c_215_n N_Y_c_446_n 0.0106382f $X=2.705 $Y=1.185 $X2=0 $Y2=0
cc_193 B1 N_Y_c_446_n 0.0251351f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_194 N_B1_c_218_n N_Y_c_446_n 0.00237053f $X=2.705 $Y=1.35 $X2=0 $Y2=0
cc_195 N_B1_M1000_g N_A_303_367#_c_503_n 0.0114565f $X=2.285 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_B1_M1006_g N_A_303_367#_c_504_n 0.0114565f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_B1_M1000_g N_VPWR_c_564_n 0.00357877f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_198 N_B1_M1006_g N_VPWR_c_564_n 0.00357877f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_199 N_B1_M1000_g N_VPWR_c_561_n 0.00537849f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_200 N_B1_M1006_g N_VPWR_c_561_n 0.00537849f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_201 N_B1_c_213_n N_VGND_c_633_n 0.00364081f $X=2.275 $Y=1.185 $X2=0 $Y2=0
cc_202 N_B1_c_215_n N_VGND_c_633_n 0.00364081f $X=2.705 $Y=1.185 $X2=0 $Y2=0
cc_203 N_B1_c_213_n N_VGND_c_638_n 0.0054574f $X=2.275 $Y=1.185 $X2=0 $Y2=0
cc_204 N_B1_c_215_n N_VGND_c_638_n 0.0054574f $X=2.705 $Y=1.185 $X2=0 $Y2=0
cc_205 N_B1_c_213_n N_VGND_c_640_n 0.00122952f $X=2.275 $Y=1.185 $X2=0 $Y2=0
cc_206 N_B1_c_213_n N_A_384_47#_c_696_n 0.0121033f $X=2.275 $Y=1.185 $X2=0 $Y2=0
cc_207 N_B1_c_215_n N_A_384_47#_c_696_n 0.0120124f $X=2.705 $Y=1.185 $X2=0 $Y2=0
cc_208 N_A2_M1011_g N_A1_c_342_n 0.0421704f $X=3.725 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_209 N_A2_M1012_g N_A1_M1009_g 0.0245418f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A2_c_269_n N_A1_M1009_g 0.0103825f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_211 N_A2_M1015_g N_A1_c_344_n 0.0269756f $X=5.015 $Y=0.655 $X2=0 $Y2=0
cc_212 N_A2_M1016_g N_A1_M1019_g 0.0269756f $X=5.015 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A2_c_269_n N_A1_M1019_g 0.010446f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_214 N_A2_M1011_g A1 0.00373094f $X=3.725 $Y=0.655 $X2=0 $Y2=0
cc_215 N_A2_c_268_n A1 0.0142774f $X=5.015 $Y=1.375 $X2=0 $Y2=0
cc_216 N_A2_c_269_n A1 0.08813f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_217 N_A2_c_270_n A1 0.0081926f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_218 N_A2_c_271_n A1 7.14113e-19 $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_219 A2 A1 0.0186394f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A2_c_273_n A1 0.00741149f $X=5.49 $Y=1.375 $X2=0 $Y2=0
cc_221 N_A2_c_268_n N_A1_c_347_n 0.0269756f $X=5.015 $Y=1.375 $X2=0 $Y2=0
cc_222 N_A2_c_269_n N_A1_c_347_n 0.00243542f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_223 N_A2_c_270_n N_A1_c_347_n 0.00108928f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_224 N_A2_c_271_n N_A1_c_347_n 0.0215588f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_225 A2 N_A1_c_347_n 4.19049e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_226 N_A2_M1011_g N_Y_c_469_n 5.8325e-19 $X=3.725 $Y=0.655 $X2=0 $Y2=0
cc_227 N_A2_M1011_g N_Y_c_446_n 0.0170458f $X=3.725 $Y=0.655 $X2=0 $Y2=0
cc_228 N_A2_c_269_n N_Y_c_446_n 0.00418135f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_229 N_A2_c_270_n N_Y_c_446_n 0.0105714f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_230 N_A2_c_271_n N_Y_c_446_n 0.00181918f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_231 N_A2_M1012_g N_A_303_367#_c_505_n 2.7414e-19 $X=3.615 $Y=2.465 $X2=0
+ $Y2=0
cc_232 N_A2_c_270_n N_A_303_367#_c_505_n 7.37441e-19 $X=3.705 $Y=1.51 $X2=0
+ $Y2=0
cc_233 N_A2_M1012_g N_A_303_367#_c_511_n 0.0109654f $X=3.615 $Y=2.465 $X2=0
+ $Y2=0
cc_234 N_A2_M1012_g N_A_303_367#_c_512_n 0.0127704f $X=3.615 $Y=2.465 $X2=0
+ $Y2=0
cc_235 N_A2_c_269_n N_A_303_367#_c_512_n 0.0288357f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_236 N_A2_c_270_n N_A_303_367#_c_512_n 0.0161105f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_237 N_A2_c_271_n N_A_303_367#_c_512_n 8.4523e-19 $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_238 N_A2_M1012_g N_A_303_367#_c_516_n 4.69865e-19 $X=3.615 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A2_M1016_g N_A_303_367#_c_517_n 0.0122129f $X=5.015 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_A2_c_269_n N_A_303_367#_c_517_n 0.0409786f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_241 N_A2_c_269_n N_A_303_367#_c_501_n 0.0155834f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_242 N_A2_c_273_n N_A_303_367#_c_501_n 6.4892e-19 $X=5.49 $Y=1.375 $X2=0 $Y2=0
cc_243 N_A2_c_274_n N_A_303_367#_c_501_n 0.00551758f $X=5.505 $Y=1.615 $X2=0
+ $Y2=0
cc_244 N_A2_c_269_n N_A_303_367#_c_522_n 0.0166768f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_245 N_A2_M1012_g N_VPWR_c_562_n 0.00416163f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A2_M1016_g N_VPWR_c_563_n 0.0161163f $X=5.015 $Y=2.465 $X2=0 $Y2=0
cc_247 N_A2_M1012_g N_VPWR_c_564_n 0.00570203f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A2_M1016_g N_VPWR_c_568_n 0.00486043f $X=5.015 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A2_M1012_g N_VPWR_c_561_n 0.0106301f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A2_M1016_g N_VPWR_c_561_n 0.00935452f $X=5.015 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A2_M1011_g N_VGND_c_631_n 0.00953649f $X=3.725 $Y=0.655 $X2=0 $Y2=0
cc_252 N_A2_M1015_g N_VGND_c_632_n 0.00662502f $X=5.015 $Y=0.655 $X2=0 $Y2=0
cc_253 N_A2_c_269_n N_VGND_c_632_n 0.00574448f $X=5.335 $Y=1.7 $X2=0 $Y2=0
cc_254 A2 N_VGND_c_632_n 0.00507585f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_255 N_A2_c_273_n N_VGND_c_632_n 0.0060872f $X=5.49 $Y=1.375 $X2=0 $Y2=0
cc_256 N_A2_M1011_g N_VGND_c_635_n 0.00547467f $X=3.725 $Y=0.655 $X2=0 $Y2=0
cc_257 N_A2_M1015_g N_VGND_c_635_n 0.00547432f $X=5.015 $Y=0.655 $X2=0 $Y2=0
cc_258 N_A2_M1011_g N_VGND_c_638_n 0.00647216f $X=3.725 $Y=0.655 $X2=0 $Y2=0
cc_259 N_A2_M1015_g N_VGND_c_638_n 0.0108612f $X=5.015 $Y=0.655 $X2=0 $Y2=0
cc_260 N_A2_M1011_g N_A_760_47#_c_707_n 0.00310894f $X=3.725 $Y=0.655 $X2=0
+ $Y2=0
cc_261 N_A2_M1015_g N_A_760_47#_c_708_n 0.0107823f $X=5.015 $Y=0.655 $X2=0 $Y2=0
cc_262 N_A1_c_342_n N_Y_c_469_n 0.00353788f $X=4.155 $Y=1.185 $X2=0 $Y2=0
cc_263 N_A1_c_347_n N_Y_c_469_n 0.00235487f $X=4.585 $Y=1.35 $X2=0 $Y2=0
cc_264 N_A1_c_342_n N_Y_c_446_n 0.00996418f $X=4.155 $Y=1.185 $X2=0 $Y2=0
cc_265 A1 N_Y_c_446_n 0.0331051f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_266 N_A1_M1009_g N_A_303_367#_c_511_n 4.33124e-19 $X=4.155 $Y=2.465 $X2=0
+ $Y2=0
cc_267 N_A1_M1009_g N_A_303_367#_c_512_n 0.0127761f $X=4.155 $Y=2.465 $X2=0
+ $Y2=0
cc_268 N_A1_M1009_g N_A_303_367#_c_516_n 0.0113428f $X=4.155 $Y=2.465 $X2=0
+ $Y2=0
cc_269 N_A1_M1019_g N_A_303_367#_c_517_n 0.0122129f $X=4.585 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_A1_M1009_g N_A_303_367#_c_522_n 2.74535e-19 $X=4.155 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A1_M1009_g N_VPWR_c_562_n 0.00266796f $X=4.155 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A1_M1009_g N_VPWR_c_563_n 7.23054e-19 $X=4.155 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A1_M1019_g N_VPWR_c_563_n 0.0143485f $X=4.585 $Y=2.465 $X2=0 $Y2=0
cc_274 N_A1_M1009_g N_VPWR_c_566_n 0.00571722f $X=4.155 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A1_M1019_g N_VPWR_c_566_n 0.00486043f $X=4.585 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A1_M1009_g N_VPWR_c_561_n 0.0105481f $X=4.155 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A1_M1019_g N_VPWR_c_561_n 0.00824727f $X=4.585 $Y=2.465 $X2=0 $Y2=0
cc_278 A1 N_VGND_c_632_n 0.00184572f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_279 N_A1_c_342_n N_VGND_c_635_n 0.00357877f $X=4.155 $Y=1.185 $X2=0 $Y2=0
cc_280 N_A1_c_344_n N_VGND_c_635_n 0.00357842f $X=4.585 $Y=1.185 $X2=0 $Y2=0
cc_281 N_A1_c_342_n N_VGND_c_638_n 0.00537654f $X=4.155 $Y=1.185 $X2=0 $Y2=0
cc_282 N_A1_c_344_n N_VGND_c_638_n 0.00537652f $X=4.585 $Y=1.185 $X2=0 $Y2=0
cc_283 N_A1_c_342_n N_A_760_47#_c_707_n 0.00990217f $X=4.155 $Y=1.185 $X2=0
+ $Y2=0
cc_284 N_A1_c_344_n N_A_760_47#_c_707_n 0.0121331f $X=4.585 $Y=1.185 $X2=0 $Y2=0
cc_285 N_A1_c_342_n N_A_760_47#_c_708_n 9.24211e-19 $X=4.155 $Y=1.185 $X2=0
+ $Y2=0
cc_286 N_A1_c_344_n N_A_760_47#_c_708_n 0.0099917f $X=4.585 $Y=1.185 $X2=0 $Y2=0
cc_287 A1 N_A_760_47#_c_708_n 0.0222258f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_288 N_A_27_367#_c_401_n N_Y_M1005_s 0.00332344f $X=1.025 $Y=2.99 $X2=0 $Y2=0
cc_289 N_A_27_367#_c_401_n Y 0.0159805f $X=1.025 $Y=2.99 $X2=0 $Y2=0
cc_290 N_A_27_367#_c_398_n N_A_303_367#_M1014_d 0.00509633f $X=1.905 $Y=2.04
+ $X2=-0.19 $Y2=1.655
cc_291 N_A_27_367#_c_408_n N_A_303_367#_M1000_s 0.00339614f $X=2.765 $Y=2.04
+ $X2=0 $Y2=0
cc_292 N_A_27_367#_c_397_n N_A_303_367#_c_499_n 0.0452321f $X=1.155 $Y=2.905
+ $X2=0 $Y2=0
cc_293 N_A_27_367#_c_398_n N_A_303_367#_c_499_n 0.0202165f $X=1.905 $Y=2.04
+ $X2=0 $Y2=0
cc_294 N_A_27_367#_M1014_s N_A_303_367#_c_503_n 0.00332344f $X=1.93 $Y=1.835
+ $X2=0 $Y2=0
cc_295 N_A_27_367#_c_409_n N_A_303_367#_c_503_n 0.0159805f $X=2.07 $Y=2.04 $X2=0
+ $Y2=0
cc_296 N_A_27_367#_c_397_n N_A_303_367#_c_500_n 0.0147157f $X=1.155 $Y=2.905
+ $X2=0 $Y2=0
cc_297 N_A_27_367#_c_408_n N_A_303_367#_c_535_n 0.0135055f $X=2.765 $Y=2.04
+ $X2=0 $Y2=0
cc_298 N_A_27_367#_M1006_d N_A_303_367#_c_504_n 0.00332344f $X=2.79 $Y=1.835
+ $X2=0 $Y2=0
cc_299 N_A_27_367#_c_412_n N_A_303_367#_c_504_n 0.0159805f $X=2.93 $Y=2.04 $X2=0
+ $Y2=0
cc_300 N_A_27_367#_c_394_n N_VPWR_c_564_n 0.0179183f $X=0.225 $Y=2.905 $X2=0
+ $Y2=0
cc_301 N_A_27_367#_c_401_n N_VPWR_c_564_n 0.0361172f $X=1.025 $Y=2.99 $X2=0
+ $Y2=0
cc_302 N_A_27_367#_c_397_n N_VPWR_c_564_n 0.0179183f $X=1.155 $Y=2.905 $X2=0
+ $Y2=0
cc_303 N_A_27_367#_M1005_d N_VPWR_c_561_n 0.00215161f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_304 N_A_27_367#_M1018_d N_VPWR_c_561_n 0.00215161f $X=0.98 $Y=1.835 $X2=0
+ $Y2=0
cc_305 N_A_27_367#_M1014_s N_VPWR_c_561_n 0.00225186f $X=1.93 $Y=1.835 $X2=0
+ $Y2=0
cc_306 N_A_27_367#_M1006_d N_VPWR_c_561_n 0.00225186f $X=2.79 $Y=1.835 $X2=0
+ $Y2=0
cc_307 N_A_27_367#_c_394_n N_VPWR_c_561_n 0.0101082f $X=0.225 $Y=2.905 $X2=0
+ $Y2=0
cc_308 N_A_27_367#_c_401_n N_VPWR_c_561_n 0.023676f $X=1.025 $Y=2.99 $X2=0 $Y2=0
cc_309 N_A_27_367#_c_397_n N_VPWR_c_561_n 0.0101082f $X=1.155 $Y=2.905 $X2=0
+ $Y2=0
cc_310 N_Y_M1005_s N_VPWR_c_561_n 0.00225186f $X=0.55 $Y=1.835 $X2=0 $Y2=0
cc_311 N_Y_c_446_n N_VGND_M1007_s 0.019321f $X=4.205 $Y=0.852 $X2=0 $Y2=0
cc_312 N_Y_c_446_n N_VGND_M1010_s 0.0142416f $X=4.205 $Y=0.852 $X2=0 $Y2=0
cc_313 N_Y_c_446_n N_VGND_c_631_n 0.0262444f $X=4.205 $Y=0.852 $X2=0 $Y2=0
cc_314 N_Y_M1003_d N_VGND_c_638_n 0.00250503f $X=0.66 $Y=0.235 $X2=0 $Y2=0
cc_315 N_Y_M1002_s N_VGND_c_638_n 0.00226546f $X=2.35 $Y=0.235 $X2=0 $Y2=0
cc_316 N_Y_M1001_d N_VGND_c_638_n 0.00225186f $X=4.23 $Y=0.235 $X2=0 $Y2=0
cc_317 N_Y_c_446_n N_VGND_c_638_n 0.0294749f $X=4.205 $Y=0.852 $X2=0 $Y2=0
cc_318 Y N_VGND_c_638_n 0.00992063f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_319 Y N_VGND_c_639_n 0.0157207f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_320 N_Y_c_446_n N_VGND_c_640_n 0.0480912f $X=4.205 $Y=0.852 $X2=0 $Y2=0
cc_321 N_Y_c_446_n N_A_384_47#_M1004_d 0.00436079f $X=4.205 $Y=0.852 $X2=-0.19
+ $Y2=-0.245
cc_322 N_Y_c_446_n N_A_384_47#_M1013_d 0.00497616f $X=4.205 $Y=0.852 $X2=0 $Y2=0
cc_323 N_Y_M1002_s N_A_384_47#_c_696_n 0.0034017f $X=2.35 $Y=0.235 $X2=0 $Y2=0
cc_324 N_Y_c_446_n N_A_384_47#_c_696_n 0.0610357f $X=4.205 $Y=0.852 $X2=0 $Y2=0
cc_325 N_Y_c_446_n N_A_760_47#_M1011_d 0.00491639f $X=4.205 $Y=0.852 $X2=-0.19
+ $Y2=-0.245
cc_326 N_Y_M1001_d N_A_760_47#_c_707_n 0.00340217f $X=4.23 $Y=0.235 $X2=0 $Y2=0
cc_327 N_Y_c_469_n N_A_760_47#_c_707_n 0.0134855f $X=4.37 $Y=0.83 $X2=0 $Y2=0
cc_328 N_Y_c_446_n N_A_760_47#_c_707_n 0.0135687f $X=4.205 $Y=0.852 $X2=0 $Y2=0
cc_329 N_A_303_367#_c_512_n N_VPWR_M1012_d 0.00590698f $X=4.22 $Y=2.04 $X2=-0.19
+ $Y2=1.655
cc_330 N_A_303_367#_c_517_n N_VPWR_M1019_d 0.00353353f $X=5.145 $Y=2.04 $X2=0
+ $Y2=0
cc_331 N_A_303_367#_c_512_n N_VPWR_c_562_n 0.022455f $X=4.22 $Y=2.04 $X2=0 $Y2=0
cc_332 N_A_303_367#_c_517_n N_VPWR_c_563_n 0.0170777f $X=5.145 $Y=2.04 $X2=0
+ $Y2=0
cc_333 N_A_303_367#_c_503_n N_VPWR_c_564_n 0.0361172f $X=2.405 $Y=2.99 $X2=0
+ $Y2=0
cc_334 N_A_303_367#_c_500_n N_VPWR_c_564_n 0.0179183f $X=1.735 $Y=2.99 $X2=0
+ $Y2=0
cc_335 N_A_303_367#_c_504_n N_VPWR_c_564_n 0.0361172f $X=3.265 $Y=2.99 $X2=0
+ $Y2=0
cc_336 N_A_303_367#_c_511_n N_VPWR_c_564_n 0.0175816f $X=3.407 $Y=2.905 $X2=0
+ $Y2=0
cc_337 N_A_303_367#_c_546_p N_VPWR_c_564_n 0.0125234f $X=2.5 $Y=2.99 $X2=0 $Y2=0
cc_338 N_A_303_367#_c_516_n N_VPWR_c_566_n 0.0143106f $X=4.37 $Y=2.48 $X2=0
+ $Y2=0
cc_339 N_A_303_367#_c_502_n N_VPWR_c_568_n 0.0174563f $X=5.23 $Y=2.48 $X2=0
+ $Y2=0
cc_340 N_A_303_367#_M1014_d N_VPWR_c_561_n 0.00215161f $X=1.515 $Y=1.835 $X2=0
+ $Y2=0
cc_341 N_A_303_367#_M1000_s N_VPWR_c_561_n 0.00223565f $X=2.36 $Y=1.835 $X2=0
+ $Y2=0
cc_342 N_A_303_367#_M1017_d N_VPWR_c_561_n 0.00255729f $X=3.22 $Y=1.835 $X2=0
+ $Y2=0
cc_343 N_A_303_367#_M1009_s N_VPWR_c_561_n 0.0041489f $X=4.23 $Y=1.835 $X2=0
+ $Y2=0
cc_344 N_A_303_367#_M1016_s N_VPWR_c_561_n 0.0040649f $X=5.09 $Y=1.835 $X2=0
+ $Y2=0
cc_345 N_A_303_367#_c_503_n N_VPWR_c_561_n 0.023676f $X=2.405 $Y=2.99 $X2=0
+ $Y2=0
cc_346 N_A_303_367#_c_500_n N_VPWR_c_561_n 0.0101082f $X=1.735 $Y=2.99 $X2=0
+ $Y2=0
cc_347 N_A_303_367#_c_504_n N_VPWR_c_561_n 0.023676f $X=3.265 $Y=2.99 $X2=0
+ $Y2=0
cc_348 N_A_303_367#_c_511_n N_VPWR_c_561_n 0.0109612f $X=3.407 $Y=2.905 $X2=0
+ $Y2=0
cc_349 N_A_303_367#_c_516_n N_VPWR_c_561_n 0.00893886f $X=4.37 $Y=2.48 $X2=0
+ $Y2=0
cc_350 N_A_303_367#_c_502_n N_VPWR_c_561_n 0.00963639f $X=5.23 $Y=2.48 $X2=0
+ $Y2=0
cc_351 N_A_303_367#_c_546_p N_VPWR_c_561_n 0.00738676f $X=2.5 $Y=2.99 $X2=0
+ $Y2=0
cc_352 N_VGND_c_638_n N_A_384_47#_M1004_d 0.00246704f $X=5.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_353 N_VGND_c_638_n N_A_384_47#_M1013_d 0.00226546f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_c_633_n N_A_384_47#_c_696_n 0.0543512f $X=3.26 $Y=0 $X2=0 $Y2=0
cc_355 N_VGND_c_638_n N_A_384_47#_c_696_n 0.0408631f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_638_n N_A_760_47#_M1011_d 0.00223577f $X=5.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_357 N_VGND_c_638_n N_A_760_47#_M1008_s 0.00223559f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_631_n N_A_760_47#_c_707_n 0.0175924f $X=3.425 $Y=0.48 $X2=0
+ $Y2=0
cc_359 N_VGND_c_635_n N_A_760_47#_c_707_n 0.0482626f $X=5.135 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_638_n N_A_760_47#_c_707_n 0.0310329f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_635_n N_A_760_47#_c_708_n 0.01906f $X=5.135 $Y=0 $X2=0 $Y2=0
cc_362 N_VGND_c_638_n N_A_760_47#_c_708_n 0.0124545f $X=5.52 $Y=0 $X2=0 $Y2=0
