* File: sky130_fd_sc_lp__sdfxbp_1.spice
* Created: Wed Sep  2 10:36:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfxbp_1.pex.spice"
.subckt sky130_fd_sc_lp__sdfxbp_1  VNB VPB SCD D SCE CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1012 A_124_119# N_SCD_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1031 N_A_196_119#_M1031_d N_SCE_M1031_g A_124_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=15.708 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1014 A_304_119# N_D_M1014_g N_A_196_119#_M1031_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=15.708 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_324_431#_M1001_g A_304_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_324_431#_M1003_d N_SCE_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_722_23#_M1005_g N_A_767_121#_M1005_s VNB NSHORT L=0.15
+ W=0.64 AD=0.273268 AS=0.1824 PD=1.67245 PS=1.85 NRD=61.872 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1021 A_1033_121# N_A_767_121#_M1021_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.179332 PD=0.63 PS=1.09755 NRD=14.28 NRS=39.276 M=1 R=2.8
+ SA=75001.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1018 N_A_722_23#_M1018_d N_A_1075_95#_M1018_g A_1033_121# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_A_196_119#_M1019_d N_A_1161_95#_M1019_g N_A_722_23#_M1018_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_1161_95#_M1013_g N_A_1075_95#_M1013_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_A_1161_95#_M1033_d N_CLK_M1033_g N_VGND_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_A_1873_497#_M1029_d N_A_1075_95#_M1029_g N_A_767_121#_M1029_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1015 A_2040_125# N_A_1161_95#_M1015_g N_A_1873_497#_M1029_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_2082_99#_M1011_g A_2040_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0988981 AS=0.0441 PD=0.859811 PS=0.63 NRD=42.132 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_2082_99#_M1007_d N_A_1873_497#_M1007_g N_VGND_M1011_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.150702 PD=1.85 PS=1.31019 NRD=0 NRS=3.744 M=1
+ R=4.26667 SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1030 N_A_2409_367#_M1030_d N_A_2082_99#_M1030_g N_VGND_M1030_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_2082_99#_M1025_g N_Q_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1239 AS=0.2226 PD=1.135 PS=2.21 NRD=2.136 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1009 N_Q_N_M1009_d N_A_2409_367#_M1009_g N_VGND_M1025_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2814 AS=0.1239 PD=2.35 PS=1.135 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1017 N_VPWR_M1017_d N_SCD_M1017_g N_A_27_483#_M1017_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1032 A_196_483# N_SCE_M1032_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1000 N_A_196_119#_M1000_d N_D_M1000_g A_196_483# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_27_483#_M1020_d N_A_324_431#_M1020_g N_A_196_119#_M1000_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_SCE_M1008_g N_A_324_431#_M1008_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1792 AS=0.3328 PD=1.84 PS=2.32 NRD=4.6098 NRS=78.4848 M=1
+ R=4.26667 SA=75000.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1004_d N_A_722_23#_M1004_g N_A_767_121#_M1004_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1792 AS=0.3399 PD=1.62 PS=2.7 NRD=0 NRS=23.443 M=1 R=5.6
+ SA=75000.3 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1023 N_A_974_425#_M1023_d N_A_767_121#_M1023_g N_VPWR_M1004_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.2562 AS=0.0896 PD=2.4 PS=0.81 NRD=260.316 NRS=74.2493 M=1
+ R=2.8 SA=75000.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1010 N_A_722_23#_M1010_d N_A_1075_95#_M1010_g N_A_196_119#_M1010_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1533 PD=0.7 PS=1.57 NRD=0 NRS=37.5088 M=1 R=2.8
+ SA=75000.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1027 N_A_974_425#_M1027_d N_A_1161_95#_M1027_g N_A_722_23#_M1010_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1449 AS=0.0588 PD=1.53 PS=0.7 NRD=37.5088 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1028 N_VPWR_M1028_d N_A_1161_95#_M1028_g N_A_1075_95#_M1028_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.18045 AS=0.1824 PD=1.405 PS=1.85 NRD=69.8562 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1016 N_A_1161_95#_M1016_d N_CLK_M1016_g N_VPWR_M1028_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.18045 PD=1.85 PS=1.405 NRD=0 NRS=69.8562 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_1873_497#_M1002_d N_A_1075_95#_M1002_g N_A_1786_497#_M1002_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.111683 AS=0.1197 PD=0.986667 PS=1.41 NRD=98.9137
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1035 N_A_767_121#_M1035_d N_A_1161_95#_M1035_g N_A_1873_497#_M1002_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2226 AS=0.223367 PD=2.21 PS=1.97333 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_A_2082_99#_M1006_g N_A_1786_497#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=46.886 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1022 N_A_2082_99#_M1022_d N_A_1873_497#_M1022_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2394 AS=0.1792 PD=2.25 PS=1.62 NRD=4.6886 NRS=0 M=1 R=5.6
+ SA=75000.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1034 N_VPWR_M1034_d N_A_2082_99#_M1034_g N_A_2409_367#_M1034_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.136185 AS=0.1696 PD=1.10147 PS=1.81 NRD=48.5605 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1024 N_Q_M1024_d N_A_2082_99#_M1024_g N_VPWR_M1034_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.268115 PD=3.05 PS=2.16853 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1026 N_Q_N_M1026_d N_A_2409_367#_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX36_noxref VNB VPB NWDIODE A=27.5647 P=33.29
c_147 VNB 0 1.73242e-19 $X=0 $Y=0
c_271 VPB 0 1.8781e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfxbp_1.pxi.spice"
*
.ends
*
*
