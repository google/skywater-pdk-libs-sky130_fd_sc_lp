* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__bufinv_16 A VGND VNB VPB VPWR Y
X0 Y a_413_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_413_49# a_63_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_413_49# a_63_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND a_413_49# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 Y a_413_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR a_63_49# a_413_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND a_413_49# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_63_49# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Y a_413_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VGND a_413_49# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 Y a_413_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 Y a_413_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 Y a_413_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 Y a_413_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VPWR a_413_49# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND a_63_49# a_413_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 Y a_413_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VPWR a_63_49# a_413_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_413_49# a_63_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 Y a_413_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VGND a_413_49# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 VGND a_413_49# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_63_49# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 Y a_413_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VPWR a_413_49# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VGND a_413_49# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 Y a_413_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 Y a_413_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 VPWR a_413_49# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_63_49# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 VGND a_413_49# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 VPWR a_63_49# a_413_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 Y a_413_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 VPWR a_413_49# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 a_413_49# a_63_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 VPWR A a_63_49# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 VGND a_63_49# a_413_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X37 VPWR a_413_49# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 VPWR a_413_49# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 Y a_413_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X40 a_63_49# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X41 VGND a_413_49# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X42 VGND A a_63_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X43 a_413_49# a_63_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X44 a_413_49# a_63_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X45 VPWR a_413_49# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X46 VPWR a_413_49# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X47 Y a_413_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X48 VGND a_63_49# a_413_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X49 Y a_413_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
