# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o21ba_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o21ba_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.210000 3.755000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.210000 3.215000 2.605000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.210000 0.895000 1.750000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.255000 1.315000 1.850000 ;
        RECT 1.065000 1.850000 1.670000 2.120000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.085000  0.700000 0.360000 1.030000 ;
      RECT 0.085000  1.030000 0.270000 1.920000 ;
      RECT 0.085000  1.920000 0.595000 2.290000 ;
      RECT 0.085000  2.290000 2.235000 2.460000 ;
      RECT 0.530000  0.085000 0.895000 1.040000 ;
      RECT 0.910000  2.630000 1.240000 3.245000 ;
      RECT 1.485000  0.085000 1.815000 0.835000 ;
      RECT 1.485000  1.005000 2.615000 1.175000 ;
      RECT 1.485000  1.175000 1.795000 1.515000 ;
      RECT 1.840000  2.630000 2.170000 3.245000 ;
      RECT 2.005000  0.255000 2.265000 1.005000 ;
      RECT 2.005000  1.345000 2.265000 1.675000 ;
      RECT 2.005000  1.675000 2.235000 2.290000 ;
      RECT 2.405000  1.855000 2.615000 3.075000 ;
      RECT 2.435000  0.255000 2.765000 0.655000 ;
      RECT 2.435000  0.655000 3.705000 0.835000 ;
      RECT 2.435000  1.175000 2.615000 1.855000 ;
      RECT 2.935000  0.085000 3.265000 0.485000 ;
      RECT 3.375000  0.835000 3.705000 1.040000 ;
      RECT 3.385000  1.920000 3.700000 3.245000 ;
      RECT 3.435000  0.255000 3.705000 0.655000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__o21ba_2
END LIBRARY
