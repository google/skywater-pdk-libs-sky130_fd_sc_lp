* File: sky130_fd_sc_lp__or3_0.pxi.spice
* Created: Fri Aug 28 11:22:58 2020
* 
x_PM_SKY130_FD_SC_LP__OR3_0%C N_C_M1001_g N_C_M1000_g N_C_c_64_n N_C_c_69_n C C
+ C N_C_c_66_n PM_SKY130_FD_SC_LP__OR3_0%C
x_PM_SKY130_FD_SC_LP__OR3_0%B N_B_M1002_g N_B_M1007_g N_B_c_101_n N_B_c_102_n B
+ B B N_B_c_106_n N_B_c_107_n PM_SKY130_FD_SC_LP__OR3_0%B
x_PM_SKY130_FD_SC_LP__OR3_0%A N_A_M1003_g N_A_M1004_g N_A_c_159_n N_A_c_164_n A
+ A N_A_c_161_n PM_SKY130_FD_SC_LP__OR3_0%A
x_PM_SKY130_FD_SC_LP__OR3_0%A_29_55# N_A_29_55#_M1001_s N_A_29_55#_M1007_d
+ N_A_29_55#_M1000_s N_A_29_55#_M1006_g N_A_29_55#_M1005_g N_A_29_55#_c_218_n
+ N_A_29_55#_c_219_n N_A_29_55#_c_210_n N_A_29_55#_c_221_n N_A_29_55#_c_222_n
+ N_A_29_55#_c_211_n N_A_29_55#_c_212_n N_A_29_55#_c_213_n N_A_29_55#_c_223_n
+ N_A_29_55#_c_224_n N_A_29_55#_c_214_n N_A_29_55#_c_215_n N_A_29_55#_c_216_n
+ PM_SKY130_FD_SC_LP__OR3_0%A_29_55#
x_PM_SKY130_FD_SC_LP__OR3_0%VPWR N_VPWR_M1003_d N_VPWR_c_296_n VPWR
+ N_VPWR_c_297_n N_VPWR_c_298_n N_VPWR_c_295_n N_VPWR_c_300_n
+ PM_SKY130_FD_SC_LP__OR3_0%VPWR
x_PM_SKY130_FD_SC_LP__OR3_0%X N_X_M1006_d N_X_M1005_d X X X X X X X N_X_c_320_n
+ X PM_SKY130_FD_SC_LP__OR3_0%X
x_PM_SKY130_FD_SC_LP__OR3_0%VGND N_VGND_M1001_d N_VGND_M1004_d N_VGND_c_339_n
+ N_VGND_c_340_n N_VGND_c_341_n VGND N_VGND_c_342_n N_VGND_c_343_n
+ N_VGND_c_344_n N_VGND_c_345_n PM_SKY130_FD_SC_LP__OR3_0%VGND
cc_1 VNB N_C_M1001_g 0.040293f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.485
cc_2 VNB N_C_c_64_n 0.029551f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.715
cc_3 VNB C 0.00830305f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_4 VNB N_C_c_66_n 0.0218585f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.245
cc_5 VNB N_B_M1002_g 0.0080888f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.485
cc_6 VNB N_B_c_101_n 0.0220598f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=2.615
cc_7 VNB N_B_c_102_n 0.028385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB B 0.00233035f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.715
cc_9 VNB B 0.00141102f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.865
cc_10 VNB B 0.00337172f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_11 VNB N_B_c_106_n 0.0258332f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.245
cc_12 VNB N_B_c_107_n 0.0156839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_M1004_g 0.0368252f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.865
cc_14 VNB N_A_c_159_n 0.0191366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A 0.00490559f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_16 VNB N_A_c_161_n 0.0157989f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.245
cc_17 VNB N_A_29_55#_M1006_g 0.058694f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.865
cc_18 VNB N_A_29_55#_c_210_n 0.0651924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_29_55#_c_211_n 0.00265598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_29_55#_c_212_n 0.00656187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_29_55#_c_213_n 0.00521361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_29_55#_c_214_n 0.00285856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_29_55#_c_215_n 0.0148318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_29_55#_c_216_n 0.00386064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_295_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB X 0.0534323f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=2.615
cc_27 VNB N_X_c_320_n 0.0166693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_339_n 0.00574374f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=2.615
cc_29 VNB N_VGND_c_340_n 0.0168921f $X=-0.19 $Y=-0.245 $X2=0.682 $Y2=1.865
cc_30 VNB N_VGND_c_341_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_31 VNB N_VGND_c_342_n 0.0212057f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.245
cc_32 VNB N_VGND_c_343_n 0.177823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_344_n 0.0167135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_345_n 0.0198298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_C_M1000_g 0.0458873f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=2.615
cc_36 VPB N_C_c_64_n 0.00481325f $X=-0.19 $Y=1.655 $X2=0.682 $Y2=1.715
cc_37 VPB N_C_c_69_n 0.0318659f $X=-0.19 $Y=1.655 $X2=0.682 $Y2=1.865
cc_38 VPB C 3.89831e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_39 VPB N_B_M1002_g 0.0426774f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.485
cc_40 VPB B 0.00413483f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_41 VPB N_A_M1003_g 0.0406247f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.485
cc_42 VPB N_A_c_159_n 0.00186984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_c_164_n 0.0217764f $X=-0.19 $Y=1.655 $X2=0.682 $Y2=1.715
cc_44 VPB A 0.00167835f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_45 VPB N_A_29_55#_M1005_g 0.0283544f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_29_55#_c_218_n 0.0247349f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.245
cc_47 VPB N_A_29_55#_c_219_n 0.0178608f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.245
cc_48 VPB N_A_29_55#_c_210_n 0.0218623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_29_55#_c_221_n 0.0183811f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.665
cc_50 VPB N_A_29_55#_c_222_n 0.0369517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_29_55#_c_223_n 0.00288783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_29_55#_c_224_n 0.0383595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_29_55#_c_214_n 4.22059e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_29_55#_c_215_n 0.00376664f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_296_n 0.0192788f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.715
cc_56 VPB N_VPWR_c_297_n 0.0533858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_298_n 0.01875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_295_n 0.0927178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_300_n 0.0112264f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.245
cc_60 VPB X 0.0371697f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=2.615
cc_61 VPB X 0.0227952f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_62 VPB X 0.0115022f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 N_C_c_64_n N_B_M1002_g 0.00774443f $X=0.682 $Y=1.715 $X2=0 $Y2=0
cc_64 N_C_c_69_n N_B_M1002_g 0.0785239f $X=0.682 $Y=1.865 $X2=0 $Y2=0
cc_65 C N_B_M1002_g 7.78255e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_66 N_C_M1001_g N_B_c_102_n 0.00583103f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_67 C N_B_c_102_n 0.00481809f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_68 N_C_M1001_g B 2.25363e-19 $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_69 C B 0.0833769f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_70 N_C_c_66_n B 2.10094e-19 $X=0.64 $Y=1.245 $X2=0 $Y2=0
cc_71 N_C_c_64_n B 2.10094e-19 $X=0.682 $Y=1.715 $X2=0 $Y2=0
cc_72 N_C_c_64_n B 7.67461e-19 $X=0.682 $Y=1.715 $X2=0 $Y2=0
cc_73 N_C_c_69_n B 0.00111118f $X=0.682 $Y=1.865 $X2=0 $Y2=0
cc_74 N_C_c_66_n N_B_c_106_n 0.0122915f $X=0.64 $Y=1.245 $X2=0 $Y2=0
cc_75 N_C_c_64_n N_B_c_107_n 0.0122915f $X=0.682 $Y=1.715 $X2=0 $Y2=0
cc_76 N_C_M1001_g N_A_29_55#_c_210_n 0.0335588f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_77 N_C_M1000_g N_A_29_55#_c_210_n 0.00473163f $X=0.88 $Y=2.615 $X2=0 $Y2=0
cc_78 C N_A_29_55#_c_210_n 0.081912f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_79 N_C_M1000_g N_A_29_55#_c_221_n 0.00967579f $X=0.88 $Y=2.615 $X2=0 $Y2=0
cc_80 N_C_M1000_g N_A_29_55#_c_222_n 0.0133379f $X=0.88 $Y=2.615 $X2=0 $Y2=0
cc_81 N_C_M1000_g N_A_29_55#_c_224_n 0.0104611f $X=0.88 $Y=2.615 $X2=0 $Y2=0
cc_82 N_C_c_69_n N_A_29_55#_c_224_n 0.0130804f $X=0.682 $Y=1.865 $X2=0 $Y2=0
cc_83 C N_A_29_55#_c_224_n 0.0247642f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_84 N_C_M1000_g N_VPWR_c_297_n 0.00465413f $X=0.88 $Y=2.615 $X2=0 $Y2=0
cc_85 N_C_M1000_g N_VPWR_c_295_n 0.00503886f $X=0.88 $Y=2.615 $X2=0 $Y2=0
cc_86 N_C_M1001_g N_VGND_c_343_n 0.010068f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_87 C N_VGND_c_343_n 0.00118332f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_88 N_C_M1001_g N_VGND_c_344_n 0.00525707f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_89 N_C_M1001_g N_VGND_c_345_n 0.0115483f $X=0.485 $Y=0.485 $X2=0 $Y2=0
cc_90 C N_VGND_c_345_n 0.02485f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_91 N_C_c_66_n N_VGND_c_345_n 9.46285e-19 $X=0.64 $Y=1.245 $X2=0 $Y2=0
cc_92 N_B_c_101_n N_A_M1004_g 0.0175882f $X=1.237 $Y=0.805 $X2=0 $Y2=0
cc_93 B N_A_M1004_g 8.28864e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_94 B N_A_M1004_g 5.14719e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_95 N_B_c_106_n N_A_M1004_g 0.00667442f $X=1.18 $Y=0.97 $X2=0 $Y2=0
cc_96 N_B_M1002_g N_A_c_159_n 0.00989004f $X=1.24 $Y=2.615 $X2=0 $Y2=0
cc_97 B N_A_c_159_n 7.2067e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_98 N_B_c_107_n N_A_c_159_n 0.00767192f $X=1.18 $Y=1.475 $X2=0 $Y2=0
cc_99 N_B_M1002_g N_A_c_164_n 0.0793505f $X=1.24 $Y=2.615 $X2=0 $Y2=0
cc_100 B N_A_c_164_n 0.00103259f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_101 N_B_M1002_g A 8.67867e-19 $X=1.24 $Y=2.615 $X2=0 $Y2=0
cc_102 B A 0.0546068f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B_c_106_n A 9.17992e-19 $X=1.18 $Y=0.97 $X2=0 $Y2=0
cc_104 B N_A_c_161_n 7.2067e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B_c_106_n N_A_c_161_n 0.00767192f $X=1.18 $Y=0.97 $X2=0 $Y2=0
cc_106 N_B_M1002_g N_A_29_55#_c_221_n 0.00220688f $X=1.24 $Y=2.615 $X2=0 $Y2=0
cc_107 N_B_M1002_g N_A_29_55#_c_222_n 0.0144337f $X=1.24 $Y=2.615 $X2=0 $Y2=0
cc_108 B N_A_29_55#_c_222_n 0.0257162f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_109 N_B_c_107_n N_A_29_55#_c_222_n 0.00107216f $X=1.18 $Y=1.475 $X2=0 $Y2=0
cc_110 N_B_c_101_n N_A_29_55#_c_211_n 0.00319289f $X=1.237 $Y=0.805 $X2=0 $Y2=0
cc_111 B N_A_29_55#_c_211_n 0.00110604f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_112 N_B_c_102_n N_A_29_55#_c_213_n 0.00137494f $X=1.237 $Y=0.955 $X2=0 $Y2=0
cc_113 B N_A_29_55#_c_213_n 0.0153978f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_114 N_B_c_106_n N_A_29_55#_c_213_n 4.55857e-19 $X=1.18 $Y=0.97 $X2=0 $Y2=0
cc_115 N_B_M1002_g N_A_29_55#_c_224_n 6.15616e-19 $X=1.24 $Y=2.615 $X2=0 $Y2=0
cc_116 B N_A_29_55#_c_216_n 0.00181963f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B_M1002_g N_VPWR_c_296_n 0.00274851f $X=1.24 $Y=2.615 $X2=0 $Y2=0
cc_118 N_B_M1002_g N_VPWR_c_297_n 0.00484506f $X=1.24 $Y=2.615 $X2=0 $Y2=0
cc_119 N_B_M1002_g N_VPWR_c_295_n 0.00503886f $X=1.24 $Y=2.615 $X2=0 $Y2=0
cc_120 N_B_c_101_n N_VGND_c_340_n 0.00545548f $X=1.237 $Y=0.805 $X2=0 $Y2=0
cc_121 N_B_c_101_n N_VGND_c_343_n 0.0113125f $X=1.237 $Y=0.805 $X2=0 $Y2=0
cc_122 N_B_c_102_n N_VGND_c_343_n 2.74929e-19 $X=1.237 $Y=0.955 $X2=0 $Y2=0
cc_123 B N_VGND_c_343_n 9.15461e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_124 N_B_c_101_n N_VGND_c_345_n 0.00368071f $X=1.237 $Y=0.805 $X2=0 $Y2=0
cc_125 N_B_c_102_n N_VGND_c_345_n 0.00292241f $X=1.237 $Y=0.955 $X2=0 $Y2=0
cc_126 B N_VGND_c_345_n 0.0202759f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_127 N_A_M1004_g N_A_29_55#_M1006_g 0.028566f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_128 A N_A_29_55#_M1006_g 3.04204e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_129 N_A_c_161_n N_A_29_55#_M1006_g 0.0167474f $X=1.75 $Y=1.36 $X2=0 $Y2=0
cc_130 N_A_M1003_g N_A_29_55#_M1005_g 0.00569538f $X=1.6 $Y=2.615 $X2=0 $Y2=0
cc_131 N_A_M1003_g N_A_29_55#_c_218_n 0.00780698f $X=1.6 $Y=2.615 $X2=0 $Y2=0
cc_132 N_A_c_164_n N_A_29_55#_c_218_n 0.00994981f $X=1.72 $Y=1.865 $X2=0 $Y2=0
cc_133 N_A_M1003_g N_A_29_55#_c_222_n 0.0154867f $X=1.6 $Y=2.615 $X2=0 $Y2=0
cc_134 N_A_c_164_n N_A_29_55#_c_222_n 0.00448187f $X=1.72 $Y=1.865 $X2=0 $Y2=0
cc_135 A N_A_29_55#_c_222_n 0.0241248f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 N_A_M1004_g N_A_29_55#_c_211_n 0.00344968f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_137 N_A_M1004_g N_A_29_55#_c_212_n 0.0139907f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_138 A N_A_29_55#_c_212_n 0.00727954f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A_c_161_n N_A_29_55#_c_212_n 0.00108035f $X=1.75 $Y=1.36 $X2=0 $Y2=0
cc_140 A N_A_29_55#_c_213_n 0.0169798f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A_c_161_n N_A_29_55#_c_213_n 0.00111374f $X=1.75 $Y=1.36 $X2=0 $Y2=0
cc_142 N_A_M1003_g N_A_29_55#_c_223_n 0.00352967f $X=1.6 $Y=2.615 $X2=0 $Y2=0
cc_143 N_A_c_164_n N_A_29_55#_c_223_n 0.00152381f $X=1.72 $Y=1.865 $X2=0 $Y2=0
cc_144 N_A_c_159_n N_A_29_55#_c_214_n 0.00152381f $X=1.72 $Y=1.685 $X2=0 $Y2=0
cc_145 N_A_c_159_n N_A_29_55#_c_215_n 0.00994981f $X=1.72 $Y=1.685 $X2=0 $Y2=0
cc_146 A N_A_29_55#_c_215_n 2.87721e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A_M1004_g N_A_29_55#_c_216_n 0.00349731f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_148 A N_A_29_55#_c_216_n 0.0492434f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A_c_161_n N_A_29_55#_c_216_n 0.00152381f $X=1.75 $Y=1.36 $X2=0 $Y2=0
cc_150 N_A_M1003_g N_VPWR_c_296_n 0.0145386f $X=1.6 $Y=2.615 $X2=0 $Y2=0
cc_151 N_A_M1003_g N_VPWR_c_297_n 0.00451101f $X=1.6 $Y=2.615 $X2=0 $Y2=0
cc_152 N_A_M1003_g N_VPWR_c_295_n 0.00473652f $X=1.6 $Y=2.615 $X2=0 $Y2=0
cc_153 N_A_M1004_g N_VGND_c_339_n 0.00171923f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_154 N_A_M1004_g N_VGND_c_340_n 0.00545548f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_155 N_A_M1004_g N_VGND_c_343_n 0.00583769f $X=1.815 $Y=0.485 $X2=0 $Y2=0
cc_156 N_A_29_55#_M1005_g N_VPWR_c_296_n 0.00490388f $X=2.37 $Y=2.725 $X2=0
+ $Y2=0
cc_157 N_A_29_55#_c_219_n N_VPWR_c_296_n 9.70101e-19 $X=2.29 $Y=2.215 $X2=0
+ $Y2=0
cc_158 N_A_29_55#_c_222_n N_VPWR_c_296_n 0.0507877f $X=2.015 $Y=2.125 $X2=0
+ $Y2=0
cc_159 N_A_29_55#_c_221_n N_VPWR_c_297_n 0.00685849f $X=0.665 $Y=2.615 $X2=0
+ $Y2=0
cc_160 N_A_29_55#_M1005_g N_VPWR_c_298_n 0.00502664f $X=2.37 $Y=2.725 $X2=0
+ $Y2=0
cc_161 N_A_29_55#_M1005_g N_VPWR_c_295_n 0.0109583f $X=2.37 $Y=2.725 $X2=0 $Y2=0
cc_162 N_A_29_55#_c_221_n N_VPWR_c_295_n 0.0103555f $X=0.665 $Y=2.615 $X2=0
+ $Y2=0
cc_163 N_A_29_55#_M1006_g X 0.0198613f $X=2.245 $Y=0.485 $X2=0 $Y2=0
cc_164 N_A_29_55#_M1005_g X 0.00653711f $X=2.37 $Y=2.725 $X2=0 $Y2=0
cc_165 N_A_29_55#_c_222_n X 0.0147515f $X=2.015 $Y=2.125 $X2=0 $Y2=0
cc_166 N_A_29_55#_c_212_n X 0.00868429f $X=2.015 $Y=0.912 $X2=0 $Y2=0
cc_167 N_A_29_55#_c_214_n X 0.0380673f $X=2.29 $Y=1.71 $X2=0 $Y2=0
cc_168 N_A_29_55#_c_215_n X 0.0166275f $X=2.29 $Y=1.71 $X2=0 $Y2=0
cc_169 N_A_29_55#_c_216_n X 0.0227876f $X=2.195 $Y=1.545 $X2=0 $Y2=0
cc_170 N_A_29_55#_M1005_g X 0.00582711f $X=2.37 $Y=2.725 $X2=0 $Y2=0
cc_171 N_A_29_55#_M1005_g X 0.00363586f $X=2.37 $Y=2.725 $X2=0 $Y2=0
cc_172 N_A_29_55#_c_219_n X 4.76781e-19 $X=2.29 $Y=2.215 $X2=0 $Y2=0
cc_173 N_A_29_55#_M1006_g N_VGND_c_339_n 0.00318537f $X=2.245 $Y=0.485 $X2=0
+ $Y2=0
cc_174 N_A_29_55#_c_212_n N_VGND_c_339_n 0.0179645f $X=2.015 $Y=0.912 $X2=0
+ $Y2=0
cc_175 N_A_29_55#_c_211_n N_VGND_c_340_n 0.0105858f $X=1.6 $Y=0.485 $X2=0 $Y2=0
cc_176 N_A_29_55#_M1006_g N_VGND_c_342_n 0.00545548f $X=2.245 $Y=0.485 $X2=0
+ $Y2=0
cc_177 N_A_29_55#_M1006_g N_VGND_c_343_n 0.0106753f $X=2.245 $Y=0.485 $X2=0
+ $Y2=0
cc_178 N_A_29_55#_c_210_n N_VGND_c_343_n 0.0104489f $X=0.27 $Y=0.485 $X2=0 $Y2=0
cc_179 N_A_29_55#_c_211_n N_VGND_c_343_n 0.00969948f $X=1.6 $Y=0.485 $X2=0 $Y2=0
cc_180 N_A_29_55#_c_212_n N_VGND_c_343_n 0.00680297f $X=2.015 $Y=0.912 $X2=0
+ $Y2=0
cc_181 N_A_29_55#_c_210_n N_VGND_c_344_n 0.013063f $X=0.27 $Y=0.485 $X2=0 $Y2=0
cc_182 N_VPWR_c_298_n X 0.0250662f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_295_n X 0.014322f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_296_n X 0.0277049f $X=2.155 $Y=2.55 $X2=0 $Y2=0
cc_185 N_X_c_320_n N_VGND_c_342_n 0.02096f $X=2.67 $Y=0.485 $X2=0 $Y2=0
cc_186 N_X_c_320_n N_VGND_c_343_n 0.017086f $X=2.67 $Y=0.485 $X2=0 $Y2=0
