# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o31ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o31ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.940000 1.425000 2.290000 1.595000 ;
        RECT 1.485000 1.595000 1.835000 1.760000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.330000 1.075000 2.985000 1.245000 ;
        RECT 0.330000 1.245000 0.660000 1.515000 ;
        RECT 2.460000 1.245000 2.985000 1.325000 ;
        RECT 2.460000 1.325000 3.670000 1.505000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.985000 1.325000 5.005000 1.695000 ;
        RECT 3.985000 1.695000 7.280000 1.865000 ;
        RECT 7.110000 1.335000 7.720000 1.535000 ;
        RECT 7.110000 1.535000 7.280000 1.695000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.240000 1.345000 6.930000 1.525000 ;
        RECT 5.435000 1.200000 6.575000 1.345000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  2.318400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.145000 2.035000 7.630000 2.215000 ;
        RECT 4.145000 2.215000 4.335000 2.735000 ;
        RECT 5.005000 2.215000 7.630000 2.240000 ;
        RECT 5.005000 2.240000 5.185000 2.725000 ;
        RECT 5.465000 0.700000 6.925000 0.995000 ;
        RECT 5.465000 0.995000 8.075000 1.030000 ;
        RECT 6.745000 1.030000 8.075000 1.165000 ;
        RECT 7.335000 2.240000 7.630000 2.715000 ;
        RECT 7.460000 1.705000 8.075000 1.875000 ;
        RECT 7.460000 1.875000 7.630000 2.035000 ;
        RECT 7.890000 1.165000 8.075000 1.705000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.205000  0.085000 0.465000 0.905000 ;
      RECT 0.205000  1.815000 1.315000 1.930000 ;
      RECT 0.205000  1.930000 3.075000 1.985000 ;
      RECT 0.205000  1.985000 0.465000 3.075000 ;
      RECT 0.635000  0.255000 0.895000 0.735000 ;
      RECT 0.635000  0.735000 3.475000 0.905000 ;
      RECT 0.635000  2.155000 0.965000 2.270000 ;
      RECT 0.635000  2.270000 2.685000 2.440000 ;
      RECT 0.635000  2.440000 0.965000 3.075000 ;
      RECT 1.065000  0.085000 1.395000 0.565000 ;
      RECT 1.135000  2.610000 1.325000 3.245000 ;
      RECT 1.145000  1.985000 2.175000 2.100000 ;
      RECT 1.495000  2.440000 1.825000 3.075000 ;
      RECT 1.565000  0.255000 1.755000 0.735000 ;
      RECT 1.925000  0.085000 2.255000 0.565000 ;
      RECT 1.995000  2.610000 2.185000 3.245000 ;
      RECT 2.005000  1.815000 3.815000 1.875000 ;
      RECT 2.005000  1.875000 3.075000 1.930000 ;
      RECT 2.355000  2.155000 2.685000 2.270000 ;
      RECT 2.355000  2.440000 2.685000 2.885000 ;
      RECT 2.355000  2.885000 3.475000 3.075000 ;
      RECT 2.425000  0.255000 2.615000 0.735000 ;
      RECT 2.785000  0.085000 3.115000 0.565000 ;
      RECT 2.855000  1.985000 3.075000 2.715000 ;
      RECT 2.865000  1.705000 3.815000 1.815000 ;
      RECT 3.245000  2.055000 3.475000 2.885000 ;
      RECT 3.275000  0.905000 3.475000 0.985000 ;
      RECT 3.275000  0.985000 5.265000 1.155000 ;
      RECT 3.285000  0.255000 3.475000 0.735000 ;
      RECT 3.645000  0.085000 3.975000 0.805000 ;
      RECT 3.645000  1.875000 3.815000 2.035000 ;
      RECT 3.645000  2.035000 3.975000 2.905000 ;
      RECT 3.645000  2.905000 5.525000 3.075000 ;
      RECT 4.155000  0.425000 4.380000 0.985000 ;
      RECT 4.505000  2.385000 4.835000 2.895000 ;
      RECT 4.505000  2.895000 5.525000 2.905000 ;
      RECT 4.550000  0.085000 4.880000 0.805000 ;
      RECT 5.065000  0.255000 7.425000 0.530000 ;
      RECT 5.065000  0.530000 5.265000 0.985000 ;
      RECT 5.355000  2.410000 7.165000 2.580000 ;
      RECT 5.355000  2.580000 5.525000 2.895000 ;
      RECT 5.695000  2.750000 5.905000 3.245000 ;
      RECT 6.555000  2.750000 6.825000 3.245000 ;
      RECT 6.995000  2.580000 7.165000 2.895000 ;
      RECT 6.995000  2.895000 8.060000 3.065000 ;
      RECT 7.095000  0.530000 7.425000 0.825000 ;
      RECT 7.605000  0.085000 7.935000 0.825000 ;
      RECT 7.800000  2.045000 8.060000 2.895000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__o31ai_4
END LIBRARY
