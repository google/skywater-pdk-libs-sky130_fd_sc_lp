* NGSPICE file created from sky130_fd_sc_lp__sdlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 VPWR a_742_107# a_1235_429# VPB phighvt w=640000u l=150000u
+  ad=1.9983e+12p pd=1.668e+07u as=1.792e+11p ps=1.84e+06u
M1001 VGND a_1235_429# GCLK VNB nshort w=840000u l=150000u
+  ad=1.1701e+12p pd=1.139e+07u as=2.352e+11p ps=2.24e+06u
M1002 a_614_133# a_282_70# a_110_70# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.809e+11p ps=3.18e+06u
M1003 VPWR CLK a_250_443# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1004 VPWR a_1235_429# GCLK VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1005 a_110_70# SCE VGND VNB nshort w=420000u l=150000u
+  ad=2.709e+11p pd=2.97e+06u as=0p ps=0u
M1006 a_1174_74# CLK VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 a_282_70# a_250_443# VPWR VPB phighvt w=640000u l=150000u
+  ad=3.136e+11p pd=2.26e+06u as=0p ps=0u
M1008 a_1235_429# a_742_107# a_1174_74# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1009 GCLK a_1235_429# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND GATE a_110_70# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_742_107# a_746_457# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1012 GCLK a_1235_429# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_742_107# a_700_133# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1014 a_614_133# a_250_443# a_110_70# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1015 a_700_133# a_282_70# a_614_133# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_742_107# a_614_133# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1017 a_110_70# GATE a_110_468# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1018 a_746_457# a_250_443# a_614_133# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_742_107# a_614_133# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1020 a_282_70# a_250_443# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1021 a_110_468# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1235_429# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND CLK a_250_443# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

