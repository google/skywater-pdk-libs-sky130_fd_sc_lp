* File: sky130_fd_sc_lp__isobufsrc_2.spice
* Created: Wed Sep  2 09:58:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__isobufsrc_2.pex.spice"
.subckt sky130_fd_sc_lp__isobufsrc_2  VNB VPB A SLEEP VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_40_131#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.182 AS=0.1113 PD=1.02333 PS=1.37 NRD=108.084 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1001_d N_SLEEP_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.364 AS=0.1176 PD=2.04667 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.8
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_40_131#_M1004_g N_X_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1004_d N_A_40_131#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_SLEEP_M1007_g N_X_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_40_131#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1003_d N_SLEEP_M1008_g N_A_283_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=4.9447 NRS=0 M=1 R=8.4
+ SA=75000.4 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1002 N_A_283_367#_M1008_s N_A_40_131#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_A_283_367#_M1005_d N_A_40_131#_M1005_g N_X_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_SLEEP_M1009_g N_A_283_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__isobufsrc_2.pxi.spice"
*
.ends
*
*
