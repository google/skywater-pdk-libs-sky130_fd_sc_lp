* File: sky130_fd_sc_lp__o21a_2.pxi.spice
* Created: Fri Aug 28 11:03:49 2020
* 
x_PM_SKY130_FD_SC_LP__O21A_2%A_86_21# N_A_86_21#_M1000_s N_A_86_21#_M1001_d
+ N_A_86_21#_c_59_n N_A_86_21#_M1004_g N_A_86_21#_M1003_g N_A_86_21#_c_61_n
+ N_A_86_21#_M1005_g N_A_86_21#_M1008_g N_A_86_21#_c_63_n N_A_86_21#_c_64_n
+ N_A_86_21#_c_65_n N_A_86_21#_c_77_p N_A_86_21#_c_95_p N_A_86_21#_c_66_n
+ N_A_86_21#_c_87_p N_A_86_21#_c_88_p N_A_86_21#_c_67_n N_A_86_21#_c_68_n
+ N_A_86_21#_c_69_n PM_SKY130_FD_SC_LP__O21A_2%A_86_21#
x_PM_SKY130_FD_SC_LP__O21A_2%B1 N_B1_M1000_g N_B1_M1001_g B1 N_B1_c_133_n
+ N_B1_c_134_n PM_SKY130_FD_SC_LP__O21A_2%B1
x_PM_SKY130_FD_SC_LP__O21A_2%A2 N_A2_M1006_g N_A2_M1009_g A2 A2 N_A2_c_168_n
+ PM_SKY130_FD_SC_LP__O21A_2%A2
x_PM_SKY130_FD_SC_LP__O21A_2%A1 N_A1_M1002_g N_A1_M1007_g A1 N_A1_c_202_n
+ N_A1_c_203_n PM_SKY130_FD_SC_LP__O21A_2%A1
x_PM_SKY130_FD_SC_LP__O21A_2%VPWR N_VPWR_M1003_s N_VPWR_M1008_s N_VPWR_M1007_d
+ N_VPWR_c_226_n N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n N_VPWR_c_230_n
+ VPWR N_VPWR_c_231_n N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_225_n
+ PM_SKY130_FD_SC_LP__O21A_2%VPWR
x_PM_SKY130_FD_SC_LP__O21A_2%X N_X_M1004_d N_X_M1003_d X X X X X X X N_X_c_269_n
+ PM_SKY130_FD_SC_LP__O21A_2%X
x_PM_SKY130_FD_SC_LP__O21A_2%VGND N_VGND_M1004_s N_VGND_M1005_s N_VGND_M1006_d
+ N_VGND_c_288_n N_VGND_c_289_n N_VGND_c_290_n N_VGND_c_291_n N_VGND_c_292_n
+ N_VGND_c_293_n VGND N_VGND_c_294_n N_VGND_c_295_n N_VGND_c_296_n
+ N_VGND_c_297_n PM_SKY130_FD_SC_LP__O21A_2%VGND
x_PM_SKY130_FD_SC_LP__O21A_2%A_392_51# N_A_392_51#_M1000_d N_A_392_51#_M1002_d
+ N_A_392_51#_c_331_n N_A_392_51#_c_332_n N_A_392_51#_c_333_n
+ N_A_392_51#_c_334_n PM_SKY130_FD_SC_LP__O21A_2%A_392_51#
cc_1 VNB N_A_86_21#_c_59_n 0.0210929f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.185
cc_2 VNB N_A_86_21#_M1003_g 0.0243375f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_3 VNB N_A_86_21#_c_61_n 0.0191409f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.185
cc_4 VNB N_A_86_21#_M1008_g 0.0082135f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_5 VNB N_A_86_21#_c_63_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.26
cc_6 VNB N_A_86_21#_c_64_n 0.00183148f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.92
cc_7 VNB N_A_86_21#_c_65_n 0.0141068f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=1.16
cc_8 VNB N_A_86_21#_c_66_n 0.0101465f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=0.42
cc_9 VNB N_A_86_21#_c_67_n 0.00586784f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.16
cc_10 VNB N_A_86_21#_c_68_n 0.0435092f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.35
cc_11 VNB N_A_86_21#_c_69_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.35
cc_12 VNB N_B1_M1000_g 0.0280604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_c_133_n 0.0296347f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_14 VNB N_B1_c_134_n 0.00234774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_M1006_g 0.0233535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A2 0.00479519f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.335
cc_17 VNB N_A2_c_168_n 0.0218524f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.26
cc_18 VNB N_A1_M1002_g 0.0274056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1007_g 0.00137316f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.185
cc_20 VNB N_A1_c_202_n 0.0552217f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=1.26
cc_21 VNB N_A1_c_203_n 0.0122352f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.26
cc_22 VNB N_VPWR_c_225_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.35
cc_23 VNB N_X_c_269_n 0.00293196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_288_n 0.0113784f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.335
cc_25 VNB N_VGND_c_289_n 0.048097f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_26 VNB N_VGND_c_290_n 0.00911982f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.185
cc_27 VNB N_VGND_c_291_n 0.00100404f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_28 VNB N_VGND_c_292_n 0.0280283f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.26
cc_29 VNB N_VGND_c_293_n 0.00463869f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.52
cc_30 VNB N_VGND_c_294_n 0.0152106f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.16
cc_31 VNB N_VGND_c_295_n 0.019138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_296_n 0.209678f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.16
cc_33 VNB N_VGND_c_297_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=2.135 $Y2=2.005
cc_34 VNB N_A_392_51#_c_331_n 0.00120843f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_35 VNB N_A_392_51#_c_332_n 0.0121897f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_36 VNB N_A_392_51#_c_333_n 0.00610995f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_37 VNB N_A_392_51#_c_334_n 0.0313753f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.26
cc_38 VPB N_A_86_21#_M1003_g 0.0265098f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_39 VPB N_A_86_21#_M1008_g 0.0224337f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_40 VPB N_A_86_21#_c_64_n 0.00394301f $X=-0.19 $Y=1.655 $X2=1.23 $Y2=1.92
cc_41 VPB N_B1_M1001_g 0.022563f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.185
cc_42 VPB N_B1_c_133_n 0.00860237f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_43 VPB N_B1_c_134_n 0.0036885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A2_M1009_g 0.0189888f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.185
cc_45 VPB A2 0.0143034f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.335
cc_46 VPB N_A2_c_168_n 0.00625343f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=1.26
cc_47 VPB N_A1_M1007_g 0.0246659f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.185
cc_48 VPB N_A1_c_203_n 0.0107005f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.26
cc_49 VPB N_VPWR_c_226_n 0.0113525f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.335
cc_50 VPB N_VPWR_c_227_n 0.0639754f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_51 VPB N_VPWR_c_228_n 0.0028356f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.655
cc_52 VPB N_VPWR_c_229_n 0.0135296f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_53 VPB N_VPWR_c_230_n 0.0483425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_231_n 0.0152106f $X=-0.19 $Y=1.655 $X2=2.005 $Y2=2.005
cc_55 VPB N_VPWR_c_232_n 0.0271101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_233_n 0.0138973f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.35
cc_57 VPB N_VPWR_c_225_n 0.0488403f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=1.35
cc_58 VPB N_X_c_269_n 0.00164967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 N_A_86_21#_c_65_n N_B1_M1000_g 0.00373845f $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_86_21#_c_67_n N_B1_M1000_g 5.36613e-19 $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_86_21#_c_68_n N_B1_M1000_g 0.00388882f $X=1.15 $Y=1.35 $X2=0 $Y2=0
cc_62 N_A_86_21#_c_64_n N_B1_M1001_g 0.00439017f $X=1.23 $Y=1.92 $X2=0 $Y2=0
cc_63 N_A_86_21#_c_77_p N_B1_M1001_g 0.0162049f $X=2.005 $Y=2.005 $X2=0 $Y2=0
cc_64 N_A_86_21#_M1008_g N_B1_c_133_n 0.00227391f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_65 N_A_86_21#_c_65_n N_B1_c_133_n 0.00595557f $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_86_21#_c_77_p N_B1_c_133_n 0.00130692f $X=2.005 $Y=2.005 $X2=0 $Y2=0
cc_67 N_A_86_21#_c_67_n N_B1_c_133_n 0.0011067f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_86_21#_c_68_n N_B1_c_133_n 0.0092217f $X=1.15 $Y=1.35 $X2=0 $Y2=0
cc_69 N_A_86_21#_c_65_n N_B1_c_134_n 0.0267489f $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A_86_21#_c_77_p N_B1_c_134_n 0.0293656f $X=2.005 $Y=2.005 $X2=0 $Y2=0
cc_71 N_A_86_21#_c_67_n N_B1_c_134_n 0.0269918f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_86_21#_c_68_n N_B1_c_134_n 6.57094e-19 $X=1.15 $Y=1.35 $X2=0 $Y2=0
cc_73 N_A_86_21#_c_87_p N_A2_M1009_g 0.00346817f $X=2.135 $Y=2.09 $X2=0 $Y2=0
cc_74 N_A_86_21#_c_88_p N_A2_M1009_g 0.0193749f $X=2.1 $Y=2.45 $X2=0 $Y2=0
cc_75 N_A_86_21#_c_87_p A2 0.0147275f $X=2.135 $Y=2.09 $X2=0 $Y2=0
cc_76 N_A_86_21#_c_87_p N_A2_c_168_n 3.07128e-19 $X=2.135 $Y=2.09 $X2=0 $Y2=0
cc_77 N_A_86_21#_c_87_p N_A1_M1007_g 5.12803e-19 $X=2.135 $Y=2.09 $X2=0 $Y2=0
cc_78 N_A_86_21#_c_88_p N_A1_M1007_g 0.00298475f $X=2.1 $Y=2.45 $X2=0 $Y2=0
cc_79 N_A_86_21#_c_64_n N_VPWR_M1008_s 0.00298128f $X=1.23 $Y=1.92 $X2=0 $Y2=0
cc_80 N_A_86_21#_c_77_p N_VPWR_M1008_s 0.0134411f $X=2.005 $Y=2.005 $X2=0 $Y2=0
cc_81 N_A_86_21#_c_95_p N_VPWR_M1008_s 0.00536166f $X=1.315 $Y=2.005 $X2=0 $Y2=0
cc_82 N_A_86_21#_M1003_g N_VPWR_c_227_n 0.00741603f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_83 N_A_86_21#_M1003_g N_VPWR_c_228_n 7.66174e-19 $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_84 N_A_86_21#_M1008_g N_VPWR_c_228_n 0.0192268f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_86_21#_c_77_p N_VPWR_c_228_n 0.0373846f $X=2.005 $Y=2.005 $X2=0 $Y2=0
cc_86 N_A_86_21#_c_95_p N_VPWR_c_228_n 0.0152373f $X=1.315 $Y=2.005 $X2=0 $Y2=0
cc_87 N_A_86_21#_c_87_p N_VPWR_c_230_n 0.00499344f $X=2.135 $Y=2.09 $X2=0 $Y2=0
cc_88 N_A_86_21#_c_88_p N_VPWR_c_230_n 0.026783f $X=2.1 $Y=2.45 $X2=0 $Y2=0
cc_89 N_A_86_21#_M1003_g N_VPWR_c_231_n 0.00564131f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_90 N_A_86_21#_M1008_g N_VPWR_c_231_n 0.00486043f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_91 N_A_86_21#_c_88_p N_VPWR_c_232_n 0.015688f $X=2.1 $Y=2.45 $X2=0 $Y2=0
cc_92 N_A_86_21#_M1001_d N_VPWR_c_225_n 0.00380103f $X=1.96 $Y=1.835 $X2=0 $Y2=0
cc_93 N_A_86_21#_M1003_g N_VPWR_c_225_n 0.0110687f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_86_21#_M1008_g N_VPWR_c_225_n 0.00824727f $X=0.935 $Y=2.465 $X2=0
+ $Y2=0
cc_95 N_A_86_21#_c_88_p N_VPWR_c_225_n 0.00984745f $X=2.1 $Y=2.45 $X2=0 $Y2=0
cc_96 N_A_86_21#_c_59_n N_X_c_269_n 0.0142786f $X=0.505 $Y=1.185 $X2=0 $Y2=0
cc_97 N_A_86_21#_M1003_g N_X_c_269_n 0.0384592f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_86_21#_c_61_n N_X_c_269_n 0.00132211f $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_99 N_A_86_21#_c_63_n N_X_c_269_n 0.00619566f $X=0.505 $Y=1.26 $X2=0 $Y2=0
cc_100 N_A_86_21#_c_64_n N_X_c_269_n 0.0172141f $X=1.23 $Y=1.92 $X2=0 $Y2=0
cc_101 N_A_86_21#_c_67_n N_X_c_269_n 0.0337447f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_86_21#_c_68_n N_X_c_269_n 0.00534016f $X=1.15 $Y=1.35 $X2=0 $Y2=0
cc_103 N_A_86_21#_c_69_n N_X_c_269_n 0.0101971f $X=0.86 $Y=1.35 $X2=0 $Y2=0
cc_104 N_A_86_21#_c_67_n N_VGND_M1005_s 0.00291336f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_86_21#_c_59_n N_VGND_c_289_n 0.00682857f $X=0.505 $Y=1.185 $X2=0
+ $Y2=0
cc_106 N_A_86_21#_c_59_n N_VGND_c_290_n 7.12485e-19 $X=0.505 $Y=1.185 $X2=0
+ $Y2=0
cc_107 N_A_86_21#_c_61_n N_VGND_c_290_n 0.0130972f $X=0.935 $Y=1.185 $X2=0 $Y2=0
cc_108 N_A_86_21#_c_66_n N_VGND_c_290_n 0.0496305f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_109 N_A_86_21#_c_67_n N_VGND_c_290_n 0.0265319f $X=1.15 $Y=1.16 $X2=0 $Y2=0
cc_110 N_A_86_21#_c_68_n N_VGND_c_290_n 0.0016889f $X=1.15 $Y=1.35 $X2=0 $Y2=0
cc_111 N_A_86_21#_c_66_n N_VGND_c_292_n 0.0190529f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_112 N_A_86_21#_c_59_n N_VGND_c_294_n 0.00564131f $X=0.505 $Y=1.185 $X2=0
+ $Y2=0
cc_113 N_A_86_21#_c_61_n N_VGND_c_294_n 0.00486043f $X=0.935 $Y=1.185 $X2=0
+ $Y2=0
cc_114 N_A_86_21#_c_59_n N_VGND_c_296_n 0.0110687f $X=0.505 $Y=1.185 $X2=0 $Y2=0
cc_115 N_A_86_21#_c_61_n N_VGND_c_296_n 0.00824727f $X=0.935 $Y=1.185 $X2=0
+ $Y2=0
cc_116 N_A_86_21#_c_66_n N_VGND_c_296_n 0.0113912f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_117 N_A_86_21#_c_65_n N_A_392_51#_c_333_n 0.00995284f $X=1.505 $Y=1.16 $X2=0
+ $Y2=0
cc_118 N_B1_M1000_g N_A2_M1006_g 0.022626f $X=1.885 $Y=0.675 $X2=0 $Y2=0
cc_119 N_B1_M1001_g N_A2_M1009_g 0.0188385f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B1_c_133_n A2 0.00351184f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_121 N_B1_c_134_n A2 0.0285163f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_122 N_B1_c_133_n N_A2_c_168_n 0.0211119f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_123 N_B1_c_134_n N_A2_c_168_n 2.37249e-19 $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_124 N_B1_M1001_g N_VPWR_c_228_n 0.0194392f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B1_M1001_g N_VPWR_c_232_n 0.00486043f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B1_M1001_g N_VPWR_c_225_n 0.0082726f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B1_M1000_g N_VGND_c_290_n 0.00318815f $X=1.885 $Y=0.675 $X2=0 $Y2=0
cc_128 N_B1_M1000_g N_VGND_c_291_n 0.00110103f $X=1.885 $Y=0.675 $X2=0 $Y2=0
cc_129 N_B1_M1000_g N_VGND_c_292_n 0.00565115f $X=1.885 $Y=0.675 $X2=0 $Y2=0
cc_130 N_B1_M1000_g N_VGND_c_296_n 0.0119838f $X=1.885 $Y=0.675 $X2=0 $Y2=0
cc_131 N_B1_M1000_g N_A_392_51#_c_333_n 9.70773e-19 $X=1.885 $Y=0.675 $X2=0
+ $Y2=0
cc_132 N_A2_M1006_g N_A1_M1002_g 0.0199943f $X=2.315 $Y=0.675 $X2=0 $Y2=0
cc_133 N_A2_M1009_g N_A1_M1007_g 0.0568391f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_134 A2 N_A1_M1007_g 0.00394011f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_135 A2 N_A1_c_202_n 0.00676517f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A2_c_168_n N_A1_c_202_n 0.0217817f $X=2.335 $Y=1.51 $X2=0 $Y2=0
cc_137 A2 N_A1_c_203_n 0.0304592f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A2_M1009_g N_VPWR_c_228_n 0.00141541f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A2_M1009_g N_VPWR_c_230_n 0.00456699f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A2_M1009_g N_VPWR_c_232_n 0.0054895f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A2_M1009_g N_VPWR_c_225_n 0.0101742f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A2_M1006_g N_VGND_c_291_n 0.00956826f $X=2.315 $Y=0.675 $X2=0 $Y2=0
cc_143 N_A2_M1006_g N_VGND_c_292_n 0.00544562f $X=2.315 $Y=0.675 $X2=0 $Y2=0
cc_144 N_A2_M1006_g N_VGND_c_296_n 0.00951556f $X=2.315 $Y=0.675 $X2=0 $Y2=0
cc_145 N_A2_M1006_g N_A_392_51#_c_332_n 0.0140338f $X=2.315 $Y=0.675 $X2=0 $Y2=0
cc_146 A2 N_A_392_51#_c_332_n 0.0396557f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A2_c_168_n N_A_392_51#_c_332_n 0.00313303f $X=2.335 $Y=1.51 $X2=0 $Y2=0
cc_148 A2 N_A_392_51#_c_333_n 0.0132025f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_149 N_A2_c_168_n N_A_392_51#_c_333_n 0.00108693f $X=2.335 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A1_M1007_g N_VPWR_c_230_n 0.0319225f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A1_c_202_n N_VPWR_c_230_n 0.00147549f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_152 N_A1_c_203_n N_VPWR_c_230_n 0.0222559f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_153 N_A1_M1007_g N_VPWR_c_232_n 0.00486043f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A1_M1007_g N_VPWR_c_225_n 0.00848326f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A1_M1002_g N_VGND_c_291_n 0.0101494f $X=2.785 $Y=0.675 $X2=0 $Y2=0
cc_156 N_A1_M1002_g N_VGND_c_295_n 0.00544562f $X=2.785 $Y=0.675 $X2=0 $Y2=0
cc_157 N_A1_M1002_g N_VGND_c_296_n 0.0104285f $X=2.785 $Y=0.675 $X2=0 $Y2=0
cc_158 N_A1_M1002_g N_A_392_51#_c_332_n 0.0189639f $X=2.785 $Y=0.675 $X2=0 $Y2=0
cc_159 N_A1_c_202_n N_A_392_51#_c_332_n 0.00866875f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_160 N_A1_c_203_n N_A_392_51#_c_332_n 0.0221394f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_161 N_VPWR_c_225_n N_X_M1003_d 0.00380103f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_162 N_VPWR_c_227_n N_X_c_269_n 0.0460757f $X=0.29 $Y=1.98 $X2=0 $Y2=0
cc_163 N_VPWR_c_231_n N_X_c_269_n 0.0150063f $X=0.985 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VPWR_c_225_n N_X_c_269_n 0.00950443f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_165 N_VPWR_c_225_n A_478_367# 0.0137053f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_166 N_X_c_269_n N_VGND_c_289_n 0.0309728f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_167 N_X_c_269_n N_VGND_c_294_n 0.0150063f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_168 N_X_M1004_d N_VGND_c_296_n 0.00380103f $X=0.58 $Y=0.235 $X2=0 $Y2=0
cc_169 N_X_c_269_n N_VGND_c_296_n 0.00950443f $X=0.72 $Y=0.42 $X2=0 $Y2=0
cc_170 N_VGND_c_292_n N_A_392_51#_c_331_n 0.0144039f $X=2.385 $Y=0 $X2=0 $Y2=0
cc_171 N_VGND_c_296_n N_A_392_51#_c_331_n 0.00944728f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_172 N_VGND_M1006_d N_A_392_51#_c_332_n 0.00218982f $X=2.39 $Y=0.255 $X2=0
+ $Y2=0
cc_173 N_VGND_c_291_n N_A_392_51#_c_332_n 0.017285f $X=2.55 $Y=0.4 $X2=0 $Y2=0
cc_174 N_VGND_c_295_n N_A_392_51#_c_334_n 0.0185207f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_175 N_VGND_c_296_n N_A_392_51#_c_334_n 0.010808f $X=3.12 $Y=0 $X2=0 $Y2=0
