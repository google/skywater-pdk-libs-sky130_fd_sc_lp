* File: sky130_fd_sc_lp__dlrtn_2.pex.spice
* Created: Fri Aug 28 10:26:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRTN_2%D 3 7 9 10 11 12 13 14 19
c40 9 0 3.55661e-20 $X=0.55 $Y=0.88
r41 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.55
+ $Y=1.045 $X2=0.55 $Y2=1.045
r42 13 14 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.65 $Y=1.295
+ $X2=0.65 $Y2=1.665
r43 13 20 7.78678 $w=3.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.65 $Y=1.295
+ $X2=0.65 $Y2=1.045
r44 12 20 3.73765 $w=3.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.65 $Y=0.925
+ $X2=0.65 $Y2=1.045
r45 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.55 $Y=1.385
+ $X2=0.55 $Y2=1.045
r46 10 11 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.385
+ $X2=0.55 $Y2=1.55
r47 9 19 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=0.88
+ $X2=0.55 $Y2=1.045
r48 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.6 $Y=0.56 $X2=0.6
+ $Y2=0.88
r49 3 11 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=0.495 $Y=2.64
+ $X2=0.495 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%GATE_N 3 6 9 10 11 12 13 14 19
c49 12 0 3.55661e-20 $X=1.2 $Y=0.925
c50 9 0 1.07576e-19 $X=1.09 $Y=0.88
r51 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.09
+ $Y=1.045 $X2=1.09 $Y2=1.045
r52 13 14 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.665
r53 13 20 9.93485 $w=2.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.045
r54 12 20 4.76873 $w=2.88e-07 $l=1.2e-07 $layer=LI1_cond $X=1.15 $Y=0.925
+ $X2=1.15 $Y2=1.045
r55 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.09 $Y=1.385
+ $X2=1.09 $Y2=1.045
r56 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.385
+ $X2=1.09 $Y2=1.55
r57 9 19 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=0.88
+ $X2=1.09 $Y2=1.045
r58 6 11 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=1.18 $Y=2.64
+ $X2=1.18 $Y2=1.55
r59 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.03 $Y=0.56 $X2=1.03
+ $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%A_31_464# 1 2 9 13 17 18 20 23 25 28 29 30
+ 32 33 34 37 38 43 45
c114 34 0 1.93583e-19 $X=1.985 $Y=2.51
c115 9 0 3.63575e-20 $X=2.695 $Y=0.835
r116 40 43 6.91466 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.2 $Y=0.532
+ $X2=0.365 $Y2=0.532
r117 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.745
+ $Y=1.68 $X2=2.745 $Y2=1.68
r118 35 37 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=2.745 $Y=2.425
+ $X2=2.745 $Y2=1.68
r119 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.58 $Y=2.51
+ $X2=2.745 $Y2=2.425
r120 33 34 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.58 $Y=2.51
+ $X2=1.985 $Y2=2.51
r121 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.9 $Y=2.595
+ $X2=1.985 $Y2=2.51
r122 31 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.9 $Y=2.595
+ $X2=1.9 $Y2=2.81
r123 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.815 $Y=2.895
+ $X2=1.9 $Y2=2.81
r124 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.815 $Y=2.895
+ $X2=1.145 $Y2=2.895
r125 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=2.81
+ $X2=1.145 $Y2=2.895
r126 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.06 $Y=2.13
+ $X2=1.06 $Y2=2.81
r127 26 45 2.49072 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.41 $Y=2.045
+ $X2=0.262 $Y2=2.045
r128 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=2.045
+ $X2=1.06 $Y2=2.13
r129 25 26 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.975 $Y=2.045
+ $X2=0.41 $Y2=2.045
r130 21 45 3.95216 $w=2.32e-07 $l=8.5e-08 $layer=LI1_cond $X=0.262 $Y=2.13
+ $X2=0.262 $Y2=2.045
r131 21 23 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=0.262 $Y=2.13
+ $X2=0.262 $Y2=2.465
r132 20 45 3.95216 $w=2.32e-07 $l=1.11781e-07 $layer=LI1_cond $X=0.2 $Y=1.96
+ $X2=0.262 $Y2=2.045
r133 19 40 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.2 $Y=0.67 $X2=0.2
+ $Y2=0.532
r134 19 20 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=0.2 $Y=0.67
+ $X2=0.2 $Y2=1.96
r135 17 38 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.745 $Y=2.02
+ $X2=2.745 $Y2=1.68
r136 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=2.02
+ $X2=2.745 $Y2=2.185
r137 16 38 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.515
+ $X2=2.745 $Y2=1.68
r138 13 18 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.835 $Y=2.685
+ $X2=2.835 $Y2=2.185
r139 9 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.695 $Y=0.835
+ $X2=2.695 $Y2=1.515
r140 2 23 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.155
+ $Y=2.32 $X2=0.28 $Y2=2.465
r141 1 43 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.24
+ $Y=0.35 $X2=0.365 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%A_372_397# 1 2 9 13 14 16 19 20 22 23 25 27
+ 28 31 32 45
c107 20 0 3.63575e-20 $X=2.985 $Y=0.377
r108 35 36 18.905 $w=2.42e-07 $l=3.75e-07 $layer=LI1_cond $X=2.017 $Y=0.835
+ $X2=2.017 $Y2=1.21
r109 31 32 6.58732 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.985 $Y=2.15
+ $X2=1.985 $Y2=1.995
r110 28 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=2.04
+ $X2=3.285 $Y2=2.205
r111 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.285
+ $Y=2.04 $X2=3.285 $Y2=2.04
r112 25 37 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=1.21
+ $X2=2.9 $Y2=1.21
r113 25 27 33.0219 $w=2.58e-07 $l=7.45e-07 $layer=LI1_cond $X=3.25 $Y=1.295
+ $X2=3.25 $Y2=2.04
r114 23 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=0.35
+ $X2=3.505 $Y2=0.515
r115 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.505
+ $Y=0.35 $X2=3.505 $Y2=0.35
r116 20 22 24.46 $w=2.43e-07 $l=5.2e-07 $layer=LI1_cond $X=2.985 $Y=0.377
+ $X2=3.505 $Y2=0.377
r117 19 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=1.125
+ $X2=2.9 $Y2=1.21
r118 18 20 7.11011 $w=2.45e-07 $l=1.5995e-07 $layer=LI1_cond $X=2.9 $Y=0.5
+ $X2=2.985 $Y2=0.377
r119 18 19 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.9 $Y=0.5 $X2=2.9
+ $Y2=1.125
r120 17 36 2.80567 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.15 $Y=1.21
+ $X2=2.017 $Y2=1.21
r121 16 37 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=1.21
+ $X2=2.9 $Y2=1.21
r122 16 17 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.815 $Y=1.21
+ $X2=2.15 $Y2=1.21
r123 14 36 4.36371 $w=2.42e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.037 $Y=1.295
+ $X2=2.017 $Y2=1.21
r124 14 32 35.8538 $w=2.23e-07 $l=7e-07 $layer=LI1_cond $X=2.037 $Y=1.295
+ $X2=2.037 $Y2=1.995
r125 13 45 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.555 $Y=0.835
+ $X2=3.555 $Y2=0.515
r126 9 42 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.195 $Y=2.685
+ $X2=3.195 $Y2=2.205
r127 2 31 600 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.985 $X2=1.985 $Y2=2.15
r128 1 35 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.625 $X2=2.05 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%A_221_70# 1 2 8 9 10 11 13 14 15 17 20 23 25
+ 26 30 33 36 42 45 46 48 52 54 55
c130 45 0 1.48338e-19 $X=1.66 $Y=1.32
c131 36 0 1.07576e-19 $X=1.465 $Y=0.505
c132 13 0 1.93583e-19 $X=2.22 $Y=1.75
r133 50 52 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.41 $Y=2.465
+ $X2=1.55 $Y2=2.465
r134 48 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=2.3
+ $X2=1.55 $Y2=2.465
r135 48 55 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.55 $Y=2.3
+ $X2=1.55 $Y2=1.825
r136 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.66
+ $Y=1.32 $X2=1.66 $Y2=1.32
r137 43 55 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.61 $Y=1.68
+ $X2=1.61 $Y2=1.825
r138 43 45 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=1.61 $Y=1.68
+ $X2=1.61 $Y2=1.32
r139 42 54 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=1.61 $Y=1.3
+ $X2=1.61 $Y2=1.155
r140 42 45 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=1.61 $Y=1.3 $X2=1.61
+ $Y2=1.32
r141 40 54 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.55 $Y=0.67
+ $X2=1.55 $Y2=1.155
r142 36 40 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.465 $Y=0.505
+ $X2=1.55 $Y2=0.67
r143 36 38 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.465 $Y=0.505
+ $X2=1.245 $Y2=0.505
r144 34 46 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.66 $Y=1.675
+ $X2=1.66 $Y2=1.32
r145 32 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.66 $Y=1.305
+ $X2=1.66 $Y2=1.32
r146 32 33 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=1.66 $Y=1.305
+ $X2=1.66 $Y2=1.23
r147 28 30 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3.74 $Y=1.665
+ $X2=3.74 $Y2=2.575
r148 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.665 $Y=1.59
+ $X2=3.74 $Y2=1.665
r149 26 27 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.665 $Y=1.59
+ $X2=3.3 $Y2=1.59
r150 23 27 107.956 $w=2e-07 $l=5.43875e-07 $layer=POLY_cond $X=3.055 $Y=1.155
+ $X2=3.3 $Y2=1.59
r151 23 25 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.055 $Y=1.155
+ $X2=3.055 $Y2=0.835
r152 22 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.055 $Y=0.255
+ $X2=3.055 $Y2=0.835
r153 18 20 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.295 $Y=1.825
+ $X2=2.295 $Y2=2.685
r154 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.265 $Y=1.155
+ $X2=2.265 $Y2=0.835
r155 14 34 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.825 $Y=1.75
+ $X2=1.66 $Y2=1.675
r156 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.22 $Y=1.75
+ $X2=2.295 $Y2=1.825
r157 13 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.22 $Y=1.75
+ $X2=1.825 $Y2=1.75
r158 12 33 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.23
+ $X2=1.66 $Y2=1.23
r159 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.19 $Y=1.23
+ $X2=2.265 $Y2=1.155
r160 11 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.19 $Y=1.23
+ $X2=1.825 $Y2=1.23
r161 9 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.98 $Y=0.18
+ $X2=3.055 $Y2=0.255
r162 9 10 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=2.98 $Y=0.18
+ $X2=1.825 $Y2=0.18
r163 8 33 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.75 $Y=1.155
+ $X2=1.66 $Y2=1.23
r164 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.75 $Y=0.255
+ $X2=1.825 $Y2=0.18
r165 7 8 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.75 $Y=0.255 $X2=1.75
+ $Y2=1.155
r166 2 50 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.255
+ $Y=2.32 $X2=1.41 $Y2=2.465
r167 1 38 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.105
+ $Y=0.35 $X2=1.245 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%A_776_99# 1 2 7 9 14 18 22 26 30 34 36 40 43
+ 47 50 52 56 57 59 63 67 69 70 72
r134 74 76 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.805 $Y=1.46
+ $X2=6.235 $Y2=1.46
r135 63 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=2.025
+ $X2=4.19 $Y2=2.19
r136 63 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=2.025
+ $X2=4.19 $Y2=1.86
r137 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.19
+ $Y=2.025 $X2=4.19 $Y2=2.025
r138 59 62 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.19 $Y=1.805
+ $X2=4.19 $Y2=2.025
r139 57 76 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=6.45 $Y=1.46
+ $X2=6.235 $Y2=1.46
r140 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.46 $X2=6.45 $Y2=1.46
r141 54 56 36.494 $w=2.68e-07 $l=8.55e-07 $layer=LI1_cond $X=6.48 $Y=2.315
+ $X2=6.48 $Y2=1.46
r142 53 70 4.16724 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=5.54 $Y=2.4
+ $X2=5.282 $Y2=2.4
r143 52 54 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=6.345 $Y=2.4
+ $X2=6.48 $Y2=2.315
r144 52 53 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=6.345 $Y=2.4
+ $X2=5.54 $Y2=2.4
r145 48 70 2.64909 $w=3.62e-07 $l=1.898e-07 $layer=LI1_cond $X=5.13 $Y=2.485
+ $X2=5.282 $Y2=2.4
r146 48 50 22.4459 $w=2.08e-07 $l=4.25e-07 $layer=LI1_cond $X=5.13 $Y=2.485
+ $X2=5.13 $Y2=2.91
r147 45 70 2.64909 $w=3.62e-07 $l=8.5e-08 $layer=LI1_cond $X=5.282 $Y=2.315
+ $X2=5.282 $Y2=2.4
r148 45 47 7.78032 $w=5.13e-07 $l=3.35e-07 $layer=LI1_cond $X=5.282 $Y=2.315
+ $X2=5.282 $Y2=1.98
r149 44 69 2.79095 $w=3.42e-07 $l=1.07912e-07 $layer=LI1_cond $X=5.282 $Y=1.89
+ $X2=5.23 $Y2=1.805
r150 44 47 2.09023 $w=5.13e-07 $l=9e-08 $layer=LI1_cond $X=5.282 $Y=1.89
+ $X2=5.282 $Y2=1.98
r151 43 69 2.79095 $w=3.42e-07 $l=2.64102e-07 $layer=LI1_cond $X=5.005 $Y=1.72
+ $X2=5.23 $Y2=1.805
r152 42 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=1.195
+ $X2=5.005 $Y2=1.11
r153 42 43 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=5.005 $Y=1.195
+ $X2=5.005 $Y2=1.72
r154 38 67 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.65 $Y=1.11
+ $X2=5.005 $Y2=1.11
r155 38 40 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=4.65 $Y=1.025
+ $X2=4.65 $Y2=0.42
r156 37 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=1.805
+ $X2=4.19 $Y2=1.805
r157 36 69 3.95098 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=4.92 $Y=1.805
+ $X2=5.23 $Y2=1.805
r158 36 37 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.92 $Y=1.805
+ $X2=4.355 $Y2=1.805
r159 32 34 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=3.955 $Y=1.23
+ $X2=4.1 $Y2=1.23
r160 28 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.235 $Y=1.625
+ $X2=6.235 $Y2=1.46
r161 28 30 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.235 $Y=1.625
+ $X2=6.235 $Y2=2.465
r162 24 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.235 $Y=1.295
+ $X2=6.235 $Y2=1.46
r163 24 26 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=6.235 $Y=1.295
+ $X2=6.235 $Y2=0.655
r164 20 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.805 $Y=1.625
+ $X2=5.805 $Y2=1.46
r165 20 22 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.805 $Y=1.625
+ $X2=5.805 $Y2=2.465
r166 16 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.805 $Y=1.295
+ $X2=5.805 $Y2=1.46
r167 16 18 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.805 $Y=1.295
+ $X2=5.805 $Y2=0.655
r168 14 73 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=4.1 $Y=2.575
+ $X2=4.1 $Y2=2.19
r169 10 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.1 $Y=1.305
+ $X2=4.1 $Y2=1.23
r170 10 72 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.1 $Y=1.305
+ $X2=4.1 $Y2=1.86
r171 7 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.955 $Y=1.155
+ $X2=3.955 $Y2=1.23
r172 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.955 $Y=1.155
+ $X2=3.955 $Y2=0.835
r173 2 50 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.835 $X2=5.12 $Y2=2.91
r174 2 47 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.98
+ $Y=1.835 $X2=5.12 $Y2=1.98
r175 1 40 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=4.565
+ $Y=0.235 $X2=4.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%A_626_125# 1 2 9 13 15 16 17 22 27 31 32 34
r93 31 32 8.46329 $w=4.53e-07 $l=1.35e-07 $layer=LI1_cond $X=3.492 $Y=2.51
+ $X2=3.492 $Y2=2.375
r94 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=1.455 $X2=4.575 $Y2=1.455
r95 25 34 1.03991 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=1.457
+ $X2=3.635 $Y2=1.457
r96 25 27 51.258 $w=1.83e-07 $l=8.55e-07 $layer=LI1_cond $X=3.72 $Y=1.457
+ $X2=4.575 $Y2=1.457
r97 23 34 5.53942 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=3.635 $Y=1.55
+ $X2=3.635 $Y2=1.457
r98 23 32 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.635 $Y=1.55
+ $X2=3.635 $Y2=2.375
r99 22 34 5.53942 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=3.635 $Y=1.365
+ $X2=3.635 $Y2=1.457
r100 21 22 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.635 $Y=0.955
+ $X2=3.635 $Y2=1.365
r101 17 21 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=3.55 $Y=0.812
+ $X2=3.635 $Y2=0.955
r102 17 19 8.49168 $w=2.83e-07 $l=2.1e-07 $layer=LI1_cond $X=3.55 $Y=0.812
+ $X2=3.34 $Y2=0.812
r103 15 28 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=4.83 $Y=1.455
+ $X2=4.575 $Y2=1.455
r104 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.83 $Y=1.455
+ $X2=4.905 $Y2=1.455
r105 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=1.62
+ $X2=4.905 $Y2=1.455
r106 11 13 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=4.905 $Y=1.62
+ $X2=4.905 $Y2=2.465
r107 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=1.29
+ $X2=4.905 $Y2=1.455
r108 7 9 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=4.905 $Y=1.29
+ $X2=4.905 $Y2=0.655
r109 2 31 300 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=2 $X=3.27
+ $Y=2.365 $X2=3.43 $Y2=2.51
r110 1 19 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.625 $X2=3.34 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%RESET_B 3 6 8 10 11 18 21
c46 6 0 1.55618e-19 $X=5.335 $Y=2.465
r47 14 18 6.2424 $w=2.38e-07 $l=1.3e-07 $layer=LI1_cond $X=5.065 $Y=0.685
+ $X2=5.065 $Y2=0.555
r48 11 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.355 $Y=1.35
+ $X2=5.355 $Y2=1.515
r49 11 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.355 $Y=1.35
+ $X2=5.355 $Y2=1.185
r50 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.355
+ $Y=1.35 $X2=5.355 $Y2=1.35
r51 8 14 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.39 $Y=0.77
+ $X2=5.065 $Y2=0.77
r52 8 10 21.9407 $w=2.58e-07 $l=4.95e-07 $layer=LI1_cond $X=5.39 $Y=0.855
+ $X2=5.39 $Y2=1.35
r53 6 22 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.335 $Y=2.465
+ $X2=5.335 $Y2=1.515
r54 3 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.265 $Y=0.655
+ $X2=5.265 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%VPWR 1 2 3 4 5 18 22 27 30 34 36 38 41 43 45
+ 50 58 66 71 77 80 83 86 90
c103 30 0 1.55618e-19 $X=4.69 $Y=2.145
r104 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r105 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r106 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r107 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r108 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 75 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r110 75 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r111 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r112 72 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=3.33
+ $X2=5.57 $Y2=3.33
r113 72 74 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.735 $Y=3.33
+ $X2=6 $Y2=3.33
r114 71 89 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=6.285 $Y=3.33
+ $X2=6.502 $Y2=3.33
r115 71 74 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.285 $Y=3.33
+ $X2=6 $Y2=3.33
r116 70 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r117 70 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r118 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r119 67 83 13.7128 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.502 $Y2=3.33
r120 67 69 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=5.04 $Y2=3.33
r121 66 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.57 $Y2=3.33
r122 66 69 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r124 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 62 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r126 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r127 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r128 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=3.33
+ $X2=2.565 $Y2=3.33
r129 59 61 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.73 $Y=3.33
+ $X2=3.12 $Y2=3.33
r130 58 83 13.7128 $w=1.7e-07 $l=3.52e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=4.502 $Y2=3.33
r131 58 64 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.15 $Y=3.33 $X2=4.08
+ $Y2=3.33
r132 57 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r134 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r135 54 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r136 53 56 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r137 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 51 77 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.692 $Y2=3.33
r139 51 53 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 50 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.565 $Y2=3.33
r141 50 56 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r143 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r144 45 77 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.692 $Y2=3.33
r145 45 47 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.24 $Y2=3.33
r146 43 65 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r147 43 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r148 41 42 6.12241 $w=7.03e-07 $l=1.6e-07 $layer=LI1_cond $X=4.502 $Y=2.57
+ $X2=4.502 $Y2=2.41
r149 36 89 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=6.45 $Y=3.245
+ $X2=6.502 $Y2=3.33
r150 36 38 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.45 $Y=3.245
+ $X2=6.45 $Y2=2.78
r151 32 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=3.245
+ $X2=5.57 $Y2=3.33
r152 32 34 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.57 $Y=3.245
+ $X2=5.57 $Y2=2.78
r153 30 42 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.69 $Y=2.145
+ $X2=4.69 $Y2=2.41
r154 25 83 2.87722 $w=7.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.502 $Y=3.245
+ $X2=4.502 $Y2=3.33
r155 25 27 5.00487 $w=7.03e-07 $l=2.95e-07 $layer=LI1_cond $X=4.502 $Y=3.245
+ $X2=4.502 $Y2=2.95
r156 24 41 3.25741 $w=7.03e-07 $l=1.92e-07 $layer=LI1_cond $X=4.502 $Y=2.762
+ $X2=4.502 $Y2=2.57
r157 24 27 3.18954 $w=7.03e-07 $l=1.88e-07 $layer=LI1_cond $X=4.502 $Y=2.762
+ $X2=4.502 $Y2=2.95
r158 20 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=3.245
+ $X2=2.565 $Y2=3.33
r159 20 22 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.565 $Y=3.245
+ $X2=2.565 $Y2=2.88
r160 16 77 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=3.245
+ $X2=0.692 $Y2=3.33
r161 16 18 39.9514 $w=2.23e-07 $l=7.8e-07 $layer=LI1_cond $X=0.692 $Y=3.245
+ $X2=0.692 $Y2=2.465
r162 5 38 600 $w=1.7e-07 $l=1.01258e-06 $layer=licon1_PDIFF $count=1 $X=6.31
+ $Y=1.835 $X2=6.45 $Y2=2.78
r163 4 34 600 $w=1.7e-07 $l=1.02187e-06 $layer=licon1_PDIFF $count=1 $X=5.41
+ $Y=1.835 $X2=5.57 $Y2=2.78
r164 3 41 300 $w=1.7e-07 $l=6.08933e-07 $layer=licon1_PDIFF $count=2 $X=4.175
+ $Y=2.365 $X2=4.69 $Y2=2.57
r165 3 30 600 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=2.365 $X2=4.69 $Y2=2.145
r166 3 27 600 $w=1.7e-07 $l=8.02185e-07 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=2.365 $X2=4.69 $Y2=2.95
r167 2 22 600 $w=1.7e-07 $l=6.0469e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=2.365 $X2=2.565 $Y2=2.88
r168 1 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=2.32 $X2=0.71 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%Q 1 2 7 8 9 10 11 18
r19 10 11 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=6.01 $Y=1.665
+ $X2=6.01 $Y2=1.98
r20 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=6.01 $Y=1.295
+ $X2=6.01 $Y2=1.665
r21 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=6.01 $Y=0.925 $X2=6.01
+ $Y2=1.295
r22 7 8 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=6.01 $Y=0.555 $X2=6.01
+ $Y2=0.925
r23 7 18 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=6.01 $Y=0.555
+ $X2=6.01 $Y2=0.42
r24 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.88
+ $Y=1.835 $X2=6.02 $Y2=1.98
r25 1 18 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.88
+ $Y=0.235 $X2=6.02 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_2%VGND 1 2 3 4 5 20 24 26 30 34 36 38 40 42 50
+ 55 61 64 67 70 74
r96 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r97 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r98 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r99 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r100 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r101 59 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r102 59 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r103 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r104 56 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=0 $X2=5.52
+ $Y2=0
r105 56 58 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.685 $Y=0 $X2=6
+ $Y2=0
r106 55 73 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=6.285 $Y=0
+ $X2=6.502 $Y2=0
r107 55 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.285 $Y=0 $X2=6
+ $Y2=0
r108 54 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r109 54 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r110 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r111 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.17
+ $Y2=0
r112 51 53 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=5.04 $Y2=0
r113 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=0 $X2=5.52
+ $Y2=0
r114 50 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.355 $Y=0
+ $X2=5.04 $Y2=0
r115 49 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r116 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r117 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r118 46 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r119 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r120 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r121 43 61 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=0.82
+ $Y2=0
r122 43 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=1.2
+ $Y2=0
r123 42 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.48
+ $Y2=0
r124 42 48 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.16 $Y2=0
r125 40 68 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r126 40 65 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.64
+ $Y2=0
r127 36 73 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=6.45 $Y=0.085
+ $X2=6.502 $Y2=0
r128 36 38 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.45 $Y=0.085
+ $X2=6.45 $Y2=0.38
r129 32 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.52 $Y2=0
r130 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.52 $Y2=0.38
r131 28 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0
r132 28 30 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=4.17 $Y=0.085
+ $X2=4.17 $Y2=0.835
r133 27 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=0 $X2=2.48
+ $Y2=0
r134 26 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.17
+ $Y2=0
r135 26 27 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.005 $Y=0
+ $X2=2.645 $Y2=0
r136 22 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0
r137 22 24 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0.835
r138 18 61 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=0.085
+ $X2=0.82 $Y2=0
r139 18 20 20.1678 $w=2.38e-07 $l=4.2e-07 $layer=LI1_cond $X=0.82 $Y=0.085
+ $X2=0.82 $Y2=0.505
r140 5 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.31
+ $Y=0.235 $X2=6.45 $Y2=0.38
r141 4 34 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.235 $X2=5.52 $Y2=0.38
r142 3 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.625 $X2=4.17 $Y2=0.835
r143 2 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.34
+ $Y=0.625 $X2=2.48 $Y2=0.835
r144 1 20 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.675
+ $Y=0.35 $X2=0.815 $Y2=0.505
.ends

