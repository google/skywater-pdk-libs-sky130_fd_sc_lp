* File: sky130_fd_sc_lp__a31o_m.pex.spice
* Created: Fri Aug 28 09:59:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31O_M%A_86_172# 1 2 8 9 10 13 16 19 20 22 25 29 31
+ 34 36 37 38 40
c88 31 0 1.78365e-19 $X=3.05 $Y=0.945
r89 40 41 17.7696 $w=2.3e-07 $l=3.35e-07 $layer=LI1_cond $X=2.8 $Y=2.835
+ $X2=3.135 $Y2=2.835
r90 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.595
+ $Y=1.025 $X2=0.595 $Y2=1.025
r91 34 41 2.50919 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=2.67
+ $X2=3.135 $Y2=2.835
r92 33 34 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=3.135 $Y=1.03
+ $X2=3.135 $Y2=2.67
r93 32 38 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.375 $Y=0.945
+ $X2=2.27 $Y2=0.945
r94 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.05 $Y=0.945
+ $X2=3.135 $Y2=1.03
r95 31 32 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.05 $Y=0.945
+ $X2=2.375 $Y2=0.945
r96 27 38 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.27 $Y=0.86
+ $X2=2.27 $Y2=0.945
r97 27 29 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=2.27 $Y=0.86
+ $X2=2.27 $Y2=0.605
r98 26 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=0.945
+ $X2=0.595 $Y2=0.945
r99 25 38 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.165 $Y=0.945
+ $X2=2.27 $Y2=0.945
r100 25 26 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=2.165 $Y=0.945
+ $X2=0.68 $Y2=0.945
r101 21 37 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.595 $Y=1.365
+ $X2=0.595 $Y2=1.025
r102 21 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.365
+ $X2=0.595 $Y2=1.53
r103 20 37 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.595 $Y=1.01
+ $X2=0.595 $Y2=1.025
r104 19 20 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.67 $Y=0.86
+ $X2=0.67 $Y2=1.01
r105 14 16 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.865 $Y=2.31
+ $X2=0.865 $Y2=2.77
r106 13 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.835 $Y=0.54
+ $X2=0.835 $Y2=0.86
r107 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.79 $Y=2.235
+ $X2=0.865 $Y2=2.31
r108 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.79 $Y=2.235
+ $X2=0.58 $Y2=2.235
r109 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.505 $Y=2.16
+ $X2=0.58 $Y2=2.235
r110 8 22 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.505 $Y=2.16
+ $X2=0.505 $Y2=1.53
r111 2 40 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.66
+ $Y=2.56 $X2=2.8 $Y2=2.835
r112 1 29 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.13
+ $Y=0.33 $X2=2.27 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_M%A3 7 9 11 13 14 15 18 20 21 22 23 24 25 31
c62 22 0 1.4401e-19 $X=1.2 $Y=1.295
c63 21 0 1.24166e-19 $X=1.26 $Y=2.31
c64 13 0 1.40505e-19 $X=1.135 $Y=1.25
c65 7 0 1.42572e-19 $X=1.295 $Y=2.77
r66 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.135
+ $Y=1.415 $X2=1.135 $Y2=1.415
r67 24 25 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.167 $Y=2.035
+ $X2=1.167 $Y2=2.405
r68 23 24 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.167 $Y=1.665
+ $X2=1.167 $Y2=2.035
r69 23 32 12.26 $w=2.33e-07 $l=2.5e-07 $layer=LI1_cond $X=1.167 $Y=1.665
+ $X2=1.167 $Y2=1.415
r70 22 32 5.88482 $w=2.33e-07 $l=1.2e-07 $layer=LI1_cond $X=1.167 $Y=1.295
+ $X2=1.167 $Y2=1.415
r71 20 21 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.26 $Y=2.16
+ $X2=1.26 $Y2=2.31
r72 16 18 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.195 $Y=0.935
+ $X2=1.335 $Y2=0.935
r73 15 20 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.225 $Y=1.92
+ $X2=1.225 $Y2=2.16
r74 14 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.135 $Y=1.755
+ $X2=1.135 $Y2=1.415
r75 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.755
+ $X2=1.135 $Y2=1.92
r76 13 31 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=1.25
+ $X2=1.135 $Y2=1.415
r77 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=0.86
+ $X2=1.335 $Y2=0.935
r78 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.335 $Y=0.86
+ $X2=1.335 $Y2=0.54
r79 7 21 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.295 $Y=2.77
+ $X2=1.295 $Y2=2.31
r80 1 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.195 $Y=1.01
+ $X2=1.195 $Y2=0.935
r81 1 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.195 $Y=1.01
+ $X2=1.195 $Y2=1.25
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_M%A2 3 7 11 12 13 14 15 20
c47 13 0 1.40505e-19 $X=1.68 $Y=1.295
c48 3 0 2.70616e-19 $X=1.695 $Y=0.54
r49 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.675
+ $Y=1.415 $X2=1.675 $Y2=1.415
r50 14 15 23.4494 $w=1.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.677 $Y=1.665
+ $X2=1.677 $Y2=2.035
r51 14 21 15.8442 $w=1.73e-07 $l=2.5e-07 $layer=LI1_cond $X=1.677 $Y=1.665
+ $X2=1.677 $Y2=1.415
r52 13 21 7.60519 $w=1.73e-07 $l=1.2e-07 $layer=LI1_cond $X=1.677 $Y=1.295
+ $X2=1.677 $Y2=1.415
r53 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.675 $Y=1.755
+ $X2=1.675 $Y2=1.415
r54 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.755
+ $X2=1.675 $Y2=1.92
r55 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.25
+ $X2=1.675 $Y2=1.415
r56 7 12 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.725 $Y=2.77
+ $X2=1.725 $Y2=1.92
r57 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.695 $Y=0.54
+ $X2=1.695 $Y2=1.25
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_M%A1 3 8 10 11 13 14 15 16 17 18 23
c53 23 0 1.78365e-19 $X=2.215 $Y=1.415
c54 16 0 1.26606e-19 $X=2.16 $Y=1.295
c55 13 0 1.32474e-19 $X=2.215 $Y=1.25
r56 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.215
+ $Y=1.415 $X2=2.215 $Y2=1.415
r57 17 18 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.187 $Y=1.665
+ $X2=2.187 $Y2=2.035
r58 17 24 12.8049 $w=2.23e-07 $l=2.5e-07 $layer=LI1_cond $X=2.187 $Y=1.665
+ $X2=2.187 $Y2=1.415
r59 16 24 6.14636 $w=2.23e-07 $l=1.2e-07 $layer=LI1_cond $X=2.187 $Y=1.295
+ $X2=2.187 $Y2=1.415
r60 14 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.215 $Y=1.755
+ $X2=2.215 $Y2=1.415
r61 14 15 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.755
+ $X2=2.215 $Y2=1.92
r62 13 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.25
+ $X2=2.215 $Y2=1.415
r63 11 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.125 $Y=1.01
+ $X2=2.125 $Y2=1.25
r64 10 11 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.09 $Y=0.86
+ $X2=2.09 $Y2=1.01
r65 8 15 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=2.155 $Y=2.77
+ $X2=2.155 $Y2=1.92
r66 3 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.055 $Y=0.54
+ $X2=2.055 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_M%B1 1 3 6 12 15 16 18 19 20 21 22 28
c47 19 0 1.32474e-19 $X=2.64 $Y=1.295
r48 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.785
+ $Y=1.805 $X2=2.785 $Y2=1.805
r49 21 22 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.712 $Y=2.035
+ $X2=2.712 $Y2=2.405
r50 21 29 8.41466 $w=3.13e-07 $l=2.3e-07 $layer=LI1_cond $X=2.712 $Y=2.035
+ $X2=2.712 $Y2=1.805
r51 20 29 5.12197 $w=3.13e-07 $l=1.4e-07 $layer=LI1_cond $X=2.712 $Y=1.665
+ $X2=2.712 $Y2=1.805
r52 19 20 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.712 $Y=1.295
+ $X2=2.712 $Y2=1.665
r53 18 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.64
+ $X2=2.785 $Y2=1.805
r54 15 28 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.785 $Y=2.16
+ $X2=2.785 $Y2=1.805
r55 15 16 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.73 $Y=2.16
+ $X2=2.73 $Y2=2.31
r56 10 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.485 $Y=0.935
+ $X2=2.695 $Y2=0.935
r57 8 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.695 $Y=1.01
+ $X2=2.695 $Y2=0.935
r58 8 18 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.695 $Y=1.01
+ $X2=2.695 $Y2=1.64
r59 6 16 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.585 $Y=2.77
+ $X2=2.585 $Y2=2.31
r60 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.485 $Y=0.86
+ $X2=2.485 $Y2=0.935
r61 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.485 $Y=0.86
+ $X2=2.485 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_M%X 1 2 7 8 11 17 20
c28 11 0 1.24166e-19 $X=0.65 $Y=2.705
r29 19 20 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.24 $Y=1.71
+ $X2=0.24 $Y2=0.925
r30 14 20 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.24 $Y=0.68
+ $X2=0.24 $Y2=0.925
r31 13 17 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.24 $Y=0.515
+ $X2=0.62 $Y2=0.515
r32 13 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.515
+ $X2=0.24 $Y2=0.68
r33 9 11 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=0.64 $Y=1.88
+ $X2=0.64 $Y2=2.705
r34 8 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.325 $Y=1.795
+ $X2=0.24 $Y2=1.71
r35 7 9 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.545 $Y=1.795
+ $X2=0.64 $Y2=1.88
r36 7 8 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.545 $Y=1.795
+ $X2=0.325 $Y2=1.795
r37 2 11 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.525
+ $Y=2.56 $X2=0.65 $Y2=2.705
r38 1 17 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.495
+ $Y=0.33 $X2=0.62 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_M%VPWR 1 2 9 13 16 17 19 20 21 34 35
r40 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r43 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 21 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 19 28 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 19 20 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.93 $Y2=3.33
r50 18 31 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 18 20 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.93 $Y2=3.33
r52 16 24 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=1.08 $Y2=3.33
r54 15 28 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=1.08 $Y2=3.33
r56 11 20 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=3.33
r57 11 13 23.933 $w=1.88e-07 $l=4.1e-07 $layer=LI1_cond $X=1.93 $Y=3.245
+ $X2=1.93 $Y2=2.835
r58 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=3.245 $X2=1.08
+ $Y2=3.33
r59 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.08 $Y=3.245 $X2=1.08
+ $Y2=2.835
r60 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.8
+ $Y=2.56 $X2=1.94 $Y2=2.835
r61 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.94
+ $Y=2.56 $X2=1.08 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_M%A_274_512# 1 2 9 10 12 14 15 20
c33 14 0 1.42572e-19 $X=1.51 $Y=2.835
r34 17 20 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=2.29 $Y=2.775 $X2=2.37
+ $Y2=2.775
r35 14 15 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.53 $Y=2.835
+ $X2=1.53 $Y2=2.67
r36 12 17 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.29 $Y=2.67 $X2=2.29
+ $Y2=2.775
r37 11 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.29 $Y=2.49
+ $X2=2.29 $Y2=2.67
r38 9 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.205 $Y=2.405
+ $X2=2.29 $Y2=2.49
r39 9 10 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.205 $Y=2.405
+ $X2=1.635 $Y2=2.405
r40 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.55 $Y=2.49
+ $X2=1.635 $Y2=2.405
r41 7 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.55 $Y=2.49 $X2=1.55
+ $Y2=2.67
r42 2 20 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=2.23
+ $Y=2.56 $X2=2.37 $Y2=2.775
r43 1 14 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.37
+ $Y=2.56 $X2=1.51 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_M%VGND 1 2 9 11 15 17 19 26 27 30 33
r35 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r36 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r37 27 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r38 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 24 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=2.7
+ $Y2=0
r40 24 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.805 $Y=0 $X2=3.12
+ $Y2=0
r41 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r42 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r44 19 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r45 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r46 17 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r47 13 33 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=0.085 $X2=2.7
+ $Y2=0
r48 13 15 20.5974 $w=2.08e-07 $l=3.9e-07 $layer=LI1_cond $X=2.7 $Y=0.085 $X2=2.7
+ $Y2=0.475
r49 12 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r50 11 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.7
+ $Y2=0
r51 11 12 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.595 $Y=0
+ $X2=1.235 $Y2=0
r52 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r53 7 9 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0.475
r54 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.56
+ $Y=0.33 $X2=2.7 $Y2=0.475
r55 1 9 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.33 $X2=1.07 $Y2=0.475
.ends

