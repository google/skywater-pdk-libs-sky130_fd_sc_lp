* File: sky130_fd_sc_lp__nand3_m.pex.spice
* Created: Fri Aug 28 10:49:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3_M%C 2 5 9 13 15 18 20 21 22 23 29
r36 22 23 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r37 21 22 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r38 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.295
r39 20 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r40 16 18 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=0.36 $Y=1.845
+ $X2=0.5 $Y2=1.845
r41 14 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.005
r42 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.51
r43 13 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.99
+ $X2=0.27 $Y2=1.005
r44 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.345 $Y=0.84
+ $X2=0.345 $Y2=0.99
r45 9 12 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.51 $Y=0.445
+ $X2=0.51 $Y2=0.84
r46 3 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.5 $Y=1.92 $X2=0.5
+ $Y2=1.845
r47 3 5 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.5 $Y=1.92 $X2=0.5
+ $Y2=2.52
r48 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=1.77 $X2=0.36
+ $Y2=1.845
r49 2 15 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=0.36 $Y=1.77 $X2=0.36
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_M%B 3 7 9 10 11 16
c38 16 0 1.44794e-19 $X=0.84 $Y=1.365
r39 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.365
+ $X2=0.84 $Y2=1.53
r40 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.365
+ $X2=0.84 $Y2=1.2
r41 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.84
+ $Y=1.365 $X2=0.84 $Y2=1.365
r42 11 17 11.9218 $w=2.88e-07 $l=3e-07 $layer=LI1_cond $X=0.78 $Y=1.665 $X2=0.78
+ $Y2=1.365
r43 10 17 2.78176 $w=2.88e-07 $l=7e-08 $layer=LI1_cond $X=0.78 $Y=1.295 $X2=0.78
+ $Y2=1.365
r44 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.78 $Y=0.925
+ $X2=0.78 $Y2=1.295
r45 7 19 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=0.93 $Y=2.52 $X2=0.93
+ $Y2=1.53
r46 3 18 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.9 $Y=0.445 $X2=0.9
+ $Y2=1.2
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_M%A 3 7 11 12 13 14 15 20
r34 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.38
+ $Y=1.005 $X2=1.38 $Y2=1.005
r35 14 15 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.29 $Y=1.295
+ $X2=1.29 $Y2=1.665
r36 14 21 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=1.29 $Y=1.295
+ $X2=1.29 $Y2=1.005
r37 13 21 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=1.29 $Y=0.925 $X2=1.29
+ $Y2=1.005
r38 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.38 $Y=1.345
+ $X2=1.38 $Y2=1.005
r39 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.345
+ $X2=1.38 $Y2=1.51
r40 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=0.84
+ $X2=1.38 $Y2=1.005
r41 7 12 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.36 $Y=2.52
+ $X2=1.36 $Y2=1.51
r42 3 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.29 $Y=0.445
+ $X2=1.29 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_M%VPWR 1 2 7 9 13 16 17 18 25 26
r27 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 23 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 20 29 3.64449 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r32 20 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 18 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 18 23 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 16 22 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=3.33 $X2=0.72
+ $Y2=3.33
r36 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=1.145 $Y2=3.33
r37 15 25 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.145 $Y2=3.33
r39 11 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=3.33
r40 11 13 37.4978 $w=2.08e-07 $l=7.1e-07 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=2.535
r41 7 29 3.2707 $w=2.1e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.195 $Y2=3.33
r42 7 9 37.4978 $w=2.08e-07 $l=7.1e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.285 $Y2=2.535
r43 2 13 600 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=2.31 $X2=1.145 $Y2=2.535
r44 1 9 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.31 $X2=0.285 $Y2=2.535
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_M%Y 1 2 3 10 15 16 17 24 30 35
c39 24 0 1.44794e-19 $X=1.47 $Y=2.035
r40 17 24 2.87242 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.642 $Y=2.035
+ $X2=1.47 $Y2=2.035
r41 17 35 10.7135 $w=5.13e-07 $l=4.05e-07 $layer=LI1_cond $X=1.642 $Y=2.12
+ $X2=1.642 $Y2=2.525
r42 16 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.2 $Y=2.035 $X2=1.47
+ $Y2=2.035
r43 16 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=0.82 $Y2=2.035
r44 15 25 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.715 $Y=2.035
+ $X2=0.82 $Y2=2.035
r45 15 30 14.5716 $w=3.78e-07 $l=4.05e-07 $layer=LI1_cond $X=0.715 $Y=2.12
+ $X2=0.715 $Y2=2.525
r46 14 17 54.288 $w=2.88e-07 $l=1.335e-06 $layer=LI1_cond $X=1.73 $Y=0.615
+ $X2=1.73 $Y2=1.95
r47 10 14 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.645 $Y=0.51
+ $X2=1.73 $Y2=0.615
r48 10 12 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=1.645 $Y=0.51
+ $X2=1.505 $Y2=0.51
r49 3 35 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=2.31 $X2=1.575 $Y2=2.525
r50 2 30 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=2.31 $X2=0.715 $Y2=2.525
r51 1 12 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.365
+ $Y=0.235 $X2=1.505 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_M%VGND 1 4 6 8 15 16
r23 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r24 15 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r25 13 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r26 12 15 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r27 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r28 10 19 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.23
+ $Y2=0
r29 10 12 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.72
+ $Y2=0
r30 8 16 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r31 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r32 4 19 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.23 $Y2=0
r33 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.38
r34 1 6 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.235 $X2=0.295 $Y2=0.38
.ends

