* File: sky130_fd_sc_lp__nand4b_m.pxi.spice
* Created: Wed Sep  2 10:06:31 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4B_M%A_N N_A_N_M1005_g N_A_N_M1003_g N_A_N_c_68_n
+ N_A_N_c_69_n A_N A_N A_N A_N A_N N_A_N_c_71_n PM_SKY130_FD_SC_LP__NAND4B_M%A_N
x_PM_SKY130_FD_SC_LP__NAND4B_M%D N_D_M1008_g N_D_M1004_g N_D_c_108_n N_D_c_109_n
+ N_D_c_110_n N_D_c_111_n N_D_c_115_n D D D N_D_c_113_n
+ PM_SKY130_FD_SC_LP__NAND4B_M%D
x_PM_SKY130_FD_SC_LP__NAND4B_M%C N_C_M1009_g N_C_M1000_g N_C_c_157_n N_C_c_158_n
+ N_C_c_159_n C C C N_C_c_161_n PM_SKY130_FD_SC_LP__NAND4B_M%C
x_PM_SKY130_FD_SC_LP__NAND4B_M%B N_B_M1006_g N_B_M1001_g N_B_c_198_n N_B_c_205_n
+ N_B_c_199_n N_B_c_200_n N_B_c_201_n B B B N_B_c_203_n
+ PM_SKY130_FD_SC_LP__NAND4B_M%B
x_PM_SKY130_FD_SC_LP__NAND4B_M%A_35_392# N_A_35_392#_M1003_s N_A_35_392#_M1005_s
+ N_A_35_392#_c_245_n N_A_35_392#_M1002_g N_A_35_392#_M1007_g
+ N_A_35_392#_c_248_n N_A_35_392#_c_243_n N_A_35_392#_c_244_n
+ N_A_35_392#_c_250_n N_A_35_392#_c_251_n PM_SKY130_FD_SC_LP__NAND4B_M%A_35_392#
x_PM_SKY130_FD_SC_LP__NAND4B_M%VPWR N_VPWR_M1005_d N_VPWR_M1000_d N_VPWR_M1002_d
+ N_VPWR_c_298_n N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n
+ N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_306_n VPWR
+ N_VPWR_c_307_n N_VPWR_c_297_n PM_SKY130_FD_SC_LP__NAND4B_M%VPWR
x_PM_SKY130_FD_SC_LP__NAND4B_M%Y N_Y_M1007_d N_Y_M1004_d N_Y_M1006_d N_Y_c_333_n
+ Y Y Y Y N_Y_c_337_n Y Y N_Y_c_343_n N_Y_c_356_n PM_SKY130_FD_SC_LP__NAND4B_M%Y
x_PM_SKY130_FD_SC_LP__NAND4B_M%VGND N_VGND_M1003_d N_VGND_c_382_n VGND
+ N_VGND_c_383_n N_VGND_c_384_n N_VGND_c_385_n PM_SKY130_FD_SC_LP__NAND4B_M%VGND
cc_1 VNB N_A_N_M1005_g 0.00859671f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.17
cc_2 VNB N_A_N_M1003_g 0.0250152f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.47
cc_3 VNB N_A_N_c_68_n 0.0265001f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.36
cc_4 VNB N_A_N_c_69_n 0.0207068f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.51
cc_5 VNB A_N 0.00397518f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_A_N_c_71_n 0.0187305f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.005
cc_7 VNB N_D_c_108_n 0.0175775f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.36
cc_8 VNB N_D_c_109_n 0.0230616f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.36
cc_9 VNB N_D_c_110_n 0.0167307f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.51
cc_10 VNB N_D_c_111_n 0.0112453f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_11 VNB D 0.00125221f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_12 VNB N_D_c_113_n 0.0167415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C_M1000_g 0.00995715f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.47
cc_14 VNB N_C_c_157_n 0.0163949f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.012
cc_15 VNB N_C_c_158_n 0.0230536f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.36
cc_16 VNB N_C_c_159_n 0.0158492f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.36
cc_17 VNB C 6.93262e-19 $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.51
cc_18 VNB N_C_c_161_n 0.0163629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B_c_198_n 0.0106802f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.012
cc_20 VNB N_B_c_199_n 0.0174079f $X=-0.19 $Y=-0.245 $X2=0.627 $Y2=1.51
cc_21 VNB N_B_c_200_n 0.0209292f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_22 VNB N_B_c_201_n 0.015299f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_23 VNB B 0.00570518f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_24 VNB N_B_c_203_n 0.0153262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_35_392#_M1007_g 0.070228f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_26 VNB N_A_35_392#_c_243_n 0.0497479f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.005
cc_27 VNB N_A_35_392#_c_244_n 0.00851174f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=0.84
cc_28 VNB N_VPWR_c_297_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_333_n 0.0109413f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_30 VNB Y 0.0101834f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_31 VNB Y 0.00472097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB Y 0.0633392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_337_n 0.00714201f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.665
cc_34 VNB N_VGND_c_382_n 0.00544905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_383_n 0.0729881f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_36 VNB N_VGND_c_384_n 0.236026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_385_n 0.0246766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_N_M1005_g 0.0297459f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.17
cc_39 VPB A_N 0.00564998f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_40 VPB N_D_c_111_n 0.00228753f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_41 VPB N_D_c_115_n 0.0270591f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_42 VPB N_C_M1000_g 0.0248656f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.47
cc_43 VPB N_B_c_198_n 0.00210941f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.012
cc_44 VPB N_B_c_205_n 0.0251677f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.36
cc_45 VPB N_A_35_392#_c_245_n 0.124654f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.47
cc_46 VPB N_A_35_392#_M1002_g 0.0409646f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.51
cc_47 VPB N_A_35_392#_M1007_g 0.00272119f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_48 VPB N_A_35_392#_c_248_n 0.0225618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_35_392#_c_243_n 0.0495943f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.005
cc_50 VPB N_A_35_392#_c_250_n 0.0226765f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.665
cc_51 VPB N_A_35_392#_c_251_n 0.0433123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_298_n 0.0286202f $X=-0.19 $Y=1.655 $X2=0.627 $Y2=1.51
cc_53 VPB N_VPWR_c_299_n 0.0293529f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_54 VPB N_VPWR_c_300_n 0.0420147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_301_n 0.0277576f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.005
cc_56 VPB N_VPWR_c_302_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.005
cc_57 VPB N_VPWR_c_303_n 0.0218935f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=0.84
cc_58 VPB N_VPWR_c_304_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.925
cc_59 VPB N_VPWR_c_305_n 0.0218935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_306_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.295
cc_61 VPB N_VPWR_c_307_n 0.0169405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_297_n 0.0947645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB Y 0.00308243f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_64 VPB Y 0.017566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_Y_c_337_n 0.00581829f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.665
cc_66 N_A_N_M1003_g N_D_c_108_n 0.00746253f $X=0.545 $Y=0.47 $X2=0 $Y2=0
cc_67 N_A_N_c_68_n N_D_c_109_n 0.0128127f $X=0.627 $Y=1.36 $X2=0 $Y2=0
cc_68 N_A_N_c_69_n N_D_c_110_n 0.0128127f $X=0.627 $Y=1.51 $X2=0 $Y2=0
cc_69 N_A_N_M1005_g N_D_c_111_n 0.00434583f $X=0.515 $Y=2.17 $X2=0 $Y2=0
cc_70 N_A_N_c_69_n N_D_c_111_n 0.00170624f $X=0.627 $Y=1.51 $X2=0 $Y2=0
cc_71 A_N N_D_c_111_n 0.00222172f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_72 N_A_N_M1005_g N_D_c_115_n 0.00600442f $X=0.515 $Y=2.17 $X2=0 $Y2=0
cc_73 A_N N_D_c_115_n 0.00328117f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_74 N_A_N_M1003_g D 0.00226132f $X=0.545 $Y=0.47 $X2=0 $Y2=0
cc_75 A_N D 0.0320704f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_76 N_A_N_c_71_n D 0.00190534f $X=0.65 $Y=1.005 $X2=0 $Y2=0
cc_77 N_A_N_M1003_g N_D_c_113_n 0.00137394f $X=0.545 $Y=0.47 $X2=0 $Y2=0
cc_78 A_N N_D_c_113_n 0.00240821f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_79 N_A_N_c_71_n N_D_c_113_n 0.0128127f $X=0.65 $Y=1.005 $X2=0 $Y2=0
cc_80 N_A_N_M1003_g N_A_35_392#_c_243_n 0.0177745f $X=0.545 $Y=0.47 $X2=0 $Y2=0
cc_81 N_A_N_c_69_n N_A_35_392#_c_243_n 0.0185364f $X=0.627 $Y=1.51 $X2=0 $Y2=0
cc_82 A_N N_A_35_392#_c_243_n 0.102366f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_83 N_A_N_M1003_g N_A_35_392#_c_244_n 0.00429189f $X=0.545 $Y=0.47 $X2=0 $Y2=0
cc_84 N_A_N_M1005_g N_A_35_392#_c_250_n 0.00506965f $X=0.515 $Y=2.17 $X2=0 $Y2=0
cc_85 A_N N_A_35_392#_c_250_n 0.0149489f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_86 N_A_N_M1005_g N_A_35_392#_c_251_n 0.00234487f $X=0.515 $Y=2.17 $X2=0 $Y2=0
cc_87 A_N N_A_35_392#_c_251_n 0.0049095f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_88 A_N N_VPWR_M1005_d 0.0053976f $X=0.635 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_89 N_A_N_M1005_g N_VPWR_c_298_n 0.00120183f $X=0.515 $Y=2.17 $X2=0 $Y2=0
cc_90 A_N N_VPWR_c_298_n 0.030321f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_91 N_A_N_M1005_g Y 5.85846e-19 $X=0.515 $Y=2.17 $X2=0 $Y2=0
cc_92 A_N Y 0.00967627f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_93 A_N N_Y_c_343_n 0.0102913f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_94 N_A_N_M1003_g N_VGND_c_382_n 0.00307951f $X=0.545 $Y=0.47 $X2=0 $Y2=0
cc_95 A_N N_VGND_c_382_n 0.00721374f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_96 N_A_N_c_71_n N_VGND_c_382_n 0.00140441f $X=0.65 $Y=1.005 $X2=0 $Y2=0
cc_97 N_A_N_M1003_g N_VGND_c_384_n 0.00952361f $X=0.545 $Y=0.47 $X2=0 $Y2=0
cc_98 A_N N_VGND_c_384_n 0.00422616f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_99 N_A_N_M1003_g N_VGND_c_385_n 0.00530222f $X=0.545 $Y=0.47 $X2=0 $Y2=0
cc_100 N_D_c_111_n N_C_M1000_g 0.0112097f $X=1.282 $Y=1.7 $X2=0 $Y2=0
cc_101 N_D_c_115_n N_C_M1000_g 0.0204913f $X=1.282 $Y=1.85 $X2=0 $Y2=0
cc_102 N_D_c_108_n N_C_c_157_n 0.0204582f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_103 D N_C_c_157_n 0.00300949f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_104 N_D_c_109_n N_C_c_158_n 0.0204582f $X=1.19 $Y=1.295 $X2=0 $Y2=0
cc_105 N_D_c_110_n N_C_c_159_n 0.0204582f $X=1.19 $Y=1.46 $X2=0 $Y2=0
cc_106 N_D_c_108_n C 0.00300949f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_107 D C 0.0574798f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_108 N_D_c_113_n N_C_c_161_n 0.0204582f $X=1.19 $Y=0.955 $X2=0 $Y2=0
cc_109 N_D_c_115_n N_A_35_392#_c_245_n 0.00582844f $X=1.282 $Y=1.85 $X2=0 $Y2=0
cc_110 D N_A_35_392#_c_243_n 0.00600246f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_111 D N_A_35_392#_c_244_n 0.00224109f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_112 N_D_c_110_n N_VPWR_c_298_n 0.00283068f $X=1.19 $Y=1.46 $X2=0 $Y2=0
cc_113 N_D_c_115_n N_VPWR_c_298_n 0.00358825f $X=1.282 $Y=1.85 $X2=0 $Y2=0
cc_114 N_D_c_110_n Y 0.00251364f $X=1.19 $Y=1.46 $X2=0 $Y2=0
cc_115 N_D_c_111_n Y 0.00667194f $X=1.282 $Y=1.7 $X2=0 $Y2=0
cc_116 N_D_c_115_n Y 0.00769865f $X=1.282 $Y=1.85 $X2=0 $Y2=0
cc_117 D Y 0.01652f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_118 N_D_c_115_n N_Y_c_343_n 0.0106992f $X=1.282 $Y=1.85 $X2=0 $Y2=0
cc_119 D N_VGND_M1003_d 0.00447568f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_120 N_D_c_108_n N_VGND_c_382_n 0.00592481f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_121 D N_VGND_c_382_n 0.00732421f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_122 N_D_c_108_n N_VGND_c_383_n 0.00380846f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_123 D N_VGND_c_383_n 0.00849572f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_124 N_D_c_108_n N_VGND_c_384_n 0.00576022f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_125 D N_VGND_c_384_n 0.0104566f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_126 N_C_M1000_g N_B_c_198_n 0.0100634f $X=1.715 $Y=2.17 $X2=0 $Y2=0
cc_127 N_C_M1000_g N_B_c_205_n 0.018573f $X=1.715 $Y=2.17 $X2=0 $Y2=0
cc_128 N_C_c_157_n N_B_c_199_n 0.0216015f $X=1.73 $Y=0.79 $X2=0 $Y2=0
cc_129 C N_B_c_199_n 0.00115329f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_130 N_C_c_158_n N_B_c_200_n 0.0142529f $X=1.73 $Y=1.295 $X2=0 $Y2=0
cc_131 N_C_c_159_n N_B_c_201_n 0.0142529f $X=1.73 $Y=1.46 $X2=0 $Y2=0
cc_132 N_C_c_157_n B 4.29236e-19 $X=1.73 $Y=0.79 $X2=0 $Y2=0
cc_133 C B 0.0618559f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_134 N_C_c_161_n B 0.00336481f $X=1.73 $Y=0.955 $X2=0 $Y2=0
cc_135 C N_B_c_203_n 6.94997e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 N_C_c_161_n N_B_c_203_n 0.0142529f $X=1.73 $Y=0.955 $X2=0 $Y2=0
cc_137 N_C_M1000_g N_A_35_392#_c_245_n 0.00582844f $X=1.715 $Y=2.17 $X2=0 $Y2=0
cc_138 N_C_M1000_g N_VPWR_c_299_n 0.00308284f $X=1.715 $Y=2.17 $X2=0 $Y2=0
cc_139 N_C_M1000_g Y 0.00278125f $X=1.715 $Y=2.17 $X2=0 $Y2=0
cc_140 N_C_c_159_n Y 0.00222012f $X=1.73 $Y=1.46 $X2=0 $Y2=0
cc_141 C Y 0.0076422f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_142 N_C_M1000_g N_Y_c_337_n 0.0113891f $X=1.715 $Y=2.17 $X2=0 $Y2=0
cc_143 N_C_c_159_n N_Y_c_337_n 0.00294516f $X=1.73 $Y=1.46 $X2=0 $Y2=0
cc_144 C N_Y_c_337_n 0.015671f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_145 N_C_M1000_g N_Y_c_343_n 0.00998842f $X=1.715 $Y=2.17 $X2=0 $Y2=0
cc_146 N_C_M1000_g N_Y_c_356_n 9.1742e-19 $X=1.715 $Y=2.17 $X2=0 $Y2=0
cc_147 N_C_c_157_n N_VGND_c_383_n 0.00380846f $X=1.73 $Y=0.79 $X2=0 $Y2=0
cc_148 C N_VGND_c_383_n 0.00849572f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_149 N_C_c_157_n N_VGND_c_384_n 0.00547146f $X=1.73 $Y=0.79 $X2=0 $Y2=0
cc_150 C N_VGND_c_384_n 0.0104566f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_151 C A_343_52# 0.0036372f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_152 N_B_c_205_n N_A_35_392#_c_245_n 0.00582844f $X=2.162 $Y=1.85 $X2=0 $Y2=0
cc_153 N_B_c_205_n N_A_35_392#_M1002_g 0.013709f $X=2.162 $Y=1.85 $X2=0 $Y2=0
cc_154 N_B_c_198_n N_A_35_392#_M1007_g 0.00792027f $X=2.162 $Y=1.7 $X2=0 $Y2=0
cc_155 N_B_c_199_n N_A_35_392#_M1007_g 0.0204501f $X=2.27 $Y=0.79 $X2=0 $Y2=0
cc_156 B N_A_35_392#_M1007_g 0.00550012f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_157 N_B_c_203_n N_A_35_392#_M1007_g 0.0416548f $X=2.27 $Y=0.955 $X2=0 $Y2=0
cc_158 N_B_c_205_n N_A_35_392#_c_248_n 0.00802233f $X=2.162 $Y=1.85 $X2=0 $Y2=0
cc_159 N_B_c_205_n N_VPWR_c_299_n 0.00308284f $X=2.162 $Y=1.85 $X2=0 $Y2=0
cc_160 N_B_c_199_n N_Y_c_333_n 3.26047e-19 $X=2.27 $Y=0.79 $X2=0 $Y2=0
cc_161 B N_Y_c_333_n 0.00803123f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_162 N_B_c_198_n Y 0.003388f $X=2.162 $Y=1.7 $X2=0 $Y2=0
cc_163 N_B_c_205_n Y 8.02895e-19 $X=2.162 $Y=1.85 $X2=0 $Y2=0
cc_164 N_B_c_201_n Y 0.00522402f $X=2.27 $Y=1.46 $X2=0 $Y2=0
cc_165 B Y 0.0184503f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_166 B Y 0.0218223f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_167 N_B_c_198_n N_Y_c_337_n 0.00382735f $X=2.162 $Y=1.7 $X2=0 $Y2=0
cc_168 N_B_c_205_n N_Y_c_337_n 0.00721397f $X=2.162 $Y=1.85 $X2=0 $Y2=0
cc_169 B N_Y_c_337_n 0.00816878f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_170 N_B_c_205_n N_Y_c_343_n 9.2663e-19 $X=2.162 $Y=1.85 $X2=0 $Y2=0
cc_171 N_B_c_205_n N_Y_c_356_n 0.0108955f $X=2.162 $Y=1.85 $X2=0 $Y2=0
cc_172 N_B_c_199_n N_VGND_c_383_n 0.00379643f $X=2.27 $Y=0.79 $X2=0 $Y2=0
cc_173 B N_VGND_c_383_n 0.00897195f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_174 N_B_c_199_n N_VGND_c_384_n 0.00585672f $X=2.27 $Y=0.79 $X2=0 $Y2=0
cc_175 B N_VGND_c_384_n 0.0114764f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_176 B A_451_52# 0.00431126f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_177 N_A_35_392#_c_245_n N_VPWR_c_298_n 0.0186861f $X=2.5 $Y=2.975 $X2=0 $Y2=0
cc_178 N_A_35_392#_c_243_n N_VPWR_c_298_n 0.00734437f $X=0.3 $Y=2.105 $X2=0
+ $Y2=0
cc_179 N_A_35_392#_c_250_n N_VPWR_c_298_n 0.0244122f $X=0.72 $Y=2.885 $X2=0
+ $Y2=0
cc_180 N_A_35_392#_c_251_n N_VPWR_c_298_n 0.00442186f $X=0.72 $Y=2.885 $X2=0
+ $Y2=0
cc_181 N_A_35_392#_c_245_n N_VPWR_c_299_n 0.0229941f $X=2.5 $Y=2.975 $X2=0 $Y2=0
cc_182 N_A_35_392#_M1002_g N_VPWR_c_299_n 0.0099747f $X=2.575 $Y=2.17 $X2=0
+ $Y2=0
cc_183 N_A_35_392#_M1002_g N_VPWR_c_300_n 0.027543f $X=2.575 $Y=2.17 $X2=0 $Y2=0
cc_184 N_A_35_392#_c_248_n N_VPWR_c_300_n 0.00247229f $X=2.72 $Y=1.775 $X2=0
+ $Y2=0
cc_185 N_A_35_392#_c_250_n N_VPWR_c_301_n 0.0365559f $X=0.72 $Y=2.885 $X2=0
+ $Y2=0
cc_186 N_A_35_392#_c_251_n N_VPWR_c_301_n 0.0109209f $X=0.72 $Y=2.885 $X2=0
+ $Y2=0
cc_187 N_A_35_392#_c_245_n N_VPWR_c_303_n 0.0203319f $X=2.5 $Y=2.975 $X2=0 $Y2=0
cc_188 N_A_35_392#_c_245_n N_VPWR_c_305_n 0.0197672f $X=2.5 $Y=2.975 $X2=0 $Y2=0
cc_189 N_A_35_392#_c_250_n N_VPWR_c_297_n 0.0239192f $X=0.72 $Y=2.885 $X2=0
+ $Y2=0
cc_190 N_A_35_392#_c_251_n N_VPWR_c_297_n 0.0519155f $X=0.72 $Y=2.885 $X2=0
+ $Y2=0
cc_191 N_A_35_392#_M1007_g N_Y_c_333_n 0.00465527f $X=2.72 $Y=0.47 $X2=0 $Y2=0
cc_192 N_A_35_392#_c_248_n Y 0.00105949f $X=2.72 $Y=1.775 $X2=0 $Y2=0
cc_193 N_A_35_392#_M1007_g Y 0.034193f $X=2.72 $Y=0.47 $X2=0 $Y2=0
cc_194 N_A_35_392#_c_248_n Y 0.0129264f $X=2.72 $Y=1.775 $X2=0 $Y2=0
cc_195 N_A_35_392#_c_245_n N_Y_c_343_n 0.00521995f $X=2.5 $Y=2.975 $X2=0 $Y2=0
cc_196 N_A_35_392#_c_245_n N_Y_c_356_n 0.00512826f $X=2.5 $Y=2.975 $X2=0 $Y2=0
cc_197 N_A_35_392#_M1002_g N_Y_c_356_n 0.013473f $X=2.575 $Y=2.17 $X2=0 $Y2=0
cc_198 N_A_35_392#_c_248_n N_Y_c_356_n 0.0055077f $X=2.72 $Y=1.775 $X2=0 $Y2=0
cc_199 N_A_35_392#_M1007_g N_VGND_c_383_n 0.00529003f $X=2.72 $Y=0.47 $X2=0
+ $Y2=0
cc_200 N_A_35_392#_M1007_g N_VGND_c_384_n 0.0109774f $X=2.72 $Y=0.47 $X2=0 $Y2=0
cc_201 N_A_35_392#_c_244_n N_VGND_c_384_n 0.0112283f $X=0.33 $Y=0.535 $X2=0
+ $Y2=0
cc_202 N_A_35_392#_c_244_n N_VGND_c_385_n 0.00970844f $X=0.33 $Y=0.535 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_298_n Y 0.002025f $X=1.07 $Y=2.235 $X2=0 $Y2=0
cc_204 N_VPWR_c_300_n Y 0.00949357f $X=2.79 $Y=2.235 $X2=0 $Y2=0
cc_205 N_VPWR_c_299_n N_Y_c_337_n 0.0087613f $X=1.93 $Y=2.235 $X2=0 $Y2=0
cc_206 N_Y_c_333_n N_VGND_c_383_n 0.0124474f $X=3.12 $Y=0.535 $X2=0 $Y2=0
cc_207 N_Y_c_333_n N_VGND_c_384_n 0.0144952f $X=3.12 $Y=0.535 $X2=0 $Y2=0
