* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfxtp_1 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 a_1157_449# a_1201_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1051_125# a_823_47# a_1137_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_319_123# a_78_123# a_441_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_1459_449# a_628_123# a_1664_65# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND CLK a_628_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_628_123# a_823_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_1657_383# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_1459_449# a_823_47# a_1615_495# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_1657_383# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND a_78_123# a_247_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_319_123# a_628_123# a_1051_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_1051_125# a_1201_99# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 a_1201_99# a_628_123# a_1459_449# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X13 a_1137_125# a_1201_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND a_1051_125# a_1201_99# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 a_464_123# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR a_628_123# a_823_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_1615_495# a_1657_383# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_78_123# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_78_123# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1051_125# a_628_123# a_1157_449# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_319_123# a_823_47# a_1051_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_247_123# D a_319_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_319_123# SCE a_464_123# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_1459_449# a_1657_383# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 a_1201_99# a_823_47# a_1459_449# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND a_1459_449# a_1657_383# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 a_441_491# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_1664_65# a_1657_383# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR SCE a_283_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_283_491# D a_319_123# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 VPWR CLK a_628_123# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
