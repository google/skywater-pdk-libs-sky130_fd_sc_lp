* File: sky130_fd_sc_lp__mux4_m.spice
* Created: Wed Sep  2 10:02:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux4_m.pex.spice"
.subckt sky130_fd_sc_lp__mux4_m  VNB VPB A2 A3 A1 S0 A0 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A0	A0
* S0	S0
* A1	A1
* A3	A3
* A2	A2
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_S0_M1014_g N_A_59_463#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1001 A_273_126# N_A2_M1001_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75000.7 SB=75003.1
+ A=0.063 P=1.14 MULT=1
MM1020 N_A_345_126#_M1020_d N_A_59_463#_M1020_g A_273_126# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1006 A_453_126# N_S0_M1006_g N_A_345_126#_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A3_M1003_g A_453_126# VNB NSHORT L=0.15 W=0.42
+ AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=7.14 NRS=14.28 M=1 R=2.8 SA=75002
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1022 A_616_126# N_A1_M1022_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.06405 PD=0.63 PS=0.725 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.4 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1015 N_A_688_126#_M1015_d N_S0_M1015_g A_616_126# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1016 A_774_126# N_A_59_463#_M1016_g N_A_688_126#_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A0_M1009_g A_774_126# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1018 N_A_1184_171#_M1018_d N_A_1118_37#_M1018_g N_A_688_126#_M1018_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.2247 PD=0.7 PS=1.91 NRD=0 NRS=77.136 M=1
+ R=2.8 SA=75000.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1021 N_A_345_126#_M1021_d N_S1_M1021_g N_A_1184_171#_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_S1_M1025_g N_A_1118_37#_M1025_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_X_M1008_d N_A_1184_171#_M1008_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1023 N_VPWR_M1023_d N_S0_M1023_g N_A_59_463#_M1023_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.10605 AS=0.1113 PD=0.925 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75004 A=0.063 P=1.14 MULT=1
MM1024 A_273_463# N_A2_M1024_g N_VPWR_M1023_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.10605 PD=0.63 PS=0.925 NRD=23.443 NRS=105.533 M=1 R=2.8
+ SA=75000.8 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1000 N_A_345_126#_M1000_d N_S0_M1000_g A_273_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1013 A_431_463# N_A_59_463#_M1013_g N_A_345_126#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A3_M1007_g A_431_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=0.99 PS=0.63 NRD=2.3443 NRS=23.443 M=1 R=2.8 SA=75002
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1011 A_647_463# N_A1_M1011_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=0.99 NRD=23.443 NRS=133.665 M=1 R=2.8
+ SA=75002.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1004 N_A_688_126#_M1004_d N_A_59_463#_M1004_g A_647_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75003.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1017 A_805_463# N_S0_M1017_g N_A_688_126#_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75003.5
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_VPWR_M1019_d N_A0_M1019_g A_805_463# VPB PHIGHVT L=0.15 W=0.42 AD=0.168
+ AS=0.0441 PD=1.64 PS=0.63 NRD=63.3158 NRS=23.443 M=1 R=2.8 SA=75003.9
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1012 N_A_1184_171#_M1012_d N_S1_M1012_g N_A_688_126#_M1012_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.2247 PD=0.7 PS=1.91 NRD=0 NRS=126.632 M=1 R=2.8
+ SA=75000.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_345_126#_M1005_d N_A_1118_37#_M1005_g N_A_1184_171#_M1012_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_S1_M1010_g N_A_1118_37#_M1010_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_1184_171#_M1002_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX26_noxref VNB VPB NWDIODE A=15.9271 P=20.81
c_88 VNB 0 1.4009e-19 $X=0 $Y=0
c_175 VPB 0 6.53158e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__mux4_m.pxi.spice"
*
.ends
*
*
