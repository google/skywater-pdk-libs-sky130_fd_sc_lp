# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__clkbuf_16
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__clkbuf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.008000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.125000 1.815000 1.455000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  3.763200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2.685000 1.920000 9.035000 2.150000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.125000  0.085000 0.420000 0.610000 ;
      RECT 0.125000  1.875000 0.420000 3.245000 ;
      RECT 0.590000  0.280000 0.840000 0.775000 ;
      RECT 0.590000  0.775000 2.550000 0.945000 ;
      RECT 0.590000  1.685000 2.200000 1.855000 ;
      RECT 0.590000  1.855000 0.855000 3.075000 ;
      RECT 1.010000  0.085000 1.290000 0.605000 ;
      RECT 1.025000  2.025000 1.290000 3.245000 ;
      RECT 1.460000  0.280000 1.705000 0.775000 ;
      RECT 1.460000  1.855000 1.710000 3.075000 ;
      RECT 1.875000  0.085000 2.550000 0.605000 ;
      RECT 1.880000  2.025000 2.550000 3.245000 ;
      RECT 1.985000  0.945000 2.550000 1.535000 ;
      RECT 1.985000  1.535000 2.200000 1.685000 ;
      RECT 2.720000  0.275000 2.935000 3.055000 ;
      RECT 3.105000  0.085000 3.415000 0.605000 ;
      RECT 3.105000  1.205000 3.415000 1.535000 ;
      RECT 3.105000  1.875000 3.415000 3.245000 ;
      RECT 3.585000  0.275000 3.795000 3.055000 ;
      RECT 3.965000  0.085000 4.275000 0.605000 ;
      RECT 3.965000  1.205000 4.275000 1.535000 ;
      RECT 3.965000  1.875000 4.275000 3.245000 ;
      RECT 4.445000  0.275000 4.655000 3.055000 ;
      RECT 4.825000  0.085000 5.135000 0.605000 ;
      RECT 4.825000  1.205000 5.135000 1.535000 ;
      RECT 4.825000  1.875000 5.135000 3.245000 ;
      RECT 5.305000  0.275000 5.515000 3.055000 ;
      RECT 5.685000  0.085000 5.995000 0.605000 ;
      RECT 5.685000  1.205000 5.995000 1.535000 ;
      RECT 5.685000  1.875000 5.995000 3.245000 ;
      RECT 6.165000  0.275000 6.375000 3.055000 ;
      RECT 6.545000  0.085000 6.850000 0.605000 ;
      RECT 6.545000  1.205000 6.850000 1.535000 ;
      RECT 6.545000  1.875000 6.850000 3.245000 ;
      RECT 7.020000  0.275000 7.235000 3.055000 ;
      RECT 7.405000  0.085000 7.715000 0.605000 ;
      RECT 7.405000  1.205000 7.715000 1.535000 ;
      RECT 7.405000  1.875000 7.715000 3.245000 ;
      RECT 7.885000  0.275000 8.095000 3.055000 ;
      RECT 8.265000  0.085000 8.575000 0.605000 ;
      RECT 8.265000  1.205000 8.575000 1.535000 ;
      RECT 8.265000  1.875000 8.575000 3.245000 ;
      RECT 8.745000  0.275000 8.955000 3.055000 ;
      RECT 9.125000  0.085000 9.445000 0.605000 ;
      RECT 9.125000  1.875000 9.445000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.020000  1.210000 2.190000 1.380000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.380000  1.210000 2.550000 1.380000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 2.745000  1.950000 2.915000 2.120000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.180000  1.210000 3.350000 1.380000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.605000  1.950000 3.775000 2.120000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.040000  1.210000 4.210000 1.380000 ;
      RECT 4.465000  1.950000 4.635000 2.120000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.900000  1.210000 5.070000 1.380000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.325000  1.950000 5.495000 2.120000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.760000  1.210000 5.930000 1.380000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.185000  1.950000 6.355000 2.120000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.615000  1.210000 6.785000 1.380000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.045000  1.950000 7.215000 2.120000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.480000  1.210000 7.650000 1.380000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 7.905000  1.950000 8.075000 2.120000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.340000  1.210000 8.510000 1.380000 ;
      RECT 8.765000  1.950000 8.935000 2.120000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
    LAYER met1 ;
      RECT 1.960000 1.180000 8.610000 1.410000 ;
  END
END sky130_fd_sc_lp__clkbuf_16
