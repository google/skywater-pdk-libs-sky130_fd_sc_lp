* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1542_428# a_223_119# a_1698_163# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1911_119# a_1542_428# a_1746_137# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 VPWR a_1746_137# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND CLK_N a_113_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_223_119# a_113_57# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_463_449# a_223_119# a_549_449# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_2618_131# a_1746_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VPWR CLK_N a_113_57# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_1698_163# a_1746_137# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_789_78# a_1191_21# a_1018_60# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 VGND SET_B a_1911_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 Q_N a_1746_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND SET_B a_1018_60# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 a_223_119# a_113_57# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VPWR a_789_78# a_1447_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 a_1447_379# a_223_119# a_1542_428# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 a_1447_119# a_113_57# a_1542_428# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 a_2048_428# a_1191_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 VPWR a_2618_131# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VPWR SET_B a_789_78# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 a_1644_506# a_1746_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_1119_379# a_1191_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 a_549_449# a_113_57# a_705_104# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_789_78# a_1447_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 VGND a_1746_137# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_1746_137# a_1542_428# a_2048_428# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X26 a_1018_60# a_549_449# a_789_78# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 a_1746_137# a_1191_21# a_1911_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 a_705_104# a_789_78# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1191_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_549_449# a_223_119# a_709_449# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_709_449# a_789_78# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 Q a_2618_131# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 a_1191_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VGND D a_463_449# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VPWR SET_B a_1746_137# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X36 Q_N a_1746_137# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X37 VGND a_2618_131# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 a_463_449# a_113_57# a_549_449# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X39 a_2618_131# a_1746_137# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VPWR D a_463_449# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X41 a_1542_428# a_113_57# a_1644_506# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X42 Q a_2618_131# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X43 a_789_78# a_549_449# a_1119_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
.ends
