# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__clkinv_16
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__clkinv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  5.544000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.715000 1.180000 10.525000 1.410000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  5.174400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.735000 1.920000 10.485000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.320000  1.835000  0.580000 3.245000 ;
      RECT  0.590000  1.160000  2.305000 1.625000 ;
      RECT  0.755000  1.835000  1.010000 3.055000 ;
      RECT  1.180000  1.835000  1.440000 3.245000 ;
      RECT  1.615000  1.835000  1.870000 3.055000 ;
      RECT  2.035000  0.085000  2.305000 0.725000 ;
      RECT  2.040000  1.835000  2.300000 3.245000 ;
      RECT  2.475000  0.395000  2.730000 3.055000 ;
      RECT  2.900000  0.085000  3.165000 0.725000 ;
      RECT  2.900000  1.160000  3.165000 1.625000 ;
      RECT  2.900000  1.835000  3.160000 3.245000 ;
      RECT  3.335000  0.395000  3.590000 3.055000 ;
      RECT  3.760000  0.085000  4.025000 0.725000 ;
      RECT  3.760000  1.160000  4.025000 1.625000 ;
      RECT  3.760000  1.835000  4.020000 3.245000 ;
      RECT  4.195000  0.395000  4.450000 3.055000 ;
      RECT  4.620000  0.085000  4.885000 0.725000 ;
      RECT  4.620000  1.160000  4.885000 1.625000 ;
      RECT  4.620000  1.835000  4.880000 3.245000 ;
      RECT  5.050000  1.885000  5.310000 3.055000 ;
      RECT  5.055000  0.395000  5.310000 1.885000 ;
      RECT  5.480000  0.085000  5.745000 0.725000 ;
      RECT  5.480000  1.160000  5.745000 1.625000 ;
      RECT  5.480000  1.835000  5.740000 3.245000 ;
      RECT  5.915000  0.395000  6.170000 3.055000 ;
      RECT  6.340000  0.085000  6.605000 0.725000 ;
      RECT  6.340000  1.160000  6.605000 1.625000 ;
      RECT  6.340000  1.835000  6.600000 3.245000 ;
      RECT  6.775000  0.395000  7.030000 3.055000 ;
      RECT  7.200000  0.085000  7.465000 0.725000 ;
      RECT  7.200000  1.160000  7.465000 1.625000 ;
      RECT  7.200000  1.835000  7.460000 3.245000 ;
      RECT  7.635000  0.395000  7.890000 3.055000 ;
      RECT  8.060000  0.085000  8.325000 0.725000 ;
      RECT  8.060000  1.160000  8.325000 1.625000 ;
      RECT  8.060000  1.835000  8.320000 3.245000 ;
      RECT  8.495000  0.395000  8.750000 3.055000 ;
      RECT  8.920000  0.085000  9.185000 0.725000 ;
      RECT  8.920000  1.160000 10.545000 1.625000 ;
      RECT  8.920000  1.835000  9.180000 3.245000 ;
      RECT  9.355000  1.835000  9.610000 3.055000 ;
      RECT  9.780000  1.835000 10.040000 3.245000 ;
      RECT 10.210000  1.835000 10.470000 3.055000 ;
      RECT 10.640000  1.835000 10.895000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  0.775000  1.210000  0.945000 1.380000 ;
      RECT  0.795000  1.950000  0.965000 2.120000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.135000  1.210000  1.305000 1.380000 ;
      RECT  1.495000  1.210000  1.665000 1.380000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  1.655000  1.950000  1.825000 2.120000 ;
      RECT  1.855000  1.210000  2.025000 1.380000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.515000  1.950000  2.685000 2.120000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  2.950000  1.210000  3.120000 1.380000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.375000  1.950000  3.545000 2.120000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.805000  1.210000  3.975000 1.380000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.235000  1.950000  4.405000 2.120000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.670000  1.210000  4.840000 1.380000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.095000  1.950000  5.265000 2.120000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.525000  1.210000  5.695000 1.380000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  5.955000  1.950000  6.125000 2.120000 ;
      RECT  6.390000  1.210000  6.560000 1.380000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.815000  1.950000  6.985000 2.120000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.250000  1.210000  7.420000 1.380000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.675000  1.950000  7.845000 2.120000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.110000  1.210000  8.280000 1.380000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.535000  1.950000  8.705000 2.120000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.215000  1.210000  9.385000 1.380000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.395000  1.950000  9.565000 2.120000 ;
      RECT  9.575000  1.210000  9.745000 1.380000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT  9.935000  1.210000 10.105000 1.380000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.255000  1.950000 10.425000 2.120000 ;
      RECT 10.295000  1.210000 10.465000 1.380000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_lp__clkinv_16
