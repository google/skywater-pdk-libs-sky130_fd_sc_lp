* File: sky130_fd_sc_lp__and2_4.pex.spice
* Created: Wed Sep  2 09:30:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2_4%A 1 3 4 6 7 11
c24 11 0 5.95137e-20 $X=0.29 $Y=1.46
r25 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.46 $X2=0.29 $Y2=1.46
r26 7 11 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=1.46
r27 4 10 51.8702 $w=3.82e-07 $l=3.26795e-07 $layer=POLY_cond $X=0.475 $Y=1.725
+ $X2=0.337 $Y2=1.46
r28 4 6 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.475 $Y=1.725
+ $X2=0.475 $Y2=2.465
r29 1 10 53.132 $w=3.82e-07 $l=3.37009e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.337 $Y2=1.46
r30 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_4%B 3 7 9 12 13
c41 13 0 5.2957e-20 $X=0.925 $Y=1.51
c42 12 0 1.28502e-19 $X=0.925 $Y=1.51
c43 7 0 5.95137e-20 $X=0.905 $Y=2.465
r44 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.675
r45 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.925 $Y2=1.345
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.51 $X2=0.925 $Y2=1.51
r47 9 13 5.55884 $w=4.23e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=1.537
+ $X2=0.925 $Y2=1.537
r48 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.905 $Y=2.465
+ $X2=0.905 $Y2=1.675
r49 3 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.835 $Y=0.655
+ $X2=0.835 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_4%A_27_47# 1 2 9 13 17 21 25 29 33 37 41 43 44
+ 45 47 49 52 54 60 65 72
c114 45 0 1.28502e-19 $X=0.69 $Y=2.1
c115 9 0 5.2957e-20 $X=1.41 $Y=0.655
r116 69 70 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.84 $Y=1.5
+ $X2=2.27 $Y2=1.5
r117 61 72 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.52 $Y=1.5 $X2=2.7
+ $Y2=1.5
r118 61 70 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.52 $Y=1.5
+ $X2=2.27 $Y2=1.5
r119 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.5 $X2=2.52 $Y2=1.5
r120 58 69 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.5 $Y=1.5 $X2=1.84
+ $Y2=1.5
r121 58 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.5 $Y=1.5 $X2=1.41
+ $Y2=1.5
r122 57 60 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=1.5 $Y=1.505
+ $X2=2.52 $Y2=1.505
r123 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.5 $Y=1.5
+ $X2=1.5 $Y2=1.5
r124 55 65 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=1.505
+ $X2=1.275 $Y2=1.505
r125 55 57 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=1.36 $Y=1.505
+ $X2=1.5 $Y2=1.505
r126 53 65 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.275 $Y=1.605
+ $X2=1.275 $Y2=1.505
r127 53 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.275 $Y=1.605
+ $X2=1.275 $Y2=1.93
r128 52 65 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.275 $Y=1.405
+ $X2=1.275 $Y2=1.505
r129 51 52 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.275 $Y=1.155
+ $X2=1.275 $Y2=1.405
r130 50 64 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.785 $Y=2.015
+ $X2=0.69 $Y2=2.015
r131 49 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.19 $Y=2.015
+ $X2=1.275 $Y2=1.93
r132 49 50 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.19 $Y=2.015
+ $X2=0.785 $Y2=2.015
r133 45 64 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.1 $X2=0.69
+ $Y2=2.015
r134 45 47 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=0.69 $Y=2.1
+ $X2=0.69 $Y2=2.91
r135 43 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.19 $Y=1.07
+ $X2=1.275 $Y2=1.155
r136 43 44 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.19 $Y=1.07
+ $X2=0.425 $Y2=1.07
r137 39 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.985
+ $X2=0.425 $Y2=1.07
r138 39 41 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=0.26 $Y=0.985
+ $X2=0.26 $Y2=0.42
r139 35 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.665
+ $X2=2.7 $Y2=1.5
r140 35 37 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.7 $Y=1.665 $X2=2.7
+ $Y2=2.465
r141 31 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.335
+ $X2=2.7 $Y2=1.5
r142 31 33 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.7 $Y=1.335
+ $X2=2.7 $Y2=0.655
r143 27 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.665
+ $X2=2.27 $Y2=1.5
r144 27 29 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.27 $Y=1.665
+ $X2=2.27 $Y2=2.465
r145 23 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.335
+ $X2=2.27 $Y2=1.5
r146 23 25 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.27 $Y=1.335
+ $X2=2.27 $Y2=0.655
r147 19 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=1.665
+ $X2=1.84 $Y2=1.5
r148 19 21 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.84 $Y=1.665
+ $X2=1.84 $Y2=2.465
r149 15 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.84 $Y=1.335
+ $X2=1.84 $Y2=1.5
r150 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.84 $Y=1.335
+ $X2=1.84 $Y2=0.655
r151 11 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.665
+ $X2=1.41 $Y2=1.5
r152 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.41 $Y=1.665
+ $X2=1.41 $Y2=2.465
r153 7 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.335
+ $X2=1.41 $Y2=1.5
r154 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.41 $Y=1.335
+ $X2=1.41 $Y2=0.655
r155 2 64 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.095
r156 2 47 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.91
r157 1 41 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_4%VPWR 1 2 3 4 13 15 21 25 31 36 37 38 39 40 41
+ 43 57 62
r53 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 54 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 48 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.155 $Y2=3.33
r59 48 50 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 47 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 47 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r62 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 44 59 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r64 44 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 43 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=1.155 $Y2=3.33
r66 43 46 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=0.72
+ $Y2=3.33
r67 41 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 41 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 41 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 39 53 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.915 $Y2=3.33
r72 38 56 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=3.08 $Y=3.33 $X2=3.12
+ $Y2=3.33
r73 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=2.915 $Y2=3.33
r74 36 50 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=2.055 $Y2=3.33
r76 35 53 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.22 $Y=3.33
+ $X2=2.64 $Y2=3.33
r77 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=3.33
+ $X2=2.055 $Y2=3.33
r78 31 34 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.915 $Y=2.2
+ $X2=2.915 $Y2=2.95
r79 29 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=3.33
r80 29 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=2.95
r81 25 28 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.2
+ $X2=2.055 $Y2=2.97
r82 23 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=3.33
r83 23 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.055 $Y=3.245
+ $X2=2.055 $Y2=2.97
r84 19 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=3.245
+ $X2=1.155 $Y2=3.33
r85 19 21 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=1.155 $Y=3.245
+ $X2=1.155 $Y2=2.385
r86 15 18 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.26 $Y=2.005
+ $X2=0.26 $Y2=2.95
r87 13 59 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r88 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r89 4 34 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.915 $Y2=2.95
r90 4 31 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.835 $X2=2.915 $Y2=2.2
r91 3 28 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.97
r92 3 25 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=1.835 $X2=2.055 $Y2=2.2
r93 2 21 300 $w=1.7e-07 $l=6.31467e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=1.835 $X2=1.155 $Y2=2.385
r94 1 18 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r95 1 15 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41 42
+ 44 45 49 51
r60 49 51 1.70732 $w=4.03e-07 $l=6e-08 $layer=LI1_cond $X=3.057 $Y=1.235
+ $X2=3.057 $Y2=1.295
r61 44 49 2.49209 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.057 $Y=1.15
+ $X2=3.057 $Y2=1.235
r62 44 45 10.187 $w=4.03e-07 $l=3.58e-07 $layer=LI1_cond $X=3.057 $Y=1.307
+ $X2=3.057 $Y2=1.665
r63 44 51 0.341465 $w=4.03e-07 $l=1.2e-08 $layer=LI1_cond $X=3.057 $Y=1.307
+ $X2=3.057 $Y2=1.295
r64 43 45 3.13009 $w=4.03e-07 $l=1.1e-07 $layer=LI1_cond $X=3.057 $Y=1.775
+ $X2=3.057 $Y2=1.665
r65 40 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.58 $Y=1.86
+ $X2=2.485 $Y2=1.86
r66 39 43 8.41448 $w=1.7e-07 $l=2.40778e-07 $layer=LI1_cond $X=2.855 $Y=1.86
+ $X2=3.057 $Y2=1.775
r67 39 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.855 $Y=1.86
+ $X2=2.58 $Y2=1.86
r68 38 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.58 $Y=1.15
+ $X2=2.485 $Y2=1.15
r69 37 44 5.92239 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=2.855 $Y=1.15
+ $X2=3.057 $Y2=1.15
r70 37 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.855 $Y=1.15
+ $X2=2.58 $Y2=1.15
r71 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.485 $Y=1.98
+ $X2=2.485 $Y2=2.91
r72 31 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=1.945
+ $X2=2.485 $Y2=1.86
r73 31 33 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=2.485 $Y=1.945
+ $X2=2.485 $Y2=1.98
r74 27 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=1.065
+ $X2=2.485 $Y2=1.15
r75 27 29 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=2.485 $Y=1.065
+ $X2=2.485 $Y2=0.42
r76 25 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.39 $Y=1.86
+ $X2=2.485 $Y2=1.86
r77 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.39 $Y=1.86
+ $X2=1.72 $Y2=1.86
r78 23 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.39 $Y=1.15
+ $X2=2.485 $Y2=1.15
r79 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.39 $Y=1.15
+ $X2=1.72 $Y2=1.15
r80 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.625 $Y=1.98
+ $X2=1.625 $Y2=2.91
r81 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.625 $Y=1.945
+ $X2=1.72 $Y2=1.86
r82 17 19 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=1.625 $Y=1.945
+ $X2=1.625 $Y2=1.98
r83 13 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.625 $Y=1.065
+ $X2=1.72 $Y2=1.15
r84 13 15 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=1.625 $Y=1.065
+ $X2=1.625 $Y2=0.42
r85 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.835 $X2=2.485 $Y2=2.91
r86 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.345
+ $Y=1.835 $X2=2.485 $Y2=1.98
r87 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=2.91
r88 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.835 $X2=1.625 $Y2=1.98
r89 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.345
+ $Y=0.235 $X2=2.485 $Y2=0.42
r90 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.235 $X2=1.625 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_4%VGND 1 2 3 12 16 20 23 24 25 26 27 28 30 44
+ 46
r49 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r51 41 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r52 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r53 35 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r54 35 37 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.68
+ $Y2=0
r55 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r56 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r58 30 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.72
+ $Y2=0
r59 28 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r60 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r61 28 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r62 26 40 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.64
+ $Y2=0
r63 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.915
+ $Y2=0
r64 25 43 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.12
+ $Y2=0
r65 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.915
+ $Y2=0
r66 23 37 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.68
+ $Y2=0
r67 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.055
+ $Y2=0
r68 22 40 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.64
+ $Y2=0
r69 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.055
+ $Y2=0
r70 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0
r71 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.38
r72 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0
r73 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.055 $Y=0.085
+ $X2=2.055 $Y2=0.38
r74 10 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r75 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.36
r76 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.775
+ $Y=0.235 $X2=2.915 $Y2=0.38
r77 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.915
+ $Y=0.235 $X2=2.055 $Y2=0.38
r78 1 12 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.235 $X2=1.12 $Y2=0.36
.ends

