# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux4_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__mux4_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.215000 1.140000 4.725000 1.390000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 1.145000 3.685000 1.760000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.550000 1.930000 1.110000 2.190000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.340000 1.930000 2.845000 2.130000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.470000 1.375000 1.290000 1.580000 ;
        RECT 0.470000 1.580000 1.460000 1.760000 ;
        RECT 1.290000 1.760000 1.460000 1.940000 ;
        RECT 1.290000 1.940000 1.680000 2.190000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.660000 0.780000 7.115000 1.825000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.285000 0.280000 7.585000 2.675000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.115000  1.025000 0.725000 1.035000 ;
      RECT 0.115000  1.035000 1.655000 1.195000 ;
      RECT 0.115000  1.195000 1.820000 1.205000 ;
      RECT 0.115000  1.205000 0.300000 2.360000 ;
      RECT 0.115000  2.360000 1.305000 2.530000 ;
      RECT 0.115000  2.530000 0.445000 2.905000 ;
      RECT 0.465000  0.640000 0.725000 1.025000 ;
      RECT 0.615000  2.700000 0.945000 3.245000 ;
      RECT 0.895000  0.085000 1.225000 0.865000 ;
      RECT 1.135000  2.530000 1.305000 2.905000 ;
      RECT 1.135000  2.905000 2.500000 3.075000 ;
      RECT 1.485000  1.205000 1.820000 1.365000 ;
      RECT 1.560000  2.475000 2.160000 2.735000 ;
      RECT 1.630000  1.365000 1.820000 1.685000 ;
      RECT 1.825000  0.640000 2.325000 0.970000 ;
      RECT 1.990000  0.970000 2.325000 1.015000 ;
      RECT 1.990000  1.015000 2.160000 2.475000 ;
      RECT 2.330000  2.300000 3.535000 2.470000 ;
      RECT 2.330000  2.470000 2.500000 2.905000 ;
      RECT 2.655000  0.085000 2.985000 0.970000 ;
      RECT 2.670000  2.640000 2.920000 3.245000 ;
      RECT 3.275000  1.930000 4.900000 2.160000 ;
      RECT 3.275000  2.160000 3.535000 2.300000 ;
      RECT 3.455000  2.640000 3.875000 2.920000 ;
      RECT 3.545000  0.640000 4.035000 0.970000 ;
      RECT 3.705000  2.330000 5.250000 2.500000 ;
      RECT 3.705000  2.500000 3.875000 2.640000 ;
      RECT 3.865000  0.970000 4.035000 1.560000 ;
      RECT 3.865000  1.560000 5.250000 1.730000 ;
      RECT 4.300000  2.670000 4.630000 3.245000 ;
      RECT 4.335000  0.085000 4.665000 0.970000 ;
      RECT 4.920000  2.500000 5.250000 2.840000 ;
      RECT 4.950000  0.670000 5.250000 1.560000 ;
      RECT 5.080000  1.730000 5.250000 2.330000 ;
      RECT 5.145000  0.255000 6.690000 0.500000 ;
      RECT 5.420000  0.670000 5.640000 1.005000 ;
      RECT 5.420000  1.005000 5.610000 2.905000 ;
      RECT 5.420000  2.905000 6.745000 3.075000 ;
      RECT 5.780000  1.175000 6.140000 1.345000 ;
      RECT 5.780000  1.345000 5.950000 2.460000 ;
      RECT 5.780000  2.460000 6.110000 2.735000 ;
      RECT 5.810000  0.670000 6.140000 1.175000 ;
      RECT 6.120000  1.525000 6.490000 1.855000 ;
      RECT 6.300000  1.855000 6.490000 2.060000 ;
      RECT 6.300000  2.060000 6.630000 2.390000 ;
      RECT 6.310000  0.500000 6.690000 0.610000 ;
      RECT 6.310000  0.610000 6.490000 1.525000 ;
      RECT 6.415000  2.780000 6.745000 2.905000 ;
      RECT 6.800000  1.995000 7.095000 2.615000 ;
      RECT 6.860000  0.085000 7.115000 0.610000 ;
      RECT 6.880000  2.615000 7.095000 2.675000 ;
      RECT 6.915000  2.675000 7.095000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  0.840000 2.245000 1.010000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  0.840000 6.085000 1.010000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
    LAYER met1 ;
      RECT 2.015000 0.810000 2.305000 0.855000 ;
      RECT 2.015000 0.855000 6.145000 0.995000 ;
      RECT 2.015000 0.995000 2.305000 1.040000 ;
      RECT 5.855000 0.810000 6.145000 0.855000 ;
      RECT 5.855000 0.995000 6.145000 1.040000 ;
  END
END sky130_fd_sc_lp__mux4_0
END LIBRARY
