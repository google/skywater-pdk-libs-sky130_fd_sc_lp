# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrbn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.210000 2.255000 1.580000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.573300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765000 1.815000 9.515000 3.075000 ;
        RECT 9.010000 0.290000 9.515000 1.140000 ;
        RECT 9.055000 1.140000 9.515000 1.815000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.835000 0.595000 8.095000 1.850000 ;
        RECT 7.835000 1.850000 8.115000 3.075000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.905000 1.170000 6.650000 1.760000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.480000 2.175000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.105000  0.085000 0.435000 0.670000 ;
      RECT 0.150000  2.345000 0.480000 3.245000 ;
      RECT 0.605000  0.340000 0.830000 0.670000 ;
      RECT 0.660000  0.670000 0.830000 1.505000 ;
      RECT 0.660000  1.505000 1.065000 2.175000 ;
      RECT 0.660000  2.175000 0.850000 2.775000 ;
      RECT 0.660000  2.775000 1.735000 3.075000 ;
      RECT 1.035000  0.280000 1.365000 0.760000 ;
      RECT 1.035000  0.760000 1.630000 1.030000 ;
      RECT 1.245000  1.030000 1.630000 1.040000 ;
      RECT 1.245000  1.040000 1.415000 1.775000 ;
      RECT 1.245000  1.775000 1.660000 2.455000 ;
      RECT 1.800000  0.085000 2.020000 1.040000 ;
      RECT 1.835000  1.775000 2.165000 2.435000 ;
      RECT 1.835000  2.435000 2.245000 2.605000 ;
      RECT 1.905000  2.605000 2.245000 3.245000 ;
      RECT 2.190000  0.710000 2.595000 1.040000 ;
      RECT 2.425000  0.265000 4.120000 0.435000 ;
      RECT 2.425000  0.435000 2.595000 0.710000 ;
      RECT 2.425000  1.040000 2.595000 1.775000 ;
      RECT 2.425000  1.775000 2.625000 2.445000 ;
      RECT 2.765000  0.605000 4.515000 0.775000 ;
      RECT 2.765000  0.775000 2.990000 1.210000 ;
      RECT 2.795000  1.515000 3.385000 1.685000 ;
      RECT 2.795000  1.685000 2.965000 2.430000 ;
      RECT 2.795000  2.430000 3.940000 2.705000 ;
      RECT 2.795000  2.705000 3.675000 2.710000 ;
      RECT 3.135000  1.855000 5.255000 2.025000 ;
      RECT 3.135000  2.025000 3.355000 2.260000 ;
      RECT 3.160000  0.945000 3.385000 1.515000 ;
      RECT 3.345000  2.710000 3.675000 3.075000 ;
      RECT 3.555000  0.945000 5.370000 1.175000 ;
      RECT 3.610000  2.195000 3.940000 2.430000 ;
      RECT 4.290000  0.390000 4.515000 0.605000 ;
      RECT 4.400000  2.195000 4.730000 3.245000 ;
      RECT 4.685000  0.085000 4.920000 0.720000 ;
      RECT 4.775000  1.355000 5.735000 1.685000 ;
      RECT 4.925000  2.025000 5.255000 2.260000 ;
      RECT 5.140000  0.390000 5.370000 0.945000 ;
      RECT 5.425000  1.685000 5.735000 1.930000 ;
      RECT 5.425000  1.930000 6.285000 2.100000 ;
      RECT 5.540000  0.255000 5.930000 0.830000 ;
      RECT 5.540000  0.830000 7.080000 1.000000 ;
      RECT 5.540000  1.000000 5.735000 1.355000 ;
      RECT 5.560000  2.270000 5.890000 3.245000 ;
      RECT 6.060000  2.100000 6.285000 3.075000 ;
      RECT 6.390000  0.085000 6.720000 0.660000 ;
      RECT 6.455000  1.930000 6.810000 3.245000 ;
      RECT 6.820000  1.000000 7.080000 1.515000 ;
      RECT 6.900000  0.255000 8.435000 0.425000 ;
      RECT 6.900000  0.425000 7.080000 0.830000 ;
      RECT 6.980000  1.815000 7.665000 2.485000 ;
      RECT 7.250000  0.705000 7.665000 1.035000 ;
      RECT 7.395000  1.035000 7.665000 1.815000 ;
      RECT 8.265000  0.425000 8.435000 1.260000 ;
      RECT 8.265000  1.260000 8.885000 1.590000 ;
      RECT 8.285000  1.815000 8.545000 3.245000 ;
      RECT 8.605000  0.085000 8.840000 1.090000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrbn_1
