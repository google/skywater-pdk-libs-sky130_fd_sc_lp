* NGSPICE file created from sky130_fd_sc_lp__o221ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_794_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.331e+12p pd=1.378e+07u as=8.064e+11p ps=6.32e+06u
M1001 VPWR B1 a_388_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.938e+11p ps=6.3e+06u
M1002 Y C1 a_29_69# VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=1.1172e+12p ps=9.38e+06u
M1003 a_305_65# B1 a_29_69# VNB nshort w=840000u l=150000u
+  ad=1.1508e+12p pd=1.114e+07u as=0p ps=0u
M1004 VPWR C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.0584e+12p ps=9.24e+06u
M1005 a_29_69# C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_305_65# B2 a_29_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_388_367# B2 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_794_367# A2 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_305_65# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=5.376e+11p ps=4.64e+06u
M1010 a_29_69# B1 a_305_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A1 a_305_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_305_65# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_388_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_29_69# B2 a_305_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y C1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_794_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A2 a_305_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y A2 a_794_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y B2 a_388_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

