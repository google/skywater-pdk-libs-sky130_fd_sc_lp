* File: sky130_fd_sc_lp__a32o_4.spice
* Created: Fri Aug 28 10:01:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32o_4.pex.spice"
.subckt sky130_fd_sc_lp__a32o_4  VNB VPB A3 A2 A1 B1 B2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1004 N_X_M1004_d N_A_101_21#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1014 N_X_M1004_d N_A_101_21#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1017 N_X_M1017_d N_A_101_21#_M1017_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1019 N_X_M1017_d N_A_101_21#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1932 PD=1.12 PS=1.3 NRD=0 NRS=12.852 M=1 R=5.6 SA=75001.5
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_511_47#_M1007_d N_A3_M1007_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1932 PD=1.12 PS=1.3 NRD=0 NRS=12.852 M=1 R=5.6 SA=75002.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1026 N_A_511_47#_M1007_d N_A3_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_511_47#_M1001_d N_A2_M1001_g N_A_760_47#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1008 N_A_511_47#_M1001_d N_A2_M1008_g N_A_760_47#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1015 N_A_101_21#_M1015_d N_A1_M1015_g N_A_760_47#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1020 N_A_101_21#_M1015_d N_A1_M1020_g N_A_760_47#_M1020_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_A_101_21#_M1009_d N_B1_M1009_g N_A_1208_65#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1027 N_A_101_21#_M1009_d N_B1_M1027_g N_A_1208_65#_M1027_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_B2_M1005_g N_A_1208_65#_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1005_d N_B2_M1022_g N_A_1208_65#_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A_101_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_101_21#_M1011_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1011_d N_A_101_21#_M1016_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1021_d N_A_101_21#_M1021_g N_X_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1021_d N_A3_M1002_g N_A_511_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A3_M1012_g N_A_511_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1010 N_A_511_367#_M1010_d N_A2_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1018 N_A_511_367#_M1018_d N_A2_M1018_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1006 N_A_511_367#_M1018_d N_A1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2142 PD=1.54 PS=1.6 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1023 N_A_511_367#_M1023_d N_A1_M1023_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2142 PD=1.54 PS=1.6 NRD=0 NRS=9.3772 M=1 R=8.4
+ SA=75001.5 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1024 N_A_101_21#_M1024_d N_B1_M1024_g N_A_511_367#_M1023_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=2.3443 NRS=0 M=1 R=8.4 SA=75002
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1025 N_A_101_21#_M1024_d N_B1_M1025_g N_A_511_367#_M1025_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.2709 PD=1.62 PS=1.69 NRD=10.1455 NRS=11.7215 M=1 R=8.4
+ SA=75002.5 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1003 N_A_511_367#_M1025_s N_B2_M1003_g N_A_101_21#_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2709 AS=0.1764 PD=1.69 PS=1.54 NRD=11.7215 NRS=0 M=1 R=8.4
+ SA=75003.1 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_A_511_367#_M1013_d N_B2_M1013_g N_A_101_21#_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.9271 P=20.81
*
.include "sky130_fd_sc_lp__a32o_4.pxi.spice"
*
.ends
*
*
