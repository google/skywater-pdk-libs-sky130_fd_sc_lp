* File: sky130_fd_sc_lp__dlxtp_lp2.pex.spice
* Created: Wed Sep  2 09:48:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%D 1 3 6 10 13 15 16 17 21 22
r37 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.07 $X2=0.63 $Y2=1.07
r38 16 17 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.65 $Y=1.295
+ $X2=0.65 $Y2=1.665
r39 16 22 7.0081 $w=3.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.65 $Y=1.295
+ $X2=0.65 $Y2=1.07
r40 14 21 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=0.607 $Y=1.388
+ $X2=0.607 $Y2=1.07
r41 14 15 33.9275 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.607 $Y=1.388
+ $X2=0.607 $Y2=1.575
r42 13 21 20.0215 $w=3.75e-07 $l=1.35e-07 $layer=POLY_cond $X=0.607 $Y=0.935
+ $X2=0.607 $Y2=1.07
r43 6 15 241 $w=2.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.545 $Y=2.545 $X2=0.545
+ $Y2=1.575
r44 1 13 24.6308 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=0.785
+ $X2=0.675 $Y2=0.935
r45 1 10 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.855 $Y=0.785
+ $X2=0.855 $Y2=0.495
r46 1 3 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.495 $Y=0.785
+ $X2=0.495 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%GATE 1 3 6 8 12 14 16 17 18 22
r55 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.215 $Y=1.295
+ $X2=1.215 $Y2=1.665
r56 17 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.215
+ $Y=1.34 $X2=1.215 $Y2=1.34
r57 15 22 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.215 $Y=1.325
+ $X2=1.215 $Y2=1.34
r58 15 16 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=1.215 $Y=1.325
+ $X2=1.215 $Y2=1.25
r59 14 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.215 $Y=1.68
+ $X2=1.215 $Y2=1.34
r60 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.645 $Y=1.175
+ $X2=1.645 $Y2=0.495
r61 9 16 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.25
+ $X2=1.215 $Y2=1.25
r62 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.57 $Y=1.25
+ $X2=1.645 $Y2=1.175
r63 8 9 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.57 $Y=1.25 $X2=1.38
+ $Y2=1.25
r64 4 16 13.5877 $w=2.4e-07 $l=1.04283e-07 $layer=POLY_cond $X=1.285 $Y=1.175
+ $X2=1.215 $Y2=1.25
r65 4 6 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.285 $Y=1.175
+ $X2=1.285 $Y2=0.495
r66 1 14 47.383 $w=2.95e-07 $l=3.53129e-07 $layer=POLY_cond $X=1.075 $Y=1.97
+ $X2=1.215 $Y2=1.68
r67 1 3 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.075 $Y=1.97
+ $X2=1.075 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%A_240_409# 1 2 7 8 9 11 15 19 23 27 30 36
+ 40 43 46 48 52
c116 27 0 1.40083e-19 $X=4.325 $Y=0.445
r117 52 60 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.5
+ $X2=4.235 $Y2=1.665
r118 52 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.5
+ $X2=4.235 $Y2=1.335
r119 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.235
+ $Y=1.5 $X2=4.235 $Y2=1.5
r120 48 51 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.235 $Y=1.35
+ $X2=4.235 $Y2=1.5
r121 47 57 22.8653 $w=5.27e-07 $l=2.5e-07 $layer=POLY_cond $X=2.812 $Y=1.43
+ $X2=2.812 $Y2=1.68
r122 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.915
+ $Y=1.43 $X2=2.915 $Y2=1.43
r123 44 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=1.35
+ $X2=2.915 $Y2=1.35
r124 43 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=1.35
+ $X2=4.235 $Y2=1.35
r125 43 44 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=4.07 $Y=1.35
+ $X2=3.08 $Y2=1.35
r126 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.86
+ $Y=1.77 $X2=1.86 $Y2=1.77
r127 36 39 44.5262 $w=3.28e-07 $l=1.275e-06 $layer=LI1_cond $X=1.86 $Y=0.495
+ $X2=1.86 $Y2=1.77
r128 34 39 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.86 $Y=2.025
+ $X2=1.86 $Y2=1.77
r129 30 34 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=1.695 $Y=2.15
+ $X2=1.86 $Y2=2.025
r130 30 32 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=1.695 $Y=2.15
+ $X2=1.34 $Y2=2.15
r131 29 40 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.86 $Y=1.755
+ $X2=1.86 $Y2=1.77
r132 27 59 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=4.325 $Y=0.445
+ $X2=4.325 $Y2=1.335
r133 23 60 231.062 $w=2.5e-07 $l=9.3e-07 $layer=POLY_cond $X=4.195 $Y=2.595
+ $X2=4.195 $Y2=1.665
r134 17 47 32.1846 $w=2.63e-07 $l=2.52357e-07 $layer=POLY_cond $X=2.995 $Y=1.265
+ $X2=2.812 $Y2=1.43
r135 17 19 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.995 $Y=1.265
+ $X2=2.995 $Y2=0.445
r136 13 47 32.1846 $w=2.63e-07 $l=2.46037e-07 $layer=POLY_cond $X=2.635 $Y=1.265
+ $X2=2.812 $Y2=1.43
r137 13 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.635 $Y=1.265
+ $X2=2.635 $Y2=0.445
r138 9 57 36.7095 $w=5.27e-07 $l=3.18174e-07 $layer=POLY_cond $X=2.67 $Y=1.935
+ $X2=2.812 $Y2=1.68
r139 9 11 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.67 $Y=1.935
+ $X2=2.67 $Y2=2.595
r140 8 29 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.025 $Y=1.68
+ $X2=1.86 $Y2=1.755
r141 7 57 32.7418 $w=1.5e-07 $l=2.67e-07 $layer=POLY_cond $X=2.545 $Y=1.68
+ $X2=2.812 $Y2=1.68
r142 7 8 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.545 $Y=1.68
+ $X2=2.025 $Y2=1.68
r143 2 32 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.045 $X2=1.34 $Y2=2.19
r144 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.285 $X2=1.86 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%A_27_57# 1 2 9 13 18 20 23 25 27 31 35 38
+ 39 40 47
r92 40 42 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.24 $Y=2.54
+ $X2=1.24 $Y2=2.67
r93 37 38 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=0.2 $Y=0.725 $X2=0.2
+ $Y2=2.025
r94 35 37 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.28 $Y=0.495
+ $X2=0.28 $Y2=0.725
r95 32 47 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.485 $Y=1.77
+ $X2=3.705 $Y2=1.77
r96 32 44 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.485 $Y=1.77
+ $X2=3.425 $Y2=1.77
r97 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.485
+ $Y=1.77 $X2=3.485 $Y2=1.77
r98 29 31 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=3.485 $Y=2.585
+ $X2=3.485 $Y2=1.77
r99 28 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=2.67
+ $X2=1.24 $Y2=2.67
r100 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.32 $Y=2.67
+ $X2=3.485 $Y2=2.585
r101 27 28 130.155 $w=1.68e-07 $l=1.995e-06 $layer=LI1_cond $X=3.32 $Y=2.67
+ $X2=1.325 $Y2=2.67
r102 26 39 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.54
+ $X2=0.28 $Y2=2.54
r103 25 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=2.54
+ $X2=1.24 $Y2=2.54
r104 25 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.155 $Y=2.54
+ $X2=0.445 $Y2=2.54
r105 21 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.625
+ $X2=0.28 $Y2=2.54
r106 21 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.28 $Y=2.625
+ $X2=0.28 $Y2=2.9
r107 20 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=2.19
+ $X2=0.28 $Y2=2.025
r108 18 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.455
+ $X2=0.28 $Y2=2.54
r109 18 20 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.28 $Y=2.455
+ $X2=0.28 $Y2=2.19
r110 11 47 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.935
+ $X2=3.705 $Y2=1.77
r111 11 13 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.705 $Y=1.935
+ $X2=3.705 $Y2=2.595
r112 7 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=1.605
+ $X2=3.425 $Y2=1.77
r113 7 9 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=3.425 $Y=1.605
+ $X2=3.425 $Y2=0.445
r114 2 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r115 2 20 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r116 1 35 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%A_452_419# 1 2 9 12 15 18 22 26 27 30 33
+ 34 36 37 41
c92 34 0 7.04837e-20 $X=4.775 $Y=1.39
c93 33 0 1.81936e-19 $X=4.775 $Y=1.39
r94 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.775
+ $Y=1.39 $X2=4.775 $Y2=1.39
r95 31 33 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.745 $Y=1.085
+ $X2=4.745 $Y2=1.39
r96 30 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.875 $Y=0.93
+ $X2=3.875 $Y2=0.765
r97 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.875
+ $Y=0.93 $X2=3.875 $Y2=0.93
r98 27 37 8.28018 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=3.87 $Y=0.925
+ $X2=3.71 $Y2=0.925
r99 27 29 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=3.87 $Y=0.925
+ $X2=3.875 $Y2=0.925
r100 26 31 6.88036 $w=3.2e-07 $l=2.17256e-07 $layer=LI1_cond $X=4.61 $Y=0.925
+ $X2=4.745 $Y2=1.085
r101 26 29 26.4702 $w=3.18e-07 $l=7.35e-07 $layer=LI1_cond $X=4.61 $Y=0.925
+ $X2=3.875 $Y2=0.925
r102 25 36 3.89502 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.585 $Y=1
+ $X2=2.412 $Y2=1
r103 25 37 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=2.585 $Y=1
+ $X2=3.71 $Y2=1
r104 20 36 2.82881 $w=3.37e-07 $l=8.84308e-08 $layer=LI1_cond $X=2.405 $Y=1.085
+ $X2=2.412 $Y2=1
r105 20 22 40.3355 $w=3.28e-07 $l=1.155e-06 $layer=LI1_cond $X=2.405 $Y=1.085
+ $X2=2.405 $Y2=2.24
r106 16 36 2.82881 $w=3.37e-07 $l=8.5e-08 $layer=LI1_cond $X=2.412 $Y=0.915
+ $X2=2.412 $Y2=1
r107 16 18 14.8648 $w=3.43e-07 $l=4.45e-07 $layer=LI1_cond $X=2.412 $Y=0.915
+ $X2=2.412 $Y2=0.47
r108 14 34 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.775 $Y=1.73
+ $X2=4.775 $Y2=1.39
r109 14 15 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.775 $Y=1.73
+ $X2=4.775 $Y2=1.895
r110 12 15 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=4.735 $Y=2.595
+ $X2=4.735 $Y2=1.895
r111 9 41 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.815 $Y=0.445
+ $X2=3.815 $Y2=0.765
r112 2 22 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.26
+ $Y=2.095 $X2=2.405 $Y2=2.24
r113 1 18 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.235 $X2=2.42 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%A_928_21# 1 2 7 9 10 11 16 18 19 22 26 30
+ 35 39 40 42 43 47 48 51 52 54 59 64
r123 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.8 $Y=1.2
+ $X2=6.8 $Y2=1.2
r124 54 56 7.24418 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.535 $Y=0.47
+ $X2=6.535 $Y2=0.675
r125 51 52 8.76046 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=6.352 $Y=2.24
+ $X2=6.352 $Y2=2.075
r126 48 52 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.48 $Y=1.875
+ $X2=6.48 $Y2=2.075
r127 47 58 5.8342 $w=4.89e-07 $l=2.21743e-07 $layer=LI1_cond $X=6.547 $Y=1.035
+ $X2=6.68 $Y2=1.2
r128 47 56 13.6026 $w=3.03e-07 $l=3.6e-07 $layer=LI1_cond $X=6.547 $Y=1.035
+ $X2=6.547 $Y2=0.675
r129 42 48 7.64329 $w=4.89e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.395 $Y=1.79
+ $X2=6.48 $Y2=1.875
r130 42 58 14.7198 $w=4.89e-07 $l=7.18505e-07 $layer=LI1_cond $X=6.395 $Y=1.79
+ $X2=6.68 $Y2=1.2
r131 42 43 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.395 $Y=1.79
+ $X2=5.675 $Y2=1.79
r132 40 65 67.6692 $w=4.95e-07 $l=5.05e-07 $layer=POLY_cond $X=5.427 $Y=1.37
+ $X2=5.427 $Y2=1.875
r133 40 64 46.3954 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=5.427 $Y=1.37
+ $X2=5.427 $Y2=1.205
r134 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.51
+ $Y=1.37 $X2=5.51 $Y2=1.37
r135 37 43 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=5.542 $Y=1.705
+ $X2=5.675 $Y2=1.79
r136 37 39 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=5.542 $Y=1.705
+ $X2=5.542 $Y2=1.37
r137 32 59 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.8 $Y=1.185
+ $X2=6.8 $Y2=1.2
r138 28 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.67 $Y=1.035
+ $X2=7.67 $Y2=1.11
r139 28 30 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.67 $Y=1.035
+ $X2=7.67 $Y2=0.625
r140 24 35 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=7.36 $Y=1.11
+ $X2=7.67 $Y2=1.11
r141 24 33 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=7.36 $Y=1.11 $X2=7.31
+ $Y2=1.11
r142 24 26 303.113 $w=2.5e-07 $l=1.22e-06 $layer=POLY_cond $X=7.36 $Y=1.185
+ $X2=7.36 $Y2=2.405
r143 20 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.31 $Y=1.035
+ $X2=7.31 $Y2=1.11
r144 20 22 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.31 $Y=1.035
+ $X2=7.31 $Y2=0.625
r145 19 32 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.965 $Y=1.11
+ $X2=6.8 $Y2=1.185
r146 18 33 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.235 $Y=1.11
+ $X2=7.31 $Y2=1.11
r147 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.235 $Y=1.11
+ $X2=6.965 $Y2=1.11
r148 16 65 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=5.305 $Y=2.595
+ $X2=5.305 $Y2=1.875
r149 12 64 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=5.255 $Y=0.88
+ $X2=5.255 $Y2=1.205
r150 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.18 $Y=0.805
+ $X2=5.255 $Y2=0.88
r151 10 11 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=5.18 $Y=0.805
+ $X2=4.79 $Y2=0.805
r152 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.715 $Y=0.73
+ $X2=4.79 $Y2=0.805
r153 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.715 $Y=0.73
+ $X2=4.715 $Y2=0.445
r154 2 51 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.165
+ $Y=2.095 $X2=6.305 $Y2=2.24
r155 1 54 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=6.395
+ $Y=0.235 $X2=6.535 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%A_778_47# 1 2 9 13 17 23 26 27 33 36 38 39
+ 44 45 47 48
c106 36 0 1.40083e-19 $X=5.145 $Y=0.855
c107 27 0 7.04837e-20 $X=5.06 $Y=0.44
r108 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.05
+ $Y=1.02 $X2=6.05 $Y2=1.02
r109 40 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.23 $Y=0.94
+ $X2=5.145 $Y2=0.94
r110 39 47 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.885 $Y=0.94
+ $X2=6.05 $Y2=0.94
r111 39 40 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.885 $Y=0.94
+ $X2=5.23 $Y2=0.94
r112 37 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=1.025
+ $X2=5.145 $Y2=0.94
r113 37 38 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=5.145 $Y=1.025
+ $X2=5.145 $Y2=2.075
r114 36 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=0.855
+ $X2=5.145 $Y2=0.94
r115 35 36 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.145 $Y=0.585
+ $X2=5.145 $Y2=0.855
r116 34 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.635 $Y=2.16
+ $X2=4.47 $Y2=2.16
r117 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.06 $Y=2.16
+ $X2=5.145 $Y2=2.075
r118 33 34 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.06 $Y=2.16
+ $X2=4.635 $Y2=2.16
r119 27 35 7.43784 $w=2.9e-07 $l=1.8262e-07 $layer=LI1_cond $X=5.06 $Y=0.44
+ $X2=5.145 $Y2=0.585
r120 27 29 37.7524 $w=2.88e-07 $l=9.5e-07 $layer=LI1_cond $X=5.06 $Y=0.44
+ $X2=4.11 $Y2=0.44
r121 25 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.05 $Y=1.36
+ $X2=6.05 $Y2=1.02
r122 25 26 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.05 $Y=1.36
+ $X2=6.05 $Y2=1.525
r123 22 48 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.05 $Y=1.005
+ $X2=6.05 $Y2=1.02
r124 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.05 $Y=0.93
+ $X2=6.32 $Y2=0.93
r125 19 22 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.96 $Y=0.93 $X2=6.05
+ $Y2=0.93
r126 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.32 $Y=0.855
+ $X2=6.32 $Y2=0.93
r127 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=6.32 $Y=0.855
+ $X2=6.32 $Y2=0.445
r128 13 26 265.845 $w=2.5e-07 $l=1.07e-06 $layer=POLY_cond $X=6.04 $Y=2.595
+ $X2=6.04 $Y2=1.525
r129 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.96 $Y=0.855
+ $X2=5.96 $Y2=0.93
r130 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=5.96 $Y=0.855
+ $X2=5.96 $Y2=0.445
r131 2 44 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.32
+ $Y=2.095 $X2=4.47 $Y2=2.24
r132 1 29 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=3.89
+ $Y=0.235 $X2=4.11 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%VPWR 1 2 3 4 17 21 27 31 33 41 46 53 54 57
+ 60 67 70
r76 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r77 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r78 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r79 60 63 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.015 $Y=3.02
+ $X2=3.015 $Y2=3.33
r80 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 54 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=6.96 $Y2=3.33
r82 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r83 51 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.26 $Y=3.33
+ $X2=7.095 $Y2=3.33
r84 51 53 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.26 $Y=3.33
+ $X2=7.92 $Y2=3.33
r85 50 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r86 50 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r87 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r88 47 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.74 $Y=3.33
+ $X2=5.575 $Y2=3.33
r89 47 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.74 $Y=3.33 $X2=6
+ $Y2=3.33
r90 46 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.93 $Y=3.33
+ $X2=7.095 $Y2=3.33
r91 46 49 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=6.93 $Y=3.33 $X2=6
+ $Y2=3.33
r92 45 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r94 42 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=3.33
+ $X2=3.015 $Y2=3.33
r95 42 44 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=3.18 $Y=3.33
+ $X2=5.04 $Y2=3.33
r96 41 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.41 $Y=3.33
+ $X2=5.575 $Y2=3.33
r97 41 44 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.41 $Y=3.33 $X2=5.04
+ $Y2=3.33
r98 40 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r99 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 37 40 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 37 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 36 39 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r104 34 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r105 34 36 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r106 33 63 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=3.33
+ $X2=3.015 $Y2=3.33
r107 33 39 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.85 $Y=3.33
+ $X2=2.64 $Y2=3.33
r108 31 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 31 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r110 27 30 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.095 $Y=2.05
+ $X2=7.095 $Y2=2.76
r111 25 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=3.245
+ $X2=7.095 $Y2=3.33
r112 25 30 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=7.095 $Y=3.245
+ $X2=7.095 $Y2=2.76
r113 21 24 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=5.575 $Y=2.24
+ $X2=5.575 $Y2=2.95
r114 19 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=3.245
+ $X2=5.575 $Y2=3.33
r115 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.575 $Y=3.245
+ $X2=5.575 $Y2=2.95
r116 15 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r117 15 17 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.895
r118 4 30 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.95
+ $Y=1.905 $X2=7.095 $Y2=2.76
r119 4 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.95
+ $Y=1.905 $X2=7.095 $Y2=2.05
r120 3 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=2.095 $X2=5.575 $Y2=2.95
r121 3 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=2.095 $X2=5.575 $Y2=2.24
r122 2 60 600 $w=1.7e-07 $l=1.02914e-06 $layer=licon1_PDIFF $count=1 $X=2.795
+ $Y=2.095 $X2=3.015 $Y2=3.02
r123 1 17 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%Q 1 2 7 8 9 10 11 12 13 21
r20 13 35 0.304088 $w=5.88e-07 $l=1.5e-08 $layer=LI1_cond $X=7.755 $Y=2.775
+ $X2=7.755 $Y2=2.76
r21 12 35 7.19674 $w=5.88e-07 $l=3.55e-07 $layer=LI1_cond $X=7.755 $Y=2.405
+ $X2=7.755 $Y2=2.76
r22 12 31 7.19674 $w=5.88e-07 $l=3.55e-07 $layer=LI1_cond $X=7.755 $Y=2.405
+ $X2=7.755 $Y2=2.05
r23 11 31 0.304088 $w=5.88e-07 $l=1.5e-08 $layer=LI1_cond $X=7.755 $Y=2.035
+ $X2=7.755 $Y2=2.05
r24 10 11 7.50083 $w=5.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.755 $Y=1.665
+ $X2=7.755 $Y2=2.035
r25 9 10 7.50083 $w=5.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.755 $Y=1.295
+ $X2=7.755 $Y2=1.665
r26 8 9 7.50083 $w=5.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.755 $Y=0.925
+ $X2=7.755 $Y2=1.295
r27 8 21 3.85178 $w=5.88e-07 $l=1.9e-07 $layer=LI1_cond $X=7.755 $Y=0.925
+ $X2=7.755 $Y2=0.735
r28 7 21 3.77996 $w=5.9e-07 $l=1.8e-07 $layer=LI1_cond $X=7.755 $Y=0.555
+ $X2=7.755 $Y2=0.735
r29 2 35 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=7.485
+ $Y=1.905 $X2=7.625 $Y2=2.76
r30 2 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.485
+ $Y=1.905 $X2=7.625 $Y2=2.05
r31 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.745
+ $Y=0.415 $X2=7.885 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_LP2%VGND 1 2 3 4 15 17 21 25 29 31 33 38 46 53
+ 54 57 60 63 66
r97 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r98 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r99 60 61 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r100 58 61 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r101 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r102 54 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=6.96
+ $Y2=0
r103 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r104 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.26 $Y=0 $X2=7.095
+ $Y2=0
r105 51 53 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.26 $Y=0 $X2=7.92
+ $Y2=0
r106 50 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r107 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r108 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r109 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.74 $Y=0 $X2=5.575
+ $Y2=0
r110 47 49 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.74 $Y=0 $X2=6
+ $Y2=0
r111 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.93 $Y=0 $X2=7.095
+ $Y2=0
r112 46 49 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=6.93 $Y=0 $X2=6
+ $Y2=0
r113 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r114 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r115 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r116 41 44 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r117 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r118 39 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.21
+ $Y2=0
r119 39 41 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.6
+ $Y2=0
r120 38 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.575
+ $Y2=0
r121 38 44 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.41 $Y=0 $X2=5.04
+ $Y2=0
r122 36 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r123 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r124 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r125 33 35 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r126 31 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r127 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r128 27 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.095 $Y=0.085
+ $X2=7.095 $Y2=0
r129 27 29 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=7.095 $Y=0.085
+ $X2=7.095 $Y2=0.625
r130 23 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0
r131 23 25 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0.445
r132 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r133 19 21 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.445
r134 18 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r135 17 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.21
+ $Y2=0
r136 17 18 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=3.045 $Y=0
+ $X2=1.235 $Y2=0
r137 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r138 13 15 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.495
r139 4 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.95
+ $Y=0.415 $X2=7.095 $Y2=0.625
r140 3 25 182 $w=1.7e-07 $l=8.83784e-07 $layer=licon1_NDIFF $count=1 $X=4.79
+ $Y=0.235 $X2=5.575 $Y2=0.445
r141 2 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.235 $X2=3.21 $Y2=0.445
r142 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.285 $X2=1.07 $Y2=0.495
.ends

