* File: sky130_fd_sc_lp__dlxtp_lp2.spice
* Created: Wed Sep  2 09:48:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxtp_lp2.pex.spice"
.subckt sky130_fd_sc_lp__dlxtp_lp2  VNB VPB D GATE VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1009 A_114_57# N_D_M1009_g N_A_27_57#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_D_M1002_g A_114_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1011 A_272_57# N_GATE_M1011_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_240_409#_M1012_d N_GATE_M1012_g A_272_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 A_542_47# N_A_240_409#_M1017_g N_A_452_419#_M1017_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_240_409#_M1010_g A_542_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1018 A_700_47# N_A_27_57#_M1018_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1021 N_A_778_47#_M1021_d N_A_452_419#_M1021_g A_700_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1000 A_880_47# N_A_240_409#_M1000_g N_A_778_47#_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75001.9 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_928_21#_M1005_g A_880_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.22995 AS=0.0504 PD=1.515 PS=0.66 NRD=184.284 NRS=18.564 M=1 R=2.8
+ SA=75002.3 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1022 A_1207_47# N_A_778_47#_M1022_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.22995 PD=0.63 PS=1.515 NRD=14.28 NRS=48.564 M=1 R=2.8
+ SA=75003.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_928_21#_M1001_d N_A_778_47#_M1001_g A_1207_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75003.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_1477_83# N_A_928_21#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_Q_M1008_d N_A_928_21#_M1008_g A_1477_83# VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_D_M1004_g N_A_27_57#_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1014 N_A_240_409#_M1014_d N_GATE_M1014_g N_VPWR_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1013 N_VPWR_M1013_d N_A_240_409#_M1013_g N_A_452_419#_M1013_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.40265 AS=0.285 PD=1.855 PS=2.57 NRD=16.7253 NRS=0 M=1 R=4
+ SA=125000 SB=125004 A=0.25 P=2.5 MULT=1
MM1003 A_766_419# N_A_27_57#_M1003_g N_VPWR_M1013_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.40265 PD=1.24 PS=1.855 NRD=12.7853 NRS=84.6903 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1015 N_A_778_47#_M1015_d N_A_240_409#_M1015_g A_766_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.145 AS=0.12 PD=1.29 PS=1.24 NRD=1.9503 NRS=12.7853 M=1 R=4 SA=125002
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1019 A_972_419# N_A_452_419#_M1019_g N_A_778_47#_M1015_d VPB PHIGHVT L=0.25
+ W=1 AD=0.16 AS=0.145 PD=1.32 PS=1.29 NRD=20.6653 NRS=0 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1016 N_VPWR_M1016_d N_A_928_21#_M1016_g A_972_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.2425 AS=0.16 PD=1.485 PS=1.32 NRD=0.9653 NRS=20.6653 M=1 R=4 SA=125003
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1020 N_A_928_21#_M1020_d N_A_778_47#_M1020_g N_VPWR_M1016_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.2425 PD=2.57 PS=1.485 NRD=0 NRS=39.4 M=1 R=4 SA=125004
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1007 N_Q_M1007_d N_A_928_21#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX23_noxref VNB VPB NWDIODE A=15.9271 P=20.81
c_137 VPB 0 1.81936e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlxtp_lp2.pxi.spice"
*
.ends
*
*
