* File: sky130_fd_sc_lp__or2_m.pex.spice
* Created: Wed Sep  2 10:29:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2_M%B 2 3 5 6 8 12 15 18 20 21 25
r40 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.295
r41 20 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=0.93 $X2=0.27 $Y2=0.93
r42 16 18 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.36 $Y=1.8
+ $X2=0.655 $Y2=1.8
r43 14 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.27
+ $X2=0.27 $Y2=0.93
r44 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.27
+ $X2=0.27 $Y2=1.435
r45 10 25 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.915
+ $X2=0.27 $Y2=0.93
r46 10 12 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=0.27 $Y=0.84
+ $X2=0.585 $Y2=0.84
r47 6 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.655 $Y=1.875
+ $X2=0.655 $Y2=1.8
r48 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.655 $Y=1.875
+ $X2=0.655 $Y2=2.195
r49 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.585 $Y=0.765
+ $X2=0.585 $Y2=0.84
r50 3 5 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.585 $Y=0.765
+ $X2=0.585 $Y2=0.445
r51 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=1.725
+ $X2=0.36 $Y2=1.8
r52 2 15 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.36 $Y=1.725
+ $X2=0.36 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_M%A 3 7 9 12 13
c36 13 0 1.71584e-19 $X=0.86 $Y=1.32
c37 7 0 4.4852e-21 $X=1.015 $Y=2.195
r38 12 15 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.892 $Y=1.32
+ $X2=0.892 $Y2=1.485
r39 12 14 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.892 $Y=1.32
+ $X2=0.892 $Y2=1.155
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.86
+ $Y=1.32 $X2=0.86 $Y2=1.32
r41 9 13 7.9627 $w=1.93e-07 $l=1.4e-07 $layer=LI1_cond $X=0.72 $Y=1.307 $X2=0.86
+ $Y2=1.307
r42 7 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.015 $Y=2.195
+ $X2=1.015 $Y2=1.485
r43 3 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.015 $Y=0.445
+ $X2=1.015 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_M%A_63_397# 1 2 7 11 14 17 22 24 25 26 29 34 35
c65 11 0 1.71584e-19 $X=1.445 $Y=0.445
r66 33 34 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=2.02
+ $X2=0.945 $Y2=2.02
r67 31 33 7.39394 $w=5.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.44 $Y=2.02
+ $X2=0.78 $Y2=2.02
r68 28 29 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.29 $Y=0.895
+ $X2=1.29 $Y2=1.745
r69 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.205 $Y=1.83
+ $X2=1.29 $Y2=1.745
r70 26 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.205 $Y=1.83
+ $X2=0.945 $Y2=1.83
r71 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.205 $Y=0.81
+ $X2=1.29 $Y2=0.895
r72 24 25 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.205 $Y=0.81
+ $X2=0.905 $Y2=0.81
r73 20 25 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.8 $Y=0.725
+ $X2=0.905 $Y2=0.81
r74 20 22 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=0.8 $Y=0.725 $X2=0.8
+ $Y2=0.51
r75 18 35 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.78 $Y=2.94 $X2=0.78
+ $Y2=2.85
r76 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.78
+ $Y=2.94 $X2=0.78 $Y2=2.94
r77 15 33 3.72573 $w=3.3e-07 $l=2.75e-07 $layer=LI1_cond $X=0.78 $Y=2.295
+ $X2=0.78 $Y2=2.02
r78 15 17 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=0.78 $Y=2.295
+ $X2=0.78 $Y2=2.94
r79 11 14 897.34 $w=1.5e-07 $l=1.75e-06 $layer=POLY_cond $X=1.445 $Y=0.445
+ $X2=1.445 $Y2=2.195
r80 9 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.445 $Y=2.775
+ $X2=1.445 $Y2=2.195
r81 8 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=2.85
+ $X2=0.78 $Y2=2.85
r82 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.37 $Y=2.85
+ $X2=1.445 $Y2=2.775
r83 7 8 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=1.37 $Y=2.85
+ $X2=0.945 $Y2=2.85
r84 2 31 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.315
+ $Y=1.985 $X2=0.44 $Y2=2.13
r85 1 22 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.235 $X2=0.8 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_M%VPWR 1 6 8 10 17 18 21
c23 18 0 4.4852e-21 $X=1.68 $Y=3.33
r24 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r25 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r26 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 15 21 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.23 $Y2=3.33
r28 15 17 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 10 21 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=1.23 $Y2=3.33
r31 10 12 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.125 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 8 13 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 4 21 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r35 4 6 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.26
r36 1 6 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.985 $X2=1.23 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_M%X 1 2 7 8 9 10 11 12 13
r14 12 13 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=2.405
+ $X2=1.66 $Y2=2.775
r15 12 34 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.66 $Y=2.405
+ $X2=1.66 $Y2=2.13
r16 11 34 5.01732 $w=2.08e-07 $l=9.5e-08 $layer=LI1_cond $X=1.66 $Y=2.035
+ $X2=1.66 $Y2=2.13
r17 10 11 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=1.665
+ $X2=1.66 $Y2=2.035
r18 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=1.295
+ $X2=1.66 $Y2=1.665
r19 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=0.925 $X2=1.66
+ $Y2=1.295
r20 7 8 21.9177 $w=2.08e-07 $l=4.15e-07 $layer=LI1_cond $X=1.66 $Y=0.51 $X2=1.66
+ $Y2=0.925
r21 2 34 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.985 $X2=1.66 $Y2=2.13
r22 1 7 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.235 $X2=1.66 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_M%VGND 1 2 7 9 11 15 17 21 22 28
r33 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r34 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 22 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r36 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r37 19 28 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.23
+ $Y2=0
r38 19 21 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.68
+ $Y2=0
r39 17 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r40 17 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r41 13 28 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0
r42 13 15 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0.38
r43 12 25 3.60924 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=0 $X2=0.237
+ $Y2=0
r44 11 28 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.23
+ $Y2=0
r45 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=0.475
+ $Y2=0
r46 7 25 3.30595 $w=2.1e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.237 $Y2=0
r47 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.37 $Y2=0.38
r48 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.38
r49 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.38
.ends

