* File: sky130_fd_sc_lp__sleep_sergate_plv_28.pex.spice
* Created: Fri Aug 28 11:32:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_28%SLEEP 2 4 5 6 8 9 10 12 13 14
+ 16 17 19 21 23 24 25 26 27 34
r80 26 27 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=2.035
+ $X2=8.52 $Y2=2.405
r81 25 26 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=1.665
+ $X2=8.52 $Y2=2.035
r82 24 25 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=1.295
+ $X2=8.52 $Y2=1.665
r83 23 24 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=0.925
+ $X2=8.52 $Y2=1.295
r84 23 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.42
+ $Y=0.965 $X2=8.42 $Y2=0.965
r85 22 34 56.9555 $w=4.15e-07 $l=4.25e-07 $layer=POLY_cond $X=8.377 $Y=1.39
+ $X2=8.377 $Y2=0.965
r86 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=8.205 $Y=1.97
+ $X2=8.205 $Y2=2.25
r87 17 19 1148.77 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=0.98 $Y=2.755
+ $X2=4.555 $Y2=2.755
r88 14 16 1833.14 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=0.98 $Y=2.325
+ $X2=4.555 $Y2=2.325
r89 13 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.13 $Y=2.325
+ $X2=8.205 $Y2=2.25
r90 13 16 1833.14 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=8.13 $Y=2.325
+ $X2=4.555 $Y2=2.325
r91 10 12 1833.14 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=0.98 $Y=1.895
+ $X2=4.555 $Y2=1.895
r92 9 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.13 $Y=1.895
+ $X2=8.205 $Y2=1.97
r93 9 12 1833.14 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=8.13 $Y=1.895
+ $X2=4.555 $Y2=1.895
r94 6 8 1833.14 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=0.98 $Y=1.465
+ $X2=4.555 $Y2=1.465
r95 5 22 35.4752 $w=1.5e-07 $l=2.41607e-07 $layer=POLY_cond $X=8.17 $Y=1.465
+ $X2=8.377 $Y2=1.39
r96 5 8 1853.65 $w=1.5e-07 $l=3.615e-06 $layer=POLY_cond $X=8.17 $Y=1.465
+ $X2=4.555 $Y2=1.465
r97 4 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=2.68
+ $X2=0.98 $Y2=2.755
r98 3 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=2.4
+ $X2=0.98 $Y2=2.325
r99 3 4 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.905 $Y=2.4 $X2=0.905
+ $Y2=2.68
r100 2 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=1.82
+ $X2=0.98 $Y2=1.895
r101 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=1.54
+ $X2=0.98 $Y2=1.465
r102 1 2 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.905 $Y=1.54
+ $X2=0.905 $Y2=1.82
.ends

.subckt PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_28%VIRTPWR 1 2 3 10 14 15 33 69 72
+ 75 78 80 98 102 103 110 111 116 120 125 126
c115 126 0 1.43534e-19 $X=6.51 $Y=3.33
c116 120 0 1.43534e-19 $X=4.955 $Y=3.33
c117 116 0 1.43534e-19 $X=3.4 $Y=3.33
c118 15 0 3.89769e-19 $X=0 $Y=3.085
c119 2 0 2.72043e-19 $X=1.055 $Y=1.97
c120 1 0 1.0636e-20 $X=1.055 $Y=1.085
r121 120 125 0.0432039 $w=4.9e-07 $l=1.55e-07 $layer=MET1_cond $X=4.955 $Y=3.33
+ $X2=4.8 $Y2=3.33
r122 109 130 0.213232 $w=4.9e-07 $l=7.65e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.155 $Y2=3.33
r123 108 110 9.36939 $w=5.73e-07 $l=1.35e-07 $layer=LI1_cond $X=7.92 $Y=3.127
+ $X2=8.055 $Y2=3.127
r124 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r125 106 108 2.80818 $w=5.73e-07 $l=1.35e-07 $layer=LI1_cond $X=7.785 $Y=3.127
+ $X2=7.92 $Y2=3.127
r126 102 110 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=8.055 $Y2=3.33
r127 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r128 95 98 34.5733 $w=2.58e-07 $l=7.8e-07 $layer=LI1_cond $X=7.005 $Y=2.11
+ $X2=7.785 $Y2=2.11
r129 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.005 $Y=2.11
+ $X2=7.005 $Y2=2.11
r130 92 95 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=5.45 $Y=2.11
+ $X2=7.005 $Y2=2.11
r131 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.45 $Y=2.11
+ $X2=5.45 $Y2=2.11
r132 89 92 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.895 $Y=2.11
+ $X2=5.45 $Y2=2.11
r133 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.895 $Y=2.11
+ $X2=3.895 $Y2=2.11
r134 86 89 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=2.34 $Y=2.11
+ $X2=3.895 $Y2=2.11
r135 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.34 $Y=2.11
+ $X2=2.34 $Y2=2.11
r136 83 86 44.9896 $w=2.58e-07 $l=1.015e-06 $layer=LI1_cond $X=1.325 $Y=2.11
+ $X2=2.34 $Y2=2.11
r137 78 96 0.175043 $w=6.45e-07 $l=8.6e-07 $layer=MET1_cond $X=6.832 $Y=1.25
+ $X2=6.832 $Y2=2.11
r138 77 80 34.5733 $w=2.58e-07 $l=7.8e-07 $layer=LI1_cond $X=7.005 $Y=1.25
+ $X2=7.785 $Y2=1.25
r139 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.005 $Y=1.25
+ $X2=7.005 $Y2=1.25
r140 75 93 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=5.267 $Y=1.25
+ $X2=5.267 $Y2=2.11
r141 74 77 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=5.45 $Y=1.25
+ $X2=7.005 $Y2=1.25
r142 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.45 $Y=1.25
+ $X2=5.45 $Y2=1.25
r143 72 90 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=3.712 $Y=1.25
+ $X2=3.712 $Y2=2.11
r144 71 74 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.895 $Y=1.25
+ $X2=5.45 $Y2=1.25
r145 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.895 $Y=1.25
+ $X2=3.895 $Y2=1.25
r146 69 87 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=2.157 $Y=1.25
+ $X2=2.157 $Y2=2.11
r147 68 71 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=2.34 $Y=1.25
+ $X2=3.895 $Y2=1.25
r148 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.34 $Y=1.25
+ $X2=2.34 $Y2=1.25
r149 65 68 44.9896 $w=2.58e-07 $l=1.015e-06 $layer=LI1_cond $X=1.325 $Y=1.25
+ $X2=2.34 $Y2=1.25
r150 63 96 0.175043 $w=6.45e-07 $l=8.6e-07 $layer=MET1_cond $X=6.832 $Y=2.97
+ $X2=6.832 $Y2=2.11
r151 62 63 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.005 $Y=2.97
+ $X2=7.005 $Y2=2.97
r152 60 126 0.00836204 $w=4.9e-07 $l=3e-08 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.51 $Y2=3.33
r153 59 62 10.9207 $w=5.73e-07 $l=5.25e-07 $layer=LI1_cond $X=6.48 $Y=3.127
+ $X2=7.005 $Y2=3.127
r154 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r155 56 59 19.9693 $w=5.73e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=3.127
+ $X2=6.48 $Y2=3.127
r156 54 93 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=5.267 $Y=2.97
+ $X2=5.267 $Y2=2.11
r157 53 56 1.4561 $w=5.73e-07 $l=7e-08 $layer=LI1_cond $X=5.45 $Y=3.127 $X2=5.52
+ $Y2=3.127
r158 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.45 $Y=2.97
+ $X2=5.45 $Y2=2.97
r159 51 125 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.8 $Y2=3.33
r160 50 53 18.5132 $w=5.73e-07 $l=8.9e-07 $layer=LI1_cond $X=4.56 $Y=3.127
+ $X2=5.45 $Y2=3.127
r161 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r162 48 90 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=3.712 $Y=2.97
+ $X2=3.712 $Y2=2.11
r163 47 50 13.8329 $w=5.73e-07 $l=6.65e-07 $layer=LI1_cond $X=3.895 $Y=3.127
+ $X2=4.56 $Y2=3.127
r164 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.895 $Y=2.97
+ $X2=3.895 $Y2=2.97
r165 45 116 0.0780457 $w=4.9e-07 $l=2.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.4 $Y2=3.33
r166 44 47 16.1211 $w=5.73e-07 $l=7.75e-07 $layer=LI1_cond $X=3.12 $Y=3.127
+ $X2=3.895 $Y2=3.127
r167 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r168 41 44 16.2251 $w=5.73e-07 $l=7.8e-07 $layer=LI1_cond $X=2.34 $Y=3.127
+ $X2=3.12 $Y2=3.127
r169 39 87 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=2.157 $Y=2.97
+ $X2=2.157 $Y2=2.11
r170 39 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.34 $Y=2.97
+ $X2=2.34 $Y2=2.97
r171 38 41 7.48849 $w=5.73e-07 $l=3.6e-07 $layer=LI1_cond $X=1.98 $Y=3.127
+ $X2=2.34 $Y2=3.127
r172 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.98 $Y=2.97
+ $X2=1.98 $Y2=2.97
r173 36 111 0.0459912 $w=4.9e-07 $l=1.65e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.845 $Y2=3.33
r174 35 38 6.24041 $w=5.73e-07 $l=3e-07 $layer=LI1_cond $X=1.68 $Y=3.127
+ $X2=1.98 $Y2=3.127
r175 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r176 33 106 0.353623 $w=5.73e-07 $l=1.7e-08 $layer=LI1_cond $X=7.768 $Y=3.127
+ $X2=7.785 $Y2=3.127
r177 33 62 15.8714 $w=5.73e-07 $l=7.63e-07 $layer=LI1_cond $X=7.768 $Y=3.127
+ $X2=7.005 $Y2=3.127
r178 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r179 15 126 0.0661031 $w=4.9e-07 $l=3.22e-07 $layer=MET1_cond $X=6.832 $Y=3.33
+ $X2=6.51 $Y2=3.33
r180 15 130 0.0661031 $w=4.9e-07 $l=3.23e-07 $layer=MET1_cond $X=6.832 $Y=3.33
+ $X2=7.155 $Y2=3.33
r181 15 120 0.0644858 $w=4.9e-07 $l=3.12e-07 $layer=MET1_cond $X=5.267 $Y=3.33
+ $X2=4.955 $Y2=3.33
r182 15 127 0.0644858 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=5.267 $Y=3.33
+ $X2=5.58 $Y2=3.33
r183 15 116 0.0644858 $w=4.9e-07 $l=3.12e-07 $layer=MET1_cond $X=3.712 $Y=3.33
+ $X2=3.4 $Y2=3.33
r184 15 121 0.0644858 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=3.712 $Y=3.33
+ $X2=4.025 $Y2=3.33
r185 15 111 0.0644858 $w=4.9e-07 $l=3.12e-07 $layer=MET1_cond $X=2.157 $Y=3.33
+ $X2=1.845 $Y2=3.33
r186 15 117 0.0644858 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=2.157 $Y=3.33
+ $X2=2.47 $Y2=3.33
r187 15 63 0.044502 $w=1.29e-06 $l=1.15e-07 $layer=MET1_cond $X=6.832 $Y=3.085
+ $X2=6.832 $Y2=2.97
r188 15 54 0.0448765 $w=1.25e-06 $l=1.15e-07 $layer=MET1_cond $X=5.267 $Y=3.085
+ $X2=5.267 $Y2=2.97
r189 15 48 0.0448765 $w=1.25e-06 $l=1.15e-07 $layer=MET1_cond $X=3.712 $Y=3.085
+ $X2=3.712 $Y2=2.97
r190 15 39 0.0448765 $w=1.25e-06 $l=1.15e-07 $layer=MET1_cond $X=2.157 $Y=3.085
+ $X2=2.157 $Y2=2.97
r191 15 103 0.2071 $w=4.9e-07 $l=7.43e-07 $layer=MET1_cond $X=8.137 $Y=3.33
+ $X2=8.88 $Y2=3.33
r192 15 109 0.0604854 $w=4.9e-07 $l=2.17e-07 $layer=MET1_cond $X=8.137 $Y=3.33
+ $X2=7.92 $Y2=3.33
r193 15 60 0.12125 $w=4.9e-07 $l=4.35e-07 $layer=MET1_cond $X=6.045 $Y=3.33
+ $X2=6.48 $Y2=3.33
r194 15 127 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=6.045 $Y=3.33
+ $X2=5.58 $Y2=3.33
r195 15 51 0.0195114 $w=4.9e-07 $l=7e-08 $layer=MET1_cond $X=4.49 $Y=3.33
+ $X2=4.56 $Y2=3.33
r196 15 121 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=4.49 $Y=3.33
+ $X2=4.025 $Y2=3.33
r197 15 45 0.0515659 $w=4.9e-07 $l=1.85e-07 $layer=MET1_cond $X=2.935 $Y=3.33
+ $X2=3.12 $Y2=3.33
r198 15 117 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=2.935 $Y=3.33
+ $X2=2.47 $Y2=3.33
r199 15 36 0.211281 $w=4.9e-07 $l=7.58e-07 $layer=MET1_cond $X=0.922 $Y=3.33
+ $X2=1.68 $Y2=3.33
r200 15 31 0.0563044 $w=4.9e-07 $l=2.02e-07 $layer=MET1_cond $X=0.922 $Y=3.33
+ $X2=0.72 $Y2=3.33
r201 15 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r202 14 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r203 13 14 12.1776 $w=5.73e-07 $l=2.7e-07 $layer=LI1_cond $X=1.325 $Y=3.127
+ $X2=1.055 $Y2=3.127
r204 10 35 7.03086 $w=5.73e-07 $l=3.38e-07 $layer=LI1_cond $X=1.342 $Y=3.127
+ $X2=1.68 $Y2=3.127
r205 10 13 0.353623 $w=5.73e-07 $l=1.7e-08 $layer=LI1_cond $X=1.342 $Y=3.127
+ $X2=1.325 $Y2=3.127
r206 3 106 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.83 $X2=7.785 $Y2=2.97
r207 3 13 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.83 $X2=1.325 $Y2=2.97
r208 2 98 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.97 $X2=7.785 $Y2=2.11
r209 2 83 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.97 $X2=1.325 $Y2=2.11
r210 1 80 60 $w=1.7e-07 $l=6.812e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.085 $X2=7.785 $Y2=1.25
r211 1 65 60 $w=1.7e-07 $l=3.4271e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.085 $X2=1.325 $Y2=1.25
.ends

.subckt PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_28%VPWR 1 2 7 25 45 50 56 62 68 74
+ 75
c108 75 0 1.0636e-20 $X=7.775 $Y=1.68
c109 68 0 9.06808e-20 $X=6.2 $Y=1.68
c110 62 0 9.06808e-20 $X=4.645 $Y=1.68
c111 56 0 9.06808e-20 $X=3.09 $Y=1.68
r112 74 75 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=7.775 $Y=1.68
+ $X2=7.775 $Y2=1.68
r113 69 75 0.0591216 $w=3.33e-06 $l=1.575e-06 $layer=MET2_cond $X=6.2 $Y=1.665
+ $X2=7.775 $Y2=1.665
r114 68 69 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=6.2 $Y=1.68 $X2=6.2
+ $Y2=1.68
r115 63 69 0.0583709 $w=3.33e-06 $l=1.555e-06 $layer=MET2_cond $X=4.645 $Y=1.665
+ $X2=6.2 $Y2=1.665
r116 62 63 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=4.645 $Y=1.68
+ $X2=4.645 $Y2=1.68
r117 56 57 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=3.09 $Y=1.68
+ $X2=3.09 $Y2=1.68
r118 51 57 0.0579955 $w=3.33e-06 $l=1.545e-06 $layer=MET2_cond $X=1.545 $Y=1.665
+ $X2=3.09 $Y2=1.665
r119 50 51 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=1.545 $Y=1.68
+ $X2=1.545 $Y2=1.68
r120 47 74 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=7.62 $Y=2.54
+ $X2=7.62 $Y2=1.68
r121 45 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.8 $Y=2.54
+ $X2=7.8 $Y2=2.54
r122 43 68 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=6.045 $Y=2.54
+ $X2=6.045 $Y2=1.68
r123 42 45 69.1466 $w=2.58e-07 $l=1.56e-06 $layer=LI1_cond $X=6.225 $Y=2.54
+ $X2=7.785 $Y2=2.54
r124 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.225 $Y=2.54
+ $X2=6.225 $Y2=2.54
r125 40 62 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=4.49 $Y=2.54
+ $X2=4.49 $Y2=1.68
r126 39 42 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=4.67 $Y=2.54
+ $X2=6.225 $Y2=2.54
r127 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.67 $Y=2.54
+ $X2=4.67 $Y2=2.54
r128 37 56 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=2.935 $Y=2.54
+ $X2=2.935 $Y2=1.68
r129 36 39 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.115 $Y=2.54
+ $X2=4.67 $Y2=2.54
r130 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.115 $Y=2.54
+ $X2=3.115 $Y2=2.54
r131 34 50 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=1.38 $Y=2.54
+ $X2=1.38 $Y2=1.68
r132 33 36 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=1.56 $Y=2.54
+ $X2=3.115 $Y2=2.54
r133 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.56 $Y=2.54
+ $X2=1.56 $Y2=2.54
r134 30 33 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=1.325 $Y=2.54
+ $X2=1.56 $Y2=2.54
r135 25 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.8 $Y=1.68
+ $X2=7.8 $Y2=1.68
r136 22 25 69.1466 $w=2.58e-07 $l=1.56e-06 $layer=LI1_cond $X=6.225 $Y=1.68
+ $X2=7.785 $Y2=1.68
r137 22 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.225 $Y=1.68
+ $X2=6.225 $Y2=1.68
r138 19 22 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=4.67 $Y=1.68
+ $X2=6.225 $Y2=1.68
r139 19 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.67 $Y=1.68
+ $X2=4.67 $Y2=1.68
r140 16 19 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.115 $Y=1.68
+ $X2=4.67 $Y2=1.68
r141 16 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.115 $Y=1.68
+ $X2=3.115 $Y2=1.68
r142 13 16 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=1.56 $Y=1.68
+ $X2=3.115 $Y2=1.68
r143 13 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.56 $Y=1.68
+ $X2=1.56 $Y2=1.68
r144 10 13 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=1.325 $Y=1.68
+ $X2=1.56 $Y2=1.68
r145 7 63 0.00319069 $w=3.33e-06 $l=8.5e-08 $layer=MET2_cond $X=4.56 $Y=1.665
+ $X2=4.645 $Y2=1.665
r146 7 57 0.0551802 $w=3.33e-06 $l=1.47e-06 $layer=MET2_cond $X=4.56 $Y=1.665
+ $X2=3.09 $Y2=1.665
r147 2 45 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.4 $X2=7.785 $Y2=2.54
r148 2 30 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.4 $X2=1.325 $Y2=2.54
r149 1 25 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.54 $X2=7.785 $Y2=1.68
r150 1 10 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.54 $X2=1.325 $Y2=1.68
.ends

