* File: sky130_fd_sc_lp__o31ai_4.pxi.spice
* Created: Wed Sep  2 10:25:28 2020
* 
x_PM_SKY130_FD_SC_LP__O31AI_4%A2 N_A2_M1004_g N_A2_M1012_g N_A2_M1007_g
+ N_A2_M1020_g N_A2_M1011_g N_A2_M1030_g N_A2_M1024_g N_A2_M1031_g N_A2_c_125_n
+ N_A2_c_126_n N_A2_c_127_n A2 N_A2_c_128_n N_A2_c_129_n N_A2_c_130_n
+ N_A2_c_131_n PM_SKY130_FD_SC_LP__O31AI_4%A2
x_PM_SKY130_FD_SC_LP__O31AI_4%A1 N_A1_M1010_g N_A1_M1001_g N_A1_M1016_g
+ N_A1_M1009_g N_A1_M1027_g N_A1_M1013_g N_A1_M1029_g N_A1_M1026_g N_A1_c_255_n
+ A1 N_A1_c_237_n N_A1_c_238_n N_A1_c_244_n PM_SKY130_FD_SC_LP__O31AI_4%A1
x_PM_SKY130_FD_SC_LP__O31AI_4%A3 N_A3_c_326_n N_A3_M1005_g N_A3_c_336_n
+ N_A3_M1006_g N_A3_c_327_n N_A3_M1017_g N_A3_c_337_n N_A3_M1015_g N_A3_c_338_n
+ N_A3_M1018_g N_A3_c_328_n N_A3_M1019_g N_A3_M1022_g N_A3_M1028_g N_A3_c_340_n
+ N_A3_c_331_n N_A3_c_332_n N_A3_c_333_n N_A3_c_334_n N_A3_c_346_n N_A3_c_342_n
+ A3 A3 N_A3_c_335_n PM_SKY130_FD_SC_LP__O31AI_4%A3
x_PM_SKY130_FD_SC_LP__O31AI_4%B1 N_B1_c_466_n N_B1_M1000_g N_B1_M1008_g
+ N_B1_M1014_g N_B1_c_467_n N_B1_M1002_g N_B1_M1023_g N_B1_c_468_n N_B1_M1003_g
+ N_B1_M1025_g N_B1_c_469_n N_B1_M1021_g N_B1_c_478_n B1 B1 B1 N_B1_c_462_n
+ N_B1_c_463_n N_B1_c_464_n B1 B1 N_B1_c_465_n PM_SKY130_FD_SC_LP__O31AI_4%B1
x_PM_SKY130_FD_SC_LP__O31AI_4%A_49_367# N_A_49_367#_M1012_s N_A_49_367#_M1020_s
+ N_A_49_367#_M1031_s N_A_49_367#_M1015_s N_A_49_367#_M1028_s
+ N_A_49_367#_c_551_n N_A_49_367#_c_552_n N_A_49_367#_c_553_n
+ N_A_49_367#_c_583_n N_A_49_367#_c_554_n N_A_49_367#_c_555_n
+ N_A_49_367#_c_574_n N_A_49_367#_c_575_n N_A_49_367#_c_605_n
+ N_A_49_367#_c_607_n N_A_49_367#_c_610_n N_A_49_367#_c_611_n
+ N_A_49_367#_c_621_n N_A_49_367#_c_624_n N_A_49_367#_c_612_n
+ N_A_49_367#_c_613_n N_A_49_367#_c_627_n N_A_49_367#_c_556_n
+ N_A_49_367#_c_557_n N_A_49_367#_c_558_n N_A_49_367#_c_559_n
+ N_A_49_367#_c_560_n N_A_49_367#_c_579_n N_A_49_367#_c_615_n
+ PM_SKY130_FD_SC_LP__O31AI_4%A_49_367#
x_PM_SKY130_FD_SC_LP__O31AI_4%A_132_367# N_A_132_367#_M1012_d
+ N_A_132_367#_M1009_d N_A_132_367#_M1026_d N_A_132_367#_M1030_d
+ N_A_132_367#_c_700_n N_A_132_367#_c_708_n N_A_132_367#_c_710_n
+ N_A_132_367#_c_701_n N_A_132_367#_c_702_n N_A_132_367#_c_743_p
+ N_A_132_367#_c_733_n N_A_132_367#_c_704_n N_A_132_367#_c_715_n
+ N_A_132_367#_c_705_n PM_SKY130_FD_SC_LP__O31AI_4%A_132_367#
x_PM_SKY130_FD_SC_LP__O31AI_4%VPWR N_VPWR_M1001_s N_VPWR_M1013_s N_VPWR_M1000_d
+ N_VPWR_M1003_d N_VPWR_c_756_n N_VPWR_c_757_n N_VPWR_c_758_n N_VPWR_c_759_n
+ N_VPWR_c_760_n N_VPWR_c_761_n N_VPWR_c_762_n N_VPWR_c_763_n VPWR
+ N_VPWR_c_764_n N_VPWR_c_765_n N_VPWR_c_766_n N_VPWR_c_755_n N_VPWR_c_768_n
+ N_VPWR_c_769_n PM_SKY130_FD_SC_LP__O31AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O31AI_4%Y N_Y_M1008_s N_Y_M1023_s N_Y_M1006_d N_Y_M1018_d
+ N_Y_M1002_s N_Y_M1021_s N_Y_c_882_n N_Y_c_886_n N_Y_c_872_n N_Y_c_893_n
+ N_Y_c_875_n N_Y_c_876_n N_Y_c_873_n N_Y_c_907_n N_Y_c_909_n N_Y_c_924_n
+ N_Y_c_874_n N_Y_c_910_n Y PM_SKY130_FD_SC_LP__O31AI_4%Y
x_PM_SKY130_FD_SC_LP__O31AI_4%VGND N_VGND_M1004_d N_VGND_M1010_d N_VGND_M1027_d
+ N_VGND_M1007_d N_VGND_M1024_d N_VGND_M1017_s N_VGND_M1022_s N_VGND_c_970_n
+ N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n N_VGND_c_974_n N_VGND_c_975_n
+ N_VGND_c_976_n N_VGND_c_977_n N_VGND_c_978_n N_VGND_c_979_n N_VGND_c_980_n
+ N_VGND_c_981_n N_VGND_c_982_n N_VGND_c_983_n VGND N_VGND_c_984_n
+ N_VGND_c_985_n N_VGND_c_986_n N_VGND_c_987_n N_VGND_c_988_n N_VGND_c_989_n
+ N_VGND_c_990_n PM_SKY130_FD_SC_LP__O31AI_4%VGND
x_PM_SKY130_FD_SC_LP__O31AI_4%A_132_47# N_A_132_47#_M1004_s N_A_132_47#_M1016_s
+ N_A_132_47#_M1029_s N_A_132_47#_M1011_s N_A_132_47#_M1005_d
+ N_A_132_47#_M1019_d N_A_132_47#_M1014_d N_A_132_47#_M1025_d
+ N_A_132_47#_c_1098_n N_A_132_47#_c_1101_n N_A_132_47#_c_1102_n
+ N_A_132_47#_c_1164_n N_A_132_47#_c_1103_n N_A_132_47#_c_1171_n
+ N_A_132_47#_c_1104_n N_A_132_47#_c_1178_n N_A_132_47#_c_1094_n
+ N_A_132_47#_c_1182_n N_A_132_47#_c_1095_n N_A_132_47#_c_1186_n
+ N_A_132_47#_c_1135_n N_A_132_47#_c_1111_n N_A_132_47#_c_1112_n
+ N_A_132_47#_c_1096_n N_A_132_47#_c_1097_n N_A_132_47#_c_1131_n
+ PM_SKY130_FD_SC_LP__O31AI_4%A_132_47#
cc_1 VNB N_A2_M1012_g 0.0114093f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_2 VNB N_A2_M1007_g 0.0180956f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=0.655
cc_3 VNB N_A2_M1020_g 0.0036256f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=2.465
cc_4 VNB N_A2_M1011_g 0.0194542f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=0.655
cc_5 VNB N_A2_M1030_g 0.00350909f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=2.465
cc_6 VNB N_A2_M1024_g 0.0190452f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=0.655
cc_7 VNB N_A2_M1031_g 0.00361688f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=2.465
cc_8 VNB N_A2_c_125_n 0.00142948f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.42
cc_9 VNB N_A2_c_126_n 0.00617583f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.16
cc_10 VNB N_A2_c_127_n 0.0447194f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_11 VNB N_A2_c_128_n 0.0196625f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_12 VNB N_A2_c_129_n 0.055593f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.42
cc_13 VNB N_A2_c_130_n 0.0233857f $X=-0.19 $Y=-0.245 $X2=2.46 $Y2=1.29
cc_14 VNB N_A2_c_131_n 0.00993616f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=1.29
cc_15 VNB N_A1_M1010_g 0.0229223f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.655
cc_16 VNB N_A1_M1016_g 0.0227036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_M1027_g 0.0226825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1029_g 0.0228866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_237_n 0.0656156f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=1.42
cc_20 VNB N_A1_c_238_n 0.00166466f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.42
cc_21 VNB N_A3_c_326_n 0.0153693f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.185
cc_22 VNB N_A3_c_327_n 0.0161428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A3_c_328_n 0.0162405f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=1.255
cc_24 VNB N_A3_M1022_g 0.0250536f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=2.465
cc_25 VNB N_A3_M1028_g 0.00297794f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=0.655
cc_26 VNB N_A3_c_331_n 0.00115099f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=2.465
cc_27 VNB N_A3_c_332_n 0.00149609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A3_c_333_n 0.00444461f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.16
cc_29 VNB N_A3_c_334_n 0.0348294f $X=-0.19 $Y=-0.245 $X2=2.985 $Y2=1.415
cc_30 VNB N_A3_c_335_n 0.0780756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B1_M1008_g 0.0203527f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_32 VNB N_B1_M1014_g 0.0197434f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=0.655
cc_33 VNB N_B1_M1023_g 0.0232398f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=0.655
cc_34 VNB N_B1_M1025_g 0.0231501f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.255
cc_35 VNB N_B1_c_462_n 0.112209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B1_c_463_n 0.00477502f $X=-0.19 $Y=-0.245 $X2=2.46 $Y2=1.29
cc_37 VNB N_B1_c_464_n 0.00255845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_B1_c_465_n 0.00238763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_755_n 0.342803f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.29
cc_40 VNB N_Y_c_872_n 0.020881f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.415
cc_41 VNB N_Y_c_873_n 0.024272f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_42 VNB N_Y_c_874_n 0.00262772f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.42
cc_43 VNB N_VGND_c_970_n 0.0137379f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=2.465
cc_44 VNB N_VGND_c_971_n 0.0311599f $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.255
cc_45 VNB N_VGND_c_972_n 3.20903e-19 $X=-0.19 $Y=-0.245 $X2=3.595 $Y2=1.585
cc_46 VNB N_VGND_c_973_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=2.46 $Y2=1.16
cc_47 VNB N_VGND_c_974_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.42
cc_48 VNB N_VGND_c_975_n 3.16879e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_976_n 0.0156709f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_50 VNB N_VGND_c_977_n 0.00497373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_978_n 0.0157256f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_52 VNB N_VGND_c_979_n 0.0285917f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.42
cc_53 VNB N_VGND_c_980_n 0.011684f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=1.42
cc_54 VNB N_VGND_c_981_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=1.42
cc_55 VNB N_VGND_c_982_n 0.0123027f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=1.42
cc_56 VNB N_VGND_c_983_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.42
cc_57 VNB N_VGND_c_984_n 0.0148035f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=1.29
cc_58 VNB N_VGND_c_985_n 0.011684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_986_n 0.0638174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_987_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_988_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_989_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_990_n 0.397298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_132_47#_c_1094_n 0.00790484f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_65 VNB N_A_132_47#_c_1095_n 0.00699782f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=1.42
cc_66 VNB N_A_132_47#_c_1096_n 0.00235487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_132_47#_c_1097_n 0.00176355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VPB N_A2_M1012_g 0.0276354f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_69 VPB N_A2_M1020_g 0.0198907f $X=-0.19 $Y=1.655 $X2=2.735 $Y2=2.465
cc_70 VPB N_A2_M1030_g 0.018695f $X=-0.19 $Y=1.655 $X2=3.165 $Y2=2.465
cc_71 VPB N_A2_M1031_g 0.0188314f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=2.465
cc_72 VPB N_A1_M1001_g 0.0188328f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A1_M1009_g 0.0183595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A1_M1013_g 0.0183595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A1_M1026_g 0.0188084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A1_c_237_n 0.0114717f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=1.42
cc_77 VPB N_A1_c_244_n 0.00260254f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=1.29
cc_78 VPB N_A3_c_336_n 0.0159302f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.515
cc_79 VPB N_A3_c_337_n 0.0152515f $X=-0.19 $Y=1.655 $X2=2.735 $Y2=0.655
cc_80 VPB N_A3_c_338_n 0.0153124f $X=-0.19 $Y=1.655 $X2=2.735 $Y2=2.465
cc_81 VPB N_A3_M1028_g 0.024782f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=0.655
cc_82 VPB N_A3_c_340_n 0.00433217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A3_c_331_n 3.96555e-19 $X=-0.19 $Y=1.655 $X2=3.595 $Y2=2.465
cc_84 VPB N_A3_c_342_n 2.38801e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A3_c_335_n 0.0176733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_B1_c_466_n 0.0173033f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.185
cc_87 VPB N_B1_c_467_n 0.0172424f $X=-0.19 $Y=1.655 $X2=2.735 $Y2=1.585
cc_88 VPB N_B1_c_468_n 0.0170203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_B1_c_469_n 0.017943f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=0.655
cc_90 VPB N_B1_c_462_n 0.0395428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_49_367#_c_551_n 0.0134383f $X=-0.19 $Y=1.655 $X2=3.165 $Y2=1.255
cc_92 VPB N_A_49_367#_c_552_n 0.0412714f $X=-0.19 $Y=1.655 $X2=3.165 $Y2=0.655
cc_93 VPB N_A_49_367#_c_553_n 0.00526475f $X=-0.19 $Y=1.655 $X2=3.165 $Y2=1.585
cc_94 VPB N_A_49_367#_c_554_n 0.00465395f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=1.255
cc_95 VPB N_A_49_367#_c_555_n 0.00555102f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=1.585
cc_96 VPB N_A_49_367#_c_556_n 0.00747154f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=1.42
cc_97 VPB N_A_49_367#_c_557_n 0.0323199f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=1.42
cc_98 VPB N_A_49_367#_c_558_n 0.00154417f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_49_367#_c_559_n 0.00154417f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=1.29
cc_100 VPB N_A_49_367#_c_560_n 0.0030295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_756_n 0.00422004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_757_n 0.00421457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_758_n 0.00441053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_759_n 0.00474504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_760_n 0.0817628f $X=-0.19 $Y=1.655 $X2=3.595 $Y2=2.465
cc_106 VPB N_VPWR_c_761_n 0.00401293f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_762_n 0.018332f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.16
cc_108 VPB N_VPWR_c_763_n 0.00516688f $X=-0.19 $Y=1.655 $X2=2.985 $Y2=1.415
cc_109 VPB N_VPWR_c_764_n 0.0325227f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=1.42
cc_110 VPB N_VPWR_c_765_n 0.017949f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.35
cc_111 VPB N_VPWR_c_766_n 0.0342149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_755_n 0.0502682f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=1.29
cc_113 VPB N_VPWR_c_768_n 0.00362205f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=1.29
cc_114 VPB N_VPWR_c_769_n 0.00362168f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_Y_c_875_n 0.0110796f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.16
cc_116 VPB N_Y_c_876_n 0.00145457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_Y_c_873_n 0.00248763f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.35
cc_118 N_A2_c_126_n N_A1_M1010_g 0.00134267f $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A2_c_128_n N_A1_M1010_g 0.0207824f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_120 N_A2_c_130_n N_A1_M1010_g 0.0105073f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_121 N_A2_M1012_g N_A1_M1001_g 0.0207824f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A2_c_130_n N_A1_M1016_g 0.0105073f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_123 N_A2_c_130_n N_A1_M1027_g 0.0105539f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_124 N_A2_M1007_g N_A1_M1029_g 0.0206156f $X=2.735 $Y=0.655 $X2=0 $Y2=0
cc_125 N_A2_c_130_n N_A1_M1029_g 0.0116297f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_126 N_A2_c_131_n N_A1_M1029_g 0.00627287f $X=2.985 $Y=1.29 $X2=0 $Y2=0
cc_127 N_A2_M1020_g N_A1_M1026_g 0.0206156f $X=2.735 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A2_c_129_n N_A1_c_255_n 6.04026e-19 $X=3.595 $Y=1.42 $X2=0 $Y2=0
cc_129 N_A2_c_131_n N_A1_c_255_n 0.00695325f $X=2.985 $Y=1.29 $X2=0 $Y2=0
cc_130 N_A2_c_127_n N_A1_c_237_n 0.0207824f $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_131 N_A2_c_129_n N_A1_c_237_n 0.0206156f $X=3.595 $Y=1.42 $X2=0 $Y2=0
cc_132 N_A2_c_130_n N_A1_c_237_n 0.00734707f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_133 N_A2_c_126_n N_A1_c_238_n 0.00475906f $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A2_c_127_n N_A1_c_238_n 8.33436e-19 $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_135 N_A2_c_130_n N_A1_c_238_n 0.0917602f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_136 N_A2_M1024_g N_A3_c_326_n 0.0217324f $X=3.595 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A2_M1031_g N_A3_c_336_n 0.0217324f $X=3.595 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A2_c_125_n N_A3_c_346_n 0.00915758f $X=3.505 $Y=1.42 $X2=0 $Y2=0
cc_139 N_A2_c_129_n N_A3_c_346_n 0.00145772f $X=3.595 $Y=1.42 $X2=0 $Y2=0
cc_140 N_A2_c_125_n N_A3_c_335_n 8.15696e-19 $X=3.505 $Y=1.42 $X2=0 $Y2=0
cc_141 N_A2_c_129_n N_A3_c_335_n 0.0217324f $X=3.595 $Y=1.42 $X2=0 $Y2=0
cc_142 N_A2_c_126_n N_A_49_367#_c_551_n 0.00757151f $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A2_c_127_n N_A_49_367#_c_551_n 9.89047e-19 $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_144 N_A2_M1012_g N_A_49_367#_c_553_n 0.0133075f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A2_c_126_n N_A_49_367#_c_553_n 0.0091803f $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A2_c_127_n N_A_49_367#_c_553_n 2.7848e-19 $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_147 N_A2_c_130_n N_A_49_367#_c_553_n 0.00910548f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_148 N_A2_M1020_g N_A_49_367#_c_554_n 0.0132346f $X=2.735 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A2_c_130_n N_A_49_367#_c_554_n 0.00483805f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_150 N_A2_c_131_n N_A_49_367#_c_554_n 0.01963f $X=2.985 $Y=1.29 $X2=0 $Y2=0
cc_151 N_A2_M1030_g N_A_49_367#_c_555_n 0.0143704f $X=3.165 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A2_M1031_g N_A_49_367#_c_555_n 0.0133056f $X=3.595 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A2_c_125_n N_A_49_367#_c_555_n 0.0368147f $X=3.505 $Y=1.42 $X2=0 $Y2=0
cc_154 N_A2_c_129_n N_A_49_367#_c_555_n 0.00241702f $X=3.595 $Y=1.42 $X2=0 $Y2=0
cc_155 N_A2_M1031_g N_A_49_367#_c_574_n 0.00900613f $X=3.595 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A2_M1031_g N_A_49_367#_c_575_n 0.001827f $X=3.595 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A2_M1020_g N_A_49_367#_c_560_n 0.00348079f $X=2.735 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A2_c_129_n N_A_49_367#_c_560_n 0.00252923f $X=3.595 $Y=1.42 $X2=0 $Y2=0
cc_159 N_A2_c_131_n N_A_49_367#_c_560_n 0.0160966f $X=2.985 $Y=1.29 $X2=0 $Y2=0
cc_160 N_A2_M1030_g N_A_49_367#_c_579_n 7.09092e-19 $X=3.165 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A2_M1031_g N_A_49_367#_c_579_n 0.00380694f $X=3.595 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A2_M1012_g N_A_132_367#_c_700_n 0.0069508f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A2_M1020_g N_A_132_367#_c_701_n 0.00643436f $X=2.735 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A2_M1020_g N_A_132_367#_c_702_n 0.011012f $X=2.735 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A2_M1030_g N_A_132_367#_c_702_n 0.012842f $X=3.165 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A2_M1012_g N_A_132_367#_c_704_n 0.00336941f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A2_M1020_g N_A_132_367#_c_705_n 0.00321327f $X=2.735 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A2_M1030_g N_A_132_367#_c_705_n 5.99202e-19 $X=3.165 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A2_M1020_g N_VPWR_c_760_n 0.00357842f $X=2.735 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A2_M1030_g N_VPWR_c_760_n 0.00357877f $X=3.165 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A2_M1031_g N_VPWR_c_760_n 0.00547432f $X=3.595 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A2_M1012_g N_VPWR_c_764_n 0.0054895f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A2_M1012_g N_VPWR_c_755_n 0.0109595f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A2_M1020_g N_VPWR_c_755_n 0.00537652f $X=2.735 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A2_M1030_g N_VPWR_c_755_n 0.0053512f $X=3.165 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A2_M1031_g N_VPWR_c_755_n 0.00990114f $X=3.595 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A2_c_126_n N_VGND_M1004_d 0.00342207f $X=0.495 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A2_c_126_n N_VGND_c_971_n 0.0111207f $X=0.495 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A2_c_127_n N_VGND_c_971_n 7.7301e-19 $X=0.495 $Y=1.35 $X2=0 $Y2=0
cc_180 N_A2_c_128_n N_VGND_c_971_n 0.00318541f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_181 N_A2_c_128_n N_VGND_c_972_n 4.78045e-19 $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_182 N_A2_M1007_g N_VGND_c_973_n 5.37623e-19 $X=2.735 $Y=0.655 $X2=0 $Y2=0
cc_183 N_A2_M1007_g N_VGND_c_974_n 0.00758038f $X=2.735 $Y=0.655 $X2=0 $Y2=0
cc_184 N_A2_M1011_g N_VGND_c_974_n 0.00758038f $X=3.165 $Y=0.655 $X2=0 $Y2=0
cc_185 N_A2_M1024_g N_VGND_c_974_n 5.37623e-19 $X=3.595 $Y=0.655 $X2=0 $Y2=0
cc_186 N_A2_M1011_g N_VGND_c_975_n 5.86e-19 $X=3.165 $Y=0.655 $X2=0 $Y2=0
cc_187 N_A2_M1024_g N_VGND_c_975_n 0.00984813f $X=3.595 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A2_M1007_g N_VGND_c_980_n 0.00365202f $X=2.735 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A2_M1011_g N_VGND_c_982_n 0.00365202f $X=3.165 $Y=0.655 $X2=0 $Y2=0
cc_190 N_A2_M1024_g N_VGND_c_982_n 0.00486043f $X=3.595 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A2_c_128_n N_VGND_c_984_n 0.0054895f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_192 N_A2_M1007_g N_VGND_c_990_n 0.00434777f $X=2.735 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A2_M1011_g N_VGND_c_990_n 0.00432244f $X=3.165 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A2_M1024_g N_VGND_c_990_n 0.00824727f $X=3.595 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A2_c_128_n N_VGND_c_990_n 0.0108123f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_196 N_A2_c_126_n N_A_132_47#_c_1098_n 0.00195985f $X=0.495 $Y=1.16 $X2=0
+ $Y2=0
cc_197 N_A2_c_128_n N_A_132_47#_c_1098_n 0.00214998f $X=0.495 $Y=1.185 $X2=0
+ $Y2=0
cc_198 N_A2_c_130_n N_A_132_47#_c_1098_n 0.0162855f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_199 N_A2_c_128_n N_A_132_47#_c_1101_n 0.00539306f $X=0.495 $Y=1.185 $X2=0
+ $Y2=0
cc_200 N_A2_c_130_n N_A_132_47#_c_1102_n 0.0402256f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_201 N_A2_c_130_n N_A_132_47#_c_1103_n 0.0402256f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_202 N_A2_M1007_g N_A_132_47#_c_1104_n 0.0098539f $X=2.735 $Y=0.655 $X2=0
+ $Y2=0
cc_203 N_A2_M1011_g N_A_132_47#_c_1104_n 0.0112123f $X=3.165 $Y=0.655 $X2=0
+ $Y2=0
cc_204 N_A2_c_125_n N_A_132_47#_c_1104_n 0.00808839f $X=3.505 $Y=1.42 $X2=0
+ $Y2=0
cc_205 N_A2_c_129_n N_A_132_47#_c_1104_n 6.93716e-19 $X=3.595 $Y=1.42 $X2=0
+ $Y2=0
cc_206 N_A2_c_131_n N_A_132_47#_c_1104_n 0.0247296f $X=2.985 $Y=1.29 $X2=0 $Y2=0
cc_207 N_A2_M1024_g N_A_132_47#_c_1094_n 0.0125739f $X=3.595 $Y=0.655 $X2=0
+ $Y2=0
cc_208 N_A2_c_125_n N_A_132_47#_c_1094_n 0.0134448f $X=3.505 $Y=1.42 $X2=0 $Y2=0
cc_209 N_A2_c_130_n N_A_132_47#_c_1111_n 0.0145842f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_210 N_A2_c_130_n N_A_132_47#_c_1112_n 0.0154311f $X=2.46 $Y=1.29 $X2=0 $Y2=0
cc_211 N_A2_M1011_g N_A_132_47#_c_1096_n 7.32965e-19 $X=3.165 $Y=0.655 $X2=0
+ $Y2=0
cc_212 N_A2_c_125_n N_A_132_47#_c_1096_n 0.0160068f $X=3.505 $Y=1.42 $X2=0 $Y2=0
cc_213 N_A2_c_129_n N_A_132_47#_c_1096_n 0.00253619f $X=3.595 $Y=1.42 $X2=0
+ $Y2=0
cc_214 N_A2_c_131_n N_A_132_47#_c_1096_n 0.00463835f $X=2.985 $Y=1.29 $X2=0
+ $Y2=0
cc_215 N_A1_M1001_g N_A_49_367#_c_553_n 0.0100694f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A1_c_238_n N_A_49_367#_c_553_n 0.0115189f $X=1.485 $Y=1.592 $X2=0 $Y2=0
cc_217 N_A1_M1009_g N_A_49_367#_c_583_n 0.00993792f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_218 N_A1_M1013_g N_A_49_367#_c_583_n 0.00993792f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_219 N_A1_c_255_n N_A_49_367#_c_583_n 0.00558926f $X=2.125 $Y=1.51 $X2=0 $Y2=0
cc_220 N_A1_c_237_n N_A_49_367#_c_583_n 5.64665e-19 $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_221 N_A1_c_238_n N_A_49_367#_c_583_n 0.00558926f $X=1.485 $Y=1.592 $X2=0
+ $Y2=0
cc_222 N_A1_c_244_n N_A_49_367#_c_583_n 0.0227178f $X=1.835 $Y=1.592 $X2=0 $Y2=0
cc_223 N_A1_M1026_g N_A_49_367#_c_554_n 0.0110492f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A1_c_255_n N_A_49_367#_c_554_n 0.00655505f $X=2.125 $Y=1.51 $X2=0 $Y2=0
cc_225 N_A1_M1001_g N_A_49_367#_c_558_n 3.30232e-19 $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_226 N_A1_M1009_g N_A_49_367#_c_558_n 8.61679e-19 $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_227 N_A1_c_237_n N_A_49_367#_c_558_n 0.0024237f $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A1_c_238_n N_A_49_367#_c_558_n 0.0103829f $X=1.485 $Y=1.592 $X2=0 $Y2=0
cc_229 N_A1_M1013_g N_A_49_367#_c_559_n 8.61679e-19 $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_230 N_A1_M1026_g N_A_49_367#_c_559_n 3.30232e-19 $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_231 N_A1_c_255_n N_A_49_367#_c_559_n 0.0103829f $X=2.125 $Y=1.51 $X2=0 $Y2=0
cc_232 N_A1_c_237_n N_A_49_367#_c_559_n 0.0024237f $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_233 N_A1_M1001_g N_A_132_367#_c_700_n 0.00784446f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_234 N_A1_M1001_g N_A_132_367#_c_708_n 0.0122718f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_235 N_A1_M1009_g N_A_132_367#_c_708_n 0.01115f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A1_M1013_g N_A_132_367#_c_710_n 0.01115f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A1_M1026_g N_A_132_367#_c_710_n 0.0122718f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_238 N_A1_M1026_g N_A_132_367#_c_701_n 0.00785158f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A1_M1001_g N_A_132_367#_c_704_n 0.00330971f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_A1_M1009_g N_A_132_367#_c_704_n 0.0012135f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_241 N_A1_M1001_g N_A_132_367#_c_715_n 5.66402e-19 $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_242 N_A1_M1009_g N_A_132_367#_c_715_n 0.0100813f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_243 N_A1_M1013_g N_A_132_367#_c_715_n 0.0100813f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_244 N_A1_M1026_g N_A_132_367#_c_715_n 5.66402e-19 $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_245 N_A1_M1013_g N_A_132_367#_c_705_n 0.00115947f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_246 N_A1_M1026_g N_A_132_367#_c_705_n 0.00330971f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_A1_M1001_g N_VPWR_c_756_n 0.00333429f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A1_M1009_g N_VPWR_c_756_n 0.0020641f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A1_M1013_g N_VPWR_c_757_n 0.0020641f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A1_M1026_g N_VPWR_c_757_n 0.00333429f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A1_M1026_g N_VPWR_c_760_n 0.00547432f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_252 N_A1_M1001_g N_VPWR_c_764_n 0.0054895f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_253 N_A1_M1009_g N_VPWR_c_765_n 0.0054895f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_254 N_A1_M1013_g N_VPWR_c_765_n 0.0054895f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_255 N_A1_M1001_g N_VPWR_c_755_n 0.00989836f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_256 N_A1_M1009_g N_VPWR_c_755_n 0.00987303f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A1_M1013_g N_VPWR_c_755_n 0.00987303f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A1_M1026_g N_VPWR_c_755_n 0.0098613f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A1_M1010_g N_VGND_c_972_n 0.00773856f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_260 N_A1_M1016_g N_VGND_c_972_n 0.00758038f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_261 N_A1_M1027_g N_VGND_c_972_n 5.37623e-19 $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_262 N_A1_M1016_g N_VGND_c_973_n 5.37623e-19 $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_263 N_A1_M1027_g N_VGND_c_973_n 0.00758038f $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_264 N_A1_M1029_g N_VGND_c_973_n 0.00758038f $X=2.305 $Y=0.655 $X2=0 $Y2=0
cc_265 N_A1_M1029_g N_VGND_c_974_n 5.37623e-19 $X=2.305 $Y=0.655 $X2=0 $Y2=0
cc_266 N_A1_M1029_g N_VGND_c_980_n 0.00365202f $X=2.305 $Y=0.655 $X2=0 $Y2=0
cc_267 N_A1_M1010_g N_VGND_c_984_n 0.00365202f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_268 N_A1_M1016_g N_VGND_c_985_n 0.00365202f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_269 N_A1_M1027_g N_VGND_c_985_n 0.00365202f $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_270 N_A1_M1010_g N_VGND_c_990_n 0.00434777f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_271 N_A1_M1016_g N_VGND_c_990_n 0.00432244f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_272 N_A1_M1027_g N_VGND_c_990_n 0.00432244f $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_273 N_A1_M1029_g N_VGND_c_990_n 0.00434777f $X=2.305 $Y=0.655 $X2=0 $Y2=0
cc_274 N_A1_M1010_g N_A_132_47#_c_1102_n 0.00990046f $X=1.015 $Y=0.655 $X2=0
+ $Y2=0
cc_275 N_A1_M1016_g N_A_132_47#_c_1102_n 0.00990046f $X=1.445 $Y=0.655 $X2=0
+ $Y2=0
cc_276 N_A1_M1027_g N_A_132_47#_c_1103_n 0.00990046f $X=1.875 $Y=0.655 $X2=0
+ $Y2=0
cc_277 N_A1_M1029_g N_A_132_47#_c_1103_n 0.00990046f $X=2.305 $Y=0.655 $X2=0
+ $Y2=0
cc_278 N_A3_c_338_n N_B1_c_466_n 0.018702f $X=4.885 $Y=1.725 $X2=-0.19
+ $Y2=-0.245
cc_279 N_A3_c_340_n N_B1_c_466_n 0.00823282f $X=7.11 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_280 N_A3_c_328_n N_B1_M1008_g 0.0195803f $X=4.955 $Y=1.185 $X2=0 $Y2=0
cc_281 N_A3_c_340_n N_B1_c_467_n 0.00827107f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_282 N_A3_c_340_n N_B1_c_468_n 0.00816755f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_283 N_A3_M1022_g N_B1_M1025_g 0.0230499f $X=7.475 $Y=0.655 $X2=0 $Y2=0
cc_284 N_A3_c_340_n N_B1_c_469_n 0.00768636f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_285 N_A3_c_332_n N_B1_c_478_n 0.0142669f $X=7.28 $Y=1.435 $X2=0 $Y2=0
cc_286 N_A3_M1028_g N_B1_c_462_n 0.0358729f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A3_c_340_n N_B1_c_462_n 0.0472875f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_288 N_A3_c_331_n N_B1_c_462_n 0.0100888f $X=7.195 $Y=1.695 $X2=0 $Y2=0
cc_289 N_A3_c_332_n N_B1_c_462_n 0.00604522f $X=7.28 $Y=1.435 $X2=0 $Y2=0
cc_290 N_A3_c_334_n N_B1_c_462_n 0.0169989f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_291 N_A3_c_342_n N_B1_c_462_n 0.00190876f $X=5.005 $Y=1.595 $X2=0 $Y2=0
cc_292 N_A3_c_335_n N_B1_c_462_n 0.0483637f $X=4.885 $Y=1.455 $X2=0 $Y2=0
cc_293 N_A3_c_340_n N_B1_c_463_n 0.0938151f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_294 N_A3_c_340_n N_B1_c_464_n 0.0249652f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_295 N_A3_c_342_n N_B1_c_464_n 0.0124869f $X=5.005 $Y=1.595 $X2=0 $Y2=0
cc_296 N_A3_c_335_n N_B1_c_464_n 0.00147404f $X=4.885 $Y=1.455 $X2=0 $Y2=0
cc_297 N_A3_c_332_n N_B1_c_465_n 3.26445e-19 $X=7.28 $Y=1.435 $X2=0 $Y2=0
cc_298 N_A3_c_346_n N_A_49_367#_M1015_s 0.00162309f $X=4.735 $Y=1.595 $X2=0
+ $Y2=0
cc_299 N_A3_c_346_n N_A_49_367#_c_555_n 0.0140819f $X=4.735 $Y=1.595 $X2=0 $Y2=0
cc_300 N_A3_c_335_n N_A_49_367#_c_555_n 0.0014302f $X=4.885 $Y=1.455 $X2=0 $Y2=0
cc_301 N_A3_c_336_n N_A_49_367#_c_574_n 0.00891749f $X=4.025 $Y=1.725 $X2=0
+ $Y2=0
cc_302 N_A3_c_337_n N_A_49_367#_c_574_n 5.82232e-19 $X=4.455 $Y=1.725 $X2=0
+ $Y2=0
cc_303 N_A3_c_336_n N_A_49_367#_c_575_n 0.00284964f $X=4.025 $Y=1.725 $X2=0
+ $Y2=0
cc_304 N_A3_c_336_n N_A_49_367#_c_605_n 0.0105205f $X=4.025 $Y=1.725 $X2=0 $Y2=0
cc_305 N_A3_c_337_n N_A_49_367#_c_605_n 0.0105205f $X=4.455 $Y=1.725 $X2=0 $Y2=0
cc_306 N_A3_c_336_n N_A_49_367#_c_607_n 5.0443e-19 $X=4.025 $Y=1.725 $X2=0 $Y2=0
cc_307 N_A3_c_337_n N_A_49_367#_c_607_n 0.00724644f $X=4.455 $Y=1.725 $X2=0
+ $Y2=0
cc_308 N_A3_c_338_n N_A_49_367#_c_607_n 0.00729178f $X=4.885 $Y=1.725 $X2=0
+ $Y2=0
cc_309 N_A3_c_338_n N_A_49_367#_c_610_n 0.0107439f $X=4.885 $Y=1.725 $X2=0 $Y2=0
cc_310 N_A3_c_338_n N_A_49_367#_c_611_n 5.0844e-19 $X=4.885 $Y=1.725 $X2=0 $Y2=0
cc_311 N_A3_M1028_g N_A_49_367#_c_612_n 6.0375e-19 $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_312 N_A3_M1028_g N_A_49_367#_c_613_n 0.0106978f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_313 N_A3_c_336_n N_A_49_367#_c_579_n 0.00331073f $X=4.025 $Y=1.725 $X2=0
+ $Y2=0
cc_314 N_A3_c_337_n N_A_49_367#_c_615_n 7.56199e-19 $X=4.455 $Y=1.725 $X2=0
+ $Y2=0
cc_315 N_A3_c_338_n N_A_49_367#_c_615_n 6.03807e-19 $X=4.885 $Y=1.725 $X2=0
+ $Y2=0
cc_316 N_A3_c_340_n N_VPWR_M1000_d 0.00464606f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_317 N_A3_c_340_n N_VPWR_M1003_d 0.00421982f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_318 N_A3_c_336_n N_VPWR_c_760_n 0.00357842f $X=4.025 $Y=1.725 $X2=0 $Y2=0
cc_319 N_A3_c_337_n N_VPWR_c_760_n 0.00357842f $X=4.455 $Y=1.725 $X2=0 $Y2=0
cc_320 N_A3_c_338_n N_VPWR_c_760_n 0.00357842f $X=4.885 $Y=1.725 $X2=0 $Y2=0
cc_321 N_A3_M1028_g N_VPWR_c_766_n 0.00359964f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A3_c_336_n N_VPWR_c_755_n 0.00537652f $X=4.025 $Y=1.725 $X2=0 $Y2=0
cc_323 N_A3_c_337_n N_VPWR_c_755_n 0.00535118f $X=4.455 $Y=1.725 $X2=0 $Y2=0
cc_324 N_A3_c_338_n N_VPWR_c_755_n 0.00537847f $X=4.885 $Y=1.725 $X2=0 $Y2=0
cc_325 N_A3_M1028_g N_VPWR_c_755_n 0.00659593f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_326 N_A3_c_346_n N_Y_M1006_d 0.0018284f $X=4.735 $Y=1.595 $X2=0 $Y2=0
cc_327 N_A3_c_340_n N_Y_M1018_d 0.00176461f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_328 N_A3_c_340_n N_Y_M1002_s 0.00176891f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_329 N_A3_c_340_n N_Y_M1021_s 7.51328e-19 $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_330 N_A3_c_337_n N_Y_c_882_n 0.0125619f $X=4.455 $Y=1.725 $X2=0 $Y2=0
cc_331 N_A3_c_338_n N_Y_c_882_n 0.0125125f $X=4.885 $Y=1.725 $X2=0 $Y2=0
cc_332 N_A3_c_346_n N_Y_c_882_n 0.0355274f $X=4.735 $Y=1.595 $X2=0 $Y2=0
cc_333 N_A3_c_335_n N_Y_c_882_n 4.97251e-19 $X=4.885 $Y=1.455 $X2=0 $Y2=0
cc_334 N_A3_c_340_n N_Y_c_886_n 0.118594f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_335 N_A3_c_333_n N_Y_c_886_n 0.00189518f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_336 N_A3_M1022_g N_Y_c_872_n 0.0161057f $X=7.475 $Y=0.655 $X2=0 $Y2=0
cc_337 N_A3_c_340_n N_Y_c_872_n 0.00494665f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_338 N_A3_c_332_n N_Y_c_872_n 0.0139851f $X=7.28 $Y=1.435 $X2=0 $Y2=0
cc_339 N_A3_c_333_n N_Y_c_872_n 0.0316716f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_340 N_A3_c_334_n N_Y_c_872_n 0.00496258f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_341 N_A3_M1028_g N_Y_c_893_n 0.00809207f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_342 N_A3_M1028_g N_Y_c_875_n 0.0093624f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_343 N_A3_c_333_n N_Y_c_875_n 0.00618094f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_344 N_A3_c_334_n N_Y_c_875_n 2.43542e-19 $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_345 N_A3_M1028_g N_Y_c_876_n 0.00353134f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_346 N_A3_c_340_n N_Y_c_876_n 0.0141755f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_347 N_A3_c_333_n N_Y_c_876_n 0.0135464f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_348 N_A3_c_334_n N_Y_c_876_n 0.00291923f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_349 N_A3_M1022_g N_Y_c_873_n 0.00314509f $X=7.475 $Y=0.655 $X2=0 $Y2=0
cc_350 N_A3_M1028_g N_Y_c_873_n 0.00231132f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_351 N_A3_c_340_n N_Y_c_873_n 3.29223e-19 $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_352 N_A3_c_331_n N_Y_c_873_n 0.00489499f $X=7.195 $Y=1.695 $X2=0 $Y2=0
cc_353 N_A3_c_333_n N_Y_c_873_n 0.0157834f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_354 N_A3_c_334_n N_Y_c_873_n 0.0056433f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_355 N_A3_c_346_n N_Y_c_907_n 0.0146785f $X=4.735 $Y=1.595 $X2=0 $Y2=0
cc_356 N_A3_c_335_n N_Y_c_907_n 5.59398e-19 $X=4.885 $Y=1.455 $X2=0 $Y2=0
cc_357 N_A3_c_340_n N_Y_c_909_n 0.0135217f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_358 N_A3_M1028_g N_Y_c_910_n 0.00318133f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_359 N_A3_c_333_n N_Y_c_910_n 0.00453424f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_360 N_A3_c_334_n N_Y_c_910_n 0.00159968f $X=7.555 $Y=1.44 $X2=0 $Y2=0
cc_361 N_A3_M1028_g Y 0.00748344f $X=7.635 $Y=2.465 $X2=0 $Y2=0
cc_362 N_A3_c_326_n N_VGND_c_975_n 0.0114092f $X=4.025 $Y=1.185 $X2=0 $Y2=0
cc_363 N_A3_c_327_n N_VGND_c_975_n 0.00106269f $X=4.455 $Y=1.185 $X2=0 $Y2=0
cc_364 N_A3_c_326_n N_VGND_c_976_n 0.00486043f $X=4.025 $Y=1.185 $X2=0 $Y2=0
cc_365 N_A3_c_327_n N_VGND_c_976_n 0.00585385f $X=4.455 $Y=1.185 $X2=0 $Y2=0
cc_366 N_A3_c_327_n N_VGND_c_977_n 0.0016985f $X=4.455 $Y=1.185 $X2=0 $Y2=0
cc_367 N_A3_c_328_n N_VGND_c_977_n 0.00326196f $X=4.955 $Y=1.185 $X2=0 $Y2=0
cc_368 N_A3_M1022_g N_VGND_c_979_n 0.0158569f $X=7.475 $Y=0.655 $X2=0 $Y2=0
cc_369 N_A3_c_328_n N_VGND_c_986_n 0.00583607f $X=4.955 $Y=1.185 $X2=0 $Y2=0
cc_370 N_A3_M1022_g N_VGND_c_986_n 0.0054895f $X=7.475 $Y=0.655 $X2=0 $Y2=0
cc_371 N_A3_c_326_n N_VGND_c_990_n 0.00835506f $X=4.025 $Y=1.185 $X2=0 $Y2=0
cc_372 N_A3_c_327_n N_VGND_c_990_n 0.0108286f $X=4.455 $Y=1.185 $X2=0 $Y2=0
cc_373 N_A3_c_328_n N_VGND_c_990_n 0.0106841f $X=4.955 $Y=1.185 $X2=0 $Y2=0
cc_374 N_A3_M1022_g N_VGND_c_990_n 0.0110886f $X=7.475 $Y=0.655 $X2=0 $Y2=0
cc_375 N_A3_c_326_n N_A_132_47#_c_1094_n 0.0142444f $X=4.025 $Y=1.185 $X2=0
+ $Y2=0
cc_376 N_A3_c_346_n N_A_132_47#_c_1094_n 0.0128082f $X=4.735 $Y=1.595 $X2=0
+ $Y2=0
cc_377 N_A3_c_327_n N_A_132_47#_c_1095_n 0.0133867f $X=4.455 $Y=1.185 $X2=0
+ $Y2=0
cc_378 N_A3_c_328_n N_A_132_47#_c_1095_n 0.0143793f $X=4.955 $Y=1.185 $X2=0
+ $Y2=0
cc_379 N_A3_c_340_n N_A_132_47#_c_1095_n 0.00851148f $X=7.11 $Y=1.78 $X2=0 $Y2=0
cc_380 N_A3_c_346_n N_A_132_47#_c_1095_n 0.0477041f $X=4.735 $Y=1.595 $X2=0
+ $Y2=0
cc_381 N_A3_c_335_n N_A_132_47#_c_1095_n 0.00510687f $X=4.885 $Y=1.455 $X2=0
+ $Y2=0
cc_382 N_A3_c_327_n N_A_132_47#_c_1097_n 9.43578e-19 $X=4.455 $Y=1.185 $X2=0
+ $Y2=0
cc_383 N_A3_c_346_n N_A_132_47#_c_1097_n 0.0196395f $X=4.735 $Y=1.595 $X2=0
+ $Y2=0
cc_384 N_A3_c_335_n N_A_132_47#_c_1097_n 0.00304738f $X=4.885 $Y=1.455 $X2=0
+ $Y2=0
cc_385 N_A3_M1022_g N_A_132_47#_c_1131_n 0.00674724f $X=7.475 $Y=0.655 $X2=0
+ $Y2=0
cc_386 N_B1_c_466_n N_A_49_367#_c_607_n 5.50549e-19 $X=5.315 $Y=1.725 $X2=0
+ $Y2=0
cc_387 N_B1_c_466_n N_A_49_367#_c_610_n 0.0112675f $X=5.315 $Y=1.725 $X2=0 $Y2=0
cc_388 N_B1_c_466_n N_A_49_367#_c_611_n 0.00833397f $X=5.315 $Y=1.725 $X2=0
+ $Y2=0
cc_389 N_B1_c_467_n N_A_49_367#_c_611_n 0.00299888f $X=6.015 $Y=1.725 $X2=0
+ $Y2=0
cc_390 N_B1_c_467_n N_A_49_367#_c_621_n 0.0135152f $X=6.015 $Y=1.725 $X2=0 $Y2=0
cc_391 N_B1_c_468_n N_A_49_367#_c_621_n 0.0133892f $X=6.445 $Y=1.725 $X2=0 $Y2=0
cc_392 N_B1_c_469_n N_A_49_367#_c_621_n 0.00804271f $X=7.105 $Y=1.725 $X2=0
+ $Y2=0
cc_393 N_B1_c_466_n N_A_49_367#_c_624_n 0.00559242f $X=5.315 $Y=1.725 $X2=0
+ $Y2=0
cc_394 N_B1_c_469_n N_A_49_367#_c_612_n 0.00977976f $X=7.105 $Y=1.725 $X2=0
+ $Y2=0
cc_395 N_B1_c_469_n N_A_49_367#_c_613_n 0.00322972f $X=7.105 $Y=1.725 $X2=0
+ $Y2=0
cc_396 N_B1_c_469_n N_A_49_367#_c_627_n 0.0048058f $X=7.105 $Y=1.725 $X2=0 $Y2=0
cc_397 N_B1_c_466_n N_VPWR_c_758_n 0.00315355f $X=5.315 $Y=1.725 $X2=0 $Y2=0
cc_398 N_B1_c_467_n N_VPWR_c_758_n 0.0019369f $X=6.015 $Y=1.725 $X2=0 $Y2=0
cc_399 N_B1_c_468_n N_VPWR_c_759_n 0.00441134f $X=6.445 $Y=1.725 $X2=0 $Y2=0
cc_400 N_B1_c_469_n N_VPWR_c_759_n 0.0041162f $X=7.105 $Y=1.725 $X2=0 $Y2=0
cc_401 N_B1_c_466_n N_VPWR_c_760_n 0.00357828f $X=5.315 $Y=1.725 $X2=0 $Y2=0
cc_402 N_B1_c_467_n N_VPWR_c_762_n 0.00441213f $X=6.015 $Y=1.725 $X2=0 $Y2=0
cc_403 N_B1_c_468_n N_VPWR_c_762_n 0.00441213f $X=6.445 $Y=1.725 $X2=0 $Y2=0
cc_404 N_B1_c_469_n N_VPWR_c_766_n 0.00359777f $X=7.105 $Y=1.725 $X2=0 $Y2=0
cc_405 N_B1_c_466_n N_VPWR_c_755_n 0.00604193f $X=5.315 $Y=1.725 $X2=0 $Y2=0
cc_406 N_B1_c_467_n N_VPWR_c_755_n 0.00660777f $X=6.015 $Y=1.725 $X2=0 $Y2=0
cc_407 N_B1_c_468_n N_VPWR_c_755_n 0.00665666f $X=6.445 $Y=1.725 $X2=0 $Y2=0
cc_408 N_B1_c_469_n N_VPWR_c_755_n 0.00621299f $X=7.105 $Y=1.725 $X2=0 $Y2=0
cc_409 N_B1_c_466_n N_Y_c_886_n 0.0125241f $X=5.315 $Y=1.725 $X2=0 $Y2=0
cc_410 N_B1_c_467_n N_Y_c_886_n 0.0108153f $X=6.015 $Y=1.725 $X2=0 $Y2=0
cc_411 N_B1_c_468_n N_Y_c_886_n 0.010663f $X=6.445 $Y=1.725 $X2=0 $Y2=0
cc_412 N_B1_c_469_n N_Y_c_886_n 0.0139249f $X=7.105 $Y=1.725 $X2=0 $Y2=0
cc_413 N_B1_c_462_n N_Y_c_886_n 0.0040141f $X=7.045 $Y=1.495 $X2=0 $Y2=0
cc_414 N_B1_M1025_g N_Y_c_872_n 0.0128907f $X=7.045 $Y=0.655 $X2=0 $Y2=0
cc_415 N_B1_c_462_n N_Y_c_872_n 2.41526e-19 $X=7.045 $Y=1.495 $X2=0 $Y2=0
cc_416 N_B1_c_469_n N_Y_c_893_n 0.00300376f $X=7.105 $Y=1.725 $X2=0 $Y2=0
cc_417 N_B1_c_469_n N_Y_c_876_n 2.43046e-19 $X=7.105 $Y=1.725 $X2=0 $Y2=0
cc_418 N_B1_c_462_n N_Y_c_876_n 5.34872e-19 $X=7.045 $Y=1.495 $X2=0 $Y2=0
cc_419 N_B1_M1014_g N_Y_c_924_n 0.0127021f $X=5.815 $Y=0.655 $X2=0 $Y2=0
cc_420 N_B1_M1023_g N_Y_c_924_n 0.0126112f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_421 N_B1_c_478_n N_Y_c_924_n 0.00783301f $X=6.765 $Y=1.43 $X2=0 $Y2=0
cc_422 N_B1_c_462_n N_Y_c_924_n 0.00652786f $X=7.045 $Y=1.495 $X2=0 $Y2=0
cc_423 N_B1_c_463_n N_Y_c_924_n 0.0685395f $X=6.413 $Y=1.362 $X2=0 $Y2=0
cc_424 N_B1_c_464_n N_Y_c_924_n 0.00873366f $X=5.597 $Y=1.362 $X2=0 $Y2=0
cc_425 N_B1_M1023_g N_Y_c_874_n 0.00292787f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_426 N_B1_c_478_n N_Y_c_874_n 0.0137637f $X=6.765 $Y=1.43 $X2=0 $Y2=0
cc_427 N_B1_c_462_n N_Y_c_874_n 0.0036317f $X=7.045 $Y=1.495 $X2=0 $Y2=0
cc_428 N_B1_c_469_n Y 0.00629589f $X=7.105 $Y=1.725 $X2=0 $Y2=0
cc_429 N_B1_M1008_g N_VGND_c_986_n 0.00357877f $X=5.385 $Y=0.655 $X2=0 $Y2=0
cc_430 N_B1_M1014_g N_VGND_c_986_n 0.00357877f $X=5.815 $Y=0.655 $X2=0 $Y2=0
cc_431 N_B1_M1023_g N_VGND_c_986_n 0.00357877f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_432 N_B1_M1025_g N_VGND_c_986_n 0.00359361f $X=7.045 $Y=0.655 $X2=0 $Y2=0
cc_433 N_B1_M1008_g N_VGND_c_990_n 0.00537654f $X=5.385 $Y=0.655 $X2=0 $Y2=0
cc_434 N_B1_M1014_g N_VGND_c_990_n 0.0053512f $X=5.815 $Y=0.655 $X2=0 $Y2=0
cc_435 N_B1_M1023_g N_VGND_c_990_n 0.00609634f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_436 N_B1_M1025_g N_VGND_c_990_n 0.00611257f $X=7.045 $Y=0.655 $X2=0 $Y2=0
cc_437 N_B1_M1008_g N_A_132_47#_c_1095_n 0.00253514f $X=5.385 $Y=0.655 $X2=0
+ $Y2=0
cc_438 N_B1_c_462_n N_A_132_47#_c_1095_n 7.40386e-19 $X=7.045 $Y=1.495 $X2=0
+ $Y2=0
cc_439 N_B1_c_464_n N_A_132_47#_c_1095_n 0.00187112f $X=5.597 $Y=1.362 $X2=0
+ $Y2=0
cc_440 N_B1_M1008_g N_A_132_47#_c_1135_n 0.0149103f $X=5.385 $Y=0.655 $X2=0
+ $Y2=0
cc_441 N_B1_M1014_g N_A_132_47#_c_1135_n 0.0103812f $X=5.815 $Y=0.655 $X2=0
+ $Y2=0
cc_442 N_B1_M1023_g N_A_132_47#_c_1135_n 0.0128053f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_443 N_B1_M1025_g N_A_132_47#_c_1135_n 0.0137488f $X=7.045 $Y=0.655 $X2=0
+ $Y2=0
cc_444 N_B1_c_464_n N_A_132_47#_c_1135_n 6.68218e-19 $X=5.597 $Y=1.362 $X2=0
+ $Y2=0
cc_445 N_B1_M1025_g N_A_132_47#_c_1131_n 0.0107542f $X=7.045 $Y=0.655 $X2=0
+ $Y2=0
cc_446 N_A_49_367#_c_553_n N_A_132_367#_M1012_d 0.00176461f $X=1.145 $Y=1.9
+ $X2=-0.19 $Y2=1.655
cc_447 N_A_49_367#_c_583_n N_A_132_367#_M1009_d 0.00333177f $X=2.005 $Y=2.015
+ $X2=0 $Y2=0
cc_448 N_A_49_367#_c_554_n N_A_132_367#_M1026_d 0.00176461f $X=2.855 $Y=1.9
+ $X2=0 $Y2=0
cc_449 N_A_49_367#_c_555_n N_A_132_367#_M1030_d 0.00180746f $X=3.645 $Y=1.79
+ $X2=0 $Y2=0
cc_450 N_A_49_367#_c_553_n N_A_132_367#_c_708_n 0.00560614f $X=1.145 $Y=1.9
+ $X2=0 $Y2=0
cc_451 N_A_49_367#_c_583_n N_A_132_367#_c_708_n 0.00843866f $X=2.005 $Y=2.015
+ $X2=0 $Y2=0
cc_452 N_A_49_367#_c_558_n N_A_132_367#_c_708_n 0.012604f $X=1.23 $Y=1.9 $X2=0
+ $Y2=0
cc_453 N_A_49_367#_c_583_n N_A_132_367#_c_710_n 0.00843866f $X=2.005 $Y=2.015
+ $X2=0 $Y2=0
cc_454 N_A_49_367#_c_554_n N_A_132_367#_c_710_n 0.00560614f $X=2.855 $Y=1.9
+ $X2=0 $Y2=0
cc_455 N_A_49_367#_c_559_n N_A_132_367#_c_710_n 0.012604f $X=2.09 $Y=1.9 $X2=0
+ $Y2=0
cc_456 N_A_49_367#_M1020_s N_A_132_367#_c_702_n 0.00333487f $X=2.81 $Y=1.835
+ $X2=0 $Y2=0
cc_457 N_A_49_367#_c_560_n N_A_132_367#_c_702_n 0.0127906f $X=2.95 $Y=1.98 $X2=0
+ $Y2=0
cc_458 N_A_49_367#_c_555_n N_A_132_367#_c_733_n 0.0129403f $X=3.645 $Y=1.79
+ $X2=0 $Y2=0
cc_459 N_A_49_367#_c_553_n N_A_132_367#_c_704_n 0.0170777f $X=1.145 $Y=1.9 $X2=0
+ $Y2=0
cc_460 N_A_49_367#_c_583_n N_A_132_367#_c_715_n 0.01723f $X=2.005 $Y=2.015 $X2=0
+ $Y2=0
cc_461 N_A_49_367#_c_554_n N_A_132_367#_c_705_n 0.0170777f $X=2.855 $Y=1.9 $X2=0
+ $Y2=0
cc_462 N_A_49_367#_c_558_n N_VPWR_M1001_s 0.0017933f $X=1.23 $Y=1.9 $X2=-0.19
+ $Y2=1.655
cc_463 N_A_49_367#_c_559_n N_VPWR_M1013_s 0.0017933f $X=2.09 $Y=1.9 $X2=0 $Y2=0
cc_464 N_A_49_367#_c_610_n N_VPWR_M1000_d 0.00248565f $X=5.355 $Y=2.985 $X2=0
+ $Y2=0
cc_465 N_A_49_367#_c_611_n N_VPWR_M1000_d 0.00373691f $X=5.44 $Y=2.895 $X2=0
+ $Y2=0
cc_466 N_A_49_367#_c_621_n N_VPWR_M1000_d 0.0106007f $X=6.995 $Y=2.495 $X2=0
+ $Y2=0
cc_467 N_A_49_367#_c_624_n N_VPWR_M1000_d 8.30889e-19 $X=5.525 $Y=2.495 $X2=0
+ $Y2=0
cc_468 N_A_49_367#_c_621_n N_VPWR_M1003_d 0.0108514f $X=6.995 $Y=2.495 $X2=0
+ $Y2=0
cc_469 N_A_49_367#_c_610_n N_VPWR_c_758_n 0.0148558f $X=5.355 $Y=2.985 $X2=0
+ $Y2=0
cc_470 N_A_49_367#_c_611_n N_VPWR_c_758_n 0.0106649f $X=5.44 $Y=2.895 $X2=0
+ $Y2=0
cc_471 N_A_49_367#_c_621_n N_VPWR_c_758_n 0.0147195f $X=6.995 $Y=2.495 $X2=0
+ $Y2=0
cc_472 N_A_49_367#_c_621_n N_VPWR_c_759_n 0.0194424f $X=6.995 $Y=2.495 $X2=0
+ $Y2=0
cc_473 N_A_49_367#_c_574_n N_VPWR_c_760_n 0.0189946f $X=3.81 $Y=2.905 $X2=0
+ $Y2=0
cc_474 N_A_49_367#_c_605_n N_VPWR_c_760_n 0.0298674f $X=4.505 $Y=2.99 $X2=0
+ $Y2=0
cc_475 N_A_49_367#_c_610_n N_VPWR_c_760_n 0.0392276f $X=5.355 $Y=2.985 $X2=0
+ $Y2=0
cc_476 N_A_49_367#_c_621_n N_VPWR_c_760_n 0.00232298f $X=6.995 $Y=2.495 $X2=0
+ $Y2=0
cc_477 N_A_49_367#_c_615_n N_VPWR_c_760_n 0.0190758f $X=4.67 $Y=2.985 $X2=0
+ $Y2=0
cc_478 N_A_49_367#_c_621_n N_VPWR_c_762_n 0.00740781f $X=6.995 $Y=2.495 $X2=0
+ $Y2=0
cc_479 N_A_49_367#_c_552_n N_VPWR_c_764_n 0.0178111f $X=0.37 $Y=2.91 $X2=0 $Y2=0
cc_480 N_A_49_367#_c_621_n N_VPWR_c_766_n 0.00218717f $X=6.995 $Y=2.495 $X2=0
+ $Y2=0
cc_481 N_A_49_367#_c_613_n N_VPWR_c_766_n 0.0329772f $X=7.8 $Y=2.98 $X2=0 $Y2=0
cc_482 N_A_49_367#_c_627_n N_VPWR_c_766_n 0.00978398f $X=7.165 $Y=2.98 $X2=0
+ $Y2=0
cc_483 N_A_49_367#_c_556_n N_VPWR_c_766_n 0.0172312f $X=7.93 $Y=2.895 $X2=0
+ $Y2=0
cc_484 N_A_49_367#_M1012_s N_VPWR_c_755_n 0.00371702f $X=0.245 $Y=1.835 $X2=0
+ $Y2=0
cc_485 N_A_49_367#_M1020_s N_VPWR_c_755_n 0.00225186f $X=2.81 $Y=1.835 $X2=0
+ $Y2=0
cc_486 N_A_49_367#_M1031_s N_VPWR_c_755_n 0.00223559f $X=3.67 $Y=1.835 $X2=0
+ $Y2=0
cc_487 N_A_49_367#_M1015_s N_VPWR_c_755_n 0.00223559f $X=4.53 $Y=1.835 $X2=0
+ $Y2=0
cc_488 N_A_49_367#_M1028_s N_VPWR_c_755_n 0.0025316f $X=7.71 $Y=1.835 $X2=0
+ $Y2=0
cc_489 N_A_49_367#_c_552_n N_VPWR_c_755_n 0.0100304f $X=0.37 $Y=2.91 $X2=0 $Y2=0
cc_490 N_A_49_367#_c_574_n N_VPWR_c_755_n 0.0124451f $X=3.81 $Y=2.905 $X2=0
+ $Y2=0
cc_491 N_A_49_367#_c_605_n N_VPWR_c_755_n 0.0187823f $X=4.505 $Y=2.99 $X2=0
+ $Y2=0
cc_492 N_A_49_367#_c_610_n N_VPWR_c_755_n 0.0249202f $X=5.355 $Y=2.985 $X2=0
+ $Y2=0
cc_493 N_A_49_367#_c_621_n N_VPWR_c_755_n 0.0261479f $X=6.995 $Y=2.495 $X2=0
+ $Y2=0
cc_494 N_A_49_367#_c_613_n N_VPWR_c_755_n 0.0228986f $X=7.8 $Y=2.98 $X2=0 $Y2=0
cc_495 N_A_49_367#_c_627_n N_VPWR_c_755_n 0.00594933f $X=7.165 $Y=2.98 $X2=0
+ $Y2=0
cc_496 N_A_49_367#_c_556_n N_VPWR_c_755_n 0.0100602f $X=7.93 $Y=2.895 $X2=0
+ $Y2=0
cc_497 N_A_49_367#_c_615_n N_VPWR_c_755_n 0.0124594f $X=4.67 $Y=2.985 $X2=0
+ $Y2=0
cc_498 N_A_49_367#_c_605_n N_Y_M1006_d 0.00332344f $X=4.505 $Y=2.99 $X2=0 $Y2=0
cc_499 N_A_49_367#_c_610_n N_Y_M1018_d 0.00332931f $X=5.355 $Y=2.985 $X2=0 $Y2=0
cc_500 N_A_49_367#_c_621_n N_Y_M1002_s 0.00495692f $X=6.995 $Y=2.495 $X2=0 $Y2=0
cc_501 N_A_49_367#_c_613_n N_Y_M1021_s 0.00660142f $X=7.8 $Y=2.98 $X2=0 $Y2=0
cc_502 N_A_49_367#_M1015_s N_Y_c_882_n 0.003357f $X=4.53 $Y=1.835 $X2=0 $Y2=0
cc_503 N_A_49_367#_c_607_n N_Y_c_882_n 0.0171647f $X=4.67 $Y=2.47 $X2=0 $Y2=0
cc_504 N_A_49_367#_c_610_n N_Y_c_886_n 0.00255653f $X=5.355 $Y=2.985 $X2=0 $Y2=0
cc_505 N_A_49_367#_c_621_n N_Y_c_886_n 0.0986844f $X=6.995 $Y=2.495 $X2=0 $Y2=0
cc_506 N_A_49_367#_c_624_n N_Y_c_886_n 0.00911135f $X=5.525 $Y=2.495 $X2=0 $Y2=0
cc_507 N_A_49_367#_c_613_n N_Y_c_886_n 0.00292862f $X=7.8 $Y=2.98 $X2=0 $Y2=0
cc_508 N_A_49_367#_M1028_s N_Y_c_875_n 0.00395918f $X=7.71 $Y=1.835 $X2=0 $Y2=0
cc_509 N_A_49_367#_c_557_n N_Y_c_875_n 0.0225797f $X=7.895 $Y=2.21 $X2=0 $Y2=0
cc_510 N_A_49_367#_c_605_n N_Y_c_907_n 0.0126631f $X=4.505 $Y=2.99 $X2=0 $Y2=0
cc_511 N_A_49_367#_c_610_n N_Y_c_909_n 0.0127285f $X=5.355 $Y=2.985 $X2=0 $Y2=0
cc_512 N_A_49_367#_c_557_n N_Y_c_910_n 0.0157939f $X=7.895 $Y=2.21 $X2=0 $Y2=0
cc_513 N_A_49_367#_c_621_n Y 0.0138951f $X=6.995 $Y=2.495 $X2=0 $Y2=0
cc_514 N_A_49_367#_c_612_n Y 0.00986538f $X=7.08 $Y=2.895 $X2=0 $Y2=0
cc_515 N_A_49_367#_c_613_n Y 0.0167688f $X=7.8 $Y=2.98 $X2=0 $Y2=0
cc_516 N_A_49_367#_c_557_n Y 0.0358652f $X=7.895 $Y=2.21 $X2=0 $Y2=0
cc_517 N_A_49_367#_c_555_n N_A_132_47#_c_1094_n 0.00541068f $X=3.645 $Y=1.79
+ $X2=0 $Y2=0
cc_518 N_A_132_367#_c_708_n N_VPWR_M1001_s 0.00343709f $X=1.495 $Y=2.355
+ $X2=0.585 $Y2=1.185
cc_519 N_A_132_367#_c_710_n N_VPWR_M1013_s 0.00343709f $X=2.355 $Y=2.355
+ $X2=0.585 $Y2=0.655
cc_520 N_A_132_367#_c_708_n N_VPWR_c_756_n 0.0135055f $X=1.495 $Y=2.355 $X2=0
+ $Y2=0
cc_521 N_A_132_367#_c_710_n N_VPWR_c_757_n 0.0135055f $X=2.355 $Y=2.355 $X2=0
+ $Y2=0
cc_522 N_A_132_367#_c_701_n N_VPWR_c_760_n 0.01906f $X=2.52 $Y=2.885 $X2=3.595
+ $Y2=2.465
cc_523 N_A_132_367#_c_702_n N_VPWR_c_760_n 0.0317835f $X=3.245 $Y=2.98 $X2=3.595
+ $Y2=2.465
cc_524 N_A_132_367#_c_743_p N_VPWR_c_760_n 0.0139427f $X=3.36 $Y=2.885 $X2=3.595
+ $Y2=2.465
cc_525 N_A_132_367#_c_700_n N_VPWR_c_764_n 0.0189236f $X=0.8 $Y=2.95 $X2=3.505
+ $Y2=1.42
cc_526 N_A_132_367#_c_715_n N_VPWR_c_765_n 0.0189236f $X=1.66 $Y=2.435 $X2=0.495
+ $Y2=1.35
cc_527 N_A_132_367#_M1012_d N_VPWR_c_755_n 0.00223559f $X=0.66 $Y=1.835 $X2=2.64
+ $Y2=1.29
cc_528 N_A_132_367#_M1009_d N_VPWR_c_755_n 0.00223559f $X=1.52 $Y=1.835 $X2=2.64
+ $Y2=1.29
cc_529 N_A_132_367#_M1026_d N_VPWR_c_755_n 0.00223559f $X=2.38 $Y=1.835 $X2=2.64
+ $Y2=1.29
cc_530 N_A_132_367#_M1030_d N_VPWR_c_755_n 0.00373407f $X=3.24 $Y=1.835 $X2=2.64
+ $Y2=1.29
cc_531 N_A_132_367#_c_700_n N_VPWR_c_755_n 0.0123859f $X=0.8 $Y=2.95 $X2=2.64
+ $Y2=1.29
cc_532 N_A_132_367#_c_701_n N_VPWR_c_755_n 0.0124545f $X=2.52 $Y=2.885 $X2=2.64
+ $Y2=1.29
cc_533 N_A_132_367#_c_702_n N_VPWR_c_755_n 0.019774f $X=3.245 $Y=2.98 $X2=2.64
+ $Y2=1.29
cc_534 N_A_132_367#_c_743_p N_VPWR_c_755_n 0.00893659f $X=3.36 $Y=2.885 $X2=2.64
+ $Y2=1.29
cc_535 N_A_132_367#_c_715_n N_VPWR_c_755_n 0.0123859f $X=1.66 $Y=2.435 $X2=2.64
+ $Y2=1.29
cc_536 N_VPWR_c_755_n N_Y_M1006_d 0.00225186f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_537 N_VPWR_c_755_n N_Y_M1018_d 0.00225186f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_538 N_VPWR_c_755_n N_Y_M1002_s 0.00373122f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_539 N_VPWR_c_755_n N_Y_M1021_s 0.00305989f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_540 N_VPWR_M1000_d N_Y_c_886_n 0.0107998f $X=5.39 $Y=1.835 $X2=0 $Y2=0
cc_541 N_VPWR_M1003_d N_Y_c_886_n 0.0095684f $X=6.52 $Y=1.835 $X2=0 $Y2=0
cc_542 N_Y_c_872_n N_VGND_M1022_s 0.00377044f $X=7.89 $Y=1.08 $X2=0 $Y2=0
cc_543 N_Y_c_872_n N_VGND_c_979_n 0.027093f $X=7.89 $Y=1.08 $X2=0 $Y2=0
cc_544 N_Y_M1008_s N_VGND_c_990_n 0.00225186f $X=5.46 $Y=0.235 $X2=0 $Y2=0
cc_545 N_Y_M1023_s N_VGND_c_990_n 0.00532502f $X=6.32 $Y=0.235 $X2=0 $Y2=0
cc_546 N_Y_c_924_n N_A_132_47#_M1014_d 0.00334677f $X=6.745 $Y=0.932 $X2=0 $Y2=0
cc_547 N_Y_c_872_n N_A_132_47#_M1025_d 0.00176461f $X=7.89 $Y=1.08 $X2=0 $Y2=0
cc_548 N_Y_M1008_s N_A_132_47#_c_1135_n 0.00337742f $X=5.46 $Y=0.235 $X2=0 $Y2=0
cc_549 N_Y_M1023_s N_A_132_47#_c_1135_n 0.0152875f $X=6.32 $Y=0.235 $X2=0 $Y2=0
cc_550 N_Y_c_872_n N_A_132_47#_c_1135_n 0.00387227f $X=7.89 $Y=1.08 $X2=0 $Y2=0
cc_551 N_Y_c_924_n N_A_132_47#_c_1135_n 0.0872087f $X=6.745 $Y=0.932 $X2=0 $Y2=0
cc_552 N_Y_c_872_n N_A_132_47#_c_1131_n 0.0168339f $X=7.89 $Y=1.08 $X2=0 $Y2=0
cc_553 N_VGND_c_990_n N_A_132_47#_M1004_s 0.00245017f $X=7.92 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_554 N_VGND_c_990_n N_A_132_47#_M1016_s 0.00266476f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_555 N_VGND_c_990_n N_A_132_47#_M1029_s 0.00266476f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_556 N_VGND_c_990_n N_A_132_47#_M1011_s 0.00400238f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_557 N_VGND_c_990_n N_A_132_47#_M1005_d 0.00440023f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_558 N_VGND_c_990_n N_A_132_47#_M1019_d 0.00341839f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_559 N_VGND_c_990_n N_A_132_47#_M1014_d 0.00223577f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_560 N_VGND_c_990_n N_A_132_47#_M1025_d 0.00223559f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_561 N_VGND_c_984_n N_A_132_47#_c_1101_n 0.0156443f $X=1.065 $Y=0 $X2=0 $Y2=0
cc_562 N_VGND_c_990_n N_A_132_47#_c_1101_n 0.00983564f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_563 N_VGND_M1010_d N_A_132_47#_c_1102_n 0.00335437f $X=1.09 $Y=0.235 $X2=0
+ $Y2=0
cc_564 N_VGND_c_972_n N_A_132_47#_c_1102_n 0.016459f $X=1.23 $Y=0.44 $X2=0 $Y2=0
cc_565 N_VGND_c_984_n N_A_132_47#_c_1102_n 0.00196209f $X=1.065 $Y=0 $X2=0 $Y2=0
cc_566 N_VGND_c_985_n N_A_132_47#_c_1102_n 0.00196209f $X=1.925 $Y=0 $X2=0 $Y2=0
cc_567 N_VGND_c_990_n N_A_132_47#_c_1102_n 0.00891615f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_568 N_VGND_c_985_n N_A_132_47#_c_1164_n 0.0124139f $X=1.925 $Y=0 $X2=0 $Y2=0
cc_569 N_VGND_c_990_n N_A_132_47#_c_1164_n 0.00730033f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_570 N_VGND_M1027_d N_A_132_47#_c_1103_n 0.00335437f $X=1.95 $Y=0.235 $X2=0
+ $Y2=0
cc_571 N_VGND_c_973_n N_A_132_47#_c_1103_n 0.016459f $X=2.09 $Y=0.44 $X2=0 $Y2=0
cc_572 N_VGND_c_980_n N_A_132_47#_c_1103_n 0.00196209f $X=2.785 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_c_985_n N_A_132_47#_c_1103_n 0.00196209f $X=1.925 $Y=0 $X2=0 $Y2=0
cc_574 N_VGND_c_990_n N_A_132_47#_c_1103_n 0.00891615f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_575 N_VGND_c_980_n N_A_132_47#_c_1171_n 0.0124139f $X=2.785 $Y=0 $X2=0 $Y2=0
cc_576 N_VGND_c_990_n N_A_132_47#_c_1171_n 0.00730033f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_577 N_VGND_M1007_d N_A_132_47#_c_1104_n 0.0035786f $X=2.81 $Y=0.235 $X2=0
+ $Y2=0
cc_578 N_VGND_c_974_n N_A_132_47#_c_1104_n 0.016459f $X=2.95 $Y=0.44 $X2=0 $Y2=0
cc_579 N_VGND_c_980_n N_A_132_47#_c_1104_n 0.00196209f $X=2.785 $Y=0 $X2=0 $Y2=0
cc_580 N_VGND_c_982_n N_A_132_47#_c_1104_n 0.00188649f $X=3.645 $Y=0 $X2=0 $Y2=0
cc_581 N_VGND_c_990_n N_A_132_47#_c_1104_n 0.00865724f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_582 N_VGND_c_982_n N_A_132_47#_c_1178_n 0.0124525f $X=3.645 $Y=0 $X2=0 $Y2=0
cc_583 N_VGND_c_990_n N_A_132_47#_c_1178_n 0.00730901f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_584 N_VGND_M1024_d N_A_132_47#_c_1094_n 0.00180746f $X=3.67 $Y=0.235 $X2=0
+ $Y2=0
cc_585 N_VGND_c_975_n N_A_132_47#_c_1094_n 0.0163515f $X=3.81 $Y=0.36 $X2=0
+ $Y2=0
cc_586 N_VGND_c_976_n N_A_132_47#_c_1182_n 0.00651381f $X=4.55 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_990_n N_A_132_47#_c_1182_n 0.00784653f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_M1017_s N_A_132_47#_c_1095_n 0.00256964f $X=4.53 $Y=0.235 $X2=0
+ $Y2=0
cc_589 N_VGND_c_977_n N_A_132_47#_c_1095_n 0.018397f $X=4.715 $Y=0.36 $X2=0
+ $Y2=0
cc_590 N_VGND_c_986_n N_A_132_47#_c_1186_n 0.0128782f $X=7.605 $Y=0 $X2=0 $Y2=0
cc_591 N_VGND_c_990_n N_A_132_47#_c_1186_n 0.00777554f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_592 N_VGND_c_986_n N_A_132_47#_c_1135_n 0.10693f $X=7.605 $Y=0 $X2=0 $Y2=0
cc_593 N_VGND_c_990_n N_A_132_47#_c_1135_n 0.0666928f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_c_990_n N_A_132_47#_c_1096_n 2.41233e-19 $X=7.92 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_c_986_n N_A_132_47#_c_1131_n 0.0187344f $X=7.605 $Y=0 $X2=0 $Y2=0
cc_596 N_VGND_c_990_n N_A_132_47#_c_1131_n 0.0123282f $X=7.92 $Y=0 $X2=0 $Y2=0
