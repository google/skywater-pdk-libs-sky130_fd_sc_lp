* File: sky130_fd_sc_lp__o32a_0.pex.spice
* Created: Fri Aug 28 11:17:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32A_0%A_97_309# 1 2 9 13 17 18 21 22 24 25 28 30 33
+ 34 36
r81 36 37 4.11508 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0.725
+ $X2=3.16 $Y2=0.725
r82 32 37 2.39319 $w=1.9e-07 $l=1.3e-07 $layer=LI1_cond $X=3.16 $Y=0.855
+ $X2=3.16 $Y2=0.725
r83 32 33 68.2967 $w=1.88e-07 $l=1.17e-06 $layer=LI1_cond $X=3.16 $Y=0.855
+ $X2=3.16 $Y2=2.025
r84 31 34 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=2.12
+ $X2=2.475 $Y2=2.12
r85 30 33 6.81649 $w=1.9e-07 $l=1.3435e-07 $layer=LI1_cond $X=3.065 $Y=2.12
+ $X2=3.16 $Y2=2.025
r86 30 31 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=3.065 $Y=2.12
+ $X2=2.64 $Y2=2.12
r87 26 34 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.475 $Y=2.215
+ $X2=2.475 $Y2=2.12
r88 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.475 $Y=2.215
+ $X2=2.475 $Y2=2.55
r89 24 34 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=2.12
+ $X2=2.475 $Y2=2.12
r90 24 25 87.2679 $w=1.88e-07 $l=1.495e-06 $layer=LI1_cond $X=2.31 $Y=2.12
+ $X2=0.815 $Y2=2.12
r91 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.65
+ $Y=1.71 $X2=0.65 $Y2=1.71
r92 19 25 7.03324 $w=1.9e-07 $l=1.71026e-07 $layer=LI1_cond $X=0.685 $Y=2.025
+ $X2=0.815 $Y2=2.12
r93 19 21 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.685 $Y=2.025
+ $X2=0.685 $Y2=1.71
r94 17 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.65 $Y=2.05
+ $X2=0.65 $Y2=1.71
r95 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=2.05
+ $X2=0.65 $Y2=2.215
r96 16 22 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=1.545
+ $X2=0.65 $Y2=1.71
r97 13 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.74 $Y=2.725
+ $X2=0.74 $Y2=2.215
r98 9 16 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=0.71 $Y=0.635
+ $X2=0.71 $Y2=1.545
r99 2 28 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=2.285
+ $Y=2.405 $X2=2.465 $Y2=2.55
r100 1 36 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.425 $X2=3.075 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_0%A1 3 6 9 13 14 17 19 20 21 26
c53 17 0 1.55717e-19 $X=1.43 $Y=2.17
r54 20 21 16.1342 $w=2.98e-07 $l=4.2e-07 $layer=LI1_cond $X=1.135 $Y=1.245
+ $X2=1.135 $Y2=1.665
r55 20 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.19
+ $Y=1.245 $X2=1.19 $Y2=1.245
r56 19 20 12.2927 $w=2.98e-07 $l=3.2e-07 $layer=LI1_cond $X=1.135 $Y=0.925
+ $X2=1.135 $Y2=1.245
r57 15 17 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.28 $Y=2.17
+ $X2=1.43 $Y2=2.17
r58 13 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.19 $Y=1.585
+ $X2=1.19 $Y2=1.245
r59 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.585
+ $X2=1.19 $Y2=1.75
r60 12 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.08
+ $X2=1.19 $Y2=1.245
r61 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.43 $Y=2.245
+ $X2=1.43 $Y2=2.17
r62 7 9 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.43 $Y=2.245 $X2=1.43
+ $Y2=2.725
r63 6 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.28 $Y=2.095
+ $X2=1.28 $Y2=2.17
r64 6 14 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.28 $Y=2.095
+ $X2=1.28 $Y2=1.75
r65 3 12 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.28 $Y=0.635
+ $X2=1.28 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_0%A2 3 7 11 12 13 14 18
c43 13 0 1.55717e-19 $X=1.68 $Y=1.295
r44 13 14 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.662 $Y=1.295
+ $X2=1.662 $Y2=1.665
r45 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.73
+ $Y=1.35 $X2=1.73 $Y2=1.35
r46 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.73 $Y=1.69
+ $X2=1.73 $Y2=1.35
r47 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.69
+ $X2=1.73 $Y2=1.855
r48 10 18 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.185
+ $X2=1.73 $Y2=1.35
r49 7 12 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.82 $Y=2.725
+ $X2=1.82 $Y2=1.855
r50 3 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.71 $Y=0.635
+ $X2=1.71 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_0%A3 3 7 11 12 13 14 18
r41 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.27
+ $Y=1.35 $X2=2.27 $Y2=1.35
r42 14 19 10.677 $w=3.38e-07 $l=3.15e-07 $layer=LI1_cond $X=2.185 $Y=1.665
+ $X2=2.185 $Y2=1.35
r43 13 19 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=2.185 $Y=1.295
+ $X2=2.185 $Y2=1.35
r44 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.27 $Y=1.69
+ $X2=2.27 $Y2=1.35
r45 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.69
+ $X2=2.27 $Y2=1.855
r46 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.185
+ $X2=2.27 $Y2=1.35
r47 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.36 $Y=0.635
+ $X2=2.36 $Y2=1.185
r48 3 12 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=2.21 $Y=2.725
+ $X2=2.21 $Y2=1.855
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_0%B2 3 7 11 12 13 14 18
r41 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.81
+ $Y=1.35 $X2=2.81 $Y2=1.35
r42 14 19 9.81134 $w=3.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.71 $Y=1.665
+ $X2=2.71 $Y2=1.35
r43 13 19 1.71309 $w=3.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.71 $Y=1.295
+ $X2=2.71 $Y2=1.35
r44 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.81 $Y=1.69
+ $X2=2.81 $Y2=1.35
r45 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.69
+ $X2=2.81 $Y2=1.855
r46 10 18 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.185
+ $X2=2.81 $Y2=1.35
r47 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.79 $Y=0.635
+ $X2=2.79 $Y2=1.185
r48 3 12 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=2.72 $Y=2.725
+ $X2=2.72 $Y2=1.855
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_0%B1 3 7 9 12 14 15 16 21 22 23
r32 21 24 88.3231 $w=4.6e-07 $l=5.05e-07 $layer=POLY_cond $X=3.445 $Y=1.12
+ $X2=3.445 $Y2=1.625
r33 21 23 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.445 $Y=1.12
+ $X2=3.445 $Y2=0.955
r34 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.51
+ $Y=1.12 $X2=3.51 $Y2=1.12
r35 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.59 $Y=1.665
+ $X2=3.59 $Y2=2.035
r36 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.59 $Y=1.295
+ $X2=3.59 $Y2=1.665
r37 14 22 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=3.59 $Y=1.295
+ $X2=3.59 $Y2=1.12
r38 10 12 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.11 $Y=2.17
+ $X2=3.29 $Y2=2.17
r39 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.29 $Y=2.095
+ $X2=3.29 $Y2=2.17
r40 9 24 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.29 $Y=2.095 $X2=3.29
+ $Y2=1.625
r41 7 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.29 $Y=0.635
+ $X2=3.29 $Y2=0.955
r42 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.11 $Y=2.245
+ $X2=3.11 $Y2=2.17
r43 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.11 $Y=2.245 $X2=3.11
+ $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_0%X 1 2 7 8 9 10 11 12 13 38 41
r19 41 42 3.23806 $w=6.03e-07 $l=1e-08 $layer=LI1_cond $X=0.387 $Y=2.405
+ $X2=0.387 $Y2=2.395
r20 22 33 1.29116 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.235 $Y=0.8 $X2=0.235
+ $Y2=0.635
r21 13 45 4.25053 $w=6.03e-07 $l=2.15e-07 $layer=LI1_cond $X=0.387 $Y=2.775
+ $X2=0.387 $Y2=2.56
r22 12 45 2.33285 $w=6.03e-07 $l=1.18e-07 $layer=LI1_cond $X=0.387 $Y=2.442
+ $X2=0.387 $Y2=2.56
r23 12 41 0.731486 $w=6.03e-07 $l=3.7e-08 $layer=LI1_cond $X=0.387 $Y=2.442
+ $X2=0.387 $Y2=2.405
r24 12 42 1.45976 $w=2.98e-07 $l=3.8e-08 $layer=LI1_cond $X=0.235 $Y=2.357
+ $X2=0.235 $Y2=2.395
r25 11 12 12.3696 $w=2.98e-07 $l=3.22e-07 $layer=LI1_cond $X=0.235 $Y=2.035
+ $X2=0.235 $Y2=2.357
r26 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.665
+ $X2=0.235 $Y2=2.035
r27 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.665
r28 8 9 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=0.925
+ $X2=0.235 $Y2=1.295
r29 8 22 4.80185 $w=2.98e-07 $l=1.25e-07 $layer=LI1_cond $X=0.235 $Y=0.925
+ $X2=0.235 $Y2=0.8
r30 7 38 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.24 $Y=0.635
+ $X2=0.495 $Y2=0.635
r31 7 33 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.24 $Y=0.635
+ $X2=0.235 $Y2=0.635
r32 2 45 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.4
+ $Y=2.405 $X2=0.525 $Y2=2.56
r33 1 38 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.37
+ $Y=0.425 $X2=0.495 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_0%VPWR 1 2 9 13 16 17 18 20 30 31 34
r37 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r38 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r39 28 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r40 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.085 $Y2=3.33
r42 25 27 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=1.25 $Y=3.33 $X2=3.12
+ $Y2=3.33
r43 23 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 20 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=3.33
+ $X2=1.085 $Y2=3.33
r46 20 22 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.92 $Y=3.33 $X2=0.72
+ $Y2=3.33
r47 18 28 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 18 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 16 27 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r50 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=3.33
+ $X2=3.325 $Y2=3.33
r51 15 30 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.49 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.49 $Y=3.33
+ $X2=3.325 $Y2=3.33
r53 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=3.245
+ $X2=3.325 $Y2=3.33
r54 11 13 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=3.325 $Y=3.245
+ $X2=3.325 $Y2=2.56
r55 7 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=3.245
+ $X2=1.085 $Y2=3.33
r56 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.085 $Y=3.245
+ $X2=1.085 $Y2=2.55
r57 2 13 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=3.185
+ $Y=2.405 $X2=3.325 $Y2=2.56
r58 1 9 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=0.815
+ $Y=2.405 $X2=1.085 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_0%VGND 1 2 9 13 16 17 18 24 30 31 34
r41 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 31 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r43 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.2 $Y=0 $X2=2.035
+ $Y2=0
r45 28 30 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.2 $Y=0 $X2=3.6
+ $Y2=0
r46 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=2.035
+ $Y2=0
r48 24 26 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.68
+ $Y2=0
r49 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r50 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r51 18 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r52 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r53 16 21 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.72
+ $Y2=0
r54 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.995
+ $Y2=0
r55 15 26 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.68
+ $Y2=0
r56 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=0.995
+ $Y2=0
r57 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=0.085
+ $X2=2.035 $Y2=0
r58 11 13 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.035 $Y=0.085
+ $X2=2.035 $Y2=0.565
r59 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.995 $Y=0.085
+ $X2=0.995 $Y2=0
r60 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.995 $Y=0.085
+ $X2=0.995 $Y2=0.55
r61 2 13 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.785
+ $Y=0.425 $X2=2.035 $Y2=0.565
r62 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.785
+ $Y=0.425 $X2=0.995 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_0%A_271_85# 1 2 3 11 12 13 17 18 19 22 27
r50 25 27 2.70925 $w=2.83e-07 $l=6.7e-08 $layer=LI1_cond $X=1.495 $Y=0.527
+ $X2=1.562 $Y2=0.527
r51 20 22 8.8128 $w=2.53e-07 $l=1.95e-07 $layer=LI1_cond $X=3.542 $Y=0.425
+ $X2=3.542 $Y2=0.62
r52 18 20 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=3.415 $Y=0.34
+ $X2=3.542 $Y2=0.425
r53 18 19 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.415 $Y=0.34
+ $X2=2.68 $Y2=0.34
r54 15 17 8.96345 $w=2.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.545 $Y=0.845
+ $X2=2.545 $Y2=0.635
r55 14 19 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.545 $Y=0.425
+ $X2=2.68 $Y2=0.34
r56 14 17 8.96345 $w=2.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.545 $Y=0.425
+ $X2=2.545 $Y2=0.635
r57 12 15 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.41 $Y=0.93
+ $X2=2.545 $Y2=0.845
r58 12 13 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.41 $Y=0.93
+ $X2=1.66 $Y2=0.93
r59 11 13 6.85817 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=1.562 $Y=0.845
+ $X2=1.66 $Y2=0.93
r60 10 27 2.9806 $w=1.95e-07 $l=1.43e-07 $layer=LI1_cond $X=1.562 $Y=0.67
+ $X2=1.562 $Y2=0.527
r61 10 11 9.95338 $w=1.93e-07 $l=1.75e-07 $layer=LI1_cond $X=1.562 $Y=0.67
+ $X2=1.562 $Y2=0.845
r62 3 22 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.425 $X2=3.505 $Y2=0.62
r63 2 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.425 $X2=2.575 $Y2=0.635
r64 1 25 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.355
+ $Y=0.425 $X2=1.495 $Y2=0.55
.ends

