* File: sky130_fd_sc_lp__o221a_m.pxi.spice
* Created: Wed Sep  2 10:18:45 2020
* 
x_PM_SKY130_FD_SC_LP__O221A_M%C1 N_C1_c_82_n N_C1_M1001_g N_C1_c_88_n
+ N_C1_M1010_g N_C1_c_84_n N_C1_c_89_n C1 C1 N_C1_c_86_n
+ PM_SKY130_FD_SC_LP__O221A_M%C1
x_PM_SKY130_FD_SC_LP__O221A_M%B1 N_B1_c_128_n N_B1_M1009_g N_B1_M1003_g
+ N_B1_c_125_n N_B1_c_126_n N_B1_c_130_n B1 N_B1_c_132_n N_B1_c_127_n
+ PM_SKY130_FD_SC_LP__O221A_M%B1
x_PM_SKY130_FD_SC_LP__O221A_M%B2 N_B2_M1011_g N_B2_M1005_g N_B2_c_184_n
+ N_B2_c_185_n B2 N_B2_c_188_n N_B2_c_189_n N_B2_c_186_n
+ PM_SKY130_FD_SC_LP__O221A_M%B2
x_PM_SKY130_FD_SC_LP__O221A_M%A2 N_A2_M1008_g N_A2_M1007_g N_A2_c_228_n
+ N_A2_c_233_n N_A2_c_234_n N_A2_c_229_n N_A2_c_230_n A2 A2 N_A2_c_235_n
+ N_A2_c_236_n PM_SKY130_FD_SC_LP__O221A_M%A2
x_PM_SKY130_FD_SC_LP__O221A_M%A1 N_A1_M1004_g N_A1_M1000_g N_A1_c_279_n
+ N_A1_c_280_n A1 A1 N_A1_c_281_n N_A1_c_282_n PM_SKY130_FD_SC_LP__O221A_M%A1
x_PM_SKY130_FD_SC_LP__O221A_M%A_27_179# N_A_27_179#_M1001_s N_A_27_179#_M1010_s
+ N_A_27_179#_M1011_d N_A_27_179#_M1002_g N_A_27_179#_M1006_g
+ N_A_27_179#_c_329_n N_A_27_179#_c_330_n N_A_27_179#_c_331_n
+ N_A_27_179#_c_335_n N_A_27_179#_c_368_n N_A_27_179#_c_336_n
+ N_A_27_179#_c_337_n N_A_27_179#_c_338_n N_A_27_179#_c_339_n
+ N_A_27_179#_c_340_n N_A_27_179#_c_341_n N_A_27_179#_c_332_n
+ PM_SKY130_FD_SC_LP__O221A_M%A_27_179#
x_PM_SKY130_FD_SC_LP__O221A_M%VPWR N_VPWR_M1010_d N_VPWR_M1004_d N_VPWR_c_436_n
+ N_VPWR_c_437_n VPWR N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_435_n
+ N_VPWR_c_441_n N_VPWR_c_442_n PM_SKY130_FD_SC_LP__O221A_M%VPWR
x_PM_SKY130_FD_SC_LP__O221A_M%X N_X_M1006_d N_X_M1002_d N_X_c_488_n N_X_c_489_n
+ X X X X X PM_SKY130_FD_SC_LP__O221A_M%X
x_PM_SKY130_FD_SC_LP__O221A_M%A_110_179# N_A_110_179#_M1001_d
+ N_A_110_179#_M1005_d N_A_110_179#_c_516_n N_A_110_179#_c_514_n
+ N_A_110_179#_c_515_n N_A_110_179#_c_534_n
+ PM_SKY130_FD_SC_LP__O221A_M%A_110_179#
x_PM_SKY130_FD_SC_LP__O221A_M%A_196_179# N_A_196_179#_M1009_d
+ N_A_196_179#_M1007_d N_A_196_179#_c_543_n N_A_196_179#_c_554_n
+ N_A_196_179#_c_544_n PM_SKY130_FD_SC_LP__O221A_M%A_196_179#
x_PM_SKY130_FD_SC_LP__O221A_M%VGND N_VGND_M1007_s N_VGND_M1000_d N_VGND_c_574_n
+ N_VGND_c_575_n N_VGND_c_576_n VGND N_VGND_c_577_n N_VGND_c_578_n
+ N_VGND_c_579_n N_VGND_c_580_n N_VGND_c_581_n PM_SKY130_FD_SC_LP__O221A_M%VGND
cc_1 VNB N_C1_c_82_n 0.00217846f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.415
cc_2 VNB N_C1_M1001_g 0.0224065f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.105
cc_3 VNB N_C1_c_84_n 0.0288566f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.53
cc_4 VNB C1 0.0353647f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB N_C1_c_86_n 0.0458716f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.555
cc_6 VNB N_B1_c_125_n 0.0183366f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.53
cc_7 VNB N_B1_c_126_n 0.0120613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_127_n 0.00714954f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.555
cc_9 VNB N_B2_c_184_n 0.0174245f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.53
cc_10 VNB N_B2_c_185_n 0.0138305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B2_c_186_n 0.00511639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_228_n 0.0416544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_229_n 0.0190512f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.49
cc_14 VNB N_A2_c_230_n 0.00906232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_M1000_g 0.0347467f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.565
cc_16 VNB N_A1_c_279_n 0.0214066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_280_n 0.00380125f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.53
cc_18 VNB N_A1_c_281_n 0.0155575f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_19 VNB N_A1_c_282_n 0.010249f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_20 VNB N_A_27_179#_c_329_n 0.0175239f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_21 VNB N_A_27_179#_c_330_n 0.0158457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_179#_c_331_n 0.0135674f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.555
cc_23 VNB N_A_27_179#_c_332_n 0.0487333f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_435_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.555
cc_25 VNB X 0.0496265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB X 0.0014231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_110_179#_c_514_n 0.0151209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_110_179#_c_515_n 0.00319977f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.53
cc_29 VNB N_A_196_179#_c_543_n 0.0235556f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.565
cc_30 VNB N_A_196_179#_c_544_n 0.00991882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_574_n 0.0126856f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.885
cc_32 VNB N_VGND_c_575_n 0.0158981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_576_n 0.00435083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_577_n 0.0460383f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_35 VNB N_VGND_c_578_n 0.0186844f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.72
cc_36 VNB N_VGND_c_579_n 0.207523f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.555
cc_37 VNB N_VGND_c_580_n 0.00522083f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=0.555
cc_38 VNB N_VGND_c_581_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_C1_c_82_n 0.0432186f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=2.415
cc_40 VPB N_C1_c_88_n 0.0210413f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.565
cc_41 VPB N_C1_c_89_n 0.0320105f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.49
cc_42 VPB N_B1_c_128_n 0.0137543f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.455
cc_43 VPB N_B1_M1003_g 0.0174934f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.53
cc_44 VPB N_B1_c_130_n 0.0277054f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.49
cc_45 VPB B1 0.00133536f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.47
cc_46 VPB N_B1_c_132_n 0.0341536f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B1_c_127_n 0.0101849f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=0.555
cc_48 VPB N_B2_M1011_g 0.0373801f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.105
cc_49 VPB N_B2_c_188_n 0.0350152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B2_c_189_n 0.00358734f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=2.49
cc_51 VPB N_B2_c_186_n 0.00835462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A2_M1008_g 0.0197719f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.72
cc_53 VPB N_A2_c_228_n 0.00879226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A2_c_233_n 0.0208671f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.53
cc_55 VPB N_A2_c_234_n 0.0151345f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A2_c_235_n 0.0153481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A2_c_236_n 0.014805f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=0.555
cc_58 VPB N_A1_M1004_g 0.0530308f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.72
cc_59 VPB N_A1_c_280_n 0.0117897f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.53
cc_60 VPB N_A1_c_282_n 0.00357398f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_61 VPB N_A_27_179#_M1002_g 0.035429f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.53
cc_62 VPB N_A_27_179#_c_331_n 0.0379157f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=0.555
cc_63 VPB N_A_27_179#_c_335_n 0.00763824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_27_179#_c_336_n 0.00285447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_27_179#_c_337_n 0.00647764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_27_179#_c_338_n 0.00660232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_27_179#_c_339_n 0.0397407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_27_179#_c_340_n 0.0166521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_27_179#_c_341_n 0.00174303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_27_179#_c_332_n 0.0192474f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_436_n 0.00563065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_437_n 0.00484152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_438_n 0.0389653f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_74 VPB N_VPWR_c_439_n 0.0197455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_435_n 0.0471025f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=0.555
cc_76 VPB N_VPWR_c_441_n 0.026081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_442_n 0.00362723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_X_c_488_n 0.0180781f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.53
cc_79 VPB N_X_c_489_n 0.0437387f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB X 0.00650483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 N_C1_c_82_n N_B1_c_128_n 0.00330595f $X=0.28 $Y=2.415 $X2=0 $Y2=0
cc_82 N_C1_c_89_n N_B1_M1003_g 0.0155971f $X=0.52 $Y=2.49 $X2=0 $Y2=0
cc_83 N_C1_M1001_g N_B1_c_125_n 0.0140814f $X=0.475 $Y=1.105 $X2=0 $Y2=0
cc_84 C1 N_B1_c_125_n 9.35271e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_85 N_C1_M1001_g N_B1_c_126_n 0.00535697f $X=0.475 $Y=1.105 $X2=0 $Y2=0
cc_86 N_C1_c_89_n N_B1_c_130_n 0.0083665f $X=0.52 $Y=2.49 $X2=0 $Y2=0
cc_87 N_C1_c_82_n B1 2.45426e-19 $X=0.28 $Y=2.415 $X2=0 $Y2=0
cc_88 N_C1_c_82_n N_B1_c_132_n 0.0178931f $X=0.28 $Y=2.415 $X2=0 $Y2=0
cc_89 N_C1_c_82_n N_B1_c_127_n 0.00364272f $X=0.28 $Y=2.415 $X2=0 $Y2=0
cc_90 N_C1_c_84_n N_B1_c_127_n 0.00535697f $X=0.475 $Y=1.53 $X2=0 $Y2=0
cc_91 N_C1_c_82_n N_A_27_179#_c_331_n 0.0264321f $X=0.28 $Y=2.415 $X2=0 $Y2=0
cc_92 N_C1_M1001_g N_A_27_179#_c_331_n 0.0032627f $X=0.475 $Y=1.105 $X2=0 $Y2=0
cc_93 N_C1_c_84_n N_A_27_179#_c_331_n 0.0104235f $X=0.475 $Y=1.53 $X2=0 $Y2=0
cc_94 N_C1_c_89_n N_A_27_179#_c_331_n 0.00390907f $X=0.52 $Y=2.49 $X2=0 $Y2=0
cc_95 C1 N_A_27_179#_c_331_n 0.0123749f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_96 N_C1_c_86_n N_A_27_179#_c_331_n 0.00153263f $X=0.455 $Y=0.555 $X2=0 $Y2=0
cc_97 N_C1_c_88_n N_A_27_179#_c_335_n 0.00603412f $X=0.52 $Y=2.565 $X2=0 $Y2=0
cc_98 N_C1_c_89_n N_A_27_179#_c_335_n 0.006575f $X=0.52 $Y=2.49 $X2=0 $Y2=0
cc_99 N_C1_c_88_n N_A_27_179#_c_340_n 0.0076482f $X=0.52 $Y=2.565 $X2=0 $Y2=0
cc_100 N_C1_c_89_n N_A_27_179#_c_340_n 0.0124164f $X=0.52 $Y=2.49 $X2=0 $Y2=0
cc_101 N_C1_c_88_n N_VPWR_c_436_n 0.00468973f $X=0.52 $Y=2.565 $X2=0 $Y2=0
cc_102 N_C1_c_88_n N_VPWR_c_435_n 0.00732324f $X=0.52 $Y=2.565 $X2=0 $Y2=0
cc_103 N_C1_c_88_n N_VPWR_c_441_n 0.00423721f $X=0.52 $Y=2.565 $X2=0 $Y2=0
cc_104 N_C1_c_89_n N_VPWR_c_441_n 6.13251e-19 $X=0.52 $Y=2.49 $X2=0 $Y2=0
cc_105 C1 N_A_110_179#_c_516_n 0.010764f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_106 N_C1_c_86_n N_A_110_179#_c_516_n 6.55408e-19 $X=0.455 $Y=0.555 $X2=0
+ $Y2=0
cc_107 C1 N_A_110_179#_c_514_n 0.00185174f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_108 N_C1_M1001_g N_A_110_179#_c_515_n 0.00158543f $X=0.475 $Y=1.105 $X2=0
+ $Y2=0
cc_109 N_C1_M1001_g N_A_196_179#_c_544_n 0.00155416f $X=0.475 $Y=1.105 $X2=0
+ $Y2=0
cc_110 C1 N_A_196_179#_c_544_n 0.00433532f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_111 N_C1_c_86_n N_A_196_179#_c_544_n 2.35625e-19 $X=0.455 $Y=0.555 $X2=0
+ $Y2=0
cc_112 C1 N_VGND_c_577_n 0.0264471f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_113 N_C1_c_86_n N_VGND_c_577_n 0.00697212f $X=0.455 $Y=0.555 $X2=0 $Y2=0
cc_114 C1 N_VGND_c_579_n 0.0260444f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_115 N_C1_c_86_n N_VGND_c_579_n 0.0103079f $X=0.455 $Y=0.555 $X2=0 $Y2=0
cc_116 N_B1_c_130_n N_B2_M1011_g 0.0525879f $X=1.115 $Y=2.46 $X2=0 $Y2=0
cc_117 N_B1_c_132_n N_B2_M1011_g 0.00693145f $X=0.76 $Y=2.01 $X2=0 $Y2=0
cc_118 N_B1_c_125_n N_B2_c_184_n 0.0125349f $X=0.877 $Y=1.425 $X2=0 $Y2=0
cc_119 N_B1_c_126_n N_B2_c_185_n 0.00398583f $X=0.877 $Y=1.575 $X2=0 $Y2=0
cc_120 N_B1_c_127_n N_B2_c_185_n 0.00751282f $X=0.775 $Y=1.845 $X2=0 $Y2=0
cc_121 N_B1_c_130_n N_B2_c_188_n 0.00140625f $X=1.115 $Y=2.46 $X2=0 $Y2=0
cc_122 B1 N_B2_c_188_n 2.0853e-19 $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_123 N_B1_c_132_n N_B2_c_188_n 0.0188687f $X=0.76 $Y=2.01 $X2=0 $Y2=0
cc_124 N_B1_c_127_n N_B2_c_188_n 0.00149204f $X=0.775 $Y=1.845 $X2=0 $Y2=0
cc_125 N_B1_c_130_n N_B2_c_189_n 0.00144789f $X=1.115 $Y=2.46 $X2=0 $Y2=0
cc_126 B1 N_B2_c_189_n 0.014069f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_127 N_B1_c_132_n N_B2_c_189_n 0.00362488f $X=0.76 $Y=2.01 $X2=0 $Y2=0
cc_128 N_B1_c_127_n N_B2_c_189_n 6.40721e-19 $X=0.775 $Y=1.845 $X2=0 $Y2=0
cc_129 N_B1_c_128_n N_A_27_179#_c_331_n 0.00502434f $X=0.88 $Y=2.385 $X2=0 $Y2=0
cc_130 N_B1_c_126_n N_A_27_179#_c_331_n 5.2866e-19 $X=0.877 $Y=1.575 $X2=0 $Y2=0
cc_131 N_B1_c_130_n N_A_27_179#_c_331_n 3.57058e-19 $X=1.115 $Y=2.46 $X2=0 $Y2=0
cc_132 B1 N_A_27_179#_c_331_n 0.0118667f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_133 N_B1_c_132_n N_A_27_179#_c_331_n 0.00346371f $X=0.76 $Y=2.01 $X2=0 $Y2=0
cc_134 N_B1_c_127_n N_A_27_179#_c_331_n 0.00508237f $X=0.775 $Y=1.845 $X2=0
+ $Y2=0
cc_135 N_B1_M1003_g N_A_27_179#_c_335_n 0.00784659f $X=1.115 $Y=2.885 $X2=0
+ $Y2=0
cc_136 N_B1_c_130_n N_A_27_179#_c_335_n 0.0166621f $X=1.115 $Y=2.46 $X2=0 $Y2=0
cc_137 B1 N_A_27_179#_c_335_n 0.0127716f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_138 N_B1_c_132_n N_A_27_179#_c_335_n 0.00442744f $X=0.76 $Y=2.01 $X2=0 $Y2=0
cc_139 N_B1_M1003_g N_A_27_179#_c_340_n 8.898e-19 $X=1.115 $Y=2.885 $X2=0 $Y2=0
cc_140 N_B1_M1003_g N_A_27_179#_c_341_n 0.00137063f $X=1.115 $Y=2.885 $X2=0
+ $Y2=0
cc_141 N_B1_c_130_n N_A_27_179#_c_341_n 2.54974e-19 $X=1.115 $Y=2.46 $X2=0 $Y2=0
cc_142 N_B1_M1003_g N_VPWR_c_436_n 0.00696812f $X=1.115 $Y=2.885 $X2=0 $Y2=0
cc_143 N_B1_c_130_n N_VPWR_c_436_n 9.75144e-19 $X=1.115 $Y=2.46 $X2=0 $Y2=0
cc_144 N_B1_M1003_g N_VPWR_c_438_n 0.00429465f $X=1.115 $Y=2.885 $X2=0 $Y2=0
cc_145 N_B1_M1003_g N_VPWR_c_435_n 0.00622319f $X=1.115 $Y=2.885 $X2=0 $Y2=0
cc_146 N_B1_c_125_n N_A_110_179#_c_516_n 2.1266e-19 $X=0.877 $Y=1.425 $X2=0
+ $Y2=0
cc_147 N_B1_c_125_n N_A_110_179#_c_514_n 0.00987759f $X=0.877 $Y=1.425 $X2=0
+ $Y2=0
cc_148 N_B1_c_126_n N_A_110_179#_c_514_n 0.00717469f $X=0.877 $Y=1.575 $X2=0
+ $Y2=0
cc_149 B1 N_A_110_179#_c_514_n 0.0041902f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_150 N_B1_c_126_n N_A_110_179#_c_515_n 0.00148666f $X=0.877 $Y=1.575 $X2=0
+ $Y2=0
cc_151 B1 N_A_110_179#_c_515_n 0.00784719f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_152 N_B1_c_132_n N_A_110_179#_c_515_n 0.00383502f $X=0.76 $Y=2.01 $X2=0 $Y2=0
cc_153 N_B1_c_125_n N_A_196_179#_c_544_n 0.00882041f $X=0.877 $Y=1.425 $X2=0
+ $Y2=0
cc_154 N_B1_c_125_n N_VGND_c_577_n 0.00250212f $X=0.877 $Y=1.425 $X2=0 $Y2=0
cc_155 N_B1_c_125_n N_VGND_c_579_n 0.00334041f $X=0.877 $Y=1.425 $X2=0 $Y2=0
cc_156 N_B2_M1011_g N_A2_M1008_g 0.0153515f $X=1.475 $Y=2.885 $X2=0 $Y2=0
cc_157 N_B2_c_185_n N_A2_c_228_n 0.0109471f $X=1.5 $Y=1.605 $X2=0 $Y2=0
cc_158 N_B2_c_186_n N_A2_c_228_n 0.00892089f $X=1.357 $Y=1.815 $X2=0 $Y2=0
cc_159 N_B2_M1011_g N_A2_c_233_n 0.0201196f $X=1.475 $Y=2.885 $X2=0 $Y2=0
cc_160 N_B2_c_184_n N_A2_c_230_n 0.0109471f $X=1.5 $Y=1.455 $X2=0 $Y2=0
cc_161 N_B2_c_188_n N_A2_c_235_n 0.0201196f $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_162 N_B2_c_189_n N_A2_c_235_n 2.2626e-19 $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_163 N_B2_c_188_n N_A2_c_236_n 0.0121915f $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_164 N_B2_c_189_n N_A2_c_236_n 0.0230368f $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_165 N_B2_c_188_n N_A_27_179#_c_335_n 0.00116195f $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_166 N_B2_c_189_n N_A_27_179#_c_335_n 0.00562289f $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_167 N_B2_M1011_g N_A_27_179#_c_368_n 0.012947f $X=1.475 $Y=2.885 $X2=0 $Y2=0
cc_168 N_B2_M1011_g N_A_27_179#_c_341_n 0.00807998f $X=1.475 $Y=2.885 $X2=0
+ $Y2=0
cc_169 N_B2_c_188_n N_A_27_179#_c_341_n 0.00317556f $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_170 N_B2_c_189_n N_A_27_179#_c_341_n 0.00804507f $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_171 N_B2_M1011_g N_VPWR_c_438_n 0.00369552f $X=1.475 $Y=2.885 $X2=0 $Y2=0
cc_172 N_B2_M1011_g N_VPWR_c_435_n 0.00529079f $X=1.475 $Y=2.885 $X2=0 $Y2=0
cc_173 N_B2_c_184_n N_A_110_179#_c_514_n 0.00878978f $X=1.5 $Y=1.455 $X2=0 $Y2=0
cc_174 N_B2_c_185_n N_A_110_179#_c_514_n 0.0106241f $X=1.5 $Y=1.605 $X2=0 $Y2=0
cc_175 N_B2_c_188_n N_A_110_179#_c_514_n 0.00473872f $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_176 N_B2_c_189_n N_A_110_179#_c_514_n 0.0142236f $X=1.33 $Y=1.98 $X2=0 $Y2=0
cc_177 N_B2_c_184_n N_A_196_179#_c_543_n 0.00763902f $X=1.5 $Y=1.455 $X2=0 $Y2=0
cc_178 N_B2_c_185_n N_A_196_179#_c_543_n 2.19762e-19 $X=1.5 $Y=1.605 $X2=0 $Y2=0
cc_179 N_B2_c_184_n N_A_196_179#_c_544_n 0.00709916f $X=1.5 $Y=1.455 $X2=0 $Y2=0
cc_180 N_A2_M1008_g N_A1_M1004_g 0.027156f $X=1.905 $Y=2.885 $X2=0 $Y2=0
cc_181 N_A2_c_234_n N_A1_M1004_g 0.0221427f $X=1.925 $Y=2.515 $X2=0 $Y2=0
cc_182 N_A2_c_236_n N_A1_M1004_g 0.00117881f $X=1.925 $Y=2.01 $X2=0 $Y2=0
cc_183 N_A2_c_228_n N_A1_M1000_g 0.00834015f $X=1.925 $Y=1.845 $X2=0 $Y2=0
cc_184 N_A2_c_229_n N_A1_M1000_g 0.0211344f $X=2.02 $Y=0.765 $X2=0 $Y2=0
cc_185 N_A2_c_235_n N_A1_c_279_n 0.0221427f $X=1.925 $Y=2.01 $X2=0 $Y2=0
cc_186 N_A2_c_233_n N_A1_c_280_n 0.0221427f $X=1.925 $Y=2.35 $X2=0 $Y2=0
cc_187 N_A2_c_228_n N_A1_c_281_n 0.0221427f $X=1.925 $Y=1.845 $X2=0 $Y2=0
cc_188 N_A2_c_228_n N_A1_c_282_n 0.00321697f $X=1.925 $Y=1.845 $X2=0 $Y2=0
cc_189 N_A2_M1008_g N_A_27_179#_c_368_n 0.0126392f $X=1.905 $Y=2.885 $X2=0 $Y2=0
cc_190 N_A2_c_234_n N_A_27_179#_c_368_n 0.00335335f $X=1.925 $Y=2.515 $X2=0
+ $Y2=0
cc_191 N_A2_c_236_n N_A_27_179#_c_368_n 0.0279975f $X=1.925 $Y=2.01 $X2=0 $Y2=0
cc_192 N_A2_M1008_g N_A_27_179#_c_336_n 0.0035961f $X=1.905 $Y=2.885 $X2=0 $Y2=0
cc_193 N_A2_c_233_n N_A_27_179#_c_336_n 0.00132907f $X=1.925 $Y=2.35 $X2=0 $Y2=0
cc_194 N_A2_c_236_n N_A_27_179#_c_336_n 0.0156774f $X=1.925 $Y=2.01 $X2=0 $Y2=0
cc_195 N_A2_c_235_n N_A_27_179#_c_337_n 0.00239088f $X=1.925 $Y=2.01 $X2=0 $Y2=0
cc_196 N_A2_c_236_n N_A_27_179#_c_337_n 0.0271676f $X=1.925 $Y=2.01 $X2=0 $Y2=0
cc_197 N_A2_M1008_g N_A_27_179#_c_341_n 8.27787e-19 $X=1.905 $Y=2.885 $X2=0
+ $Y2=0
cc_198 N_A2_c_236_n N_A_27_179#_c_341_n 0.00147478f $X=1.925 $Y=2.01 $X2=0 $Y2=0
cc_199 N_A2_M1008_g N_VPWR_c_438_n 0.00368123f $X=1.905 $Y=2.885 $X2=0 $Y2=0
cc_200 N_A2_M1008_g N_VPWR_c_435_n 0.00559621f $X=1.905 $Y=2.885 $X2=0 $Y2=0
cc_201 N_A2_c_228_n N_A_110_179#_c_514_n 0.00221593f $X=1.925 $Y=1.845 $X2=0
+ $Y2=0
cc_202 N_A2_c_235_n N_A_110_179#_c_514_n 5.74635e-19 $X=1.925 $Y=2.01 $X2=0
+ $Y2=0
cc_203 N_A2_c_236_n N_A_110_179#_c_514_n 0.013093f $X=1.925 $Y=2.01 $X2=0 $Y2=0
cc_204 N_A2_c_228_n N_A_110_179#_c_534_n 0.00390481f $X=1.925 $Y=1.845 $X2=0
+ $Y2=0
cc_205 N_A2_c_229_n N_A_196_179#_c_543_n 0.0080112f $X=2.02 $Y=0.765 $X2=0 $Y2=0
cc_206 N_A2_c_230_n N_A_196_179#_c_543_n 0.0100859f $X=2.02 $Y=0.915 $X2=0 $Y2=0
cc_207 N_A2_c_229_n N_A_196_179#_c_554_n 2.1266e-19 $X=2.02 $Y=0.765 $X2=0 $Y2=0
cc_208 N_A2_c_229_n N_A_196_179#_c_544_n 2.03062e-19 $X=2.02 $Y=0.765 $X2=0
+ $Y2=0
cc_209 N_A2_c_229_n N_VGND_c_574_n 0.00742523f $X=2.02 $Y=0.765 $X2=0 $Y2=0
cc_210 N_A2_c_229_n N_VGND_c_575_n 0.00414412f $X=2.02 $Y=0.765 $X2=0 $Y2=0
cc_211 N_A2_c_229_n N_VGND_c_579_n 0.00486498f $X=2.02 $Y=0.765 $X2=0 $Y2=0
cc_212 N_A1_M1004_g N_A_27_179#_M1002_g 0.0222221f $X=2.375 $Y=2.885 $X2=0 $Y2=0
cc_213 N_A1_M1000_g N_A_27_179#_c_329_n 0.0195747f $X=2.455 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A1_M1004_g N_A_27_179#_c_368_n 0.00993068f $X=2.375 $Y=2.885 $X2=0
+ $Y2=0
cc_215 N_A1_M1004_g N_A_27_179#_c_336_n 0.0102806f $X=2.375 $Y=2.885 $X2=0 $Y2=0
cc_216 N_A1_M1004_g N_A_27_179#_c_337_n 0.00434406f $X=2.375 $Y=2.885 $X2=0
+ $Y2=0
cc_217 N_A1_c_282_n N_A_27_179#_c_337_n 0.00420508f $X=2.465 $Y=1.255 $X2=0
+ $Y2=0
cc_218 N_A1_M1004_g N_A_27_179#_c_338_n 0.0113346f $X=2.375 $Y=2.885 $X2=0 $Y2=0
cc_219 N_A1_c_280_n N_A_27_179#_c_338_n 0.00127164f $X=2.465 $Y=1.76 $X2=0 $Y2=0
cc_220 N_A1_c_282_n N_A_27_179#_c_338_n 0.0293659f $X=2.465 $Y=1.255 $X2=0 $Y2=0
cc_221 N_A1_M1004_g N_A_27_179#_c_339_n 0.0213434f $X=2.375 $Y=2.885 $X2=0 $Y2=0
cc_222 N_A1_c_282_n N_A_27_179#_c_339_n 0.00262891f $X=2.465 $Y=1.255 $X2=0
+ $Y2=0
cc_223 N_A1_M1004_g N_A_27_179#_c_332_n 0.00642957f $X=2.375 $Y=2.885 $X2=0
+ $Y2=0
cc_224 N_A1_M1000_g N_A_27_179#_c_332_n 0.00781354f $X=2.455 $Y=0.445 $X2=0
+ $Y2=0
cc_225 N_A1_c_281_n N_A_27_179#_c_332_n 0.0330195f $X=2.465 $Y=1.255 $X2=0 $Y2=0
cc_226 N_A1_c_282_n N_A_27_179#_c_332_n 0.00501972f $X=2.465 $Y=1.255 $X2=0
+ $Y2=0
cc_227 N_A1_M1004_g N_VPWR_c_437_n 0.00453563f $X=2.375 $Y=2.885 $X2=0 $Y2=0
cc_228 N_A1_M1004_g N_VPWR_c_438_n 0.004984f $X=2.375 $Y=2.885 $X2=0 $Y2=0
cc_229 N_A1_M1004_g N_VPWR_c_435_n 0.00886845f $X=2.375 $Y=2.885 $X2=0 $Y2=0
cc_230 N_A1_c_282_n N_X_c_489_n 5.0653e-19 $X=2.465 $Y=1.255 $X2=0 $Y2=0
cc_231 N_A1_M1000_g X 0.00148088f $X=2.455 $Y=0.445 $X2=0 $Y2=0
cc_232 N_A1_c_281_n X 2.74948e-19 $X=2.465 $Y=1.255 $X2=0 $Y2=0
cc_233 N_A1_c_282_n X 0.0436709f $X=2.465 $Y=1.255 $X2=0 $Y2=0
cc_234 N_A1_c_279_n X 2.74948e-19 $X=2.465 $Y=1.595 $X2=0 $Y2=0
cc_235 N_A1_c_282_n N_A_110_179#_c_514_n 0.00697912f $X=2.465 $Y=1.255 $X2=0
+ $Y2=0
cc_236 N_A1_c_282_n N_A_110_179#_c_534_n 0.00840326f $X=2.465 $Y=1.255 $X2=0
+ $Y2=0
cc_237 N_A1_M1000_g N_A_196_179#_c_543_n 0.00287294f $X=2.455 $Y=0.445 $X2=0
+ $Y2=0
cc_238 N_A1_c_281_n N_A_196_179#_c_543_n 3.14764e-19 $X=2.465 $Y=1.255 $X2=0
+ $Y2=0
cc_239 N_A1_c_282_n N_A_196_179#_c_543_n 0.00281565f $X=2.465 $Y=1.255 $X2=0
+ $Y2=0
cc_240 N_A1_M1000_g N_VGND_c_574_n 7.33522e-19 $X=2.455 $Y=0.445 $X2=0 $Y2=0
cc_241 N_A1_M1000_g N_VGND_c_575_n 0.00585385f $X=2.455 $Y=0.445 $X2=0 $Y2=0
cc_242 N_A1_M1000_g N_VGND_c_576_n 0.00151442f $X=2.455 $Y=0.445 $X2=0 $Y2=0
cc_243 N_A1_c_281_n N_VGND_c_576_n 3.16663e-19 $X=2.465 $Y=1.255 $X2=0 $Y2=0
cc_244 N_A1_c_282_n N_VGND_c_576_n 0.00711076f $X=2.465 $Y=1.255 $X2=0 $Y2=0
cc_245 N_A1_M1000_g N_VGND_c_579_n 0.0107511f $X=2.455 $Y=0.445 $X2=0 $Y2=0
cc_246 N_A_27_179#_c_335_n N_VPWR_c_436_n 0.0243509f $X=1.245 $Y=2.58 $X2=0
+ $Y2=0
cc_247 N_A_27_179#_M1002_g N_VPWR_c_437_n 0.00291137f $X=2.84 $Y=2.885 $X2=0
+ $Y2=0
cc_248 N_A_27_179#_c_368_n N_VPWR_c_437_n 0.0181826f $X=2.19 $Y=2.86 $X2=0 $Y2=0
cc_249 N_A_27_179#_c_338_n N_VPWR_c_437_n 0.00691098f $X=2.825 $Y=2.135 $X2=0
+ $Y2=0
cc_250 N_A_27_179#_c_339_n N_VPWR_c_437_n 0.00120879f $X=2.825 $Y=2.135 $X2=0
+ $Y2=0
cc_251 N_A_27_179#_c_335_n N_VPWR_c_438_n 0.00424746f $X=1.245 $Y=2.58 $X2=0
+ $Y2=0
cc_252 N_A_27_179#_c_368_n N_VPWR_c_438_n 0.0418789f $X=2.19 $Y=2.86 $X2=0 $Y2=0
cc_253 N_A_27_179#_c_341_n N_VPWR_c_438_n 0.00730918f $X=1.33 $Y=2.58 $X2=0
+ $Y2=0
cc_254 N_A_27_179#_M1002_g N_VPWR_c_439_n 0.00585385f $X=2.84 $Y=2.885 $X2=0
+ $Y2=0
cc_255 N_A_27_179#_M1010_s N_VPWR_c_435_n 0.00235821f $X=0.18 $Y=2.675 $X2=0
+ $Y2=0
cc_256 N_A_27_179#_M1011_d N_VPWR_c_435_n 0.00228308f $X=1.55 $Y=2.675 $X2=0
+ $Y2=0
cc_257 N_A_27_179#_M1002_g N_VPWR_c_435_n 0.0118535f $X=2.84 $Y=2.885 $X2=0
+ $Y2=0
cc_258 N_A_27_179#_c_335_n N_VPWR_c_435_n 0.0125076f $X=1.245 $Y=2.58 $X2=0
+ $Y2=0
cc_259 N_A_27_179#_c_368_n N_VPWR_c_435_n 0.0335288f $X=2.19 $Y=2.86 $X2=0 $Y2=0
cc_260 N_A_27_179#_c_340_n N_VPWR_c_435_n 0.0115132f $X=0.305 $Y=2.58 $X2=0
+ $Y2=0
cc_261 N_A_27_179#_c_341_n N_VPWR_c_435_n 0.00624785f $X=1.33 $Y=2.58 $X2=0
+ $Y2=0
cc_262 N_A_27_179#_c_335_n N_VPWR_c_441_n 0.00283869f $X=1.245 $Y=2.58 $X2=0
+ $Y2=0
cc_263 N_A_27_179#_c_340_n N_VPWR_c_441_n 0.0106141f $X=0.305 $Y=2.58 $X2=0
+ $Y2=0
cc_264 N_A_27_179#_c_341_n A_238_535# 0.00103573f $X=1.33 $Y=2.58 $X2=-0.19
+ $Y2=-0.245
cc_265 N_A_27_179#_c_368_n A_396_535# 0.00694732f $X=2.19 $Y=2.86 $X2=-0.19
+ $Y2=-0.245
cc_266 N_A_27_179#_c_336_n A_396_535# 2.26742e-19 $X=2.275 $Y=2.695 $X2=-0.19
+ $Y2=-0.245
cc_267 N_A_27_179#_M1002_g N_X_c_488_n 5.45259e-19 $X=2.84 $Y=2.885 $X2=0 $Y2=0
cc_268 N_A_27_179#_c_336_n N_X_c_488_n 7.69639e-19 $X=2.275 $Y=2.695 $X2=0 $Y2=0
cc_269 N_A_27_179#_c_339_n N_X_c_488_n 0.00255109f $X=2.825 $Y=2.135 $X2=0 $Y2=0
cc_270 N_A_27_179#_M1002_g N_X_c_489_n 0.0120718f $X=2.84 $Y=2.885 $X2=0 $Y2=0
cc_271 N_A_27_179#_c_338_n N_X_c_489_n 0.0252087f $X=2.825 $Y=2.135 $X2=0 $Y2=0
cc_272 N_A_27_179#_c_332_n N_X_c_489_n 0.0167853f $X=2.84 $Y=1.97 $X2=0 $Y2=0
cc_273 N_A_27_179#_c_329_n X 0.00218306f $X=2.915 $Y=0.73 $X2=0 $Y2=0
cc_274 N_A_27_179#_c_330_n X 0.00642975f $X=2.915 $Y=0.88 $X2=0 $Y2=0
cc_275 N_A_27_179#_c_332_n X 0.0239315f $X=2.84 $Y=1.97 $X2=0 $Y2=0
cc_276 N_A_27_179#_c_332_n X 0.00518941f $X=2.84 $Y=1.97 $X2=0 $Y2=0
cc_277 N_A_27_179#_c_331_n N_A_110_179#_c_516_n 5.54215e-19 $X=0.26 $Y=1.17
+ $X2=0 $Y2=0
cc_278 N_A_27_179#_c_331_n N_A_110_179#_c_515_n 0.0120352f $X=0.26 $Y=1.17 $X2=0
+ $Y2=0
cc_279 N_A_27_179#_c_329_n N_VGND_c_576_n 0.00288714f $X=2.915 $Y=0.73 $X2=0
+ $Y2=0
cc_280 N_A_27_179#_c_329_n N_VGND_c_578_n 0.00585385f $X=2.915 $Y=0.73 $X2=0
+ $Y2=0
cc_281 N_A_27_179#_c_330_n N_VGND_c_578_n 8.06102e-19 $X=2.915 $Y=0.88 $X2=0
+ $Y2=0
cc_282 N_A_27_179#_c_329_n N_VGND_c_579_n 0.0117282f $X=2.915 $Y=0.73 $X2=0
+ $Y2=0
cc_283 N_A_27_179#_c_330_n N_VGND_c_579_n 9.8182e-19 $X=2.915 $Y=0.88 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_435_n A_238_535# 0.00191866f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_285 N_VPWR_c_435_n A_396_535# 0.00260882f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_286 N_VPWR_c_435_n N_X_M1002_d 0.00344799f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_287 N_VPWR_c_439_n N_X_c_488_n 0.0126729f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_288 N_VPWR_c_435_n N_X_c_488_n 0.0112063f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_289 X N_A_196_179#_c_543_n 0.00529389f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_290 X N_A_196_179#_c_554_n 2.58893e-19 $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_291 X N_VGND_c_578_n 0.0112582f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_292 N_X_M1006_d N_VGND_c_579_n 0.00264243f $X=2.96 $Y=0.235 $X2=0 $Y2=0
cc_293 X N_VGND_c_579_n 0.00974255f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_294 N_A_110_179#_c_514_n N_A_196_179#_M1009_d 0.00344211f $X=1.635 $Y=1.41
+ $X2=-0.19 $Y2=-0.245
cc_295 N_A_110_179#_c_514_n N_A_196_179#_c_543_n 0.00639579f $X=1.635 $Y=1.41
+ $X2=0 $Y2=0
cc_296 N_A_110_179#_c_534_n N_A_196_179#_c_543_n 0.0140281f $X=1.74 $Y=1.2 $X2=0
+ $Y2=0
cc_297 N_A_110_179#_c_514_n N_A_196_179#_c_544_n 0.0249115f $X=1.635 $Y=1.41
+ $X2=0 $Y2=0
cc_298 N_A_196_179#_c_543_n N_VGND_c_574_n 0.022009f $X=2.135 $Y=0.75 $X2=0
+ $Y2=0
cc_299 N_A_196_179#_c_543_n N_VGND_c_575_n 0.002793f $X=2.135 $Y=0.75 $X2=0
+ $Y2=0
cc_300 N_A_196_179#_c_554_n N_VGND_c_575_n 0.0081737f $X=2.24 $Y=0.51 $X2=0
+ $Y2=0
cc_301 N_A_196_179#_c_543_n N_VGND_c_577_n 0.00418704f $X=2.135 $Y=0.75 $X2=0
+ $Y2=0
cc_302 N_A_196_179#_c_544_n N_VGND_c_577_n 0.00608292f $X=1.215 $Y=0.75 $X2=0
+ $Y2=0
cc_303 N_A_196_179#_M1007_d N_VGND_c_579_n 0.00369956f $X=2.1 $Y=0.235 $X2=0
+ $Y2=0
cc_304 N_A_196_179#_c_543_n N_VGND_c_579_n 0.0126301f $X=2.135 $Y=0.75 $X2=0
+ $Y2=0
cc_305 N_A_196_179#_c_554_n N_VGND_c_579_n 0.00762225f $X=2.24 $Y=0.51 $X2=0
+ $Y2=0
cc_306 N_A_196_179#_c_544_n N_VGND_c_579_n 0.00957819f $X=1.215 $Y=0.75 $X2=0
+ $Y2=0
