* NGSPICE file created from sky130_fd_sc_lp__a2bb2o_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2bb2o_m A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VPWR a_85_345# X VPB phighvt w=420000u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=1.197e+11p ps=1.41e+06u
M1001 VGND A2_N a_210_125# VNB nshort w=420000u l=150000u
+  ad=3.465e+11p pd=4.17e+06u as=2.2975e+11p ps=2.03e+06u
M1002 a_85_345# a_210_125# VGND VNB nshort w=420000u l=150000u
+  ad=2.247e+11p pd=1.91e+06u as=0p ps=0u
M1003 a_223_535# A1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_210_125# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B2 a_479_429# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.289e+11p ps=2.77e+06u
M1006 VGND a_85_345# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1007 a_210_125# A2_N a_223_535# VPB phighvt w=420000u l=150000u
+  ad=1.141e+11p pd=1.41e+06u as=0p ps=0u
M1008 a_479_429# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_551_125# B2 a_85_345# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1010 VGND B1 a_551_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_479_429# a_210_125# a_85_345# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.141e+11p ps=1.41e+06u
.ends

