* NGSPICE file created from sky130_fd_sc_lp__or4b_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or4b_2 A B C D_N VGND VNB VPB VPWR X
M1000 X a_189_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=8.148e+11p ps=6.8e+06u
M1001 a_189_21# C VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=8.085e+11p ps=7.83e+06u
M1002 X a_189_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1003 a_436_385# A VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 a_616_385# C a_508_385# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.638e+11p ps=1.62e+06u
M1005 VGND B a_189_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_189_21# a_31_131# a_616_385# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 VGND a_189_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR D_N a_31_131# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 VPWR a_189_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_189_21# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_31_131# a_189_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D_N a_31_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1013 a_508_385# B a_436_385# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

