* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 VPWR A1_N a_462_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.2823e+12p pd=2.285e+07u as=7.056e+11p ps=6.16e+06u
M1001 a_218_367# a_462_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=0p ps=0u
M1002 VGND a_218_367# X VNB nshort w=840000u l=150000u
+  ad=1.7388e+12p pd=1.422e+07u as=4.704e+11p ps=4.48e+06u
M1003 a_49_47# a_462_21# a_218_367# VNB nshort w=840000u l=150000u
+  ad=9.156e+11p pd=8.9e+06u as=2.352e+11p ps=2.24e+06u
M1004 VGND A1_N a_768_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.48e+06u
M1005 VGND a_218_367# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_49_47# B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_768_47# A1_N VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_218_367# B2 a_132_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.16e+06u
M1009 VGND B1 a_49_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_218_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=0p ps=0u
M1011 VPWR B1 a_132_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A2_N a_462_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_218_367# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_49_47# B2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_218_367# a_462_21# a_49_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_462_21# A2_N a_768_47# VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1017 X a_218_367# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_218_367# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_462_21# a_218_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_462_21# A2_N VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_132_367# B2 a_218_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_462_21# A1_N VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_218_367# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND B2 a_49_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_768_47# A2_N a_462_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_132_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_218_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
