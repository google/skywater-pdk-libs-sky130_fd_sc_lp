* File: sky130_fd_sc_lp__dfxbp_2.pex.spice
* Created: Wed Sep  2 09:44:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFXBP_2%CLK 3 6 9 10 11 12 13 14 19
r29 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.045 $X2=0.385 $Y2=1.045
r30 13 14 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.295
+ $X2=0.28 $Y2=1.665
r31 13 20 7.58186 $w=3.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.28 $Y=1.295
+ $X2=0.28 $Y2=1.045
r32 12 20 3.63929 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=0.28 $Y=0.925
+ $X2=0.28 $Y2=1.045
r33 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.385
+ $X2=0.385 $Y2=1.045
r34 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.385
+ $X2=0.385 $Y2=1.55
r35 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=0.88
+ $X2=0.385 $Y2=1.045
r36 6 11 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.475 $Y=2.61
+ $X2=0.475 $Y2=1.55
r37 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.56
+ $X2=0.475 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%D 3 6 9 10 11 12 13 14 19
c38 12 0 1.23912e-19 $X=2.16 $Y=1.295
c39 6 0 1.28884e-19 $X=2.22 $Y=2.525
r40 13 14 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.125 $Y=1.665
+ $X2=2.125 $Y2=2.035
r41 12 13 16.6218 $w=2.58e-07 $l=3.75e-07 $layer=LI1_cond $X=2.125 $Y=1.29
+ $X2=2.125 $Y2=1.665
r42 12 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.16
+ $Y=1.29 $X2=2.16 $Y2=1.29
r43 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.16 $Y=1.63
+ $X2=2.16 $Y2=1.29
r44 10 11 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.63
+ $X2=2.16 $Y2=1.795
r45 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.125
+ $X2=2.16 $Y2=1.29
r46 6 11 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.22 $Y=2.525
+ $X2=2.22 $Y2=1.795
r47 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.07 $Y=0.805 $X2=2.07
+ $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%A_236_463# 1 2 9 12 15 19 21 23 25 32 34 37
+ 38 39 40 41 42 46 50 53 56 62
c167 50 0 2.13954e-20 $X=1.305 $Y=2.46
c168 38 0 1.82964e-19 $X=3.305 $Y=2.99
c169 12 0 1.05623e-19 $X=2.725 $Y=2.08
r170 55 56 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.065 $Y=1.99
+ $X2=2.99 $Y2=1.99
r171 53 55 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.29 $Y=1.99
+ $X2=3.065 $Y2=1.99
r172 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.29
+ $Y=1.99 $X2=3.29 $Y2=1.99
r173 47 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.34
+ $X2=5.215 $Y2=1.34
r174 47 59 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=5.05 $Y=1.34
+ $X2=4.93 $Y2=1.34
r175 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=1.34 $X2=5.05 $Y2=1.34
r176 44 46 52.244 $w=1.88e-07 $l=8.95e-07 $layer=LI1_cond $X=5.05 $Y=2.235
+ $X2=5.05 $Y2=1.34
r177 43 52 15.4253 $w=2.61e-07 $l=4.08228e-07 $layer=LI1_cond $X=3.475 $Y=2.32
+ $X2=3.3 $Y2=1.99
r178 42 44 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.955 $Y=2.32
+ $X2=5.05 $Y2=2.235
r179 42 43 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=4.955 $Y=2.32
+ $X2=3.475 $Y2=2.32
r180 40 43 5.45457 $w=2.61e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.39 $Y=2.405
+ $X2=3.475 $Y2=2.32
r181 40 41 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.39 $Y=2.405
+ $X2=3.39 $Y2=2.905
r182 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.305 $Y=2.99
+ $X2=3.39 $Y2=2.905
r183 38 39 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=3.305 $Y=2.99
+ $X2=2.17 $Y2=2.99
r184 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.085 $Y=2.905
+ $X2=2.17 $Y2=2.99
r185 36 37 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.085 $Y=2.47
+ $X2=2.085 $Y2=2.905
r186 35 50 2.98021 $w=1.7e-07 $l=1.69493e-07 $layer=LI1_cond $X=1.475 $Y=2.385
+ $X2=1.307 $Y2=2.382
r187 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2 $Y=2.385
+ $X2=2.085 $Y2=2.47
r188 34 35 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2 $Y=2.385
+ $X2=1.475 $Y2=2.385
r189 30 50 3.52026 $w=2.65e-07 $l=1.04283e-07 $layer=LI1_cond $X=1.345 $Y=2.295
+ $X2=1.307 $Y2=2.382
r190 30 32 66.0438 $w=2.58e-07 $l=1.49e-06 $layer=LI1_cond $X=1.345 $Y=2.295
+ $X2=1.345 $Y2=0.805
r191 23 27 56.1165 $w=2.22e-07 $l=2.69907e-07 $layer=POLY_cond $X=5.71 $Y=1.665
+ $X2=5.635 $Y2=1.43
r192 23 25 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.71 $Y=1.665
+ $X2=5.71 $Y2=2.475
r193 21 27 11.9802 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.485 $Y=1.43
+ $X2=5.635 $Y2=1.43
r194 21 62 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.485 $Y=1.43
+ $X2=5.215 $Y2=1.43
r195 17 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.93 $Y=1.175
+ $X2=4.93 $Y2=1.34
r196 17 19 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.93 $Y=1.175
+ $X2=4.93 $Y2=0.805
r197 13 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.825
+ $X2=3.065 $Y2=1.99
r198 13 15 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.065 $Y=1.825
+ $X2=3.065 $Y2=0.805
r199 12 56 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.725 $Y=2.08
+ $X2=2.99 $Y2=2.08
r200 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.65 $Y=2.155
+ $X2=2.725 $Y2=2.08
r201 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.65 $Y=2.155
+ $X2=2.65 $Y2=2.525
r202 2 50 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.18
+ $Y=2.315 $X2=1.305 $Y2=2.46
r203 1 32 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.255
+ $Y=0.595 $X2=1.38 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%A_670_93# 1 2 7 9 14 16 17 18 22 26 28 35 39
c73 28 0 1.10981e-19 $X=3.65 $Y=1.09
c74 26 0 8.34361e-20 $X=4.62 $Y=0.75
c75 16 0 1.38922e-19 $X=3.76 $Y=1.925
r76 32 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.65 $Y=1.29 $X2=3.74
+ $Y2=1.29
r77 32 36 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.65 $Y=1.29
+ $X2=3.425 $Y2=1.29
r78 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.65
+ $Y=1.29 $X2=3.65 $Y2=1.29
r79 28 31 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.65 $Y=1.09 $X2=3.65
+ $Y2=1.29
r80 24 35 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.655 $Y=1.005
+ $X2=4.62 $Y2=1.09
r81 24 26 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=4.655 $Y=1.005
+ $X2=4.655 $Y2=0.75
r82 20 35 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=1.175
+ $X2=4.62 $Y2=1.09
r83 20 22 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=4.62 $Y=1.175
+ $X2=4.62 $Y2=1.97
r84 19 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=1.09
+ $X2=3.65 $Y2=1.09
r85 18 35 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=1.09
+ $X2=4.62 $Y2=1.09
r86 18 19 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.455 $Y=1.09
+ $X2=3.815 $Y2=1.09
r87 16 17 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=3.76 $Y=1.925
+ $X2=3.76 $Y2=2.075
r88 14 17 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.78 $Y=2.525
+ $X2=3.78 $Y2=2.075
r89 10 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.74 $Y=1.455
+ $X2=3.74 $Y2=1.29
r90 10 16 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.74 $Y=1.455 $X2=3.74
+ $Y2=1.925
r91 7 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=1.125
+ $X2=3.425 $Y2=1.29
r92 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.425 $Y=1.125
+ $X2=3.425 $Y2=0.805
r93 2 22 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.845 $X2=4.62 $Y2=1.97
r94 1 35 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=4.48
+ $Y=0.595 $X2=4.62 $Y2=1.09
r95 1 26 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.48
+ $Y=0.595 $X2=4.62 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%A_537_119# 1 2 7 9 12 16 19 20 22 26 29 36
c76 36 0 1.10981e-19 $X=4.405 $Y=1.52
c77 29 0 1.38922e-19 $X=4.19 $Y=1.52
c78 7 0 8.34361e-20 $X=4.405 $Y=1.355
r79 30 36 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.19 $Y=1.52
+ $X2=4.405 $Y2=1.52
r80 29 32 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=4.155 $Y=1.52
+ $X2=4.155 $Y2=1.64
r81 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.19
+ $Y=1.52 $X2=4.19 $Y2=1.52
r82 23 26 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.855 $Y=2.57
+ $X2=2.96 $Y2=2.57
r83 21 22 2.20034 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.015 $Y=1.64
+ $X2=2.89 $Y2=1.64
r84 20 32 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.025 $Y=1.64
+ $X2=4.155 $Y2=1.64
r85 20 21 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.025 $Y=1.64
+ $X2=3.015 $Y2=1.64
r86 19 23 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=2.405
+ $X2=2.855 $Y2=2.57
r87 18 22 4.23118 $w=2.15e-07 $l=1.00995e-07 $layer=LI1_cond $X=2.855 $Y=1.725
+ $X2=2.89 $Y2=1.64
r88 18 19 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.855 $Y=1.725
+ $X2=2.855 $Y2=2.405
r89 14 22 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=1.555
+ $X2=2.89 $Y2=1.64
r90 14 16 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=2.89 $Y=1.555
+ $X2=2.89 $Y2=0.805
r91 10 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=1.685
+ $X2=4.405 $Y2=1.52
r92 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.405 $Y=1.685
+ $X2=4.405 $Y2=2.265
r93 7 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=1.355
+ $X2=4.405 $Y2=1.52
r94 7 9 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.405 $Y=1.355
+ $X2=4.405 $Y2=0.915
r95 2 26 600 $w=1.7e-07 $l=3.53483e-07 $layer=licon1_PDIFF $count=1 $X=2.725
+ $Y=2.315 $X2=2.96 $Y2=2.57
r96 1 16 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=2.685
+ $Y=0.595 $X2=2.85 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%A_110_70# 1 2 7 8 12 16 17 18 19 20 23 25 29
+ 31 35 39 42 43 44 47 50 52 53 61
c133 29 0 5.07986e-20 $X=3.27 $Y=2.705
c134 23 0 1.82889e-20 $X=2.61 $Y=0.805
r135 59 61 6.64871 $w=3.88e-07 $l=2.25e-07 $layer=LI1_cond $X=0.69 $Y=0.525
+ $X2=0.915 $Y2=0.525
r136 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=1.595 $X2=0.955 $Y2=1.595
r137 50 52 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.915 $Y=1.93
+ $X2=0.915 $Y2=1.595
r138 49 61 3.33926 $w=2.5e-07 $l=1.95e-07 $layer=LI1_cond $X=0.915 $Y=0.72
+ $X2=0.915 $Y2=0.525
r139 49 52 40.3355 $w=2.48e-07 $l=8.75e-07 $layer=LI1_cond $X=0.915 $Y=0.72
+ $X2=0.915 $Y2=1.595
r140 45 50 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.715 $Y=2.015
+ $X2=0.915 $Y2=2.015
r141 45 47 14.1997 $w=2.78e-07 $l=3.45e-07 $layer=LI1_cond $X=0.715 $Y=2.1
+ $X2=0.715 $Y2=2.445
r142 41 53 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.955 $Y=1.58
+ $X2=0.955 $Y2=1.595
r143 37 39 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.55 $Y=0.255
+ $X2=5.55 $Y2=0.805
r144 33 35 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.835 $Y=3.075
+ $X2=4.835 $Y2=2.265
r145 32 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.345 $Y=3.15
+ $X2=3.27 $Y2=3.15
r146 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.76 $Y=3.15
+ $X2=4.835 $Y2=3.075
r147 31 32 725.564 $w=1.5e-07 $l=1.415e-06 $layer=POLY_cond $X=4.76 $Y=3.15
+ $X2=3.345 $Y2=3.15
r148 27 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.27 $Y=3.075
+ $X2=3.27 $Y2=3.15
r149 27 29 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.27 $Y=3.075
+ $X2=3.27 $Y2=2.705
r150 26 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.685 $Y=0.18
+ $X2=2.61 $Y2=0.18
r151 25 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.475 $Y=0.18
+ $X2=5.55 $Y2=0.255
r152 25 26 1430.62 $w=1.5e-07 $l=2.79e-06 $layer=POLY_cond $X=5.475 $Y=0.18
+ $X2=2.685 $Y2=0.18
r153 21 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.61 $Y=0.255
+ $X2=2.61 $Y2=0.18
r154 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.61 $Y=0.255
+ $X2=2.61 $Y2=0.805
r155 19 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.535 $Y=0.18
+ $X2=2.61 $Y2=0.18
r156 19 20 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=2.535 $Y=0.18
+ $X2=1.67 $Y2=0.18
r157 17 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.195 $Y=3.15
+ $X2=3.27 $Y2=3.15
r158 17 18 820.426 $w=1.5e-07 $l=1.6e-06 $layer=POLY_cond $X=3.195 $Y=3.15
+ $X2=1.595 $Y2=3.15
r159 14 42 20.4101 $w=1.5e-07 $l=9.20598e-08 $layer=POLY_cond $X=1.595 $Y=1.43
+ $X2=1.557 $Y2=1.505
r160 14 16 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.595 $Y=1.43
+ $X2=1.595 $Y2=0.805
r161 13 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.595 $Y=0.255
+ $X2=1.67 $Y2=0.18
r162 13 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.595 $Y=0.255
+ $X2=1.595 $Y2=0.805
r163 10 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.52 $Y=3.075
+ $X2=1.595 $Y2=3.15
r164 10 12 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.52 $Y=3.075
+ $X2=1.52 $Y2=2.635
r165 9 42 20.4101 $w=1.5e-07 $l=9.16515e-08 $layer=POLY_cond $X=1.52 $Y=1.58
+ $X2=1.557 $Y2=1.505
r166 9 12 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=1.52 $Y=1.58
+ $X2=1.52 $Y2=2.635
r167 8 41 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.12 $Y=1.505
+ $X2=0.955 $Y2=1.58
r168 7 42 5.30422 $w=1.5e-07 $l=1.12e-07 $layer=POLY_cond $X=1.445 $Y=1.505
+ $X2=1.557 $Y2=1.505
r169 7 8 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.445 $Y=1.505
+ $X2=1.12 $Y2=1.505
r170 2 47 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.29 $X2=0.69 $Y2=2.445
r171 1 59 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.35 $X2=0.69 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%A_1169_93# 1 2 7 9 14 16 20 24 28 32 36 40
+ 44 47 48 49 50 53 54 56 57 60 63 65 66 71 75 80 81 84 86 98
c164 81 0 2.85281e-19 $X=7.27 $Y=1.35
c165 36 0 6.36774e-20 $X=10.035 $Y=2.465
c166 28 0 6.36774e-20 $X=9.605 $Y=2.465
r167 97 98 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=10.035 $Y=1.485
+ $X2=10.04 $Y2=1.485
r168 96 97 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=9.61 $Y=1.485
+ $X2=10.035 $Y2=1.485
r169 95 96 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=9.605 $Y=1.485
+ $X2=9.61 $Y2=1.485
r170 85 95 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=9.47 $Y=1.485
+ $X2=9.605 $Y2=1.485
r171 84 86 9.98442 $w=1.83e-07 $l=1.65e-07 $layer=LI1_cond $X=9.462 $Y=1.485
+ $X2=9.462 $Y2=1.32
r172 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.47
+ $Y=1.485 $X2=9.47 $Y2=1.485
r173 81 91 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.27 $Y=1.35 $X2=7.27
+ $Y2=1.44
r174 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.27
+ $Y=1.35 $X2=7.27 $Y2=1.35
r175 78 80 8.99792 $w=2.58e-07 $l=2.03e-07 $layer=LI1_cond $X=7.067 $Y=1.385
+ $X2=7.27 $Y2=1.385
r176 76 78 0.75352 $w=2.58e-07 $l=1.7e-08 $layer=LI1_cond $X=7.05 $Y=1.385
+ $X2=7.067 $Y2=1.385
r177 73 74 13.8993 $w=4.73e-07 $l=3.45e-07 $layer=LI1_cond $X=6.897 $Y=0.63
+ $X2=6.897 $Y2=0.975
r178 71 73 2.76987 $w=4.73e-07 $l=1.1e-07 $layer=LI1_cond $X=6.897 $Y=0.52
+ $X2=6.897 $Y2=0.63
r179 68 86 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.455 $Y=0.715
+ $X2=9.455 $Y2=1.32
r180 67 73 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=7.135 $Y=0.63
+ $X2=6.897 $Y2=0.63
r181 66 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.37 $Y=0.63
+ $X2=9.455 $Y2=0.715
r182 66 67 145.813 $w=1.68e-07 $l=2.235e-06 $layer=LI1_cond $X=9.37 $Y=0.63
+ $X2=7.135 $Y2=0.63
r183 65 75 4.07813 $w=2.37e-07 $l=1.04785e-07 $layer=LI1_cond $X=7.067 $Y=1.985
+ $X2=7.035 $Y2=2.075
r184 64 78 2.15511 $w=2.05e-07 $l=1.3e-07 $layer=LI1_cond $X=7.067 $Y=1.515
+ $X2=7.067 $Y2=1.385
r185 64 65 25.4279 $w=2.03e-07 $l=4.7e-07 $layer=LI1_cond $X=7.067 $Y=1.515
+ $X2=7.067 $Y2=1.985
r186 63 76 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.05 $Y=1.255
+ $X2=7.05 $Y2=1.385
r187 63 74 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.05 $Y=1.255
+ $X2=7.05 $Y2=0.975
r188 58 75 4.07813 $w=2.37e-07 $l=9e-08 $layer=LI1_cond $X=7.035 $Y=2.165
+ $X2=7.035 $Y2=2.075
r189 58 60 10.0305 $w=2.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.035 $Y=2.165
+ $X2=7.035 $Y2=2.4
r190 56 75 2.35733 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=6.9 $Y=2.075
+ $X2=7.035 $Y2=2.075
r191 56 57 35.4293 $w=1.78e-07 $l=5.75e-07 $layer=LI1_cond $X=6.9 $Y=2.075
+ $X2=6.325 $Y2=2.075
r192 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.16
+ $Y=1.59 $X2=6.16 $Y2=1.59
r193 51 57 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=6.16 $Y=1.985
+ $X2=6.325 $Y2=2.075
r194 51 53 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=6.16 $Y=1.985
+ $X2=6.16 $Y2=1.59
r195 48 54 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.16 $Y=1.93
+ $X2=6.16 $Y2=1.59
r196 48 49 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.93
+ $X2=6.16 $Y2=2.095
r197 47 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.425
+ $X2=6.16 $Y2=1.59
r198 42 44 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.92 $Y=1.2
+ $X2=6.07 $Y2=1.2
r199 38 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.04 $Y=1.32
+ $X2=10.04 $Y2=1.485
r200 38 40 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=10.04 $Y=1.32
+ $X2=10.04 $Y2=0.685
r201 34 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.035 $Y=1.65
+ $X2=10.035 $Y2=1.485
r202 34 36 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=10.035 $Y=1.65
+ $X2=10.035 $Y2=2.465
r203 30 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.61 $Y=1.32
+ $X2=9.61 $Y2=1.485
r204 30 32 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.61 $Y=1.32
+ $X2=9.61 $Y2=0.685
r205 26 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.605 $Y=1.65
+ $X2=9.605 $Y2=1.485
r206 26 28 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=9.605 $Y=1.65
+ $X2=9.605 $Y2=2.465
r207 22 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.925 $Y=1.515
+ $X2=7.925 $Y2=1.44
r208 22 24 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.925 $Y=1.515
+ $X2=7.925 $Y2=2.155
r209 18 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.925 $Y=1.365
+ $X2=7.925 $Y2=1.44
r210 18 20 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=7.925 $Y=1.365
+ $X2=7.925 $Y2=0.895
r211 17 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.435 $Y=1.44
+ $X2=7.27 $Y2=1.44
r212 16 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.85 $Y=1.44
+ $X2=7.925 $Y2=1.44
r213 16 17 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=7.85 $Y=1.44
+ $X2=7.435 $Y2=1.44
r214 14 49 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.22 $Y=2.465
+ $X2=6.22 $Y2=2.095
r215 10 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.07 $Y=1.275
+ $X2=6.07 $Y2=1.2
r216 10 47 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.07 $Y=1.275
+ $X2=6.07 $Y2=1.425
r217 7 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.92 $Y=1.125
+ $X2=5.92 $Y2=1.2
r218 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.92 $Y=1.125
+ $X2=5.92 $Y2=0.805
r219 2 60 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.865
+ $Y=2.255 $X2=7.005 $Y2=2.4
r220 1 71 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.685
+ $Y=0.375 $X2=6.825 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%A_982_369# 1 2 9 13 17 18 20 23 27 34 36 38
+ 39
c90 38 0 2.85281e-19 $X=6.7 $Y=1.31
r91 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.7 $Y=1.31
+ $X2=6.7 $Y2=1.31
r92 32 34 6.88026 $w=3.33e-07 $l=2e-07 $layer=LI1_cond $X=5.24 $Y=0.807 $X2=5.44
+ $Y2=0.807
r93 28 36 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.565 $Y=1.23
+ $X2=5.44 $Y2=1.23
r94 27 38 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.535 $Y=1.23
+ $X2=6.665 $Y2=1.23
r95 27 28 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=6.535 $Y=1.23
+ $X2=5.565 $Y2=1.23
r96 23 25 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=5.44 $Y=1.99
+ $X2=5.44 $Y2=2.54
r97 21 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=1.315
+ $X2=5.44 $Y2=1.23
r98 21 23 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.44 $Y=1.315
+ $X2=5.44 $Y2=1.99
r99 20 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=1.145
+ $X2=5.44 $Y2=1.23
r100 19 34 2.45311 $w=2.5e-07 $l=1.68e-07 $layer=LI1_cond $X=5.44 $Y=0.975
+ $X2=5.44 $Y2=0.807
r101 19 20 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.44 $Y=0.975
+ $X2=5.44 $Y2=1.145
r102 17 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.7 $Y=1.65 $X2=6.7
+ $Y2=1.31
r103 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=1.65
+ $X2=6.7 $Y2=1.815
r104 16 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=1.145
+ $X2=6.7 $Y2=1.31
r105 13 18 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.79 $Y=2.675
+ $X2=6.79 $Y2=1.815
r106 9 16 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.61 $Y=0.695
+ $X2=6.61 $Y2=1.145
r107 2 25 600 $w=1.7e-07 $l=9.0751e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.845 $X2=5.4 $Y2=2.54
r108 2 23 600 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.845 $X2=5.4 $Y2=1.99
r109 1 32 182 $w=1.7e-07 $l=3.23381e-07 $layer=licon1_NDIFF $count=1 $X=5.005
+ $Y=0.595 $X2=5.24 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%A_1513_137# 1 2 7 9 12 14 16 19 24 26 31 35
r64 34 35 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=8.59 $Y=1.38
+ $X2=9.02 $Y2=1.38
r65 29 34 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=8.375 $Y=1.38
+ $X2=8.59 $Y2=1.38
r66 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.375
+ $Y=1.38 $X2=8.375 $Y2=1.38
r67 26 28 11.6902 $w=6.94e-07 $l=6.65e-07 $layer=LI1_cond $X=7.71 $Y=1.26
+ $X2=8.375 $Y2=1.26
r68 24 31 7.7181 $w=3.25e-07 $l=1.65e-07 $layer=LI1_cond $X=7.71 $Y=1.815
+ $X2=7.71 $Y2=1.98
r69 23 26 7.89474 $w=2.1e-07 $l=3.65e-07 $layer=LI1_cond $X=7.71 $Y=1.625
+ $X2=7.71 $Y2=1.26
r70 23 24 10.0346 $w=2.08e-07 $l=1.9e-07 $layer=LI1_cond $X=7.71 $Y=1.625
+ $X2=7.71 $Y2=1.815
r71 17 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.02 $Y=1.545
+ $X2=9.02 $Y2=1.38
r72 17 19 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=9.02 $Y=1.545
+ $X2=9.02 $Y2=2.465
r73 14 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.02 $Y=1.215
+ $X2=9.02 $Y2=1.38
r74 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.02 $Y=1.215
+ $X2=9.02 $Y2=0.685
r75 10 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.59 $Y=1.545
+ $X2=8.59 $Y2=1.38
r76 10 12 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=8.59 $Y=1.545
+ $X2=8.59 $Y2=2.465
r77 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.59 $Y=1.215
+ $X2=8.59 $Y2=1.38
r78 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.59 $Y=1.215 $X2=8.59
+ $Y2=0.685
r79 2 31 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=7.585
+ $Y=1.835 $X2=7.71 $Y2=1.98
r80 1 26 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=7.565
+ $Y=0.685 $X2=7.71 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 42 48 52
+ 54 59 60 61 63 68 76 91 95 104 107 110 113 117
r111 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r112 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r113 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r115 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r117 99 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r118 99 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r119 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r120 96 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.48 $Y=3.33
+ $X2=9.315 $Y2=3.33
r121 96 98 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.48 $Y=3.33
+ $X2=9.84 $Y2=3.33
r122 95 116 4.31554 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=10.125 $Y=3.33
+ $X2=10.342 $Y2=3.33
r123 95 98 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.125 $Y=3.33
+ $X2=9.84 $Y2=3.33
r124 94 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r125 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r126 91 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.15 $Y=3.33
+ $X2=9.315 $Y2=3.33
r127 91 93 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.15 $Y=3.33
+ $X2=8.88 $Y2=3.33
r128 90 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r129 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r130 87 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 87 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r132 86 89 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r133 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r134 84 110 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=6.73 $Y=3.33
+ $X2=6.5 $Y2=3.33
r135 84 86 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.73 $Y=3.33
+ $X2=6.96 $Y2=3.33
r136 83 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r137 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r138 80 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r139 79 82 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=6
+ $Y2=3.33
r140 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r141 77 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.11 $Y2=3.33
r142 77 79 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 76 110 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=6.27 $Y=3.33
+ $X2=6.5 $Y2=3.33
r144 76 82 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.27 $Y=3.33 $X2=6
+ $Y2=3.33
r145 75 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r146 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r147 72 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r148 72 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r149 71 74 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r150 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r151 69 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=1.705 $Y2=3.33
r152 69 71 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=2.16 $Y2=3.33
r153 68 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=4.11 $Y2=3.33
r154 68 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=3.6 $Y2=3.33
r155 67 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r156 67 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r157 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r158 64 101 4.59118 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.202 $Y2=3.33
r159 64 66 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=1.2 $Y2=3.33
r160 63 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.58 $Y=3.33
+ $X2=1.705 $Y2=3.33
r161 63 66 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.58 $Y=3.33
+ $X2=1.2 $Y2=3.33
r162 61 83 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33 $X2=6
+ $Y2=3.33
r163 61 80 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.56 $Y2=3.33
r164 59 89 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.045 $Y=3.33
+ $X2=7.92 $Y2=3.33
r165 59 60 10.2049 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=8.045 $Y=3.33
+ $X2=8.257 $Y2=3.33
r166 58 93 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 58 60 10.2049 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=8.257 $Y2=3.33
r168 54 57 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=10.27 $Y=1.98
+ $X2=10.27 $Y2=2.95
r169 52 116 3.1223 $w=2.9e-07 $l=1.15521e-07 $layer=LI1_cond $X=10.27 $Y=3.245
+ $X2=10.342 $Y2=3.33
r170 52 57 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=10.27 $Y=3.245
+ $X2=10.27 $Y2=2.95
r171 48 51 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=9.315 $Y=1.985
+ $X2=9.315 $Y2=2.97
r172 46 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.315 $Y=3.245
+ $X2=9.315 $Y2=3.33
r173 46 51 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.315 $Y=3.245
+ $X2=9.315 $Y2=2.97
r174 42 45 11.2533 $w=4.23e-07 $l=4.15e-07 $layer=LI1_cond $X=8.257 $Y=1.98
+ $X2=8.257 $Y2=2.395
r175 40 60 1.63918 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=8.257 $Y=3.245
+ $X2=8.257 $Y2=3.33
r176 40 45 23.0489 $w=4.23e-07 $l=8.5e-07 $layer=LI1_cond $X=8.257 $Y=3.245
+ $X2=8.257 $Y2=2.395
r177 36 39 12.8708 $w=4.58e-07 $l=4.95e-07 $layer=LI1_cond $X=6.5 $Y=2.455
+ $X2=6.5 $Y2=2.95
r178 34 110 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=3.245
+ $X2=6.5 $Y2=3.33
r179 34 39 7.6705 $w=4.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.5 $Y=3.245
+ $X2=6.5 $Y2=2.95
r180 30 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=3.33
r181 30 32 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=2.67
r182 26 104 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=3.33
r183 26 28 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=2.805
r184 22 101 3.00801 $w=3.1e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.25 $Y=3.245
+ $X2=0.202 $Y2=3.33
r185 22 24 29.7405 $w=3.08e-07 $l=8e-07 $layer=LI1_cond $X=0.25 $Y=3.245
+ $X2=0.25 $Y2=2.445
r186 7 57 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=10.11
+ $Y=1.835 $X2=10.25 $Y2=2.95
r187 7 54 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.11
+ $Y=1.835 $X2=10.25 $Y2=1.98
r188 6 51 400 $w=1.7e-07 $l=1.24013e-06 $layer=licon1_PDIFF $count=1 $X=9.095
+ $Y=1.835 $X2=9.315 $Y2=2.97
r189 6 48 400 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_PDIFF $count=1 $X=9.095
+ $Y=1.835 $X2=9.315 $Y2=1.985
r190 5 45 300 $w=1.7e-07 $l=7.23602e-07 $layer=licon1_PDIFF $count=2 $X=8
+ $Y=1.835 $X2=8.375 $Y2=2.395
r191 5 42 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8
+ $Y=1.835 $X2=8.14 $Y2=1.98
r192 4 39 600 $w=1.7e-07 $l=8.2318e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=2.255 $X2=6.575 $Y2=2.95
r193 4 36 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=2.255 $X2=6.435 $Y2=2.455
r194 3 32 600 $w=1.7e-07 $l=4.65349e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=2.315 $X2=4.11 $Y2=2.67
r195 2 28 600 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=2.315 $X2=1.735 $Y2=2.805
r196 1 24 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.29 $X2=0.26 $Y2=2.445
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%A_429_119# 1 2 12 15 16
c24 15 0 1.58287e-19 $X=2.435 $Y=2.465
r25 15 16 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.472 $Y=2.465
+ $X2=2.472 $Y2=2.3
r26 10 12 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=0.79
+ $X2=2.51 $Y2=0.79
r27 7 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=0.955
+ $X2=2.51 $Y2=0.79
r28 7 16 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=2.51 $Y=0.955
+ $X2=2.51 $Y2=2.3
r29 2 15 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=2.315 $X2=2.435 $Y2=2.465
r30 1 10 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.595 $X2=2.345 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%Q_N 1 2 7 8 9 10 11 18
r19 11 32 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=8.805 $Y=2.775
+ $X2=8.805 $Y2=2.91
r20 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.805 $Y=2.405
+ $X2=8.805 $Y2=2.775
r21 9 10 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.805 $Y=1.96
+ $X2=8.805 $Y2=2.405
r22 8 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.805 $Y=1.665
+ $X2=8.805 $Y2=1.96
r23 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.805 $Y=1.295
+ $X2=8.805 $Y2=1.665
r24 7 18 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=8.805 $Y=1.295
+ $X2=8.805 $Y2=0.98
r25 2 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.665
+ $Y=1.835 $X2=8.805 $Y2=2.91
r26 2 9 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=8.665
+ $Y=1.835 $X2=8.805 $Y2=1.96
r27 1 18 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=8.665
+ $Y=0.265 $X2=8.805 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%Q 1 2 9 10 11 12 13 14 15 16 25
r22 16 43 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=9.845 $Y=2.775
+ $X2=9.845 $Y2=2.91
r23 15 16 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=9.845 $Y=2.405
+ $X2=9.845 $Y2=2.775
r24 14 15 23.3108 $w=2.18e-07 $l=4.45e-07 $layer=LI1_cond $X=9.845 $Y=1.96
+ $X2=9.845 $Y2=2.405
r25 13 14 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=9.845 $Y=1.665
+ $X2=9.845 $Y2=1.96
r26 12 13 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=9.845 $Y=1.295
+ $X2=9.845 $Y2=1.665
r27 10 11 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=9.837 $Y=0.555
+ $X2=9.837 $Y2=0.925
r28 10 25 6.62042 $w=2.33e-07 $l=1.35e-07 $layer=LI1_cond $X=9.837 $Y=0.555
+ $X2=9.837 $Y2=0.42
r29 9 12 8.11948 $w=2.18e-07 $l=1.55e-07 $layer=LI1_cond $X=9.845 $Y=1.14
+ $X2=9.845 $Y2=1.295
r30 7 11 4.80593 $w=2.33e-07 $l=9.8e-08 $layer=LI1_cond $X=9.837 $Y=1.023
+ $X2=9.837 $Y2=0.925
r31 7 9 5.80015 $w=2.33e-07 $l=1.17e-07 $layer=LI1_cond $X=9.837 $Y=1.023
+ $X2=9.837 $Y2=1.14
r32 2 43 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=2.91
r33 2 14 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=1.96
r34 1 25 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=9.685
+ $Y=0.265 $X2=9.825 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_2%VGND 1 2 3 4 5 6 7 22 24 28 32 34 36 38 39
+ 45 47 52 60 69 73 82 86 94 100 107
r108 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r109 100 103 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=9.315 $Y=0
+ $X2=9.315 $Y2=0.28
r110 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r111 95 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r112 94 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r113 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r114 87 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r115 86 91 10.2591 $w=8.78e-07 $l=7.4e-07 $layer=LI1_cond $X=3.915 $Y=0
+ $X2=3.915 $Y2=0.74
r116 86 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r117 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r118 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r119 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r120 77 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r121 77 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r122 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r123 74 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.48 $Y=0
+ $X2=9.315 $Y2=0
r124 74 76 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.48 $Y=0 $X2=9.84
+ $Y2=0
r125 73 106 4.36189 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=10.125 $Y=0
+ $X2=10.342 $Y2=0
r126 73 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.125 $Y=0
+ $X2=9.84 $Y2=0
r127 72 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r128 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r129 69 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.15 $Y=0
+ $X2=9.315 $Y2=0
r130 69 71 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.15 $Y=0 $X2=8.88
+ $Y2=0
r131 68 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r132 68 95 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=6.48 $Y2=0
r133 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r134 65 94 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=6.49 $Y=0 $X2=6.23
+ $Y2=0
r135 65 67 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=6.49 $Y=0 $X2=7.92
+ $Y2=0
r136 64 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r137 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r138 61 86 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=3.915
+ $Y2=0
r139 61 63 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.355 $Y=0
+ $X2=4.56 $Y2=0
r140 60 94 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=5.97 $Y=0 $X2=6.23
+ $Y2=0
r141 60 63 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=5.97 $Y=0 $X2=4.56
+ $Y2=0
r142 59 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r143 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r144 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r145 56 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r146 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r147 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r148 53 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.81
+ $Y2=0
r149 53 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=2.16 $Y2=0
r150 52 86 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.915
+ $Y2=0
r151 52 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.475 $Y=0
+ $X2=3.12 $Y2=0
r152 51 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r153 51 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r154 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r155 48 79 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r156 48 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r157 47 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=0 $X2=1.81
+ $Y2=0
r158 47 50 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.645 $Y=0
+ $X2=0.72 $Y2=0
r159 45 97 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=6
+ $Y2=0
r160 45 64 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=4.56
+ $Y2=0
r161 41 71 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=8.425 $Y=0
+ $X2=8.88 $Y2=0
r162 39 67 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=8.095 $Y=0
+ $X2=7.92 $Y2=0
r163 38 43 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=8.26 $Y=0 $X2=8.26
+ $Y2=0.28
r164 38 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.26 $Y=0 $X2=8.425
+ $Y2=0
r165 38 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.26 $Y=0 $X2=8.095
+ $Y2=0
r166 34 106 3.11564 $w=2.95e-07 $l=1.14782e-07 $layer=LI1_cond $X=10.272
+ $Y=0.085 $X2=10.342 $Y2=0
r167 34 36 12.6964 $w=2.93e-07 $l=3.25e-07 $layer=LI1_cond $X=10.272 $Y=0.085
+ $X2=10.272 $Y2=0.41
r168 30 94 2.17428 $w=5.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.23 $Y=0.085
+ $X2=6.23 $Y2=0
r169 30 32 10.0057 $w=5.18e-07 $l=4.35e-07 $layer=LI1_cond $X=6.23 $Y=0.085
+ $X2=6.23 $Y2=0.52
r170 26 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0
r171 26 28 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0.805
r172 22 79 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r173 22 24 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.555
r174 7 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.115
+ $Y=0.265 $X2=10.255 $Y2=0.41
r175 6 103 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=9.095
+ $Y=0.265 $X2=9.315 $Y2=0.28
r176 5 43 182 $w=1.7e-07 $l=5.18965e-07 $layer=licon1_NDIFF $count=1 $X=8
+ $Y=0.685 $X2=8.26 $Y2=0.28
r177 4 32 91 $w=1.7e-07 $l=4.3589e-07 $layer=licon1_NDIFF $count=2 $X=5.995
+ $Y=0.595 $X2=6.395 $Y2=0.52
r178 3 91 91 $w=1.7e-07 $l=7.59045e-07 $layer=licon1_NDIFF $count=2 $X=3.5
+ $Y=0.595 $X2=4.19 $Y2=0.74
r179 2 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.595 $X2=1.81 $Y2=0.805
r180 1 24 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.35 $X2=0.26 $Y2=0.555
.ends

