# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a211oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a211oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.730000 1.415000 4.715000 1.595000 ;
        RECT 4.445000 1.210000 4.715000 1.415000 ;
        RECT 4.445000 1.595000 4.715000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 1.415000 3.450000 1.595000 ;
        RECT 2.005000 1.595000 2.895000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 1.425000 1.835000 1.750000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.425000 1.750000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.125600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.255000 0.855000 1.075000 ;
        RECT 0.595000 1.075000 4.265000 1.245000 ;
        RECT 0.595000 1.245000 0.925000 2.735000 ;
        RECT 1.525000 0.255000 1.765000 1.075000 ;
        RECT 3.935000 0.595000 4.265000 1.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.165000  0.085000 0.425000 1.040000 ;
      RECT 0.165000  1.920000 0.425000 2.905000 ;
      RECT 0.165000  2.905000 2.215000 3.075000 ;
      RECT 1.025000  0.085000 1.355000 0.905000 ;
      RECT 1.095000  1.920000 1.285000 2.905000 ;
      RECT 1.455000  1.920000 4.115000 1.935000 ;
      RECT 1.455000  1.935000 3.255000 2.090000 ;
      RECT 1.455000  2.090000 1.785000 2.735000 ;
      RECT 1.935000  0.085000 2.215000 0.905000 ;
      RECT 1.955000  2.260000 2.215000 2.905000 ;
      RECT 2.405000  0.305000 2.735000 0.735000 ;
      RECT 2.405000  0.735000 3.755000 0.905000 ;
      RECT 2.565000  2.260000 2.895000 3.245000 ;
      RECT 2.915000  0.085000 3.245000 0.565000 ;
      RECT 3.065000  1.765000 4.115000 1.920000 ;
      RECT 3.065000  2.090000 3.255000 3.075000 ;
      RECT 3.425000  0.255000 4.695000 0.425000 ;
      RECT 3.425000  0.425000 3.755000 0.735000 ;
      RECT 3.425000  2.105000 3.755000 3.245000 ;
      RECT 3.925000  1.935000 4.115000 3.075000 ;
      RECT 4.285000  1.920000 4.615000 3.245000 ;
      RECT 4.435000  0.425000 4.695000 1.040000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__a211oi_2
END LIBRARY
