* File: sky130_fd_sc_lp__o32ai_0.spice
* Created: Wed Sep  2 10:26:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32ai_0.pex.spice"
.subckt sky130_fd_sc_lp__o32ai_0  VNB VPB B1 B2 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_33_82#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.1113 PD=0.77 PS=1.37 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_33_82#_M1000_d N_B2_M1000_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=0 M=1 R=2.8 SA=75000.7 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A3_M1002_g N_A_33_82#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.14175 AS=0.0588 PD=1.095 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_A_33_82#_M1005_d N_A2_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.14175 PD=0.7 PS=1.095 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A1_M1001_g N_A_33_82#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1006 A_133_491# N_B1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1728 PD=0.88 PS=1.82 NRD=19.9955 NRS=1.5366 M=1 R=4.26667
+ SA=75000.2 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1007 N_Y_M1007_d N_B2_M1007_g A_133_491# VPB PHIGHVT L=0.15 W=0.64 AD=0.1344
+ AS=0.0768 PD=1.06 PS=0.88 NRD=7.683 NRS=19.9955 M=1 R=4.26667 SA=75000.6
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1004 A_325_491# N_A3_M1004_g N_Y_M1007_d VPB PHIGHVT L=0.15 W=0.64 AD=0.1344
+ AS=0.1344 PD=1.06 PS=1.06 NRD=47.6937 NRS=35.3812 M=1 R=4.26667 SA=75001.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1008 A_439_491# N_A2_M1008_g A_325_491# VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.1344 PD=0.88 PS=1.06 NRD=19.9955 NRS=47.6937 M=1 R=4.26667 SA=75001.7
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_439_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75002.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o32ai_0.pxi.spice"
*
.ends
*
*
