* NGSPICE file created from sky130_fd_sc_lp__o31a_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o31a_0 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 a_270_55# A1 VGND VNB nshort w=420000u l=150000u
+  ad=2.688e+11p pd=2.96e+06u as=3.108e+11p ps=3.16e+06u
M1001 VPWR a_90_309# X VPB phighvt w=640000u l=150000u
+  ad=4.736e+11p pd=4.04e+06u as=1.696e+11p ps=1.81e+06u
M1002 a_354_481# A2 a_270_481# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.728e+11p ps=1.82e+06u
M1003 a_270_55# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_270_481# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_270_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B1 a_90_309# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.112e+11p ps=1.94e+06u
M1007 a_90_309# B1 a_270_55# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 VGND a_90_309# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 a_90_309# A3 a_354_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

