* File: sky130_fd_sc_lp__dlxtn_4.pxi.spice
* Created: Wed Sep  2 09:48:37 2020
* 
x_PM_SKY130_FD_SC_LP__DLXTN_4%D N_D_M1017_g N_D_M1007_g D D N_D_c_162_n
+ N_D_c_163_n PM_SKY130_FD_SC_LP__DLXTN_4%D
x_PM_SKY130_FD_SC_LP__DLXTN_4%GATE_N N_GATE_N_M1003_g N_GATE_N_c_194_n
+ N_GATE_N_M1008_g N_GATE_N_c_195_n N_GATE_N_c_196_n N_GATE_N_c_197_n
+ N_GATE_N_c_203_n N_GATE_N_c_198_n GATE_N GATE_N N_GATE_N_c_200_n
+ PM_SKY130_FD_SC_LP__DLXTN_4%GATE_N
x_PM_SKY130_FD_SC_LP__DLXTN_4%A_200_481# N_A_200_481#_M1008_d
+ N_A_200_481#_M1003_d N_A_200_481#_M1014_g N_A_200_481#_c_253_n
+ N_A_200_481#_M1023_g N_A_200_481#_M1012_g N_A_200_481#_M1005_g
+ N_A_200_481#_c_255_n N_A_200_481#_c_256_n N_A_200_481#_c_268_n
+ N_A_200_481#_c_257_n N_A_200_481#_c_269_n N_A_200_481#_c_270_n
+ N_A_200_481#_c_297_p N_A_200_481#_c_271_n N_A_200_481#_c_272_n
+ N_A_200_481#_c_258_n N_A_200_481#_c_259_n N_A_200_481#_c_260_n
+ N_A_200_481#_c_261_n N_A_200_481#_c_262_n N_A_200_481#_c_274_n
+ N_A_200_481#_c_263_n N_A_200_481#_c_264_n N_A_200_481#_c_265_n
+ PM_SKY130_FD_SC_LP__DLXTN_4%A_200_481#
x_PM_SKY130_FD_SC_LP__DLXTN_4%A_27_481# N_A_27_481#_M1007_s N_A_27_481#_M1017_s
+ N_A_27_481#_M1004_g N_A_27_481#_M1009_g N_A_27_481#_c_421_n
+ N_A_27_481#_c_427_n N_A_27_481#_c_422_n N_A_27_481#_c_429_n
+ N_A_27_481#_c_430_n N_A_27_481#_c_460_n N_A_27_481#_c_423_n
+ N_A_27_481#_c_424_n N_A_27_481#_c_431_n PM_SKY130_FD_SC_LP__DLXTN_4%A_27_481#
x_PM_SKY130_FD_SC_LP__DLXTN_4%A_310_485# N_A_310_485#_M1023_s
+ N_A_310_485#_M1014_s N_A_310_485#_M1020_g N_A_310_485#_c_502_n
+ N_A_310_485#_c_503_n N_A_310_485#_M1015_g N_A_310_485#_c_505_n
+ N_A_310_485#_c_514_n N_A_310_485#_c_506_n N_A_310_485#_c_507_n
+ N_A_310_485#_c_515_n N_A_310_485#_c_516_n N_A_310_485#_c_517_n
+ N_A_310_485#_c_521_n N_A_310_485#_c_508_n N_A_310_485#_c_509_n
+ N_A_310_485#_c_564_n N_A_310_485#_c_510_n N_A_310_485#_c_511_n
+ N_A_310_485#_c_512_n PM_SKY130_FD_SC_LP__DLXTN_4%A_310_485#
x_PM_SKY130_FD_SC_LP__DLXTN_4%A_795_423# N_A_795_423#_M1021_d
+ N_A_795_423#_M1002_d N_A_795_423#_M1013_g N_A_795_423#_M1022_g
+ N_A_795_423#_c_627_n N_A_795_423#_M1000_g N_A_795_423#_M1001_g
+ N_A_795_423#_M1010_g N_A_795_423#_M1006_g N_A_795_423#_M1016_g
+ N_A_795_423#_M1011_g N_A_795_423#_M1018_g N_A_795_423#_M1019_g
+ N_A_795_423#_c_651_n N_A_795_423#_c_636_n N_A_795_423#_c_637_n
+ N_A_795_423#_c_652_n N_A_795_423#_c_653_n N_A_795_423#_c_654_n
+ N_A_795_423#_c_638_n N_A_795_423#_c_655_n N_A_795_423#_c_639_n
+ N_A_795_423#_c_640_n N_A_795_423#_c_718_p N_A_795_423#_c_641_n
+ N_A_795_423#_c_642_n N_A_795_423#_c_658_n N_A_795_423#_c_643_n
+ N_A_795_423#_c_644_n N_A_795_423#_c_645_n
+ PM_SKY130_FD_SC_LP__DLXTN_4%A_795_423#
x_PM_SKY130_FD_SC_LP__DLXTN_4%A_609_485# N_A_609_485#_M1012_d
+ N_A_609_485#_M1020_d N_A_609_485#_c_790_n N_A_609_485#_M1021_g
+ N_A_609_485#_M1002_g N_A_609_485#_c_799_n N_A_609_485#_c_815_n
+ N_A_609_485#_c_792_n N_A_609_485#_c_793_n N_A_609_485#_c_794_n
+ N_A_609_485#_c_795_n N_A_609_485#_c_796_n N_A_609_485#_c_797_n
+ PM_SKY130_FD_SC_LP__DLXTN_4%A_609_485#
x_PM_SKY130_FD_SC_LP__DLXTN_4%VPWR N_VPWR_M1017_d N_VPWR_M1014_d N_VPWR_M1013_d
+ N_VPWR_M1001_d N_VPWR_M1006_d N_VPWR_M1019_d N_VPWR_c_891_n N_VPWR_c_892_n
+ N_VPWR_c_893_n N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n N_VPWR_c_897_n
+ N_VPWR_c_898_n N_VPWR_c_899_n N_VPWR_c_900_n N_VPWR_c_962_n N_VPWR_c_901_n
+ N_VPWR_c_902_n VPWR N_VPWR_c_903_n N_VPWR_c_904_n N_VPWR_c_905_n
+ N_VPWR_c_906_n N_VPWR_c_907_n N_VPWR_c_908_n N_VPWR_c_909_n N_VPWR_c_890_n
+ PM_SKY130_FD_SC_LP__DLXTN_4%VPWR
x_PM_SKY130_FD_SC_LP__DLXTN_4%Q N_Q_M1000_s N_Q_M1016_s N_Q_M1001_s N_Q_M1011_s
+ N_Q_c_1050_p N_Q_c_1038_n N_Q_c_1004_n N_Q_c_1005_n N_Q_c_1008_n N_Q_c_1009_n
+ Q Q Q Q N_Q_c_1051_p Q Q PM_SKY130_FD_SC_LP__DLXTN_4%Q
x_PM_SKY130_FD_SC_LP__DLXTN_4%VGND N_VGND_M1007_d N_VGND_M1023_d N_VGND_M1022_d
+ N_VGND_M1000_d N_VGND_M1010_d N_VGND_M1018_d N_VGND_c_1056_n N_VGND_c_1057_n
+ N_VGND_c_1058_n N_VGND_c_1059_n N_VGND_c_1060_n N_VGND_c_1061_n
+ N_VGND_c_1062_n N_VGND_c_1063_n N_VGND_c_1064_n VGND N_VGND_c_1065_n
+ N_VGND_c_1066_n N_VGND_c_1067_n N_VGND_c_1068_n N_VGND_c_1069_n
+ N_VGND_c_1070_n N_VGND_c_1071_n N_VGND_c_1072_n N_VGND_c_1073_n
+ PM_SKY130_FD_SC_LP__DLXTN_4%VGND
cc_1 VNB N_D_M1017_g 0.00806231f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.725
cc_2 VNB D 0.00932086f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_3 VNB N_D_c_162_n 0.0326421f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_4 VNB N_D_c_163_n 0.0219202f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.19
cc_5 VNB N_GATE_N_c_194_n 0.0174454f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.19
cc_6 VNB N_GATE_N_c_195_n 0.0213631f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_7 VNB N_GATE_N_c_196_n 0.0281964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_GATE_N_c_197_n 0.0350463f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_9 VNB N_GATE_N_c_198_n 0.0041128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB GATE_N 0.0142852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_GATE_N_c_200_n 0.0449125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_200_481#_M1014_g 0.00758528f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_13 VNB N_A_200_481#_c_253_n 0.0187337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_200_481#_M1012_g 0.0223999f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.52
cc_15 VNB N_A_200_481#_c_255_n 0.0368194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_200_481#_c_256_n 0.0178494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_200_481#_c_257_n 0.0083363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_200_481#_c_258_n 0.0135386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_200_481#_c_259_n 0.00160541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_200_481#_c_260_n 0.0026905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_200_481#_c_261_n 0.00530849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_200_481#_c_262_n 2.6117e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_200_481#_c_263_n 0.0108106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_200_481#_c_264_n 0.0320123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_200_481#_c_265_n 0.0286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_481#_M1009_g 0.0312553f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_27 VNB N_A_27_481#_c_421_n 0.0161217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_481#_c_422_n 0.0304633f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.355
cc_29 VNB N_A_27_481#_c_423_n 0.0458138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_481#_c_424_n 0.0160375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_310_485#_c_502_n 0.0348062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_310_485#_c_503_n 0.0142475f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_33 VNB N_A_310_485#_M1015_g 0.0198893f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.19
cc_34 VNB N_A_310_485#_c_505_n 0.00989603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_310_485#_c_506_n 0.0131637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_310_485#_c_507_n 0.0190857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_310_485#_c_508_n 0.00751184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_310_485#_c_509_n 0.00169266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_310_485#_c_510_n 0.00106943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_310_485#_c_511_n 0.00100838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_310_485#_c_512_n 0.016938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_795_423#_M1022_g 0.0459975f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.355
cc_43 VNB N_A_795_423#_c_627_n 0.00574572f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.19
cc_44 VNB N_A_795_423#_M1000_g 0.0245299f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.355
cc_45 VNB N_A_795_423#_M1001_g 0.00359468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_795_423#_M1010_g 0.0191829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_795_423#_M1006_g 0.00299719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_795_423#_M1016_g 0.0191586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_795_423#_M1011_g 0.0029813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_795_423#_M1018_g 0.027939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_795_423#_M1019_g 0.00472897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_795_423#_c_636_n 0.0108569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_795_423#_c_637_n 4.3079e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_795_423#_c_638_n 0.0115241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_795_423#_c_639_n 0.00454897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_795_423#_c_640_n 5.6438e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_795_423#_c_641_n 0.00682967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_795_423#_c_642_n 0.00722737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_795_423#_c_643_n 0.00109702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_795_423#_c_644_n 0.0462935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_795_423#_c_645_n 0.0868295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_609_485#_c_790_n 0.0207063f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.87
cc_63 VNB N_A_609_485#_M1002_g 0.00375148f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.355
cc_64 VNB N_A_609_485#_c_792_n 0.00442499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_609_485#_c_793_n 0.00440375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_609_485#_c_794_n 0.0109329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_609_485#_c_795_n 8.95292e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_609_485#_c_796_n 0.0118444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_609_485#_c_797_n 0.0350453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VPWR_c_890_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_Q_c_1004_n 0.00315163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_Q_c_1005_n 0.00292432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB Q 0.00100033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB Q 0.0027949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1056_n 0.023702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1057_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1058_n 0.00240575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1059_n 0.00666504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1060_n 3.22151e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1061_n 0.0125262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1062_n 0.0143133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1063_n 0.020823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1064_n 0.00471252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1065_n 0.0378138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1066_n 0.0413193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1067_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1068_n 0.0149772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1069_n 0.0256782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1070_n 0.00436092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1071_n 0.00365101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1072_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1073_n 0.397671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VPB N_D_M1017_g 0.0566206f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.725
cc_94 VPB N_GATE_N_M1003_g 0.0473134f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.725
cc_95 VPB N_GATE_N_c_195_n 0.00742177f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_96 VPB N_GATE_N_c_203_n 0.015799f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.52
cc_97 VPB N_A_200_481#_M1014_g 0.0688238f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_98 VPB N_A_200_481#_M1005_g 0.0222645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_200_481#_c_268_n 0.00968559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_200_481#_c_269_n 0.0143465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_200_481#_c_270_n 0.00287821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_200_481#_c_271_n 0.0139643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_200_481#_c_272_n 0.00138828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_200_481#_c_262_n 0.00434506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_200_481#_c_274_n 0.0334648f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_27_481#_M1004_g 0.0372644f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_107 VPB N_A_27_481#_c_421_n 0.00855093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_27_481#_c_427_n 0.0156149f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.355
cc_109 VPB N_A_27_481#_c_422_n 0.00217356f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.355
cc_110 VPB N_A_27_481#_c_429_n 0.0573078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_27_481#_c_430_n 0.0435423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_27_481#_c_431_n 0.0129748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_310_485#_M1020_g 0.0217728f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_114 VPB N_A_310_485#_c_514_n 0.0143399f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.355
cc_115 VPB N_A_310_485#_c_515_n 0.00840856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_310_485#_c_516_n 0.0229652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_310_485#_c_517_n 0.00576856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_310_485#_c_510_n 0.0315209f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_795_423#_M1013_g 0.0209238f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_120 VPB N_A_795_423#_M1001_g 0.024097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_795_423#_M1006_g 0.0183095f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_795_423#_M1011_g 0.0185006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_795_423#_M1019_g 0.0265273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_795_423#_c_651_n 0.0321968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_795_423#_c_652_n 0.00194828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_795_423#_c_653_n 0.0284836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_795_423#_c_654_n 0.00672635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_795_423#_c_655_n 0.0139987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_795_423#_c_640_n 0.00192872f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_795_423#_c_641_n 0.0103257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_795_423#_c_658_n 0.00378347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_795_423#_c_644_n 0.00707719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_609_485#_M1002_g 0.0257386f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.355
cc_134 VPB N_A_609_485#_c_799_n 0.0063368f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.355
cc_135 VPB N_A_609_485#_c_792_n 0.0092649f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_891_n 0.0105698f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.355
cc_137 VPB N_VPWR_c_892_n 0.00320896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_893_n 0.0136071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_894_n 0.00408426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_895_n 0.0174344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_896_n 0.00191385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_897_n 0.0102066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_898_n 0.0643353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_899_n 0.0352338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_900_n 0.00398926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_901_n 0.0169585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_902_n 0.00545601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_903_n 0.0177231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_904_n 0.0412666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_905_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_906_n 0.0149952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_907_n 0.00487897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_908_n 0.0130242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_909_n 0.0044352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_890_n 0.0845347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_Q_c_1008_n 0.0027739f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_Q_c_1009_n 0.0035848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB Q 5.4375e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB Q 0.00169322f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 N_D_c_163_n N_GATE_N_c_194_n 0.0102856f $X=0.525 $Y=1.19 $X2=0 $Y2=0
cc_161 N_D_M1017_g N_GATE_N_c_195_n 0.00850309f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_162 D N_GATE_N_c_195_n 0.00979217f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_163 D N_GATE_N_c_196_n 0.0108662f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_164 N_D_M1017_g N_GATE_N_c_203_n 0.0353738f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_165 D N_GATE_N_c_203_n 4.97108e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_166 D N_GATE_N_c_198_n 0.00977717f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_167 N_D_c_162_n N_GATE_N_c_198_n 0.0181282f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_168 D N_A_200_481#_c_257_n 0.0142357f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_169 D N_A_200_481#_c_263_n 0.015415f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_170 D N_A_200_481#_c_264_n 0.0011362f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_171 N_D_M1017_g N_A_27_481#_c_422_n 0.006195f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_172 D N_A_27_481#_c_422_n 0.0262102f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_173 N_D_c_162_n N_A_27_481#_c_422_n 0.00806477f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_174 N_D_c_163_n N_A_27_481#_c_422_n 0.00522007f $X=0.525 $Y=1.19 $X2=0 $Y2=0
cc_175 N_D_M1017_g N_A_27_481#_c_429_n 0.0231158f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_176 N_D_M1017_g N_A_27_481#_c_430_n 0.0174815f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_177 D N_A_27_481#_c_430_n 0.062569f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_178 N_D_c_162_n N_A_27_481#_c_430_n 0.00326718f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_179 N_D_c_162_n N_A_27_481#_c_424_n 0.00365478f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_180 N_D_c_162_n N_A_27_481#_c_431_n 0.0021982f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_181 N_D_M1017_g N_VPWR_c_891_n 0.00305293f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_182 N_D_M1017_g N_VPWR_c_903_n 0.0053602f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_183 N_D_M1017_g N_VPWR_c_890_n 0.0108605f $X=0.495 $Y=2.725 $X2=0 $Y2=0
cc_184 D N_VGND_c_1056_n 0.0183063f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_185 N_D_c_162_n N_VGND_c_1056_n 0.00100132f $X=0.525 $Y=1.355 $X2=0 $Y2=0
cc_186 N_D_c_163_n N_VGND_c_1056_n 0.00353747f $X=0.525 $Y=1.19 $X2=0 $Y2=0
cc_187 N_D_c_163_n N_VGND_c_1069_n 0.00397346f $X=0.525 $Y=1.19 $X2=0 $Y2=0
cc_188 N_D_c_163_n N_VGND_c_1073_n 0.00459866f $X=0.525 $Y=1.19 $X2=0 $Y2=0
cc_189 N_GATE_N_c_197_n N_A_200_481#_c_253_n 0.00177483f $X=1.495 $Y=1.19 $X2=0
+ $Y2=0
cc_190 N_GATE_N_c_200_n N_A_200_481#_c_253_n 0.00338013f $X=1.585 $Y=0.365 $X2=0
+ $Y2=0
cc_191 N_GATE_N_c_197_n N_A_200_481#_c_255_n 0.0153552f $X=1.495 $Y=1.19 $X2=0
+ $Y2=0
cc_192 GATE_N N_A_200_481#_c_255_n 9.94013e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_193 N_GATE_N_M1003_g N_A_200_481#_c_268_n 2.34164e-19 $X=0.925 $Y=2.725 $X2=0
+ $Y2=0
cc_194 N_GATE_N_c_203_n N_A_200_481#_c_268_n 0.00162482f $X=1.005 $Y=1.835 $X2=0
+ $Y2=0
cc_195 N_GATE_N_c_194_n N_A_200_481#_c_257_n 0.00258368f $X=1.005 $Y=1.19 $X2=0
+ $Y2=0
cc_196 N_GATE_N_c_196_n N_A_200_481#_c_257_n 0.00373396f $X=1.42 $Y=1.265 $X2=0
+ $Y2=0
cc_197 N_GATE_N_c_197_n N_A_200_481#_c_257_n 0.0153809f $X=1.495 $Y=1.19 $X2=0
+ $Y2=0
cc_198 GATE_N N_A_200_481#_c_257_n 0.046537f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_199 N_GATE_N_c_200_n N_A_200_481#_c_257_n 6.55474e-19 $X=1.585 $Y=0.365 $X2=0
+ $Y2=0
cc_200 N_GATE_N_M1003_g N_A_200_481#_c_270_n 7.32615e-19 $X=0.925 $Y=2.725 $X2=0
+ $Y2=0
cc_201 N_GATE_N_c_195_n N_A_200_481#_c_263_n 0.0011026f $X=1.005 $Y=1.76 $X2=0
+ $Y2=0
cc_202 N_GATE_N_c_197_n N_A_200_481#_c_263_n 0.00668367f $X=1.495 $Y=1.19 $X2=0
+ $Y2=0
cc_203 GATE_N N_A_200_481#_c_263_n 0.0128992f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_204 N_GATE_N_c_200_n N_A_200_481#_c_263_n 3.23921e-19 $X=1.585 $Y=0.365 $X2=0
+ $Y2=0
cc_205 N_GATE_N_c_196_n N_A_200_481#_c_264_n 0.0153552f $X=1.42 $Y=1.265 $X2=0
+ $Y2=0
cc_206 N_GATE_N_c_195_n N_A_27_481#_c_430_n 0.0051607f $X=1.005 $Y=1.76 $X2=0
+ $Y2=0
cc_207 N_GATE_N_c_196_n N_A_27_481#_c_430_n 0.0103761f $X=1.42 $Y=1.265 $X2=0
+ $Y2=0
cc_208 N_GATE_N_c_203_n N_A_27_481#_c_430_n 0.0160606f $X=1.005 $Y=1.835 $X2=0
+ $Y2=0
cc_209 N_GATE_N_M1003_g N_A_310_485#_c_515_n 0.00483989f $X=0.925 $Y=2.725 $X2=0
+ $Y2=0
cc_210 N_GATE_N_M1003_g N_A_310_485#_c_517_n 0.00479618f $X=0.925 $Y=2.725 $X2=0
+ $Y2=0
cc_211 N_GATE_N_c_197_n N_A_310_485#_c_521_n 2.19257e-19 $X=1.495 $Y=1.19 $X2=0
+ $Y2=0
cc_212 GATE_N N_A_310_485#_c_521_n 0.0266316f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_213 N_GATE_N_c_200_n N_A_310_485#_c_521_n 0.00133992f $X=1.585 $Y=0.365 $X2=0
+ $Y2=0
cc_214 N_GATE_N_c_197_n N_A_310_485#_c_509_n 0.00284979f $X=1.495 $Y=1.19 $X2=0
+ $Y2=0
cc_215 GATE_N N_A_310_485#_c_509_n 0.00203396f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_216 N_GATE_N_M1003_g N_VPWR_c_891_n 0.00264084f $X=0.925 $Y=2.725 $X2=0 $Y2=0
cc_217 N_GATE_N_M1003_g N_VPWR_c_899_n 0.0053602f $X=0.925 $Y=2.725 $X2=0 $Y2=0
cc_218 N_GATE_N_M1003_g N_VPWR_c_890_n 0.0111156f $X=0.925 $Y=2.725 $X2=0 $Y2=0
cc_219 N_GATE_N_c_194_n N_VGND_c_1056_n 0.00117505f $X=1.005 $Y=1.19 $X2=0 $Y2=0
cc_220 GATE_N N_VGND_c_1056_n 0.031333f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_221 N_GATE_N_c_200_n N_VGND_c_1056_n 0.00253261f $X=1.585 $Y=0.365 $X2=0
+ $Y2=0
cc_222 N_GATE_N_c_200_n N_VGND_c_1057_n 2.99742e-19 $X=1.585 $Y=0.365 $X2=0
+ $Y2=0
cc_223 N_GATE_N_c_194_n N_VGND_c_1065_n 0.00339706f $X=1.005 $Y=1.19 $X2=0 $Y2=0
cc_224 GATE_N N_VGND_c_1065_n 0.0454564f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_225 N_GATE_N_c_200_n N_VGND_c_1065_n 0.006386f $X=1.585 $Y=0.365 $X2=0 $Y2=0
cc_226 N_GATE_N_c_194_n N_VGND_c_1073_n 0.00383222f $X=1.005 $Y=1.19 $X2=0 $Y2=0
cc_227 GATE_N N_VGND_c_1073_n 0.0282868f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_228 N_GATE_N_c_200_n N_VGND_c_1073_n 0.00915883f $X=1.585 $Y=0.365 $X2=0
+ $Y2=0
cc_229 N_A_200_481#_M1014_g N_A_27_481#_M1004_g 0.0206332f $X=1.91 $Y=2.745
+ $X2=0 $Y2=0
cc_230 N_A_200_481#_c_269_n N_A_27_481#_M1004_g 3.4075e-19 $X=1.96 $Y=2.99 $X2=0
+ $Y2=0
cc_231 N_A_200_481#_c_297_p N_A_27_481#_M1004_g 0.00283231f $X=2.045 $Y=2.905
+ $X2=0 $Y2=0
cc_232 N_A_200_481#_c_271_n N_A_27_481#_M1004_g 0.0126793f $X=3.435 $Y=2.485
+ $X2=0 $Y2=0
cc_233 N_A_200_481#_c_253_n N_A_27_481#_M1009_g 0.0238735f $X=2.365 $Y=0.77
+ $X2=0 $Y2=0
cc_234 N_A_200_481#_M1012_g N_A_27_481#_M1009_g 0.0361902f $X=3.155 $Y=0.445
+ $X2=0 $Y2=0
cc_235 N_A_200_481#_c_258_n N_A_27_481#_M1009_g 0.00765553f $X=3.08 $Y=1.055
+ $X2=0 $Y2=0
cc_236 N_A_200_481#_c_264_n N_A_27_481#_M1009_g 0.00319845f $X=1.975 $Y=1.06
+ $X2=0 $Y2=0
cc_237 N_A_200_481#_M1014_g N_A_27_481#_c_421_n 0.0133504f $X=1.91 $Y=2.745
+ $X2=0 $Y2=0
cc_238 N_A_200_481#_c_256_n N_A_27_481#_c_421_n 0.00876245f $X=1.975 $Y=1.565
+ $X2=0 $Y2=0
cc_239 N_A_200_481#_M1014_g N_A_27_481#_c_430_n 0.0134931f $X=1.91 $Y=2.745
+ $X2=0 $Y2=0
cc_240 N_A_200_481#_c_256_n N_A_27_481#_c_430_n 0.00494514f $X=1.975 $Y=1.565
+ $X2=0 $Y2=0
cc_241 N_A_200_481#_c_268_n N_A_27_481#_c_430_n 0.0114149f $X=1.14 $Y=2.56 $X2=0
+ $Y2=0
cc_242 N_A_200_481#_c_258_n N_A_27_481#_c_430_n 0.00715569f $X=3.08 $Y=1.055
+ $X2=0 $Y2=0
cc_243 N_A_200_481#_c_263_n N_A_27_481#_c_430_n 0.0353941f $X=1.917 $Y=1.055
+ $X2=0 $Y2=0
cc_244 N_A_200_481#_M1014_g N_A_27_481#_c_460_n 7.85937e-19 $X=1.91 $Y=2.745
+ $X2=0 $Y2=0
cc_245 N_A_200_481#_c_256_n N_A_27_481#_c_460_n 2.48769e-19 $X=1.975 $Y=1.565
+ $X2=0 $Y2=0
cc_246 N_A_200_481#_c_258_n N_A_27_481#_c_460_n 0.0253742f $X=3.08 $Y=1.055
+ $X2=0 $Y2=0
cc_247 N_A_200_481#_c_260_n N_A_27_481#_c_460_n 4.22635e-19 $X=3.245 $Y=1.325
+ $X2=0 $Y2=0
cc_248 N_A_200_481#_c_261_n N_A_27_481#_c_460_n 0.00746397f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_249 N_A_200_481#_c_263_n N_A_27_481#_c_460_n 0.0136767f $X=1.917 $Y=1.055
+ $X2=0 $Y2=0
cc_250 N_A_200_481#_c_264_n N_A_27_481#_c_460_n 2.71033e-19 $X=1.975 $Y=1.06
+ $X2=0 $Y2=0
cc_251 N_A_200_481#_c_255_n N_A_27_481#_c_423_n 0.00261354f $X=2.365 $Y=0.845
+ $X2=0 $Y2=0
cc_252 N_A_200_481#_c_258_n N_A_27_481#_c_423_n 0.0177929f $X=3.08 $Y=1.055
+ $X2=0 $Y2=0
cc_253 N_A_200_481#_c_260_n N_A_27_481#_c_423_n 0.00394613f $X=3.245 $Y=1.325
+ $X2=0 $Y2=0
cc_254 N_A_200_481#_c_261_n N_A_27_481#_c_423_n 0.00328054f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_255 N_A_200_481#_c_263_n N_A_27_481#_c_423_n 0.00185634f $X=1.917 $Y=1.055
+ $X2=0 $Y2=0
cc_256 N_A_200_481#_c_264_n N_A_27_481#_c_423_n 0.0135117f $X=1.975 $Y=1.06
+ $X2=0 $Y2=0
cc_257 N_A_200_481#_c_265_n N_A_27_481#_c_423_n 0.0361902f $X=3.245 $Y=1.06
+ $X2=0 $Y2=0
cc_258 N_A_200_481#_c_269_n N_A_310_485#_M1014_s 0.00334776f $X=1.96 $Y=2.99
+ $X2=0 $Y2=0
cc_259 N_A_200_481#_M1005_g N_A_310_485#_M1020_g 0.0174045f $X=3.51 $Y=2.635
+ $X2=0 $Y2=0
cc_260 N_A_200_481#_c_271_n N_A_310_485#_M1020_g 0.0121065f $X=3.435 $Y=2.485
+ $X2=0 $Y2=0
cc_261 N_A_200_481#_c_262_n N_A_310_485#_M1020_g 7.77208e-19 $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_262 N_A_200_481#_c_261_n N_A_310_485#_c_502_n 0.014018f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_263 N_A_200_481#_c_262_n N_A_310_485#_c_502_n 0.0141749f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_264 N_A_200_481#_c_274_n N_A_310_485#_c_502_n 0.0192032f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_265 N_A_200_481#_c_258_n N_A_310_485#_c_503_n 0.00401531f $X=3.08 $Y=1.055
+ $X2=0 $Y2=0
cc_266 N_A_200_481#_c_260_n N_A_310_485#_c_503_n 3.13573e-19 $X=3.245 $Y=1.325
+ $X2=0 $Y2=0
cc_267 N_A_200_481#_c_261_n N_A_310_485#_c_503_n 0.00314455f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_268 N_A_200_481#_c_265_n N_A_310_485#_c_503_n 0.016063f $X=3.245 $Y=1.06
+ $X2=0 $Y2=0
cc_269 N_A_200_481#_M1012_g N_A_310_485#_M1015_g 0.0204508f $X=3.155 $Y=0.445
+ $X2=0 $Y2=0
cc_270 N_A_200_481#_c_261_n N_A_310_485#_c_505_n 0.00541036f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_271 N_A_200_481#_M1005_g N_A_310_485#_c_514_n 0.0119074f $X=3.51 $Y=2.635
+ $X2=0 $Y2=0
cc_272 N_A_200_481#_c_271_n N_A_310_485#_c_514_n 0.00495015f $X=3.435 $Y=2.485
+ $X2=0 $Y2=0
cc_273 N_A_200_481#_c_262_n N_A_310_485#_c_514_n 3.22261e-19 $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_274 N_A_200_481#_c_260_n N_A_310_485#_c_506_n 5.63705e-19 $X=3.245 $Y=1.325
+ $X2=0 $Y2=0
cc_275 N_A_200_481#_c_260_n N_A_310_485#_c_507_n 0.0027898f $X=3.245 $Y=1.325
+ $X2=0 $Y2=0
cc_276 N_A_200_481#_c_261_n N_A_310_485#_c_507_n 0.00187868f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_277 N_A_200_481#_M1014_g N_A_310_485#_c_515_n 0.00784864f $X=1.91 $Y=2.745
+ $X2=0 $Y2=0
cc_278 N_A_200_481#_c_268_n N_A_310_485#_c_515_n 0.0226279f $X=1.14 $Y=2.56
+ $X2=0 $Y2=0
cc_279 N_A_200_481#_c_269_n N_A_310_485#_c_515_n 0.0188656f $X=1.96 $Y=2.99
+ $X2=0 $Y2=0
cc_280 N_A_200_481#_c_272_n N_A_310_485#_c_515_n 0.00776157f $X=2.13 $Y=2.485
+ $X2=0 $Y2=0
cc_281 N_A_200_481#_M1014_g N_A_310_485#_c_516_n 0.0168084f $X=1.91 $Y=2.745
+ $X2=0 $Y2=0
cc_282 N_A_200_481#_c_271_n N_A_310_485#_c_516_n 0.0783668f $X=3.435 $Y=2.485
+ $X2=0 $Y2=0
cc_283 N_A_200_481#_c_272_n N_A_310_485#_c_516_n 0.0135705f $X=2.13 $Y=2.485
+ $X2=0 $Y2=0
cc_284 N_A_200_481#_c_262_n N_A_310_485#_c_516_n 0.0111889f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_285 N_A_200_481#_c_274_n N_A_310_485#_c_516_n 5.83169e-19 $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_286 N_A_200_481#_c_253_n N_A_310_485#_c_508_n 0.00908285f $X=2.365 $Y=0.77
+ $X2=0 $Y2=0
cc_287 N_A_200_481#_M1012_g N_A_310_485#_c_508_n 0.0117899f $X=3.155 $Y=0.445
+ $X2=0 $Y2=0
cc_288 N_A_200_481#_c_255_n N_A_310_485#_c_508_n 0.00336563f $X=2.365 $Y=0.845
+ $X2=0 $Y2=0
cc_289 N_A_200_481#_c_258_n N_A_310_485#_c_508_n 0.0619255f $X=3.08 $Y=1.055
+ $X2=0 $Y2=0
cc_290 N_A_200_481#_c_259_n N_A_310_485#_c_508_n 0.0245354f $X=3.245 $Y=1.145
+ $X2=0 $Y2=0
cc_291 N_A_200_481#_c_261_n N_A_310_485#_c_508_n 0.00722733f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_292 N_A_200_481#_c_265_n N_A_310_485#_c_508_n 0.0043813f $X=3.245 $Y=1.06
+ $X2=0 $Y2=0
cc_293 N_A_200_481#_c_255_n N_A_310_485#_c_509_n 0.00771163f $X=2.365 $Y=0.845
+ $X2=0 $Y2=0
cc_294 N_A_200_481#_c_258_n N_A_310_485#_c_509_n 0.00744773f $X=3.08 $Y=1.055
+ $X2=0 $Y2=0
cc_295 N_A_200_481#_c_263_n N_A_310_485#_c_509_n 0.00861306f $X=1.917 $Y=1.055
+ $X2=0 $Y2=0
cc_296 N_A_200_481#_c_258_n N_A_310_485#_c_564_n 0.00610558f $X=3.08 $Y=1.055
+ $X2=0 $Y2=0
cc_297 N_A_200_481#_c_261_n N_A_310_485#_c_564_n 0.0102831f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_298 N_A_200_481#_c_262_n N_A_310_485#_c_564_n 0.0241401f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_299 N_A_200_481#_c_274_n N_A_310_485#_c_564_n 5.91458e-19 $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_300 N_A_200_481#_c_262_n N_A_310_485#_c_510_n 0.00663493f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_301 N_A_200_481#_c_274_n N_A_310_485#_c_510_n 0.0119074f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_302 N_A_200_481#_M1012_g N_A_310_485#_c_511_n 6.85545e-19 $X=3.155 $Y=0.445
+ $X2=0 $Y2=0
cc_303 N_A_200_481#_c_259_n N_A_310_485#_c_511_n 0.00670294f $X=3.245 $Y=1.145
+ $X2=0 $Y2=0
cc_304 N_A_200_481#_c_261_n N_A_310_485#_c_511_n 0.00386575f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_305 N_A_200_481#_c_265_n N_A_310_485#_c_511_n 6.25161e-19 $X=3.245 $Y=1.06
+ $X2=0 $Y2=0
cc_306 N_A_200_481#_c_259_n N_A_310_485#_c_512_n 9.10309e-19 $X=3.245 $Y=1.145
+ $X2=0 $Y2=0
cc_307 N_A_200_481#_c_265_n N_A_310_485#_c_512_n 0.0214051f $X=3.245 $Y=1.06
+ $X2=0 $Y2=0
cc_308 N_A_200_481#_c_271_n N_A_795_423#_M1013_g 5.68128e-19 $X=3.435 $Y=2.485
+ $X2=0 $Y2=0
cc_309 N_A_200_481#_M1005_g N_A_795_423#_c_651_n 0.0215259f $X=3.51 $Y=2.635
+ $X2=0 $Y2=0
cc_310 N_A_200_481#_c_262_n N_A_795_423#_c_651_n 6.19391e-19 $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_311 N_A_200_481#_c_274_n N_A_795_423#_c_651_n 0.00589862f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_312 N_A_200_481#_c_274_n N_A_795_423#_c_653_n 0.00618103f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_313 N_A_200_481#_c_271_n N_A_609_485#_M1020_d 0.00311887f $X=3.435 $Y=2.485
+ $X2=0 $Y2=0
cc_314 N_A_200_481#_M1005_g N_A_609_485#_c_799_n 0.0146531f $X=3.51 $Y=2.635
+ $X2=0 $Y2=0
cc_315 N_A_200_481#_c_271_n N_A_609_485#_c_799_n 0.0374641f $X=3.435 $Y=2.485
+ $X2=0 $Y2=0
cc_316 N_A_200_481#_c_274_n N_A_609_485#_c_799_n 0.00222307f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_317 N_A_200_481#_M1005_g N_A_609_485#_c_792_n 0.00417693f $X=3.51 $Y=2.635
+ $X2=0 $Y2=0
cc_318 N_A_200_481#_c_271_n N_A_609_485#_c_792_n 0.013908f $X=3.435 $Y=2.485
+ $X2=0 $Y2=0
cc_319 N_A_200_481#_c_261_n N_A_609_485#_c_792_n 0.00622081f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_320 N_A_200_481#_c_262_n N_A_609_485#_c_792_n 0.0684716f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_321 N_A_200_481#_c_274_n N_A_609_485#_c_792_n 0.00254738f $X=3.6 $Y=2.045
+ $X2=0 $Y2=0
cc_322 N_A_200_481#_c_260_n N_A_609_485#_c_794_n 0.00315408f $X=3.245 $Y=1.325
+ $X2=0 $Y2=0
cc_323 N_A_200_481#_c_261_n N_A_609_485#_c_794_n 0.0076837f $X=3.565 $Y=1.495
+ $X2=0 $Y2=0
cc_324 N_A_200_481#_c_269_n N_VPWR_M1014_d 0.00152634f $X=1.96 $Y=2.99 $X2=0
+ $Y2=0
cc_325 N_A_200_481#_c_297_p N_VPWR_M1014_d 0.00389344f $X=2.045 $Y=2.905 $X2=0
+ $Y2=0
cc_326 N_A_200_481#_c_271_n N_VPWR_M1014_d 0.00670698f $X=3.435 $Y=2.485 $X2=0
+ $Y2=0
cc_327 N_A_200_481#_c_268_n N_VPWR_c_891_n 7.29177e-19 $X=1.14 $Y=2.56 $X2=0
+ $Y2=0
cc_328 N_A_200_481#_c_270_n N_VPWR_c_891_n 0.00251712f $X=1.305 $Y=2.99 $X2=0
+ $Y2=0
cc_329 N_A_200_481#_M1014_g N_VPWR_c_892_n 0.0027647f $X=1.91 $Y=2.745 $X2=0
+ $Y2=0
cc_330 N_A_200_481#_c_269_n N_VPWR_c_892_n 0.0142704f $X=1.96 $Y=2.99 $X2=0
+ $Y2=0
cc_331 N_A_200_481#_c_297_p N_VPWR_c_892_n 0.0123418f $X=2.045 $Y=2.905 $X2=0
+ $Y2=0
cc_332 N_A_200_481#_c_271_n N_VPWR_c_892_n 0.0156969f $X=3.435 $Y=2.485 $X2=0
+ $Y2=0
cc_333 N_A_200_481#_M1014_g N_VPWR_c_899_n 0.0033828f $X=1.91 $Y=2.745 $X2=0
+ $Y2=0
cc_334 N_A_200_481#_c_269_n N_VPWR_c_899_n 0.0538669f $X=1.96 $Y=2.99 $X2=0
+ $Y2=0
cc_335 N_A_200_481#_c_270_n N_VPWR_c_899_n 0.021506f $X=1.305 $Y=2.99 $X2=0
+ $Y2=0
cc_336 N_A_200_481#_c_271_n N_VPWR_c_899_n 0.00227783f $X=3.435 $Y=2.485 $X2=0
+ $Y2=0
cc_337 N_A_200_481#_M1005_g N_VPWR_c_904_n 7.94025e-19 $X=3.51 $Y=2.635 $X2=0
+ $Y2=0
cc_338 N_A_200_481#_c_271_n N_VPWR_c_904_n 0.00519804f $X=3.435 $Y=2.485 $X2=0
+ $Y2=0
cc_339 N_A_200_481#_M1014_g N_VPWR_c_890_n 0.00665088f $X=1.91 $Y=2.745 $X2=0
+ $Y2=0
cc_340 N_A_200_481#_c_269_n N_VPWR_c_890_n 0.0305438f $X=1.96 $Y=2.99 $X2=0
+ $Y2=0
cc_341 N_A_200_481#_c_270_n N_VPWR_c_890_n 0.0116633f $X=1.305 $Y=2.99 $X2=0
+ $Y2=0
cc_342 N_A_200_481#_c_271_n N_VPWR_c_890_n 0.0167342f $X=3.435 $Y=2.485 $X2=0
+ $Y2=0
cc_343 N_A_200_481#_c_271_n A_537_485# 0.00190305f $X=3.435 $Y=2.485 $X2=-0.19
+ $Y2=-0.245
cc_344 N_A_200_481#_c_271_n A_717_485# 0.00189254f $X=3.435 $Y=2.485 $X2=-0.19
+ $Y2=-0.245
cc_345 N_A_200_481#_c_253_n N_VGND_c_1057_n 0.00764533f $X=2.365 $Y=0.77 $X2=0
+ $Y2=0
cc_346 N_A_200_481#_M1012_g N_VGND_c_1057_n 0.00179412f $X=3.155 $Y=0.445 $X2=0
+ $Y2=0
cc_347 N_A_200_481#_c_253_n N_VGND_c_1065_n 0.0035231f $X=2.365 $Y=0.77 $X2=0
+ $Y2=0
cc_348 N_A_200_481#_c_255_n N_VGND_c_1065_n 0.00438783f $X=2.365 $Y=0.845 $X2=0
+ $Y2=0
cc_349 N_A_200_481#_M1012_g N_VGND_c_1066_n 0.0042361f $X=3.155 $Y=0.445 $X2=0
+ $Y2=0
cc_350 N_A_200_481#_c_253_n N_VGND_c_1073_n 0.00524031f $X=2.365 $Y=0.77 $X2=0
+ $Y2=0
cc_351 N_A_200_481#_M1012_g N_VGND_c_1073_n 0.00602557f $X=3.155 $Y=0.445 $X2=0
+ $Y2=0
cc_352 N_A_200_481#_c_255_n N_VGND_c_1073_n 0.00509645f $X=2.365 $Y=0.845 $X2=0
+ $Y2=0
cc_353 N_A_200_481#_c_263_n N_VGND_c_1073_n 0.00100231f $X=1.917 $Y=1.055 $X2=0
+ $Y2=0
cc_354 N_A_27_481#_c_421_n N_A_310_485#_c_503_n 0.0379344f $X=2.52 $Y=1.785
+ $X2=0 $Y2=0
cc_355 N_A_27_481#_c_460_n N_A_310_485#_c_503_n 0.00140925f $X=2.52 $Y=1.445
+ $X2=0 $Y2=0
cc_356 N_A_27_481#_M1004_g N_A_310_485#_c_514_n 0.0340287f $X=2.61 $Y=2.745
+ $X2=0 $Y2=0
cc_357 N_A_27_481#_M1004_g N_A_310_485#_c_516_n 0.0111473f $X=2.61 $Y=2.745
+ $X2=0 $Y2=0
cc_358 N_A_27_481#_c_427_n N_A_310_485#_c_516_n 0.0050701f $X=2.52 $Y=1.95 $X2=0
+ $Y2=0
cc_359 N_A_27_481#_c_430_n N_A_310_485#_c_516_n 0.0677047f $X=2.355 $Y=1.79
+ $X2=0 $Y2=0
cc_360 N_A_27_481#_c_430_n N_A_310_485#_c_517_n 0.0212104f $X=2.355 $Y=1.79
+ $X2=0 $Y2=0
cc_361 N_A_27_481#_M1009_g N_A_310_485#_c_508_n 0.0110349f $X=2.795 $Y=0.445
+ $X2=0 $Y2=0
cc_362 N_A_27_481#_c_423_n N_A_310_485#_c_508_n 8.81106e-19 $X=2.52 $Y=1.445
+ $X2=0 $Y2=0
cc_363 N_A_27_481#_c_421_n N_A_310_485#_c_564_n 3.13799e-19 $X=2.52 $Y=1.785
+ $X2=0 $Y2=0
cc_364 N_A_27_481#_c_427_n N_A_310_485#_c_564_n 0.0011595f $X=2.52 $Y=1.95 $X2=0
+ $Y2=0
cc_365 N_A_27_481#_c_430_n N_A_310_485#_c_564_n 0.012087f $X=2.355 $Y=1.79 $X2=0
+ $Y2=0
cc_366 N_A_27_481#_c_460_n N_A_310_485#_c_564_n 0.00155265f $X=2.52 $Y=1.445
+ $X2=0 $Y2=0
cc_367 N_A_27_481#_c_427_n N_A_310_485#_c_510_n 0.0340287f $X=2.52 $Y=1.95 $X2=0
+ $Y2=0
cc_368 N_A_27_481#_c_430_n N_A_310_485#_c_510_n 6.25005e-19 $X=2.355 $Y=1.79
+ $X2=0 $Y2=0
cc_369 N_A_27_481#_M1004_g N_A_609_485#_c_799_n 7.53302e-19 $X=2.61 $Y=2.745
+ $X2=0 $Y2=0
cc_370 N_A_27_481#_c_429_n N_VPWR_c_891_n 0.0014656f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_371 N_A_27_481#_c_430_n N_VPWR_c_891_n 0.00993218f $X=2.355 $Y=1.79 $X2=0
+ $Y2=0
cc_372 N_A_27_481#_M1004_g N_VPWR_c_892_n 0.0105067f $X=2.61 $Y=2.745 $X2=0
+ $Y2=0
cc_373 N_A_27_481#_c_429_n N_VPWR_c_903_n 0.0202345f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_374 N_A_27_481#_M1004_g N_VPWR_c_904_n 0.00346665f $X=2.61 $Y=2.745 $X2=0
+ $Y2=0
cc_375 N_A_27_481#_M1004_g N_VPWR_c_890_n 0.00416619f $X=2.61 $Y=2.745 $X2=0
+ $Y2=0
cc_376 N_A_27_481#_c_429_n N_VPWR_c_890_n 0.0122439f $X=0.26 $Y=2.55 $X2=0 $Y2=0
cc_377 N_A_27_481#_M1009_g N_VGND_c_1057_n 0.00877879f $X=2.795 $Y=0.445 $X2=0
+ $Y2=0
cc_378 N_A_27_481#_M1009_g N_VGND_c_1066_n 0.0035231f $X=2.795 $Y=0.445 $X2=0
+ $Y2=0
cc_379 N_A_27_481#_c_424_n N_VGND_c_1069_n 0.00604219f $X=0.34 $Y=0.845 $X2=0
+ $Y2=0
cc_380 N_A_27_481#_M1009_g N_VGND_c_1073_n 0.00400373f $X=2.795 $Y=0.445 $X2=0
+ $Y2=0
cc_381 N_A_27_481#_c_424_n N_VGND_c_1073_n 0.0107791f $X=0.34 $Y=0.845 $X2=0
+ $Y2=0
cc_382 N_A_310_485#_M1015_g N_A_795_423#_M1022_g 0.020968f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_383 N_A_310_485#_c_511_n N_A_795_423#_M1022_g 9.83513e-19 $X=3.785 $Y=0.71
+ $X2=0 $Y2=0
cc_384 N_A_310_485#_c_512_n N_A_795_423#_M1022_g 0.0328615f $X=3.785 $Y=0.98
+ $X2=0 $Y2=0
cc_385 N_A_310_485#_c_505_n N_A_795_423#_c_627_n 0.00304959f $X=3.695 $Y=1.49
+ $X2=0 $Y2=0
cc_386 N_A_310_485#_c_502_n N_A_795_423#_c_636_n 0.00304959f $X=3.62 $Y=1.565
+ $X2=0 $Y2=0
cc_387 N_A_310_485#_c_502_n N_A_795_423#_c_641_n 0.0012857f $X=3.62 $Y=1.565
+ $X2=0 $Y2=0
cc_388 N_A_310_485#_c_508_n N_A_609_485#_M1012_d 0.00287031f $X=3.62 $Y=0.71
+ $X2=-0.19 $Y2=-0.245
cc_389 N_A_310_485#_M1020_g N_A_609_485#_c_799_n 0.00502594f $X=2.97 $Y=2.745
+ $X2=0 $Y2=0
cc_390 N_A_310_485#_M1015_g N_A_609_485#_c_815_n 0.0118335f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_391 N_A_310_485#_c_508_n N_A_609_485#_c_815_n 0.0192199f $X=3.62 $Y=0.71
+ $X2=0 $Y2=0
cc_392 N_A_310_485#_c_511_n N_A_609_485#_c_815_n 0.0196013f $X=3.785 $Y=0.71
+ $X2=0 $Y2=0
cc_393 N_A_310_485#_c_512_n N_A_609_485#_c_815_n 7.18523e-19 $X=3.785 $Y=0.98
+ $X2=0 $Y2=0
cc_394 N_A_310_485#_c_505_n N_A_609_485#_c_792_n 0.00205618f $X=3.695 $Y=1.49
+ $X2=0 $Y2=0
cc_395 N_A_310_485#_c_507_n N_A_609_485#_c_792_n 6.31904e-19 $X=3.785 $Y=1.34
+ $X2=0 $Y2=0
cc_396 N_A_310_485#_M1015_g N_A_609_485#_c_793_n 3.86856e-19 $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_397 N_A_310_485#_c_511_n N_A_609_485#_c_793_n 0.0312599f $X=3.785 $Y=0.71
+ $X2=0 $Y2=0
cc_398 N_A_310_485#_c_512_n N_A_609_485#_c_793_n 0.00494658f $X=3.785 $Y=0.98
+ $X2=0 $Y2=0
cc_399 N_A_310_485#_c_505_n N_A_609_485#_c_794_n 6.3907e-19 $X=3.695 $Y=1.49
+ $X2=0 $Y2=0
cc_400 N_A_310_485#_c_507_n N_A_609_485#_c_794_n 0.00573551f $X=3.785 $Y=1.34
+ $X2=0 $Y2=0
cc_401 N_A_310_485#_c_511_n N_A_609_485#_c_794_n 0.00589379f $X=3.785 $Y=0.71
+ $X2=0 $Y2=0
cc_402 N_A_310_485#_M1020_g N_VPWR_c_892_n 0.00200675f $X=2.97 $Y=2.745 $X2=0
+ $Y2=0
cc_403 N_A_310_485#_M1020_g N_VPWR_c_904_n 0.00405543f $X=2.97 $Y=2.745 $X2=0
+ $Y2=0
cc_404 N_A_310_485#_M1020_g N_VPWR_c_890_n 0.00682237f $X=2.97 $Y=2.745 $X2=0
+ $Y2=0
cc_405 N_A_310_485#_c_508_n N_VGND_M1023_d 0.00169275f $X=3.62 $Y=0.71 $X2=0
+ $Y2=0
cc_406 N_A_310_485#_c_508_n N_VGND_c_1057_n 0.0159471f $X=3.62 $Y=0.71 $X2=0
+ $Y2=0
cc_407 N_A_310_485#_c_521_n N_VGND_c_1065_n 0.0136564f $X=2.15 $Y=0.435 $X2=0
+ $Y2=0
cc_408 N_A_310_485#_c_508_n N_VGND_c_1065_n 0.00262544f $X=3.62 $Y=0.71 $X2=0
+ $Y2=0
cc_409 N_A_310_485#_M1015_g N_VGND_c_1066_n 0.00357877f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_410 N_A_310_485#_c_508_n N_VGND_c_1066_n 0.00764761f $X=3.62 $Y=0.71 $X2=0
+ $Y2=0
cc_411 N_A_310_485#_M1023_s N_VGND_c_1073_n 0.00245903f $X=2.025 $Y=0.235 $X2=0
+ $Y2=0
cc_412 N_A_310_485#_M1015_g N_VGND_c_1073_n 0.005989f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_413 N_A_310_485#_c_521_n N_VGND_c_1073_n 0.00764688f $X=2.15 $Y=0.435 $X2=0
+ $Y2=0
cc_414 N_A_310_485#_c_508_n N_VGND_c_1073_n 0.0199092f $X=3.62 $Y=0.71 $X2=0
+ $Y2=0
cc_415 N_A_310_485#_c_508_n A_574_47# 0.00165214f $X=3.62 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_416 N_A_310_485#_c_511_n A_754_47# 0.00154654f $X=3.785 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_417 N_A_795_423#_M1022_g N_A_609_485#_c_790_n 0.0238741f $X=4.235 $Y=0.445
+ $X2=0 $Y2=0
cc_418 N_A_795_423#_c_639_n N_A_609_485#_c_790_n 0.0031023f $X=5.295 $Y=1.345
+ $X2=0 $Y2=0
cc_419 N_A_795_423#_c_636_n N_A_609_485#_M1002_g 0.00219399f $X=4.3 $Y=1.595
+ $X2=0 $Y2=0
cc_420 N_A_795_423#_c_637_n N_A_609_485#_M1002_g 3.95987e-19 $X=4.31 $Y=1.845
+ $X2=0 $Y2=0
cc_421 N_A_795_423#_c_652_n N_A_609_485#_M1002_g 3.03243e-19 $X=4.3 $Y=2.1 $X2=0
+ $Y2=0
cc_422 N_A_795_423#_c_654_n N_A_609_485#_M1002_g 0.0146001f $X=5.085 $Y=1.76
+ $X2=0 $Y2=0
cc_423 N_A_795_423#_c_655_n N_A_609_485#_M1002_g 0.00412809f $X=5.18 $Y=1.9
+ $X2=0 $Y2=0
cc_424 N_A_795_423#_c_640_n N_A_609_485#_M1002_g 0.00440107f $X=5.29 $Y=1.675
+ $X2=0 $Y2=0
cc_425 N_A_795_423#_c_641_n N_A_609_485#_M1002_g 0.0127733f $X=4.3 $Y=1.76 $X2=0
+ $Y2=0
cc_426 N_A_795_423#_M1013_g N_A_609_485#_c_799_n 0.00751866f $X=4.05 $Y=2.635
+ $X2=0 $Y2=0
cc_427 N_A_795_423#_M1022_g N_A_609_485#_c_815_n 0.00778803f $X=4.235 $Y=0.445
+ $X2=0 $Y2=0
cc_428 N_A_795_423#_M1013_g N_A_609_485#_c_792_n 0.0118674f $X=4.05 $Y=2.635
+ $X2=0 $Y2=0
cc_429 N_A_795_423#_c_627_n N_A_609_485#_c_792_n 0.00324778f $X=4.25 $Y=1.43
+ $X2=0 $Y2=0
cc_430 N_A_795_423#_c_651_n N_A_609_485#_c_792_n 0.00520299f $X=4.22 $Y=2.265
+ $X2=0 $Y2=0
cc_431 N_A_795_423#_c_637_n N_A_609_485#_c_792_n 0.0193181f $X=4.31 $Y=1.845
+ $X2=0 $Y2=0
cc_432 N_A_795_423#_c_652_n N_A_609_485#_c_792_n 0.029877f $X=4.3 $Y=2.1 $X2=0
+ $Y2=0
cc_433 N_A_795_423#_c_641_n N_A_609_485#_c_792_n 0.00815846f $X=4.3 $Y=1.76
+ $X2=0 $Y2=0
cc_434 N_A_795_423#_M1022_g N_A_609_485#_c_793_n 0.0209233f $X=4.235 $Y=0.445
+ $X2=0 $Y2=0
cc_435 N_A_795_423#_M1022_g N_A_609_485#_c_794_n 0.00249727f $X=4.235 $Y=0.445
+ $X2=0 $Y2=0
cc_436 N_A_795_423#_c_627_n N_A_609_485#_c_794_n 0.00523633f $X=4.25 $Y=1.43
+ $X2=0 $Y2=0
cc_437 N_A_795_423#_c_637_n N_A_609_485#_c_794_n 0.0132147f $X=4.31 $Y=1.845
+ $X2=0 $Y2=0
cc_438 N_A_795_423#_c_641_n N_A_609_485#_c_794_n 0.00101678f $X=4.3 $Y=1.76
+ $X2=0 $Y2=0
cc_439 N_A_795_423#_c_627_n N_A_609_485#_c_795_n 3.64484e-19 $X=4.25 $Y=1.43
+ $X2=0 $Y2=0
cc_440 N_A_795_423#_c_654_n N_A_609_485#_c_795_n 0.0238144f $X=5.085 $Y=1.76
+ $X2=0 $Y2=0
cc_441 N_A_795_423#_c_639_n N_A_609_485#_c_795_n 0.00790617f $X=5.295 $Y=1.345
+ $X2=0 $Y2=0
cc_442 N_A_795_423#_c_642_n N_A_609_485#_c_795_n 0.0107543f $X=5.137 $Y=1.075
+ $X2=0 $Y2=0
cc_443 N_A_795_423#_c_643_n N_A_609_485#_c_795_n 0.013783f $X=5.295 $Y=1.43
+ $X2=0 $Y2=0
cc_444 N_A_795_423#_c_644_n N_A_609_485#_c_795_n 2.38919e-19 $X=5.81 $Y=1.43
+ $X2=0 $Y2=0
cc_445 N_A_795_423#_M1022_g N_A_609_485#_c_796_n 0.00188779f $X=4.235 $Y=0.445
+ $X2=0 $Y2=0
cc_446 N_A_795_423#_c_627_n N_A_609_485#_c_796_n 0.00236845f $X=4.25 $Y=1.43
+ $X2=0 $Y2=0
cc_447 N_A_795_423#_c_637_n N_A_609_485#_c_796_n 0.00172158f $X=4.31 $Y=1.845
+ $X2=0 $Y2=0
cc_448 N_A_795_423#_c_654_n N_A_609_485#_c_796_n 0.0160003f $X=5.085 $Y=1.76
+ $X2=0 $Y2=0
cc_449 N_A_795_423#_c_641_n N_A_609_485#_c_796_n 0.00244398f $X=4.3 $Y=1.76
+ $X2=0 $Y2=0
cc_450 N_A_795_423#_c_627_n N_A_609_485#_c_797_n 0.00547562f $X=4.25 $Y=1.43
+ $X2=0 $Y2=0
cc_451 N_A_795_423#_c_654_n N_A_609_485#_c_797_n 0.00479409f $X=5.085 $Y=1.76
+ $X2=0 $Y2=0
cc_452 N_A_795_423#_c_639_n N_A_609_485#_c_797_n 0.00327859f $X=5.295 $Y=1.345
+ $X2=0 $Y2=0
cc_453 N_A_795_423#_c_642_n N_A_609_485#_c_797_n 0.00432167f $X=5.137 $Y=1.075
+ $X2=0 $Y2=0
cc_454 N_A_795_423#_c_643_n N_A_609_485#_c_797_n 0.00149876f $X=5.295 $Y=1.43
+ $X2=0 $Y2=0
cc_455 N_A_795_423#_c_644_n N_A_609_485#_c_797_n 0.0125427f $X=5.81 $Y=1.43
+ $X2=0 $Y2=0
cc_456 N_A_795_423#_c_654_n N_VPWR_M1013_d 0.00253128f $X=5.085 $Y=1.76 $X2=0
+ $Y2=0
cc_457 N_A_795_423#_M1013_g N_VPWR_c_894_n 0.00282633f $X=4.05 $Y=2.635 $X2=0
+ $Y2=0
cc_458 N_A_795_423#_c_652_n N_VPWR_c_894_n 0.0191203f $X=4.3 $Y=2.1 $X2=0 $Y2=0
cc_459 N_A_795_423#_c_653_n N_VPWR_c_894_n 0.00237191f $X=4.3 $Y=2.1 $X2=0 $Y2=0
cc_460 N_A_795_423#_c_654_n N_VPWR_c_894_n 0.0220026f $X=5.085 $Y=1.76 $X2=0
+ $Y2=0
cc_461 N_A_795_423#_c_655_n N_VPWR_c_894_n 0.0417649f $X=5.18 $Y=1.9 $X2=0 $Y2=0
cc_462 N_A_795_423#_M1001_g N_VPWR_c_895_n 0.00767654f $X=5.915 $Y=2.465 $X2=0
+ $Y2=0
cc_463 N_A_795_423#_c_655_n N_VPWR_c_895_n 0.0970019f $X=5.18 $Y=1.9 $X2=0 $Y2=0
cc_464 N_A_795_423#_c_718_p N_VPWR_c_895_n 0.0149606f $X=6.53 $Y=1.43 $X2=0
+ $Y2=0
cc_465 N_A_795_423#_c_658_n N_VPWR_c_895_n 0.00262627f $X=5.23 $Y=1.76 $X2=0
+ $Y2=0
cc_466 N_A_795_423#_c_644_n N_VPWR_c_895_n 0.00679391f $X=5.81 $Y=1.43 $X2=0
+ $Y2=0
cc_467 N_A_795_423#_M1001_g N_VPWR_c_896_n 7.59349e-19 $X=5.915 $Y=2.465 $X2=0
+ $Y2=0
cc_468 N_A_795_423#_M1006_g N_VPWR_c_896_n 0.0147414f $X=6.345 $Y=2.465 $X2=0
+ $Y2=0
cc_469 N_A_795_423#_M1011_g N_VPWR_c_896_n 0.00161651f $X=6.775 $Y=2.465 $X2=0
+ $Y2=0
cc_470 N_A_795_423#_M1011_g N_VPWR_c_898_n 8.12047e-19 $X=6.775 $Y=2.465 $X2=0
+ $Y2=0
cc_471 N_A_795_423#_M1019_g N_VPWR_c_898_n 0.0216233f $X=7.205 $Y=2.465 $X2=0
+ $Y2=0
cc_472 N_A_795_423#_M1013_g N_VPWR_c_962_n 0.00476356f $X=4.05 $Y=2.635 $X2=0
+ $Y2=0
cc_473 N_A_795_423#_c_651_n N_VPWR_c_962_n 0.0033152f $X=4.22 $Y=2.265 $X2=0
+ $Y2=0
cc_474 N_A_795_423#_c_652_n N_VPWR_c_962_n 0.0181368f $X=4.3 $Y=2.1 $X2=0 $Y2=0
cc_475 N_A_795_423#_c_654_n N_VPWR_c_962_n 0.00549911f $X=5.085 $Y=1.76 $X2=0
+ $Y2=0
cc_476 N_A_795_423#_c_655_n N_VPWR_c_901_n 0.0164655f $X=5.18 $Y=1.9 $X2=0 $Y2=0
cc_477 N_A_795_423#_M1013_g N_VPWR_c_904_n 0.00330087f $X=4.05 $Y=2.635 $X2=0
+ $Y2=0
cc_478 N_A_795_423#_M1001_g N_VPWR_c_905_n 0.00585385f $X=5.915 $Y=2.465 $X2=0
+ $Y2=0
cc_479 N_A_795_423#_M1006_g N_VPWR_c_905_n 0.00486043f $X=6.345 $Y=2.465 $X2=0
+ $Y2=0
cc_480 N_A_795_423#_M1011_g N_VPWR_c_906_n 0.00585385f $X=6.775 $Y=2.465 $X2=0
+ $Y2=0
cc_481 N_A_795_423#_M1019_g N_VPWR_c_906_n 0.00525069f $X=7.205 $Y=2.465 $X2=0
+ $Y2=0
cc_482 N_A_795_423#_M1013_g N_VPWR_c_890_n 0.00305932f $X=4.05 $Y=2.635 $X2=0
+ $Y2=0
cc_483 N_A_795_423#_M1001_g N_VPWR_c_890_n 0.0118221f $X=5.915 $Y=2.465 $X2=0
+ $Y2=0
cc_484 N_A_795_423#_M1006_g N_VPWR_c_890_n 0.00824727f $X=6.345 $Y=2.465 $X2=0
+ $Y2=0
cc_485 N_A_795_423#_M1011_g N_VPWR_c_890_n 0.0105224f $X=6.775 $Y=2.465 $X2=0
+ $Y2=0
cc_486 N_A_795_423#_M1019_g N_VPWR_c_890_n 0.00886509f $X=7.205 $Y=2.465 $X2=0
+ $Y2=0
cc_487 N_A_795_423#_c_655_n N_VPWR_c_890_n 0.0109746f $X=5.18 $Y=1.9 $X2=0 $Y2=0
cc_488 N_A_795_423#_M1010_g N_Q_c_1004_n 0.0132064f $X=6.315 $Y=0.655 $X2=0
+ $Y2=0
cc_489 N_A_795_423#_M1016_g N_Q_c_1004_n 0.0145206f $X=6.745 $Y=0.655 $X2=0
+ $Y2=0
cc_490 N_A_795_423#_c_718_p N_Q_c_1004_n 0.0350722f $X=6.53 $Y=1.43 $X2=0 $Y2=0
cc_491 N_A_795_423#_c_645_n N_Q_c_1004_n 0.00259366f $X=7.175 $Y=1.43 $X2=0
+ $Y2=0
cc_492 N_A_795_423#_M1000_g N_Q_c_1005_n 0.00151567f $X=5.885 $Y=0.655 $X2=0
+ $Y2=0
cc_493 N_A_795_423#_c_639_n N_Q_c_1005_n 0.00283779f $X=5.295 $Y=1.345 $X2=0
+ $Y2=0
cc_494 N_A_795_423#_c_718_p N_Q_c_1005_n 0.0181554f $X=6.53 $Y=1.43 $X2=0 $Y2=0
cc_495 N_A_795_423#_c_645_n N_Q_c_1005_n 0.00269667f $X=7.175 $Y=1.43 $X2=0
+ $Y2=0
cc_496 N_A_795_423#_M1006_g N_Q_c_1008_n 0.0137063f $X=6.345 $Y=2.465 $X2=0
+ $Y2=0
cc_497 N_A_795_423#_M1011_g N_Q_c_1008_n 0.0159576f $X=6.775 $Y=2.465 $X2=0
+ $Y2=0
cc_498 N_A_795_423#_c_718_p N_Q_c_1008_n 0.03302f $X=6.53 $Y=1.43 $X2=0 $Y2=0
cc_499 N_A_795_423#_c_645_n N_Q_c_1008_n 0.00259366f $X=7.175 $Y=1.43 $X2=0
+ $Y2=0
cc_500 N_A_795_423#_M1001_g N_Q_c_1009_n 0.00243205f $X=5.915 $Y=2.465 $X2=0
+ $Y2=0
cc_501 N_A_795_423#_c_718_p N_Q_c_1009_n 0.0181554f $X=6.53 $Y=1.43 $X2=0 $Y2=0
cc_502 N_A_795_423#_c_658_n N_Q_c_1009_n 0.00483787f $X=5.23 $Y=1.76 $X2=0 $Y2=0
cc_503 N_A_795_423#_c_645_n N_Q_c_1009_n 0.00269667f $X=7.175 $Y=1.43 $X2=0
+ $Y2=0
cc_504 N_A_795_423#_M1018_g Q 0.00286881f $X=7.175 $Y=0.655 $X2=0 $Y2=0
cc_505 N_A_795_423#_M1016_g Q 0.00227886f $X=6.745 $Y=0.655 $X2=0 $Y2=0
cc_506 N_A_795_423#_M1011_g Q 0.00236762f $X=6.775 $Y=2.465 $X2=0 $Y2=0
cc_507 N_A_795_423#_M1018_g Q 0.00239819f $X=7.175 $Y=0.655 $X2=0 $Y2=0
cc_508 N_A_795_423#_M1019_g Q 0.00230796f $X=7.205 $Y=2.465 $X2=0 $Y2=0
cc_509 N_A_795_423#_c_718_p Q 0.0130696f $X=6.53 $Y=1.43 $X2=0 $Y2=0
cc_510 N_A_795_423#_c_645_n Q 0.034985f $X=7.175 $Y=1.43 $X2=0 $Y2=0
cc_511 N_A_795_423#_M1019_g Q 0.00438093f $X=7.205 $Y=2.465 $X2=0 $Y2=0
cc_512 N_A_795_423#_M1022_g N_VGND_c_1058_n 0.00722947f $X=4.235 $Y=0.445 $X2=0
+ $Y2=0
cc_513 N_A_795_423#_M1000_g N_VGND_c_1059_n 0.00705062f $X=5.885 $Y=0.655 $X2=0
+ $Y2=0
cc_514 N_A_795_423#_c_638_n N_VGND_c_1059_n 0.069225f $X=4.995 $Y=0.42 $X2=0
+ $Y2=0
cc_515 N_A_795_423#_c_718_p N_VGND_c_1059_n 0.0147147f $X=6.53 $Y=1.43 $X2=0
+ $Y2=0
cc_516 N_A_795_423#_c_644_n N_VGND_c_1059_n 0.00597448f $X=5.81 $Y=1.43 $X2=0
+ $Y2=0
cc_517 N_A_795_423#_M1000_g N_VGND_c_1060_n 6.28227e-19 $X=5.885 $Y=0.655 $X2=0
+ $Y2=0
cc_518 N_A_795_423#_M1010_g N_VGND_c_1060_n 0.0102576f $X=6.315 $Y=0.655 $X2=0
+ $Y2=0
cc_519 N_A_795_423#_M1016_g N_VGND_c_1060_n 0.0104021f $X=6.745 $Y=0.655 $X2=0
+ $Y2=0
cc_520 N_A_795_423#_M1018_g N_VGND_c_1060_n 6.39229e-19 $X=7.175 $Y=0.655 $X2=0
+ $Y2=0
cc_521 N_A_795_423#_M1018_g N_VGND_c_1062_n 0.00699379f $X=7.175 $Y=0.655 $X2=0
+ $Y2=0
cc_522 N_A_795_423#_c_645_n N_VGND_c_1062_n 5.59349e-19 $X=7.175 $Y=1.43 $X2=0
+ $Y2=0
cc_523 N_A_795_423#_c_638_n N_VGND_c_1063_n 0.0342954f $X=4.995 $Y=0.42 $X2=0
+ $Y2=0
cc_524 N_A_795_423#_M1022_g N_VGND_c_1066_n 0.00372849f $X=4.235 $Y=0.445 $X2=0
+ $Y2=0
cc_525 N_A_795_423#_M1000_g N_VGND_c_1067_n 0.00585385f $X=5.885 $Y=0.655 $X2=0
+ $Y2=0
cc_526 N_A_795_423#_M1010_g N_VGND_c_1067_n 0.00486043f $X=6.315 $Y=0.655 $X2=0
+ $Y2=0
cc_527 N_A_795_423#_M1016_g N_VGND_c_1068_n 0.00486043f $X=6.745 $Y=0.655 $X2=0
+ $Y2=0
cc_528 N_A_795_423#_M1018_g N_VGND_c_1068_n 0.00585385f $X=7.175 $Y=0.655 $X2=0
+ $Y2=0
cc_529 N_A_795_423#_M1021_d N_VGND_c_1073_n 0.00336915f $X=4.855 $Y=0.235 $X2=0
+ $Y2=0
cc_530 N_A_795_423#_M1022_g N_VGND_c_1073_n 0.00637924f $X=4.235 $Y=0.445 $X2=0
+ $Y2=0
cc_531 N_A_795_423#_M1000_g N_VGND_c_1073_n 0.0118221f $X=5.885 $Y=0.655 $X2=0
+ $Y2=0
cc_532 N_A_795_423#_M1010_g N_VGND_c_1073_n 0.00824727f $X=6.315 $Y=0.655 $X2=0
+ $Y2=0
cc_533 N_A_795_423#_M1016_g N_VGND_c_1073_n 0.00824727f $X=6.745 $Y=0.655 $X2=0
+ $Y2=0
cc_534 N_A_795_423#_M1018_g N_VGND_c_1073_n 0.0114959f $X=7.175 $Y=0.655 $X2=0
+ $Y2=0
cc_535 N_A_795_423#_c_638_n N_VGND_c_1073_n 0.0191667f $X=4.995 $Y=0.42 $X2=0
+ $Y2=0
cc_536 N_A_609_485#_c_799_n N_VPWR_c_892_n 0.00969809f $X=3.865 $Y=2.88 $X2=0
+ $Y2=0
cc_537 N_A_609_485#_M1002_g N_VPWR_c_893_n 0.00808958f $X=4.965 $Y=2.385 $X2=0
+ $Y2=0
cc_538 N_A_609_485#_M1002_g N_VPWR_c_894_n 0.00479687f $X=4.965 $Y=2.385 $X2=0
+ $Y2=0
cc_539 N_A_609_485#_c_792_n N_VPWR_c_894_n 0.00528102f $X=3.95 $Y=2.74 $X2=0
+ $Y2=0
cc_540 N_A_609_485#_M1002_g N_VPWR_c_895_n 0.00299433f $X=4.965 $Y=2.385 $X2=0
+ $Y2=0
cc_541 N_A_609_485#_M1002_g N_VPWR_c_962_n 0.00378169f $X=4.965 $Y=2.385 $X2=0
+ $Y2=0
cc_542 N_A_609_485#_c_799_n N_VPWR_c_962_n 0.0249039f $X=3.865 $Y=2.88 $X2=0
+ $Y2=0
cc_543 N_A_609_485#_c_792_n N_VPWR_c_962_n 0.0240124f $X=3.95 $Y=2.74 $X2=0
+ $Y2=0
cc_544 N_A_609_485#_M1002_g N_VPWR_c_901_n 0.00422142f $X=4.965 $Y=2.385 $X2=0
+ $Y2=0
cc_545 N_A_609_485#_c_799_n N_VPWR_c_904_n 0.0492374f $X=3.865 $Y=2.88 $X2=0
+ $Y2=0
cc_546 N_A_609_485#_M1002_g N_VPWR_c_890_n 0.00853956f $X=4.965 $Y=2.385 $X2=0
+ $Y2=0
cc_547 N_A_609_485#_c_799_n N_VPWR_c_890_n 0.0373799f $X=3.865 $Y=2.88 $X2=0
+ $Y2=0
cc_548 N_A_609_485#_c_799_n A_717_485# 0.00586413f $X=3.865 $Y=2.88 $X2=-0.19
+ $Y2=-0.245
cc_549 N_A_609_485#_c_792_n A_717_485# 0.00339801f $X=3.95 $Y=2.74 $X2=-0.19
+ $Y2=-0.245
cc_550 N_A_609_485#_c_790_n N_VGND_c_1058_n 0.0116376f $X=4.78 $Y=1.185 $X2=0
+ $Y2=0
cc_551 N_A_609_485#_c_815_n N_VGND_c_1058_n 0.0161536f $X=4.13 $Y=0.355 $X2=0
+ $Y2=0
cc_552 N_A_609_485#_c_793_n N_VGND_c_1058_n 0.0310829f $X=4.215 $Y=1.245 $X2=0
+ $Y2=0
cc_553 N_A_609_485#_c_796_n N_VGND_c_1058_n 0.010375f $X=4.705 $Y=1.375 $X2=0
+ $Y2=0
cc_554 N_A_609_485#_c_790_n N_VGND_c_1063_n 0.00525069f $X=4.78 $Y=1.185 $X2=0
+ $Y2=0
cc_555 N_A_609_485#_c_815_n N_VGND_c_1066_n 0.0615844f $X=4.13 $Y=0.355 $X2=0
+ $Y2=0
cc_556 N_A_609_485#_M1012_d N_VGND_c_1073_n 0.00320398f $X=3.23 $Y=0.235 $X2=0
+ $Y2=0
cc_557 N_A_609_485#_c_790_n N_VGND_c_1073_n 0.0101648f $X=4.78 $Y=1.185 $X2=0
+ $Y2=0
cc_558 N_A_609_485#_c_815_n N_VGND_c_1073_n 0.0384826f $X=4.13 $Y=0.355 $X2=0
+ $Y2=0
cc_559 N_A_609_485#_c_815_n A_754_47# 0.0100285f $X=4.13 $Y=0.355 $X2=-0.19
+ $Y2=-0.245
cc_560 N_VPWR_c_890_n N_Q_M1001_s 0.0041489f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_561 N_VPWR_c_890_n N_Q_M1011_s 0.00380103f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_562 N_VPWR_c_905_n N_Q_c_1038_n 0.0136943f $X=6.395 $Y=3.33 $X2=0 $Y2=0
cc_563 N_VPWR_c_890_n N_Q_c_1038_n 0.00866972f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_564 N_VPWR_M1006_d N_Q_c_1008_n 0.00176461f $X=6.42 $Y=1.835 $X2=0 $Y2=0
cc_565 N_VPWR_c_896_n N_Q_c_1008_n 0.0152916f $X=6.56 $Y=2.19 $X2=0 $Y2=0
cc_566 N_VPWR_c_895_n N_Q_c_1009_n 0.00166212f $X=5.7 $Y=1.98 $X2=0 $Y2=0
cc_567 N_VPWR_c_898_n Q 0.0023867f $X=7.42 $Y=1.98 $X2=0 $Y2=0
cc_568 N_VPWR_c_906_n Q 0.0140491f $X=7.265 $Y=3.33 $X2=0 $Y2=0
cc_569 N_VPWR_c_890_n Q 0.0090585f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_570 N_Q_c_1004_n N_VGND_M1010_d 0.00176461f $X=6.865 $Y=1.09 $X2=0 $Y2=0
cc_571 N_Q_c_1005_n N_VGND_c_1059_n 0.00164453f $X=6.195 $Y=1.09 $X2=0 $Y2=0
cc_572 N_Q_c_1004_n N_VGND_c_1060_n 0.0170777f $X=6.865 $Y=1.09 $X2=0 $Y2=0
cc_573 Q N_VGND_c_1062_n 0.0016373f $X=6.875 $Y=0.84 $X2=0 $Y2=0
cc_574 N_Q_c_1050_p N_VGND_c_1067_n 0.0136943f $X=6.1 $Y=0.42 $X2=0 $Y2=0
cc_575 N_Q_c_1051_p N_VGND_c_1068_n 0.0135169f $X=6.96 $Y=0.42 $X2=0 $Y2=0
cc_576 N_Q_M1000_s N_VGND_c_1073_n 0.0041489f $X=5.96 $Y=0.235 $X2=0 $Y2=0
cc_577 N_Q_M1016_s N_VGND_c_1073_n 0.00432284f $X=6.82 $Y=0.235 $X2=0 $Y2=0
cc_578 N_Q_c_1050_p N_VGND_c_1073_n 0.00866972f $X=6.1 $Y=0.42 $X2=0 $Y2=0
cc_579 N_Q_c_1051_p N_VGND_c_1073_n 0.00847005f $X=6.96 $Y=0.42 $X2=0 $Y2=0
cc_580 N_VGND_c_1073_n A_574_47# 0.00241193f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
cc_581 N_VGND_c_1073_n A_754_47# 0.00313854f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
