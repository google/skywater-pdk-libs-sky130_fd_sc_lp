* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4_0 A B C D VGND VNB VPB VPWR X
X0 VPWR A a_84_58# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_84_58# A a_167_58# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_84_58# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_84_58# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR a_84_58# X VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VPWR C a_84_58# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_311_58# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_84_58# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_239_58# C a_311_58# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_167_58# B a_239_58# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
