* NGSPICE file created from sky130_fd_sc_lp__and3b_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and3b_m A_N B C VGND VNB VPB VPWR X
M1000 a_220_53# B VPWR VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=4.116e+11p ps=4.48e+06u
M1001 X a_220_53# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1002 a_304_53# a_110_53# a_220_53# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.134e+11p ps=1.38e+06u
M1003 a_376_53# B a_304_53# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1004 VPWR a_110_53# a_220_53# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND C a_376_53# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1006 a_110_53# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 VPWR C a_220_53# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_110_53# A_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1009 X a_220_53# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

