# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o22a_0
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.990000 1.170000 1.295000 1.215000 ;
        RECT 0.990000 1.215000 1.685000 1.395000 ;
        RECT 0.995000 0.265000 1.325000 0.435000 ;
        RECT 0.995000 0.435000 1.295000 0.500000 ;
        RECT 1.115000 0.500000 1.295000 1.170000 ;
        RECT 1.515000 1.395000 1.685000 2.095000 ;
        RECT 1.515000 2.095000 3.370000 2.265000 ;
        RECT 3.060000 1.935000 3.370000 2.095000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.245000 1.115000 3.755000 1.415000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 1.565000 1.345000 2.235000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 1.385000 2.735000 1.925000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.280900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.605000 0.465000 0.935000 ;
        RECT 0.085000 0.935000 0.325000 2.425000 ;
        RECT 0.085000 2.425000 0.425000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.495000  1.565000 0.665000 2.065000 ;
      RECT 0.495000  2.065000 0.765000 2.235000 ;
      RECT 0.595000  2.235000 0.765000 2.435000 ;
      RECT 0.595000  2.435000 3.745000 2.605000 ;
      RECT 0.595000  2.775000 1.735000 3.245000 ;
      RECT 0.645000  0.085000 0.825000 0.670000 ;
      RECT 0.645000  0.670000 0.945000 1.000000 ;
      RECT 1.465000  0.615000 1.685000 1.000000 ;
      RECT 1.495000  0.445000 2.695000 0.615000 ;
      RECT 1.855000  0.785000 2.185000 1.035000 ;
      RECT 1.855000  1.035000 3.075000 1.205000 ;
      RECT 2.225000  2.605000 2.555000 3.075000 ;
      RECT 2.365000  0.615000 2.695000 0.865000 ;
      RECT 2.875000  0.085000 3.205000 0.865000 ;
      RECT 2.905000  1.205000 3.075000 1.585000 ;
      RECT 2.905000  1.585000 3.745000 1.755000 ;
      RECT 3.185000  2.775000 3.515000 3.245000 ;
      RECT 3.540000  1.755000 3.745000 2.435000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__o22a_0
END LIBRARY
