* File: sky130_fd_sc_lp__nor4b_4.pxi.spice
* Created: Wed Sep  2 10:11:09 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4B_4%D_N N_D_N_M1033_g N_D_N_M1027_g D_N N_D_N_c_146_n
+ N_D_N_c_147_n PM_SKY130_FD_SC_LP__NOR4B_4%D_N
x_PM_SKY130_FD_SC_LP__NOR4B_4%A_27_367# N_A_27_367#_M1027_s N_A_27_367#_M1033_s
+ N_A_27_367#_M1004_g N_A_27_367#_M1009_g N_A_27_367#_M1005_g
+ N_A_27_367#_M1006_g N_A_27_367#_M1024_g N_A_27_367#_M1018_g
+ N_A_27_367#_M1029_g N_A_27_367#_M1031_g N_A_27_367#_c_195_n
+ N_A_27_367#_c_196_n N_A_27_367#_c_183_n N_A_27_367#_c_197_n
+ N_A_27_367#_c_184_n N_A_27_367#_c_185_n N_A_27_367#_c_186_n
+ N_A_27_367#_c_187_n N_A_27_367#_c_188_n N_A_27_367#_c_189_n
+ N_A_27_367#_c_190_n PM_SKY130_FD_SC_LP__NOR4B_4%A_27_367#
x_PM_SKY130_FD_SC_LP__NOR4B_4%C N_C_M1001_g N_C_M1008_g N_C_M1016_g N_C_M1012_g
+ N_C_M1025_g N_C_M1021_g N_C_M1030_g N_C_M1023_g C C N_C_c_311_n N_C_c_361_p C
+ N_C_c_312_n PM_SKY130_FD_SC_LP__NOR4B_4%C
x_PM_SKY130_FD_SC_LP__NOR4B_4%B N_B_M1000_g N_B_M1007_g N_B_M1003_g N_B_M1014_g
+ N_B_M1015_g N_B_M1019_g N_B_M1017_g N_B_M1026_g B B B N_B_c_394_n
+ PM_SKY130_FD_SC_LP__NOR4B_4%B
x_PM_SKY130_FD_SC_LP__NOR4B_4%A N_A_M1011_g N_A_M1002_g N_A_M1013_g N_A_M1010_g
+ N_A_M1022_g N_A_M1020_g N_A_M1028_g N_A_M1032_g A A A N_A_c_486_n N_A_c_487_n
+ N_A_c_488_n A N_A_c_489_n PM_SKY130_FD_SC_LP__NOR4B_4%A
x_PM_SKY130_FD_SC_LP__NOR4B_4%VPWR N_VPWR_M1033_d N_VPWR_M1002_d N_VPWR_M1020_d
+ N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_565_n
+ N_VPWR_c_566_n N_VPWR_c_567_n VPWR N_VPWR_c_568_n N_VPWR_c_569_n
+ N_VPWR_c_560_n N_VPWR_c_571_n PM_SKY130_FD_SC_LP__NOR4B_4%VPWR
x_PM_SKY130_FD_SC_LP__NOR4B_4%A_217_367# N_A_217_367#_M1005_s
+ N_A_217_367#_M1006_s N_A_217_367#_M1031_s N_A_217_367#_M1012_d
+ N_A_217_367#_M1023_d N_A_217_367#_c_698_n N_A_217_367#_c_673_n
+ N_A_217_367#_c_682_n N_A_217_367#_c_719_p N_A_217_367#_c_684_n
+ N_A_217_367#_c_722_p N_A_217_367#_c_686_n N_A_217_367#_c_726_p
+ N_A_217_367#_c_674_n N_A_217_367#_c_675_n N_A_217_367#_c_710_n
+ N_A_217_367#_c_712_n N_A_217_367#_c_714_n
+ PM_SKY130_FD_SC_LP__NOR4B_4%A_217_367#
x_PM_SKY130_FD_SC_LP__NOR4B_4%Y N_Y_M1004_s N_Y_M1024_s N_Y_M1001_s N_Y_M1025_s
+ N_Y_M1000_d N_Y_M1015_d N_Y_M1011_s N_Y_M1022_s N_Y_M1005_d N_Y_M1018_d
+ N_Y_c_877_p N_Y_c_733_n N_Y_c_734_n N_Y_c_759_n N_Y_c_746_n N_Y_c_747_n
+ N_Y_c_878_p N_Y_c_735_n N_Y_c_774_n N_Y_c_748_n N_Y_c_869_p N_Y_c_736_n
+ N_Y_c_737_n N_Y_c_874_p N_Y_c_738_n N_Y_c_875_p N_Y_c_833_n N_Y_c_876_p
+ N_Y_c_739_n N_Y_c_750_n N_Y_c_740_n N_Y_c_741_n N_Y_c_742_n Y Y Y Y
+ N_Y_c_805_n N_Y_c_810_n N_Y_c_745_n N_Y_c_899_p N_Y_c_879_p
+ PM_SKY130_FD_SC_LP__NOR4B_4%Y
x_PM_SKY130_FD_SC_LP__NOR4B_4%A_644_367# N_A_644_367#_M1008_s
+ N_A_644_367#_M1021_s N_A_644_367#_M1007_s N_A_644_367#_M1019_s
+ N_A_644_367#_c_906_n N_A_644_367#_c_934_n N_A_644_367#_c_905_n
+ N_A_644_367#_c_946_p N_A_644_367#_c_915_n N_A_644_367#_c_909_n
+ N_A_644_367#_c_941_n N_A_644_367#_c_919_n N_A_644_367#_c_921_n
+ PM_SKY130_FD_SC_LP__NOR4B_4%A_644_367#
x_PM_SKY130_FD_SC_LP__NOR4B_4%A_1009_367# N_A_1009_367#_M1007_d
+ N_A_1009_367#_M1014_d N_A_1009_367#_M1026_d N_A_1009_367#_M1010_s
+ N_A_1009_367#_M1032_s N_A_1009_367#_c_950_n N_A_1009_367#_c_960_n
+ N_A_1009_367#_c_951_n N_A_1009_367#_c_1012_n N_A_1009_367#_c_963_n
+ N_A_1009_367#_c_992_n N_A_1009_367#_c_952_n N_A_1009_367#_c_953_n
+ N_A_1009_367#_c_996_n N_A_1009_367#_c_954_n N_A_1009_367#_c_955_n
+ N_A_1009_367#_c_1002_n N_A_1009_367#_c_956_n
+ PM_SKY130_FD_SC_LP__NOR4B_4%A_1009_367#
x_PM_SKY130_FD_SC_LP__NOR4B_4%VGND N_VGND_M1027_d N_VGND_M1009_d N_VGND_M1029_d
+ N_VGND_M1016_d N_VGND_M1030_d N_VGND_M1003_s N_VGND_M1017_s N_VGND_M1013_d
+ N_VGND_M1028_d N_VGND_c_1015_n N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n
+ N_VGND_c_1019_n N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n
+ N_VGND_c_1023_n N_VGND_c_1024_n N_VGND_c_1025_n N_VGND_c_1026_n
+ N_VGND_c_1027_n N_VGND_c_1028_n N_VGND_c_1029_n VGND N_VGND_c_1030_n
+ N_VGND_c_1031_n N_VGND_c_1032_n N_VGND_c_1033_n N_VGND_c_1034_n
+ N_VGND_c_1035_n N_VGND_c_1036_n N_VGND_c_1037_n N_VGND_c_1038_n
+ N_VGND_c_1039_n N_VGND_c_1040_n N_VGND_c_1041_n N_VGND_c_1042_n
+ PM_SKY130_FD_SC_LP__NOR4B_4%VGND
cc_1 VNB N_D_N_M1033_g 0.00193879f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB N_D_N_M1027_g 0.0294645f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.655
cc_3 VNB N_D_N_c_146_n 0.0379134f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.46
cc_4 VNB N_D_N_c_147_n 0.0146281f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.46
cc_5 VNB N_A_27_367#_M1004_g 0.018645f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_27_367#_M1009_g 0.0184866f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.46
cc_7 VNB N_A_27_367#_M1005_g 0.00535162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_367#_M1006_g 0.00452622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_367#_M1024_g 0.0186996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_367#_M1018_g 0.00452622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_367#_M1029_g 0.0209152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_367#_M1031_g 0.00467754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_367#_c_183_n 0.0277218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_367#_c_184_n 0.00572279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_367#_c_185_n 0.00933582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_367#_c_186_n 0.00154157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_367#_c_187_n 0.00211781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_367#_c_188_n 0.00112218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_367#_c_189_n 0.00109104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_367#_c_190_n 0.130245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C_M1001_g 0.0209152f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_22 VNB N_C_M1008_g 0.00467754f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.655
cc_23 VNB N_C_M1016_g 0.0185234f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.46
cc_24 VNB N_C_M1012_g 0.00452622f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.625
cc_25 VNB N_C_M1025_g 0.0184495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C_M1021_g 0.00452622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C_M1030_g 0.0219645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C_M1023_g 0.00572192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB C 0.00690638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_c_311_n 0.0994231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C_c_312_n 0.00112218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_M1000_g 0.0280445f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_33 VNB N_B_M1003_g 0.023169f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.46
cc_34 VNB N_B_M1015_g 0.0231894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_M1017_g 0.0236356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB B 0.0023978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_394_n 0.0720172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_M1011_g 0.0203821f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_39 VNB N_A_M1002_g 0.00257131f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.655
cc_40 VNB N_A_M1013_g 0.0204771f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.46
cc_41 VNB N_A_M1010_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.625
cc_42 VNB N_A_M1022_g 0.0200495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_M1020_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_M1028_g 0.0270322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_M1032_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB A 0.0318619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_c_486_n 0.0764182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_c_487_n 0.0626476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_c_488_n 0.00179308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_c_489_n 0.00132888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VPWR_c_560_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_Y_c_733_n 0.00288059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_Y_c_734_n 0.00201249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_Y_c_735_n 0.00658468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_Y_c_736_n 0.0101794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Y_c_737_n 0.00306317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Y_c_738_n 0.00568741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Y_c_739_n 0.00172316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_Y_c_740_n 0.00227375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_Y_c_741_n 0.00145644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_Y_c_742_n 0.00232334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB Y 0.00224459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB Y 0.00145644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_Y_c_745_n 0.00674194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1015_n 0.00222256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1016_n 0.00220289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1017_n 0.00180234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1018_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1019_n 3.08929e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1020_n 3.08929e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1021_n 3.16049e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1022_n 3.16049e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1023_n 0.0339216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1024_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1025_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1026_n 0.0138364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1027_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1028_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1029_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1030_n 0.0156941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1031_n 0.01612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1032_n 0.0146078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1033_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1034_n 0.0143948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1035_n 0.439958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1036_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1037_n 0.00525267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1038_n 0.0106533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1039_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1040_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1041_n 0.016163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1042_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VPB N_D_N_M1033_g 0.0285084f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_94 VPB N_D_N_c_147_n 0.00726557f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.46
cc_95 VPB N_A_27_367#_M1005_g 0.0232962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_27_367#_M1006_g 0.0183695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_27_367#_M1018_g 0.0183695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_27_367#_M1031_g 0.0184535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_27_367#_c_195_n 0.00755006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_27_367#_c_196_n 0.0369431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_27_367#_c_197_n 0.00510572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_27_367#_c_187_n 0.00491198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_C_M1008_g 0.0184604f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.655
cc_104 VPB N_C_M1012_g 0.0183765f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.625
cc_105 VPB N_C_M1021_g 0.0183765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_C_M1023_g 0.0236789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_B_M1007_g 0.0224653f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.655
cc_108 VPB N_B_M1014_g 0.0173921f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.625
cc_109 VPB N_B_M1019_g 0.0173921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_B_M1026_g 0.0183445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB B 0.0102727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_B_c_394_n 0.0149551f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_M1002_g 0.0185418f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.655
cc_114 VPB N_A_M1010_g 0.0184123f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.625
cc_115 VPB N_A_M1020_g 0.0184123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_M1032_g 0.0243928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_561_n 0.0111769f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.46
cc_118 VPB N_VPWR_c_562_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.46
cc_119 VPB N_VPWR_c_563_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_564_n 0.144214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_565_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_566_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_567_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_568_n 0.0153759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_569_n 0.0233314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_560_n 0.0743348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_571_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_217_367#_c_673_n 0.00207782f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.665
cc_129 VPB N_A_217_367#_c_674_n 0.00181979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_217_367#_c_675_n 0.00526929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_Y_c_746_n 0.00716512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_Y_c_747_n 0.00233203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_Y_c_748_n 0.0344056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_Y_c_736_n 2.13491e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_Y_c_750_n 0.00233203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_644_367#_c_905_n 0.0116064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_1009_367#_c_950_n 0.00526929f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.665
cc_138 VPB N_A_1009_367#_c_951_n 0.00181979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_1009_367#_c_952_n 0.00290381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_1009_367#_c_953_n 0.00367337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_1009_367#_c_954_n 0.0145696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_1009_367#_c_955_n 0.0435297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_1009_367#_c_956_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 N_D_N_M1027_g N_A_27_367#_M1004_g 0.0159185f $X=0.485 $Y=0.655 $X2=0
+ $Y2=0
cc_145 N_D_N_c_146_n N_A_27_367#_c_195_n 7.41055e-19 $X=0.385 $Y=1.46 $X2=0
+ $Y2=0
cc_146 N_D_N_c_147_n N_A_27_367#_c_195_n 0.0226401f $X=0.385 $Y=1.46 $X2=0 $Y2=0
cc_147 N_D_N_M1033_g N_A_27_367#_c_197_n 0.0137783f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_D_N_c_147_n N_A_27_367#_c_197_n 0.0128665f $X=0.385 $Y=1.46 $X2=0 $Y2=0
cc_149 N_D_N_M1027_g N_A_27_367#_c_184_n 0.0143468f $X=0.485 $Y=0.655 $X2=0
+ $Y2=0
cc_150 N_D_N_c_146_n N_A_27_367#_c_184_n 0.00108293f $X=0.385 $Y=1.46 $X2=0
+ $Y2=0
cc_151 N_D_N_c_147_n N_A_27_367#_c_184_n 0.0136372f $X=0.385 $Y=1.46 $X2=0 $Y2=0
cc_152 N_D_N_c_146_n N_A_27_367#_c_185_n 0.00349977f $X=0.385 $Y=1.46 $X2=0
+ $Y2=0
cc_153 N_D_N_c_147_n N_A_27_367#_c_185_n 0.0229487f $X=0.385 $Y=1.46 $X2=0 $Y2=0
cc_154 N_D_N_M1027_g N_A_27_367#_c_186_n 0.00342474f $X=0.485 $Y=0.655 $X2=0
+ $Y2=0
cc_155 N_D_N_M1033_g N_A_27_367#_c_187_n 0.00850562f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_D_N_c_146_n N_A_27_367#_c_187_n 0.00181301f $X=0.385 $Y=1.46 $X2=0
+ $Y2=0
cc_157 N_D_N_c_147_n N_A_27_367#_c_187_n 0.0214441f $X=0.385 $Y=1.46 $X2=0 $Y2=0
cc_158 N_D_N_c_146_n N_A_27_367#_c_189_n 0.00128064f $X=0.385 $Y=1.46 $X2=0
+ $Y2=0
cc_159 N_D_N_c_147_n N_A_27_367#_c_189_n 0.013818f $X=0.385 $Y=1.46 $X2=0 $Y2=0
cc_160 N_D_N_M1027_g N_A_27_367#_c_190_n 0.0205025f $X=0.485 $Y=0.655 $X2=0
+ $Y2=0
cc_161 N_D_N_c_147_n N_A_27_367#_c_190_n 2.65069e-19 $X=0.385 $Y=1.46 $X2=0
+ $Y2=0
cc_162 N_D_N_M1033_g N_VPWR_c_561_n 0.0186436f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_163 N_D_N_M1033_g N_VPWR_c_568_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_164 N_D_N_M1033_g N_VPWR_c_560_n 0.00917987f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_165 N_D_N_M1033_g N_A_217_367#_c_673_n 0.0053647f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_D_N_M1027_g N_VGND_c_1015_n 0.0116791f $X=0.485 $Y=0.655 $X2=0 $Y2=0
cc_167 N_D_N_M1027_g N_VGND_c_1030_n 0.00486043f $X=0.485 $Y=0.655 $X2=0 $Y2=0
cc_168 N_D_N_M1027_g N_VGND_c_1035_n 0.00918921f $X=0.485 $Y=0.655 $X2=0 $Y2=0
cc_169 N_A_27_367#_M1029_g N_C_M1001_g 0.00763827f $X=2.305 $Y=0.655 $X2=0 $Y2=0
cc_170 N_A_27_367#_M1031_g N_C_M1008_g 0.0256219f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A_27_367#_c_188_n N_C_c_311_n 2.08417e-19 $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_172 N_A_27_367#_c_190_n N_C_c_311_n 0.0245335f $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_173 N_A_27_367#_c_188_n N_C_c_312_n 0.0119872f $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_174 N_A_27_367#_c_190_n N_C_c_312_n 2.08417e-19 $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_175 N_A_27_367#_c_197_n N_VPWR_M1033_d 0.00730404f $X=0.72 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A_27_367#_c_187_n N_VPWR_M1033_d 0.00155748f $X=0.822 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_177 N_A_27_367#_M1005_g N_VPWR_c_561_n 0.002302f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_27_367#_c_197_n N_VPWR_c_561_n 0.0230836f $X=0.72 $Y=2.015 $X2=0
+ $Y2=0
cc_179 N_A_27_367#_M1005_g N_VPWR_c_564_n 0.00357877f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_27_367#_M1006_g N_VPWR_c_564_n 0.00357877f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_27_367#_M1018_g N_VPWR_c_564_n 0.00357877f $X=2.285 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_27_367#_M1031_g N_VPWR_c_564_n 0.00357877f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_27_367#_c_196_n N_VPWR_c_568_n 0.0178111f $X=0.26 $Y=2.91 $X2=0 $Y2=0
cc_184 N_A_27_367#_M1033_s N_VPWR_c_560_n 0.00371702f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_185 N_A_27_367#_M1005_g N_VPWR_c_560_n 0.00665089f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A_27_367#_M1006_g N_VPWR_c_560_n 0.0053512f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_27_367#_M1018_g N_VPWR_c_560_n 0.0053512f $X=2.285 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_27_367#_M1031_g N_VPWR_c_560_n 0.00537654f $X=2.715 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_A_27_367#_c_196_n N_VPWR_c_560_n 0.0100304f $X=0.26 $Y=2.91 $X2=0 $Y2=0
cc_190 N_A_27_367#_M1005_g N_A_217_367#_c_673_n 0.00334874f $X=1.425 $Y=2.465
+ $X2=0 $Y2=0
cc_191 N_A_27_367#_c_197_n N_A_217_367#_c_673_n 0.0143312f $X=0.72 $Y=2.015
+ $X2=0 $Y2=0
cc_192 N_A_27_367#_c_187_n N_A_217_367#_c_673_n 0.00875455f $X=0.822 $Y=1.93
+ $X2=0 $Y2=0
cc_193 N_A_27_367#_c_188_n N_A_217_367#_c_673_n 0.0102637f $X=2.635 $Y=1.4 $X2=0
+ $Y2=0
cc_194 N_A_27_367#_c_190_n N_A_217_367#_c_673_n 0.00524748f $X=2.715 $Y=1.4
+ $X2=0 $Y2=0
cc_195 N_A_27_367#_M1005_g N_A_217_367#_c_682_n 0.0115031f $X=1.425 $Y=2.465
+ $X2=0 $Y2=0
cc_196 N_A_27_367#_M1006_g N_A_217_367#_c_682_n 0.0114565f $X=1.855 $Y=2.465
+ $X2=0 $Y2=0
cc_197 N_A_27_367#_M1018_g N_A_217_367#_c_684_n 0.0115031f $X=2.285 $Y=2.465
+ $X2=0 $Y2=0
cc_198 N_A_27_367#_M1031_g N_A_217_367#_c_684_n 0.0115031f $X=2.715 $Y=2.465
+ $X2=0 $Y2=0
cc_199 N_A_27_367#_M1009_g N_Y_c_733_n 0.0140118f $X=1.395 $Y=0.655 $X2=0 $Y2=0
cc_200 N_A_27_367#_M1024_g N_Y_c_733_n 0.0143795f $X=1.875 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A_27_367#_c_188_n N_Y_c_733_n 0.0469361f $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_202 N_A_27_367#_c_190_n N_Y_c_733_n 0.00391713f $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_203 N_A_27_367#_M1004_g N_Y_c_734_n 5.60107e-19 $X=0.965 $Y=0.655 $X2=0 $Y2=0
cc_204 N_A_27_367#_c_184_n N_Y_c_734_n 0.0100024f $X=0.72 $Y=1.07 $X2=0 $Y2=0
cc_205 N_A_27_367#_c_188_n N_Y_c_734_n 0.0161378f $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_206 N_A_27_367#_c_190_n N_Y_c_734_n 0.00256759f $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_207 N_A_27_367#_M1005_g N_Y_c_759_n 0.00990505f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A_27_367#_M1006_g N_Y_c_759_n 0.0106535f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A_27_367#_M1018_g N_Y_c_759_n 6.41373e-19 $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A_27_367#_M1006_g N_Y_c_746_n 0.0112007f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A_27_367#_M1018_g N_Y_c_746_n 0.0112007f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A_27_367#_c_188_n N_Y_c_746_n 0.0353087f $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_213 N_A_27_367#_c_190_n N_Y_c_746_n 0.00253405f $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_214 N_A_27_367#_M1005_g N_Y_c_747_n 0.00561586f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A_27_367#_M1006_g N_Y_c_747_n 0.00279204f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A_27_367#_c_187_n N_Y_c_747_n 0.00497405f $X=0.822 $Y=1.93 $X2=0 $Y2=0
cc_217 N_A_27_367#_c_188_n N_Y_c_747_n 0.0252825f $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_218 N_A_27_367#_c_190_n N_Y_c_747_n 0.00255521f $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_219 N_A_27_367#_M1029_g N_Y_c_735_n 0.0147947f $X=2.305 $Y=0.655 $X2=0 $Y2=0
cc_220 N_A_27_367#_c_188_n N_Y_c_735_n 0.0435831f $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_221 N_A_27_367#_c_190_n N_Y_c_735_n 0.0116986f $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_222 N_A_27_367#_M1006_g N_Y_c_774_n 6.41373e-19 $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A_27_367#_M1018_g N_Y_c_774_n 0.0106535f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_27_367#_M1031_g N_Y_c_774_n 0.0107923f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A_27_367#_M1031_g N_Y_c_748_n 0.0111542f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A_27_367#_c_188_n N_Y_c_748_n 0.0087457f $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_227 N_A_27_367#_c_190_n N_Y_c_748_n 2.44902e-19 $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_228 N_A_27_367#_c_188_n N_Y_c_739_n 0.0177519f $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_229 N_A_27_367#_c_190_n N_Y_c_739_n 0.00265365f $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_230 N_A_27_367#_M1018_g N_Y_c_750_n 0.00279204f $X=2.285 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_27_367#_M1031_g N_Y_c_750_n 0.00279204f $X=2.715 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A_27_367#_c_188_n N_Y_c_750_n 0.0252825f $X=2.635 $Y=1.4 $X2=0 $Y2=0
cc_233 N_A_27_367#_c_190_n N_Y_c_750_n 0.00255521f $X=2.715 $Y=1.4 $X2=0 $Y2=0
cc_234 N_A_27_367#_c_184_n N_VGND_M1027_d 0.00233477f $X=0.72 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_235 N_A_27_367#_M1004_g N_VGND_c_1015_n 0.00168004f $X=0.965 $Y=0.655 $X2=0
+ $Y2=0
cc_236 N_A_27_367#_c_184_n N_VGND_c_1015_n 0.0203178f $X=0.72 $Y=1.07 $X2=0
+ $Y2=0
cc_237 N_A_27_367#_c_190_n N_VGND_c_1015_n 3.67726e-19 $X=2.715 $Y=1.4 $X2=0
+ $Y2=0
cc_238 N_A_27_367#_M1004_g N_VGND_c_1016_n 5.99888e-19 $X=0.965 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_A_27_367#_M1009_g N_VGND_c_1016_n 0.00819291f $X=1.395 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_27_367#_M1024_g N_VGND_c_1016_n 0.00171412f $X=1.875 $Y=0.655 $X2=0
+ $Y2=0
cc_241 N_A_27_367#_M1024_g N_VGND_c_1017_n 6.27507e-19 $X=1.875 $Y=0.655 $X2=0
+ $Y2=0
cc_242 N_A_27_367#_M1029_g N_VGND_c_1017_n 0.0107588f $X=2.305 $Y=0.655 $X2=0
+ $Y2=0
cc_243 N_A_27_367#_c_183_n N_VGND_c_1030_n 0.0178111f $X=0.27 $Y=0.42 $X2=0
+ $Y2=0
cc_244 N_A_27_367#_M1004_g N_VGND_c_1031_n 0.00585385f $X=0.965 $Y=0.655 $X2=0
+ $Y2=0
cc_245 N_A_27_367#_M1009_g N_VGND_c_1031_n 0.00564095f $X=1.395 $Y=0.655 $X2=0
+ $Y2=0
cc_246 N_A_27_367#_M1024_g N_VGND_c_1032_n 0.00585385f $X=1.875 $Y=0.655 $X2=0
+ $Y2=0
cc_247 N_A_27_367#_M1029_g N_VGND_c_1032_n 0.00486043f $X=2.305 $Y=0.655 $X2=0
+ $Y2=0
cc_248 N_A_27_367#_M1027_s N_VGND_c_1035_n 0.00371702f $X=0.145 $Y=0.235 $X2=0
+ $Y2=0
cc_249 N_A_27_367#_M1004_g N_VGND_c_1035_n 0.0107048f $X=0.965 $Y=0.655 $X2=0
+ $Y2=0
cc_250 N_A_27_367#_M1009_g N_VGND_c_1035_n 0.00948291f $X=1.395 $Y=0.655 $X2=0
+ $Y2=0
cc_251 N_A_27_367#_M1024_g N_VGND_c_1035_n 0.0106333f $X=1.875 $Y=0.655 $X2=0
+ $Y2=0
cc_252 N_A_27_367#_M1029_g N_VGND_c_1035_n 0.00824727f $X=2.305 $Y=0.655 $X2=0
+ $Y2=0
cc_253 N_A_27_367#_c_183_n N_VGND_c_1035_n 0.0100304f $X=0.27 $Y=0.42 $X2=0
+ $Y2=0
cc_254 N_C_c_311_n N_B_M1000_g 0.00556344f $X=4.535 $Y=1.4 $X2=0 $Y2=0
cc_255 N_C_M1023_g N_B_c_394_n 0.00101774f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_256 N_C_M1008_g N_VPWR_c_564_n 0.00357877f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_257 N_C_M1012_g N_VPWR_c_564_n 0.00357877f $X=3.575 $Y=2.465 $X2=0 $Y2=0
cc_258 N_C_M1021_g N_VPWR_c_564_n 0.00357877f $X=4.005 $Y=2.465 $X2=0 $Y2=0
cc_259 N_C_M1023_g N_VPWR_c_564_n 0.00357842f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_260 N_C_M1008_g N_VPWR_c_560_n 0.00537654f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_261 N_C_M1012_g N_VPWR_c_560_n 0.0053512f $X=3.575 $Y=2.465 $X2=0 $Y2=0
cc_262 N_C_M1021_g N_VPWR_c_560_n 0.0053512f $X=4.005 $Y=2.465 $X2=0 $Y2=0
cc_263 N_C_M1023_g N_VPWR_c_560_n 0.00665087f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_264 N_C_M1008_g N_A_217_367#_c_686_n 0.0115031f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_265 N_C_M1012_g N_A_217_367#_c_686_n 0.0115031f $X=3.575 $Y=2.465 $X2=0 $Y2=0
cc_266 N_C_M1021_g N_A_217_367#_c_674_n 0.012237f $X=4.005 $Y=2.465 $X2=0 $Y2=0
cc_267 N_C_M1023_g N_A_217_367#_c_674_n 0.0111017f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_268 N_C_M1021_g N_A_217_367#_c_675_n 5.5465e-19 $X=4.005 $Y=2.465 $X2=0 $Y2=0
cc_269 N_C_M1023_g N_A_217_367#_c_675_n 0.00850024f $X=4.435 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_C_M1001_g N_Y_c_735_n 0.0146256f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_271 N_C_c_312_n N_Y_c_735_n 0.0134081f $X=3.885 $Y=1.347 $X2=0 $Y2=0
cc_272 N_C_M1008_g N_Y_c_774_n 9.67954e-19 $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_273 N_C_M1008_g N_Y_c_748_n 0.014324f $X=3.145 $Y=2.465 $X2=0 $Y2=0
cc_274 N_C_M1012_g N_Y_c_748_n 0.0105529f $X=3.575 $Y=2.465 $X2=0 $Y2=0
cc_275 N_C_M1021_g N_Y_c_748_n 0.0105539f $X=4.005 $Y=2.465 $X2=0 $Y2=0
cc_276 N_C_M1023_g N_Y_c_748_n 0.0123714f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_277 N_C_c_311_n N_Y_c_748_n 0.01449f $X=4.535 $Y=1.4 $X2=0 $Y2=0
cc_278 N_C_c_312_n N_Y_c_748_n 0.115492f $X=3.885 $Y=1.347 $X2=0 $Y2=0
cc_279 N_C_M1030_g N_Y_c_736_n 7.74296e-19 $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_280 N_C_M1023_g N_Y_c_736_n 0.00195832f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_281 C N_Y_c_736_n 0.022102f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_282 N_C_c_311_n N_Y_c_736_n 0.00307083f $X=4.535 $Y=1.4 $X2=0 $Y2=0
cc_283 N_C_M1016_g N_Y_c_740_n 0.00224236f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_284 N_C_c_311_n N_Y_c_740_n 0.00282576f $X=4.535 $Y=1.4 $X2=0 $Y2=0
cc_285 N_C_c_312_n N_Y_c_740_n 0.0160848f $X=3.885 $Y=1.347 $X2=0 $Y2=0
cc_286 C Y 0.0151777f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_287 N_C_c_311_n Y 7.34815e-19 $X=4.535 $Y=1.4 $X2=0 $Y2=0
cc_288 N_C_M1030_g Y 0.00457663f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_289 N_C_M1016_g N_Y_c_805_n 0.0111976f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_290 N_C_M1025_g N_Y_c_805_n 0.0106173f $X=3.945 $Y=0.655 $X2=0 $Y2=0
cc_291 N_C_c_311_n N_Y_c_805_n 0.00253467f $X=4.535 $Y=1.4 $X2=0 $Y2=0
cc_292 N_C_c_361_p N_Y_c_805_n 0.0112833f $X=4.022 $Y=1.347 $X2=0 $Y2=0
cc_293 N_C_c_312_n N_Y_c_805_n 0.019269f $X=3.885 $Y=1.347 $X2=0 $Y2=0
cc_294 N_C_M1030_g N_Y_c_810_n 0.0129857f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_295 C N_Y_c_810_n 0.0297806f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_296 N_C_c_311_n N_Y_c_810_n 0.0015348f $X=4.535 $Y=1.4 $X2=0 $Y2=0
cc_297 N_C_M1012_g N_A_644_367#_c_906_n 0.0114269f $X=3.575 $Y=2.465 $X2=0 $Y2=0
cc_298 N_C_M1021_g N_A_644_367#_c_906_n 0.0133021f $X=4.005 $Y=2.465 $X2=0 $Y2=0
cc_299 N_C_M1023_g N_A_644_367#_c_905_n 0.0147239f $X=4.435 $Y=2.465 $X2=0 $Y2=0
cc_300 N_C_M1008_g N_A_644_367#_c_909_n 0.00961578f $X=3.145 $Y=2.465 $X2=0
+ $Y2=0
cc_301 N_C_M1012_g N_A_644_367#_c_909_n 0.00959704f $X=3.575 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_C_M1021_g N_A_644_367#_c_909_n 5.5465e-19 $X=4.005 $Y=2.465 $X2=0 $Y2=0
cc_303 N_C_M1023_g N_A_1009_367#_c_950_n 9.94534e-19 $X=4.435 $Y=2.465 $X2=0
+ $Y2=0
cc_304 N_C_M1001_g N_VGND_c_1017_n 0.0106896f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_305 N_C_M1016_g N_VGND_c_1017_n 6.14488e-19 $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_306 N_C_M1001_g N_VGND_c_1018_n 0.00486043f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_307 N_C_M1016_g N_VGND_c_1018_n 0.00486043f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_308 N_C_M1001_g N_VGND_c_1019_n 5.67328e-19 $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_309 N_C_M1016_g N_VGND_c_1019_n 0.00996624f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_310 N_C_M1025_g N_VGND_c_1019_n 0.00995595f $X=3.945 $Y=0.655 $X2=0 $Y2=0
cc_311 N_C_M1030_g N_VGND_c_1019_n 5.66918e-19 $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_312 N_C_M1001_g N_VGND_c_1035_n 0.00824727f $X=3.085 $Y=0.655 $X2=0 $Y2=0
cc_313 N_C_M1016_g N_VGND_c_1035_n 0.00454119f $X=3.515 $Y=0.655 $X2=0 $Y2=0
cc_314 N_C_M1025_g N_VGND_c_1035_n 0.00454119f $X=3.945 $Y=0.655 $X2=0 $Y2=0
cc_315 N_C_M1030_g N_VGND_c_1035_n 0.004522f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_316 N_C_M1025_g N_VGND_c_1040_n 0.00486043f $X=3.945 $Y=0.655 $X2=0 $Y2=0
cc_317 N_C_M1030_g N_VGND_c_1040_n 0.00486043f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_318 N_C_M1025_g N_VGND_c_1041_n 5.83998e-19 $X=3.945 $Y=0.655 $X2=0 $Y2=0
cc_319 N_C_M1030_g N_VGND_c_1041_n 0.0125692f $X=4.375 $Y=0.655 $X2=0 $Y2=0
cc_320 N_B_M1017_g N_A_M1011_g 0.0240394f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_321 B N_A_M1002_g 5.33312e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_322 N_B_c_394_n N_A_M1002_g 0.0219037f $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_323 B N_A_c_486_n 6.41625e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_324 N_B_c_394_n N_A_c_486_n 0.0184638f $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_325 B N_A_c_489_n 0.0082195f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_326 N_B_c_394_n N_A_c_489_n 7.31414e-19 $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_327 N_B_M1026_g N_VPWR_c_562_n 0.00109252f $X=6.675 $Y=2.465 $X2=0 $Y2=0
cc_328 N_B_M1007_g N_VPWR_c_564_n 0.00357842f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_329 N_B_M1014_g N_VPWR_c_564_n 0.00357877f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_330 N_B_M1019_g N_VPWR_c_564_n 0.00357877f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_331 N_B_M1026_g N_VPWR_c_564_n 0.00357877f $X=6.675 $Y=2.465 $X2=0 $Y2=0
cc_332 N_B_M1007_g N_VPWR_c_560_n 0.00665087f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_333 N_B_M1014_g N_VPWR_c_560_n 0.0053512f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_334 N_B_M1019_g N_VPWR_c_560_n 0.0053512f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_335 N_B_M1026_g N_VPWR_c_560_n 0.00537654f $X=6.675 $Y=2.465 $X2=0 $Y2=0
cc_336 N_B_M1007_g N_A_217_367#_c_675_n 0.00106488f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_337 N_B_M1007_g N_Y_c_748_n 0.00103212f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_338 B N_Y_c_748_n 0.0157877f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_339 N_B_M1000_g N_Y_c_736_n 0.00458762f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_340 B N_Y_c_736_n 0.0248547f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_341 N_B_c_394_n N_Y_c_736_n 0.00123595f $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_342 N_B_M1003_g N_Y_c_737_n 0.0138758f $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_343 N_B_M1015_g N_Y_c_737_n 0.0138758f $X=6.165 $Y=0.655 $X2=0 $Y2=0
cc_344 B N_Y_c_737_n 0.0508543f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_345 N_B_c_394_n N_Y_c_737_n 0.00259007f $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_346 N_B_M1017_g N_Y_c_738_n 0.0152745f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_347 B N_Y_c_738_n 0.0112213f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_348 N_B_c_394_n N_Y_c_738_n 0.00337522f $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_349 B N_Y_c_741_n 0.0164475f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_350 N_B_c_394_n N_Y_c_741_n 0.00267671f $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_351 B Y 0.0164475f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_352 N_B_c_394_n Y 0.00267671f $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_353 N_B_M1000_g N_Y_c_745_n 0.0196361f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_354 B N_Y_c_745_n 0.0152595f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_355 N_B_M1007_g N_A_644_367#_c_905_n 0.0147239f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_356 B N_A_644_367#_c_905_n 0.0174046f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_357 N_B_c_394_n N_A_644_367#_c_905_n 2.86355e-19 $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_358 N_B_M1014_g N_A_644_367#_c_915_n 0.0133021f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_359 N_B_M1019_g N_A_644_367#_c_915_n 0.0114269f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_360 B N_A_644_367#_c_915_n 0.0391191f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_361 N_B_c_394_n N_A_644_367#_c_915_n 4.75711e-19 $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_362 B N_A_644_367#_c_919_n 0.0174054f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_363 N_B_c_394_n N_A_644_367#_c_919_n 5.36991e-19 $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_364 N_B_M1014_g N_A_644_367#_c_921_n 5.49585e-19 $X=5.815 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_B_M1019_g N_A_644_367#_c_921_n 0.00965218f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_366 N_B_M1026_g N_A_644_367#_c_921_n 0.00973616f $X=6.675 $Y=2.465 $X2=0
+ $Y2=0
cc_367 B N_A_644_367#_c_921_n 0.023857f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_368 N_B_c_394_n N_A_644_367#_c_921_n 5.36991e-19 $X=6.675 $Y=1.51 $X2=0 $Y2=0
cc_369 N_B_M1007_g N_A_1009_367#_c_950_n 0.00904346f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_370 N_B_M1014_g N_A_1009_367#_c_950_n 5.49585e-19 $X=5.815 $Y=2.465 $X2=0
+ $Y2=0
cc_371 N_B_M1007_g N_A_1009_367#_c_960_n 0.0105205f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_372 N_B_M1014_g N_A_1009_367#_c_960_n 0.012237f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_373 N_B_M1007_g N_A_1009_367#_c_951_n 5.81207e-19 $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_374 N_B_M1019_g N_A_1009_367#_c_963_n 0.0114565f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_375 N_B_M1026_g N_A_1009_367#_c_963_n 0.0114588f $X=6.675 $Y=2.465 $X2=0
+ $Y2=0
cc_376 N_B_M1026_g N_A_1009_367#_c_953_n 0.00114792f $X=6.675 $Y=2.465 $X2=0
+ $Y2=0
cc_377 B N_A_1009_367#_c_953_n 0.0123907f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_378 N_B_M1000_g N_VGND_c_1020_n 6.13597e-19 $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_379 N_B_M1003_g N_VGND_c_1020_n 0.0101747f $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_380 N_B_M1015_g N_VGND_c_1020_n 0.010177f $X=6.165 $Y=0.655 $X2=0 $Y2=0
cc_381 N_B_M1017_g N_VGND_c_1020_n 6.14008e-19 $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_382 N_B_M1015_g N_VGND_c_1021_n 6.14008e-19 $X=6.165 $Y=0.655 $X2=0 $Y2=0
cc_383 N_B_M1017_g N_VGND_c_1021_n 0.0101862f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_384 N_B_M1015_g N_VGND_c_1024_n 0.00486043f $X=6.165 $Y=0.655 $X2=0 $Y2=0
cc_385 N_B_M1017_g N_VGND_c_1024_n 0.00486043f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_386 N_B_M1000_g N_VGND_c_1033_n 0.00486043f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_387 N_B_M1003_g N_VGND_c_1033_n 0.00486043f $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_388 N_B_M1000_g N_VGND_c_1035_n 0.004522f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_389 N_B_M1003_g N_VGND_c_1035_n 0.00824727f $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_390 N_B_M1015_g N_VGND_c_1035_n 0.00824727f $X=6.165 $Y=0.655 $X2=0 $Y2=0
cc_391 N_B_M1017_g N_VGND_c_1035_n 0.00824727f $X=6.595 $Y=0.655 $X2=0 $Y2=0
cc_392 N_B_M1000_g N_VGND_c_1041_n 0.0125692f $X=5.305 $Y=0.655 $X2=0 $Y2=0
cc_393 N_B_M1003_g N_VGND_c_1041_n 5.83998e-19 $X=5.735 $Y=0.655 $X2=0 $Y2=0
cc_394 N_A_M1002_g N_VPWR_c_562_n 0.0153008f $X=7.105 $Y=2.465 $X2=0 $Y2=0
cc_395 N_A_M1010_g N_VPWR_c_562_n 0.0141279f $X=7.535 $Y=2.465 $X2=0 $Y2=0
cc_396 N_A_M1020_g N_VPWR_c_562_n 7.24342e-19 $X=7.965 $Y=2.465 $X2=0 $Y2=0
cc_397 N_A_M1010_g N_VPWR_c_563_n 7.24342e-19 $X=7.535 $Y=2.465 $X2=0 $Y2=0
cc_398 N_A_M1020_g N_VPWR_c_563_n 0.0141279f $X=7.965 $Y=2.465 $X2=0 $Y2=0
cc_399 N_A_M1032_g N_VPWR_c_563_n 0.0161027f $X=8.395 $Y=2.465 $X2=0 $Y2=0
cc_400 N_A_M1002_g N_VPWR_c_564_n 0.00486043f $X=7.105 $Y=2.465 $X2=0 $Y2=0
cc_401 N_A_M1010_g N_VPWR_c_566_n 0.00486043f $X=7.535 $Y=2.465 $X2=0 $Y2=0
cc_402 N_A_M1020_g N_VPWR_c_566_n 0.00486043f $X=7.965 $Y=2.465 $X2=0 $Y2=0
cc_403 N_A_M1032_g N_VPWR_c_569_n 0.00486043f $X=8.395 $Y=2.465 $X2=0 $Y2=0
cc_404 N_A_M1002_g N_VPWR_c_560_n 0.0082726f $X=7.105 $Y=2.465 $X2=0 $Y2=0
cc_405 N_A_M1010_g N_VPWR_c_560_n 0.00824727f $X=7.535 $Y=2.465 $X2=0 $Y2=0
cc_406 N_A_M1020_g N_VPWR_c_560_n 0.00824727f $X=7.965 $Y=2.465 $X2=0 $Y2=0
cc_407 N_A_M1032_g N_VPWR_c_560_n 0.00934593f $X=8.395 $Y=2.465 $X2=0 $Y2=0
cc_408 N_A_M1011_g N_Y_c_738_n 0.0134196f $X=7.035 $Y=0.655 $X2=0 $Y2=0
cc_409 N_A_c_489_n N_Y_c_738_n 0.0127274f $X=7.735 $Y=1.367 $X2=0 $Y2=0
cc_410 N_A_M1013_g N_Y_c_833_n 0.0135911f $X=7.495 $Y=0.655 $X2=0 $Y2=0
cc_411 N_A_M1022_g N_Y_c_833_n 0.0122595f $X=7.925 $Y=0.655 $X2=0 $Y2=0
cc_412 A N_Y_c_833_n 0.0153383f $X=8.795 $Y=1.21 $X2=0 $Y2=0
cc_413 N_A_c_486_n N_Y_c_833_n 0.00262887f $X=8.47 $Y=1.44 $X2=0 $Y2=0
cc_414 N_A_c_488_n N_Y_c_833_n 0.019322f $X=7.892 $Y=1.367 $X2=0 $Y2=0
cc_415 N_A_c_489_n N_Y_c_833_n 0.0118843f $X=7.735 $Y=1.367 $X2=0 $Y2=0
cc_416 N_A_M1011_g N_Y_c_742_n 2.96597e-19 $X=7.035 $Y=0.655 $X2=0 $Y2=0
cc_417 N_A_M1013_g N_Y_c_742_n 0.00412222f $X=7.495 $Y=0.655 $X2=0 $Y2=0
cc_418 N_A_M1022_g N_Y_c_742_n 7.60284e-19 $X=7.925 $Y=0.655 $X2=0 $Y2=0
cc_419 N_A_c_486_n N_Y_c_742_n 0.00363906f $X=8.47 $Y=1.44 $X2=0 $Y2=0
cc_420 N_A_c_489_n N_Y_c_742_n 0.0221657f $X=7.735 $Y=1.367 $X2=0 $Y2=0
cc_421 N_A_M1002_g N_A_1009_367#_c_952_n 0.0153483f $X=7.105 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_M1010_g N_A_1009_367#_c_952_n 0.0156683f $X=7.535 $Y=2.465 $X2=0
+ $Y2=0
cc_423 N_A_c_486_n N_A_1009_367#_c_952_n 0.00396342f $X=8.47 $Y=1.44 $X2=0 $Y2=0
cc_424 N_A_c_489_n N_A_1009_367#_c_952_n 0.0478599f $X=7.735 $Y=1.367 $X2=0
+ $Y2=0
cc_425 N_A_c_486_n N_A_1009_367#_c_953_n 7.49468e-19 $X=8.47 $Y=1.44 $X2=0 $Y2=0
cc_426 N_A_c_489_n N_A_1009_367#_c_953_n 0.00201686f $X=7.735 $Y=1.367 $X2=0
+ $Y2=0
cc_427 N_A_M1020_g N_A_1009_367#_c_954_n 0.0157315f $X=7.965 $Y=2.465 $X2=0
+ $Y2=0
cc_428 N_A_M1032_g N_A_1009_367#_c_954_n 0.0168713f $X=8.395 $Y=2.465 $X2=0
+ $Y2=0
cc_429 A N_A_1009_367#_c_954_n 0.0218546f $X=8.795 $Y=1.21 $X2=0 $Y2=0
cc_430 N_A_c_486_n N_A_1009_367#_c_954_n 0.00265527f $X=8.47 $Y=1.44 $X2=0 $Y2=0
cc_431 N_A_c_487_n N_A_1009_367#_c_954_n 0.00776841f $X=8.825 $Y=1.44 $X2=0
+ $Y2=0
cc_432 N_A_c_488_n N_A_1009_367#_c_954_n 0.0500405f $X=7.892 $Y=1.367 $X2=0
+ $Y2=0
cc_433 N_A_c_486_n N_A_1009_367#_c_956_n 0.0027397f $X=8.47 $Y=1.44 $X2=0 $Y2=0
cc_434 N_A_c_489_n N_A_1009_367#_c_956_n 0.0156687f $X=7.735 $Y=1.367 $X2=0
+ $Y2=0
cc_435 N_A_M1011_g N_VGND_c_1021_n 0.00947683f $X=7.035 $Y=0.655 $X2=0 $Y2=0
cc_436 N_A_M1013_g N_VGND_c_1021_n 5.86791e-19 $X=7.495 $Y=0.655 $X2=0 $Y2=0
cc_437 N_A_M1011_g N_VGND_c_1022_n 5.66286e-19 $X=7.035 $Y=0.655 $X2=0 $Y2=0
cc_438 N_A_M1013_g N_VGND_c_1022_n 0.0102049f $X=7.495 $Y=0.655 $X2=0 $Y2=0
cc_439 N_A_M1022_g N_VGND_c_1022_n 0.0100888f $X=7.925 $Y=0.655 $X2=0 $Y2=0
cc_440 N_A_M1028_g N_VGND_c_1022_n 5.75816e-19 $X=8.355 $Y=0.655 $X2=0 $Y2=0
cc_441 N_A_M1022_g N_VGND_c_1023_n 6.24191e-19 $X=7.925 $Y=0.655 $X2=0 $Y2=0
cc_442 N_A_M1028_g N_VGND_c_1023_n 0.0165374f $X=8.355 $Y=0.655 $X2=0 $Y2=0
cc_443 A N_VGND_c_1023_n 0.0256422f $X=8.795 $Y=1.21 $X2=0 $Y2=0
cc_444 N_A_c_486_n N_VGND_c_1023_n 0.00187306f $X=8.47 $Y=1.44 $X2=0 $Y2=0
cc_445 N_A_M1011_g N_VGND_c_1026_n 0.00525069f $X=7.035 $Y=0.655 $X2=0 $Y2=0
cc_446 N_A_M1013_g N_VGND_c_1026_n 0.00486043f $X=7.495 $Y=0.655 $X2=0 $Y2=0
cc_447 N_A_M1022_g N_VGND_c_1028_n 0.00486043f $X=7.925 $Y=0.655 $X2=0 $Y2=0
cc_448 N_A_M1028_g N_VGND_c_1028_n 0.00486043f $X=8.355 $Y=0.655 $X2=0 $Y2=0
cc_449 N_A_M1011_g N_VGND_c_1035_n 0.00894125f $X=7.035 $Y=0.655 $X2=0 $Y2=0
cc_450 N_A_M1013_g N_VGND_c_1035_n 0.00832343f $X=7.495 $Y=0.655 $X2=0 $Y2=0
cc_451 N_A_M1022_g N_VGND_c_1035_n 0.00824727f $X=7.925 $Y=0.655 $X2=0 $Y2=0
cc_452 N_A_M1028_g N_VGND_c_1035_n 0.00824727f $X=8.355 $Y=0.655 $X2=0 $Y2=0
cc_453 N_VPWR_c_560_n N_A_217_367#_M1005_s 0.00249949f $X=8.88 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_454 N_VPWR_c_560_n N_A_217_367#_M1006_s 0.00223565f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_560_n N_A_217_367#_M1031_s 0.00223565f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_560_n N_A_217_367#_M1012_d 0.00223564f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_560_n N_A_217_367#_M1023_d 0.00215158f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_561_n N_A_217_367#_c_698_n 0.0114889f $X=0.69 $Y=2.4 $X2=0 $Y2=0
cc_459 N_VPWR_c_564_n N_A_217_367#_c_698_n 0.0143128f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_560_n N_A_217_367#_c_698_n 0.00815375f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_561_n N_A_217_367#_c_673_n 0.039213f $X=0.69 $Y=2.4 $X2=0 $Y2=0
cc_462 N_VPWR_c_564_n N_A_217_367#_c_682_n 0.0361172f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_560_n N_A_217_367#_c_682_n 0.023676f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_464 N_VPWR_c_564_n N_A_217_367#_c_684_n 0.0361172f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_560_n N_A_217_367#_c_684_n 0.023676f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_466 N_VPWR_c_564_n N_A_217_367#_c_686_n 0.0361172f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_560_n N_A_217_367#_c_686_n 0.023676f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_468 N_VPWR_c_564_n N_A_217_367#_c_674_n 0.0539065f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_560_n N_A_217_367#_c_674_n 0.0335145f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_564_n N_A_217_367#_c_710_n 0.0125234f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_560_n N_A_217_367#_c_710_n 0.00738676f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_564_n N_A_217_367#_c_712_n 0.0125234f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_560_n N_A_217_367#_c_712_n 0.00738676f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_564_n N_A_217_367#_c_714_n 0.0129275f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_560_n N_A_217_367#_c_714_n 0.00778723f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_560_n N_Y_M1005_d 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_c_560_n N_Y_M1018_d 0.00225186f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_478 N_VPWR_c_560_n N_A_644_367#_M1008_s 0.00225186f $X=8.88 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_479 N_VPWR_c_560_n N_A_644_367#_M1021_s 0.00225186f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_560_n N_A_644_367#_M1007_s 0.00225186f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_560_n N_A_644_367#_M1019_s 0.00225186f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_560_n N_A_1009_367#_M1007_d 0.00215158f $X=8.88 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_483 N_VPWR_c_560_n N_A_1009_367#_M1014_d 0.00223562f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_560_n N_A_1009_367#_M1026_d 0.00376627f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_560_n N_A_1009_367#_M1010_s 0.00536646f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_560_n N_A_1009_367#_M1032_s 0.00371702f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_564_n N_A_1009_367#_c_960_n 0.0317578f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_560_n N_A_1009_367#_c_960_n 0.0199132f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_564_n N_A_1009_367#_c_951_n 0.021267f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_560_n N_A_1009_367#_c_951_n 0.0126613f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_564_n N_A_1009_367#_c_963_n 0.0361172f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_560_n N_A_1009_367#_c_963_n 0.023676f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_564_n N_A_1009_367#_c_992_n 0.0125234f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_560_n N_A_1009_367#_c_992_n 0.00738676f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_495 N_VPWR_M1002_d N_A_1009_367#_c_952_n 0.00182444f $X=7.18 $Y=1.835 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_562_n N_A_1009_367#_c_952_n 0.0166945f $X=7.32 $Y=2.19 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_566_n N_A_1009_367#_c_996_n 0.0124525f $X=8.015 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_560_n N_A_1009_367#_c_996_n 0.00730901f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_M1020_d N_A_1009_367#_c_954_n 0.00182444f $X=8.04 $Y=1.835 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_563_n N_A_1009_367#_c_954_n 0.0166945f $X=8.18 $Y=2.19 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_569_n N_A_1009_367#_c_955_n 0.0178111f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_560_n N_A_1009_367#_c_955_n 0.0100304f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_564_n N_A_1009_367#_c_1002_n 0.0138145f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_560_n N_A_1009_367#_c_1002_n 0.00876065f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_505 N_A_217_367#_c_682_n N_Y_M1005_d 0.00332344f $X=1.975 $Y=2.99 $X2=0 $Y2=0
cc_506 N_A_217_367#_c_684_n N_Y_M1018_d 0.00332344f $X=2.835 $Y=2.99 $X2=0 $Y2=0
cc_507 N_A_217_367#_c_682_n N_Y_c_759_n 0.0159805f $X=1.975 $Y=2.99 $X2=0 $Y2=0
cc_508 N_A_217_367#_c_719_p N_Y_c_746_n 0.0145583f $X=2.07 $Y=2.17 $X2=0 $Y2=0
cc_509 N_A_217_367#_c_673_n N_Y_c_747_n 0.00158375f $X=1.21 $Y=1.98 $X2=0 $Y2=0
cc_510 N_A_217_367#_c_684_n N_Y_c_774_n 0.0159805f $X=2.835 $Y=2.99 $X2=0 $Y2=0
cc_511 N_A_217_367#_c_722_p N_Y_c_748_n 0.0145583f $X=2.93 $Y=2.17 $X2=0 $Y2=0
cc_512 N_A_217_367#_c_686_n N_A_644_367#_M1008_s 0.00332344f $X=3.695 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_513 N_A_217_367#_c_674_n N_A_644_367#_M1021_s 0.00332344f $X=4.485 $Y=2.99
+ $X2=0 $Y2=0
cc_514 N_A_217_367#_M1012_d N_A_644_367#_c_906_n 0.00340214f $X=3.65 $Y=1.835
+ $X2=0 $Y2=0
cc_515 N_A_217_367#_c_726_p N_A_644_367#_c_906_n 0.0136211f $X=3.79 $Y=2.52
+ $X2=0 $Y2=0
cc_516 N_A_217_367#_c_674_n N_A_644_367#_c_934_n 0.0126348f $X=4.485 $Y=2.99
+ $X2=0 $Y2=0
cc_517 N_A_217_367#_M1023_d N_A_644_367#_c_905_n 0.00508977f $X=4.51 $Y=1.835
+ $X2=0 $Y2=0
cc_518 N_A_217_367#_c_675_n N_A_644_367#_c_905_n 0.0221917f $X=4.65 $Y=2.46
+ $X2=0 $Y2=0
cc_519 N_A_217_367#_c_686_n N_A_644_367#_c_909_n 0.0159805f $X=3.695 $Y=2.99
+ $X2=0 $Y2=0
cc_520 N_A_217_367#_c_675_n N_A_1009_367#_c_950_n 0.0422743f $X=4.65 $Y=2.46
+ $X2=0 $Y2=0
cc_521 N_A_217_367#_c_674_n N_A_1009_367#_c_951_n 0.0147157f $X=4.485 $Y=2.99
+ $X2=0 $Y2=0
cc_522 N_Y_c_748_n N_A_644_367#_c_906_n 0.036594f $X=4.87 $Y=1.75 $X2=0 $Y2=0
cc_523 N_Y_c_748_n N_A_644_367#_c_905_n 0.0526323f $X=4.87 $Y=1.75 $X2=0 $Y2=0
cc_524 N_Y_c_748_n N_A_644_367#_c_909_n 0.0217611f $X=4.87 $Y=1.75 $X2=0 $Y2=0
cc_525 N_Y_c_748_n N_A_644_367#_c_941_n 0.0150119f $X=4.87 $Y=1.75 $X2=0 $Y2=0
cc_526 N_Y_c_738_n N_A_1009_367#_c_953_n 0.00652243f $X=7.145 $Y=1.095 $X2=0
+ $Y2=0
cc_527 N_Y_c_733_n N_VGND_M1009_d 0.00230018f $X=1.965 $Y=1.055 $X2=0 $Y2=0
cc_528 N_Y_c_735_n N_VGND_M1029_d 0.00725728f $X=3.205 $Y=1.055 $X2=0 $Y2=0
cc_529 N_Y_c_805_n N_VGND_M1016_d 0.00365904f $X=4.065 $Y=0.94 $X2=0 $Y2=0
cc_530 Y N_VGND_M1030_d 0.00500207f $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_531 N_Y_c_810_n N_VGND_M1030_d 0.0113247f $X=4.87 $Y=0.94 $X2=0 $Y2=0
cc_532 N_Y_c_745_n N_VGND_M1030_d 0.00120318f $X=5.425 $Y=1.012 $X2=0 $Y2=0
cc_533 N_Y_c_737_n N_VGND_M1003_s 0.00176773f $X=6.285 $Y=1.095 $X2=0 $Y2=0
cc_534 N_Y_c_738_n N_VGND_M1017_s 0.00187422f $X=7.145 $Y=1.095 $X2=0 $Y2=0
cc_535 N_Y_c_833_n N_VGND_M1013_d 0.00362687f $X=8.045 $Y=0.955 $X2=0 $Y2=0
cc_536 N_Y_c_733_n N_VGND_c_1016_n 0.0179051f $X=1.965 $Y=1.055 $X2=0 $Y2=0
cc_537 N_Y_c_735_n N_VGND_c_1017_n 0.0438043f $X=3.205 $Y=1.055 $X2=0 $Y2=0
cc_538 N_Y_c_869_p N_VGND_c_1018_n 0.0124525f $X=3.3 $Y=0.42 $X2=0 $Y2=0
cc_539 N_Y_c_805_n N_VGND_c_1019_n 0.0168833f $X=4.065 $Y=0.94 $X2=0 $Y2=0
cc_540 N_Y_c_737_n N_VGND_c_1020_n 0.0171443f $X=6.285 $Y=1.095 $X2=0 $Y2=0
cc_541 N_Y_c_738_n N_VGND_c_1021_n 0.0171962f $X=7.145 $Y=1.095 $X2=0 $Y2=0
cc_542 N_Y_c_833_n N_VGND_c_1022_n 0.0170777f $X=8.045 $Y=0.955 $X2=0 $Y2=0
cc_543 N_Y_c_874_p N_VGND_c_1024_n 0.0124525f $X=6.38 $Y=0.42 $X2=0 $Y2=0
cc_544 N_Y_c_875_p N_VGND_c_1026_n 0.0149167f $X=7.26 $Y=0.42 $X2=0 $Y2=0
cc_545 N_Y_c_876_p N_VGND_c_1028_n 0.0124525f $X=8.14 $Y=0.42 $X2=0 $Y2=0
cc_546 N_Y_c_877_p N_VGND_c_1031_n 0.0128073f $X=1.18 $Y=0.42 $X2=0 $Y2=0
cc_547 N_Y_c_878_p N_VGND_c_1032_n 0.0135169f $X=2.09 $Y=0.42 $X2=0 $Y2=0
cc_548 N_Y_c_879_p N_VGND_c_1033_n 0.0124525f $X=5.52 $Y=0.42 $X2=0 $Y2=0
cc_549 N_Y_M1004_s N_VGND_c_1035_n 0.00501859f $X=1.04 $Y=0.235 $X2=0 $Y2=0
cc_550 N_Y_M1024_s N_VGND_c_1035_n 0.00432284f $X=1.95 $Y=0.235 $X2=0 $Y2=0
cc_551 N_Y_M1001_s N_VGND_c_1035_n 0.00408468f $X=3.16 $Y=0.235 $X2=0 $Y2=0
cc_552 N_Y_M1025_s N_VGND_c_1035_n 0.0028032f $X=4.02 $Y=0.235 $X2=0 $Y2=0
cc_553 N_Y_M1000_d N_VGND_c_1035_n 0.00408483f $X=5.38 $Y=0.235 $X2=0 $Y2=0
cc_554 N_Y_M1015_d N_VGND_c_1035_n 0.00536646f $X=6.24 $Y=0.235 $X2=0 $Y2=0
cc_555 N_Y_M1011_s N_VGND_c_1035_n 0.00525984f $X=7.11 $Y=0.235 $X2=0 $Y2=0
cc_556 N_Y_M1022_s N_VGND_c_1035_n 0.00536646f $X=8 $Y=0.235 $X2=0 $Y2=0
cc_557 N_Y_c_877_p N_VGND_c_1035_n 0.0076925f $X=1.18 $Y=0.42 $X2=0 $Y2=0
cc_558 N_Y_c_878_p N_VGND_c_1035_n 0.00847534f $X=2.09 $Y=0.42 $X2=0 $Y2=0
cc_559 N_Y_c_869_p N_VGND_c_1035_n 0.00730901f $X=3.3 $Y=0.42 $X2=0 $Y2=0
cc_560 N_Y_c_874_p N_VGND_c_1035_n 0.00730901f $X=6.38 $Y=0.42 $X2=0 $Y2=0
cc_561 N_Y_c_875_p N_VGND_c_1035_n 0.00886411f $X=7.26 $Y=0.42 $X2=0 $Y2=0
cc_562 N_Y_c_876_p N_VGND_c_1035_n 0.00730901f $X=8.14 $Y=0.42 $X2=0 $Y2=0
cc_563 N_Y_c_740_n N_VGND_c_1035_n 3.64927e-19 $X=3.3 $Y=0.93 $X2=0 $Y2=0
cc_564 Y N_VGND_c_1035_n 6.9347e-19 $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_565 N_Y_c_805_n N_VGND_c_1035_n 0.0107119f $X=4.065 $Y=0.94 $X2=0 $Y2=0
cc_566 N_Y_c_810_n N_VGND_c_1035_n 0.00641882f $X=4.87 $Y=0.94 $X2=0 $Y2=0
cc_567 N_Y_c_745_n N_VGND_c_1035_n 0.0059104f $X=5.425 $Y=1.012 $X2=0 $Y2=0
cc_568 N_Y_c_899_p N_VGND_c_1035_n 0.00730901f $X=4.16 $Y=0.42 $X2=0 $Y2=0
cc_569 N_Y_c_879_p N_VGND_c_1035_n 0.00730901f $X=5.52 $Y=0.42 $X2=0 $Y2=0
cc_570 N_Y_c_899_p N_VGND_c_1040_n 0.0124525f $X=4.16 $Y=0.42 $X2=0 $Y2=0
cc_571 Y N_VGND_c_1041_n 0.0166368f $X=4.955 $Y=0.84 $X2=0 $Y2=0
cc_572 N_Y_c_810_n N_VGND_c_1041_n 0.0308534f $X=4.87 $Y=0.94 $X2=0 $Y2=0
cc_573 N_Y_c_745_n N_VGND_c_1041_n 0.0112499f $X=5.425 $Y=1.012 $X2=0 $Y2=0
cc_574 N_A_644_367#_c_905_n N_A_1009_367#_M1007_d 0.00994881f $X=5.505 $Y=2.095
+ $X2=-0.19 $Y2=1.655
cc_575 N_A_644_367#_c_915_n N_A_1009_367#_M1014_d 0.00336413f $X=6.295 $Y=2.095
+ $X2=0 $Y2=0
cc_576 N_A_644_367#_c_905_n N_A_1009_367#_c_950_n 0.0221917f $X=5.505 $Y=2.095
+ $X2=0 $Y2=0
cc_577 N_A_644_367#_M1007_s N_A_1009_367#_c_960_n 0.00332344f $X=5.46 $Y=1.835
+ $X2=0 $Y2=0
cc_578 N_A_644_367#_c_946_p N_A_1009_367#_c_960_n 0.0126348f $X=5.6 $Y=2.57
+ $X2=0 $Y2=0
cc_579 N_A_644_367#_c_915_n N_A_1009_367#_c_1012_n 0.0136211f $X=6.295 $Y=2.095
+ $X2=0 $Y2=0
cc_580 N_A_644_367#_M1019_s N_A_1009_367#_c_963_n 0.00332344f $X=6.32 $Y=1.835
+ $X2=0 $Y2=0
cc_581 N_A_644_367#_c_921_n N_A_1009_367#_c_963_n 0.0159805f $X=6.46 $Y=2.1
+ $X2=0 $Y2=0
