* NGSPICE file created from sky130_fd_sc_lp__fahcin_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
M1000 a_364_73# B a_256_87# VNB nshort w=640000u l=150000u
+  ad=5.5115e+11p pd=4.88e+06u as=5.216e+11p ps=4.19e+06u
M1001 SUM a_1926_135# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=1.8946e+12p ps=1.185e+07u
M1002 a_29_47# a_439_47# a_555_73# VPB phighvt w=840000u l=150000u
+  ad=8.127e+11p pd=5.85e+06u as=4.69e+11p ps=2.98e+06u
M1003 VPWR CIN a_1500_63# VPB phighvt w=1e+06u l=150000u
+  ad=2.5664e+12p pd=1.462e+07u as=3.774e+11p ps=2.79e+06u
M1004 VGND B a_439_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1005 a_256_87# a_29_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_555_73# B a_29_47# VNB nshort w=640000u l=150000u
+  ad=3.481e+11p pd=2.9e+06u as=4.186e+11p ps=4.09e+06u
M1007 a_256_87# a_29_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=5.202e+11p pd=4.81e+06u as=0p ps=0u
M1008 a_1500_63# a_555_73# COUT VNB nshort w=640000u l=150000u
+  ad=3.456e+11p pd=2.36e+06u as=6.656e+11p ps=3.36e+06u
M1009 a_256_87# a_439_47# a_555_73# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_555_73# B a_256_87# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND CIN a_1500_63# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_29_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B a_439_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.591e+11p ps=3.09e+06u
M1014 a_364_73# B a_29_47# VPB phighvt w=840000u l=150000u
+  ad=4.872e+11p pd=4.52e+06u as=0p ps=0u
M1015 a_1152_389# a_439_47# VGND VNB nshort w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1016 VGND A a_29_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_1774_367# a_1883_395# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.496e+11p ps=2.46e+06u
M1018 SUM a_1926_135# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1019 a_1152_389# a_439_47# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=3.774e+11p pd=2.79e+06u as=0p ps=0u
M1020 a_1926_135# a_555_73# a_1883_395# VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=5.152e+11p ps=4.8e+06u
M1021 a_256_87# a_439_47# a_364_73# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1774_367# CIN VGND VNB nshort w=840000u l=150000u
+  ad=3.252e+11p pd=2.79e+06u as=0p ps=0u
M1023 a_1774_367# CIN VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.385e+11p pd=5.99e+06u as=0p ps=0u
M1024 a_1774_367# a_364_73# a_1926_135# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1774_367# a_1883_395# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_29_47# a_439_47# a_364_73# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 COUT a_364_73# a_1152_389# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1883_395# a_364_73# a_1926_135# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=3.52e+11p ps=2.38e+06u
M1029 a_1500_63# a_364_73# COUT VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=8.988e+11p ps=3.82e+06u
M1030 COUT a_555_73# a_1152_389# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1926_135# a_555_73# a_1774_367# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

