* File: sky130_fd_sc_lp__or2b_2.spice
* Created: Fri Aug 28 11:22:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2b_2.pex.spice"
.subckt sky130_fd_sc_lp__or2b_2  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_B_N_M1001_g N_A_27_49#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.118433 AS=0.1113 PD=0.926667 PS=1.37 NRD=24.276 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_191_254#_M1000_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.236867 PD=1.12 PS=1.85333 NRD=0 NRS=12.132 M=1 R=5.6 SA=75000.5
+ SB=75001.4 A=0.126 P=1.98 MULT=1
MM1003 N_X_M1000_d N_A_191_254#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.262067 PD=1.12 PS=1.92667 NRD=0 NRS=12.132 M=1 R=5.6 SA=75000.9
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1004 N_A_191_254#_M1004_d N_A_M1004_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.131033 PD=0.81 PS=0.963333 NRD=0 NRS=73.416 M=1 R=2.8
+ SA=75001.3 SB=75001 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_27_49#_M1009_g N_A_191_254#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.2373 AS=0.0819 PD=1.97 PS=0.81 NRD=85.704 NRS=31.428 M=1 R=2.8
+ SA=75001.9 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_B_N_M1005_g N_A_27_49#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09135 AS=0.1197 PD=0.8 PS=1.41 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1005_d N_A_191_254#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.27405 AS=0.1764 PD=2.4 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4 SB=75001
+ A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A_191_254#_M1008_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.1764 PD=2.955 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 A_479_367# N_A_M1006_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.1302 PD=0.63 PS=0.985 NRD=23.443 NRS=119.599 M=1 R=2.8 SA=75002
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_191_254#_M1007_d N_A_27_49#_M1007_g A_479_367# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75002.3 SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__or2b_2.pxi.spice"
*
.ends
*
*
