* File: sky130_fd_sc_lp__clkinvlp_4.pxi.spice
* Created: Wed Sep  2 09:41:19 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINVLP_4%A N_A_M1007_g N_A_M1000_g N_A_M1001_g
+ N_A_M1002_g N_A_M1003_g N_A_M1004_g N_A_M1006_g N_A_M1005_g A A N_A_c_48_n
+ PM_SKY130_FD_SC_LP__CLKINVLP_4%A
x_PM_SKY130_FD_SC_LP__CLKINVLP_4%VPWR N_VPWR_M1000_s N_VPWR_M1002_s
+ N_VPWR_M1005_s N_VPWR_c_109_n N_VPWR_c_110_n N_VPWR_c_111_n N_VPWR_c_112_n
+ N_VPWR_c_113_n N_VPWR_c_114_n N_VPWR_c_115_n VPWR N_VPWR_c_116_n
+ N_VPWR_c_108_n N_VPWR_c_118_n PM_SKY130_FD_SC_LP__CLKINVLP_4%VPWR
x_PM_SKY130_FD_SC_LP__CLKINVLP_4%Y N_Y_M1001_d N_Y_M1000_d N_Y_M1004_d
+ N_Y_c_147_n N_Y_c_150_n N_Y_c_148_n Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__CLKINVLP_4%Y
x_PM_SKY130_FD_SC_LP__CLKINVLP_4%VGND N_VGND_M1007_s N_VGND_M1006_s
+ N_VGND_c_188_n N_VGND_c_189_n N_VGND_c_190_n VGND N_VGND_c_191_n
+ N_VGND_c_192_n N_VGND_c_193_n N_VGND_c_194_n
+ PM_SKY130_FD_SC_LP__CLKINVLP_4%VGND
cc_1 VNB N_A_M1007_g 0.0369914f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.61
cc_2 VNB N_A_M1000_g 0.00506355f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.48
cc_3 VNB N_A_M1001_g 0.0244485f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.61
cc_4 VNB N_A_M1002_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.48
cc_5 VNB N_A_M1003_g 0.0275159f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=0.61
cc_6 VNB N_A_M1004_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.48
cc_7 VNB N_A_M1006_g 0.0394314f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=0.61
cc_8 VNB N_A_M1005_g 0.00795919f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.48
cc_9 VNB A 0.0243288f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_A_c_48_n 0.151635f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.407
cc_11 VNB N_VPWR_c_108_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.407
cc_12 VNB N_Y_c_147_n 0.00479344f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.61
cc_13 VNB N_Y_c_148_n 0.00345438f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.48
cc_14 VNB Y 0.00674419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_188_n 0.0111239f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.48
cc_16 VNB N_VGND_c_189_n 0.0257259f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.235
cc_17 VNB N_VGND_c_190_n 0.0255131f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.565
cc_18 VNB N_VGND_c_191_n 0.0340106f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.235
cc_19 VNB N_VGND_c_192_n 0.0299875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_193_n 0.214098f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.235
cc_21 VNB N_VGND_c_194_n 0.00589254f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.48
cc_22 VPB N_A_M1000_g 0.0435143f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.48
cc_23 VPB N_A_M1002_g 0.0340581f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.48
cc_24 VPB N_A_M1004_g 0.0340581f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.48
cc_25 VPB N_A_M1005_g 0.0461397f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.48
cc_26 VPB A 0.00764565f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_27 VPB N_VPWR_c_109_n 0.0112117f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.61
cc_28 VPB N_VPWR_c_110_n 0.0508745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_111_n 0.0199224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_112_n 0.00678226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_113_n 0.0608249f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=0.61
cc_32 VPB N_VPWR_c_114_n 0.0199224f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.48
cc_33 VPB N_VPWR_c_115_n 0.00598038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_116_n 0.0128037f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.407
cc_35 VPB N_VPWR_c_108_n 0.057395f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.407
cc_36 VPB N_VPWR_c_118_n 0.00577233f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=1.407
cc_37 VPB N_Y_c_150_n 0.00232136f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.48
cc_38 VPB Y 0.00232136f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=0.61
cc_39 N_A_M1000_g N_VPWR_c_110_n 0.0235557f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_40 N_A_M1002_g N_VPWR_c_110_n 8.05893e-19 $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_41 A N_VPWR_c_110_n 0.0288185f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_42 N_A_c_48_n N_VPWR_c_110_n 0.00122665f $X=1.625 $Y=1.407 $X2=0 $Y2=0
cc_43 N_A_M1000_g N_VPWR_c_111_n 0.00687065f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_44 N_A_M1002_g N_VPWR_c_111_n 0.00687065f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_45 N_A_M1000_g N_VPWR_c_112_n 8.05893e-19 $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_46 N_A_M1002_g N_VPWR_c_112_n 0.0225326f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_47 N_A_M1004_g N_VPWR_c_112_n 0.0225326f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_48 N_A_M1005_g N_VPWR_c_112_n 8.05893e-19 $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_49 N_A_c_48_n N_VPWR_c_112_n 0.00233601f $X=1.625 $Y=1.407 $X2=0 $Y2=0
cc_50 N_A_M1004_g N_VPWR_c_113_n 8.05893e-19 $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_51 N_A_M1005_g N_VPWR_c_113_n 0.0244443f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_52 N_A_M1004_g N_VPWR_c_114_n 0.00687065f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_53 N_A_M1005_g N_VPWR_c_114_n 0.00687065f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_54 N_A_M1000_g N_VPWR_c_108_n 0.0129282f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_55 N_A_M1002_g N_VPWR_c_108_n 0.0129282f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_56 N_A_M1004_g N_VPWR_c_108_n 0.0129282f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_57 N_A_M1005_g N_VPWR_c_108_n 0.0129282f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_58 N_A_c_48_n N_Y_c_147_n 0.104708f $X=1.625 $Y=1.407 $X2=0 $Y2=0
cc_59 N_A_M1002_g N_Y_c_150_n 0.00197414f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_60 N_A_M1004_g N_Y_c_150_n 0.0308281f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_61 N_A_M1005_g N_Y_c_150_n 0.0411856f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_62 N_A_M1007_g N_Y_c_148_n 0.0034335f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_63 N_A_M1001_g N_Y_c_148_n 0.0116329f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_64 N_A_M1003_g N_Y_c_148_n 0.00898912f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_65 N_A_M1006_g N_Y_c_148_n 0.00126558f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_66 N_A_c_48_n N_Y_c_148_n 0.00225966f $X=1.625 $Y=1.407 $X2=0 $Y2=0
cc_67 N_A_M1007_g Y 0.00909638f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_68 N_A_M1001_g Y 0.0117107f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_69 N_A_M1003_g Y 0.0078929f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_70 A Y 0.0102621f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 A Y 0.026482f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_c_48_n Y 0.0182148f $X=1.625 $Y=1.407 $X2=0 $Y2=0
cc_73 N_A_M1000_g Y 0.0347043f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_74 N_A_M1002_g Y 0.0308281f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_75 N_A_M1004_g Y 0.00197414f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_76 A Y 0.0161123f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_48_n Y 3.96106e-19 $X=1.625 $Y=1.407 $X2=0 $Y2=0
cc_78 N_A_M1007_g N_VGND_c_189_n 0.0121806f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_79 N_A_M1001_g N_VGND_c_189_n 0.0010716f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_80 A N_VGND_c_189_n 0.016704f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_c_48_n N_VGND_c_189_n 0.00118321f $X=1.625 $Y=1.407 $X2=0 $Y2=0
cc_82 N_A_M1003_g N_VGND_c_190_n 0.00194234f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_83 N_A_M1006_g N_VGND_c_190_n 0.0147015f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_84 N_A_c_48_n N_VGND_c_190_n 0.00181815f $X=1.625 $Y=1.407 $X2=0 $Y2=0
cc_85 N_A_M1007_g N_VGND_c_191_n 0.00407525f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_86 N_A_M1001_g N_VGND_c_191_n 0.00306316f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_87 N_A_M1003_g N_VGND_c_191_n 0.00460068f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_88 N_A_M1006_g N_VGND_c_191_n 0.00407525f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_89 N_A_M1007_g N_VGND_c_193_n 0.00774993f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_90 N_A_M1001_g N_VGND_c_193_n 0.00413202f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_91 N_A_M1003_g N_VGND_c_193_n 0.00874311f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_92 N_A_M1006_g N_VGND_c_193_n 0.00774993f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_93 N_VPWR_c_112_n N_Y_c_147_n 0.0145538f $X=1.32 $Y=2.125 $X2=0 $Y2=0
cc_94 N_VPWR_c_112_n N_Y_c_150_n 0.0685263f $X=1.32 $Y=2.125 $X2=0 $Y2=0
cc_95 N_VPWR_c_113_n N_Y_c_150_n 0.0685263f $X=2.38 $Y=2.125 $X2=0 $Y2=0
cc_96 N_VPWR_c_114_n N_Y_c_150_n 0.0157615f $X=2.215 $Y=3.33 $X2=0 $Y2=0
cc_97 N_VPWR_c_108_n N_Y_c_150_n 0.0120285f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_98 N_VPWR_c_110_n Y 0.0685263f $X=0.26 $Y=2.125 $X2=0 $Y2=0
cc_99 N_VPWR_c_111_n Y 0.0157615f $X=1.155 $Y=3.33 $X2=0 $Y2=0
cc_100 N_VPWR_c_112_n Y 0.0685263f $X=1.32 $Y=2.125 $X2=0 $Y2=0
cc_101 N_VPWR_c_108_n Y 0.0120285f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_102 N_Y_c_148_n N_VGND_c_189_n 0.0330838f $X=1.05 $Y=0.545 $X2=0 $Y2=0
cc_103 N_Y_c_147_n N_VGND_c_190_n 0.0119351f $X=1.685 $Y=1.4 $X2=0 $Y2=0
cc_104 N_Y_c_148_n N_VGND_c_190_n 0.0161046f $X=1.05 $Y=0.545 $X2=0 $Y2=0
cc_105 N_Y_c_148_n N_VGND_c_191_n 0.0291015f $X=1.05 $Y=0.545 $X2=0 $Y2=0
cc_106 N_Y_c_148_n N_VGND_c_193_n 0.0211357f $X=1.05 $Y=0.545 $X2=0 $Y2=0
cc_107 N_Y_c_148_n A_268_67# 0.00418236f $X=1.05 $Y=0.545 $X2=-0.19 $Y2=-0.245
cc_108 Y A_268_67# 0.00148246f $X=0.635 $Y=0.84 $X2=-0.19 $Y2=-0.245
