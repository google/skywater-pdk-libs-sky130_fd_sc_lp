* File: sky130_fd_sc_lp__xnor2_4.pex.spice
* Created: Wed Sep  2 10:40:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XNOR2_4%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 65 66 67 68 71 72 74 77 78 83 86 88 89 105 120
c262 120 0 1.29663e-19 $X=7.885 $Y=1.51
c263 63 0 9.6647e-20 $X=7.885 $Y=0.745
c264 59 0 1.99483e-19 $X=7.85 $Y=2.465
c265 51 0 1.29745e-19 $X=7.42 $Y=2.465
c266 27 0 1.19078e-19 $X=3.645 $Y=2.465
r267 119 120 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.85 $Y=1.51
+ $X2=7.885 $Y2=1.51
r268 116 117 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.42 $Y=1.51
+ $X2=7.455 $Y2=1.51
r269 115 116 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=7.025 $Y=1.51
+ $X2=7.42 $Y2=1.51
r270 114 115 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.99 $Y=1.51
+ $X2=7.025 $Y2=1.51
r271 110 112 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.515 $Y=1.51
+ $X2=6.56 $Y2=1.51
r272 104 105 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.455 $Y=1.51
+ $X2=1.495 $Y2=1.51
r273 102 104 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.29 $Y=1.51
+ $X2=1.455 $Y2=1.51
r274 102 103 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.29
+ $Y=1.51 $X2=1.29 $Y2=1.51
r275 100 102 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.025 $Y=1.51
+ $X2=1.29 $Y2=1.51
r276 99 100 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=1.025 $Y2=1.51
r277 97 99 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=0.61 $Y=1.51
+ $X2=0.905 $Y2=1.51
r278 97 98 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.51 $X2=0.61 $Y2=1.51
r279 95 97 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.515 $Y=1.51
+ $X2=0.61 $Y2=1.51
r280 93 95 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.475 $Y=1.51
+ $X2=0.515 $Y2=1.51
r281 89 103 4.30969 $w=5.05e-07 $l=1.78746e-07 $layer=LI1_cond $X=1.285 $Y=1.665
+ $X2=1.427 $Y2=1.582
r282 88 89 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.582
+ $X2=1.2 $Y2=1.582
r283 88 98 3.78414 $w=3.33e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.582
+ $X2=0.61 $Y2=1.582
r284 86 87 8.01992 $w=2.51e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=1.85
+ $X2=3.665 $Y2=2.015
r285 84 119 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=7.705 $Y=1.51
+ $X2=7.85 $Y2=1.51
r286 84 117 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=7.705 $Y=1.51
+ $X2=7.455 $Y2=1.51
r287 83 84 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.705
+ $Y=1.51 $X2=7.705 $Y2=1.51
r288 81 114 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=6.685 $Y=1.51
+ $X2=6.99 $Y2=1.51
r289 81 112 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.685 $Y=1.51
+ $X2=6.56 $Y2=1.51
r290 80 83 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.685 $Y=1.51
+ $X2=7.705 $Y2=1.51
r291 80 81 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.685
+ $Y=1.51 $X2=6.685 $Y2=1.51
r292 78 80 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.475 $Y=1.51
+ $X2=6.685 $Y2=1.51
r293 76 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.39 $Y=1.595
+ $X2=6.475 $Y2=1.51
r294 76 77 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.39 $Y=1.595
+ $X2=6.39 $Y2=1.765
r295 75 86 3.01842 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.83 $Y=1.85
+ $X2=3.665 $Y2=1.85
r296 74 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.305 $Y=1.85
+ $X2=6.39 $Y2=1.765
r297 74 75 161.471 $w=1.68e-07 $l=2.475e-06 $layer=LI1_cond $X=6.305 $Y=1.85
+ $X2=3.83 $Y2=1.85
r298 72 109 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.51
+ $X2=3.665 $Y2=1.675
r299 72 108 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.51
+ $X2=3.665 $Y2=1.345
r300 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.665
+ $Y=1.51 $X2=3.665 $Y2=1.51
r301 69 86 3.87119 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=1.765
+ $X2=3.665 $Y2=1.85
r302 69 71 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.665 $Y=1.765
+ $X2=3.665 $Y2=1.51
r303 67 87 3.01842 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.5 $Y=2.015
+ $X2=3.665 $Y2=2.015
r304 67 68 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=3.5 $Y=2.015
+ $X2=1.57 $Y2=2.015
r305 66 68 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=1.427 $Y=1.93
+ $X2=1.57 $Y2=2.015
r306 65 103 3.2179 $w=2.85e-07 $l=1.68e-07 $layer=LI1_cond $X=1.427 $Y=1.75
+ $X2=1.427 $Y2=1.582
r307 65 66 7.27859 $w=2.83e-07 $l=1.8e-07 $layer=LI1_cond $X=1.427 $Y=1.75
+ $X2=1.427 $Y2=1.93
r308 61 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.885 $Y=1.345
+ $X2=7.885 $Y2=1.51
r309 61 63 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.885 $Y=1.345
+ $X2=7.885 $Y2=0.745
r310 57 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.85 $Y=1.675
+ $X2=7.85 $Y2=1.51
r311 57 59 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.85 $Y=1.675
+ $X2=7.85 $Y2=2.465
r312 53 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.455 $Y=1.345
+ $X2=7.455 $Y2=1.51
r313 53 55 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.455 $Y=1.345
+ $X2=7.455 $Y2=0.745
r314 49 116 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.42 $Y=1.675
+ $X2=7.42 $Y2=1.51
r315 49 51 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.42 $Y=1.675
+ $X2=7.42 $Y2=2.465
r316 45 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.345
+ $X2=7.025 $Y2=1.51
r317 45 47 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.025 $Y=1.345
+ $X2=7.025 $Y2=0.745
r318 41 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.99 $Y=1.675
+ $X2=6.99 $Y2=1.51
r319 41 43 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.99 $Y=1.675
+ $X2=6.99 $Y2=2.465
r320 37 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.56 $Y=1.675
+ $X2=6.56 $Y2=1.51
r321 37 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.56 $Y=1.675
+ $X2=6.56 $Y2=2.465
r322 33 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.515 $Y=1.345
+ $X2=6.515 $Y2=1.51
r323 33 35 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.515 $Y=1.345
+ $X2=6.515 $Y2=0.745
r324 31 108 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.685 $Y=0.745
+ $X2=3.685 $Y2=1.345
r325 27 109 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.645 $Y=2.465
+ $X2=3.645 $Y2=1.675
r326 21 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.675
+ $X2=1.495 $Y2=1.51
r327 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.495 $Y=1.675
+ $X2=1.495 $Y2=2.465
r328 17 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.345
+ $X2=1.455 $Y2=1.51
r329 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.455 $Y=1.345
+ $X2=1.455 $Y2=0.745
r330 13 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.025 $Y=1.345
+ $X2=1.025 $Y2=1.51
r331 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.025 $Y=1.345
+ $X2=1.025 $Y2=0.745
r332 9 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.905 $Y2=1.51
r333 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.905 $Y2=2.465
r334 5 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.345
+ $X2=0.515 $Y2=1.51
r335 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.515 $Y=1.345 $X2=0.515
+ $Y2=0.745
r336 1 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.675
+ $X2=0.475 $Y2=1.51
r337 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=1.675
+ $X2=0.475 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_4%B 3 7 11 15 19 23 27 31 33 35 38 40 42 45 47
+ 49 52 54 56 59 61 66 69 70 75 87 100 101
c214 75 0 3.09595e-19 $X=8.4 $Y=1.665
c215 66 0 1.19078e-19 $X=2.995 $Y=1.51
c216 27 0 7.53043e-20 $X=3.175 $Y=0.745
r217 101 102 4.52279 $w=3.73e-07 $l=3.5e-08 $layer=POLY_cond $X=9.57 $Y=1.535
+ $X2=9.605 $Y2=1.535
r218 100 104 36.3463 $w=3.23e-07 $l=1.025e-06 $layer=LI1_cond $X=9.425 $Y=1.587
+ $X2=8.4 $Y2=1.587
r219 99 101 18.7373 $w=3.73e-07 $l=1.45e-07 $layer=POLY_cond $X=9.425 $Y=1.535
+ $X2=9.57 $Y2=1.535
r220 99 100 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.425
+ $Y=1.51 $X2=9.425 $Y2=1.51
r221 97 99 32.3056 $w=3.73e-07 $l=2.5e-07 $layer=POLY_cond $X=9.175 $Y=1.535
+ $X2=9.425 $Y2=1.535
r222 96 97 4.52279 $w=3.73e-07 $l=3.5e-08 $layer=POLY_cond $X=9.14 $Y=1.535
+ $X2=9.175 $Y2=1.535
r223 95 96 51.0429 $w=3.73e-07 $l=3.95e-07 $layer=POLY_cond $X=8.745 $Y=1.535
+ $X2=9.14 $Y2=1.535
r224 94 95 4.52279 $w=3.73e-07 $l=3.5e-08 $layer=POLY_cond $X=8.71 $Y=1.535
+ $X2=8.745 $Y2=1.535
r225 92 94 39.4129 $w=3.73e-07 $l=3.05e-07 $layer=POLY_cond $X=8.405 $Y=1.535
+ $X2=8.71 $Y2=1.535
r226 92 104 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.405
+ $Y=1.51 $X2=8.405 $Y2=1.51
r227 90 92 11.63 $w=3.73e-07 $l=9e-08 $layer=POLY_cond $X=8.315 $Y=1.535
+ $X2=8.405 $Y2=1.535
r228 89 90 4.52279 $w=3.73e-07 $l=3.5e-08 $layer=POLY_cond $X=8.28 $Y=1.535
+ $X2=8.315 $Y2=1.535
r229 87 88 5.93231 $w=3.25e-07 $l=4e-08 $layer=POLY_cond $X=3.175 $Y=1.51
+ $X2=3.215 $Y2=1.51
r230 84 85 5.93231 $w=3.25e-07 $l=4e-08 $layer=POLY_cond $X=2.745 $Y=1.51
+ $X2=2.785 $Y2=1.51
r231 80 82 5.93231 $w=3.25e-07 $l=4e-08 $layer=POLY_cond $X=2.315 $Y=1.51
+ $X2=2.355 $Y2=1.51
r232 78 80 57.84 $w=3.25e-07 $l=3.9e-07 $layer=POLY_cond $X=1.925 $Y=1.51
+ $X2=2.315 $Y2=1.51
r233 77 78 5.93231 $w=3.25e-07 $l=4e-08 $layer=POLY_cond $X=1.885 $Y=1.51
+ $X2=1.925 $Y2=1.51
r234 75 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r235 73 80 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.315
+ $Y=1.51 $X2=2.315 $Y2=1.51
r236 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.665
r237 70 72 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=1.665
+ $X2=2.16 $Y2=1.665
r238 69 75 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r239 69 70 7.36385 $w=1.4e-07 $l=5.95e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=2.305 $Y2=1.665
r240 67 87 26.6954 $w=3.25e-07 $l=1.8e-07 $layer=POLY_cond $X=2.995 $Y=1.51
+ $X2=3.175 $Y2=1.51
r241 67 85 31.1446 $w=3.25e-07 $l=2.1e-07 $layer=POLY_cond $X=2.995 $Y=1.51
+ $X2=2.785 $Y2=1.51
r242 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.995
+ $Y=1.51 $X2=2.995 $Y2=1.51
r243 64 84 13.3477 $w=3.25e-07 $l=9e-08 $layer=POLY_cond $X=2.655 $Y=1.51
+ $X2=2.745 $Y2=1.51
r244 64 82 44.4923 $w=3.25e-07 $l=3e-07 $layer=POLY_cond $X=2.655 $Y=1.51
+ $X2=2.355 $Y2=1.51
r245 63 66 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.655 $Y=1.582
+ $X2=2.995 $Y2=1.582
r246 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.655
+ $Y=1.51 $X2=2.655 $Y2=1.51
r247 61 73 9.65663 $w=3.35e-07 $l=2.5e-07 $layer=LI1_cond $X=2.41 $Y=1.582
+ $X2=2.16 $Y2=1.582
r248 61 63 8.42831 $w=3.33e-07 $l=2.45e-07 $layer=LI1_cond $X=2.41 $Y=1.582
+ $X2=2.655 $Y2=1.582
r249 57 102 24.162 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.605 $Y=1.345
+ $X2=9.605 $Y2=1.535
r250 57 59 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=9.605 $Y=1.345
+ $X2=9.605 $Y2=0.745
r251 54 101 24.162 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.57 $Y=1.725
+ $X2=9.57 $Y2=1.535
r252 54 56 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.57 $Y=1.725
+ $X2=9.57 $Y2=2.465
r253 50 97 24.162 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.175 $Y=1.345
+ $X2=9.175 $Y2=1.535
r254 50 52 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=9.175 $Y=1.345
+ $X2=9.175 $Y2=0.745
r255 47 96 24.162 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.14 $Y=1.725
+ $X2=9.14 $Y2=1.535
r256 47 49 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.14 $Y=1.725
+ $X2=9.14 $Y2=2.465
r257 43 95 24.162 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.745 $Y=1.345
+ $X2=8.745 $Y2=1.535
r258 43 45 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.745 $Y=1.345
+ $X2=8.745 $Y2=0.745
r259 40 94 24.162 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.71 $Y=1.725
+ $X2=8.71 $Y2=1.535
r260 40 42 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.71 $Y=1.725
+ $X2=8.71 $Y2=2.465
r261 36 90 24.162 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.315 $Y=1.345
+ $X2=8.315 $Y2=1.535
r262 36 38 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.315 $Y=1.345
+ $X2=8.315 $Y2=0.745
r263 33 89 24.162 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.28 $Y=1.725
+ $X2=8.28 $Y2=1.535
r264 33 35 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.28 $Y=1.725
+ $X2=8.28 $Y2=2.465
r265 29 88 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.675
+ $X2=3.215 $Y2=1.51
r266 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.215 $Y=1.675
+ $X2=3.215 $Y2=2.465
r267 25 87 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.175 $Y=1.345
+ $X2=3.175 $Y2=1.51
r268 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.175 $Y=1.345
+ $X2=3.175 $Y2=0.745
r269 21 85 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.675
+ $X2=2.785 $Y2=1.51
r270 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.785 $Y=1.675
+ $X2=2.785 $Y2=2.465
r271 17 84 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.345
+ $X2=2.745 $Y2=1.51
r272 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.745 $Y=1.345
+ $X2=2.745 $Y2=0.745
r273 13 82 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.675
+ $X2=2.355 $Y2=1.51
r274 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.355 $Y=1.675
+ $X2=2.355 $Y2=2.465
r275 9 80 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=1.345
+ $X2=2.315 $Y2=1.51
r276 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.315 $Y=1.345
+ $X2=2.315 $Y2=0.745
r277 5 78 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.675
+ $X2=1.925 $Y2=1.51
r278 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.925 $Y=1.675
+ $X2=1.925 $Y2=2.465
r279 1 77 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.345
+ $X2=1.885 $Y2=1.51
r280 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.885 $Y=1.345 $X2=1.885
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_4%A_808_39# 1 2 3 4 5 6 21 25 29 33 37 39 40
+ 43 47 51 61 65 69 70 73 75 79 83 85 87 91 95 97 99 102 106 107 108 114 116 117
+ 119 129
c231 114 0 9.6647e-20 $X=8.53 $Y=1.16
c232 108 0 2.85944e-19 $X=7.67 $Y=1.86
c233 107 0 1.29663e-19 $X=6.135 $Y=1.335
c234 69 0 4.60864e-20 $X=7.54 $Y=1.86
c235 43 0 3.12942e-20 $X=5.485 $Y=0.745
r236 123 124 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=4.545 $Y=1.5
+ $X2=4.985 $Y2=1.5
r237 112 113 4.62437 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=2.005
+ $X2=7.67 $Y2=2.09
r238 111 112 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=7.67 $Y=1.96
+ $X2=7.67 $Y2=2.005
r239 108 111 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=7.67 $Y=1.86
+ $X2=7.67 $Y2=1.96
r240 105 129 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=5.905 $Y=1.5
+ $X2=6.13 $Y2=1.5
r241 105 127 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.905 $Y=1.5
+ $X2=5.7 $Y2=1.5
r242 104 107 11.072 $w=4.98e-07 $l=2.3e-07 $layer=LI1_cond $X=5.905 $Y=1.335
+ $X2=6.135 $Y2=1.335
r243 104 106 12.2681 $w=4.98e-07 $l=2.8e-07 $layer=LI1_cond $X=5.905 $Y=1.335
+ $X2=5.625 $Y2=1.335
r244 104 105 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.905
+ $Y=1.5 $X2=5.905 $Y2=1.5
r245 101 102 34.8352 $w=2.18e-07 $l=6.65e-07 $layer=LI1_cond $X=9.88 $Y=1.255
+ $X2=9.88 $Y2=1.92
r246 100 117 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=9.555 $Y=1.16
+ $X2=9.39 $Y2=1.16
r247 99 101 6.86407 $w=1.9e-07 $l=1.50167e-07 $layer=LI1_cond $X=9.77 $Y=1.16
+ $X2=9.88 $Y2=1.255
r248 99 100 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=9.77 $Y=1.16
+ $X2=9.555 $Y2=1.16
r249 98 119 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.45 $Y=2.005
+ $X2=9.355 $Y2=2.005
r250 97 102 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=9.77 $Y=2.005
+ $X2=9.88 $Y2=1.92
r251 97 98 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.77 $Y=2.005
+ $X2=9.45 $Y2=2.005
r252 93 119 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.355 $Y=2.09
+ $X2=9.355 $Y2=2.005
r253 93 95 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=9.355 $Y=2.09
+ $X2=9.355 $Y2=2.45
r254 89 117 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=9.39 $Y=1.065
+ $X2=9.39 $Y2=1.16
r255 89 91 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=9.39 $Y=1.065
+ $X2=9.39 $Y2=0.7
r256 88 114 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=1.16
+ $X2=8.53 $Y2=1.16
r257 87 117 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=9.225 $Y=1.16
+ $X2=9.39 $Y2=1.16
r258 87 88 30.9378 $w=1.88e-07 $l=5.3e-07 $layer=LI1_cond $X=9.225 $Y=1.16
+ $X2=8.695 $Y2=1.16
r259 86 116 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.59 $Y=2.005
+ $X2=8.495 $Y2=2.005
r260 85 119 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.26 $Y=2.005
+ $X2=9.355 $Y2=2.005
r261 85 86 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.26 $Y=2.005
+ $X2=8.59 $Y2=2.005
r262 81 116 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.495 $Y=2.09
+ $X2=8.495 $Y2=2.005
r263 81 83 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=8.495 $Y=2.09
+ $X2=8.495 $Y2=2.45
r264 77 114 0.718145 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=8.53 $Y=1.065
+ $X2=8.53 $Y2=1.16
r265 77 79 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=8.53 $Y=1.065
+ $X2=8.53 $Y2=0.7
r266 76 112 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.8 $Y=2.005
+ $X2=7.67 $Y2=2.005
r267 75 116 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.4 $Y=2.005
+ $X2=8.495 $Y2=2.005
r268 75 76 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.4 $Y=2.005 $X2=7.8
+ $Y2=2.005
r269 73 113 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.635 $Y=2.45
+ $X2=7.635 $Y2=2.09
r270 69 108 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.54 $Y=1.86
+ $X2=7.67 $Y2=1.86
r271 69 70 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.54 $Y=1.86
+ $X2=6.87 $Y2=1.86
r272 65 67 48.6587 $w=2.23e-07 $l=9.5e-07 $layer=LI1_cond $X=6.757 $Y=1.96
+ $X2=6.757 $Y2=2.91
r273 63 70 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=6.757 $Y=1.945
+ $X2=6.87 $Y2=1.86
r274 63 65 0.768295 $w=2.23e-07 $l=1.5e-08 $layer=LI1_cond $X=6.757 $Y=1.945
+ $X2=6.757 $Y2=1.96
r275 61 114 8.26956 $w=1.8e-07 $l=1.69926e-07 $layer=LI1_cond $X=8.365 $Y=1.17
+ $X2=8.53 $Y2=1.16
r276 61 107 145.487 $w=1.68e-07 $l=2.23e-06 $layer=LI1_cond $X=8.365 $Y=1.17
+ $X2=6.135 $Y2=1.17
r277 60 127 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=5.565 $Y=1.5
+ $X2=5.7 $Y2=1.5
r278 60 125 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.565 $Y=1.5
+ $X2=5.485 $Y2=1.5
r279 59 106 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.565 $Y=1.5
+ $X2=5.625 $Y2=1.5
r280 59 60 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.565
+ $Y=1.5 $X2=5.565 $Y2=1.5
r281 56 123 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.205 $Y=1.5
+ $X2=4.545 $Y2=1.5
r282 56 120 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.205 $Y=1.5
+ $X2=4.115 $Y2=1.5
r283 55 59 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.205 $Y=1.5
+ $X2=5.565 $Y2=1.5
r284 55 56 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.205
+ $Y=1.5 $X2=4.205 $Y2=1.5
r285 49 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.13 $Y=1.665
+ $X2=6.13 $Y2=1.5
r286 49 51 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=6.13 $Y=1.665
+ $X2=6.13 $Y2=2.465
r287 45 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.7 $Y=1.665
+ $X2=5.7 $Y2=1.5
r288 45 47 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.7 $Y=1.665 $X2=5.7
+ $Y2=2.465
r289 41 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.485 $Y=1.335
+ $X2=5.485 $Y2=1.5
r290 41 43 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.485 $Y=1.335
+ $X2=5.485 $Y2=0.745
r291 40 124 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.06 $Y=1.5
+ $X2=4.985 $Y2=1.5
r292 39 125 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.41 $Y=1.5
+ $X2=5.485 $Y2=1.5
r293 39 40 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=5.41 $Y=1.5
+ $X2=5.06 $Y2=1.5
r294 35 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.335
+ $X2=4.985 $Y2=1.5
r295 35 37 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.985 $Y=1.335
+ $X2=4.985 $Y2=0.745
r296 31 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.545 $Y=1.665
+ $X2=4.545 $Y2=1.5
r297 31 33 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.545 $Y=1.665
+ $X2=4.545 $Y2=2.465
r298 27 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.545 $Y=1.335
+ $X2=4.545 $Y2=1.5
r299 27 29 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.545 $Y=1.335
+ $X2=4.545 $Y2=0.745
r300 23 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.115 $Y=1.665
+ $X2=4.115 $Y2=1.5
r301 23 25 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.115 $Y=1.665
+ $X2=4.115 $Y2=2.465
r302 19 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.115 $Y=1.335
+ $X2=4.115 $Y2=1.5
r303 19 21 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.115 $Y=1.335
+ $X2=4.115 $Y2=0.745
r304 6 119 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=9.215
+ $Y=1.835 $X2=9.355 $Y2=2.005
r305 6 95 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=9.215
+ $Y=1.835 $X2=9.355 $Y2=2.45
r306 5 116 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=8.355
+ $Y=1.835 $X2=8.495 $Y2=2.005
r307 5 83 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=8.355
+ $Y=1.835 $X2=8.495 $Y2=2.45
r308 4 111 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.495
+ $Y=1.835 $X2=7.635 $Y2=1.96
r309 4 73 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=7.495
+ $Y=1.835 $X2=7.635 $Y2=2.45
r310 3 67 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.635
+ $Y=1.835 $X2=6.775 $Y2=2.91
r311 3 65 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=6.635
+ $Y=1.835 $X2=6.775 $Y2=1.96
r312 2 91 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=9.25
+ $Y=0.325 $X2=9.39 $Y2=0.7
r313 1 79 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=8.39
+ $Y=0.325 $X2=8.53 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 44 48 52
+ 56 58 60 63 64 66 67 68 69 70 72 84 95 100 109 116 125 128 132
r158 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r159 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r160 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r161 116 119 6.30269 $w=8.33e-07 $l=4.4e-07 $layer=LI1_cond $X=5.232 $Y=2.53
+ $X2=5.232 $Y2=2.97
r162 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r163 109 112 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=3.065
+ $X2=1.2 $Y2=3.33
r164 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r165 104 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r166 104 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r168 101 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=8.925 $Y2=3.33
r169 101 103 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=9.36 $Y2=3.33
r170 100 131 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=9.62 $Y=3.33
+ $X2=9.85 $Y2=3.33
r171 100 103 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.62 $Y=3.33
+ $X2=9.36 $Y2=3.33
r172 99 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r173 99 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r174 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r175 96 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.23 $Y=3.33
+ $X2=8.065 $Y2=3.33
r176 96 98 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.23 $Y=3.33
+ $X2=8.4 $Y2=3.33
r177 95 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.76 $Y=3.33
+ $X2=8.925 $Y2=3.33
r178 95 98 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.76 $Y=3.33
+ $X2=8.4 $Y2=3.33
r179 94 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r180 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r181 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r182 91 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r183 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r184 88 90 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.65 $Y=3.33 $X2=6
+ $Y2=3.33
r185 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r186 84 88 10.4966 $w=1.7e-07 $l=4.18e-07 $layer=LI1_cond $X=5.232 $Y=3.33
+ $X2=5.65 $Y2=3.33
r187 84 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r188 84 119 5.15675 $w=8.33e-07 $l=3.6e-07 $layer=LI1_cond $X=5.232 $Y=3.33
+ $X2=5.232 $Y2=2.97
r189 84 86 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.815 $Y=3.33
+ $X2=4.56 $Y2=3.33
r190 83 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r191 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r192 80 83 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r193 80 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r194 79 82 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r195 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r196 77 112 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.2 $Y2=3.33
r197 77 79 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.68 $Y2=3.33
r198 76 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r199 76 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r200 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r201 73 106 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r202 73 75 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r203 72 112 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.2 $Y2=3.33
r204 72 75 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.72 $Y2=3.33
r205 70 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r206 70 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r207 68 93 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.04 $Y=3.33 $X2=6.96
+ $Y2=3.33
r208 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.04 $Y=3.33
+ $X2=7.205 $Y2=3.33
r209 66 90 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.25 $Y=3.33 $X2=6
+ $Y2=3.33
r210 66 67 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.25 $Y=3.33
+ $X2=6.36 $Y2=3.33
r211 65 93 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=6.47 $Y=3.33
+ $X2=6.96 $Y2=3.33
r212 65 67 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.47 $Y=3.33
+ $X2=6.36 $Y2=3.33
r213 63 82 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=3.6 $Y2=3.33
r214 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=3.88 $Y2=3.33
r215 62 86 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.56 $Y2=3.33
r216 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=3.88 $Y2=3.33
r217 58 131 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=9.785 $Y=3.245
+ $X2=9.85 $Y2=3.33
r218 58 60 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=9.785 $Y=3.245
+ $X2=9.785 $Y2=2.365
r219 54 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.925 $Y=3.245
+ $X2=8.925 $Y2=3.33
r220 54 56 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=8.925 $Y=3.245
+ $X2=8.925 $Y2=2.365
r221 50 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.065 $Y=3.245
+ $X2=8.065 $Y2=3.33
r222 50 52 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=8.065 $Y=3.245
+ $X2=8.065 $Y2=2.365
r223 49 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=3.33
+ $X2=7.205 $Y2=3.33
r224 48 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.9 $Y=3.33
+ $X2=8.065 $Y2=3.33
r225 48 49 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.9 $Y=3.33
+ $X2=7.37 $Y2=3.33
r226 44 47 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=7.205 $Y=2.21
+ $X2=7.205 $Y2=2.97
r227 42 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.205 $Y=3.245
+ $X2=7.205 $Y2=3.33
r228 42 47 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.205 $Y=3.245
+ $X2=7.205 $Y2=2.97
r229 38 41 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=6.36 $Y=2.29
+ $X2=6.36 $Y2=2.97
r230 36 67 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.36 $Y=3.245
+ $X2=6.36 $Y2=3.33
r231 36 41 14.4055 $w=2.18e-07 $l=2.75e-07 $layer=LI1_cond $X=6.36 $Y=3.245
+ $X2=6.36 $Y2=2.97
r232 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=3.33
r233 32 34 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=2.745
r234 28 106 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r235 28 30 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.365
r236 9 60 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=9.645
+ $Y=1.835 $X2=9.785 $Y2=2.365
r237 8 56 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=8.785
+ $Y=1.835 $X2=8.925 $Y2=2.365
r238 7 52 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=7.925
+ $Y=1.835 $X2=8.065 $Y2=2.365
r239 6 47 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=7.065
+ $Y=1.835 $X2=7.205 $Y2=2.97
r240 6 44 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=7.065
+ $Y=1.835 $X2=7.205 $Y2=2.21
r241 5 41 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.835 $X2=6.345 $Y2=2.97
r242 5 38 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=1.835 $X2=6.345 $Y2=2.29
r243 4 119 300 $w=1.7e-07 $l=1.26729e-06 $layer=licon1_PDIFF $count=2 $X=4.62
+ $Y=1.835 $X2=4.9 $Y2=2.97
r244 4 116 300 $w=1.7e-07 $l=1.16164e-06 $layer=licon1_PDIFF $count=2 $X=4.62
+ $Y=1.835 $X2=5.485 $Y2=2.53
r245 3 34 600 $w=1.7e-07 $l=9.86762e-07 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.835 $X2=3.88 $Y2=2.745
r246 2 109 600 $w=1.7e-07 $l=1.33548e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.2 $Y2=3.065
r247 1 30 300 $w=1.7e-07 $l=5.89194e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_4%A_110_367# 1 2 3 4 15 19 24 27
r37 26 27 8.81087 $w=3.38e-07 $l=1.75e-07 $layer=LI1_cond $X=1.71 $Y=2.79
+ $X2=1.535 $Y2=2.79
r38 24 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.865 $Y=2.705
+ $X2=1.535 $Y2=2.705
r39 22 24 8.8114 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.69 $Y=2.785
+ $X2=0.865 $Y2=2.785
r40 17 19 29.15 $w=3.38e-07 $l=8.6e-07 $layer=LI1_cond $X=2.57 $Y=2.79 $X2=3.43
+ $Y2=2.79
r41 15 26 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=2.79
+ $X2=1.71 $Y2=2.79
r42 15 17 23.5573 $w=3.38e-07 $l=6.95e-07 $layer=LI1_cond $X=1.875 $Y=2.79
+ $X2=2.57 $Y2=2.79
r43 4 19 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=1.835 $X2=3.43 $Y2=2.795
r44 3 17 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.835 $X2=2.57 $Y2=2.795
r45 2 26 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.835 $X2=1.71 $Y2=2.795
r46 1 22 600 $w=1.7e-07 $l=1.0176e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_4%Y 1 2 3 4 5 6 20 21 22 23 24 26 27 28 35 37
+ 39 43 45 47 49 52 53 64 71
r143 71 72 1.27814 $w=4.78e-07 $l=4.5e-08 $layer=LI1_cond $X=4.405 $Y=2.405
+ $X2=4.405 $Y2=2.45
r144 67 68 3.48856 $w=4.78e-07 $l=1.4e-07 $layer=LI1_cond $X=4.405 $Y=2.22
+ $X2=4.405 $Y2=2.36
r145 64 67 0.747549 $w=4.78e-07 $l=3e-08 $layer=LI1_cond $X=4.405 $Y=2.19
+ $X2=4.405 $Y2=2.22
r146 53 60 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.43 $Y=2.775
+ $X2=4.43 $Y2=2.56
r147 52 71 0.498366 $w=4.78e-07 $l=2e-08 $layer=LI1_cond $X=4.405 $Y=2.385
+ $X2=4.405 $Y2=2.405
r148 52 68 0.622958 $w=4.78e-07 $l=2.5e-08 $layer=LI1_cond $X=4.405 $Y=2.385
+ $X2=4.405 $Y2=2.36
r149 52 60 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=4.43 $Y=2.47 $X2=4.43
+ $Y2=2.56
r150 52 72 0.53602 $w=4.28e-07 $l=2e-08 $layer=LI1_cond $X=4.43 $Y=2.47 $X2=4.43
+ $Y2=2.45
r151 45 51 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=2.275
+ $X2=5.95 $Y2=2.19
r152 45 47 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=5.95 $Y=2.275
+ $X2=5.95 $Y2=2.55
r153 41 43 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=5.27 $Y=1.075
+ $X2=5.27 $Y2=0.68
r154 40 64 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=4.645 $Y=2.19
+ $X2=4.405 $Y2=2.19
r155 39 51 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.82 $Y=2.19
+ $X2=5.95 $Y2=2.19
r156 39 40 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=5.82 $Y=2.19
+ $X2=4.645 $Y2=2.19
r157 38 49 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.435 $Y=1.16
+ $X2=4.335 $Y2=1.16
r158 37 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.105 $Y=1.16
+ $X2=5.27 $Y2=1.075
r159 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.105 $Y=1.16
+ $X2=4.435 $Y2=1.16
r160 33 49 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.335 $Y=1.075
+ $X2=4.335 $Y2=1.16
r161 33 35 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=4.335 $Y=1.075
+ $X2=4.335 $Y2=0.77
r162 30 32 52.9899 $w=1.78e-07 $l=8.6e-07 $layer=LI1_cond $X=2.14 $Y=2.36 $X2=3
+ $Y2=2.36
r163 28 30 63.1566 $w=1.78e-07 $l=1.025e-06 $layer=LI1_cond $X=1.115 $Y=2.36
+ $X2=2.14 $Y2=2.36
r164 27 68 6.54597 $w=1.8e-07 $l=2.4e-07 $layer=LI1_cond $X=4.165 $Y=2.36
+ $X2=4.405 $Y2=2.36
r165 27 32 71.7828 $w=1.78e-07 $l=1.165e-06 $layer=LI1_cond $X=4.165 $Y=2.36
+ $X2=3 $Y2=2.36
r166 26 28 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.03 $Y=2.27
+ $X2=1.115 $Y2=2.36
r167 25 26 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.03 $Y=2.09
+ $X2=1.03 $Y2=2.27
r168 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.945 $Y=2.005
+ $X2=1.03 $Y2=2.09
r169 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.945 $Y=2.005
+ $X2=0.275 $Y2=2.005
r170 21 49 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.235 $Y=1.16
+ $X2=4.335 $Y2=1.16
r171 21 22 258.353 $w=1.68e-07 $l=3.96e-06 $layer=LI1_cond $X=4.235 $Y=1.16
+ $X2=0.275 $Y2=1.16
r172 20 24 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.185 $Y=1.92
+ $X2=0.275 $Y2=2.005
r173 19 22 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.185 $Y=1.245
+ $X2=0.275 $Y2=1.16
r174 19 20 41.5909 $w=1.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.185 $Y=1.245
+ $X2=0.185 $Y2=1.92
r175 6 51 600 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=5.775
+ $Y=1.835 $X2=5.915 $Y2=2.19
r176 6 47 300 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_PDIFF $count=2 $X=5.775
+ $Y=1.835 $X2=5.915 $Y2=2.55
r177 5 67 600 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=4.19
+ $Y=1.835 $X2=4.33 $Y2=2.22
r178 5 60 300 $w=1.7e-07 $l=7.91912e-07 $layer=licon1_PDIFF $count=2 $X=4.19
+ $Y=1.835 $X2=4.33 $Y2=2.56
r179 4 32 600 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.835 $X2=3 $Y2=2.365
r180 3 30 600 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.835 $X2=2.14 $Y2=2.365
r181 2 43 91 $w=1.7e-07 $l=4.47856e-07 $layer=licon1_NDIFF $count=2 $X=5.06
+ $Y=0.325 $X2=5.27 $Y2=0.68
r182 1 35 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=4.19
+ $Y=0.325 $X2=4.33 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_4%A_31_65# 1 2 3 4 5 6 7 24 26 27 30 32 36 38
+ 42 44 49 50 51 54 56 60 63 65 67 68
c120 68 0 3.12942e-20 $X=4.77 $Y=0.345
c121 51 0 7.53043e-20 $X=4.065 $Y=0.345
r122 58 60 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.77 $Y=0.425
+ $X2=5.77 $Y2=0.47
r123 57 68 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.935 $Y=0.34
+ $X2=4.77 $Y2=0.345
r124 56 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.605 $Y=0.34
+ $X2=5.77 $Y2=0.425
r125 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.605 $Y=0.34
+ $X2=4.935 $Y2=0.34
r126 52 68 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.77 $Y=0.435
+ $X2=4.77 $Y2=0.345
r127 52 54 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.77 $Y=0.435
+ $X2=4.77 $Y2=0.45
r128 50 68 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=0.345
+ $X2=4.77 $Y2=0.345
r129 50 51 33.2727 $w=1.78e-07 $l=5.4e-07 $layer=LI1_cond $X=4.605 $Y=0.345
+ $X2=4.065 $Y2=0.345
r130 47 49 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.9 $Y=0.735
+ $X2=3.9 $Y2=0.45
r131 46 51 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.9 $Y=0.435
+ $X2=4.065 $Y2=0.345
r132 46 49 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.9 $Y=0.435
+ $X2=3.9 $Y2=0.45
r133 45 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.055 $Y=0.82
+ $X2=2.96 $Y2=0.82
r134 44 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.735 $Y=0.82
+ $X2=3.9 $Y2=0.735
r135 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.735 $Y=0.82
+ $X2=3.055 $Y2=0.82
r136 40 67 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.96 $Y=0.735
+ $X2=2.96 $Y2=0.82
r137 40 42 16.6364 $w=1.88e-07 $l=2.85e-07 $layer=LI1_cond $X=2.96 $Y=0.735
+ $X2=2.96 $Y2=0.45
r138 39 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.195 $Y=0.82
+ $X2=2.1 $Y2=0.82
r139 38 67 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.865 $Y=0.82
+ $X2=2.96 $Y2=0.82
r140 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.865 $Y=0.82
+ $X2=2.195 $Y2=0.82
r141 34 65 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=0.735
+ $X2=2.1 $Y2=0.82
r142 34 36 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=2.1 $Y=0.735
+ $X2=2.1 $Y2=0.48
r143 33 63 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.335 $Y=0.82
+ $X2=1.245 $Y2=0.82
r144 32 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.005 $Y=0.82
+ $X2=2.1 $Y2=0.82
r145 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=0.82
+ $X2=1.335 $Y2=0.82
r146 28 63 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.735
+ $X2=1.245 $Y2=0.82
r147 28 30 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=1.245 $Y=0.735
+ $X2=1.245 $Y2=0.48
r148 26 63 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.155 $Y=0.82
+ $X2=1.245 $Y2=0.82
r149 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.155 $Y=0.82
+ $X2=0.465 $Y2=0.82
r150 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.3 $Y=0.735
+ $X2=0.465 $Y2=0.82
r151 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.3 $Y=0.735
+ $X2=0.3 $Y2=0.46
r152 7 60 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.56
+ $Y=0.325 $X2=5.77 $Y2=0.47
r153 6 54 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=4.62
+ $Y=0.325 $X2=4.77 $Y2=0.45
r154 5 49 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.76
+ $Y=0.325 $X2=3.9 $Y2=0.45
r155 4 67 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.325 $X2=2.96 $Y2=0.82
r156 4 42 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.325 $X2=2.96 $Y2=0.45
r157 3 65 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.325 $X2=2.1 $Y2=0.82
r158 3 36 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.325 $X2=2.1 $Y2=0.48
r159 2 63 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.325 $X2=1.24 $Y2=0.82
r160 2 30 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.325 $X2=1.24 $Y2=0.48
r161 1 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.325 $X2=0.3 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_4%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 50 51 53 54 55 57 62 87 88 91 94
r157 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r158 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r159 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r160 85 88 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r161 84 87 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r162 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r163 82 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r164 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r165 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r166 78 79 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r167 75 78 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6.48
+ $Y2=0
r168 75 76 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r169 73 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r170 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r171 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r172 70 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r173 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r174 67 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.67
+ $Y2=0
r175 67 69 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.835 $Y=0
+ $X2=2.16 $Y2=0
r176 66 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r177 66 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r178 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r179 63 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.8
+ $Y2=0
r180 63 65 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.2
+ $Y2=0
r181 62 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=0 $X2=1.67
+ $Y2=0
r182 62 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.505 $Y=0 $X2=1.2
+ $Y2=0
r183 60 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r184 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r185 57 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.8
+ $Y2=0
r186 57 59 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=0
+ $X2=0.24 $Y2=0
r187 55 79 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r188 55 76 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=3.6
+ $Y2=0
r189 53 81 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.505 $Y=0 $X2=7.44
+ $Y2=0
r190 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.505 $Y=0 $X2=7.67
+ $Y2=0
r191 52 84 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.835 $Y=0 $X2=7.92
+ $Y2=0
r192 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.835 $Y=0 $X2=7.67
+ $Y2=0
r193 50 78 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.635 $Y=0
+ $X2=6.48 $Y2=0
r194 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.635 $Y=0 $X2=6.8
+ $Y2=0
r195 49 81 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=6.965 $Y=0
+ $X2=7.44 $Y2=0
r196 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.965 $Y=0 $X2=6.8
+ $Y2=0
r197 47 72 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.225 $Y=0
+ $X2=3.12 $Y2=0
r198 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.39
+ $Y2=0
r199 46 75 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.6
+ $Y2=0
r200 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.39
+ $Y2=0
r201 44 69 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.365 $Y=0
+ $X2=2.16 $Y2=0
r202 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.53
+ $Y2=0
r203 43 72 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.695 $Y=0
+ $X2=3.12 $Y2=0
r204 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.53
+ $Y2=0
r205 39 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=0.085
+ $X2=7.67 $Y2=0
r206 39 41 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.67 $Y=0.085
+ $X2=7.67 $Y2=0.45
r207 35 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.8 $Y=0.085 $X2=6.8
+ $Y2=0
r208 35 37 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=6.8 $Y=0.085
+ $X2=6.8 $Y2=0.45
r209 31 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.39 $Y2=0
r210 31 33 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.39 $Y=0.085
+ $X2=3.39 $Y2=0.45
r211 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0
r212 27 29 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.53 $Y=0.085
+ $X2=2.53 $Y2=0.45
r213 23 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r214 23 25 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.45
r215 19 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0
r216 19 21 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.8 $Y=0.085
+ $X2=0.8 $Y2=0.45
r217 6 41 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=7.53
+ $Y=0.325 $X2=7.67 $Y2=0.45
r218 5 37 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=6.59
+ $Y=0.325 $X2=6.8 $Y2=0.45
r219 4 33 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.325 $X2=3.39 $Y2=0.45
r220 3 29 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.325 $X2=2.53 $Y2=0.45
r221 2 25 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.325 $X2=1.67 $Y2=0.45
r222 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.325 $X2=0.8 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR2_4%A_1235_65# 1 2 3 4 5 18 20 21 24 26 29 30 31
+ 34 36 40 43 46
r72 38 40 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=9.855 $Y=0.425
+ $X2=9.855 $Y2=0.73
r73 37 46 5.52892 $w=1.75e-07 $l=9.74679e-08 $layer=LI1_cond $X=9.055 $Y=0.34
+ $X2=8.96 $Y2=0.345
r74 36 38 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.725 $Y=0.34
+ $X2=9.855 $Y2=0.425
r75 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.725 $Y=0.34
+ $X2=9.055 $Y2=0.34
r76 32 46 1.04816 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=8.96 $Y=0.435 $X2=8.96
+ $Y2=0.345
r77 32 34 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=8.96 $Y=0.435
+ $X2=8.96 $Y2=0.73
r78 30 46 5.52892 $w=1.75e-07 $l=9.5e-08 $layer=LI1_cond $X=8.865 $Y=0.345
+ $X2=8.96 $Y2=0.345
r79 30 31 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=8.865 $Y=0.345
+ $X2=8.195 $Y2=0.345
r80 29 45 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.1 $Y=0.745 $X2=8.1
+ $Y2=0.83
r81 28 31 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=8.1 $Y=0.435
+ $X2=8.195 $Y2=0.345
r82 28 29 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=8.1 $Y=0.435 $X2=8.1
+ $Y2=0.745
r83 27 43 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.335 $Y=0.83 $X2=7.235
+ $Y2=0.83
r84 26 45 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.005 $Y=0.83 $X2=8.1
+ $Y2=0.83
r85 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.005 $Y=0.83
+ $X2=7.335 $Y2=0.83
r86 22 43 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.235 $Y=0.745
+ $X2=7.235 $Y2=0.83
r87 22 24 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=7.235 $Y=0.745
+ $X2=7.235 $Y2=0.45
r88 20 43 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.135 $Y=0.83 $X2=7.235
+ $Y2=0.83
r89 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.135 $Y=0.83
+ $X2=6.465 $Y2=0.83
r90 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.3 $Y=0.745
+ $X2=6.465 $Y2=0.83
r91 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.3 $Y=0.745
+ $X2=6.3 $Y2=0.47
r92 5 40 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=9.68
+ $Y=0.325 $X2=9.82 $Y2=0.73
r93 4 34 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=8.82
+ $Y=0.325 $X2=8.96 $Y2=0.73
r94 3 45 182 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_NDIFF $count=1 $X=7.96
+ $Y=0.325 $X2=8.1 $Y2=0.75
r95 2 43 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=7.1
+ $Y=0.325 $X2=7.24 $Y2=0.83
r96 2 24 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=7.1
+ $Y=0.325 $X2=7.24 $Y2=0.45
r97 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.175
+ $Y=0.325 $X2=6.3 $Y2=0.47
.ends

