* File: sky130_fd_sc_lp__dfstp_4.pex.spice
* Created: Wed Sep  2 09:44:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFSTP_4%CLK 3 5 8 10 11 12 13 14 15 22 24
r39 22 24 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.602 $Y=1.19
+ $X2=0.602 $Y2=1.025
r40 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.625
+ $Y=1.19 $X2=0.625 $Y2=1.19
r41 14 15 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.672 $Y=1.665
+ $X2=0.672 $Y2=2.035
r42 13 14 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.672 $Y=1.295
+ $X2=0.672 $Y2=1.665
r43 13 23 4.24584 $w=2.83e-07 $l=1.05e-07 $layer=LI1_cond $X=0.672 $Y=1.295
+ $X2=0.672 $Y2=1.19
r44 12 23 10.7157 $w=2.83e-07 $l=2.65e-07 $layer=LI1_cond $X=0.672 $Y=0.925
+ $X2=0.672 $Y2=1.19
r45 11 12 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.672 $Y=0.555
+ $X2=0.672 $Y2=0.925
r46 8 10 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.645 $Y=2.645
+ $X2=0.645 $Y2=1.695
r47 5 10 40.5548 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.602 $Y=1.508
+ $X2=0.602 $Y2=1.695
r48 4 22 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.602 $Y=1.212
+ $X2=0.602 $Y2=1.19
r49 4 5 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.602 $Y=1.212
+ $X2=0.602 $Y2=1.508
r50 3 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.49 $Y=0.705
+ $X2=0.49 $Y2=1.025
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%D 3 4 5 7 9 10 12 13 16 18
c52 18 0 1.90265e-19 $X=1.865 $Y=1.915
c53 16 0 1.87691e-19 $X=1.865 $Y=2.08
c54 13 0 1.95278e-19 $X=2.16 $Y=2.035
r55 16 19 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.865 $Y=2.08
+ $X2=1.865 $Y2=2.13
r56 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=2.08
+ $X2=1.865 $Y2=1.915
r57 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=2.08 $X2=1.865 $Y2=2.08
r58 13 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.16 $Y=2.08
+ $X2=1.865 $Y2=2.08
r59 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.515 $Y=2.205
+ $X2=2.515 $Y2=2.525
r60 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.305 $Y=1.125
+ $X2=2.305 $Y2=0.805
r61 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=2.13
+ $X2=1.865 $Y2=2.13
r62 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.44 $Y=2.13
+ $X2=2.515 $Y2=2.205
r63 5 6 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.44 $Y=2.13 $X2=2.03
+ $Y2=2.13
r64 3 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.23 $Y=1.2
+ $X2=2.305 $Y2=1.125
r65 3 4 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.23 $Y=1.2 $X2=2.03
+ $Y2=1.2
r66 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.955 $Y=1.275
+ $X2=2.03 $Y2=1.2
r67 1 18 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.955 $Y=1.275
+ $X2=1.955 $Y2=1.915
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_230_465# 1 2 7 11 15 19 23 26 29 32 38 42
+ 46 47 48 51 54 57 63 64
c173 64 0 9.13638e-20 $X=6.16 $Y=1.51
c174 63 0 7.15321e-20 $X=5.845 $Y=1.51
c175 57 0 5.22509e-20 $X=2.435 $Y=1.56
c176 48 0 1.95278e-19 $X=1.825 $Y=1.295
c177 47 0 1.41563e-20 $X=5.375 $Y=1.295
c178 38 0 8.79279e-20 $X=1.515 $Y=2.805
r179 62 64 63.5272 $w=2.39e-07 $l=3.15e-07 $layer=POLY_cond $X=5.845 $Y=1.51
+ $X2=6.16 $Y2=1.51
r180 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.845
+ $Y=1.51 $X2=5.845 $Y2=1.51
r181 55 63 8.41672 $w=4.43e-07 $l=3.25e-07 $layer=LI1_cond $X=5.52 $Y=1.372
+ $X2=5.845 $Y2=1.372
r182 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r183 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=1.295
+ $X2=1.68 $Y2=1.295
r184 48 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.825 $Y=1.295
+ $X2=1.68 $Y2=1.295
r185 47 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=5.52 $Y2=1.295
r186 47 48 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=1.825 $Y2=1.295
r187 45 51 5.68738 $w=3.83e-07 $l=1.9e-07 $layer=LI1_cond $X=1.622 $Y=1.485
+ $X2=1.622 $Y2=1.295
r188 45 46 4.89178 $w=2.77e-07 $l=1.3e-07 $layer=LI1_cond $X=1.622 $Y=1.485
+ $X2=1.622 $Y2=1.615
r189 44 51 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=1.622 $Y=0.935
+ $X2=1.622 $Y2=1.295
r190 42 44 6.23421 $w=4.38e-07 $l=2.3e-07 $layer=LI1_cond $X=1.595 $Y=0.705
+ $X2=1.595 $Y2=0.935
r191 36 38 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.29 $Y=2.805
+ $X2=1.515 $Y2=2.805
r192 33 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.435 $Y=1.65
+ $X2=2.435 $Y2=1.56
r193 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=1.65 $X2=2.435 $Y2=1.65
r194 30 46 1.57815 $w=2.6e-07 $l=1.93e-07 $layer=LI1_cond $X=1.815 $Y=1.615
+ $X2=1.622 $Y2=1.615
r195 30 32 27.4813 $w=2.58e-07 $l=6.2e-07 $layer=LI1_cond $X=1.815 $Y=1.615
+ $X2=2.435 $Y2=1.615
r196 29 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=2.64
+ $X2=1.515 $Y2=2.805
r197 28 46 4.89178 $w=2.77e-07 $l=1.75528e-07 $layer=LI1_cond $X=1.515 $Y=1.745
+ $X2=1.622 $Y2=1.615
r198 28 29 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.515 $Y=1.745
+ $X2=1.515 $Y2=2.64
r199 25 26 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.945 $Y=1.56
+ $X2=3.165 $Y2=1.56
r200 21 64 37.3096 $w=2.39e-07 $l=1.85e-07 $layer=POLY_cond $X=6.345 $Y=1.51
+ $X2=6.16 $Y2=1.51
r201 21 23 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=6.345 $Y=1.525
+ $X2=6.345 $Y2=2.245
r202 17 64 13.6804 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.345
+ $X2=6.16 $Y2=1.51
r203 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.16 $Y=1.345
+ $X2=6.16 $Y2=0.555
r204 13 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=1.485
+ $X2=3.165 $Y2=1.56
r205 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.165 $Y=1.485
+ $X2=3.165 $Y2=0.805
r206 9 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.945 $Y=1.635
+ $X2=2.945 $Y2=1.56
r207 9 11 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2.945 $Y=1.635
+ $X2=2.945 $Y2=2.525
r208 8 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.56
+ $X2=2.435 $Y2=1.56
r209 7 25 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.87 $Y=1.56
+ $X2=2.945 $Y2=1.56
r210 7 8 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.87 $Y=1.56 $X2=2.6
+ $Y2=1.56
r211 2 36 600 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=2.325 $X2=1.29 $Y2=2.805
r212 1 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.36
+ $Y=0.495 $X2=1.5 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_690_93# 1 2 7 9 14 16 19 21 25 29 36 37 42
+ 45
c84 45 0 1.2803e-19 $X=3.825 $Y=1.825
c85 25 0 1.67044e-19 $X=4.28 $Y=0.45
c86 21 0 9.72951e-20 $X=4.115 $Y=1.07
r87 36 37 9.63527 $w=3.53e-07 $l=2e-07 $layer=LI1_cond $X=4.482 $Y=2.525
+ $X2=4.482 $Y2=2.325
r88 33 42 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.645 $Y=1.29
+ $X2=3.735 $Y2=1.29
r89 33 39 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=3.645 $Y=1.29
+ $X2=3.525 $Y2=1.29
r90 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.645
+ $Y=1.29 $X2=3.645 $Y2=1.29
r91 29 32 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.645 $Y=1.07
+ $X2=3.645 $Y2=1.29
r92 27 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.39 $Y=2.155
+ $X2=4.39 $Y2=2.325
r93 23 25 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=4.28 $Y=0.985
+ $X2=4.28 $Y2=0.45
r94 22 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=1.07
+ $X2=3.645 $Y2=1.07
r95 21 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.115 $Y=1.07
+ $X2=4.28 $Y2=0.985
r96 21 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.115 $Y=1.07
+ $X2=3.81 $Y2=1.07
r97 19 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.99
+ $X2=3.825 $Y2=2.155
r98 19 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.99
+ $X2=3.825 $Y2=1.825
r99 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.99 $X2=3.825 $Y2=1.99
r100 16 27 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.305 $Y=2.025
+ $X2=4.39 $Y2=2.155
r101 16 18 21.2759 $w=2.58e-07 $l=4.8e-07 $layer=LI1_cond $X=4.305 $Y=2.025
+ $X2=3.825 $Y2=2.025
r102 14 46 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.735 $Y=2.525
+ $X2=3.735 $Y2=2.155
r103 10 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.735 $Y=1.455
+ $X2=3.735 $Y2=1.29
r104 10 45 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.735 $Y=1.455
+ $X2=3.735 $Y2=1.825
r105 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=1.125
+ $X2=3.525 $Y2=1.29
r106 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.525 $Y=1.125
+ $X2=3.525 $Y2=0.805
r107 2 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.355
+ $Y=2.315 $X2=4.495 $Y2=2.525
r108 1 25 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.235 $X2=4.28 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%SET_B 3 7 8 10 11 12 13 15 19 20 23 27 29 30
+ 31 32 33 34 35 45
c116 35 0 2.63443e-19 $X=8.4 $Y=1.665
c117 30 0 4.32671e-20 $X=6.35 $Y=1.63
c118 20 0 2.78495e-19 $X=4.945 $Y=0.94
c119 19 0 7.49068e-20 $X=4.945 $Y=0.94
r120 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.905
+ $Y=1.41 $X2=7.905 $Y2=1.41
r121 34 35 11.2572 $w=5.08e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=1.58
+ $X2=8.4 $Y2=1.58
r122 34 50 0.351788 $w=5.08e-07 $l=1.5e-08 $layer=LI1_cond $X=7.92 $Y=1.58
+ $X2=7.905 $Y2=1.58
r123 33 50 10.9054 $w=5.08e-07 $l=4.65e-07 $layer=LI1_cond $X=7.44 $Y=1.58
+ $X2=7.905 $Y2=1.58
r124 32 33 11.2572 $w=5.08e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.58
+ $X2=7.44 $Y2=1.58
r125 31 32 11.2572 $w=5.08e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.58
+ $X2=6.96 $Y2=1.58
r126 30 31 3.04883 $w=5.08e-07 $l=1.3e-07 $layer=LI1_cond $X=6.35 $Y=1.58
+ $X2=6.48 $Y2=1.58
r127 29 30 9.69611 $w=5.08e-07 $l=1.7e-07 $layer=LI1_cond $X=6.18 $Y=1.63
+ $X2=6.35 $Y2=1.63
r128 27 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.73 $Y=1.99
+ $X2=4.73 $Y2=2.155
r129 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.73
+ $Y=1.99 $X2=4.73 $Y2=1.99
r130 23 26 5.42222 $w=3.15e-07 $l=3.09175e-07 $layer=LI1_cond $X=4.977 $Y=1.85
+ $X2=4.73 $Y2=1.99
r131 23 29 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=5.11 $Y=1.85
+ $X2=6.18 $Y2=1.85
r132 20 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.945 $Y=0.94
+ $X2=4.945 $Y2=0.775
r133 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.945
+ $Y=0.94 $X2=4.945 $Y2=0.94
r134 17 23 3.50625 $w=4.65e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.877 $Y=1.765
+ $X2=4.977 $Y2=1.85
r135 17 19 21.2207 $w=4.63e-07 $l=8.25e-07 $layer=LI1_cond $X=4.877 $Y=1.765
+ $X2=4.877 $Y2=0.94
r136 13 49 72.9565 $w=5.53e-07 $l=6.29623e-07 $layer=POLY_cond $X=8.375 $Y=1.915
+ $X2=8.095 $Y2=1.41
r137 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.375 $Y=1.915
+ $X2=8.375 $Y2=2.495
r138 11 49 30.5063 $w=5.53e-07 $l=5.00275e-07 $layer=POLY_cond $X=7.74 $Y=1.06
+ $X2=8.095 $Y2=1.41
r139 11 12 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.74 $Y=1.06
+ $X2=7.5 $Y2=1.06
r140 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.425 $Y=0.985
+ $X2=7.5 $Y2=1.06
r141 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.425 $Y=0.985
+ $X2=7.425 $Y2=0.665
r142 7 45 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.855 $Y=0.445
+ $X2=4.855 $Y2=0.775
r143 3 43 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.71 $Y=2.525
+ $X2=4.71 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_562_119# 1 2 9 13 15 18 21 23 24 25 27 28
+ 30 33 38 41 42 44 46 55
c136 46 0 1.2803e-19 $X=4.3 $Y=1.42
c137 44 0 1.22064e-19 $X=3.215 $Y=1.64
c138 38 0 1.31402e-19 $X=3.215 $Y=0.75
c139 21 0 1.62847e-19 $X=5.395 $Y=2.315
r140 54 55 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.495 $Y=1.42
+ $X2=4.57 $Y2=1.42
r141 47 54 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.3 $Y=1.42
+ $X2=4.495 $Y2=1.42
r142 47 51 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.3 $Y=1.42 $X2=4.28
+ $Y2=1.42
r143 46 49 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.3 $Y=1.42 $X2=4.3
+ $Y2=1.64
r144 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.3
+ $Y=1.42 $X2=4.3 $Y2=1.42
r145 41 42 11.479 $w=2.63e-07 $l=2.3e-07 $layer=LI1_cond $X=3.167 $Y=2.525
+ $X2=3.167 $Y2=2.295
r146 36 38 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.95 $Y=0.75
+ $X2=3.215 $Y2=0.75
r147 34 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=1.64
+ $X2=3.215 $Y2=1.64
r148 33 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=1.64
+ $X2=4.3 $Y2=1.64
r149 33 34 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.135 $Y=1.64
+ $X2=3.3 $Y2=1.64
r150 31 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=1.725
+ $X2=3.215 $Y2=1.64
r151 31 42 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.215 $Y=1.725
+ $X2=3.215 $Y2=2.295
r152 30 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=1.555
+ $X2=3.215 $Y2=1.64
r153 29 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=0.915
+ $X2=3.215 $Y2=0.75
r154 29 30 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.215 $Y=0.915
+ $X2=3.215 $Y2=1.555
r155 25 27 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.8 $Y=0.985
+ $X2=5.8 $Y2=0.555
r156 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.725 $Y=1.06
+ $X2=5.8 $Y2=0.985
r157 23 24 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.725 $Y=1.06
+ $X2=5.47 $Y2=1.06
r158 19 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.395 $Y=1.585
+ $X2=5.395 $Y2=1.51
r159 19 21 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=5.395 $Y=1.585
+ $X2=5.395 $Y2=2.315
r160 18 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.395 $Y=1.435
+ $X2=5.395 $Y2=1.51
r161 17 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.395 $Y=1.135
+ $X2=5.47 $Y2=1.06
r162 17 18 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=5.395 $Y=1.135
+ $X2=5.395 $Y2=1.435
r163 15 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.32 $Y=1.51
+ $X2=5.395 $Y2=1.51
r164 15 55 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.32 $Y=1.51
+ $X2=4.57 $Y2=1.51
r165 11 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.495 $Y=1.255
+ $X2=4.495 $Y2=1.42
r166 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.495 $Y=1.255
+ $X2=4.495 $Y2=0.445
r167 7 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.28 $Y=1.585
+ $X2=4.28 $Y2=1.42
r168 7 9 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.28 $Y=1.585 $X2=4.28
+ $Y2=2.525
r169 2 41 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=2.315 $X2=3.16 $Y2=2.525
r170 1 36 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.595 $X2=2.95 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_30_99# 1 2 8 12 13 14 18 19 20 23 27 29 33
+ 38 39 40 43 47 51 53 57 58 60
c138 57 0 1.90265e-19 $X=1.165 $Y=1.66
c139 43 0 1.19092e-19 $X=6.87 $Y=1.85
c140 38 0 4.32671e-20 $X=6.87 $Y=2.455
c141 33 0 7.15321e-20 $X=6.705 $Y=0.665
c142 23 0 1.75661e-19 $X=2.735 $Y=0.805
c143 12 0 8.79279e-20 $X=1.075 $Y=2.645
r144 58 62 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.66
+ $X2=1.18 $Y2=1.495
r145 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.165
+ $Y=1.66 $X2=1.165 $Y2=1.66
r146 55 57 28.3678 $w=2.58e-07 $l=6.4e-07 $layer=LI1_cond $X=1.13 $Y=2.3
+ $X2=1.13 $Y2=1.66
r147 54 60 3.08518 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.525 $Y=2.385
+ $X2=0.347 $Y2=2.385
r148 53 55 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1 $Y=2.385
+ $X2=1.13 $Y2=2.3
r149 53 54 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1 $Y=2.385
+ $X2=0.525 $Y2=2.385
r150 51 60 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=0.347 $Y=2.47
+ $X2=0.347 $Y2=2.385
r151 45 60 3.43356 $w=2.72e-07 $l=1.19143e-07 $layer=LI1_cond $X=0.265 $Y=2.3
+ $X2=0.347 $Y2=2.385
r152 45 47 93.1053 $w=1.88e-07 $l=1.595e-06 $layer=LI1_cond $X=0.265 $Y=2.3
+ $X2=0.265 $Y2=0.705
r153 41 43 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.705 $Y=1.85
+ $X2=6.87 $Y2=1.85
r154 36 38 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.87 $Y=3.075
+ $X2=6.87 $Y2=2.455
r155 35 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.87 $Y=1.925
+ $X2=6.87 $Y2=1.85
r156 35 38 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.87 $Y=1.925
+ $X2=6.87 $Y2=2.455
r157 31 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.705 $Y=1.775
+ $X2=6.705 $Y2=1.85
r158 31 33 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=6.705 $Y=1.775
+ $X2=6.705 $Y2=0.665
r159 30 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.45 $Y=3.15
+ $X2=3.375 $Y2=3.15
r160 29 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.795 $Y=3.15
+ $X2=6.87 $Y2=3.075
r161 29 30 1715.2 $w=1.5e-07 $l=3.345e-06 $layer=POLY_cond $X=6.795 $Y=3.15
+ $X2=3.45 $Y2=3.15
r162 25 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.375 $Y=3.075
+ $X2=3.375 $Y2=3.15
r163 25 27 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.375 $Y=3.075
+ $X2=3.375 $Y2=2.525
r164 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.735 $Y=0.255
+ $X2=2.735 $Y2=0.805
r165 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.66 $Y=0.18
+ $X2=2.735 $Y2=0.255
r166 19 20 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=2.66 $Y=0.18
+ $X2=1.36 $Y2=0.18
r167 18 62 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.285 $Y=0.705
+ $X2=1.285 $Y2=1.495
r168 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.285 $Y=0.255
+ $X2=1.36 $Y2=0.18
r169 15 18 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.285 $Y=0.255
+ $X2=1.285 $Y2=0.705
r170 13 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.3 $Y=3.15
+ $X2=3.375 $Y2=3.15
r171 13 14 1102.45 $w=1.5e-07 $l=2.15e-06 $layer=POLY_cond $X=3.3 $Y=3.15
+ $X2=1.15 $Y2=3.15
r172 12 39 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.075 $Y=2.645
+ $X2=1.075 $Y2=2.165
r173 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.075 $Y=3.075
+ $X2=1.15 $Y2=3.15
r174 10 12 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.075 $Y=3.075
+ $X2=1.075 $Y2=2.645
r175 8 39 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.18 $Y=1.985
+ $X2=1.18 $Y2=2.165
r176 7 58 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.18 $Y=1.675
+ $X2=1.18 $Y2=1.66
r177 7 8 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.18 $Y=1.675
+ $X2=1.18 $Y2=1.985
r178 2 51 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.285
+ $Y=2.325 $X2=0.41 $Y2=2.47
r179 1 47 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.495 $X2=0.275 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_1398_65# 1 2 9 11 12 14 15 16 19 21 23 27
+ 29 30 33 36
c92 19 0 1.28829e-19 $X=7.945 $Y=2.495
r93 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.61 $Y=2.6
+ $X2=9.61 $Y2=2.6
r94 33 35 24.2352 $w=3.38e-07 $l=7.15e-07 $layer=LI1_cond $X=9.605 $Y=1.885
+ $X2=9.605 $Y2=2.6
r95 31 33 49.1483 $w=3.38e-07 $l=1.45e-06 $layer=LI1_cond $X=9.605 $Y=0.435
+ $X2=9.605 $Y2=1.885
r96 29 31 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=9.435 $Y=0.35
+ $X2=9.605 $Y2=0.435
r97 29 30 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=9.435 $Y=0.35
+ $X2=8.575 $Y2=0.35
r98 25 30 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=8.445 $Y=0.435
+ $X2=8.575 $Y2=0.35
r99 25 27 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=8.445 $Y=0.435
+ $X2=8.445 $Y2=0.62
r100 24 36 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=9.61 $Y=3.075
+ $X2=9.61 $Y2=2.6
r101 22 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.02 $Y=3.15
+ $X2=7.945 $Y2=3.15
r102 21 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=9.445 $Y=3.15
+ $X2=9.61 $Y2=3.075
r103 21 22 730.691 $w=1.5e-07 $l=1.425e-06 $layer=POLY_cond $X=9.445 $Y=3.15
+ $X2=8.02 $Y2=3.15
r104 17 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.945 $Y=3.075
+ $X2=7.945 $Y2=3.15
r105 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.945 $Y=3.075
+ $X2=7.945 $Y2=2.495
r106 15 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.87 $Y=3.15
+ $X2=7.945 $Y2=3.15
r107 15 16 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.87 $Y=3.15
+ $X2=7.53 $Y2=3.15
r108 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.455 $Y=3.075
+ $X2=7.53 $Y2=3.15
r109 13 14 789.66 $w=1.5e-07 $l=1.54e-06 $layer=POLY_cond $X=7.455 $Y=1.535
+ $X2=7.455 $Y2=3.075
r110 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.38 $Y=1.46
+ $X2=7.455 $Y2=1.535
r111 11 12 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.38 $Y=1.46
+ $X2=7.14 $Y2=1.46
r112 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.065 $Y=1.385
+ $X2=7.14 $Y2=1.46
r113 7 9 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=7.065 $Y=1.385
+ $X2=7.065 $Y2=0.665
r114 2 33 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=9.41
+ $Y=1.675 $X2=9.55 $Y2=1.885
r115 1 27 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=8.27
+ $Y=0.455 $X2=8.41 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_1247_47# 1 2 3 10 12 13 14 18 19 21 22 26
+ 30 32 33 36 39 40 44 47 48 50 51 53 58 60 64
c121 22 0 3.92666e-20 $X=10.21 $Y=1.49
c122 10 0 1.34614e-19 $X=8.195 $Y=0.345
r123 59 60 5.33595 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=8.745 $Y=1.08
+ $X2=8.655 $Y2=1.08
r124 53 56 3.77163 $w=2.73e-07 $l=9e-08 $layer=LI1_cond $X=6.657 $Y=2.1
+ $X2=6.657 $Y2=2.19
r125 51 65 87.4515 $w=4.75e-07 $l=5.05e-07 $layer=POLY_cond $X=9.172 $Y=0.7
+ $X2=9.172 $Y2=1.205
r126 51 64 47.6426 $w=4.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.172 $Y=0.7
+ $X2=9.172 $Y2=0.535
r127 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.1 $Y=0.7
+ $X2=9.1 $Y2=0.7
r128 48 59 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=9.1 $Y=1.08
+ $X2=8.745 $Y2=1.08
r129 48 50 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=9.1 $Y=0.955
+ $X2=9.1 $Y2=0.7
r130 47 58 3.58051 $w=2.6e-07 $l=1.18427e-07 $layer=LI1_cond $X=8.745 $Y=2.015
+ $X2=8.665 $Y2=2.1
r131 46 59 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=8.745 $Y=1.205
+ $X2=8.745 $Y2=1.08
r132 46 47 49.9091 $w=1.78e-07 $l=8.1e-07 $layer=LI1_cond $X=8.745 $Y=1.205
+ $X2=8.745 $Y2=2.015
r133 42 58 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.665 $Y=2.185
+ $X2=8.665 $Y2=2.1
r134 42 44 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=8.665 $Y=2.185
+ $X2=8.665 $Y2=2.495
r135 41 53 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=6.795 $Y=2.1
+ $X2=6.657 $Y2=2.1
r136 40 58 2.90867 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.495 $Y=2.1
+ $X2=8.665 $Y2=2.1
r137 40 41 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=8.495 $Y=2.1
+ $X2=6.795 $Y2=2.1
r138 39 60 127.219 $w=1.68e-07 $l=1.95e-06 $layer=LI1_cond $X=6.705 $Y=1.04
+ $X2=8.655 $Y2=1.04
r139 34 39 9.18857 $w=1.7e-07 $l=2.87374e-07 $layer=LI1_cond $X=6.457 $Y=0.955
+ $X2=6.705 $Y2=1.04
r140 34 36 13.6522 $w=4.93e-07 $l=5.65e-07 $layer=LI1_cond $X=6.457 $Y=0.955
+ $X2=6.457 $Y2=0.39
r141 28 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.285 $Y=1.565
+ $X2=10.285 $Y2=1.49
r142 28 30 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=10.285 $Y=1.565
+ $X2=10.285 $Y2=2.465
r143 24 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.285 $Y=1.415
+ $X2=10.285 $Y2=1.49
r144 24 26 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=10.285 $Y=1.415
+ $X2=10.285 $Y2=0.665
r145 23 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.41 $Y=1.49
+ $X2=9.335 $Y2=1.49
r146 22 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.21 $Y=1.49
+ $X2=10.285 $Y2=1.49
r147 22 23 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=10.21 $Y=1.49
+ $X2=9.41 $Y2=1.49
r148 19 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.335 $Y=1.565
+ $X2=9.335 $Y2=1.49
r149 19 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.335 $Y=1.565
+ $X2=9.335 $Y2=1.885
r150 18 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.335 $Y=1.415
+ $X2=9.335 $Y2=1.49
r151 18 65 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.335 $Y=1.415
+ $X2=9.335 $Y2=1.205
r152 15 64 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.01 $Y=0.345
+ $X2=9.01 $Y2=0.535
r153 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.935 $Y=0.27
+ $X2=9.01 $Y2=0.345
r154 13 14 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=8.935 $Y=0.27
+ $X2=8.27 $Y2=0.27
r155 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.195 $Y=0.345
+ $X2=8.27 $Y2=0.27
r156 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.195 $Y=0.345
+ $X2=8.195 $Y2=0.665
r157 3 44 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.45
+ $Y=2.285 $X2=8.59 $Y2=2.495
r158 2 56 600 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_PDIFF $count=1 $X=6.42
+ $Y=2.035 $X2=6.63 $Y2=2.19
r159 1 36 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=6.235
+ $Y=0.235 $X2=6.375 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_1989_49# 1 2 9 13 17 21 25 29 33 37 41 45
+ 54 57 64
c95 54 0 3.92666e-20 $X=11.81 $Y=1.51
r96 61 62 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=11.145 $Y=1.51
+ $X2=11.575 $Y2=1.51
r97 55 64 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=11.81 $Y=1.51
+ $X2=12.005 $Y2=1.51
r98 55 62 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=11.81 $Y=1.51
+ $X2=11.575 $Y2=1.51
r99 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.81
+ $Y=1.51 $X2=11.81 $Y2=1.51
r100 52 61 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=10.79 $Y=1.51
+ $X2=11.145 $Y2=1.51
r101 52 58 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.79 $Y=1.51
+ $X2=10.715 $Y2=1.51
r102 51 54 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=10.79 $Y=1.51
+ $X2=11.81 $Y2=1.51
r103 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.79
+ $Y=1.51 $X2=10.79 $Y2=1.51
r104 49 57 2.87242 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.205 $Y=1.51
+ $X2=10.075 $Y2=1.51
r105 49 51 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=10.205 $Y=1.51
+ $X2=10.79 $Y2=1.51
r106 45 47 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=10.075 $Y=1.98
+ $X2=10.075 $Y2=2.91
r107 43 57 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=10.075 $Y=1.595
+ $X2=10.075 $Y2=1.51
r108 43 45 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=10.075 $Y=1.595
+ $X2=10.075 $Y2=1.98
r109 39 57 3.6114 $w=2.57e-07 $l=8.6487e-08 $layer=LI1_cond $X=10.072 $Y=1.425
+ $X2=10.075 $Y2=1.51
r110 39 41 45.4198 $w=2.53e-07 $l=1.005e-06 $layer=LI1_cond $X=10.072 $Y=1.425
+ $X2=10.072 $Y2=0.42
r111 35 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.005 $Y=1.675
+ $X2=12.005 $Y2=1.51
r112 35 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=12.005 $Y=1.675
+ $X2=12.005 $Y2=2.465
r113 31 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.005 $Y=1.345
+ $X2=12.005 $Y2=1.51
r114 31 33 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=12.005 $Y=1.345
+ $X2=12.005 $Y2=0.665
r115 27 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.575 $Y=1.675
+ $X2=11.575 $Y2=1.51
r116 27 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.575 $Y=1.675
+ $X2=11.575 $Y2=2.465
r117 23 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.575 $Y=1.345
+ $X2=11.575 $Y2=1.51
r118 23 25 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=11.575 $Y=1.345
+ $X2=11.575 $Y2=0.665
r119 19 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.145 $Y=1.675
+ $X2=11.145 $Y2=1.51
r120 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.145 $Y=1.675
+ $X2=11.145 $Y2=2.465
r121 15 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.145 $Y=1.345
+ $X2=11.145 $Y2=1.51
r122 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=11.145 $Y=1.345
+ $X2=11.145 $Y2=0.665
r123 11 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.715 $Y=1.675
+ $X2=10.715 $Y2=1.51
r124 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.715 $Y=1.675
+ $X2=10.715 $Y2=2.465
r125 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.715 $Y=1.345
+ $X2=10.715 $Y2=1.51
r126 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=10.715 $Y=1.345
+ $X2=10.715 $Y2=0.665
r127 2 47 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=9.945
+ $Y=1.835 $X2=10.07 $Y2=2.91
r128 2 45 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.945
+ $Y=1.835 $X2=10.07 $Y2=1.98
r129 1 41 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=9.945
+ $Y=0.245 $X2=10.07 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 32 36 40 42 46 52 56
+ 60 66 70 72 77 78 80 81 83 84 85 87 92 116 120 126 129 132 135 138 142
c163 36 0 5.22509e-20 $X=2.3 $Y=2.55
r164 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r165 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r166 135 136 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r167 133 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r168 132 133 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r169 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r170 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r171 124 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r172 124 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r173 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r174 121 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.525 $Y=3.33
+ $X2=11.36 $Y2=3.33
r175 121 123 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=11.525 $Y=3.33
+ $X2=11.76 $Y2=3.33
r176 120 141 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=12.055 $Y=3.33
+ $X2=12.267 $Y2=3.33
r177 120 123 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.055 $Y=3.33
+ $X2=11.76 $Y2=3.33
r178 119 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r179 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r180 116 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.195 $Y=3.33
+ $X2=11.36 $Y2=3.33
r181 116 118 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.195 $Y=3.33
+ $X2=10.8 $Y2=3.33
r182 115 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r183 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r184 112 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r185 111 114 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r186 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r187 109 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r188 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r189 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r190 105 106 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r191 103 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r192 102 105 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.92 $Y2=3.33
r193 102 103 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r194 100 135 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.145 $Y2=3.33
r195 100 102 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.52 $Y2=3.33
r196 99 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r197 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r198 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r199 96 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r200 95 98 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r201 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r202 93 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.3 $Y2=3.33
r203 93 95 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.64 $Y2=3.33
r204 92 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=3.33
+ $X2=3.97 $Y2=3.33
r205 92 98 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.805 $Y=3.33
+ $X2=3.6 $Y2=3.33
r206 91 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r207 91 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r208 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r209 88 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.86 $Y2=3.33
r210 88 90 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 87 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=3.33
+ $X2=2.3 $Y2=3.33
r212 87 90 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.135 $Y=3.33 $X2=1.2
+ $Y2=3.33
r213 85 106 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=7.92 $Y2=3.33
r214 85 103 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=5.52 $Y2=3.33
r215 83 114 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=10.375 $Y=3.33
+ $X2=10.32 $Y2=3.33
r216 83 84 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=10.375 $Y=3.33
+ $X2=10.502 $Y2=3.33
r217 82 118 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.63 $Y=3.33
+ $X2=10.8 $Y2=3.33
r218 82 84 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=10.63 $Y=3.33
+ $X2=10.502 $Y2=3.33
r219 80 108 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.005 $Y=3.33
+ $X2=8.88 $Y2=3.33
r220 80 81 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.005 $Y=3.33
+ $X2=9.135 $Y2=3.33
r221 79 111 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=9.265 $Y=3.33
+ $X2=9.36 $Y2=3.33
r222 79 81 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.265 $Y=3.33
+ $X2=9.135 $Y2=3.33
r223 77 105 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.995 $Y=3.33
+ $X2=7.92 $Y2=3.33
r224 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.995 $Y=3.33
+ $X2=8.16 $Y2=3.33
r225 76 108 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=8.325 $Y=3.33
+ $X2=8.88 $Y2=3.33
r226 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.325 $Y=3.33
+ $X2=8.16 $Y2=3.33
r227 72 75 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=12.22 $Y=2.19
+ $X2=12.22 $Y2=2.95
r228 70 141 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=12.22 $Y=3.245
+ $X2=12.267 $Y2=3.33
r229 70 75 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=12.22 $Y=3.245
+ $X2=12.22 $Y2=2.95
r230 66 69 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=11.36 $Y=2.19
+ $X2=11.36 $Y2=2.97
r231 64 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.36 $Y=3.245
+ $X2=11.36 $Y2=3.33
r232 64 69 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=11.36 $Y=3.245
+ $X2=11.36 $Y2=2.97
r233 60 63 44.7419 $w=2.53e-07 $l=9.9e-07 $layer=LI1_cond $X=10.502 $Y=1.96
+ $X2=10.502 $Y2=2.95
r234 58 84 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=10.502 $Y=3.245
+ $X2=10.502 $Y2=3.33
r235 58 63 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=10.502 $Y=3.245
+ $X2=10.502 $Y2=2.95
r236 54 81 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.135 $Y=3.245
+ $X2=9.135 $Y2=3.33
r237 54 56 60.2816 $w=2.58e-07 $l=1.36e-06 $layer=LI1_cond $X=9.135 $Y=3.245
+ $X2=9.135 $Y2=1.885
r238 50 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.16 $Y=3.245
+ $X2=8.16 $Y2=3.33
r239 50 52 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=8.16 $Y=3.245
+ $X2=8.16 $Y2=2.495
r240 46 49 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=5.145 $Y=2.27
+ $X2=5.145 $Y2=2.61
r241 44 135 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=3.33
r242 44 49 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=5.145 $Y=3.245
+ $X2=5.145 $Y2=2.61
r243 43 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=3.33
+ $X2=3.97 $Y2=3.33
r244 42 135 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.015 $Y=3.33
+ $X2=5.145 $Y2=3.33
r245 42 43 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=5.015 $Y=3.33
+ $X2=4.135 $Y2=3.33
r246 38 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=3.245
+ $X2=3.97 $Y2=3.33
r247 38 40 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=3.97 $Y=3.245
+ $X2=3.97 $Y2=2.525
r248 34 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=3.245
+ $X2=2.3 $Y2=3.33
r249 34 36 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.3 $Y=3.245
+ $X2=2.3 $Y2=2.55
r250 30 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=3.245
+ $X2=0.86 $Y2=3.33
r251 30 32 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.86 $Y=3.245
+ $X2=0.86 $Y2=2.765
r252 9 75 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=12.08
+ $Y=1.835 $X2=12.22 $Y2=2.95
r253 9 72 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=12.08
+ $Y=1.835 $X2=12.22 $Y2=2.19
r254 8 69 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=11.22
+ $Y=1.835 $X2=11.36 $Y2=2.97
r255 8 66 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=11.22
+ $Y=1.835 $X2=11.36 $Y2=2.19
r256 7 63 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=10.36
+ $Y=1.835 $X2=10.5 $Y2=2.95
r257 7 60 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=10.36
+ $Y=1.835 $X2=10.5 $Y2=1.96
r258 6 56 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=8.995
+ $Y=1.675 $X2=9.12 $Y2=1.885
r259 5 52 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.02
+ $Y=2.285 $X2=8.16 $Y2=2.495
r260 4 49 600 $w=1.7e-07 $l=5.22063e-07 $layer=licon1_PDIFF $count=1 $X=4.785
+ $Y=2.315 $X2=5.18 $Y2=2.61
r261 4 46 600 $w=1.7e-07 $l=4.16893e-07 $layer=licon1_PDIFF $count=1 $X=4.785
+ $Y=2.315 $X2=5.18 $Y2=2.27
r262 3 40 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=2.315 $X2=3.97 $Y2=2.525
r263 2 36 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.175
+ $Y=2.405 $X2=2.3 $Y2=2.55
r264 1 32 600 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=2.325 $X2=0.86 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_476_119# 1 2 9 13 19 21 22
c48 22 0 1.87691e-19 $X=2.792 $Y=2.085
c49 21 0 4.42586e-20 $X=2.792 $Y=1.915
r50 21 22 9.32577 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.792 $Y=1.915
+ $X2=2.792 $Y2=2.085
r51 15 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=1.255
+ $X2=2.865 $Y2=1.17
r52 15 21 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.865 $Y=1.255
+ $X2=2.865 $Y2=1.915
r53 13 22 22.0467 $w=2.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.75 $Y=2.525
+ $X2=2.75 $Y2=2.085
r54 7 19 22.3775 $w=1.68e-07 $l=3.43e-07 $layer=LI1_cond $X=2.522 $Y=1.17
+ $X2=2.865 $Y2=1.17
r55 7 9 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=2.522 $Y=1.085
+ $X2=2.522 $Y2=0.805
r56 2 13 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=2.315 $X2=2.73 $Y2=2.525
r57 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.595 $X2=2.52 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_1094_379# 1 2 9 11 13
c27 11 0 1.62847e-19 $X=5.775 $Y=2.965
r28 11 13 77.9136 $w=1.98e-07 $l=1.405e-06 $layer=LI1_cond $X=5.775 $Y=2.965
+ $X2=7.18 $Y2=2.965
r29 7 11 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=5.61 $Y=2.865
+ $X2=5.775 $Y2=2.965
r30 7 9 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=5.61 $Y=2.865
+ $X2=5.61 $Y2=2.25
r31 2 13 600 $w=1.7e-07 $l=1.03586e-06 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=2.035 $X2=7.18 $Y2=2.96
r32 1 9 300 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=2 $X=5.47
+ $Y=1.895 $X2=5.61 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%A_1201_407# 1 2 9 11 12 14
c29 11 0 1.19092e-19 $X=7.565 $Y=2.61
r30 14 16 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=7.695 $Y=2.52
+ $X2=7.695 $Y2=2.61
r31 11 16 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.565 $Y=2.61
+ $X2=7.695 $Y2=2.61
r32 11 12 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=7.565 $Y=2.61
+ $X2=6.295 $Y2=2.61
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.13 $Y=2.525
+ $X2=6.295 $Y2=2.61
r34 7 9 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.13 $Y=2.525 $X2=6.13
+ $Y2=2.245
r35 2 14 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=7.605
+ $Y=2.285 $X2=7.73 $Y2=2.52
r36 1 9 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=6.005
+ $Y=2.035 $X2=6.13 $Y2=2.245
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%Q 1 2 3 4 15 19 23 24 25 26 29 33 37 39 41
+ 42 44 47 49
c60 37 0 7.44113e-20 $X=12.145 $Y=1.16
r61 47 49 2.35192 $w=2.43e-07 $l=5e-08 $layer=LI1_cond $X=12.267 $Y=1.245
+ $X2=12.267 $Y2=1.295
r62 44 47 2.91961 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=12.267 $Y=1.16
+ $X2=12.267 $Y2=1.245
r63 44 49 0.799654 $w=2.43e-07 $l=1.7e-08 $layer=LI1_cond $X=12.267 $Y=1.312
+ $X2=12.267 $Y2=1.295
r64 43 44 21.3084 $w=2.43e-07 $l=4.53e-07 $layer=LI1_cond $X=12.267 $Y=1.765
+ $X2=12.267 $Y2=1.312
r65 40 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=11.885 $Y=1.85
+ $X2=11.79 $Y2=1.85
r66 39 43 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=12.145 $Y=1.85
+ $X2=12.267 $Y2=1.765
r67 39 40 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.145 $Y=1.85
+ $X2=11.885 $Y2=1.85
r68 38 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=11.885 $Y=1.16
+ $X2=11.79 $Y2=1.16
r69 37 44 4.1905 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=12.145 $Y=1.16
+ $X2=12.267 $Y2=1.16
r70 37 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.145 $Y=1.16
+ $X2=11.885 $Y2=1.16
r71 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=11.79 $Y=1.98
+ $X2=11.79 $Y2=2.91
r72 31 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.79 $Y=1.935
+ $X2=11.79 $Y2=1.85
r73 31 33 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=11.79 $Y=1.935
+ $X2=11.79 $Y2=1.98
r74 27 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.79 $Y=1.075
+ $X2=11.79 $Y2=1.16
r75 27 29 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=11.79 $Y=1.075
+ $X2=11.79 $Y2=0.42
r76 25 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=11.695 $Y=1.85
+ $X2=11.79 $Y2=1.85
r77 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.695 $Y=1.85
+ $X2=11.025 $Y2=1.85
r78 23 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=11.695 $Y=1.16
+ $X2=11.79 $Y2=1.16
r79 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.695 $Y=1.16
+ $X2=11.025 $Y2=1.16
r80 19 21 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=10.912 $Y=1.98
+ $X2=10.912 $Y2=2.91
r81 17 26 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=10.912 $Y=1.935
+ $X2=11.025 $Y2=1.85
r82 17 19 2.30489 $w=2.23e-07 $l=4.5e-08 $layer=LI1_cond $X=10.912 $Y=1.935
+ $X2=10.912 $Y2=1.98
r83 13 24 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=10.912 $Y=1.075
+ $X2=11.025 $Y2=1.16
r84 13 15 33.5489 $w=2.23e-07 $l=6.55e-07 $layer=LI1_cond $X=10.912 $Y=1.075
+ $X2=10.912 $Y2=0.42
r85 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=11.65
+ $Y=1.835 $X2=11.79 $Y2=2.91
r86 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.65
+ $Y=1.835 $X2=11.79 $Y2=1.98
r87 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.79
+ $Y=1.835 $X2=10.93 $Y2=2.91
r88 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.79
+ $Y=1.835 $X2=10.93 $Y2=1.98
r89 2 29 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=11.65
+ $Y=0.245 $X2=11.79 $Y2=0.42
r90 1 15 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=10.79
+ $Y=0.245 $X2=10.93 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_4%VGND 1 2 3 4 5 6 7 8 27 31 33 37 41 45 49 51
+ 53 56 57 59 60 61 67 71 76 91 95 101 104 112 116 119 123
c156 112 0 1.6457e-20 $X=5.585 $Y=0.38
c157 8 0 7.44113e-20 $X=12.08 $Y=0.245
r158 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r159 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r160 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r161 112 114 1.1361 $w=6.98e-07 $l=6.5e-08 $layer=LI1_cond $X=5.327 $Y=0.38
+ $X2=5.327 $Y2=0.445
r162 108 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r163 107 112 6.64183 $w=6.98e-07 $l=3.8e-07 $layer=LI1_cond $X=5.327 $Y=0
+ $X2=5.327 $Y2=0.38
r164 107 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r165 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r166 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r167 102 105 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=3.6 $Y2=0
r168 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r169 99 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r170 99 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r171 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r172 96 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.525 $Y=0
+ $X2=11.36 $Y2=0
r173 96 98 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=11.525 $Y=0
+ $X2=11.76 $Y2=0
r174 95 122 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=12.267 $Y2=0
r175 95 98 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=11.76 $Y2=0
r176 94 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r177 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r178 91 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.195 $Y=0
+ $X2=11.36 $Y2=0
r179 91 93 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.195 $Y=0
+ $X2=10.8 $Y2=0
r180 90 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r181 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r182 87 90 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=10.32 $Y2=0
r183 87 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r184 86 89 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=10.32
+ $Y2=0
r185 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r186 84 116 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.145 $Y=0
+ $X2=7.81 $Y2=0
r187 84 86 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.145 $Y=0 $X2=8.4
+ $Y2=0
r188 83 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r189 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r190 80 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r191 79 82 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=0 $X2=7.44
+ $Y2=0
r192 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r193 77 107 9.30268 $w=1.7e-07 $l=4.23e-07 $layer=LI1_cond $X=5.75 $Y=0
+ $X2=5.327 $Y2=0
r194 77 79 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=6
+ $Y2=0
r195 76 116 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=7.81 $Y2=0
r196 76 82 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.475 $Y=0 $X2=7.44
+ $Y2=0
r197 75 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r198 75 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r199 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r200 72 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=0
+ $X2=3.74 $Y2=0
r201 72 74 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.905 $Y=0
+ $X2=4.56 $Y2=0
r202 71 107 9.30268 $w=1.7e-07 $l=4.22e-07 $layer=LI1_cond $X=4.905 $Y=0
+ $X2=5.327 $Y2=0
r203 71 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.905 $Y=0 $X2=4.56
+ $Y2=0
r204 70 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r205 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r206 67 101 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=2.105 $Y2=0
r207 67 69 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=1.68 $Y2=0
r208 65 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r209 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r210 61 83 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=6.24 $Y=0 $X2=7.44
+ $Y2=0
r211 61 80 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=0 $X2=6
+ $Y2=0
r212 59 89 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=10.37 $Y=0 $X2=10.32
+ $Y2=0
r213 59 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.37 $Y=0 $X2=10.5
+ $Y2=0
r214 58 93 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.63 $Y=0 $X2=10.8
+ $Y2=0
r215 58 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.63 $Y=0 $X2=10.5
+ $Y2=0
r216 56 64 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0
+ $X2=0.72 $Y2=0
r217 56 57 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.095
+ $Y2=0
r218 55 69 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=1.68 $Y2=0
r219 55 57 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.095
+ $Y2=0
r220 51 122 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=12.22 $Y=0.085
+ $X2=12.267 $Y2=0
r221 51 53 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=12.22 $Y=0.085
+ $X2=12.22 $Y2=0.39
r222 47 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.36 $Y=0.085
+ $X2=11.36 $Y2=0
r223 47 49 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=11.36 $Y=0.085
+ $X2=11.36 $Y2=0.39
r224 43 60 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0
r225 43 45 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=10.5 $Y=0.085
+ $X2=10.5 $Y2=0.39
r226 39 116 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0
r227 39 41 10.1756 $w=6.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0.655
r228 35 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=0.085
+ $X2=3.74 $Y2=0
r229 35 37 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.74 $Y=0.085
+ $X2=3.74 $Y2=0.72
r230 34 101 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.105 $Y2=0
r231 33 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=0
+ $X2=3.74 $Y2=0
r232 33 34 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.575 $Y=0
+ $X2=2.225 $Y2=0
r233 29 101 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r234 29 31 34.5733 $w=2.38e-07 $l=7.2e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.805
r235 25 57 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=0.085
+ $X2=1.095 $Y2=0
r236 25 27 32.4779 $w=2.18e-07 $l=6.2e-07 $layer=LI1_cond $X=1.095 $Y=0.085
+ $X2=1.095 $Y2=0.705
r237 8 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.08
+ $Y=0.245 $X2=12.22 $Y2=0.39
r238 7 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.22
+ $Y=0.245 $X2=11.36 $Y2=0.39
r239 6 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.36
+ $Y=0.245 $X2=10.5 $Y2=0.39
r240 5 41 91 $w=1.7e-07 $l=5.71314e-07 $layer=licon1_NDIFF $count=2 $X=7.5
+ $Y=0.455 $X2=7.98 $Y2=0.655
r241 4 114 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.235 $X2=5.07 $Y2=0.445
r242 4 112 91 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_NDIFF $count=2 $X=4.93
+ $Y=0.235 $X2=5.585 $Y2=0.38
r243 3 37 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.6
+ $Y=0.595 $X2=3.74 $Y2=0.72
r244 2 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.595 $X2=2.09 $Y2=0.805
r245 1 27 182 $w=1.7e-07 $l=6.00895e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.495 $X2=1.07 $Y2=0.705
.ends

