* File: sky130_fd_sc_lp__o32a_1.pxi.spice
* Created: Fri Aug 28 11:17:17 2020
* 
x_PM_SKY130_FD_SC_LP__O32A_1%A_88_269# N_A_88_269#_M1000_d N_A_88_269#_M1007_d
+ N_A_88_269#_M1009_g N_A_88_269#_M1004_g N_A_88_269#_c_66_n N_A_88_269#_c_76_p
+ N_A_88_269#_c_132_p N_A_88_269#_c_89_p N_A_88_269#_c_108_p N_A_88_269#_c_100_p
+ N_A_88_269#_c_67_n N_A_88_269#_c_68_n N_A_88_269#_c_69_n N_A_88_269#_c_94_p
+ N_A_88_269#_c_104_p PM_SKY130_FD_SC_LP__O32A_1%A_88_269#
x_PM_SKY130_FD_SC_LP__O32A_1%A1 N_A1_M1006_g N_A1_M1010_g A1 A1 N_A1_c_154_n
+ N_A1_c_155_n PM_SKY130_FD_SC_LP__O32A_1%A1
x_PM_SKY130_FD_SC_LP__O32A_1%A2 N_A2_M1001_g N_A2_M1008_g A2 A2 N_A2_c_193_n
+ N_A2_c_194_n PM_SKY130_FD_SC_LP__O32A_1%A2
x_PM_SKY130_FD_SC_LP__O32A_1%A3 N_A3_M1007_g N_A3_c_228_n N_A3_M1003_g A3 A3
+ N_A3_c_230_n PM_SKY130_FD_SC_LP__O32A_1%A3
x_PM_SKY130_FD_SC_LP__O32A_1%B2 N_B2_M1000_g N_B2_M1002_g B2 N_B2_c_267_n
+ N_B2_c_268_n PM_SKY130_FD_SC_LP__O32A_1%B2
x_PM_SKY130_FD_SC_LP__O32A_1%B1 N_B1_c_305_n N_B1_M1011_g N_B1_M1005_g B1 B1 B1
+ N_B1_c_308_n PM_SKY130_FD_SC_LP__O32A_1%B1
x_PM_SKY130_FD_SC_LP__O32A_1%X N_X_M1004_s N_X_M1009_s N_X_c_339_n N_X_c_340_n
+ N_X_c_336_n X X N_X_c_337_n X PM_SKY130_FD_SC_LP__O32A_1%X
x_PM_SKY130_FD_SC_LP__O32A_1%VPWR N_VPWR_M1009_d N_VPWR_M1005_d N_VPWR_c_361_n
+ N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n VPWR
+ N_VPWR_c_366_n N_VPWR_c_360_n PM_SKY130_FD_SC_LP__O32A_1%VPWR
x_PM_SKY130_FD_SC_LP__O32A_1%VGND N_VGND_M1004_d N_VGND_M1001_d N_VGND_c_409_n
+ N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n VGND N_VGND_c_413_n
+ N_VGND_c_414_n N_VGND_c_415_n PM_SKY130_FD_SC_LP__O32A_1%VGND
x_PM_SKY130_FD_SC_LP__O32A_1%A_250_69# N_A_250_69#_M1006_d N_A_250_69#_M1003_d
+ N_A_250_69#_M1011_d N_A_250_69#_c_450_n N_A_250_69#_c_460_n
+ N_A_250_69#_c_457_n N_A_250_69#_c_451_n N_A_250_69#_c_452_n
+ N_A_250_69#_c_453_n PM_SKY130_FD_SC_LP__O32A_1%A_250_69#
cc_1 VNB N_A_88_269#_M1004_g 0.0254059f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.765
cc_2 VNB N_A_88_269#_c_66_n 4.2869e-19 $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.93
cc_3 VNB N_A_88_269#_c_67_n 0.00337162f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=1.93
cc_4 VNB N_A_88_269#_c_68_n 0.0279242f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.51
cc_5 VNB N_A_88_269#_c_69_n 0.00644348f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.495
cc_6 VNB N_A1_M1010_g 0.00138691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB A1 0.00570663f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.465
cc_8 VNB N_A1_c_154_n 0.0310924f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.765
cc_9 VNB N_A1_c_155_n 0.0171353f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.645
cc_10 VNB N_A2_M1008_g 0.00131622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A2 0.00508855f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.465
cc_12 VNB N_A2_c_193_n 0.0331995f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.765
cc_13 VNB N_A2_c_194_n 0.0182078f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.645
cc_14 VNB N_A3_M1007_g 0.0014022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_c_228_n 0.0186807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A3 0.00557487f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.465
cc_17 VNB N_A3_c_230_n 0.0326476f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.015
cc_18 VNB N_B2_M1000_g 0.0200388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B2_c_267_n 0.0264797f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.765
cc_20 VNB N_B2_c_268_n 0.00324317f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.765
cc_21 VNB N_B1_c_305_n 0.0197725f $X=-0.19 $Y=-0.245 $X2=2.88 $Y2=0.345
cc_22 VNB N_B1_M1005_g 0.00137508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB B1 0.0215197f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.465
cc_24 VNB N_B1_c_308_n 0.0483409f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.015
cc_25 VNB N_X_c_336_n 0.0232051f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=1.645
cc_26 VNB N_X_c_337_n 0.0332721f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.995
cc_27 VNB X 0.0134875f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=1.175
cc_28 VNB N_VPWR_c_360_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.51
cc_29 VNB N_VGND_c_409_n 0.00810141f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.465
cc_30 VNB N_VGND_c_410_n 0.0154877f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.345
cc_31 VNB N_VGND_c_411_n 0.0224375f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.765
cc_32 VNB N_VGND_c_412_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_413_n 0.038345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_414_n 0.226232f $X=-0.19 $Y=-0.245 $X2=3.09 $Y2=2.015
cc_35 VNB N_VGND_c_415_n 0.017378f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.495
cc_36 VNB N_A_250_69#_c_450_n 0.00244555f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.765
cc_37 VNB N_A_250_69#_c_451_n 0.0123614f $X=-0.19 $Y=-0.245 $X2=2.562 $Y2=2.95
cc_38 VNB N_A_250_69#_c_452_n 0.00239286f $X=-0.19 $Y=-0.245 $X2=2.39 $Y2=2.95
cc_39 VNB N_A_250_69#_c_453_n 0.0230363f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.72
cc_40 VPB N_A_88_269#_M1009_g 0.0242977f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.465
cc_41 VPB N_A_88_269#_c_66_n 0.00146206f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=1.93
cc_42 VPB N_A_88_269#_c_67_n 0.0012959f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=1.93
cc_43 VPB N_A_88_269#_c_68_n 0.00736583f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.51
cc_44 VPB N_A1_M1010_g 0.021178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB A1 0.00255005f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.465
cc_46 VPB N_A2_M1008_g 0.0201502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB A2 0.00290499f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.465
cc_48 VPB N_A3_M1007_g 0.0226039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB A3 0.00329127f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.465
cc_50 VPB N_B2_M1002_g 0.0208994f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.675
cc_51 VPB N_B2_c_267_n 0.00744913f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=0.765
cc_52 VPB N_B2_c_268_n 0.00374531f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=0.765
cc_53 VPB N_B1_M1005_g 0.0206287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB B1 0.0230163f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.465
cc_55 VPB N_X_c_339_n 0.0508238f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.345
cc_56 VPB N_X_c_340_n 0.0148526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_X_c_336_n 0.00785558f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=1.645
cc_58 VPB N_VPWR_c_361_n 0.00561645f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.465
cc_59 VPB N_VPWR_c_362_n 0.0122537f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.345
cc_60 VPB N_VPWR_c_363_n 0.0340705f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=0.765
cc_61 VPB N_VPWR_c_364_n 0.0231511f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=1.93
cc_62 VPB N_VPWR_c_365_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.015
cc_63 VPB N_VPWR_c_366_n 0.0629107f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=0.72
cc_64 VPB N_VPWR_c_360_n 0.0483424f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.51
cc_65 N_A_88_269#_M1009_g N_A1_M1010_g 0.0374687f $X=0.69 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_88_269#_c_66_n N_A1_M1010_g 0.0036314f $X=0.815 $Y=1.93 $X2=0 $Y2=0
cc_67 N_A_88_269#_c_76_p N_A1_M1010_g 0.0158624f $X=2.215 $Y=2.015 $X2=0 $Y2=0
cc_68 N_A_88_269#_c_68_n N_A1_M1010_g 0.00138148f $X=0.605 $Y=1.51 $X2=0 $Y2=0
cc_69 N_A_88_269#_M1009_g A1 2.18647e-19 $X=0.69 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_88_269#_M1004_g A1 0.00197622f $X=0.695 $Y=0.765 $X2=0 $Y2=0
cc_71 N_A_88_269#_c_66_n A1 0.00861942f $X=0.815 $Y=1.93 $X2=0 $Y2=0
cc_72 N_A_88_269#_c_76_p A1 0.0183362f $X=2.215 $Y=2.015 $X2=0 $Y2=0
cc_73 N_A_88_269#_c_68_n A1 3.7042e-19 $X=0.605 $Y=1.51 $X2=0 $Y2=0
cc_74 N_A_88_269#_c_69_n A1 0.0241626f $X=0.815 $Y=1.495 $X2=0 $Y2=0
cc_75 N_A_88_269#_M1004_g N_A1_c_154_n 0.0205945f $X=0.695 $Y=0.765 $X2=0 $Y2=0
cc_76 N_A_88_269#_c_76_p N_A1_c_154_n 0.00335962f $X=2.215 $Y=2.015 $X2=0 $Y2=0
cc_77 N_A_88_269#_c_69_n N_A1_c_154_n 0.00196255f $X=0.815 $Y=1.495 $X2=0 $Y2=0
cc_78 N_A_88_269#_M1004_g N_A1_c_155_n 0.0128218f $X=0.695 $Y=0.765 $X2=0 $Y2=0
cc_79 N_A_88_269#_c_76_p N_A2_M1008_g 0.0153706f $X=2.215 $Y=2.015 $X2=0 $Y2=0
cc_80 N_A_88_269#_c_89_p N_A2_M1008_g 0.00472922f $X=2.39 $Y=2.95 $X2=0 $Y2=0
cc_81 N_A_88_269#_c_76_p A2 0.0208962f $X=2.215 $Y=2.015 $X2=0 $Y2=0
cc_82 N_A_88_269#_c_76_p N_A2_c_193_n 0.00190192f $X=2.215 $Y=2.015 $X2=0 $Y2=0
cc_83 N_A_88_269#_c_76_p N_A3_M1007_g 0.0105324f $X=2.215 $Y=2.015 $X2=0 $Y2=0
cc_84 N_A_88_269#_c_89_p N_A3_M1007_g 0.023734f $X=2.39 $Y=2.95 $X2=0 $Y2=0
cc_85 N_A_88_269#_c_94_p N_A3_M1007_g 0.00103564f $X=2.39 $Y=2.015 $X2=0 $Y2=0
cc_86 N_A_88_269#_c_76_p A3 0.0133528f $X=2.215 $Y=2.015 $X2=0 $Y2=0
cc_87 N_A_88_269#_c_94_p A3 0.0110683f $X=2.39 $Y=2.015 $X2=0 $Y2=0
cc_88 N_A_88_269#_c_94_p N_A3_c_230_n 0.00393327f $X=2.39 $Y=2.015 $X2=0 $Y2=0
cc_89 N_A_88_269#_c_67_n N_B2_M1000_g 0.00340574f $X=3.175 $Y=1.93 $X2=0 $Y2=0
cc_90 N_A_88_269#_c_89_p N_B2_M1002_g 0.0201749f $X=2.39 $Y=2.95 $X2=0 $Y2=0
cc_91 N_A_88_269#_c_100_p N_B2_M1002_g 0.0124101f $X=3.09 $Y=2.015 $X2=0 $Y2=0
cc_92 N_A_88_269#_c_94_p N_B2_M1002_g 0.00118965f $X=2.39 $Y=2.015 $X2=0 $Y2=0
cc_93 N_A_88_269#_c_67_n N_B2_c_267_n 0.00648263f $X=3.175 $Y=1.93 $X2=0 $Y2=0
cc_94 N_A_88_269#_c_94_p N_B2_c_267_n 0.00118218f $X=2.39 $Y=2.015 $X2=0 $Y2=0
cc_95 N_A_88_269#_c_104_p N_B2_c_267_n 0.00479029f $X=3.08 $Y=1.175 $X2=0 $Y2=0
cc_96 N_A_88_269#_c_100_p N_B2_c_268_n 6.93626e-19 $X=3.09 $Y=2.015 $X2=0 $Y2=0
cc_97 N_A_88_269#_c_67_n N_B2_c_268_n 0.0314886f $X=3.175 $Y=1.93 $X2=0 $Y2=0
cc_98 N_A_88_269#_c_94_p N_B2_c_268_n 0.0297407f $X=2.39 $Y=2.015 $X2=0 $Y2=0
cc_99 N_A_88_269#_c_108_p N_B1_c_305_n 0.00478669f $X=3.065 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_88_269#_c_67_n N_B1_c_305_n 0.00327491f $X=3.175 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_88_269#_c_104_p N_B1_c_305_n 0.00645728f $X=3.08 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_88_269#_c_89_p N_B1_M1005_g 0.00310236f $X=2.39 $Y=2.95 $X2=0 $Y2=0
cc_103 N_A_88_269#_c_100_p N_B1_M1005_g 0.00496459f $X=3.09 $Y=2.015 $X2=0 $Y2=0
cc_104 N_A_88_269#_c_67_n N_B1_M1005_g 0.00506996f $X=3.175 $Y=1.93 $X2=0 $Y2=0
cc_105 N_A_88_269#_c_89_p B1 6.55082e-19 $X=2.39 $Y=2.95 $X2=0 $Y2=0
cc_106 N_A_88_269#_c_100_p B1 0.0133537f $X=3.09 $Y=2.015 $X2=0 $Y2=0
cc_107 N_A_88_269#_c_67_n B1 0.0502856f $X=3.175 $Y=1.93 $X2=0 $Y2=0
cc_108 N_A_88_269#_c_67_n N_B1_c_308_n 0.00748906f $X=3.175 $Y=1.93 $X2=0 $Y2=0
cc_109 N_A_88_269#_M1009_g N_X_c_340_n 0.00332321f $X=0.69 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A_88_269#_c_66_n N_X_c_340_n 0.00469872f $X=0.815 $Y=1.93 $X2=0 $Y2=0
cc_111 N_A_88_269#_c_68_n N_X_c_340_n 0.00287432f $X=0.605 $Y=1.51 $X2=0 $Y2=0
cc_112 N_A_88_269#_c_69_n N_X_c_340_n 0.00997021f $X=0.815 $Y=1.495 $X2=0 $Y2=0
cc_113 N_A_88_269#_M1009_g N_X_c_336_n 0.00159211f $X=0.69 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A_88_269#_M1004_g N_X_c_336_n 0.00338369f $X=0.695 $Y=0.765 $X2=0 $Y2=0
cc_115 N_A_88_269#_c_66_n N_X_c_336_n 0.00404815f $X=0.815 $Y=1.93 $X2=0 $Y2=0
cc_116 N_A_88_269#_c_68_n N_X_c_336_n 0.00289787f $X=0.605 $Y=1.51 $X2=0 $Y2=0
cc_117 N_A_88_269#_c_69_n N_X_c_336_n 0.0226832f $X=0.815 $Y=1.495 $X2=0 $Y2=0
cc_118 N_A_88_269#_M1004_g N_X_c_337_n 0.0030598f $X=0.695 $Y=0.765 $X2=0 $Y2=0
cc_119 N_A_88_269#_c_68_n X 0.00359431f $X=0.605 $Y=1.51 $X2=0 $Y2=0
cc_120 N_A_88_269#_c_69_n X 0.0114278f $X=0.815 $Y=1.495 $X2=0 $Y2=0
cc_121 N_A_88_269#_c_66_n N_VPWR_M1009_d 0.00117769f $X=0.815 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_88_269#_c_76_p N_VPWR_M1009_d 0.00723526f $X=2.215 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_88_269#_c_132_p N_VPWR_M1009_d 8.41722e-19 $X=0.9 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_88_269#_M1009_g N_VPWR_c_361_n 0.00816333f $X=0.69 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_88_269#_c_76_p N_VPWR_c_361_n 0.0172929f $X=2.215 $Y=2.015 $X2=0
+ $Y2=0
cc_126 N_A_88_269#_c_132_p N_VPWR_c_361_n 0.00678672f $X=0.9 $Y=2.015 $X2=0
+ $Y2=0
cc_127 N_A_88_269#_c_89_p N_VPWR_c_363_n 0.0286478f $X=2.39 $Y=2.95 $X2=0 $Y2=0
cc_128 N_A_88_269#_M1009_g N_VPWR_c_364_n 0.00585385f $X=0.69 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_A_88_269#_c_89_p N_VPWR_c_366_n 0.0445342f $X=2.39 $Y=2.95 $X2=0 $Y2=0
cc_130 N_A_88_269#_M1007_d N_VPWR_c_360_n 0.00505717f $X=2.25 $Y=1.835 $X2=0
+ $Y2=0
cc_131 N_A_88_269#_M1009_g N_VPWR_c_360_n 0.0121002f $X=0.69 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_A_88_269#_c_89_p N_VPWR_c_360_n 0.0264619f $X=2.39 $Y=2.95 $X2=0 $Y2=0
cc_133 N_A_88_269#_c_76_p A_264_367# 0.0140113f $X=2.215 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_134 N_A_88_269#_c_76_p A_358_367# 0.0131285f $X=2.215 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A_88_269#_c_100_p A_604_367# 0.0046148f $X=3.09 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_88_269#_c_67_n A_604_367# 0.00103702f $X=3.175 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A_88_269#_M1004_g N_VGND_c_409_n 0.00338181f $X=0.695 $Y=0.765 $X2=0
+ $Y2=0
cc_138 N_A_88_269#_c_69_n N_VGND_c_409_n 0.00566627f $X=0.815 $Y=1.495 $X2=0
+ $Y2=0
cc_139 N_A_88_269#_M1004_g N_VGND_c_411_n 0.00480781f $X=0.695 $Y=0.765 $X2=0
+ $Y2=0
cc_140 N_A_88_269#_M1004_g N_VGND_c_414_n 0.00969511f $X=0.695 $Y=0.765 $X2=0
+ $Y2=0
cc_141 N_A_88_269#_M1000_d N_A_250_69#_c_451_n 0.00250873f $X=2.88 $Y=0.345
+ $X2=0 $Y2=0
cc_142 N_A_88_269#_c_108_p N_A_250_69#_c_451_n 0.0198504f $X=3.065 $Y=0.72 $X2=0
+ $Y2=0
cc_143 N_A1_M1010_g N_A2_M1008_g 0.0657736f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_144 A1 N_A2_M1008_g 3.50715e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_145 A1 A2 0.0447637f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A1_c_154_n A2 0.0014248f $X=1.155 $Y=1.46 $X2=0 $Y2=0
cc_147 N_A1_c_155_n A2 2.3177e-19 $X=1.15 $Y=1.295 $X2=0 $Y2=0
cc_148 N_A1_c_154_n N_A2_c_193_n 0.0214254f $X=1.155 $Y=1.46 $X2=0 $Y2=0
cc_149 A1 N_A2_c_194_n 0.00133483f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_150 N_A1_c_155_n N_A2_c_194_n 0.0167608f $X=1.15 $Y=1.295 $X2=0 $Y2=0
cc_151 N_A1_M1010_g N_VPWR_c_361_n 0.00808177f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A1_M1010_g N_VPWR_c_366_n 0.00585385f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A1_M1010_g N_VPWR_c_360_n 0.0112675f $X=1.245 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A1_c_154_n N_VGND_c_409_n 0.00307332f $X=1.155 $Y=1.46 $X2=0 $Y2=0
cc_155 N_A1_c_155_n N_VGND_c_409_n 0.00175009f $X=1.15 $Y=1.295 $X2=0 $Y2=0
cc_156 N_A1_c_155_n N_VGND_c_410_n 0.00480781f $X=1.15 $Y=1.295 $X2=0 $Y2=0
cc_157 N_A1_c_155_n N_VGND_c_414_n 0.00945063f $X=1.15 $Y=1.295 $X2=0 $Y2=0
cc_158 N_A1_c_155_n N_VGND_c_415_n 3.91165e-19 $X=1.15 $Y=1.295 $X2=0 $Y2=0
cc_159 N_A1_c_155_n N_A_250_69#_c_450_n 3.72339e-19 $X=1.15 $Y=1.295 $X2=0 $Y2=0
cc_160 A1 N_A_250_69#_c_457_n 0.0059253f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_161 N_A1_c_154_n N_A_250_69#_c_457_n 2.19594e-19 $X=1.155 $Y=1.46 $X2=0 $Y2=0
cc_162 N_A2_M1008_g N_A3_M1007_g 0.0666343f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_163 A2 N_A3_M1007_g 3.94569e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A2_c_194_n N_A3_c_228_n 0.0118618f $X=1.71 $Y=1.295 $X2=0 $Y2=0
cc_165 N_A2_M1008_g A3 4.30812e-19 $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_166 A2 A3 0.0445838f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_167 N_A2_c_193_n A3 0.00207333f $X=1.725 $Y=1.46 $X2=0 $Y2=0
cc_168 N_A2_c_194_n A3 2.5317e-19 $X=1.71 $Y=1.295 $X2=0 $Y2=0
cc_169 A2 N_A3_c_230_n 3.23461e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A2_c_193_n N_A3_c_230_n 0.0206395f $X=1.725 $Y=1.46 $X2=0 $Y2=0
cc_171 N_A2_M1008_g N_VPWR_c_366_n 0.00585385f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A2_M1008_g N_VPWR_c_360_n 0.0112127f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A2_c_194_n N_VGND_c_410_n 0.00401871f $X=1.71 $Y=1.295 $X2=0 $Y2=0
cc_174 N_A2_c_194_n N_VGND_c_414_n 0.00775088f $X=1.71 $Y=1.295 $X2=0 $Y2=0
cc_175 N_A2_c_194_n N_VGND_c_415_n 0.00963058f $X=1.71 $Y=1.295 $X2=0 $Y2=0
cc_176 N_A2_c_194_n N_A_250_69#_c_450_n 3.53182e-19 $X=1.71 $Y=1.295 $X2=0 $Y2=0
cc_177 A2 N_A_250_69#_c_460_n 0.022686f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A2_c_193_n N_A_250_69#_c_460_n 0.00238843f $X=1.725 $Y=1.46 $X2=0 $Y2=0
cc_179 N_A2_c_194_n N_A_250_69#_c_460_n 0.0133633f $X=1.71 $Y=1.295 $X2=0 $Y2=0
cc_180 N_A3_c_228_n N_B2_M1000_g 0.0183633f $X=2.375 $Y=1.295 $X2=0 $Y2=0
cc_181 A3 N_B2_M1000_g 7.11376e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A3_M1007_g N_B2_M1002_g 0.00724472f $X=2.175 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A3_M1007_g N_B2_c_267_n 0.00132475f $X=2.175 $Y=2.465 $X2=0 $Y2=0
cc_184 A3 N_B2_c_267_n 3.8851e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A3_c_230_n N_B2_c_267_n 0.0174225f $X=2.375 $Y=1.46 $X2=0 $Y2=0
cc_186 N_A3_M1007_g N_B2_c_268_n 4.28968e-19 $X=2.175 $Y=2.465 $X2=0 $Y2=0
cc_187 A3 N_B2_c_268_n 0.0339458f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A3_c_230_n N_B2_c_268_n 0.00189044f $X=2.375 $Y=1.46 $X2=0 $Y2=0
cc_189 N_A3_M1007_g N_VPWR_c_366_n 0.00533769f $X=2.175 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A3_M1007_g N_VPWR_c_360_n 0.0103949f $X=2.175 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A3_c_228_n N_VGND_c_413_n 0.00401871f $X=2.375 $Y=1.295 $X2=0 $Y2=0
cc_192 N_A3_c_228_n N_VGND_c_414_n 0.00775088f $X=2.375 $Y=1.295 $X2=0 $Y2=0
cc_193 N_A3_c_228_n N_VGND_c_415_n 0.00948429f $X=2.375 $Y=1.295 $X2=0 $Y2=0
cc_194 N_A3_c_228_n N_A_250_69#_c_460_n 0.0156609f $X=2.375 $Y=1.295 $X2=0 $Y2=0
cc_195 A3 N_A_250_69#_c_460_n 0.0262772f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A3_c_230_n N_A_250_69#_c_460_n 0.00101095f $X=2.375 $Y=1.46 $X2=0 $Y2=0
cc_197 N_A3_c_228_n N_A_250_69#_c_452_n 7.38449e-19 $X=2.375 $Y=1.295 $X2=0
+ $Y2=0
cc_198 N_B2_M1000_g N_B1_c_305_n 0.0152938f $X=2.805 $Y=0.765 $X2=-0.19
+ $Y2=-0.245
cc_199 N_B2_M1002_g N_B1_M1005_g 0.0562145f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_200 N_B2_c_267_n N_B1_c_308_n 0.0562145f $X=2.825 $Y=1.51 $X2=0 $Y2=0
cc_201 N_B2_c_268_n N_B1_c_308_n 3.37791e-19 $X=2.825 $Y=1.51 $X2=0 $Y2=0
cc_202 N_B2_M1002_g N_VPWR_c_363_n 0.00335008f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B2_M1002_g N_VPWR_c_366_n 0.00526178f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B2_M1002_g N_VPWR_c_360_n 0.009938f $X=2.945 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B2_M1000_g N_VGND_c_413_n 0.0029147f $X=2.805 $Y=0.765 $X2=0 $Y2=0
cc_206 N_B2_M1000_g N_VGND_c_414_n 0.00403486f $X=2.805 $Y=0.765 $X2=0 $Y2=0
cc_207 N_B2_M1000_g N_VGND_c_415_n 3.79187e-19 $X=2.805 $Y=0.765 $X2=0 $Y2=0
cc_208 N_B2_c_267_n N_A_250_69#_c_460_n 0.00127925f $X=2.825 $Y=1.51 $X2=0 $Y2=0
cc_209 N_B2_c_268_n N_A_250_69#_c_460_n 0.00904262f $X=2.825 $Y=1.51 $X2=0 $Y2=0
cc_210 N_B2_M1000_g N_A_250_69#_c_451_n 0.012143f $X=2.805 $Y=0.765 $X2=0 $Y2=0
cc_211 N_B2_M1000_g N_A_250_69#_c_452_n 8.15578e-19 $X=2.805 $Y=0.765 $X2=0
+ $Y2=0
cc_212 B1 N_VPWR_M1005_d 0.00790348f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_213 N_B1_M1005_g N_VPWR_c_363_n 0.0229577f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_214 B1 N_VPWR_c_363_n 0.0220472f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_215 N_B1_c_308_n N_VPWR_c_363_n 0.00152745f $X=3.525 $Y=1.46 $X2=0 $Y2=0
cc_216 N_B1_M1005_g N_VPWR_c_366_n 0.00486043f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_217 N_B1_M1005_g N_VPWR_c_360_n 0.00818711f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B1_c_305_n N_VGND_c_413_n 0.0029147f $X=3.305 $Y=1.295 $X2=0 $Y2=0
cc_219 N_B1_c_305_n N_VGND_c_414_n 0.00425623f $X=3.305 $Y=1.295 $X2=0 $Y2=0
cc_220 N_B1_c_305_n N_A_250_69#_c_451_n 0.0130808f $X=3.305 $Y=1.295 $X2=0 $Y2=0
cc_221 B1 N_A_250_69#_c_453_n 0.0246705f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_222 N_B1_c_308_n N_A_250_69#_c_453_n 0.00185801f $X=3.525 $Y=1.46 $X2=0 $Y2=0
cc_223 N_X_c_339_n N_VPWR_c_364_n 0.0335583f $X=0.455 $Y=2.91 $X2=0 $Y2=0
cc_224 N_X_M1009_s N_VPWR_c_360_n 0.00423245f $X=0.33 $Y=1.835 $X2=0 $Y2=0
cc_225 N_X_c_339_n N_VPWR_c_360_n 0.0183839f $X=0.455 $Y=2.91 $X2=0 $Y2=0
cc_226 N_X_c_337_n N_VGND_c_409_n 0.0299267f $X=0.48 $Y=0.49 $X2=0 $Y2=0
cc_227 N_X_c_337_n N_VGND_c_411_n 0.0254358f $X=0.48 $Y=0.49 $X2=0 $Y2=0
cc_228 N_X_c_337_n N_VGND_c_414_n 0.0192268f $X=0.48 $Y=0.49 $X2=0 $Y2=0
cc_229 N_VPWR_c_360_n A_264_367# 0.0137053f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_230 N_VPWR_c_360_n A_358_367# 0.0132771f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_231 N_VPWR_c_360_n A_604_367# 0.00899413f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_232 N_VGND_c_409_n N_A_250_69#_c_450_n 0.0243612f $X=0.935 $Y=0.47 $X2=0
+ $Y2=0
cc_233 N_VGND_c_410_n N_A_250_69#_c_450_n 0.0115876f $X=1.655 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_414_n N_A_250_69#_c_450_n 0.00807296f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_415_n N_A_250_69#_c_450_n 0.0180362f $X=1.68 $Y=0 $X2=0 $Y2=0
cc_236 N_VGND_M1001_d N_A_250_69#_c_460_n 0.016221f $X=1.68 $Y=0.345 $X2=0 $Y2=0
cc_237 N_VGND_c_415_n N_A_250_69#_c_460_n 0.0447396f $X=1.68 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_c_413_n N_A_250_69#_c_451_n 0.0642364f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_239 N_VGND_c_414_n N_A_250_69#_c_451_n 0.0358316f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_c_413_n N_A_250_69#_c_452_n 0.0168464f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_414_n N_A_250_69#_c_452_n 0.00913626f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_242 N_VGND_c_415_n N_A_250_69#_c_452_n 0.0112909f $X=1.68 $Y=0 $X2=0 $Y2=0
