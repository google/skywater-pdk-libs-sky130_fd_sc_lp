* File: sky130_fd_sc_lp__o2111ai_m.pxi.spice
* Created: Fri Aug 28 11:01:28 2020
* 
x_PM_SKY130_FD_SC_LP__O2111AI_M%D1 N_D1_c_72_n N_D1_c_73_n N_D1_c_74_n
+ N_D1_M1002_g N_D1_c_75_n N_D1_M1003_g N_D1_c_76_n N_D1_c_81_n D1 D1 D1 D1
+ N_D1_c_78_n PM_SKY130_FD_SC_LP__O2111AI_M%D1
x_PM_SKY130_FD_SC_LP__O2111AI_M%C1 N_C1_M1009_g N_C1_M1004_g N_C1_c_121_n
+ N_C1_c_124_n N_C1_c_125_n N_C1_c_126_n C1 C1 C1 C1 C1 N_C1_c_123_n
+ PM_SKY130_FD_SC_LP__O2111AI_M%C1
x_PM_SKY130_FD_SC_LP__O2111AI_M%B1 N_B1_M1005_g N_B1_M1006_g N_B1_c_181_n
+ N_B1_c_182_n B1 B1 B1 N_B1_c_179_n PM_SKY130_FD_SC_LP__O2111AI_M%B1
x_PM_SKY130_FD_SC_LP__O2111AI_M%A2 N_A2_M1007_g N_A2_M1001_g N_A2_c_222_n
+ N_A2_c_227_n A2 A2 A2 N_A2_c_224_n PM_SKY130_FD_SC_LP__O2111AI_M%A2
x_PM_SKY130_FD_SC_LP__O2111AI_M%A1 N_A1_M1008_g N_A1_M1000_g N_A1_c_269_n
+ N_A1_c_264_n N_A1_c_265_n A1 A1 A1 A1 N_A1_c_267_n
+ PM_SKY130_FD_SC_LP__O2111AI_M%A1
x_PM_SKY130_FD_SC_LP__O2111AI_M%VPWR N_VPWR_M1002_s N_VPWR_M1009_d
+ N_VPWR_M1008_d N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n
+ N_VPWR_c_304_n N_VPWR_c_305_n VPWR N_VPWR_c_306_n N_VPWR_c_307_n
+ N_VPWR_c_299_n N_VPWR_c_309_n PM_SKY130_FD_SC_LP__O2111AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O2111AI_M%Y N_Y_M1003_s N_Y_M1002_d N_Y_M1006_d
+ N_Y_c_343_n N_Y_c_344_n N_Y_c_346_n Y Y Y N_Y_c_349_n Y
+ PM_SKY130_FD_SC_LP__O2111AI_M%Y
x_PM_SKY130_FD_SC_LP__O2111AI_M%A_357_50# N_A_357_50#_M1005_d
+ N_A_357_50#_M1000_d N_A_357_50#_c_399_n N_A_357_50#_c_400_n
+ N_A_357_50#_c_401_n N_A_357_50#_c_402_n
+ PM_SKY130_FD_SC_LP__O2111AI_M%A_357_50#
x_PM_SKY130_FD_SC_LP__O2111AI_M%VGND N_VGND_M1007_d N_VGND_c_425_n
+ N_VGND_c_426_n N_VGND_c_427_n VGND N_VGND_c_428_n N_VGND_c_429_n
+ PM_SKY130_FD_SC_LP__O2111AI_M%VGND
cc_1 VNB N_D1_c_72_n 0.0114615f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.08
cc_2 VNB N_D1_c_73_n 0.0248401f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.855
cc_3 VNB N_D1_c_74_n 0.0182337f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.855
cc_4 VNB N_D1_c_75_n 0.0198376f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.78
cc_5 VNB N_D1_c_76_n 0.0188187f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.45
cc_6 VNB D1 0.0106325f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_7 VNB N_D1_c_78_n 0.0266412f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.945
cc_8 VNB N_C1_M1004_g 0.0321819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C1_c_121_n 0.0256237f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.93
cc_10 VNB C1 0.00389884f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=2.155
cc_11 VNB N_C1_c_123_n 0.0262822f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.945
cc_12 VNB N_B1_M1005_g 0.051823f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.855
cc_13 VNB B1 0.0106035f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.285
cc_14 VNB N_B1_c_179_n 0.0136116f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_15 VNB N_A2_M1007_g 0.0392157f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.855
cc_16 VNB N_A2_c_222_n 0.0197933f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.46
cc_17 VNB A2 0.00115904f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.285
cc_18 VNB N_A2_c_224_n 0.0170341f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_19 VNB N_A1_M1000_g 0.021924f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=2.885
cc_20 VNB N_A1_c_264_n 0.0220612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_265_n 0.0426653f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_22 VNB A1 0.0193098f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_23 VNB N_A1_c_267_n 0.0125346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_299_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.035
cc_25 VNB N_Y_c_343_n 0.0510671f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.46
cc_26 VNB N_Y_c_344_n 0.0255917f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.155
cc_27 VNB N_A_357_50#_c_399_n 0.00133101f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.78
cc_28 VNB N_A_357_50#_c_400_n 0.0180103f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.46
cc_29 VNB N_A_357_50#_c_401_n 0.00918778f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.93
cc_30 VNB N_A_357_50#_c_402_n 0.00300716f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=2.155
cc_31 VNB N_VGND_c_425_n 0.00533876f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=2.885
cc_32 VNB N_VGND_c_426_n 0.0645149f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.78
cc_33 VNB N_VGND_c_427_n 0.00401228f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=0.46
cc_34 VNB N_VGND_c_428_n 0.0283878f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_35 VNB N_VGND_c_429_n 0.229372f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_36 VPB N_D1_c_72_n 0.0251751f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.08
cc_37 VPB N_D1_M1002_g 0.0383839f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=2.885
cc_38 VPB N_D1_c_81_n 0.0245356f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=2.155
cc_39 VPB D1 0.00850737f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_40 VPB N_C1_c_124_n 0.016875f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.45
cc_41 VPB N_C1_c_125_n 0.0280654f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=2.155
cc_42 VPB N_C1_c_126_n 0.0269947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB C1 0.00276239f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=2.155
cc_44 VPB N_C1_c_123_n 0.00131911f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.945
cc_45 VPB N_B1_M1006_g 0.0334862f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=2.885
cc_46 VPB N_B1_c_181_n 0.023306f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=0.46
cc_47 VPB N_B1_c_182_n 0.0160194f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.93
cc_48 VPB N_B1_c_179_n 0.00272988f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_49 VPB N_A2_M1001_g 0.0464234f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=2.885
cc_50 VPB N_A2_c_222_n 0.00409533f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=0.46
cc_51 VPB N_A2_c_227_n 0.0187231f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.93
cc_52 VPB A2 0.00489505f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.285
cc_53 VPB N_A1_M1008_g 0.040065f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.855
cc_54 VPB N_A1_c_269_n 0.077999f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.45
cc_55 VPB A1 0.0153829f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_56 VPB N_A1_c_267_n 0.0107424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_300_n 0.0142813f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=0.46
cc_58 VPB N_VPWR_c_301_n 0.00485511f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.93
cc_59 VPB N_VPWR_c_302_n 0.00494119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_303_n 0.0126648f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_61 VPB N_VPWR_c_304_n 0.024626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_305_n 0.00401108f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_306_n 0.0250527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_307_n 0.0174178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_299_n 0.0629016f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.035
cc_66 VPB N_VPWR_c_309_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_Y_c_343_n 0.0321979f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=0.46
cc_68 VPB N_Y_c_346_n 0.0106168f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=2.155
cc_69 VPB Y 0.0274458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB Y 0.0131778f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_71 VPB N_Y_c_349_n 0.0135773f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=0.945
cc_72 N_D1_c_75_n N_C1_M1004_g 0.0505824f $X=0.99 $Y=0.78 $X2=0 $Y2=0
cc_73 D1 N_C1_M1004_g 6.8772e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_74 N_D1_c_78_n N_C1_M1004_g 0.00362761f $X=0.58 $Y=0.945 $X2=0 $Y2=0
cc_75 N_D1_c_73_n N_C1_c_121_n 0.00667458f $X=0.915 $Y=0.855 $X2=0 $Y2=0
cc_76 D1 N_C1_c_121_n 0.00496107f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_77 N_D1_c_78_n N_C1_c_121_n 0.0123075f $X=0.58 $Y=0.945 $X2=0 $Y2=0
cc_78 N_D1_c_72_n N_C1_c_124_n 0.0123075f $X=0.67 $Y=2.08 $X2=0 $Y2=0
cc_79 N_D1_c_72_n N_C1_c_125_n 0.00686479f $X=0.67 $Y=2.08 $X2=0 $Y2=0
cc_80 N_D1_c_81_n N_C1_c_125_n 0.0157653f $X=0.85 $Y=2.155 $X2=0 $Y2=0
cc_81 D1 N_C1_c_125_n 8.75728e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_82 N_D1_M1002_g N_C1_c_126_n 0.0309382f $X=0.85 $Y=2.885 $X2=0 $Y2=0
cc_83 N_D1_c_72_n C1 8.04522e-19 $X=0.67 $Y=2.08 $X2=0 $Y2=0
cc_84 N_D1_c_75_n C1 0.00504103f $X=0.99 $Y=0.78 $X2=0 $Y2=0
cc_85 N_D1_c_81_n C1 2.76198e-19 $X=0.85 $Y=2.155 $X2=0 $Y2=0
cc_86 D1 C1 0.0764462f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_87 N_D1_c_78_n C1 0.00147148f $X=0.58 $Y=0.945 $X2=0 $Y2=0
cc_88 N_D1_c_76_n N_C1_c_123_n 0.0123075f $X=0.58 $Y=1.45 $X2=0 $Y2=0
cc_89 N_D1_M1002_g N_VPWR_c_301_n 0.00690632f $X=0.85 $Y=2.885 $X2=0 $Y2=0
cc_90 N_D1_M1002_g N_VPWR_c_304_n 0.00375793f $X=0.85 $Y=2.885 $X2=0 $Y2=0
cc_91 N_D1_M1002_g N_VPWR_c_299_n 0.00689964f $X=0.85 $Y=2.885 $X2=0 $Y2=0
cc_92 N_D1_c_72_n N_Y_c_343_n 0.00367353f $X=0.67 $Y=2.08 $X2=0 $Y2=0
cc_93 N_D1_c_74_n N_Y_c_343_n 0.0169123f $X=0.745 $Y=0.855 $X2=0 $Y2=0
cc_94 N_D1_M1002_g N_Y_c_343_n 0.00224546f $X=0.85 $Y=2.885 $X2=0 $Y2=0
cc_95 N_D1_c_75_n N_Y_c_343_n 0.00393299f $X=0.99 $Y=0.78 $X2=0 $Y2=0
cc_96 N_D1_c_81_n N_Y_c_343_n 0.00367332f $X=0.85 $Y=2.155 $X2=0 $Y2=0
cc_97 D1 N_Y_c_343_n 0.0986931f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_98 N_D1_c_74_n N_Y_c_344_n 0.00532783f $X=0.745 $Y=0.855 $X2=0 $Y2=0
cc_99 N_D1_c_75_n N_Y_c_344_n 0.010835f $X=0.99 $Y=0.78 $X2=0 $Y2=0
cc_100 D1 N_Y_c_344_n 0.0189367f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_101 N_D1_M1002_g Y 0.0327939f $X=0.85 $Y=2.885 $X2=0 $Y2=0
cc_102 N_D1_c_81_n Y 0.00516985f $X=0.85 $Y=2.155 $X2=0 $Y2=0
cc_103 D1 Y 0.0233645f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_104 N_D1_c_73_n N_VGND_c_426_n 0.00222659f $X=0.915 $Y=0.855 $X2=0 $Y2=0
cc_105 N_D1_c_75_n N_VGND_c_426_n 0.00570116f $X=0.99 $Y=0.78 $X2=0 $Y2=0
cc_106 N_D1_c_73_n N_VGND_c_429_n 0.00233389f $X=0.915 $Y=0.855 $X2=0 $Y2=0
cc_107 N_D1_c_75_n N_VGND_c_429_n 0.0119156f $X=0.99 $Y=0.78 $X2=0 $Y2=0
cc_108 D1 N_VGND_c_429_n 0.00263639f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_109 N_C1_M1004_g N_B1_M1005_g 0.0721357f $X=1.35 $Y=0.46 $X2=0 $Y2=0
cc_110 C1 N_B1_M1005_g 0.00299884f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_111 N_C1_c_123_n N_B1_M1005_g 0.00862156f $X=1.15 $Y=1.335 $X2=0 $Y2=0
cc_112 N_C1_c_125_n N_B1_M1006_g 0.00797157f $X=1.245 $Y=2.41 $X2=0 $Y2=0
cc_113 N_C1_c_126_n N_B1_M1006_g 0.0224409f $X=1.245 $Y=2.56 $X2=0 $Y2=0
cc_114 N_C1_c_124_n N_B1_c_181_n 0.00946567f $X=1.15 $Y=1.84 $X2=0 $Y2=0
cc_115 N_C1_c_125_n N_B1_c_181_n 0.0185999f $X=1.245 $Y=2.41 $X2=0 $Y2=0
cc_116 N_C1_c_121_n B1 6.25096e-19 $X=1.205 $Y=1.29 $X2=0 $Y2=0
cc_117 N_C1_c_125_n B1 8.87589e-19 $X=1.245 $Y=2.41 $X2=0 $Y2=0
cc_118 C1 B1 0.0514933f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_119 N_C1_c_123_n B1 0.00287473f $X=1.15 $Y=1.335 $X2=0 $Y2=0
cc_120 C1 N_B1_c_179_n 0.00206011f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_121 N_C1_c_123_n N_B1_c_179_n 0.00946567f $X=1.15 $Y=1.335 $X2=0 $Y2=0
cc_122 N_C1_c_126_n N_VPWR_c_302_n 0.00288714f $X=1.245 $Y=2.56 $X2=0 $Y2=0
cc_123 N_C1_c_126_n N_VPWR_c_304_n 0.00435108f $X=1.245 $Y=2.56 $X2=0 $Y2=0
cc_124 N_C1_c_126_n N_VPWR_c_299_n 0.00599853f $X=1.245 $Y=2.56 $X2=0 $Y2=0
cc_125 N_C1_c_124_n Y 0.00308999f $X=1.15 $Y=1.84 $X2=0 $Y2=0
cc_126 N_C1_c_125_n Y 0.0018761f $X=1.245 $Y=2.41 $X2=0 $Y2=0
cc_127 N_C1_c_126_n Y 0.00399346f $X=1.245 $Y=2.56 $X2=0 $Y2=0
cc_128 C1 Y 0.00826963f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_129 N_C1_c_124_n N_Y_c_349_n 5.8207e-19 $X=1.15 $Y=1.84 $X2=0 $Y2=0
cc_130 N_C1_c_125_n N_Y_c_349_n 0.00417383f $X=1.245 $Y=2.41 $X2=0 $Y2=0
cc_131 N_C1_c_126_n N_Y_c_349_n 0.0119205f $X=1.245 $Y=2.56 $X2=0 $Y2=0
cc_132 C1 N_Y_c_349_n 0.0079389f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_133 C1 A_213_50# 0.00139886f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_134 C1 N_A_357_50#_c_399_n 0.00489879f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_135 C1 N_A_357_50#_c_401_n 0.0058747f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_136 N_C1_M1004_g N_VGND_c_426_n 0.00559135f $X=1.35 $Y=0.46 $X2=0 $Y2=0
cc_137 C1 N_VGND_c_426_n 0.00477283f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_138 N_C1_M1004_g N_VGND_c_429_n 0.0101967f $X=1.35 $Y=0.46 $X2=0 $Y2=0
cc_139 C1 N_VGND_c_429_n 0.007402f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_140 N_B1_M1005_g N_A2_M1007_g 0.048454f $X=1.71 $Y=0.46 $X2=0 $Y2=0
cc_141 N_B1_M1006_g N_A2_M1001_g 0.032997f $X=1.71 $Y=2.885 $X2=0 $Y2=0
cc_142 N_B1_c_182_n N_A2_M1001_g 0.0135626f $X=1.69 $Y=2.2 $X2=0 $Y2=0
cc_143 B1 N_A2_c_222_n 0.00195213f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_B1_c_179_n N_A2_c_222_n 0.0135626f $X=1.69 $Y=1.695 $X2=0 $Y2=0
cc_145 N_B1_c_181_n N_A2_c_227_n 0.0135626f $X=1.69 $Y=2.035 $X2=0 $Y2=0
cc_146 N_B1_M1005_g A2 3.63816e-19 $X=1.71 $Y=0.46 $X2=0 $Y2=0
cc_147 B1 A2 0.0554443f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_148 N_B1_c_179_n A2 0.00202068f $X=1.69 $Y=1.695 $X2=0 $Y2=0
cc_149 B1 N_A2_c_224_n 0.00213788f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_150 N_B1_M1006_g N_VPWR_c_302_n 0.00288714f $X=1.71 $Y=2.885 $X2=0 $Y2=0
cc_151 N_B1_M1006_g N_VPWR_c_306_n 0.00435108f $X=1.71 $Y=2.885 $X2=0 $Y2=0
cc_152 N_B1_M1006_g N_VPWR_c_299_n 0.00599853f $X=1.71 $Y=2.885 $X2=0 $Y2=0
cc_153 N_B1_M1006_g Y 0.00153267f $X=1.71 $Y=2.885 $X2=0 $Y2=0
cc_154 N_B1_c_182_n Y 0.00100459f $X=1.69 $Y=2.2 $X2=0 $Y2=0
cc_155 B1 Y 0.00259002f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B1_M1006_g N_Y_c_349_n 0.0152561f $X=1.71 $Y=2.885 $X2=0 $Y2=0
cc_157 N_B1_c_182_n N_Y_c_349_n 0.00412199f $X=1.69 $Y=2.2 $X2=0 $Y2=0
cc_158 B1 N_Y_c_349_n 0.0210678f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_159 N_B1_M1005_g N_A_357_50#_c_399_n 8.59822e-19 $X=1.71 $Y=0.46 $X2=0 $Y2=0
cc_160 N_B1_M1005_g N_A_357_50#_c_401_n 0.0025826f $X=1.71 $Y=0.46 $X2=0 $Y2=0
cc_161 B1 N_A_357_50#_c_401_n 0.00210798f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B1_M1005_g N_VGND_c_426_n 0.00570116f $X=1.71 $Y=0.46 $X2=0 $Y2=0
cc_163 N_B1_M1005_g N_VGND_c_429_n 0.0106903f $X=1.71 $Y=0.46 $X2=0 $Y2=0
cc_164 N_A2_M1007_g N_A1_M1000_g 0.0235637f $X=2.14 $Y=0.46 $X2=0 $Y2=0
cc_165 N_A2_M1001_g N_A1_c_269_n 0.0745228f $X=2.14 $Y=2.885 $X2=0 $Y2=0
cc_166 N_A2_c_227_n N_A1_c_269_n 0.0116837f $X=2.23 $Y=1.88 $X2=0 $Y2=0
cc_167 A2 N_A1_c_269_n 7.8118e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_168 N_A2_M1007_g N_A1_c_265_n 0.00840749f $X=2.14 $Y=0.46 $X2=0 $Y2=0
cc_169 A2 N_A1_c_265_n 6.66405e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A2_c_224_n N_A1_c_265_n 0.0116837f $X=2.23 $Y=1.375 $X2=0 $Y2=0
cc_171 N_A2_M1001_g A1 0.00195666f $X=2.14 $Y=2.885 $X2=0 $Y2=0
cc_172 A2 A1 0.0553677f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A2_c_224_n A1 0.00476259f $X=2.23 $Y=1.375 $X2=0 $Y2=0
cc_174 N_A2_c_222_n N_A1_c_267_n 0.0116837f $X=2.23 $Y=1.715 $X2=0 $Y2=0
cc_175 N_A2_M1001_g N_VPWR_c_303_n 0.0019051f $X=2.14 $Y=2.885 $X2=0 $Y2=0
cc_176 N_A2_M1001_g N_VPWR_c_306_n 0.0037962f $X=2.14 $Y=2.885 $X2=0 $Y2=0
cc_177 N_A2_M1001_g N_VPWR_c_299_n 0.00535384f $X=2.14 $Y=2.885 $X2=0 $Y2=0
cc_178 N_A2_M1001_g Y 0.0185143f $X=2.14 $Y=2.885 $X2=0 $Y2=0
cc_179 A2 Y 0.012686f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A2_M1001_g N_Y_c_349_n 2.28537e-19 $X=2.14 $Y=2.885 $X2=0 $Y2=0
cc_181 N_A2_M1007_g N_A_357_50#_c_399_n 9.4709e-19 $X=2.14 $Y=0.46 $X2=0 $Y2=0
cc_182 N_A2_M1007_g N_A_357_50#_c_400_n 0.0128333f $X=2.14 $Y=0.46 $X2=0 $Y2=0
cc_183 A2 N_A_357_50#_c_400_n 0.0118697f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A2_c_224_n N_A_357_50#_c_400_n 0.00351131f $X=2.23 $Y=1.375 $X2=0 $Y2=0
cc_185 N_A2_M1007_g N_VGND_c_425_n 0.00280554f $X=2.14 $Y=0.46 $X2=0 $Y2=0
cc_186 N_A2_M1007_g N_VGND_c_426_n 0.00426948f $X=2.14 $Y=0.46 $X2=0 $Y2=0
cc_187 N_A2_M1007_g N_VGND_c_429_n 0.00599235f $X=2.14 $Y=0.46 $X2=0 $Y2=0
cc_188 N_A1_M1008_g N_VPWR_c_303_n 0.010326f $X=2.5 $Y=2.885 $X2=0 $Y2=0
cc_189 N_A1_c_269_n N_VPWR_c_303_n 0.00127879f $X=2.8 $Y=2.12 $X2=0 $Y2=0
cc_190 A1 N_VPWR_c_303_n 0.013632f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_191 N_A1_M1008_g N_VPWR_c_306_n 0.00486043f $X=2.5 $Y=2.885 $X2=0 $Y2=0
cc_192 N_A1_M1008_g N_VPWR_c_299_n 0.00818711f $X=2.5 $Y=2.885 $X2=0 $Y2=0
cc_193 A1 N_VPWR_c_299_n 0.00194381f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A1_M1008_g Y 0.00629968f $X=2.5 $Y=2.885 $X2=0 $Y2=0
cc_195 A1 Y 0.00878512f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A1_M1000_g N_A_357_50#_c_400_n 0.00735288f $X=2.57 $Y=0.46 $X2=0 $Y2=0
cc_197 N_A1_c_264_n N_A_357_50#_c_400_n 0.0137094f $X=2.71 $Y=0.895 $X2=0 $Y2=0
cc_198 A1 N_A_357_50#_c_400_n 0.0180004f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_199 N_A1_c_267_n N_A_357_50#_c_400_n 5.18908e-19 $X=2.8 $Y=1.765 $X2=0 $Y2=0
cc_200 N_A1_M1000_g N_A_357_50#_c_402_n 0.0020107f $X=2.57 $Y=0.46 $X2=0 $Y2=0
cc_201 N_A1_M1000_g N_VGND_c_425_n 0.00280554f $X=2.57 $Y=0.46 $X2=0 $Y2=0
cc_202 N_A1_M1000_g N_VGND_c_428_n 0.00426948f $X=2.57 $Y=0.46 $X2=0 $Y2=0
cc_203 N_A1_M1000_g N_VGND_c_429_n 0.00704947f $X=2.57 $Y=0.46 $X2=0 $Y2=0
cc_204 N_VPWR_c_299_n N_Y_M1002_d 0.00247873f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_c_299_n N_Y_M1006_d 0.00251033f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_206 N_VPWR_c_301_n N_Y_c_346_n 0.00271309f $X=0.37 $Y=2.95 $X2=0 $Y2=0
cc_207 N_VPWR_c_299_n N_Y_c_346_n 0.00498685f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_208 N_VPWR_M1002_s Y 0.00804398f $X=0.245 $Y=2.675 $X2=0 $Y2=0
cc_209 N_VPWR_c_301_n Y 0.0223766f $X=0.37 $Y=2.95 $X2=0 $Y2=0
cc_210 N_VPWR_c_304_n Y 0.0204774f $X=1.39 $Y=3.33 $X2=0 $Y2=0
cc_211 N_VPWR_c_299_n Y 0.025825f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_306_n Y 0.0149241f $X=2.55 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_299_n Y 0.0147121f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_c_302_n N_Y_c_349_n 0.0145132f $X=1.495 $Y=2.97 $X2=0 $Y2=0
cc_215 N_VPWR_c_304_n N_Y_c_349_n 0.00332233f $X=1.39 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_306_n N_Y_c_349_n 0.00332233f $X=2.55 $Y=3.33 $X2=0 $Y2=0
cc_217 N_VPWR_c_299_n N_Y_c_349_n 0.0114916f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_218 N_VPWR_c_299_n A_443_535# 0.0079978f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_219 N_Y_c_344_n N_VGND_c_426_n 0.0367543f $X=0.64 $Y=0.435 $X2=0 $Y2=0
cc_220 N_Y_c_344_n N_VGND_c_429_n 0.0227079f $X=0.64 $Y=0.435 $X2=0 $Y2=0
cc_221 N_A_357_50#_c_400_n N_VGND_c_425_n 0.0140142f $X=2.68 $Y=0.825 $X2=0
+ $Y2=0
cc_222 N_A_357_50#_c_399_n N_VGND_c_426_n 0.00775159f $X=1.925 $Y=0.525 $X2=0
+ $Y2=0
cc_223 N_A_357_50#_c_400_n N_VGND_c_426_n 0.00296079f $X=2.68 $Y=0.825 $X2=0
+ $Y2=0
cc_224 N_A_357_50#_c_400_n N_VGND_c_428_n 0.00296079f $X=2.68 $Y=0.825 $X2=0
+ $Y2=0
cc_225 N_A_357_50#_c_402_n N_VGND_c_428_n 0.00815096f $X=2.785 $Y=0.525 $X2=0
+ $Y2=0
cc_226 N_A_357_50#_c_399_n N_VGND_c_429_n 0.00758036f $X=1.925 $Y=0.525 $X2=0
+ $Y2=0
cc_227 N_A_357_50#_c_400_n N_VGND_c_429_n 0.0109527f $X=2.68 $Y=0.825 $X2=0
+ $Y2=0
cc_228 N_A_357_50#_c_402_n N_VGND_c_429_n 0.00758036f $X=2.785 $Y=0.525 $X2=0
+ $Y2=0
