* File: sky130_fd_sc_lp__mux2_4.pxi.spice
* Created: Fri Aug 28 10:44:04 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2_4%S N_S_c_101_n N_S_M1013_g N_S_c_102_n N_S_M1007_g
+ N_S_c_103_n N_S_M1004_g N_S_M1009_g N_S_c_110_n N_S_c_111_n N_S_c_112_n S S
+ N_S_c_106_n N_S_c_114_n S PM_SKY130_FD_SC_LP__MUX2_4%S
x_PM_SKY130_FD_SC_LP__MUX2_4%A_41_367# N_A_41_367#_M1007_s N_A_41_367#_M1013_s
+ N_A_41_367#_c_202_n N_A_41_367#_M1017_g N_A_41_367#_M1008_g
+ N_A_41_367#_c_196_n N_A_41_367#_c_203_n N_A_41_367#_c_197_n
+ N_A_41_367#_c_198_n N_A_41_367#_c_199_n N_A_41_367#_c_200_n
+ N_A_41_367#_c_205_n N_A_41_367#_c_201_n PM_SKY130_FD_SC_LP__MUX2_4%A_41_367#
x_PM_SKY130_FD_SC_LP__MUX2_4%A0 N_A0_c_251_n N_A0_M1010_g N_A0_M1005_g A0 A0 A0
+ N_A0_c_254_n PM_SKY130_FD_SC_LP__MUX2_4%A0
x_PM_SKY130_FD_SC_LP__MUX2_4%A1 N_A1_M1002_g N_A1_M1011_g A1 A1 N_A1_c_294_n
+ N_A1_c_295_n PM_SKY130_FD_SC_LP__MUX2_4%A1
x_PM_SKY130_FD_SC_LP__MUX2_4%A_359_47# N_A_359_47#_M1010_d N_A_359_47#_M1005_d
+ N_A_359_47#_M1000_g N_A_359_47#_M1003_g N_A_359_47#_M1001_g
+ N_A_359_47#_M1006_g N_A_359_47#_M1014_g N_A_359_47#_M1012_g
+ N_A_359_47#_M1015_g N_A_359_47#_M1016_g N_A_359_47#_c_351_n
+ N_A_359_47#_c_343_n N_A_359_47#_c_355_n N_A_359_47#_c_373_n
+ N_A_359_47#_c_334_n N_A_359_47#_c_335_n N_A_359_47#_c_336_n
+ N_A_359_47#_c_337_n N_A_359_47#_c_367_n N_A_359_47#_c_338_n
+ PM_SKY130_FD_SC_LP__MUX2_4%A_359_47#
x_PM_SKY130_FD_SC_LP__MUX2_4%VPWR N_VPWR_M1013_d N_VPWR_M1009_d N_VPWR_M1006_s
+ N_VPWR_M1016_s N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_470_n
+ N_VPWR_c_471_n N_VPWR_c_472_n N_VPWR_c_473_n N_VPWR_c_474_n VPWR
+ N_VPWR_c_475_n N_VPWR_c_476_n N_VPWR_c_477_n N_VPWR_c_466_n N_VPWR_c_479_n
+ N_VPWR_c_480_n PM_SKY130_FD_SC_LP__MUX2_4%VPWR
x_PM_SKY130_FD_SC_LP__MUX2_4%A_210_367# N_A_210_367#_M1017_d
+ N_A_210_367#_M1002_d N_A_210_367#_c_543_n N_A_210_367#_c_544_n
+ N_A_210_367#_c_545_n N_A_210_367#_c_546_n
+ PM_SKY130_FD_SC_LP__MUX2_4%A_210_367#
x_PM_SKY130_FD_SC_LP__MUX2_4%A_317_367# N_A_317_367#_M1005_s
+ N_A_317_367#_M1009_s N_A_317_367#_c_572_n N_A_317_367#_c_573_n
+ N_A_317_367#_c_574_n N_A_317_367#_c_575_n
+ PM_SKY130_FD_SC_LP__MUX2_4%A_317_367#
x_PM_SKY130_FD_SC_LP__MUX2_4%X N_X_M1000_s N_X_M1014_s N_X_M1003_d N_X_M1012_d
+ N_X_c_661_p N_X_c_647_n N_X_c_602_n N_X_c_603_n N_X_c_609_n N_X_c_610_n
+ N_X_c_658_p N_X_c_651_n N_X_c_604_n N_X_c_611_n N_X_c_605_n N_X_c_606_n
+ N_X_c_613_n N_X_c_607_n X X PM_SKY130_FD_SC_LP__MUX2_4%X
x_PM_SKY130_FD_SC_LP__MUX2_4%VGND N_VGND_M1007_d N_VGND_M1004_d N_VGND_M1001_d
+ N_VGND_M1015_d N_VGND_c_668_n N_VGND_c_669_n N_VGND_c_670_n N_VGND_c_671_n
+ N_VGND_c_672_n N_VGND_c_673_n VGND N_VGND_c_674_n N_VGND_c_675_n
+ N_VGND_c_676_n N_VGND_c_677_n N_VGND_c_678_n N_VGND_c_679_n N_VGND_c_680_n
+ PM_SKY130_FD_SC_LP__MUX2_4%VGND
cc_1 VNB N_S_c_101_n 0.0553896f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.665
cc_2 VNB N_S_c_102_n 0.0211359f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.185
cc_3 VNB N_S_c_103_n 0.0183752f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=1.185
cc_4 VNB N_S_M1009_g 0.00843967f $X=-0.19 $Y=-0.245 $X2=3.305 $Y2=2.465
cc_5 VNB S 0.00313482f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.21
cc_6 VNB N_S_c_106_n 0.0559523f $X=-0.19 $Y=-0.245 $X2=3.07 $Y2=1.35
cc_7 VNB N_A_41_367#_M1008_g 0.0200101f $X=-0.19 $Y=-0.245 $X2=3.305 $Y2=2.465
cc_8 VNB N_A_41_367#_c_196_n 0.0419242f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.5
cc_9 VNB N_A_41_367#_c_197_n 0.00253996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_41_367#_c_198_n 0.00116838f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=1.35
cc_11 VNB N_A_41_367#_c_199_n 0.0431341f $X=-0.19 $Y=-0.245 $X2=3.07 $Y2=1.35
cc_12 VNB N_A_41_367#_c_200_n 0.0159702f $X=-0.19 $Y=-0.245 $X2=3.07 $Y2=1.35
cc_13 VNB N_A_41_367#_c_201_n 0.0234793f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.295
cc_14 VNB N_A0_c_251_n 0.0168132f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.665
cc_15 VNB N_A0_M1005_g 0.00814441f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.655
cc_16 VNB A0 0.00669262f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=1.185
cc_17 VNB N_A0_c_254_n 0.035532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1002_g 0.00869358f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_19 VNB A1 0.0118191f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=0.655
cc_20 VNB N_A1_c_294_n 0.0281524f $X=-0.19 $Y=-0.245 $X2=3.305 $Y2=2.465
cc_21 VNB N_A1_c_295_n 0.0182444f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.695
cc_22 VNB N_A_359_47#_M1000_g 0.0255228f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=0.655
cc_23 VNB N_A_359_47#_M1001_g 0.0222563f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.5
cc_24 VNB N_A_359_47#_M1014_g 0.0222627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_359_47#_M1015_g 0.0284456f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.695
cc_26 VNB N_A_359_47#_c_334_n 0.00281505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_359_47#_c_335_n 4.00689e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_359_47#_c_336_n 0.00170445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_359_47#_c_337_n 0.083014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_359_47#_c_338_n 0.0010634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_466_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_602_n 0.00304705f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.58
cc_33 VNB N_X_c_603_n 0.00292895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_604_n 0.00960778f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.637
cc_35 VNB N_X_c_605_n 0.0214627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_606_n 0.00177181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_607_n 0.00865274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB X 0.0366274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_668_n 7.65996e-19 $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.695
cc_40 VNB N_VGND_c_669_n 3.18577e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_670_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.78
cc_42 VNB N_VGND_c_671_n 0.0043908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_672_n 0.0133822f $X=-0.19 $Y=-0.245 $X2=0.617 $Y2=1.5
cc_44 VNB N_VGND_c_673_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.825 $Y2=1.35
cc_45 VNB N_VGND_c_674_n 0.0230618f $X=-0.19 $Y=-0.245 $X2=3.07 $Y2=1.35
cc_46 VNB N_VGND_c_675_n 0.0162846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_676_n 0.2988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_677_n 0.00642167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_678_n 0.0401645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_679_n 0.0137706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_680_n 0.00432782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VPB N_S_c_101_n 0.00605561f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.665
cc_53 VPB N_S_M1013_g 0.0228083f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_54 VPB N_S_M1009_g 0.0244412f $X=-0.19 $Y=1.655 $X2=3.305 $Y2=2.465
cc_55 VPB N_S_c_110_n 5.70274e-19 $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.5
cc_56 VPB N_S_c_111_n 0.0290118f $X=-0.19 $Y=1.655 $X2=2.905 $Y2=1.78
cc_57 VPB N_S_c_112_n 0.00130528f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.78
cc_58 VPB S 5.34441e-19 $X=-0.19 $Y=1.655 $X2=3.035 $Y2=1.21
cc_59 VPB N_S_c_114_n 0.00137123f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=1.695
cc_60 VPB N_A_41_367#_c_202_n 0.0193752f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.655
cc_61 VPB N_A_41_367#_c_203_n 0.0370647f $X=-0.19 $Y=1.655 $X2=3.035 $Y2=1.21
cc_62 VPB N_A_41_367#_c_199_n 0.0176542f $X=-0.19 $Y=1.655 $X2=3.07 $Y2=1.35
cc_63 VPB N_A_41_367#_c_205_n 0.00693948f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=1.695
cc_64 VPB N_A_41_367#_c_201_n 0.0163286f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=1.295
cc_65 VPB N_A0_M1005_g 0.0234666f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.655
cc_66 VPB N_A1_M1002_g 0.0239037f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_67 VPB N_A_359_47#_M1003_g 0.0192683f $X=-0.19 $Y=1.655 $X2=3.305 $Y2=2.465
cc_68 VPB N_A_359_47#_M1006_g 0.0183494f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.78
cc_69 VPB N_A_359_47#_M1012_g 0.0183546f $X=-0.19 $Y=1.655 $X2=3.07 $Y2=1.35
cc_70 VPB N_A_359_47#_M1016_g 0.0222269f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=1.637
cc_71 VPB N_A_359_47#_c_343_n 0.00679109f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_359_47#_c_335_n 0.00235585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_359_47#_c_337_n 0.016032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_467_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.695
cc_75 VPB N_VPWR_c_468_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.78
cc_76 VPB N_VPWR_c_469_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_470_n 0.0415892f $X=-0.19 $Y=1.655 $X2=3.07 $Y2=1.35
cc_78 VPB N_VPWR_c_471_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_472_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=1.637
cc_80 VPB N_VPWR_c_473_n 0.0130339f $X=-0.19 $Y=1.655 $X2=3.12 $Y2=1.665
cc_81 VPB N_VPWR_c_474_n 0.00510842f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=1.78
cc_82 VPB N_VPWR_c_475_n 0.0168978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_476_n 0.0562379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_477_n 0.0134401f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_466_n 0.0613816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_479_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_480_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_210_367#_c_543_n 0.00898706f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=0.655
cc_89 VPB N_A_210_367#_c_544_n 5.42696e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_210_367#_c_545_n 0.0027126f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.5
cc_91 VPB N_A_210_367#_c_546_n 0.00991302f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.5
cc_92 VPB N_A_317_367#_c_572_n 0.00454007f $X=-0.19 $Y=1.655 $X2=2.825 $Y2=0.655
cc_93 VPB N_A_317_367#_c_573_n 0.00681061f $X=-0.19 $Y=1.655 $X2=3.305 $Y2=1.515
cc_94 VPB N_A_317_367#_c_574_n 0.00239611f $X=-0.19 $Y=1.655 $X2=3.305 $Y2=2.465
cc_95 VPB N_A_317_367#_c_575_n 0.00725438f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.5
cc_96 VPB N_X_c_609_n 0.00304538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_X_c_610_n 0.0020802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_X_c_611_n 0.0231306f $X=-0.19 $Y=1.655 $X2=3.12 $Y2=1.665
cc_99 VPB N_X_c_605_n 0.00531654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_X_c_613_n 0.00134754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 N_S_c_111_n N_A_41_367#_c_202_n 0.0127841f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_102 N_S_c_102_n N_A_41_367#_M1008_g 0.0315361f $X=0.8 $Y=1.185 $X2=0 $Y2=0
cc_103 N_S_c_101_n N_A_41_367#_c_197_n 6.81252e-19 $X=0.545 $Y=1.665 $X2=0 $Y2=0
cc_104 N_S_c_102_n N_A_41_367#_c_197_n 0.0159639f $X=0.8 $Y=1.185 $X2=0 $Y2=0
cc_105 N_S_c_111_n N_A_41_367#_c_197_n 0.0116973f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_106 N_S_c_101_n N_A_41_367#_c_198_n 0.00132042f $X=0.545 $Y=1.665 $X2=0 $Y2=0
cc_107 N_S_c_102_n N_A_41_367#_c_198_n 0.00269174f $X=0.8 $Y=1.185 $X2=0 $Y2=0
cc_108 N_S_c_110_n N_A_41_367#_c_198_n 0.00710109f $X=0.525 $Y=1.5 $X2=0 $Y2=0
cc_109 N_S_c_111_n N_A_41_367#_c_198_n 0.0245092f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_110 N_S_c_101_n N_A_41_367#_c_199_n 0.0183286f $X=0.545 $Y=1.665 $X2=0 $Y2=0
cc_111 N_S_M1013_g N_A_41_367#_c_199_n 0.0199271f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_112 N_S_c_110_n N_A_41_367#_c_199_n 0.00245993f $X=0.525 $Y=1.5 $X2=0 $Y2=0
cc_113 N_S_c_111_n N_A_41_367#_c_199_n 0.0174893f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_114 N_S_c_101_n N_A_41_367#_c_200_n 0.0122935f $X=0.545 $Y=1.665 $X2=0 $Y2=0
cc_115 N_S_c_110_n N_A_41_367#_c_200_n 0.0216315f $X=0.525 $Y=1.5 $X2=0 $Y2=0
cc_116 N_S_c_111_n N_A_41_367#_c_200_n 3.57946e-19 $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_117 N_S_c_101_n N_A_41_367#_c_205_n 0.00217836f $X=0.545 $Y=1.665 $X2=0 $Y2=0
cc_118 N_S_c_101_n N_A_41_367#_c_201_n 0.0136097f $X=0.545 $Y=1.665 $X2=0 $Y2=0
cc_119 N_S_M1013_g N_A_41_367#_c_201_n 0.00522086f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_120 N_S_c_110_n N_A_41_367#_c_201_n 0.026649f $X=0.525 $Y=1.5 $X2=0 $Y2=0
cc_121 N_S_c_112_n N_A_41_367#_c_201_n 0.0128704f $X=0.69 $Y=1.78 $X2=0 $Y2=0
cc_122 N_S_c_111_n N_A0_M1005_g 0.0167596f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_123 N_S_c_111_n A0 0.0264079f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_124 N_S_c_111_n N_A0_c_254_n 0.00138973f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_125 N_S_c_111_n N_A1_M1002_g 0.0124865f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_126 S N_A1_M1002_g 0.00465606f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_127 N_S_c_111_n A1 0.0502907f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_128 S A1 0.0261322f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_129 N_S_c_106_n A1 0.00279768f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_130 N_S_c_111_n N_A1_c_294_n 0.00122433f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_131 S N_A1_c_294_n 2.23674e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_132 N_S_c_106_n N_A1_c_294_n 0.0435327f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_133 N_S_c_103_n N_A1_c_295_n 0.0435327f $X=2.825 $Y=1.185 $X2=0 $Y2=0
cc_134 N_S_c_111_n N_A_359_47#_M1005_d 0.00176891f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_135 N_S_c_103_n N_A_359_47#_M1000_g 0.00869442f $X=2.825 $Y=1.185 $X2=0 $Y2=0
cc_136 S N_A_359_47#_M1000_g 4.22911e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_137 N_S_c_106_n N_A_359_47#_M1000_g 0.00592825f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_138 N_S_M1009_g N_A_359_47#_M1003_g 0.0328136f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_139 N_S_c_103_n N_A_359_47#_c_351_n 0.00252433f $X=2.825 $Y=1.185 $X2=0 $Y2=0
cc_140 N_S_M1009_g N_A_359_47#_c_343_n 0.0202837f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_141 N_S_c_106_n N_A_359_47#_c_343_n 0.00121958f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_142 N_S_c_114_n N_A_359_47#_c_343_n 0.023855f $X=3.08 $Y=1.695 $X2=0 $Y2=0
cc_143 N_S_c_103_n N_A_359_47#_c_355_n 0.0145795f $X=2.825 $Y=1.185 $X2=0 $Y2=0
cc_144 N_S_c_111_n N_A_359_47#_c_355_n 0.00419173f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_145 S N_A_359_47#_c_355_n 0.0255284f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_146 N_S_c_106_n N_A_359_47#_c_355_n 0.0120075f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_147 N_S_c_103_n N_A_359_47#_c_334_n 0.00243731f $X=2.825 $Y=1.185 $X2=0 $Y2=0
cc_148 S N_A_359_47#_c_334_n 0.0161222f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_149 N_S_c_106_n N_A_359_47#_c_334_n 0.00115354f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_150 N_S_M1009_g N_A_359_47#_c_335_n 0.0026042f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_151 S N_A_359_47#_c_335_n 0.00840631f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_152 N_S_c_114_n N_A_359_47#_c_335_n 0.0126411f $X=3.08 $Y=1.695 $X2=0 $Y2=0
cc_153 S N_A_359_47#_c_337_n 2.29508e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_154 N_S_c_106_n N_A_359_47#_c_337_n 0.0185262f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_155 N_S_c_111_n N_A_359_47#_c_367_n 0.0555546f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_156 S N_A_359_47#_c_338_n 0.015201f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_157 N_S_c_106_n N_A_359_47#_c_338_n 0.00144735f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_158 N_S_c_111_n N_VPWR_M1013_d 0.00161579f $X=2.905 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_159 N_S_c_101_n N_VPWR_c_467_n 2.2435e-19 $X=0.545 $Y=1.665 $X2=0 $Y2=0
cc_160 N_S_M1013_g N_VPWR_c_467_n 0.0173896f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_161 N_S_c_111_n N_VPWR_c_467_n 0.0141975f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_162 N_S_c_112_n N_VPWR_c_467_n 0.00310396f $X=0.69 $Y=1.78 $X2=0 $Y2=0
cc_163 N_S_M1009_g N_VPWR_c_468_n 0.0128318f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_164 N_S_M1013_g N_VPWR_c_475_n 0.00486043f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_165 N_S_M1009_g N_VPWR_c_476_n 0.00486043f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_166 N_S_M1013_g N_VPWR_c_466_n 0.00923967f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_167 N_S_M1009_g N_VPWR_c_466_n 0.00954696f $X=3.305 $Y=2.465 $X2=0 $Y2=0
cc_168 N_S_c_111_n N_A_210_367#_M1017_d 0.00221108f $X=2.905 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_169 N_S_c_111_n N_A_210_367#_M1002_d 0.00235291f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_170 N_S_c_111_n N_A_210_367#_c_543_n 0.0202162f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_171 N_S_c_111_n N_A_317_367#_M1005_s 0.00229936f $X=2.905 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_172 N_S_c_114_n N_A_317_367#_M1009_s 0.00244702f $X=3.08 $Y=1.695 $X2=0 $Y2=0
cc_173 N_S_c_111_n N_A_317_367#_c_572_n 0.0202647f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_174 N_S_c_111_n N_A_317_367#_c_573_n 0.00280043f $X=2.905 $Y=1.78 $X2=0 $Y2=0
cc_175 N_S_c_102_n N_VGND_c_668_n 0.0195226f $X=0.8 $Y=1.185 $X2=0 $Y2=0
cc_176 N_S_c_102_n N_VGND_c_674_n 0.00564095f $X=0.8 $Y=1.185 $X2=0 $Y2=0
cc_177 N_S_c_102_n N_VGND_c_676_n 0.0107826f $X=0.8 $Y=1.185 $X2=0 $Y2=0
cc_178 N_S_c_103_n N_VGND_c_676_n 0.00447364f $X=2.825 $Y=1.185 $X2=0 $Y2=0
cc_179 N_S_c_103_n N_VGND_c_678_n 0.00486043f $X=2.825 $Y=1.185 $X2=0 $Y2=0
cc_180 N_S_c_103_n N_VGND_c_679_n 0.014644f $X=2.825 $Y=1.185 $X2=0 $Y2=0
cc_181 N_A_41_367#_M1008_g N_A0_c_251_n 0.0426261f $X=1.36 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_41_367#_c_198_n N_A0_c_251_n 3.83942e-19 $X=1.25 $Y=1.43 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_41_367#_c_199_n N_A0_M1005_g 0.00765399f $X=1.25 $Y=1.43 $X2=0 $Y2=0
cc_184 N_A_41_367#_M1008_g A0 0.0100339f $X=1.36 $Y=0.655 $X2=0 $Y2=0
cc_185 N_A_41_367#_c_197_n A0 0.0140973f $X=1.085 $Y=1.07 $X2=0 $Y2=0
cc_186 N_A_41_367#_c_198_n A0 0.0291342f $X=1.25 $Y=1.43 $X2=0 $Y2=0
cc_187 N_A_41_367#_c_199_n N_A0_c_254_n 0.0426261f $X=1.25 $Y=1.43 $X2=0 $Y2=0
cc_188 N_A_41_367#_c_202_n N_VPWR_c_467_n 0.0173862f $X=0.975 $Y=1.725 $X2=0
+ $Y2=0
cc_189 N_A_41_367#_c_203_n N_VPWR_c_475_n 0.0231876f $X=0.33 $Y=2.91 $X2=0 $Y2=0
cc_190 N_A_41_367#_c_202_n N_VPWR_c_476_n 0.00486043f $X=0.975 $Y=1.725 $X2=0
+ $Y2=0
cc_191 N_A_41_367#_M1013_s N_VPWR_c_466_n 0.00371702f $X=0.205 $Y=1.835 $X2=0
+ $Y2=0
cc_192 N_A_41_367#_c_202_n N_VPWR_c_466_n 0.00954696f $X=0.975 $Y=1.725 $X2=0
+ $Y2=0
cc_193 N_A_41_367#_c_203_n N_VPWR_c_466_n 0.0129463f $X=0.33 $Y=2.91 $X2=0 $Y2=0
cc_194 N_A_41_367#_c_199_n N_A_210_367#_c_543_n 0.00142237f $X=1.25 $Y=1.43
+ $X2=0 $Y2=0
cc_195 N_A_41_367#_c_197_n N_VGND_M1007_d 0.00341868f $X=1.085 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_41_367#_M1008_g N_VGND_c_668_n 0.0239221f $X=1.36 $Y=0.655 $X2=0
+ $Y2=0
cc_197 N_A_41_367#_c_197_n N_VGND_c_668_n 0.0290545f $X=1.085 $Y=1.07 $X2=0
+ $Y2=0
cc_198 N_A_41_367#_c_199_n N_VGND_c_668_n 7.47969e-19 $X=1.25 $Y=1.43 $X2=0
+ $Y2=0
cc_199 N_A_41_367#_c_196_n N_VGND_c_674_n 0.0421773f $X=0.585 $Y=0.42 $X2=0
+ $Y2=0
cc_200 N_A_41_367#_M1007_s N_VGND_c_676_n 0.00302127f $X=0.46 $Y=0.235 $X2=0
+ $Y2=0
cc_201 N_A_41_367#_M1008_g N_VGND_c_676_n 0.00695146f $X=1.36 $Y=0.655 $X2=0
+ $Y2=0
cc_202 N_A_41_367#_c_196_n N_VGND_c_676_n 0.0236376f $X=0.585 $Y=0.42 $X2=0
+ $Y2=0
cc_203 N_A_41_367#_M1008_g N_VGND_c_678_n 0.00407992f $X=1.36 $Y=0.655 $X2=0
+ $Y2=0
cc_204 N_A0_M1005_g N_A1_M1002_g 0.062731f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_205 A0 A1 0.0270396f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_206 N_A0_c_254_n A1 0.00239461f $X=1.925 $Y=1.35 $X2=0 $Y2=0
cc_207 A0 N_A1_c_294_n 3.52813e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_208 N_A0_c_254_n N_A1_c_294_n 0.0206179f $X=1.925 $Y=1.35 $X2=0 $Y2=0
cc_209 N_A0_c_251_n N_A1_c_295_n 0.0109388f $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_210 A0 N_A1_c_295_n 0.00376431f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_211 A0 N_A_359_47#_M1010_d 0.00807818f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_212 N_A0_c_251_n N_A_359_47#_c_351_n 0.0039705f $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_213 A0 N_A_359_47#_c_351_n 0.040361f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_214 N_A0_c_251_n N_A_359_47#_c_373_n 6.39834e-19 $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_215 A0 N_A_359_47#_c_373_n 0.0138417f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_216 N_A0_M1005_g N_A_359_47#_c_367_n 0.00386074f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_217 N_A0_M1005_g N_VPWR_c_476_n 0.00357877f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A0_M1005_g N_VPWR_c_466_n 0.00684889f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A0_M1005_g N_A_210_367#_c_543_n 0.00406957f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_220 N_A0_M1005_g N_A_210_367#_c_545_n 2.88213e-19 $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_221 N_A0_M1005_g N_A_210_367#_c_546_n 0.0120816f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_222 N_A0_M1005_g N_A_317_367#_c_573_n 0.0105188f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_223 N_A0_c_251_n N_VGND_c_668_n 0.00224066f $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_224 A0 N_VGND_c_668_n 0.0273347f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_225 N_A0_c_251_n N_VGND_c_676_n 0.00595922f $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_226 A0 N_VGND_c_676_n 0.0110452f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_227 N_A0_c_251_n N_VGND_c_678_n 0.00375793f $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_228 A0 N_VGND_c_678_n 0.011392f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_229 A0 A_287_47# 0.00754813f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_230 N_A1_c_295_n N_A_359_47#_c_351_n 0.0174308f $X=2.375 $Y=1.185 $X2=0 $Y2=0
cc_231 N_A1_M1002_g N_A_359_47#_c_343_n 0.0103388f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_232 A1 N_A_359_47#_c_355_n 0.0118505f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_233 N_A1_c_295_n N_A_359_47#_c_355_n 0.00199054f $X=2.375 $Y=1.185 $X2=0
+ $Y2=0
cc_234 A1 N_A_359_47#_c_373_n 0.0342358f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_235 N_A1_c_294_n N_A_359_47#_c_373_n 0.00453156f $X=2.375 $Y=1.35 $X2=0 $Y2=0
cc_236 N_A1_c_295_n N_A_359_47#_c_373_n 0.00424005f $X=2.375 $Y=1.185 $X2=0
+ $Y2=0
cc_237 N_A1_M1002_g N_A_359_47#_c_367_n 0.00624864f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_238 N_A1_M1002_g N_VPWR_c_476_n 0.00357877f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A1_M1002_g N_VPWR_c_466_n 0.00667818f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A1_M1002_g N_A_210_367#_c_545_n 0.00200444f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_241 N_A1_M1002_g N_A_210_367#_c_546_n 0.00698156f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_242 N_A1_M1002_g N_A_317_367#_c_573_n 0.0133246f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_243 N_A1_M1002_g N_A_317_367#_c_575_n 0.00635247f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_244 N_A1_c_295_n N_VGND_c_676_n 0.00585922f $X=2.375 $Y=1.185 $X2=0 $Y2=0
cc_245 N_A1_c_295_n N_VGND_c_678_n 0.00374367f $X=2.375 $Y=1.185 $X2=0 $Y2=0
cc_246 N_A1_c_295_n N_VGND_c_679_n 0.00240485f $X=2.375 $Y=1.185 $X2=0 $Y2=0
cc_247 N_A_359_47#_c_343_n N_VPWR_M1009_d 0.00252989f $X=3.425 $Y=2.125 $X2=0
+ $Y2=0
cc_248 N_A_359_47#_c_335_n N_VPWR_M1009_d 5.24721e-19 $X=3.537 $Y=2.035 $X2=0
+ $Y2=0
cc_249 N_A_359_47#_M1003_g N_VPWR_c_468_n 0.01186f $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A_359_47#_M1006_g N_VPWR_c_468_n 6.28154e-19 $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_251 N_A_359_47#_c_343_n N_VPWR_c_468_n 0.0133508f $X=3.425 $Y=2.125 $X2=0
+ $Y2=0
cc_252 N_A_359_47#_M1003_g N_VPWR_c_469_n 7.27171e-19 $X=3.735 $Y=2.465 $X2=0
+ $Y2=0
cc_253 N_A_359_47#_M1006_g N_VPWR_c_469_n 0.0143393f $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_254 N_A_359_47#_M1012_g N_VPWR_c_469_n 0.0143393f $X=4.595 $Y=2.465 $X2=0
+ $Y2=0
cc_255 N_A_359_47#_M1016_g N_VPWR_c_469_n 7.27171e-19 $X=5.025 $Y=2.465 $X2=0
+ $Y2=0
cc_256 N_A_359_47#_M1012_g N_VPWR_c_470_n 7.42371e-19 $X=4.595 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_A_359_47#_M1016_g N_VPWR_c_470_n 0.0157104f $X=5.025 $Y=2.465 $X2=0
+ $Y2=0
cc_258 N_A_359_47#_M1003_g N_VPWR_c_471_n 0.00486043f $X=3.735 $Y=2.465 $X2=0
+ $Y2=0
cc_259 N_A_359_47#_M1006_g N_VPWR_c_471_n 0.00486043f $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_260 N_A_359_47#_M1012_g N_VPWR_c_473_n 0.00486043f $X=4.595 $Y=2.465 $X2=0
+ $Y2=0
cc_261 N_A_359_47#_M1016_g N_VPWR_c_473_n 0.00486043f $X=5.025 $Y=2.465 $X2=0
+ $Y2=0
cc_262 N_A_359_47#_M1005_d N_VPWR_c_466_n 0.00225186f $X=2 $Y=1.835 $X2=0 $Y2=0
cc_263 N_A_359_47#_M1003_g N_VPWR_c_466_n 0.00824727f $X=3.735 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A_359_47#_M1006_g N_VPWR_c_466_n 0.00824727f $X=4.165 $Y=2.465 $X2=0
+ $Y2=0
cc_265 N_A_359_47#_M1012_g N_VPWR_c_466_n 0.00824727f $X=4.595 $Y=2.465 $X2=0
+ $Y2=0
cc_266 N_A_359_47#_M1016_g N_VPWR_c_466_n 0.00824727f $X=5.025 $Y=2.465 $X2=0
+ $Y2=0
cc_267 N_A_359_47#_c_343_n N_A_210_367#_M1002_d 0.00583293f $X=3.425 $Y=2.125
+ $X2=0 $Y2=0
cc_268 N_A_359_47#_M1005_d N_A_210_367#_c_546_n 0.00357898f $X=2 $Y=1.835 $X2=0
+ $Y2=0
cc_269 N_A_359_47#_c_343_n N_A_317_367#_M1009_s 0.00503349f $X=3.425 $Y=2.125
+ $X2=0 $Y2=0
cc_270 N_A_359_47#_M1005_d N_A_317_367#_c_573_n 0.0037055f $X=2 $Y=1.835 $X2=0
+ $Y2=0
cc_271 N_A_359_47#_c_343_n N_A_317_367#_c_573_n 0.0277572f $X=3.425 $Y=2.125
+ $X2=0 $Y2=0
cc_272 N_A_359_47#_c_367_n N_A_317_367#_c_573_n 0.0160615f $X=2.305 $Y=2.185
+ $X2=0 $Y2=0
cc_273 N_A_359_47#_c_343_n N_A_317_367#_c_575_n 0.0204038f $X=3.425 $Y=2.125
+ $X2=0 $Y2=0
cc_274 N_A_359_47#_M1001_g N_X_c_602_n 0.0138111f $X=4.095 $Y=0.655 $X2=0 $Y2=0
cc_275 N_A_359_47#_M1014_g N_X_c_602_n 0.0141287f $X=4.525 $Y=0.655 $X2=0 $Y2=0
cc_276 N_A_359_47#_c_336_n N_X_c_602_n 0.0469272f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_277 N_A_359_47#_c_337_n N_X_c_602_n 0.00273301f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_278 N_A_359_47#_M1000_g N_X_c_603_n 0.00137282f $X=3.665 $Y=0.655 $X2=0 $Y2=0
cc_279 N_A_359_47#_c_334_n N_X_c_603_n 0.0132011f $X=3.51 $Y=1.405 $X2=0 $Y2=0
cc_280 N_A_359_47#_c_336_n N_X_c_603_n 0.0170082f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_281 N_A_359_47#_c_337_n N_X_c_603_n 0.00283411f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_282 N_A_359_47#_M1006_g N_X_c_609_n 0.0130035f $X=4.165 $Y=2.465 $X2=0 $Y2=0
cc_283 N_A_359_47#_M1012_g N_X_c_609_n 0.0131657f $X=4.595 $Y=2.465 $X2=0 $Y2=0
cc_284 N_A_359_47#_c_336_n N_X_c_609_n 0.0469271f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_285 N_A_359_47#_c_337_n N_X_c_609_n 0.00276559f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_286 N_A_359_47#_M1003_g N_X_c_610_n 7.14036e-19 $X=3.735 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A_359_47#_c_335_n N_X_c_610_n 0.00595425f $X=3.537 $Y=2.035 $X2=0 $Y2=0
cc_288 N_A_359_47#_c_336_n N_X_c_610_n 0.015388f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_289 N_A_359_47#_c_337_n N_X_c_610_n 0.00286879f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_290 N_A_359_47#_M1015_g N_X_c_604_n 0.016842f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_291 N_A_359_47#_c_336_n N_X_c_604_n 0.028847f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_292 N_A_359_47#_c_337_n N_X_c_604_n 0.00638615f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_293 N_A_359_47#_M1016_g N_X_c_611_n 0.0150697f $X=5.025 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A_359_47#_c_336_n N_X_c_611_n 0.0270525f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_295 N_A_359_47#_c_337_n N_X_c_611_n 0.0044365f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_296 N_A_359_47#_M1015_g N_X_c_605_n 0.00262569f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_297 N_A_359_47#_M1016_g N_X_c_605_n 0.00253816f $X=5.025 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A_359_47#_c_336_n N_X_c_605_n 0.0137813f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_299 N_A_359_47#_c_337_n N_X_c_605_n 0.00757919f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_300 N_A_359_47#_c_336_n N_X_c_606_n 0.0182232f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_301 N_A_359_47#_c_337_n N_X_c_606_n 0.00283411f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_302 N_A_359_47#_c_336_n N_X_c_613_n 0.0145779f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_303 N_A_359_47#_c_337_n N_X_c_613_n 0.00286879f $X=5.115 $Y=1.5 $X2=0 $Y2=0
cc_304 N_A_359_47#_M1015_g X 0.00334511f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_305 N_A_359_47#_c_355_n N_VGND_M1004_d 0.0148334f $X=3.425 $Y=0.945 $X2=0
+ $Y2=0
cc_306 N_A_359_47#_c_334_n N_VGND_M1004_d 6.92714e-19 $X=3.51 $Y=1.405 $X2=0
+ $Y2=0
cc_307 N_A_359_47#_M1000_g N_VGND_c_669_n 6.38741e-19 $X=3.665 $Y=0.655 $X2=0
+ $Y2=0
cc_308 N_A_359_47#_M1001_g N_VGND_c_669_n 0.0113089f $X=4.095 $Y=0.655 $X2=0
+ $Y2=0
cc_309 N_A_359_47#_M1014_g N_VGND_c_669_n 0.0113454f $X=4.525 $Y=0.655 $X2=0
+ $Y2=0
cc_310 N_A_359_47#_M1015_g N_VGND_c_669_n 6.45202e-19 $X=4.955 $Y=0.655 $X2=0
+ $Y2=0
cc_311 N_A_359_47#_M1014_g N_VGND_c_670_n 0.00486043f $X=4.525 $Y=0.655 $X2=0
+ $Y2=0
cc_312 N_A_359_47#_M1015_g N_VGND_c_670_n 0.00585385f $X=4.955 $Y=0.655 $X2=0
+ $Y2=0
cc_313 N_A_359_47#_M1015_g N_VGND_c_671_n 0.00335315f $X=4.955 $Y=0.655 $X2=0
+ $Y2=0
cc_314 N_A_359_47#_M1000_g N_VGND_c_672_n 0.00564095f $X=3.665 $Y=0.655 $X2=0
+ $Y2=0
cc_315 N_A_359_47#_M1001_g N_VGND_c_672_n 0.00486043f $X=4.095 $Y=0.655 $X2=0
+ $Y2=0
cc_316 N_A_359_47#_M1010_d N_VGND_c_676_n 0.01122f $X=1.795 $Y=0.235 $X2=0 $Y2=0
cc_317 N_A_359_47#_M1000_g N_VGND_c_676_n 0.00943408f $X=3.665 $Y=0.655 $X2=0
+ $Y2=0
cc_318 N_A_359_47#_M1001_g N_VGND_c_676_n 0.00824727f $X=4.095 $Y=0.655 $X2=0
+ $Y2=0
cc_319 N_A_359_47#_M1014_g N_VGND_c_676_n 0.00824727f $X=4.525 $Y=0.655 $X2=0
+ $Y2=0
cc_320 N_A_359_47#_M1015_g N_VGND_c_676_n 0.0118221f $X=4.955 $Y=0.655 $X2=0
+ $Y2=0
cc_321 N_A_359_47#_c_351_n N_VGND_c_676_n 0.0165136f $X=2.25 $Y=0.36 $X2=0 $Y2=0
cc_322 N_A_359_47#_c_355_n N_VGND_c_676_n 0.0130501f $X=3.425 $Y=0.945 $X2=0
+ $Y2=0
cc_323 N_A_359_47#_c_351_n N_VGND_c_678_n 0.0288329f $X=2.25 $Y=0.36 $X2=0 $Y2=0
cc_324 N_A_359_47#_M1000_g N_VGND_c_679_n 0.0103758f $X=3.665 $Y=0.655 $X2=0
+ $Y2=0
cc_325 N_A_359_47#_M1001_g N_VGND_c_679_n 5.69019e-19 $X=4.095 $Y=0.655 $X2=0
+ $Y2=0
cc_326 N_A_359_47#_c_351_n N_VGND_c_679_n 0.0201164f $X=2.25 $Y=0.36 $X2=0 $Y2=0
cc_327 N_A_359_47#_c_355_n N_VGND_c_679_n 0.0487492f $X=3.425 $Y=0.945 $X2=0
+ $Y2=0
cc_328 N_A_359_47#_c_355_n A_508_47# 0.00298571f $X=3.425 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_329 N_VPWR_c_466_n N_A_210_367#_M1017_d 0.00368223f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_330 N_VPWR_c_466_n N_A_210_367#_M1002_d 0.00215176f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_476_n N_A_210_367#_c_544_n 0.0179183f $X=3.355 $Y=3.33 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_466_n N_A_210_367#_c_544_n 0.0101082f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_476_n N_A_210_367#_c_546_n 0.0810516f $X=3.355 $Y=3.33 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_466_n N_A_210_367#_c_546_n 0.0505225f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_335 N_VPWR_c_466_n N_A_317_367#_M1005_s 0.0021598f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_336 N_VPWR_c_466_n N_A_317_367#_M1009_s 0.00371702f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_476_n N_A_317_367#_c_573_n 0.00331372f $X=3.355 $Y=3.33 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_466_n N_A_317_367#_c_573_n 0.00732526f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_476_n N_A_317_367#_c_575_n 0.0178299f $X=3.355 $Y=3.33 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_466_n N_A_317_367#_c_575_n 0.0100343f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_466_n N_X_M1003_d 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_342 N_VPWR_c_466_n N_X_M1012_d 0.00571434f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_343 N_VPWR_c_471_n N_X_c_647_n 0.0124525f $X=4.215 $Y=3.33 $X2=0 $Y2=0
cc_344 N_VPWR_c_466_n N_X_c_647_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_345 N_VPWR_M1006_s N_X_c_609_n 0.00176461f $X=4.24 $Y=1.835 $X2=0 $Y2=0
cc_346 N_VPWR_c_469_n N_X_c_609_n 0.0170777f $X=4.38 $Y=2.18 $X2=0 $Y2=0
cc_347 N_VPWR_c_473_n N_X_c_651_n 0.0120977f $X=5.075 $Y=3.33 $X2=0 $Y2=0
cc_348 N_VPWR_c_466_n N_X_c_651_n 0.00691495f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_349 N_VPWR_M1016_s N_X_c_611_n 0.00262981f $X=5.1 $Y=1.835 $X2=0 $Y2=0
cc_350 N_VPWR_c_470_n N_X_c_611_n 0.0220026f $X=5.24 $Y=2.18 $X2=0 $Y2=0
cc_351 N_A_210_367#_c_546_n N_A_317_367#_M1005_s 0.00495471f $X=2.405 $Y=2.96
+ $X2=-0.19 $Y2=1.655
cc_352 N_A_210_367#_c_543_n N_A_317_367#_c_572_n 0.034871f $X=1.19 $Y=2.22 $X2=0
+ $Y2=0
cc_353 N_A_210_367#_M1002_d N_A_317_367#_c_573_n 0.00575811f $X=2.43 $Y=1.835
+ $X2=0 $Y2=0
cc_354 N_A_210_367#_c_545_n N_A_317_367#_c_573_n 0.0192788f $X=2.57 $Y=2.95
+ $X2=0 $Y2=0
cc_355 N_A_210_367#_c_546_n N_A_317_367#_c_573_n 0.0220826f $X=2.405 $Y=2.96
+ $X2=0 $Y2=0
cc_356 N_A_210_367#_c_543_n N_A_317_367#_c_574_n 0.0181294f $X=1.19 $Y=2.22
+ $X2=0 $Y2=0
cc_357 N_A_210_367#_c_546_n N_A_317_367#_c_574_n 0.0190344f $X=2.405 $Y=2.96
+ $X2=0 $Y2=0
cc_358 N_A_210_367#_c_545_n N_A_317_367#_c_575_n 0.0180679f $X=2.57 $Y=2.95
+ $X2=0 $Y2=0
cc_359 N_X_c_602_n N_VGND_M1001_d 0.00176461f $X=4.645 $Y=1.15 $X2=0 $Y2=0
cc_360 N_X_c_604_n N_VGND_M1015_d 0.00310671f $X=5.435 $Y=1.15 $X2=0 $Y2=0
cc_361 N_X_c_602_n N_VGND_c_669_n 0.0170777f $X=4.645 $Y=1.15 $X2=0 $Y2=0
cc_362 N_X_c_658_p N_VGND_c_670_n 0.0136943f $X=4.74 $Y=0.42 $X2=0 $Y2=0
cc_363 N_X_c_604_n N_VGND_c_671_n 0.0144005f $X=5.435 $Y=1.15 $X2=0 $Y2=0
cc_364 X N_VGND_c_671_n 0.0389663f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_365 N_X_c_661_p N_VGND_c_672_n 0.0131621f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_366 X N_VGND_c_675_n 0.00857001f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_367 N_X_M1000_s N_VGND_c_676_n 0.00467071f $X=3.74 $Y=0.235 $X2=0 $Y2=0
cc_368 N_X_M1014_s N_VGND_c_676_n 0.0041489f $X=4.6 $Y=0.235 $X2=0 $Y2=0
cc_369 N_X_c_661_p N_VGND_c_676_n 0.00808656f $X=3.88 $Y=0.42 $X2=0 $Y2=0
cc_370 N_X_c_658_p N_VGND_c_676_n 0.00866972f $X=4.74 $Y=0.42 $X2=0 $Y2=0
cc_371 X N_VGND_c_676_n 0.00803447f $X=5.435 $Y=0.47 $X2=0 $Y2=0
cc_372 N_VGND_c_676_n A_287_47# 0.00695948f $X=5.52 $Y=0 $X2=-0.19 $Y2=-0.245
cc_373 N_VGND_c_676_n A_508_47# 0.00314438f $X=5.52 $Y=0 $X2=-0.19 $Y2=-0.245
