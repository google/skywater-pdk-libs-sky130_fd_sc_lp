* File: sky130_fd_sc_lp__or2b_1.pxi.spice
* Created: Fri Aug 28 11:22:10 2020
* 
x_PM_SKY130_FD_SC_LP__OR2B_1%B_N N_B_N_M1006_g N_B_N_c_66_n N_B_N_c_67_n
+ N_B_N_c_68_n N_B_N_M1000_g N_B_N_c_69_n B_N B_N B_N N_B_N_c_72_n
+ PM_SKY130_FD_SC_LP__OR2B_1%B_N
x_PM_SKY130_FD_SC_LP__OR2B_1%A_27_535# N_A_27_535#_M1000_s N_A_27_535#_M1006_s
+ N_A_27_535#_c_106_n N_A_27_535#_c_114_n N_A_27_535#_c_107_n
+ N_A_27_535#_M1003_g N_A_27_535#_c_116_n N_A_27_535#_M1004_g
+ N_A_27_535#_c_109_n N_A_27_535#_c_110_n N_A_27_535#_c_119_n
+ N_A_27_535#_c_111_n N_A_27_535#_c_112_n N_A_27_535#_c_120_n
+ N_A_27_535#_c_121_n N_A_27_535#_c_122_n N_A_27_535#_c_123_n
+ PM_SKY130_FD_SC_LP__OR2B_1%A_27_535#
x_PM_SKY130_FD_SC_LP__OR2B_1%A N_A_M1005_g N_A_M1007_g N_A_c_189_n A A
+ N_A_c_192_n PM_SKY130_FD_SC_LP__OR2B_1%A
x_PM_SKY130_FD_SC_LP__OR2B_1%A_224_382# N_A_224_382#_M1003_d
+ N_A_224_382#_M1004_s N_A_224_382#_M1001_g N_A_224_382#_M1002_g
+ N_A_224_382#_c_232_n N_A_224_382#_c_233_n N_A_224_382#_c_234_n
+ N_A_224_382#_c_235_n N_A_224_382#_c_240_n N_A_224_382#_c_236_n
+ N_A_224_382#_c_237_n PM_SKY130_FD_SC_LP__OR2B_1%A_224_382#
x_PM_SKY130_FD_SC_LP__OR2B_1%VPWR N_VPWR_M1006_d N_VPWR_M1005_d N_VPWR_c_289_n
+ N_VPWR_c_290_n VPWR N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n
+ N_VPWR_c_288_n N_VPWR_c_295_n N_VPWR_c_296_n PM_SKY130_FD_SC_LP__OR2B_1%VPWR
x_PM_SKY130_FD_SC_LP__OR2B_1%X N_X_M1002_d N_X_M1001_d X X X X X X X N_X_c_328_n
+ X PM_SKY130_FD_SC_LP__OR2B_1%X
x_PM_SKY130_FD_SC_LP__OR2B_1%VGND N_VGND_M1000_d N_VGND_M1007_d N_VGND_c_343_n
+ N_VGND_c_344_n VGND N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n
+ N_VGND_c_348_n N_VGND_c_349_n N_VGND_c_350_n PM_SKY130_FD_SC_LP__OR2B_1%VGND
cc_1 VNB N_B_N_M1006_g 0.0128423f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_2 VNB N_B_N_c_66_n 0.02779f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.85
cc_3 VNB N_B_N_c_67_n 0.0182574f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.85
cc_4 VNB N_B_N_c_68_n 0.0206032f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.775
cc_5 VNB N_B_N_c_69_n 0.0194121f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.445
cc_6 VNB B_N 0.0110542f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_7 VNB B_N 0.00115202f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_B_N_c_72_n 0.0288487f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.94
cc_9 VNB N_A_27_535#_c_106_n 0.00717241f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.775
cc_10 VNB N_A_27_535#_c_107_n 0.016828f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.455
cc_11 VNB N_A_27_535#_M1003_g 0.0648518f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_12 VNB N_A_27_535#_c_109_n 0.00325641f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.94
cc_13 VNB N_A_27_535#_c_110_n 0.0515072f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.94
cc_14 VNB N_A_27_535#_c_111_n 0.0166068f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.94
cc_15 VNB N_A_27_535#_c_112_n 0.0130624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_M1005_g 0.031392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_M1007_g 0.0190979f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.775
cc_18 VNB N_A_c_189_n 0.0121131f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.925
cc_19 VNB N_A_224_382#_M1001_g 0.00774477f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.455
cc_20 VNB N_A_224_382#_c_232_n 0.00619551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_224_382#_c_233_n 0.00247405f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.94
cc_22 VNB N_A_224_382#_c_234_n 0.0066068f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.475
cc_23 VNB N_A_224_382#_c_235_n 0.0369761f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=0.925
cc_24 VNB N_A_224_382#_c_236_n 0.00402415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_224_382#_c_237_n 0.0202792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_288_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_328_n 0.0624645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_343_n 0.00471205f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.455
cc_29 VNB N_VGND_c_344_n 0.00700266f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_30 VNB N_VGND_c_345_n 0.0306569f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.94
cc_31 VNB N_VGND_c_346_n 0.0171343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_347_n 0.0153476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_348_n 0.172525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_349_n 0.00439895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_350_n 0.00617187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_B_N_M1006_g 0.0752131f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_37 VPB B_N 0.00525072f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_38 VPB N_A_27_535#_c_106_n 0.00896473f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=0.775
cc_39 VPB N_A_27_535#_c_114_n 0.0446738f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=0.455
cc_40 VPB N_A_27_535#_c_107_n 0.00941559f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=0.455
cc_41 VPB N_A_27_535#_c_116_n 0.0193671f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_42 VPB N_A_27_535#_c_109_n 0.0026256f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.94
cc_43 VPB N_A_27_535#_c_110_n 0.0360718f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.94
cc_44 VPB N_A_27_535#_c_119_n 0.0210677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_27_535#_c_120_n 0.0131023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_27_535#_c_121_n 0.00348275f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_27_535#_c_122_n 0.0461443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_27_535#_c_123_n 0.0122038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_M1005_g 0.0312172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB A 0.00674954f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.28
cc_51 VPB N_A_c_192_n 0.0432937f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.94
cc_52 VPB N_A_224_382#_M1001_g 0.0257567f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=0.455
cc_53 VPB N_A_224_382#_c_233_n 0.00334f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.94
cc_54 VPB N_A_224_382#_c_240_n 0.00469529f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=0.94
cc_55 VPB N_VPWR_c_289_n 0.00513962f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=0.455
cc_56 VPB N_VPWR_c_290_n 0.0167609f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_57 VPB N_VPWR_c_291_n 0.017249f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.94
cc_58 VPB N_VPWR_c_292_n 0.0320985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_293_n 0.0166266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_288_n 0.0649044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_295_n 0.00468717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_296_n 0.00530076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB X 0.0550654f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.28
cc_64 VPB N_X_c_328_n 0.00889774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 N_B_N_M1006_g N_A_27_535#_c_106_n 0.0422431f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_66 N_B_N_c_66_n N_A_27_535#_c_106_n 0.00490563f $X=0.945 $Y=0.85 $X2=0 $Y2=0
cc_67 B_N N_A_27_535#_c_106_n 0.0113512f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_68 B_N N_A_27_535#_c_114_n 0.00118588f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_69 N_B_N_c_68_n N_A_27_535#_M1003_g 0.0197976f $X=1.02 $Y=0.775 $X2=0 $Y2=0
cc_70 B_N N_A_27_535#_M1003_g 0.00590079f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_71 B_N N_A_27_535#_M1003_g 0.00177345f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_72 N_B_N_c_72_n N_A_27_535#_M1003_g 0.00565342f $X=0.535 $Y=0.94 $X2=0 $Y2=0
cc_73 B_N N_A_27_535#_c_116_n 3.74435e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_74 N_B_N_M1006_g N_A_27_535#_c_110_n 0.0275024f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_75 N_B_N_c_67_n N_A_27_535#_c_110_n 0.0171698f $X=0.7 $Y=0.85 $X2=0 $Y2=0
cc_76 N_B_N_c_68_n N_A_27_535#_c_110_n 0.00307339f $X=1.02 $Y=0.775 $X2=0 $Y2=0
cc_77 B_N N_A_27_535#_c_110_n 0.0545498f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_78 B_N N_A_27_535#_c_110_n 0.0301977f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_79 N_B_N_M1006_g N_A_27_535#_c_119_n 0.00404342f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_80 N_B_N_c_67_n N_A_27_535#_c_112_n 0.00698512f $X=0.7 $Y=0.85 $X2=0 $Y2=0
cc_81 N_B_N_c_68_n N_A_27_535#_c_112_n 0.00445262f $X=1.02 $Y=0.775 $X2=0 $Y2=0
cc_82 B_N N_A_27_535#_c_112_n 0.0366577f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_83 N_B_N_M1006_g N_A_27_535#_c_120_n 0.016144f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_84 B_N N_A_27_535#_c_120_n 0.0173693f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_85 N_B_N_M1006_g N_A_27_535#_c_121_n 5.51458e-19 $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_86 B_N N_A_224_382#_c_232_n 0.0136148f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_87 B_N N_A_224_382#_c_233_n 0.00948089f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_88 B_N N_A_224_382#_c_236_n 0.0103058f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_89 B_N N_A_224_382#_c_236_n 0.0018464f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_90 N_B_N_M1006_g N_VPWR_c_289_n 0.00514375f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_91 N_B_N_M1006_g N_VPWR_c_291_n 0.00585385f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_92 N_B_N_M1006_g N_VPWR_c_288_n 0.00854432f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_93 N_B_N_c_68_n N_VGND_c_343_n 0.00283475f $X=1.02 $Y=0.775 $X2=0 $Y2=0
cc_94 N_B_N_c_68_n N_VGND_c_345_n 0.0053901f $X=1.02 $Y=0.775 $X2=0 $Y2=0
cc_95 N_B_N_c_68_n N_VGND_c_348_n 0.0111236f $X=1.02 $Y=0.775 $X2=0 $Y2=0
cc_96 N_A_27_535#_c_114_n N_A_M1005_g 0.00230327f $X=0.97 $Y=2.625 $X2=0 $Y2=0
cc_97 N_A_27_535#_c_109_n N_A_M1005_g 0.0468809f $X=1.455 $Y=1.65 $X2=0 $Y2=0
cc_98 N_A_27_535#_c_120_n N_A_M1005_g 5.22607e-19 $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_27_535#_c_121_n N_A_M1005_g 2.06646e-19 $X=1.14 $Y=2.79 $X2=0 $Y2=0
cc_100 N_A_27_535#_M1003_g N_A_M1007_g 0.0125409f $X=1.45 $Y=0.455 $X2=0 $Y2=0
cc_101 N_A_27_535#_M1003_g N_A_c_189_n 0.0417983f $X=1.45 $Y=0.455 $X2=0 $Y2=0
cc_102 N_A_27_535#_c_114_n A 9.00669e-19 $X=0.97 $Y=2.625 $X2=0 $Y2=0
cc_103 N_A_27_535#_c_116_n A 0.0021965f $X=1.46 $Y=1.725 $X2=0 $Y2=0
cc_104 N_A_27_535#_c_120_n A 0.0127532f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A_27_535#_c_121_n A 0.0258657f $X=1.14 $Y=2.79 $X2=0 $Y2=0
cc_106 N_A_27_535#_c_122_n A 0.00119812f $X=1.14 $Y=2.79 $X2=0 $Y2=0
cc_107 N_A_27_535#_c_116_n N_A_c_192_n 0.00111921f $X=1.46 $Y=1.725 $X2=0 $Y2=0
cc_108 N_A_27_535#_c_121_n N_A_c_192_n 0.00118009f $X=1.14 $Y=2.79 $X2=0 $Y2=0
cc_109 N_A_27_535#_c_122_n N_A_c_192_n 0.0206627f $X=1.14 $Y=2.79 $X2=0 $Y2=0
cc_110 N_A_27_535#_M1003_g N_A_224_382#_c_232_n 0.0085458f $X=1.45 $Y=0.455
+ $X2=0 $Y2=0
cc_111 N_A_27_535#_M1003_g N_A_224_382#_c_233_n 6.27537e-19 $X=1.45 $Y=0.455
+ $X2=0 $Y2=0
cc_112 N_A_27_535#_c_109_n N_A_224_382#_c_233_n 0.00374381f $X=1.455 $Y=1.65
+ $X2=0 $Y2=0
cc_113 N_A_27_535#_c_114_n N_A_224_382#_c_240_n 0.0103571f $X=0.97 $Y=2.625
+ $X2=0 $Y2=0
cc_114 N_A_27_535#_c_107_n N_A_224_382#_c_240_n 0.0104042f $X=1.375 $Y=1.65
+ $X2=0 $Y2=0
cc_115 N_A_27_535#_c_116_n N_A_224_382#_c_240_n 0.0174363f $X=1.46 $Y=1.725
+ $X2=0 $Y2=0
cc_116 N_A_27_535#_c_120_n N_A_224_382#_c_240_n 0.0194524f $X=0.975 $Y=2.465
+ $X2=0 $Y2=0
cc_117 N_A_27_535#_c_122_n N_A_224_382#_c_240_n 9.55916e-19 $X=1.14 $Y=2.79
+ $X2=0 $Y2=0
cc_118 N_A_27_535#_M1003_g N_A_224_382#_c_236_n 0.00531413f $X=1.45 $Y=0.455
+ $X2=0 $Y2=0
cc_119 N_A_27_535#_c_120_n N_VPWR_c_289_n 0.0174947f $X=0.975 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_27_535#_c_121_n N_VPWR_c_289_n 0.0178318f $X=1.14 $Y=2.79 $X2=0 $Y2=0
cc_121 N_A_27_535#_c_122_n N_VPWR_c_289_n 0.00204931f $X=1.14 $Y=2.79 $X2=0
+ $Y2=0
cc_122 N_A_27_535#_c_119_n N_VPWR_c_291_n 0.0170468f $X=0.26 $Y=2.885 $X2=0
+ $Y2=0
cc_123 N_A_27_535#_c_121_n N_VPWR_c_292_n 0.0122174f $X=1.14 $Y=2.79 $X2=0 $Y2=0
cc_124 N_A_27_535#_c_122_n N_VPWR_c_292_n 0.00442206f $X=1.14 $Y=2.79 $X2=0
+ $Y2=0
cc_125 N_A_27_535#_M1006_s N_VPWR_c_288_n 0.00221783f $X=0.135 $Y=2.675 $X2=0
+ $Y2=0
cc_126 N_A_27_535#_c_119_n N_VPWR_c_288_n 0.0116351f $X=0.26 $Y=2.885 $X2=0
+ $Y2=0
cc_127 N_A_27_535#_c_120_n N_VPWR_c_288_n 0.0118802f $X=0.975 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_A_27_535#_c_121_n N_VPWR_c_288_n 0.0115782f $X=1.14 $Y=2.79 $X2=0 $Y2=0
cc_129 N_A_27_535#_c_122_n N_VPWR_c_288_n 0.00275076f $X=1.14 $Y=2.79 $X2=0
+ $Y2=0
cc_130 N_A_27_535#_M1003_g N_VGND_c_343_n 0.00167516f $X=1.45 $Y=0.455 $X2=0
+ $Y2=0
cc_131 N_A_27_535#_c_111_n N_VGND_c_345_n 0.0114393f $X=0.28 $Y=0.447 $X2=0
+ $Y2=0
cc_132 N_A_27_535#_c_112_n N_VGND_c_345_n 0.0362311f $X=0.805 $Y=0.455 $X2=0
+ $Y2=0
cc_133 N_A_27_535#_M1003_g N_VGND_c_346_n 0.00575161f $X=1.45 $Y=0.455 $X2=0
+ $Y2=0
cc_134 N_A_27_535#_M1000_s N_VGND_c_348_n 0.00214766f $X=0.68 $Y=0.245 $X2=0
+ $Y2=0
cc_135 N_A_27_535#_M1003_g N_VGND_c_348_n 0.0106647f $X=1.45 $Y=0.455 $X2=0
+ $Y2=0
cc_136 N_A_27_535#_c_111_n N_VGND_c_348_n 0.00745041f $X=0.28 $Y=0.447 $X2=0
+ $Y2=0
cc_137 N_A_27_535#_c_112_n N_VGND_c_348_n 0.0256541f $X=0.805 $Y=0.455 $X2=0
+ $Y2=0
cc_138 N_A_M1005_g N_A_224_382#_M1001_g 0.0214797f $X=1.82 $Y=2.045 $X2=0 $Y2=0
cc_139 N_A_M1005_g N_A_224_382#_c_232_n 0.00584282f $X=1.82 $Y=2.045 $X2=0 $Y2=0
cc_140 N_A_M1007_g N_A_224_382#_c_232_n 0.0011878f $X=1.88 $Y=0.455 $X2=0 $Y2=0
cc_141 N_A_c_189_n N_A_224_382#_c_232_n 0.00351014f $X=1.85 $Y=0.955 $X2=0 $Y2=0
cc_142 N_A_M1005_g N_A_224_382#_c_233_n 0.00743217f $X=1.82 $Y=2.045 $X2=0 $Y2=0
cc_143 N_A_M1005_g N_A_224_382#_c_234_n 0.0184856f $X=1.82 $Y=2.045 $X2=0 $Y2=0
cc_144 N_A_c_189_n N_A_224_382#_c_234_n 0.00246912f $X=1.85 $Y=0.955 $X2=0 $Y2=0
cc_145 N_A_M1005_g N_A_224_382#_c_235_n 0.0213482f $X=1.82 $Y=2.045 $X2=0 $Y2=0
cc_146 A N_A_224_382#_c_240_n 0.013187f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_147 N_A_c_192_n N_A_224_382#_c_240_n 6.34652e-19 $X=1.82 $Y=2.79 $X2=0 $Y2=0
cc_148 N_A_M1005_g N_A_224_382#_c_236_n 0.00438576f $X=1.82 $Y=2.045 $X2=0 $Y2=0
cc_149 N_A_M1005_g N_A_224_382#_c_237_n 0.00405575f $X=1.82 $Y=2.045 $X2=0 $Y2=0
cc_150 N_A_M1007_g N_A_224_382#_c_237_n 0.0104793f $X=1.88 $Y=0.455 $X2=0 $Y2=0
cc_151 N_A_M1005_g N_VPWR_c_290_n 0.0113561f $X=1.82 $Y=2.045 $X2=0 $Y2=0
cc_152 A N_VPWR_c_290_n 0.0496084f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_153 A N_VPWR_c_292_n 0.010049f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_154 N_A_c_192_n N_VPWR_c_292_n 0.00506192f $X=1.82 $Y=2.79 $X2=0 $Y2=0
cc_155 A N_VPWR_c_288_n 0.00949318f $X=1.595 $Y=2.32 $X2=0 $Y2=0
cc_156 N_A_c_192_n N_VPWR_c_288_n 0.00375854f $X=1.82 $Y=2.79 $X2=0 $Y2=0
cc_157 N_A_M1005_g N_VGND_c_344_n 6.65525e-19 $X=1.82 $Y=2.045 $X2=0 $Y2=0
cc_158 N_A_M1007_g N_VGND_c_344_n 0.00520522f $X=1.88 $Y=0.455 $X2=0 $Y2=0
cc_159 N_A_M1007_g N_VGND_c_346_n 0.00575161f $X=1.88 $Y=0.455 $X2=0 $Y2=0
cc_160 N_A_M1007_g N_VGND_c_348_n 0.0108714f $X=1.88 $Y=0.455 $X2=0 $Y2=0
cc_161 N_A_c_189_n N_VGND_c_348_n 9.39959e-19 $X=1.85 $Y=0.955 $X2=0 $Y2=0
cc_162 N_A_224_382#_M1001_g N_VPWR_c_290_n 0.0230628f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_224_382#_c_233_n N_VPWR_c_290_n 0.00275739f $X=1.635 $Y=1.88 $X2=0
+ $Y2=0
cc_164 N_A_224_382#_c_234_n N_VPWR_c_290_n 0.0196818f $X=2.27 $Y=1.36 $X2=0
+ $Y2=0
cc_165 N_A_224_382#_c_235_n N_VPWR_c_290_n 0.00358941f $X=2.27 $Y=1.36 $X2=0
+ $Y2=0
cc_166 N_A_224_382#_M1001_g N_VPWR_c_293_n 0.00486043f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_224_382#_M1001_g N_VPWR_c_288_n 0.00923188f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_224_382#_c_240_n A_307_367# 0.00100994f $X=1.245 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_224_382#_M1001_g X 0.00335524f $X=2.345 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_224_382#_c_235_n X 5.95802e-19 $X=2.27 $Y=1.36 $X2=0 $Y2=0
cc_171 N_A_224_382#_M1001_g N_X_c_328_n 0.0112229f $X=2.345 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A_224_382#_c_234_n N_X_c_328_n 0.0271104f $X=2.27 $Y=1.36 $X2=0 $Y2=0
cc_173 N_A_224_382#_c_237_n N_X_c_328_n 0.0159898f $X=2.292 $Y=1.195 $X2=0 $Y2=0
cc_174 N_A_224_382#_c_232_n N_VGND_c_344_n 0.0248689f $X=1.665 $Y=0.455 $X2=0
+ $Y2=0
cc_175 N_A_224_382#_c_234_n N_VGND_c_344_n 0.0292369f $X=2.27 $Y=1.36 $X2=0
+ $Y2=0
cc_176 N_A_224_382#_c_235_n N_VGND_c_344_n 0.00530449f $X=2.27 $Y=1.36 $X2=0
+ $Y2=0
cc_177 N_A_224_382#_c_237_n N_VGND_c_344_n 0.0155923f $X=2.292 $Y=1.195 $X2=0
+ $Y2=0
cc_178 N_A_224_382#_c_232_n N_VGND_c_346_n 0.0113468f $X=1.665 $Y=0.455 $X2=0
+ $Y2=0
cc_179 N_A_224_382#_c_237_n N_VGND_c_347_n 0.00477554f $X=2.292 $Y=1.195 $X2=0
+ $Y2=0
cc_180 N_A_224_382#_M1003_d N_VGND_c_348_n 0.00325517f $X=1.525 $Y=0.245 $X2=0
+ $Y2=0
cc_181 N_A_224_382#_c_232_n N_VGND_c_348_n 0.00871125f $X=1.665 $Y=0.455 $X2=0
+ $Y2=0
cc_182 N_A_224_382#_c_237_n N_VGND_c_348_n 0.00919076f $X=2.292 $Y=1.195 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_288_n N_X_M1001_d 0.00371702f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_290_n X 0.0482852f $X=2.075 $Y=1.98 $X2=0 $Y2=0
cc_185 N_VPWR_c_293_n X 0.0228292f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_186 N_VPWR_c_288_n X 0.0127519f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_187 N_X_c_328_n N_VGND_c_347_n 0.018528f $X=2.62 $Y=0.42 $X2=0 $Y2=0
cc_188 N_X_M1002_d N_VGND_c_348_n 0.00368844f $X=2.48 $Y=0.245 $X2=0 $Y2=0
cc_189 N_X_c_328_n N_VGND_c_348_n 0.0104192f $X=2.62 $Y=0.42 $X2=0 $Y2=0
