* File: sky130_fd_sc_lp__dlrtp_4.pxi.spice
* Created: Fri Aug 28 10:27:19 2020
* 
x_PM_SKY130_FD_SC_LP__DLRTP_4%D N_D_M1001_g N_D_c_170_n N_D_M1006_g N_D_c_172_n
+ D D D D D N_D_c_175_n N_D_c_176_n D PM_SKY130_FD_SC_LP__DLRTP_4%D
x_PM_SKY130_FD_SC_LP__DLRTP_4%GATE N_GATE_c_210_n N_GATE_M1022_g N_GATE_M1025_g
+ N_GATE_c_212_n N_GATE_c_213_n GATE GATE GATE GATE N_GATE_c_215_n
+ PM_SKY130_FD_SC_LP__DLRTP_4%GATE
x_PM_SKY130_FD_SC_LP__DLRTP_4%A_267_464# N_A_267_464#_M1025_d
+ N_A_267_464#_M1022_d N_A_267_464#_c_258_n N_A_267_464#_c_259_n
+ N_A_267_464#_c_260_n N_A_267_464#_M1002_g N_A_267_464#_c_261_n
+ N_A_267_464#_M1000_g N_A_267_464#_M1020_g N_A_267_464#_M1017_g
+ N_A_267_464#_c_265_n N_A_267_464#_c_266_n N_A_267_464#_c_267_n
+ N_A_267_464#_c_280_n N_A_267_464#_c_268_n N_A_267_464#_c_269_n
+ N_A_267_464#_c_270_n N_A_267_464#_c_271_n N_A_267_464#_c_272_n
+ N_A_267_464#_c_273_n N_A_267_464#_c_274_n N_A_267_464#_c_275_n
+ N_A_267_464#_c_276_n N_A_267_464#_c_277_n
+ PM_SKY130_FD_SC_LP__DLRTP_4%A_267_464#
x_PM_SKY130_FD_SC_LP__DLRTP_4%A_49_70# N_A_49_70#_M1001_s N_A_49_70#_M1006_s
+ N_A_49_70#_c_417_n N_A_49_70#_M1012_g N_A_49_70#_M1004_g N_A_49_70#_c_419_n
+ N_A_49_70#_c_425_n N_A_49_70#_c_436_n N_A_49_70#_c_426_n N_A_49_70#_c_427_n
+ N_A_49_70#_c_428_n N_A_49_70#_c_429_n N_A_49_70#_c_420_n N_A_49_70#_c_421_n
+ N_A_49_70#_c_422_n PM_SKY130_FD_SC_LP__DLRTP_4%A_49_70#
x_PM_SKY130_FD_SC_LP__DLRTP_4%A_414_47# N_A_414_47#_M1002_s N_A_414_47#_M1000_s
+ N_A_414_47#_M1009_g N_A_414_47#_M1016_g N_A_414_47#_c_513_n
+ N_A_414_47#_c_514_n N_A_414_47#_c_544_n N_A_414_47#_c_515_n
+ N_A_414_47#_c_516_n N_A_414_47#_c_517_n N_A_414_47#_c_518_n
+ N_A_414_47#_c_523_n N_A_414_47#_c_524_n N_A_414_47#_c_525_n
+ N_A_414_47#_c_526_n N_A_414_47#_c_519_n N_A_414_47#_c_520_n
+ N_A_414_47#_c_528_n N_A_414_47#_c_529_n PM_SKY130_FD_SC_LP__DLRTP_4%A_414_47#
x_PM_SKY130_FD_SC_LP__DLRTP_4%A_857_21# N_A_857_21#_M1013_s N_A_857_21#_M1014_d
+ N_A_857_21#_c_644_n N_A_857_21#_M1024_g N_A_857_21#_M1010_g
+ N_A_857_21#_c_657_n N_A_857_21#_M1008_g N_A_857_21#_c_645_n
+ N_A_857_21#_M1003_g N_A_857_21#_c_658_n N_A_857_21#_M1015_g
+ N_A_857_21#_c_646_n N_A_857_21#_M1005_g N_A_857_21#_c_659_n
+ N_A_857_21#_M1018_g N_A_857_21#_c_647_n N_A_857_21#_M1011_g
+ N_A_857_21#_c_660_n N_A_857_21#_M1023_g N_A_857_21#_c_648_n
+ N_A_857_21#_M1019_g N_A_857_21#_c_649_n N_A_857_21#_c_661_n
+ N_A_857_21#_c_662_n N_A_857_21#_c_663_n N_A_857_21#_c_683_n
+ N_A_857_21#_c_650_n N_A_857_21#_c_689_p N_A_857_21#_c_686_p
+ N_A_857_21#_c_753_p N_A_857_21#_c_714_p N_A_857_21#_c_651_n
+ N_A_857_21#_c_652_n N_A_857_21#_c_769_p N_A_857_21#_c_725_p
+ N_A_857_21#_c_653_n N_A_857_21#_c_654_n N_A_857_21#_c_655_n
+ PM_SKY130_FD_SC_LP__DLRTP_4%A_857_21#
x_PM_SKY130_FD_SC_LP__DLRTP_4%A_671_47# N_A_671_47#_M1009_d N_A_671_47#_M1020_d
+ N_A_671_47#_c_821_n N_A_671_47#_c_822_n N_A_671_47#_c_823_n
+ N_A_671_47#_c_824_n N_A_671_47#_c_825_n N_A_671_47#_M1013_g
+ N_A_671_47#_c_834_n N_A_671_47#_M1014_g N_A_671_47#_c_837_n
+ N_A_671_47#_c_835_n N_A_671_47#_c_826_n N_A_671_47#_c_846_n
+ N_A_671_47#_c_827_n N_A_671_47#_c_828_n N_A_671_47#_c_829_n
+ N_A_671_47#_c_830_n N_A_671_47#_c_855_n N_A_671_47#_c_831_n
+ N_A_671_47#_c_832_n PM_SKY130_FD_SC_LP__DLRTP_4%A_671_47#
x_PM_SKY130_FD_SC_LP__DLRTP_4%RESET_B N_RESET_B_M1007_g N_RESET_B_M1021_g
+ RESET_B RESET_B RESET_B N_RESET_B_c_938_n N_RESET_B_c_939_n
+ PM_SKY130_FD_SC_LP__DLRTP_4%RESET_B
x_PM_SKY130_FD_SC_LP__DLRTP_4%VPWR N_VPWR_M1006_d N_VPWR_M1000_d N_VPWR_M1010_d
+ N_VPWR_M1007_d N_VPWR_M1015_s N_VPWR_M1023_s N_VPWR_c_986_n N_VPWR_c_987_n
+ N_VPWR_c_988_n N_VPWR_c_989_n N_VPWR_c_990_n N_VPWR_c_991_n N_VPWR_c_992_n
+ N_VPWR_c_993_n N_VPWR_c_994_n VPWR N_VPWR_c_995_n N_VPWR_c_996_n
+ N_VPWR_c_997_n N_VPWR_c_998_n N_VPWR_c_999_n N_VPWR_c_1000_n N_VPWR_c_1001_n
+ N_VPWR_c_1002_n N_VPWR_c_985_n PM_SKY130_FD_SC_LP__DLRTP_4%VPWR
x_PM_SKY130_FD_SC_LP__DLRTP_4%Q N_Q_M1003_d N_Q_M1011_d N_Q_M1008_d N_Q_M1018_d
+ N_Q_c_1134_n N_Q_c_1092_n N_Q_c_1098_n N_Q_c_1099_n N_Q_c_1093_n N_Q_c_1094_n
+ N_Q_c_1095_n N_Q_c_1138_n N_Q_c_1100_n Q Q PM_SKY130_FD_SC_LP__DLRTP_4%Q
x_PM_SKY130_FD_SC_LP__DLRTP_4%VGND N_VGND_M1001_d N_VGND_M1002_d N_VGND_M1024_d
+ N_VGND_M1021_d N_VGND_M1005_s N_VGND_M1019_s N_VGND_c_1154_n N_VGND_c_1155_n
+ N_VGND_c_1156_n N_VGND_c_1157_n N_VGND_c_1158_n N_VGND_c_1159_n
+ N_VGND_c_1160_n N_VGND_c_1161_n N_VGND_c_1162_n VGND N_VGND_c_1163_n
+ N_VGND_c_1164_n N_VGND_c_1165_n N_VGND_c_1166_n N_VGND_c_1167_n
+ N_VGND_c_1168_n N_VGND_c_1169_n N_VGND_c_1170_n N_VGND_c_1171_n
+ N_VGND_c_1172_n PM_SKY130_FD_SC_LP__DLRTP_4%VGND
cc_1 VNB N_D_c_170_n 0.0234588f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.363
cc_2 VNB N_D_M1006_g 0.00602934f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_3 VNB N_D_c_172_n 0.0216329f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.55
cc_4 VNB D 8.16722e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB D 0.00235627f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_D_c_175_n 0.0214688f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_7 VNB N_D_c_176_n 0.0227023f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=0.88
cc_8 VNB N_GATE_c_210_n 0.0174047f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.88
cc_9 VNB N_GATE_M1022_g 0.00528957f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.56
cc_10 VNB N_GATE_c_212_n 0.0222961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_GATE_c_213_n 0.0232171f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.55
cc_12 VNB GATE 0.00819805f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_13 VNB N_GATE_c_215_n 0.0163851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_267_464#_c_258_n 0.0216449f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_15 VNB N_A_267_464#_c_259_n 0.0210588f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_16 VNB N_A_267_464#_c_260_n 0.0203385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_267_464#_c_261_n 0.023481f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_18 VNB N_A_267_464#_M1000_g 7.34616e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_267_464#_M1020_g 0.00233989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_267_464#_M1017_g 0.0295526f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_21 VNB N_A_267_464#_c_265_n 0.0092194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_267_464#_c_266_n 0.00495479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_267_464#_c_267_n 0.0274767f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.965
cc_24 VNB N_A_267_464#_c_268_n 0.0191013f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.035
cc_25 VNB N_A_267_464#_c_269_n 0.00133745f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.902
cc_26 VNB N_A_267_464#_c_270_n 0.00410061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_267_464#_c_271_n 7.42849e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_267_464#_c_272_n 9.75862e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_267_464#_c_273_n 0.0151017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_267_464#_c_274_n 0.00125452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_267_464#_c_275_n 0.0346245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_267_464#_c_276_n 0.00343068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_267_464#_c_277_n 0.0320748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_49_70#_c_417_n 0.00597403f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_35 VNB N_A_49_70#_M1012_g 0.0379096f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_36 VNB N_A_49_70#_c_419_n 0.0592959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_49_70#_c_420_n 0.00243056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_49_70#_c_421_n 0.0220135f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.665
cc_39 VNB N_A_49_70#_c_422_n 0.0111948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_414_47#_M1009_g 0.0236944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_414_47#_c_513_n 0.0156945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_414_47#_c_514_n 0.00487002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_414_47#_c_515_n 0.0114319f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.045
cc_44 VNB N_A_414_47#_c_516_n 0.0120226f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_45 VNB N_A_414_47#_c_517_n 0.00909023f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_46 VNB N_A_414_47#_c_518_n 0.00355905f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=0.88
cc_47 VNB N_A_414_47#_c_519_n 0.00344051f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.665
cc_48 VNB N_A_414_47#_c_520_n 0.0306673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_857_21#_c_644_n 0.0178455f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_50 VNB N_A_857_21#_c_645_n 0.0164206f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_857_21#_c_646_n 0.0173233f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_52 VNB N_A_857_21#_c_647_n 0.0173053f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.84
cc_53 VNB N_A_857_21#_c_648_n 0.0197006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_857_21#_c_649_n 0.0134227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_857_21#_c_650_n 0.00138081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_857_21#_c_651_n 0.00118879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_857_21#_c_652_n 4.64928e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_857_21#_c_653_n 0.0010166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_857_21#_c_654_n 0.0355567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_857_21#_c_655_n 0.0732176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_671_47#_c_821_n 0.0582477f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_62 VNB N_A_671_47#_c_822_n 0.0327582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_671_47#_c_823_n 0.00995698f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.55
cc_64 VNB N_A_671_47#_c_824_n 0.0118398f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_65 VNB N_A_671_47#_c_825_n 0.0147854f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_66 VNB N_A_671_47#_c_826_n 0.0122487f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_67 VNB N_A_671_47#_c_827_n 0.00160875f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.555
cc_68 VNB N_A_671_47#_c_828_n 0.0030201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_671_47#_c_829_n 0.0117491f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.987
cc_70 VNB N_A_671_47#_c_830_n 0.0355337f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.295
cc_71 VNB N_A_671_47#_c_831_n 0.00434093f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.925
cc_72 VNB N_A_671_47#_c_832_n 0.00659665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_RESET_B_M1007_g 3.97806e-19 $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.56
cc_74 VNB RESET_B 0.00521677f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_75 VNB N_RESET_B_c_938_n 0.0338036f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_76 VNB N_RESET_B_c_939_n 0.0171443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VPWR_c_985_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_Q_c_1092_n 0.00211134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_Q_c_1093_n 0.00243449f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_80 VNB N_Q_c_1094_n 0.00195287f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=0.88
cc_81 VNB N_Q_c_1095_n 0.0022743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB Q 0.0129987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB Q 0.0219117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1154_n 0.00797237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1155_n 0.002833f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.045
cc_86 VNB N_VGND_c_1156_n 0.010113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1157_n 0.00317786f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.987
cc_88 VNB N_VGND_c_1158_n 0.00715738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1159_n 0.0150197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1160_n 0.0314892f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.902
cc_91 VNB N_VGND_c_1161_n 0.0302977f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.925
cc_92 VNB N_VGND_c_1162_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1163_n 0.0360874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1164_n 0.0380679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1165_n 0.0350656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1166_n 0.0159998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1167_n 0.0159657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1168_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1169_n 0.00583882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1170_n 0.0059813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1171_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1172_n 0.444062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VPB N_D_M1006_g 0.055239f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.64
cc_104 VPB D 0.00560473f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_105 VPB N_GATE_M1022_g 0.0502117f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.56
cc_106 VPB GATE 0.00915375f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_107 VPB N_A_267_464#_M1000_g 0.0526669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_267_464#_M1020_g 0.0464944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_267_464#_c_280_n 0.0147639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_267_464#_c_271_n 0.00323064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_267_464#_c_272_n 0.0511566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_49_70#_M1004_g 0.0219298f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_113 VPB N_A_49_70#_c_419_n 0.0325279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_49_70#_c_425_n 0.0104445f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.045
cc_115 VPB N_A_49_70#_c_426_n 0.0247024f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.555
cc_116 VPB N_A_49_70#_c_427_n 0.001675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_49_70#_c_428_n 0.0030263f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.84
cc_118 VPB N_A_49_70#_c_429_n 0.0293387f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.987
cc_119 VPB N_A_49_70#_c_420_n 0.0119654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_49_70#_c_421_n 0.0542075f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.665
cc_121 VPB N_A_414_47#_M1016_g 0.0183504f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_122 VPB N_A_414_47#_c_518_n 0.00408273f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=0.88
cc_123 VPB N_A_414_47#_c_523_n 0.0162211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_414_47#_c_524_n 8.66281e-19 $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.555
cc_125 VPB N_A_414_47#_c_525_n 0.0022396f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_414_47#_c_526_n 0.00593147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_414_47#_c_519_n 0.0130225f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.665
cc_128 VPB N_A_414_47#_c_528_n 0.036305f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.925
cc_129 VPB N_A_414_47#_c_529_n 0.00267949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_857_21#_M1010_g 0.021918f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_131 VPB N_A_857_21#_c_657_n 0.01643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_857_21#_c_658_n 0.0152002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_857_21#_c_659_n 0.015197f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.555
cc_134 VPB N_A_857_21#_c_660_n 0.0186488f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.295
cc_135 VPB N_A_857_21#_c_661_n 0.00333919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_857_21#_c_662_n 0.0367893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_857_21#_c_663_n 0.00420734f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_857_21#_c_652_n 0.00110232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_857_21#_c_654_n 0.0170152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_857_21#_c_655_n 0.0221186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_671_47#_c_824_n 0.00973013f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_142 VPB N_A_671_47#_c_834_n 0.0207962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_671_47#_c_835_n 0.00605292f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.045
cc_144 VPB N_A_671_47#_c_830_n 0.00773475f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.295
cc_145 VPB N_RESET_B_M1007_g 0.0192636f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.56
cc_146 VPB RESET_B 0.00118525f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.64
cc_147 VPB N_VPWR_c_986_n 0.00543707f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.045
cc_148 VPB N_VPWR_c_987_n 0.00859155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_988_n 0.0121674f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.84
cc_150 VPB N_VPWR_c_989_n 0.00431365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_990_n 3.16879e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_991_n 0.0141676f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.925
cc_153 VPB N_VPWR_c_992_n 0.0419756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_993_n 0.0463215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_994_n 0.00381736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_995_n 0.0515085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_996_n 0.014796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_997_n 0.0154186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_998_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_999_n 0.02506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1000_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1001_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1002_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_985_n 0.112422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_Q_c_1098_n 0.0031952f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.045
cc_166 VPB N_Q_c_1099_n 0.00209769f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.045
cc_167 VPB N_Q_c_1100_n 0.0148421f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.035
cc_168 VPB Q 0.00467239f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 N_D_c_172_n N_GATE_c_210_n 0.0140295f $X=0.697 $Y=1.55 $X2=-0.19
+ $Y2=-0.245
cc_170 N_D_M1006_g N_GATE_M1022_g 0.0258826f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_171 D N_GATE_M1022_g 0.00165826f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_172 D N_GATE_c_212_n 0.00314813f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_173 N_D_c_176_n N_GATE_c_212_n 0.00746628f $X=0.697 $Y=0.88 $X2=0 $Y2=0
cc_174 N_D_c_170_n N_GATE_c_213_n 0.0140295f $X=0.697 $Y=1.363 $X2=0 $Y2=0
cc_175 D N_GATE_c_213_n 3.71975e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_176 N_D_M1006_g GATE 0.0014688f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_177 D GATE 0.102427f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_178 N_D_c_175_n GATE 0.00390713f $X=0.72 $Y=1.045 $X2=0 $Y2=0
cc_179 D N_GATE_c_215_n 3.71975e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_180 N_D_c_175_n N_GATE_c_215_n 0.0140295f $X=0.72 $Y=1.045 $X2=0 $Y2=0
cc_181 D N_A_49_70#_c_419_n 0.113039f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_182 N_D_c_176_n N_A_49_70#_c_419_n 0.0402501f $X=0.697 $Y=0.88 $X2=0 $Y2=0
cc_183 N_D_M1006_g N_A_49_70#_c_425_n 0.0147197f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_184 D N_A_49_70#_c_425_n 0.0206645f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_185 N_D_M1006_g N_A_49_70#_c_436_n 0.00128408f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_186 N_D_M1006_g N_A_49_70#_c_427_n 4.23593e-19 $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_187 N_D_M1006_g N_A_49_70#_c_429_n 2.2485e-19 $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_188 N_D_M1006_g N_VPWR_c_986_n 0.0103896f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_189 N_D_M1006_g N_VPWR_c_999_n 0.00413917f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_190 N_D_M1006_g N_VPWR_c_985_n 0.00422746f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_191 D N_VGND_M1001_d 0.00451906f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_192 D N_VGND_c_1154_n 0.0147113f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_193 N_D_c_176_n N_VGND_c_1154_n 0.00455991f $X=0.697 $Y=0.88 $X2=0 $Y2=0
cc_194 D N_VGND_c_1161_n 0.00433101f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_195 N_D_c_176_n N_VGND_c_1161_n 0.00441982f $X=0.697 $Y=0.88 $X2=0 $Y2=0
cc_196 D N_VGND_c_1172_n 0.00590997f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_197 D N_VGND_c_1172_n 0.00272067f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_198 N_D_c_175_n N_VGND_c_1172_n 2.83568e-19 $X=0.72 $Y=1.045 $X2=0 $Y2=0
cc_199 N_D_c_176_n N_VGND_c_1172_n 0.00854955f $X=0.697 $Y=0.88 $X2=0 $Y2=0
cc_200 N_GATE_c_210_n N_A_267_464#_c_259_n 0.00374353f $X=1.26 $Y=1.55 $X2=0
+ $Y2=0
cc_201 N_GATE_M1022_g N_A_267_464#_c_259_n 0.0251057f $X=1.26 $Y=2.64 $X2=0
+ $Y2=0
cc_202 GATE N_A_267_464#_c_259_n 0.00172444f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_203 N_GATE_M1022_g N_A_267_464#_c_280_n 0.00147561f $X=1.26 $Y=2.64 $X2=0
+ $Y2=0
cc_204 N_GATE_c_212_n N_A_267_464#_c_270_n 0.00349721f $X=1.26 $Y=0.88 $X2=0
+ $Y2=0
cc_205 GATE N_A_267_464#_c_270_n 0.00250243f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_206 N_GATE_c_215_n N_A_267_464#_c_270_n 0.00130974f $X=1.26 $Y=1.045 $X2=0
+ $Y2=0
cc_207 N_GATE_M1022_g N_A_267_464#_c_271_n 0.0072293f $X=1.26 $Y=2.64 $X2=0
+ $Y2=0
cc_208 N_GATE_c_213_n N_A_267_464#_c_271_n 0.00740982f $X=1.26 $Y=1.385 $X2=0
+ $Y2=0
cc_209 N_GATE_c_212_n N_A_267_464#_c_273_n 0.00458297f $X=1.26 $Y=0.88 $X2=0
+ $Y2=0
cc_210 GATE N_A_267_464#_c_273_n 0.102672f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_211 N_GATE_c_215_n N_A_267_464#_c_273_n 0.00740982f $X=1.26 $Y=1.045 $X2=0
+ $Y2=0
cc_212 N_GATE_M1022_g N_A_49_70#_c_425_n 0.00590121f $X=1.26 $Y=2.64 $X2=0 $Y2=0
cc_213 GATE N_A_49_70#_c_425_n 0.0170432f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_214 N_GATE_M1022_g N_A_49_70#_c_436_n 0.0173951f $X=1.26 $Y=2.64 $X2=0 $Y2=0
cc_215 N_GATE_M1022_g N_A_49_70#_c_426_n 0.0104857f $X=1.26 $Y=2.64 $X2=0 $Y2=0
cc_216 N_GATE_M1022_g N_A_49_70#_c_427_n 0.00294468f $X=1.26 $Y=2.64 $X2=0 $Y2=0
cc_217 N_GATE_c_212_n N_A_414_47#_c_514_n 0.00258531f $X=1.26 $Y=0.88 $X2=0
+ $Y2=0
cc_218 N_GATE_M1022_g N_A_414_47#_c_526_n 0.00165917f $X=1.26 $Y=2.64 $X2=0
+ $Y2=0
cc_219 N_GATE_M1022_g N_VPWR_c_986_n 0.00159208f $X=1.26 $Y=2.64 $X2=0 $Y2=0
cc_220 N_GATE_M1022_g N_VPWR_c_993_n 0.00278223f $X=1.26 $Y=2.64 $X2=0 $Y2=0
cc_221 N_GATE_M1022_g N_VPWR_c_985_n 0.00360368f $X=1.26 $Y=2.64 $X2=0 $Y2=0
cc_222 N_GATE_c_212_n N_VGND_c_1154_n 0.00350603f $X=1.26 $Y=0.88 $X2=0 $Y2=0
cc_223 GATE N_VGND_c_1154_n 0.0100853f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_224 N_GATE_c_215_n N_VGND_c_1154_n 4.53926e-19 $X=1.26 $Y=1.045 $X2=0 $Y2=0
cc_225 N_GATE_c_212_n N_VGND_c_1163_n 0.00449875f $X=1.26 $Y=0.88 $X2=0 $Y2=0
cc_226 N_GATE_c_212_n N_VGND_c_1172_n 0.00513312f $X=1.26 $Y=0.88 $X2=0 $Y2=0
cc_227 GATE N_VGND_c_1172_n 0.00627207f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_228 N_A_267_464#_c_261_n N_A_49_70#_c_417_n 0.00509239f $X=2.41 $Y=1.49 $X2=0
+ $Y2=0
cc_229 N_A_267_464#_c_260_n N_A_49_70#_M1012_g 0.0163409f $X=2.41 $Y=0.765 $X2=0
+ $Y2=0
cc_230 N_A_267_464#_c_261_n N_A_49_70#_M1012_g 0.00498675f $X=2.41 $Y=1.49 $X2=0
+ $Y2=0
cc_231 N_A_267_464#_c_268_n N_A_49_70#_M1012_g 0.01221f $X=3.745 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_267_464#_c_274_n N_A_49_70#_M1012_g 0.00133252f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_233 N_A_267_464#_c_275_n N_A_49_70#_M1012_g 0.0162866f $X=2.41 $Y=0.93 $X2=0
+ $Y2=0
cc_234 N_A_267_464#_M1000_g N_A_49_70#_M1004_g 0.00699574f $X=2.41 $Y=2.665
+ $X2=0 $Y2=0
cc_235 N_A_267_464#_M1020_g N_A_49_70#_M1004_g 0.0483867f $X=3.54 $Y=2.665 $X2=0
+ $Y2=0
cc_236 N_A_267_464#_c_280_n N_A_49_70#_c_425_n 0.0139615f $X=1.63 $Y=2.3 $X2=0
+ $Y2=0
cc_237 N_A_267_464#_c_280_n N_A_49_70#_c_436_n 0.0143208f $X=1.63 $Y=2.3 $X2=0
+ $Y2=0
cc_238 N_A_267_464#_M1022_d N_A_49_70#_c_426_n 0.0035559f $X=1.335 $Y=2.32 $X2=0
+ $Y2=0
cc_239 N_A_267_464#_M1000_g N_A_49_70#_c_426_n 0.0162421f $X=2.41 $Y=2.665 $X2=0
+ $Y2=0
cc_240 N_A_267_464#_c_280_n N_A_49_70#_c_426_n 0.0169481f $X=1.63 $Y=2.3 $X2=0
+ $Y2=0
cc_241 N_A_267_464#_M1000_g N_A_49_70#_c_428_n 0.00600044f $X=2.41 $Y=2.665
+ $X2=0 $Y2=0
cc_242 N_A_267_464#_c_266_n N_A_49_70#_c_420_n 0.00600044f $X=2.41 $Y=1.565
+ $X2=0 $Y2=0
cc_243 N_A_267_464#_c_266_n N_A_49_70#_c_421_n 0.0406487f $X=2.41 $Y=1.565 $X2=0
+ $Y2=0
cc_244 N_A_267_464#_c_267_n N_A_49_70#_c_421_n 0.0483867f $X=3.82 $Y=1.54 $X2=0
+ $Y2=0
cc_245 N_A_267_464#_c_266_n N_A_49_70#_c_422_n 0.00509239f $X=2.41 $Y=1.565
+ $X2=0 $Y2=0
cc_246 N_A_267_464#_c_267_n N_A_49_70#_c_422_n 5.34943e-19 $X=3.82 $Y=1.54 $X2=0
+ $Y2=0
cc_247 N_A_267_464#_c_274_n N_A_414_47#_M1002_s 9.34767e-19 $X=2.41 $Y=0.74
+ $X2=-0.19 $Y2=-0.245
cc_248 N_A_267_464#_M1017_g N_A_414_47#_M1009_g 0.020338f $X=3.82 $Y=0.445 $X2=0
+ $Y2=0
cc_249 N_A_267_464#_c_268_n N_A_414_47#_M1009_g 0.0119368f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_250 N_A_267_464#_c_269_n N_A_414_47#_M1009_g 5.77214e-19 $X=3.83 $Y=1.065
+ $X2=0 $Y2=0
cc_251 N_A_267_464#_M1020_g N_A_414_47#_M1016_g 0.0136861f $X=3.54 $Y=2.665
+ $X2=0 $Y2=0
cc_252 N_A_267_464#_c_260_n N_A_414_47#_c_513_n 0.00431025f $X=2.41 $Y=0.765
+ $X2=0 $Y2=0
cc_253 N_A_267_464#_c_261_n N_A_414_47#_c_513_n 0.00306068f $X=2.41 $Y=1.49
+ $X2=0 $Y2=0
cc_254 N_A_267_464#_c_270_n N_A_414_47#_c_513_n 0.0141964f $X=1.63 $Y=0.532
+ $X2=0 $Y2=0
cc_255 N_A_267_464#_c_273_n N_A_414_47#_c_513_n 0.0379715f $X=1.755 $Y=1.535
+ $X2=0 $Y2=0
cc_256 N_A_267_464#_c_274_n N_A_414_47#_c_513_n 0.0270931f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_257 N_A_267_464#_c_275_n N_A_414_47#_c_513_n 0.00839331f $X=2.41 $Y=0.93
+ $X2=0 $Y2=0
cc_258 N_A_267_464#_c_270_n N_A_414_47#_c_514_n 0.00745055f $X=1.63 $Y=0.532
+ $X2=0 $Y2=0
cc_259 N_A_267_464#_c_260_n N_A_414_47#_c_544_n 0.00265059f $X=2.41 $Y=0.765
+ $X2=0 $Y2=0
cc_260 N_A_267_464#_c_274_n N_A_414_47#_c_544_n 0.00620102f $X=2.41 $Y=0.74
+ $X2=0 $Y2=0
cc_261 N_A_267_464#_c_275_n N_A_414_47#_c_544_n 3.75239e-19 $X=2.41 $Y=0.93
+ $X2=0 $Y2=0
cc_262 N_A_267_464#_c_261_n N_A_414_47#_c_515_n 0.0170042f $X=2.41 $Y=1.49 $X2=0
+ $Y2=0
cc_263 N_A_267_464#_c_268_n N_A_414_47#_c_515_n 0.026537f $X=3.745 $Y=0.74 $X2=0
+ $Y2=0
cc_264 N_A_267_464#_c_275_n N_A_414_47#_c_515_n 0.00220684f $X=2.41 $Y=0.93
+ $X2=0 $Y2=0
cc_265 N_A_267_464#_c_258_n N_A_414_47#_c_516_n 9.63653e-19 $X=2.335 $Y=1.565
+ $X2=0 $Y2=0
cc_266 N_A_267_464#_c_259_n N_A_414_47#_c_516_n 0.00909879f $X=1.965 $Y=1.565
+ $X2=0 $Y2=0
cc_267 N_A_267_464#_c_271_n N_A_414_47#_c_516_n 0.00547332f $X=1.8 $Y=1.655
+ $X2=0 $Y2=0
cc_268 N_A_267_464#_c_273_n N_A_414_47#_c_516_n 0.0136254f $X=1.755 $Y=1.535
+ $X2=0 $Y2=0
cc_269 N_A_267_464#_c_274_n N_A_414_47#_c_516_n 0.0243902f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_270 N_A_267_464#_c_275_n N_A_414_47#_c_516_n 7.97049e-19 $X=2.41 $Y=0.93
+ $X2=0 $Y2=0
cc_271 N_A_267_464#_c_267_n N_A_414_47#_c_517_n 5.41413e-19 $X=3.82 $Y=1.54
+ $X2=0 $Y2=0
cc_272 N_A_267_464#_c_268_n N_A_414_47#_c_517_n 0.0248926f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_273 N_A_267_464#_c_269_n N_A_414_47#_c_517_n 0.0042396f $X=3.83 $Y=1.065
+ $X2=0 $Y2=0
cc_274 N_A_267_464#_c_274_n N_A_414_47#_c_517_n 7.57195e-19 $X=2.41 $Y=0.74
+ $X2=0 $Y2=0
cc_275 N_A_267_464#_c_276_n N_A_414_47#_c_517_n 0.014627f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_276 N_A_267_464#_c_277_n N_A_414_47#_c_517_n 0.00291068f $X=3.91 $Y=1.16
+ $X2=0 $Y2=0
cc_277 N_A_267_464#_c_265_n N_A_414_47#_c_518_n 0.00274103f $X=3.82 $Y=1.465
+ $X2=0 $Y2=0
cc_278 N_A_267_464#_c_267_n N_A_414_47#_c_518_n 0.00948465f $X=3.82 $Y=1.54
+ $X2=0 $Y2=0
cc_279 N_A_267_464#_M1020_g N_A_414_47#_c_523_n 0.0143369f $X=3.54 $Y=2.665
+ $X2=0 $Y2=0
cc_280 N_A_267_464#_M1020_g N_A_414_47#_c_525_n 7.25841e-19 $X=3.54 $Y=2.665
+ $X2=0 $Y2=0
cc_281 N_A_267_464#_c_280_n N_A_414_47#_c_526_n 0.0139209f $X=1.63 $Y=2.3 $X2=0
+ $Y2=0
cc_282 N_A_267_464#_c_258_n N_A_414_47#_c_519_n 0.0113719f $X=2.335 $Y=1.565
+ $X2=0 $Y2=0
cc_283 N_A_267_464#_c_261_n N_A_414_47#_c_519_n 0.00511279f $X=2.41 $Y=1.49
+ $X2=0 $Y2=0
cc_284 N_A_267_464#_M1000_g N_A_414_47#_c_519_n 0.00955934f $X=2.41 $Y=2.665
+ $X2=0 $Y2=0
cc_285 N_A_267_464#_c_280_n N_A_414_47#_c_519_n 0.00997914f $X=1.63 $Y=2.3 $X2=0
+ $Y2=0
cc_286 N_A_267_464#_c_271_n N_A_414_47#_c_519_n 0.045227f $X=1.8 $Y=1.655 $X2=0
+ $Y2=0
cc_287 N_A_267_464#_c_272_n N_A_414_47#_c_519_n 0.00380799f $X=1.8 $Y=1.655
+ $X2=0 $Y2=0
cc_288 N_A_267_464#_c_273_n N_A_414_47#_c_519_n 0.0064102f $X=1.755 $Y=1.535
+ $X2=0 $Y2=0
cc_289 N_A_267_464#_M1017_g N_A_414_47#_c_520_n 0.021138f $X=3.82 $Y=0.445 $X2=0
+ $Y2=0
cc_290 N_A_267_464#_c_267_n N_A_414_47#_c_520_n 0.00467018f $X=3.82 $Y=1.54
+ $X2=0 $Y2=0
cc_291 N_A_267_464#_c_268_n N_A_414_47#_c_520_n 0.0043813f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_292 N_A_267_464#_c_269_n N_A_414_47#_c_520_n 5.8936e-19 $X=3.83 $Y=1.065
+ $X2=0 $Y2=0
cc_293 N_A_267_464#_c_276_n N_A_414_47#_c_520_n 2.39094e-19 $X=3.91 $Y=1.16
+ $X2=0 $Y2=0
cc_294 N_A_267_464#_M1020_g N_A_414_47#_c_528_n 0.0203599f $X=3.54 $Y=2.665
+ $X2=0 $Y2=0
cc_295 N_A_267_464#_c_267_n N_A_414_47#_c_528_n 0.0037305f $X=3.82 $Y=1.54 $X2=0
+ $Y2=0
cc_296 N_A_267_464#_c_277_n N_A_414_47#_c_528_n 0.00287195f $X=3.91 $Y=1.16
+ $X2=0 $Y2=0
cc_297 N_A_267_464#_M1020_g N_A_414_47#_c_529_n 2.99505e-19 $X=3.54 $Y=2.665
+ $X2=0 $Y2=0
cc_298 N_A_267_464#_M1017_g N_A_857_21#_c_644_n 0.0218947f $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_299 N_A_267_464#_c_268_n N_A_857_21#_c_644_n 4.39223e-19 $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_300 N_A_267_464#_c_269_n N_A_857_21#_c_649_n 2.17156e-19 $X=3.83 $Y=1.065
+ $X2=0 $Y2=0
cc_301 N_A_267_464#_M1017_g N_A_857_21#_c_654_n 0.00168987f $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_302 N_A_267_464#_c_265_n N_A_857_21#_c_654_n 0.00602995f $X=3.82 $Y=1.465
+ $X2=0 $Y2=0
cc_303 N_A_267_464#_c_269_n N_A_857_21#_c_654_n 3.10192e-19 $X=3.83 $Y=1.065
+ $X2=0 $Y2=0
cc_304 N_A_267_464#_c_276_n N_A_857_21#_c_654_n 2.55416e-19 $X=3.91 $Y=1.16
+ $X2=0 $Y2=0
cc_305 N_A_267_464#_c_277_n N_A_857_21#_c_654_n 0.0140616f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_306 N_A_267_464#_M1017_g N_A_671_47#_c_837_n 0.00945998f $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_307 N_A_267_464#_c_268_n N_A_671_47#_c_837_n 0.0310228f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_308 N_A_267_464#_c_276_n N_A_671_47#_c_837_n 0.00394891f $X=3.91 $Y=1.16
+ $X2=0 $Y2=0
cc_309 N_A_267_464#_c_277_n N_A_671_47#_c_837_n 0.00274166f $X=3.91 $Y=1.16
+ $X2=0 $Y2=0
cc_310 N_A_267_464#_M1020_g N_A_671_47#_c_835_n 0.0159106f $X=3.54 $Y=2.665
+ $X2=0 $Y2=0
cc_311 N_A_267_464#_c_267_n N_A_671_47#_c_826_n 0.00860187f $X=3.82 $Y=1.54
+ $X2=0 $Y2=0
cc_312 N_A_267_464#_c_268_n N_A_671_47#_c_826_n 4.91022e-19 $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_313 N_A_267_464#_c_276_n N_A_671_47#_c_826_n 0.0236141f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_314 N_A_267_464#_c_277_n N_A_671_47#_c_826_n 0.00169953f $X=3.91 $Y=1.16
+ $X2=0 $Y2=0
cc_315 N_A_267_464#_M1020_g N_A_671_47#_c_846_n 0.0010673f $X=3.54 $Y=2.665
+ $X2=0 $Y2=0
cc_316 N_A_267_464#_c_267_n N_A_671_47#_c_846_n 0.00871468f $X=3.82 $Y=1.54
+ $X2=0 $Y2=0
cc_317 N_A_267_464#_c_268_n N_A_671_47#_c_846_n 0.00484635f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_318 N_A_267_464#_M1017_g N_A_671_47#_c_827_n 0.00386958f $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_319 N_A_267_464#_c_268_n N_A_671_47#_c_827_n 0.0059341f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_320 N_A_267_464#_M1017_g N_A_671_47#_c_828_n 3.65583e-19 $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_321 N_A_267_464#_c_269_n N_A_671_47#_c_828_n 0.00764797f $X=3.83 $Y=1.065
+ $X2=0 $Y2=0
cc_322 N_A_267_464#_c_276_n N_A_671_47#_c_828_n 0.0172132f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_323 N_A_267_464#_c_277_n N_A_671_47#_c_828_n 0.0015645f $X=3.91 $Y=1.16 $X2=0
+ $Y2=0
cc_324 N_A_267_464#_M1020_g N_A_671_47#_c_855_n 0.005142f $X=3.54 $Y=2.665 $X2=0
+ $Y2=0
cc_325 N_A_267_464#_M1017_g N_A_671_47#_c_831_n 6.20052e-19 $X=3.82 $Y=0.445
+ $X2=0 $Y2=0
cc_326 N_A_267_464#_c_268_n N_A_671_47#_c_831_n 0.00881515f $X=3.745 $Y=0.74
+ $X2=0 $Y2=0
cc_327 N_A_267_464#_c_269_n N_A_671_47#_c_831_n 0.0054701f $X=3.83 $Y=1.065
+ $X2=0 $Y2=0
cc_328 N_A_267_464#_c_265_n N_A_671_47#_c_832_n 0.00352373f $X=3.82 $Y=1.465
+ $X2=0 $Y2=0
cc_329 N_A_267_464#_c_277_n N_A_671_47#_c_832_n 2.79863e-19 $X=3.91 $Y=1.16
+ $X2=0 $Y2=0
cc_330 N_A_267_464#_M1000_g N_VPWR_c_987_n 0.00197993f $X=2.41 $Y=2.665 $X2=0
+ $Y2=0
cc_331 N_A_267_464#_M1000_g N_VPWR_c_993_n 0.0029147f $X=2.41 $Y=2.665 $X2=0
+ $Y2=0
cc_332 N_A_267_464#_M1020_g N_VPWR_c_995_n 0.0029147f $X=3.54 $Y=2.665 $X2=0
+ $Y2=0
cc_333 N_A_267_464#_M1000_g N_VPWR_c_985_n 0.00443422f $X=2.41 $Y=2.665 $X2=0
+ $Y2=0
cc_334 N_A_267_464#_M1020_g N_VPWR_c_985_n 0.00425026f $X=3.54 $Y=2.665 $X2=0
+ $Y2=0
cc_335 N_A_267_464#_c_274_n N_VGND_M1002_d 0.00135161f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_336 N_A_267_464#_c_260_n N_VGND_c_1155_n 0.00432564f $X=2.41 $Y=0.765 $X2=0
+ $Y2=0
cc_337 N_A_267_464#_c_268_n N_VGND_c_1155_n 0.0202264f $X=3.745 $Y=0.74 $X2=0
+ $Y2=0
cc_338 N_A_267_464#_c_274_n N_VGND_c_1155_n 0.00263585f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_339 N_A_267_464#_c_260_n N_VGND_c_1163_n 0.00417244f $X=2.41 $Y=0.765 $X2=0
+ $Y2=0
cc_340 N_A_267_464#_c_270_n N_VGND_c_1163_n 0.0122448f $X=1.63 $Y=0.532 $X2=0
+ $Y2=0
cc_341 N_A_267_464#_c_274_n N_VGND_c_1163_n 0.00301785f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_342 N_A_267_464#_M1017_g N_VGND_c_1164_n 0.00359964f $X=3.82 $Y=0.445 $X2=0
+ $Y2=0
cc_343 N_A_267_464#_c_268_n N_VGND_c_1164_n 0.00943729f $X=3.745 $Y=0.74 $X2=0
+ $Y2=0
cc_344 N_A_267_464#_c_260_n N_VGND_c_1172_n 0.0072946f $X=2.41 $Y=0.765 $X2=0
+ $Y2=0
cc_345 N_A_267_464#_M1017_g N_VGND_c_1172_n 0.00590845f $X=3.82 $Y=0.445 $X2=0
+ $Y2=0
cc_346 N_A_267_464#_c_268_n N_VGND_c_1172_n 0.0165312f $X=3.745 $Y=0.74 $X2=0
+ $Y2=0
cc_347 N_A_267_464#_c_270_n N_VGND_c_1172_n 0.0130827f $X=1.63 $Y=0.532 $X2=0
+ $Y2=0
cc_348 N_A_267_464#_c_274_n N_VGND_c_1172_n 0.00499201f $X=2.41 $Y=0.74 $X2=0
+ $Y2=0
cc_349 N_A_267_464#_c_268_n A_779_47# 2.00183e-19 $X=3.745 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_350 N_A_49_70#_c_426_n N_A_414_47#_M1000_s 0.00258276f $X=2.495 $Y=2.99 $X2=0
+ $Y2=0
cc_351 N_A_49_70#_M1012_g N_A_414_47#_M1009_g 0.0363025f $X=2.92 $Y=0.445 $X2=0
+ $Y2=0
cc_352 N_A_49_70#_c_417_n N_A_414_47#_c_515_n 0.00470675f $X=2.905 $Y=1.315
+ $X2=0 $Y2=0
cc_353 N_A_49_70#_M1012_g N_A_414_47#_c_515_n 0.00418676f $X=2.92 $Y=0.445 $X2=0
+ $Y2=0
cc_354 N_A_49_70#_c_420_n N_A_414_47#_c_515_n 0.0422498f $X=2.86 $Y=1.66 $X2=0
+ $Y2=0
cc_355 N_A_49_70#_c_421_n N_A_414_47#_c_515_n 0.0118457f $X=2.86 $Y=1.66 $X2=0
+ $Y2=0
cc_356 N_A_49_70#_c_422_n N_A_414_47#_c_515_n 0.00493111f $X=2.975 $Y=1.495
+ $X2=0 $Y2=0
cc_357 N_A_49_70#_M1012_g N_A_414_47#_c_517_n 0.00125671f $X=2.92 $Y=0.445 $X2=0
+ $Y2=0
cc_358 N_A_49_70#_M1004_g N_A_414_47#_c_518_n 0.0139532f $X=3.18 $Y=2.665 $X2=0
+ $Y2=0
cc_359 N_A_49_70#_c_428_n N_A_414_47#_c_518_n 0.00507115f $X=2.58 $Y=2.905 $X2=0
+ $Y2=0
cc_360 N_A_49_70#_c_420_n N_A_414_47#_c_518_n 0.0446709f $X=2.86 $Y=1.66 $X2=0
+ $Y2=0
cc_361 N_A_49_70#_c_421_n N_A_414_47#_c_518_n 0.0174135f $X=2.86 $Y=1.66 $X2=0
+ $Y2=0
cc_362 N_A_49_70#_c_422_n N_A_414_47#_c_518_n 0.00397617f $X=2.975 $Y=1.495
+ $X2=0 $Y2=0
cc_363 N_A_49_70#_M1004_g N_A_414_47#_c_524_n 0.00435293f $X=3.18 $Y=2.665 $X2=0
+ $Y2=0
cc_364 N_A_49_70#_c_426_n N_A_414_47#_c_526_n 0.018445f $X=2.495 $Y=2.99 $X2=0
+ $Y2=0
cc_365 N_A_49_70#_c_420_n N_A_414_47#_c_519_n 0.0651598f $X=2.86 $Y=1.66 $X2=0
+ $Y2=0
cc_366 N_A_49_70#_c_421_n N_A_414_47#_c_519_n 2.85733e-19 $X=2.86 $Y=1.66 $X2=0
+ $Y2=0
cc_367 N_A_49_70#_c_417_n N_A_414_47#_c_520_n 0.0363025f $X=2.905 $Y=1.315 $X2=0
+ $Y2=0
cc_368 N_A_49_70#_c_421_n N_A_414_47#_c_520_n 0.00278165f $X=2.86 $Y=1.66 $X2=0
+ $Y2=0
cc_369 N_A_49_70#_c_421_n N_A_671_47#_c_835_n 6.44795e-19 $X=2.86 $Y=1.66 $X2=0
+ $Y2=0
cc_370 N_A_49_70#_M1004_g N_A_671_47#_c_855_n 2.87829e-19 $X=3.18 $Y=2.665 $X2=0
+ $Y2=0
cc_371 N_A_49_70#_c_425_n N_VPWR_M1006_d 0.00669513f $X=1.065 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_372 N_A_49_70#_c_436_n N_VPWR_M1006_d 0.00491256f $X=1.15 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_373 N_A_49_70#_c_427_n N_VPWR_M1006_d 5.2468e-19 $X=1.235 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_374 N_A_49_70#_c_426_n N_VPWR_M1000_d 7.72915e-19 $X=2.495 $Y=2.99 $X2=0
+ $Y2=0
cc_375 N_A_49_70#_c_428_n N_VPWR_M1000_d 0.00776157f $X=2.58 $Y=2.905 $X2=0
+ $Y2=0
cc_376 N_A_49_70#_c_425_n N_VPWR_c_986_n 0.015111f $X=1.065 $Y=2.385 $X2=0 $Y2=0
cc_377 N_A_49_70#_c_436_n N_VPWR_c_986_n 0.0197836f $X=1.15 $Y=2.905 $X2=0 $Y2=0
cc_378 N_A_49_70#_c_427_n N_VPWR_c_986_n 0.0145681f $X=1.235 $Y=2.99 $X2=0 $Y2=0
cc_379 N_A_49_70#_c_429_n N_VPWR_c_986_n 0.0122299f $X=0.37 $Y=2.465 $X2=0 $Y2=0
cc_380 N_A_49_70#_M1004_g N_VPWR_c_987_n 0.00383052f $X=3.18 $Y=2.665 $X2=0
+ $Y2=0
cc_381 N_A_49_70#_c_426_n N_VPWR_c_987_n 0.0142667f $X=2.495 $Y=2.99 $X2=0 $Y2=0
cc_382 N_A_49_70#_c_428_n N_VPWR_c_987_n 0.0419022f $X=2.58 $Y=2.905 $X2=0 $Y2=0
cc_383 N_A_49_70#_c_420_n N_VPWR_c_987_n 0.0166691f $X=2.86 $Y=1.66 $X2=0 $Y2=0
cc_384 N_A_49_70#_c_421_n N_VPWR_c_987_n 0.00195037f $X=2.86 $Y=1.66 $X2=0 $Y2=0
cc_385 N_A_49_70#_c_426_n N_VPWR_c_993_n 0.0925345f $X=2.495 $Y=2.99 $X2=0 $Y2=0
cc_386 N_A_49_70#_c_427_n N_VPWR_c_993_n 0.012011f $X=1.235 $Y=2.99 $X2=0 $Y2=0
cc_387 N_A_49_70#_M1004_g N_VPWR_c_995_n 0.00418602f $X=3.18 $Y=2.665 $X2=0
+ $Y2=0
cc_388 N_A_49_70#_c_429_n N_VPWR_c_999_n 0.0114959f $X=0.37 $Y=2.465 $X2=0 $Y2=0
cc_389 N_A_49_70#_M1004_g N_VPWR_c_985_n 0.00776521f $X=3.18 $Y=2.665 $X2=0
+ $Y2=0
cc_390 N_A_49_70#_c_425_n N_VPWR_c_985_n 0.0113549f $X=1.065 $Y=2.385 $X2=0
+ $Y2=0
cc_391 N_A_49_70#_c_426_n N_VPWR_c_985_n 0.052832f $X=2.495 $Y=2.99 $X2=0 $Y2=0
cc_392 N_A_49_70#_c_427_n N_VPWR_c_985_n 0.00638043f $X=1.235 $Y=2.99 $X2=0
+ $Y2=0
cc_393 N_A_49_70#_c_429_n N_VPWR_c_985_n 0.00983801f $X=0.37 $Y=2.465 $X2=0
+ $Y2=0
cc_394 N_A_49_70#_M1012_g N_VGND_c_1155_n 0.00957712f $X=2.92 $Y=0.445 $X2=0
+ $Y2=0
cc_395 N_A_49_70#_c_419_n N_VGND_c_1161_n 0.00911408f $X=0.37 $Y=0.56 $X2=0
+ $Y2=0
cc_396 N_A_49_70#_M1012_g N_VGND_c_1164_n 0.00355956f $X=2.92 $Y=0.445 $X2=0
+ $Y2=0
cc_397 N_A_49_70#_M1012_g N_VGND_c_1172_n 0.00406467f $X=2.92 $Y=0.445 $X2=0
+ $Y2=0
cc_398 N_A_49_70#_c_419_n N_VGND_c_1172_n 0.00889983f $X=0.37 $Y=0.56 $X2=0
+ $Y2=0
cc_399 N_A_414_47#_M1016_g N_A_857_21#_M1010_g 0.0381454f $X=4.065 $Y=2.555
+ $X2=0 $Y2=0
cc_400 N_A_414_47#_c_523_n N_A_857_21#_M1010_g 2.74173e-19 $X=4.04 $Y=2.98 $X2=0
+ $Y2=0
cc_401 N_A_414_47#_c_525_n N_A_857_21#_M1010_g 0.0100652f $X=4.125 $Y=2.885
+ $X2=0 $Y2=0
cc_402 N_A_414_47#_c_525_n N_A_857_21#_c_661_n 0.00778881f $X=4.125 $Y=2.885
+ $X2=0 $Y2=0
cc_403 N_A_414_47#_c_528_n N_A_857_21#_c_661_n 3.57016e-19 $X=3.99 $Y=2.02 $X2=0
+ $Y2=0
cc_404 N_A_414_47#_c_529_n N_A_857_21#_c_661_n 0.0259018f $X=4.125 $Y=2.02 $X2=0
+ $Y2=0
cc_405 N_A_414_47#_c_528_n N_A_857_21#_c_662_n 0.0206007f $X=3.99 $Y=2.02 $X2=0
+ $Y2=0
cc_406 N_A_414_47#_c_529_n N_A_857_21#_c_662_n 0.00189557f $X=4.125 $Y=2.02
+ $X2=0 $Y2=0
cc_407 N_A_414_47#_c_525_n N_A_857_21#_c_683_n 0.0134342f $X=4.125 $Y=2.885
+ $X2=0 $Y2=0
cc_408 N_A_414_47#_c_523_n N_A_671_47#_M1020_d 0.00258609f $X=4.04 $Y=2.98 $X2=0
+ $Y2=0
cc_409 N_A_414_47#_M1009_g N_A_671_47#_c_837_n 0.00339307f $X=3.28 $Y=0.445
+ $X2=0 $Y2=0
cc_410 N_A_414_47#_M1016_g N_A_671_47#_c_835_n 0.00135725f $X=4.065 $Y=2.555
+ $X2=0 $Y2=0
cc_411 N_A_414_47#_c_518_n N_A_671_47#_c_835_n 0.0506113f $X=3.29 $Y=2.885 $X2=0
+ $Y2=0
cc_412 N_A_414_47#_c_525_n N_A_671_47#_c_835_n 0.0089648f $X=4.125 $Y=2.885
+ $X2=0 $Y2=0
cc_413 N_A_414_47#_c_528_n N_A_671_47#_c_835_n 0.00201101f $X=3.99 $Y=2.02 $X2=0
+ $Y2=0
cc_414 N_A_414_47#_c_529_n N_A_671_47#_c_835_n 0.0246834f $X=4.125 $Y=2.02 $X2=0
+ $Y2=0
cc_415 N_A_414_47#_c_528_n N_A_671_47#_c_826_n 0.00508165f $X=3.99 $Y=2.02 $X2=0
+ $Y2=0
cc_416 N_A_414_47#_c_529_n N_A_671_47#_c_826_n 0.0204364f $X=4.125 $Y=2.02 $X2=0
+ $Y2=0
cc_417 N_A_414_47#_c_518_n N_A_671_47#_c_846_n 0.0129658f $X=3.29 $Y=2.885 $X2=0
+ $Y2=0
cc_418 N_A_414_47#_M1016_g N_A_671_47#_c_855_n 0.00247873f $X=4.065 $Y=2.555
+ $X2=0 $Y2=0
cc_419 N_A_414_47#_c_518_n N_A_671_47#_c_855_n 0.0231987f $X=3.29 $Y=2.885 $X2=0
+ $Y2=0
cc_420 N_A_414_47#_c_523_n N_A_671_47#_c_855_n 0.0184108f $X=4.04 $Y=2.98 $X2=0
+ $Y2=0
cc_421 N_A_414_47#_c_525_n N_A_671_47#_c_855_n 0.0243014f $X=4.125 $Y=2.885
+ $X2=0 $Y2=0
cc_422 N_A_414_47#_c_528_n N_A_671_47#_c_855_n 0.00176126f $X=3.99 $Y=2.02 $X2=0
+ $Y2=0
cc_423 N_A_414_47#_c_518_n N_VPWR_c_987_n 0.0390846f $X=3.29 $Y=2.885 $X2=0
+ $Y2=0
cc_424 N_A_414_47#_c_524_n N_VPWR_c_987_n 0.0152264f $X=3.375 $Y=2.98 $X2=0
+ $Y2=0
cc_425 N_A_414_47#_M1016_g N_VPWR_c_995_n 6.25023e-19 $X=4.065 $Y=2.555 $X2=0
+ $Y2=0
cc_426 N_A_414_47#_c_523_n N_VPWR_c_995_n 0.0548529f $X=4.04 $Y=2.98 $X2=0 $Y2=0
cc_427 N_A_414_47#_c_524_n N_VPWR_c_995_n 0.0119421f $X=3.375 $Y=2.98 $X2=0
+ $Y2=0
cc_428 N_A_414_47#_c_523_n N_VPWR_c_985_n 0.0309798f $X=4.04 $Y=2.98 $X2=0 $Y2=0
cc_429 N_A_414_47#_c_524_n N_VPWR_c_985_n 0.00637045f $X=3.375 $Y=2.98 $X2=0
+ $Y2=0
cc_430 N_A_414_47#_c_518_n A_651_469# 0.00538426f $X=3.29 $Y=2.885 $X2=-0.19
+ $Y2=-0.245
cc_431 N_A_414_47#_c_523_n A_651_469# 0.00123754f $X=4.04 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_432 N_A_414_47#_c_525_n A_828_469# 0.00445924f $X=4.125 $Y=2.885 $X2=-0.19
+ $Y2=-0.245
cc_433 N_A_414_47#_M1009_g N_VGND_c_1155_n 0.00192097f $X=3.28 $Y=0.445 $X2=0
+ $Y2=0
cc_434 N_A_414_47#_c_514_n N_VGND_c_1163_n 0.0102395f $X=2.065 $Y=0.385 $X2=0
+ $Y2=0
cc_435 N_A_414_47#_c_544_n N_VGND_c_1163_n 0.0144341f $X=2.195 $Y=0.39 $X2=0
+ $Y2=0
cc_436 N_A_414_47#_M1009_g N_VGND_c_1164_n 0.00428022f $X=3.28 $Y=0.445 $X2=0
+ $Y2=0
cc_437 N_A_414_47#_M1002_s N_VGND_c_1172_n 0.00215649f $X=2.07 $Y=0.235 $X2=0
+ $Y2=0
cc_438 N_A_414_47#_M1009_g N_VGND_c_1172_n 0.00619329f $X=3.28 $Y=0.445 $X2=0
+ $Y2=0
cc_439 N_A_414_47#_c_514_n N_VGND_c_1172_n 0.00651219f $X=2.065 $Y=0.385 $X2=0
+ $Y2=0
cc_440 N_A_414_47#_c_544_n N_VGND_c_1172_n 0.0107418f $X=2.195 $Y=0.39 $X2=0
+ $Y2=0
cc_441 N_A_857_21#_c_649_n N_A_671_47#_c_821_n 0.0259756f $X=4.44 $Y=0.84 $X2=0
+ $Y2=0
cc_442 N_A_857_21#_c_650_n N_A_671_47#_c_821_n 0.00766216f $X=5.125 $Y=0.525
+ $X2=0 $Y2=0
cc_443 N_A_857_21#_c_686_p N_A_671_47#_c_821_n 0.0025711f $X=5.23 $Y=0.955 $X2=0
+ $Y2=0
cc_444 N_A_857_21#_c_650_n N_A_671_47#_c_822_n 0.00361283f $X=5.125 $Y=0.525
+ $X2=0 $Y2=0
cc_445 N_A_857_21#_c_644_n N_A_671_47#_c_823_n 0.0161376f $X=4.36 $Y=0.765 $X2=0
+ $Y2=0
cc_446 N_A_857_21#_c_689_p N_A_671_47#_c_824_n 2.65883e-19 $X=6.055 $Y=0.955
+ $X2=0 $Y2=0
cc_447 N_A_857_21#_c_686_p N_A_671_47#_c_824_n 0.00450469f $X=5.23 $Y=0.955
+ $X2=0 $Y2=0
cc_448 N_A_857_21#_c_689_p N_A_671_47#_c_825_n 0.0135066f $X=6.055 $Y=0.955
+ $X2=0 $Y2=0
cc_449 N_A_857_21#_c_661_n N_A_671_47#_c_834_n 0.00384418f $X=4.53 $Y=2.02 $X2=0
+ $Y2=0
cc_450 N_A_857_21#_c_662_n N_A_671_47#_c_834_n 0.00613116f $X=4.53 $Y=2.02 $X2=0
+ $Y2=0
cc_451 N_A_857_21#_c_663_n N_A_671_47#_c_834_n 0.0158536f $X=5.46 $Y=2.375 $X2=0
+ $Y2=0
cc_452 N_A_857_21#_c_654_n N_A_671_47#_c_835_n 0.00440452f $X=4.53 $Y=1.855
+ $X2=0 $Y2=0
cc_453 N_A_857_21#_c_644_n N_A_671_47#_c_827_n 0.00287104f $X=4.36 $Y=0.765
+ $X2=0 $Y2=0
cc_454 N_A_857_21#_c_649_n N_A_671_47#_c_828_n 0.00313888f $X=4.44 $Y=0.84 $X2=0
+ $Y2=0
cc_455 N_A_857_21#_c_686_p N_A_671_47#_c_828_n 0.00425805f $X=5.23 $Y=0.955
+ $X2=0 $Y2=0
cc_456 N_A_857_21#_c_654_n N_A_671_47#_c_828_n 0.0108271f $X=4.53 $Y=1.855 $X2=0
+ $Y2=0
cc_457 N_A_857_21#_c_661_n N_A_671_47#_c_829_n 0.0186675f $X=4.53 $Y=2.02 $X2=0
+ $Y2=0
cc_458 N_A_857_21#_c_662_n N_A_671_47#_c_829_n 0.00127867f $X=4.53 $Y=2.02 $X2=0
+ $Y2=0
cc_459 N_A_857_21#_c_663_n N_A_671_47#_c_829_n 0.00981764f $X=5.46 $Y=2.375
+ $X2=0 $Y2=0
cc_460 N_A_857_21#_c_686_p N_A_671_47#_c_829_n 0.00196596f $X=5.23 $Y=0.955
+ $X2=0 $Y2=0
cc_461 N_A_857_21#_c_654_n N_A_671_47#_c_829_n 0.0111425f $X=4.53 $Y=1.855 $X2=0
+ $Y2=0
cc_462 N_A_857_21#_c_663_n N_A_671_47#_c_830_n 0.00987099f $X=5.46 $Y=2.375
+ $X2=0 $Y2=0
cc_463 N_A_857_21#_c_686_p N_A_671_47#_c_830_n 7.95229e-19 $X=5.23 $Y=0.955
+ $X2=0 $Y2=0
cc_464 N_A_857_21#_c_654_n N_A_671_47#_c_830_n 0.0246756f $X=4.53 $Y=1.855 $X2=0
+ $Y2=0
cc_465 N_A_857_21#_c_644_n N_A_671_47#_c_831_n 0.00496249f $X=4.36 $Y=0.765
+ $X2=0 $Y2=0
cc_466 N_A_857_21#_c_649_n N_A_671_47#_c_831_n 0.00550064f $X=4.44 $Y=0.84 $X2=0
+ $Y2=0
cc_467 N_A_857_21#_c_650_n N_A_671_47#_c_831_n 0.00400505f $X=5.125 $Y=0.525
+ $X2=0 $Y2=0
cc_468 N_A_857_21#_c_686_p N_A_671_47#_c_831_n 7.40577e-19 $X=5.23 $Y=0.955
+ $X2=0 $Y2=0
cc_469 N_A_857_21#_c_661_n N_A_671_47#_c_832_n 0.00307618f $X=4.53 $Y=2.02 $X2=0
+ $Y2=0
cc_470 N_A_857_21#_c_654_n N_A_671_47#_c_832_n 0.00806147f $X=4.53 $Y=1.855
+ $X2=0 $Y2=0
cc_471 N_A_857_21#_c_714_p N_RESET_B_M1007_g 0.0133444f $X=6.055 $Y=2.375 $X2=0
+ $Y2=0
cc_472 N_A_857_21#_c_652_n N_RESET_B_M1007_g 0.00490576f $X=6.14 $Y=2.29 $X2=0
+ $Y2=0
cc_473 N_A_857_21#_c_655_n N_RESET_B_M1007_g 0.0381315f $X=7.565 $Y=1.525 $X2=0
+ $Y2=0
cc_474 N_A_857_21#_M1014_d RESET_B 0.001837f $X=5.415 $Y=1.835 $X2=0 $Y2=0
cc_475 N_A_857_21#_c_661_n RESET_B 0.00706929f $X=4.53 $Y=2.02 $X2=0 $Y2=0
cc_476 N_A_857_21#_c_662_n RESET_B 0.00104042f $X=4.53 $Y=2.02 $X2=0 $Y2=0
cc_477 N_A_857_21#_c_663_n RESET_B 0.0075073f $X=5.46 $Y=2.375 $X2=0 $Y2=0
cc_478 N_A_857_21#_c_689_p RESET_B 0.0416126f $X=6.055 $Y=0.955 $X2=0 $Y2=0
cc_479 N_A_857_21#_c_714_p RESET_B 0.0113922f $X=6.055 $Y=2.375 $X2=0 $Y2=0
cc_480 N_A_857_21#_c_651_n RESET_B 0.015246f $X=6.142 $Y=1.405 $X2=0 $Y2=0
cc_481 N_A_857_21#_c_652_n RESET_B 0.0314981f $X=6.14 $Y=2.29 $X2=0 $Y2=0
cc_482 N_A_857_21#_c_725_p RESET_B 0.0149669f $X=5.56 $Y=2.375 $X2=0 $Y2=0
cc_483 N_A_857_21#_c_653_n RESET_B 0.0148938f $X=6.142 $Y=1.49 $X2=0 $Y2=0
cc_484 N_A_857_21#_c_655_n RESET_B 0.00104582f $X=7.565 $Y=1.525 $X2=0 $Y2=0
cc_485 N_A_857_21#_c_645_n N_RESET_B_c_938_n 4.66546e-19 $X=6.28 $Y=1.325 $X2=0
+ $Y2=0
cc_486 N_A_857_21#_c_689_p N_RESET_B_c_938_n 7.00203e-19 $X=6.055 $Y=0.955 $X2=0
+ $Y2=0
cc_487 N_A_857_21#_c_714_p N_RESET_B_c_938_n 0.00154058f $X=6.055 $Y=2.375 $X2=0
+ $Y2=0
cc_488 N_A_857_21#_c_651_n N_RESET_B_c_938_n 5.51765e-19 $X=6.142 $Y=1.405 $X2=0
+ $Y2=0
cc_489 N_A_857_21#_c_652_n N_RESET_B_c_938_n 4.22693e-19 $X=6.14 $Y=2.29 $X2=0
+ $Y2=0
cc_490 N_A_857_21#_c_653_n N_RESET_B_c_938_n 0.00120117f $X=6.142 $Y=1.49 $X2=0
+ $Y2=0
cc_491 N_A_857_21#_c_655_n N_RESET_B_c_938_n 0.0199142f $X=7.565 $Y=1.525 $X2=0
+ $Y2=0
cc_492 N_A_857_21#_c_645_n N_RESET_B_c_939_n 0.02987f $X=6.28 $Y=1.325 $X2=0
+ $Y2=0
cc_493 N_A_857_21#_c_689_p N_RESET_B_c_939_n 0.0156563f $X=6.055 $Y=0.955 $X2=0
+ $Y2=0
cc_494 N_A_857_21#_c_651_n N_RESET_B_c_939_n 0.0043224f $X=6.142 $Y=1.405 $X2=0
+ $Y2=0
cc_495 N_A_857_21#_c_663_n N_VPWR_M1010_d 0.0187028f $X=5.46 $Y=2.375 $X2=0
+ $Y2=0
cc_496 N_A_857_21#_c_683_n N_VPWR_M1010_d 0.00542699f $X=4.695 $Y=2.375 $X2=0
+ $Y2=0
cc_497 N_A_857_21#_c_714_p N_VPWR_M1007_d 0.00727695f $X=6.055 $Y=2.375 $X2=0
+ $Y2=0
cc_498 N_A_857_21#_c_652_n N_VPWR_M1007_d 0.00443626f $X=6.14 $Y=2.29 $X2=0
+ $Y2=0
cc_499 N_A_857_21#_M1010_g N_VPWR_c_988_n 0.00735647f $X=4.44 $Y=2.555 $X2=0
+ $Y2=0
cc_500 N_A_857_21#_c_663_n N_VPWR_c_988_n 0.0218816f $X=5.46 $Y=2.375 $X2=0
+ $Y2=0
cc_501 N_A_857_21#_c_657_n N_VPWR_c_989_n 0.00250495f $X=6.275 $Y=1.725 $X2=0
+ $Y2=0
cc_502 N_A_857_21#_c_714_p N_VPWR_c_989_n 0.0203005f $X=6.055 $Y=2.375 $X2=0
+ $Y2=0
cc_503 N_A_857_21#_c_657_n N_VPWR_c_990_n 7.48224e-19 $X=6.275 $Y=1.725 $X2=0
+ $Y2=0
cc_504 N_A_857_21#_c_658_n N_VPWR_c_990_n 0.0146036f $X=6.705 $Y=1.725 $X2=0
+ $Y2=0
cc_505 N_A_857_21#_c_659_n N_VPWR_c_990_n 0.0145005f $X=7.135 $Y=1.725 $X2=0
+ $Y2=0
cc_506 N_A_857_21#_c_660_n N_VPWR_c_990_n 7.3e-19 $X=7.565 $Y=1.725 $X2=0 $Y2=0
cc_507 N_A_857_21#_c_659_n N_VPWR_c_992_n 7.3e-19 $X=7.135 $Y=1.725 $X2=0 $Y2=0
cc_508 N_A_857_21#_c_660_n N_VPWR_c_992_n 0.0156867f $X=7.565 $Y=1.725 $X2=0
+ $Y2=0
cc_509 N_A_857_21#_M1010_g N_VPWR_c_995_n 0.00448383f $X=4.44 $Y=2.555 $X2=0
+ $Y2=0
cc_510 N_A_857_21#_c_753_p N_VPWR_c_996_n 0.0128073f $X=5.555 $Y=2.465 $X2=0
+ $Y2=0
cc_511 N_A_857_21#_c_657_n N_VPWR_c_997_n 0.00585385f $X=6.275 $Y=1.725 $X2=0
+ $Y2=0
cc_512 N_A_857_21#_c_658_n N_VPWR_c_997_n 0.00486043f $X=6.705 $Y=1.725 $X2=0
+ $Y2=0
cc_513 N_A_857_21#_c_659_n N_VPWR_c_998_n 0.00486043f $X=7.135 $Y=1.725 $X2=0
+ $Y2=0
cc_514 N_A_857_21#_c_660_n N_VPWR_c_998_n 0.00486043f $X=7.565 $Y=1.725 $X2=0
+ $Y2=0
cc_515 N_A_857_21#_M1014_d N_VPWR_c_985_n 0.00501859f $X=5.415 $Y=1.835 $X2=0
+ $Y2=0
cc_516 N_A_857_21#_M1010_g N_VPWR_c_985_n 0.00486331f $X=4.44 $Y=2.555 $X2=0
+ $Y2=0
cc_517 N_A_857_21#_c_657_n N_VPWR_c_985_n 0.0108678f $X=6.275 $Y=1.725 $X2=0
+ $Y2=0
cc_518 N_A_857_21#_c_658_n N_VPWR_c_985_n 0.00824727f $X=6.705 $Y=1.725 $X2=0
+ $Y2=0
cc_519 N_A_857_21#_c_659_n N_VPWR_c_985_n 0.00824727f $X=7.135 $Y=1.725 $X2=0
+ $Y2=0
cc_520 N_A_857_21#_c_660_n N_VPWR_c_985_n 0.00824727f $X=7.565 $Y=1.725 $X2=0
+ $Y2=0
cc_521 N_A_857_21#_c_753_p N_VPWR_c_985_n 0.00769778f $X=5.555 $Y=2.465 $X2=0
+ $Y2=0
cc_522 N_A_857_21#_c_645_n N_Q_c_1092_n 7.57727e-19 $X=6.28 $Y=1.325 $X2=0 $Y2=0
cc_523 N_A_857_21#_c_646_n N_Q_c_1092_n 8.15613e-19 $X=6.71 $Y=1.325 $X2=0 $Y2=0
cc_524 N_A_857_21#_c_658_n N_Q_c_1098_n 0.0130971f $X=6.705 $Y=1.725 $X2=0 $Y2=0
cc_525 N_A_857_21#_c_659_n N_Q_c_1098_n 0.0136555f $X=7.135 $Y=1.725 $X2=0 $Y2=0
cc_526 N_A_857_21#_c_769_p N_Q_c_1098_n 0.0411721f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_527 N_A_857_21#_c_655_n N_Q_c_1098_n 0.00280751f $X=7.565 $Y=1.525 $X2=0
+ $Y2=0
cc_528 N_A_857_21#_c_657_n N_Q_c_1099_n 7.38449e-19 $X=6.275 $Y=1.725 $X2=0
+ $Y2=0
cc_529 N_A_857_21#_c_652_n N_Q_c_1099_n 0.00993784f $X=6.14 $Y=2.29 $X2=0 $Y2=0
cc_530 N_A_857_21#_c_769_p N_Q_c_1099_n 0.0153303f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_531 N_A_857_21#_c_655_n N_Q_c_1099_n 0.00292686f $X=7.565 $Y=1.525 $X2=0
+ $Y2=0
cc_532 N_A_857_21#_c_646_n N_Q_c_1093_n 0.0132586f $X=6.71 $Y=1.325 $X2=0 $Y2=0
cc_533 N_A_857_21#_c_647_n N_Q_c_1093_n 0.01372f $X=7.14 $Y=1.325 $X2=0 $Y2=0
cc_534 N_A_857_21#_c_769_p N_Q_c_1093_n 0.0383296f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_535 N_A_857_21#_c_655_n N_Q_c_1093_n 0.00258025f $X=7.565 $Y=1.525 $X2=0
+ $Y2=0
cc_536 N_A_857_21#_c_645_n N_Q_c_1094_n 2.43521e-19 $X=6.28 $Y=1.325 $X2=0 $Y2=0
cc_537 N_A_857_21#_c_651_n N_Q_c_1094_n 0.00716655f $X=6.142 $Y=1.405 $X2=0
+ $Y2=0
cc_538 N_A_857_21#_c_769_p N_Q_c_1094_n 0.0181554f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_539 N_A_857_21#_c_655_n N_Q_c_1094_n 0.00268325f $X=7.565 $Y=1.525 $X2=0
+ $Y2=0
cc_540 N_A_857_21#_c_647_n N_Q_c_1095_n 8.9451e-19 $X=7.14 $Y=1.325 $X2=0 $Y2=0
cc_541 N_A_857_21#_c_648_n N_Q_c_1095_n 8.30973e-19 $X=7.57 $Y=1.325 $X2=0 $Y2=0
cc_542 N_A_857_21#_c_660_n N_Q_c_1100_n 0.0140138f $X=7.565 $Y=1.725 $X2=0 $Y2=0
cc_543 N_A_857_21#_c_655_n N_Q_c_1100_n 0.00162117f $X=7.565 $Y=1.525 $X2=0
+ $Y2=0
cc_544 N_A_857_21#_c_648_n Q 0.0118478f $X=7.57 $Y=1.325 $X2=0 $Y2=0
cc_545 N_A_857_21#_c_655_n Q 0.001296f $X=7.565 $Y=1.525 $X2=0 $Y2=0
cc_546 N_A_857_21#_c_659_n Q 5.44902e-19 $X=7.135 $Y=1.725 $X2=0 $Y2=0
cc_547 N_A_857_21#_c_647_n Q 0.0025678f $X=7.14 $Y=1.325 $X2=0 $Y2=0
cc_548 N_A_857_21#_c_660_n Q 7.78943e-19 $X=7.565 $Y=1.725 $X2=0 $Y2=0
cc_549 N_A_857_21#_c_648_n Q 0.0038143f $X=7.57 $Y=1.325 $X2=0 $Y2=0
cc_550 N_A_857_21#_c_769_p Q 0.0141537f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_551 N_A_857_21#_c_655_n Q 0.0372739f $X=7.565 $Y=1.525 $X2=0 $Y2=0
cc_552 N_A_857_21#_c_689_p N_VGND_M1021_d 0.00454173f $X=6.055 $Y=0.955 $X2=0
+ $Y2=0
cc_553 N_A_857_21#_c_651_n N_VGND_M1021_d 0.00186325f $X=6.142 $Y=1.405 $X2=0
+ $Y2=0
cc_554 N_A_857_21#_c_644_n N_VGND_c_1156_n 0.00322069f $X=4.36 $Y=0.765 $X2=0
+ $Y2=0
cc_555 N_A_857_21#_c_649_n N_VGND_c_1156_n 0.00234948f $X=4.44 $Y=0.84 $X2=0
+ $Y2=0
cc_556 N_A_857_21#_c_650_n N_VGND_c_1156_n 0.0107283f $X=5.125 $Y=0.525 $X2=0
+ $Y2=0
cc_557 N_A_857_21#_c_645_n N_VGND_c_1157_n 0.00818956f $X=6.28 $Y=1.325 $X2=0
+ $Y2=0
cc_558 N_A_857_21#_c_646_n N_VGND_c_1157_n 4.59734e-19 $X=6.71 $Y=1.325 $X2=0
+ $Y2=0
cc_559 N_A_857_21#_c_650_n N_VGND_c_1157_n 0.00410912f $X=5.125 $Y=0.525 $X2=0
+ $Y2=0
cc_560 N_A_857_21#_c_689_p N_VGND_c_1157_n 0.0180641f $X=6.055 $Y=0.955 $X2=0
+ $Y2=0
cc_561 N_A_857_21#_c_646_n N_VGND_c_1158_n 0.00251973f $X=6.71 $Y=1.325 $X2=0
+ $Y2=0
cc_562 N_A_857_21#_c_647_n N_VGND_c_1158_n 0.00245995f $X=7.14 $Y=1.325 $X2=0
+ $Y2=0
cc_563 N_A_857_21#_c_647_n N_VGND_c_1160_n 4.9918e-19 $X=7.14 $Y=1.325 $X2=0
+ $Y2=0
cc_564 N_A_857_21#_c_648_n N_VGND_c_1160_n 0.0113375f $X=7.57 $Y=1.325 $X2=0
+ $Y2=0
cc_565 N_A_857_21#_c_644_n N_VGND_c_1164_n 0.00445911f $X=4.36 $Y=0.765 $X2=0
+ $Y2=0
cc_566 N_A_857_21#_c_650_n N_VGND_c_1165_n 0.00891671f $X=5.125 $Y=0.525 $X2=0
+ $Y2=0
cc_567 N_A_857_21#_c_645_n N_VGND_c_1166_n 0.00386543f $X=6.28 $Y=1.325 $X2=0
+ $Y2=0
cc_568 N_A_857_21#_c_646_n N_VGND_c_1166_n 0.00465548f $X=6.71 $Y=1.325 $X2=0
+ $Y2=0
cc_569 N_A_857_21#_c_647_n N_VGND_c_1167_n 0.00465548f $X=7.14 $Y=1.325 $X2=0
+ $Y2=0
cc_570 N_A_857_21#_c_648_n N_VGND_c_1167_n 0.00386543f $X=7.57 $Y=1.325 $X2=0
+ $Y2=0
cc_571 N_A_857_21#_c_644_n N_VGND_c_1172_n 0.00662787f $X=4.36 $Y=0.765 $X2=0
+ $Y2=0
cc_572 N_A_857_21#_c_645_n N_VGND_c_1172_n 0.0076141f $X=6.28 $Y=1.325 $X2=0
+ $Y2=0
cc_573 N_A_857_21#_c_646_n N_VGND_c_1172_n 0.00914385f $X=6.71 $Y=1.325 $X2=0
+ $Y2=0
cc_574 N_A_857_21#_c_647_n N_VGND_c_1172_n 0.00914385f $X=7.14 $Y=1.325 $X2=0
+ $Y2=0
cc_575 N_A_857_21#_c_648_n N_VGND_c_1172_n 0.0076141f $X=7.57 $Y=1.325 $X2=0
+ $Y2=0
cc_576 N_A_857_21#_c_650_n N_VGND_c_1172_n 0.00680157f $X=5.125 $Y=0.525 $X2=0
+ $Y2=0
cc_577 N_A_857_21#_c_689_p A_1083_73# 0.0118207f $X=6.055 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_578 N_A_671_47#_c_824_n N_RESET_B_M1007_g 0.0369628f $X=5.265 $Y=1.65 $X2=0
+ $Y2=0
cc_579 N_A_671_47#_c_821_n RESET_B 5.64669e-19 $X=4.85 $Y=1.315 $X2=0 $Y2=0
cc_580 N_A_671_47#_c_824_n RESET_B 0.00903561f $X=5.265 $Y=1.65 $X2=0 $Y2=0
cc_581 N_A_671_47#_c_825_n RESET_B 0.00718309f $X=5.34 $Y=0.255 $X2=0 $Y2=0
cc_582 N_A_671_47#_c_834_n RESET_B 0.0194591f $X=5.34 $Y=1.725 $X2=0 $Y2=0
cc_583 N_A_671_47#_c_829_n RESET_B 0.0204784f $X=4.89 $Y=1.48 $X2=0 $Y2=0
cc_584 N_A_671_47#_c_830_n RESET_B 0.00118304f $X=4.89 $Y=1.48 $X2=0 $Y2=0
cc_585 N_A_671_47#_c_824_n N_RESET_B_c_938_n 0.00455934f $X=5.265 $Y=1.65 $X2=0
+ $Y2=0
cc_586 N_A_671_47#_c_825_n N_RESET_B_c_938_n 0.00129249f $X=5.34 $Y=0.255 $X2=0
+ $Y2=0
cc_587 N_A_671_47#_c_829_n N_RESET_B_c_938_n 2.38485e-19 $X=4.89 $Y=1.48 $X2=0
+ $Y2=0
cc_588 N_A_671_47#_c_830_n N_RESET_B_c_938_n 0.00363765f $X=4.89 $Y=1.48 $X2=0
+ $Y2=0
cc_589 N_A_671_47#_c_822_n N_RESET_B_c_939_n 0.0359806f $X=5.265 $Y=0.18 $X2=0
+ $Y2=0
cc_590 N_A_671_47#_c_834_n N_VPWR_c_988_n 0.0129067f $X=5.34 $Y=1.725 $X2=0
+ $Y2=0
cc_591 N_A_671_47#_c_834_n N_VPWR_c_996_n 0.00486043f $X=5.34 $Y=1.725 $X2=0
+ $Y2=0
cc_592 N_A_671_47#_c_834_n N_VPWR_c_985_n 0.0082726f $X=5.34 $Y=1.725 $X2=0
+ $Y2=0
cc_593 N_A_671_47#_c_837_n N_VGND_c_1155_n 0.00695402f $X=4.085 $Y=0.375 $X2=0
+ $Y2=0
cc_594 N_A_671_47#_c_823_n N_VGND_c_1156_n 0.00864157f $X=4.925 $Y=0.18 $X2=0
+ $Y2=0
cc_595 N_A_671_47#_c_822_n N_VGND_c_1157_n 0.00399361f $X=5.265 $Y=0.18 $X2=0
+ $Y2=0
cc_596 N_A_671_47#_c_837_n N_VGND_c_1164_n 0.0460912f $X=4.085 $Y=0.375 $X2=0
+ $Y2=0
cc_597 N_A_671_47#_c_831_n N_VGND_c_1164_n 0.00218966f $X=4.34 $Y=0.81 $X2=0
+ $Y2=0
cc_598 N_A_671_47#_c_823_n N_VGND_c_1165_n 0.0214712f $X=4.925 $Y=0.18 $X2=0
+ $Y2=0
cc_599 N_A_671_47#_M1009_d N_VGND_c_1172_n 0.00347107f $X=3.355 $Y=0.235 $X2=0
+ $Y2=0
cc_600 N_A_671_47#_c_822_n N_VGND_c_1172_n 0.0245037f $X=5.265 $Y=0.18 $X2=0
+ $Y2=0
cc_601 N_A_671_47#_c_823_n N_VGND_c_1172_n 0.010142f $X=4.925 $Y=0.18 $X2=0
+ $Y2=0
cc_602 N_A_671_47#_c_837_n N_VGND_c_1172_n 0.0303761f $X=4.085 $Y=0.375 $X2=0
+ $Y2=0
cc_603 N_A_671_47#_c_831_n N_VGND_c_1172_n 0.00357682f $X=4.34 $Y=0.81 $X2=0
+ $Y2=0
cc_604 N_A_671_47#_c_837_n A_779_47# 0.00691306f $X=4.085 $Y=0.375 $X2=-0.19
+ $Y2=-0.245
cc_605 N_A_671_47#_c_827_n A_779_47# 0.00258734f $X=4.175 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_606 N_RESET_B_M1007_g N_VPWR_c_988_n 5.88023e-19 $X=5.77 $Y=2.465 $X2=0 $Y2=0
cc_607 N_RESET_B_M1007_g N_VPWR_c_989_n 0.00257861f $X=5.77 $Y=2.465 $X2=0 $Y2=0
cc_608 N_RESET_B_M1007_g N_VPWR_c_996_n 0.00585385f $X=5.77 $Y=2.465 $X2=0 $Y2=0
cc_609 N_RESET_B_M1007_g N_VPWR_c_985_n 0.0108521f $X=5.77 $Y=2.465 $X2=0 $Y2=0
cc_610 N_RESET_B_c_939_n N_VGND_c_1157_n 0.0118504f $X=5.79 $Y=1.315 $X2=0 $Y2=0
cc_611 N_RESET_B_c_939_n N_VGND_c_1165_n 0.00386543f $X=5.79 $Y=1.315 $X2=0
+ $Y2=0
cc_612 N_RESET_B_c_939_n N_VGND_c_1172_n 0.00762996f $X=5.79 $Y=1.315 $X2=0
+ $Y2=0
cc_613 N_VPWR_c_985_n N_Q_M1008_d 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_614 N_VPWR_c_985_n N_Q_M1018_d 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_615 N_VPWR_c_997_n N_Q_c_1134_n 0.0124525f $X=6.755 $Y=3.33 $X2=0 $Y2=0
cc_616 N_VPWR_c_985_n N_Q_c_1134_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_617 N_VPWR_M1015_s N_Q_c_1098_n 0.00176461f $X=6.78 $Y=1.835 $X2=0 $Y2=0
cc_618 N_VPWR_c_990_n N_Q_c_1098_n 0.0170777f $X=6.92 $Y=2.17 $X2=0 $Y2=0
cc_619 N_VPWR_c_998_n N_Q_c_1138_n 0.0124525f $X=7.615 $Y=3.33 $X2=0 $Y2=0
cc_620 N_VPWR_c_985_n N_Q_c_1138_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_621 N_VPWR_M1023_s N_Q_c_1100_n 0.00267816f $X=7.64 $Y=1.835 $X2=0 $Y2=0
cc_622 N_VPWR_c_992_n N_Q_c_1100_n 0.0243971f $X=7.78 $Y=2.17 $X2=0 $Y2=0
cc_623 N_Q_c_1093_n N_VGND_M1005_s 0.00176461f $X=7.225 $Y=1.15 $X2=0 $Y2=0
cc_624 Q N_VGND_M1019_s 0.00277226f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_625 N_Q_c_1092_n N_VGND_c_1157_n 0.0132986f $X=6.495 $Y=0.52 $X2=0 $Y2=0
cc_626 N_Q_c_1092_n N_VGND_c_1158_n 7.14495e-19 $X=6.495 $Y=0.52 $X2=0 $Y2=0
cc_627 N_Q_c_1093_n N_VGND_c_1158_n 0.0135055f $X=7.225 $Y=1.15 $X2=0 $Y2=0
cc_628 N_Q_c_1095_n N_VGND_c_1158_n 0.00150838f $X=7.355 $Y=0.51 $X2=0 $Y2=0
cc_629 N_Q_c_1095_n N_VGND_c_1160_n 0.0228841f $X=7.355 $Y=0.51 $X2=0 $Y2=0
cc_630 Q N_VGND_c_1160_n 0.0243971f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_631 N_Q_c_1092_n N_VGND_c_1166_n 0.00975472f $X=6.495 $Y=0.52 $X2=0 $Y2=0
cc_632 N_Q_c_1095_n N_VGND_c_1167_n 0.010154f $X=7.355 $Y=0.51 $X2=0 $Y2=0
cc_633 N_Q_c_1092_n N_VGND_c_1172_n 0.00821134f $X=6.495 $Y=0.52 $X2=0 $Y2=0
cc_634 N_Q_c_1095_n N_VGND_c_1172_n 0.00826079f $X=7.355 $Y=0.51 $X2=0 $Y2=0
cc_635 N_VGND_c_1172_n A_599_47# 0.00250288f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
cc_636 N_VGND_c_1172_n A_779_47# 0.00324826f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
