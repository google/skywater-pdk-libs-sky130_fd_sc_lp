* NGSPICE file created from sky130_fd_sc_lp__or2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or2b_2 A B_N VGND VNB VPB VPWR X
M1000 X a_191_254# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=9.857e+11p ps=7.64e+06u
M1001 VGND B_N a_27_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1002 VPWR a_191_254# X VPB phighvt w=1.26e+06u l=150000u
+  ad=8.862e+11p pd=7.14e+06u as=3.528e+11p ps=3.08e+06u
M1003 VGND a_191_254# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_191_254# A VGND VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1005 VPWR B_N a_27_49# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1006 a_479_367# A VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 a_191_254# a_27_49# a_479_367# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 X a_191_254# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_49# a_191_254# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

