* NGSPICE file created from sky130_fd_sc_lp__dlxbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_214_136# a_354_47# VPB phighvt w=640000u l=150000u
+  ad=2.3303e+12p pd=1.783e+07u as=1.696e+11p ps=1.81e+06u
M1001 a_547_47# a_45_136# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.7475e+12p ps=1.394e+07u
M1002 a_737_47# a_354_47# a_619_47# VNB nshort w=420000u l=150000u
+  ad=1.428e+11p pd=1.52e+06u as=1.877e+11p ps=1.74e+06u
M1003 VPWR a_1138_153# Q_N VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1004 Q a_805_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1005 VPWR a_805_21# a_769_491# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_769_491# a_214_136# a_619_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.221e+11p ps=2.06e+06u
M1007 VGND a_1138_153# Q_N VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1008 Q a_805_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1009 VPWR a_805_21# a_1138_153# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1010 VGND a_214_136# a_354_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 VPWR D a_45_136# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.048e+11p ps=1.92e+06u
M1012 a_805_21# a_619_47# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1013 a_214_136# GATE_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1014 VGND D a_45_136# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1015 Q_N a_1138_153# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_805_21# a_619_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1017 VGND a_805_21# a_737_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_805_21# a_1138_153# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1019 a_214_136# GATE_N VPWR VPB phighvt w=640000u l=150000u
+  ad=3.459e+11p pd=2.7e+06u as=0p ps=0u
M1020 a_619_47# a_354_47# a_589_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1021 VPWR a_805_21# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_619_47# a_214_136# a_547_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_589_491# a_45_136# VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Q_N a_1138_153# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_805_21# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

