# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__clkinvlp_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__clkinvlp_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  5.650000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.075000 1.180000 8.545000 1.410000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.010000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.575000 1.920000 8.355000 2.150000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 9.120000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 9.310000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.095000  0.085000 0.425000 0.775000 ;
      RECT 0.095000  1.960000 0.425000 3.245000 ;
      RECT 0.100000  1.105000 0.455000 1.780000 ;
      RECT 0.625000  0.315000 1.215000 0.780000 ;
      RECT 0.625000  0.780000 0.955000 1.010000 ;
      RECT 0.625000  1.010000 0.905000 1.735000 ;
      RECT 0.625000  1.735000 0.955000 3.000000 ;
      RECT 1.075000  1.180000 2.265000 1.565000 ;
      RECT 1.155000  1.960000 1.485000 3.245000 ;
      RECT 1.675000  0.085000 2.005000 0.775000 ;
      RECT 1.685000  1.920000 2.015000 3.000000 ;
      RECT 2.215000  1.960000 2.545000 3.245000 ;
      RECT 2.465000  0.445000 2.795000 1.195000 ;
      RECT 2.465000  1.195000 3.075000 1.565000 ;
      RECT 2.745000  1.565000 3.075000 3.000000 ;
      RECT 3.255000  0.085000 3.585000 0.775000 ;
      RECT 3.275000  1.180000 3.710000 1.565000 ;
      RECT 3.275000  1.960000 3.605000 3.245000 ;
      RECT 3.805000  1.805000 4.135000 3.000000 ;
      RECT 3.880000  1.195000 4.375000 1.565000 ;
      RECT 3.880000  1.565000 4.135000 1.805000 ;
      RECT 4.045000  0.445000 4.375000 1.195000 ;
      RECT 4.335000  1.960000 4.665000 3.245000 ;
      RECT 4.655000  1.180000 5.380000 1.565000 ;
      RECT 4.835000  0.085000 5.165000 0.775000 ;
      RECT 4.865000  1.920000 5.195000 3.000000 ;
      RECT 5.395000  1.960000 5.725000 3.245000 ;
      RECT 5.625000  0.445000 5.955000 1.195000 ;
      RECT 5.625000  1.195000 6.190000 1.565000 ;
      RECT 5.895000  1.565000 6.190000 1.875000 ;
      RECT 5.895000  1.875000 6.255000 3.000000 ;
      RECT 6.370000  1.180000 6.700000 1.565000 ;
      RECT 6.415000  0.085000 6.745000 0.775000 ;
      RECT 6.455000  1.960000 6.785000 3.245000 ;
      RECT 6.985000  1.195000 7.535000 1.565000 ;
      RECT 6.985000  1.565000 7.315000 3.000000 ;
      RECT 7.205000  0.445000 7.535000 1.195000 ;
      RECT 7.515000  1.960000 7.845000 3.245000 ;
      RECT 7.705000  1.180000 8.715000 1.565000 ;
      RECT 7.995000  0.085000 8.325000 0.775000 ;
      RECT 8.045000  1.920000 8.375000 3.000000 ;
      RECT 8.575000  1.960000 8.905000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  1.210000 0.325000 1.380000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  1.950000 0.805000 2.120000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  1.210000 1.285000 1.380000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  1.210000 1.765000 1.380000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 1.765000  1.950000 1.935000 2.120000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  1.210000 2.245000 1.380000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 2.825000  1.950000 2.995000 2.120000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  1.210000 3.685000 1.380000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.885000  1.950000 4.055000 2.120000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  1.210000 5.125000 1.380000 ;
      RECT 4.955000  1.950000 5.125000 2.120000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  1.950000 6.085000 2.120000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  1.210000 6.565000 1.380000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.065000  1.950000 7.235000 2.120000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  1.210000 8.005000 1.380000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.125000  1.950000 8.295000 2.120000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  1.210000 8.485000 1.380000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_lp__clkinvlp_16
END LIBRARY
