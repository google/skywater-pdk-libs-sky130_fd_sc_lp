* File: sky130_fd_sc_lp__o21ai_4.pxi.spice
* Created: Wed Sep  2 10:16:13 2020
* 
x_PM_SKY130_FD_SC_LP__O21AI_4%A1 N_A1_c_87_n N_A1_M1011_g N_A1_M1006_g
+ N_A1_c_89_n N_A1_M1015_g N_A1_M1012_g N_A1_c_91_n N_A1_M1019_g N_A1_M1013_g
+ N_A1_M1020_g N_A1_M1022_g N_A1_c_94_n N_A1_c_95_n N_A1_c_96_n A1 A1 A1 A1
+ N_A1_c_97_n N_A1_c_98_n N_A1_c_99_n N_A1_c_100_n
+ PM_SKY130_FD_SC_LP__O21AI_4%A1
x_PM_SKY130_FD_SC_LP__O21AI_4%A2 N_A2_M1004_g N_A2_M1001_g N_A2_M1008_g
+ N_A2_M1005_g N_A2_M1016_g N_A2_M1010_g N_A2_M1018_g N_A2_M1021_g A2 A2 A2
+ N_A2_c_203_n PM_SKY130_FD_SC_LP__O21AI_4%A2
x_PM_SKY130_FD_SC_LP__O21AI_4%B1 N_B1_c_284_n N_B1_M1000_g N_B1_M1002_g
+ N_B1_c_286_n N_B1_M1003_g N_B1_M1007_g N_B1_c_288_n N_B1_M1009_g N_B1_M1017_g
+ N_B1_c_290_n N_B1_M1014_g N_B1_M1023_g B1 B1 B1 N_B1_c_293_n
+ PM_SKY130_FD_SC_LP__O21AI_4%B1
x_PM_SKY130_FD_SC_LP__O21AI_4%VPWR N_VPWR_M1006_d N_VPWR_M1012_d N_VPWR_M1020_d
+ N_VPWR_M1007_s N_VPWR_M1023_s N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n
+ N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n VPWR
+ N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n
+ N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_353_n PM_SKY130_FD_SC_LP__O21AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O21AI_4%A_115_367# N_A_115_367#_M1006_s
+ N_A_115_367#_M1013_s N_A_115_367#_M1005_d N_A_115_367#_M1021_d
+ N_A_115_367#_c_460_n N_A_115_367#_c_441_n N_A_115_367#_c_442_n
+ N_A_115_367#_c_465_n N_A_115_367#_c_452_n N_A_115_367#_c_476_p
+ N_A_115_367#_c_454_n N_A_115_367#_c_478_p N_A_115_367#_c_471_n
+ PM_SKY130_FD_SC_LP__O21AI_4%A_115_367#
x_PM_SKY130_FD_SC_LP__O21AI_4%Y N_Y_M1000_d N_Y_M1009_d N_Y_M1001_s N_Y_M1010_s
+ N_Y_M1002_d N_Y_M1017_d N_Y_c_494_n N_Y_c_488_n N_Y_c_532_n N_Y_c_481_n
+ N_Y_c_482_n N_Y_c_483_n N_Y_c_538_n N_Y_c_502_n N_Y_c_493_n N_Y_c_484_n Y
+ PM_SKY130_FD_SC_LP__O21AI_4%Y
x_PM_SKY130_FD_SC_LP__O21AI_4%A_32_47# N_A_32_47#_M1011_s N_A_32_47#_M1015_s
+ N_A_32_47#_M1004_s N_A_32_47#_M1016_s N_A_32_47#_M1022_s N_A_32_47#_M1003_s
+ N_A_32_47#_M1014_s N_A_32_47#_c_560_n N_A_32_47#_c_564_n N_A_32_47#_c_561_n
+ N_A_32_47#_c_610_p N_A_32_47#_c_570_n N_A_32_47#_c_613_p N_A_32_47#_c_573_n
+ N_A_32_47#_c_616_p N_A_32_47#_c_574_n N_A_32_47#_c_588_n N_A_32_47#_c_578_n
+ N_A_32_47#_c_562_n N_A_32_47#_c_580_n N_A_32_47#_c_582_n N_A_32_47#_c_583_n
+ PM_SKY130_FD_SC_LP__O21AI_4%A_32_47#
x_PM_SKY130_FD_SC_LP__O21AI_4%VGND N_VGND_M1011_d N_VGND_M1019_d N_VGND_M1008_d
+ N_VGND_M1018_d N_VGND_c_639_n N_VGND_c_640_n N_VGND_c_641_n N_VGND_c_642_n
+ N_VGND_c_643_n N_VGND_c_644_n N_VGND_c_645_n N_VGND_c_646_n N_VGND_c_647_n
+ N_VGND_c_648_n VGND N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n
+ N_VGND_c_652_n PM_SKY130_FD_SC_LP__O21AI_4%VGND
cc_1 VNB N_A1_c_87_n 0.0218823f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_2 VNB N_A1_M1006_g 0.0111859f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_3 VNB N_A1_c_89_n 0.0159814f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.185
cc_4 VNB N_A1_M1012_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.465
cc_5 VNB N_A1_c_91_n 0.0155545f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_6 VNB N_A1_M1013_g 0.00730151f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.465
cc_7 VNB N_A1_M1020_g 0.00769966f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=2.465
cc_8 VNB N_A1_c_94_n 0.0240154f $X=-0.19 $Y=-0.245 $X2=3.445 $Y2=1.16
cc_9 VNB N_A1_c_95_n 0.00251498f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=1.16
cc_10 VNB N_A1_c_96_n 0.0323821f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=1.35
cc_11 VNB N_A1_c_97_n 0.0887232f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.35
cc_12 VNB N_A1_c_98_n 0.0157708f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=1.185
cc_13 VNB N_A1_c_99_n 0.0123404f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.295
cc_14 VNB N_A1_c_100_n 0.00641466f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=1.295
cc_15 VNB N_A2_M1004_g 0.0220385f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_16 VNB N_A2_M1008_g 0.022674f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.515
cc_17 VNB N_A2_M1016_g 0.0227036f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.465
cc_18 VNB N_A2_M1018_g 0.0227913f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=0.655
cc_19 VNB A2 0.00316813f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=1.35
cc_20 VNB N_A2_c_203_n 0.0632941f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.35
cc_21 VNB N_B1_c_284_n 0.0164f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_22 VNB N_B1_M1002_g 0.00701446f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_23 VNB N_B1_c_286_n 0.0162039f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.185
cc_24 VNB N_B1_M1007_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=2.465
cc_25 VNB N_B1_c_288_n 0.0162015f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_26 VNB N_B1_M1017_g 0.00663861f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.465
cc_27 VNB N_B1_c_290_n 0.0192832f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.515
cc_28 VNB N_B1_M1023_g 0.00774528f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=0.655
cc_29 VNB B1 0.00149192f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=1.16
cc_30 VNB N_B1_c_293_n 0.0769828f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.35
cc_31 VNB N_VPWR_c_353_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_481_n 0.0148033f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=1.16
cc_33 VNB N_Y_c_482_n 0.00307882f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_Y_c_483_n 0.003947f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_35 VNB N_Y_c_484_n 0.00589876f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.35
cc_36 VNB Y 0.0292025f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=1.185
cc_37 VNB N_A_32_47#_c_560_n 0.0233935f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=2.465
cc_38 VNB N_A_32_47#_c_561_n 0.00757813f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=0.655
cc_39 VNB N_A_32_47#_c_562_n 0.0121795f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.35
cc_40 VNB N_VGND_c_639_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.185
cc_41 VNB N_VGND_c_640_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.465
cc_42 VNB N_VGND_c_641_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=2.465
cc_43 VNB N_VGND_c_642_n 0.00274151f $X=-0.19 $Y=-0.245 $X2=3.55 $Y2=0.655
cc_44 VNB N_VGND_c_643_n 0.0123027f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=1.16
cc_45 VNB N_VGND_c_644_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=1.16
cc_46 VNB N_VGND_c_645_n 0.011684f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=1.35
cc_47 VNB N_VGND_c_646_n 0.00436716f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=1.35
cc_48 VNB N_VGND_c_647_n 0.011684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_648_n 0.0051069f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_50 VNB N_VGND_c_649_n 0.0161714f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_51 VNB N_VGND_c_650_n 0.0551225f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=1.362
cc_52 VNB N_VGND_c_651_n 0.289354f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.362
cc_53 VNB N_VGND_c_652_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.362
cc_54 VPB N_A1_M1006_g 0.0269287f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_55 VPB N_A1_M1012_g 0.018914f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.465
cc_56 VPB N_A1_M1013_g 0.0191417f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.465
cc_57 VPB N_A1_M1020_g 0.0202192f $X=-0.19 $Y=1.655 $X2=3.51 $Y2=2.465
cc_58 VPB N_A2_M1001_g 0.0190209f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A2_M1005_g 0.0180507f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=1.185
cc_60 VPB N_A2_M1010_g 0.0180542f $X=-0.19 $Y=1.655 $X2=3.51 $Y2=2.465
cc_61 VPB N_A2_M1021_g 0.0182305f $X=-0.19 $Y=1.655 $X2=3.57 $Y2=1.16
cc_62 VPB A2 0.0095727f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=1.35
cc_63 VPB N_A2_c_203_n 0.0121773f $X=-0.19 $Y=1.655 $X2=1.31 $Y2=1.35
cc_64 VPB N_B1_M1002_g 0.0185106f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_65 VPB N_B1_M1007_g 0.0180695f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=2.465
cc_66 VPB N_B1_M1017_g 0.0180695f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.465
cc_67 VPB N_B1_M1023_g 0.0227978f $X=-0.19 $Y=1.655 $X2=3.55 $Y2=0.655
cc_68 VPB N_VPWR_c_354_n 0.0114848f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=0.655
cc_69 VPB N_VPWR_c_355_n 0.055719f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=1.515
cc_70 VPB N_VPWR_c_356_n 4.06898e-19 $X=-0.19 $Y=1.655 $X2=3.51 $Y2=2.465
cc_71 VPB N_VPWR_c_357_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=1.825 $Y2=1.16
cc_72 VPB N_VPWR_c_358_n 3.12649e-19 $X=-0.19 $Y=1.655 $X2=3.53 $Y2=1.35
cc_73 VPB N_VPWR_c_359_n 0.0108182f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_74 VPB N_VPWR_c_360_n 0.0412093f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_75 VPB N_VPWR_c_361_n 0.0149824f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.35
cc_76 VPB N_VPWR_c_362_n 0.0514145f $X=-0.19 $Y=1.655 $X2=1.31 $Y2=1.35
cc_77 VPB N_VPWR_c_363_n 0.0133881f $X=-0.19 $Y=1.655 $X2=3.53 $Y2=1.35
cc_78 VPB N_VPWR_c_364_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_365_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_366_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_367_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_353_n 0.0454562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A_115_367#_c_441_n 0.00626995f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.465
cc_84 VPB N_A_115_367#_c_442_n 0.00244447f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.465
cc_85 VPB N_Y_c_483_n 0.00821092f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_86 VPB N_Y_c_484_n 0.0132668f $X=-0.19 $Y=1.655 $X2=1.31 $Y2=1.35
cc_87 N_A1_c_91_n N_A2_M1004_g 0.0310833f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_88 N_A1_c_94_n N_A2_M1004_g 0.00488235f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A1_c_97_n N_A2_M1004_g 0.0182178f $X=1.36 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A1_c_100_n N_A2_M1004_g 0.00879766f $X=1.825 $Y=1.295 $X2=0 $Y2=0
cc_91 N_A1_c_94_n N_A2_M1008_g 0.0105539f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A1_c_100_n N_A2_M1008_g 5.64968e-19 $X=1.825 $Y=1.295 $X2=0 $Y2=0
cc_93 N_A1_c_94_n N_A2_M1016_g 0.0105539f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A1_c_94_n N_A2_M1018_g 0.0102909f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A1_c_95_n N_A2_M1018_g 0.00118562f $X=3.57 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A1_c_96_n N_A2_M1018_g 0.0217495f $X=3.53 $Y=1.35 $X2=0 $Y2=0
cc_97 N_A1_c_98_n N_A2_M1018_g 0.0274869f $X=3.53 $Y=1.185 $X2=0 $Y2=0
cc_98 N_A1_M1013_g A2 5.87554e-19 $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A1_M1020_g A2 0.00450157f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A1_c_94_n A2 0.0910584f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A1_c_95_n A2 0.00736506f $X=3.57 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A1_c_96_n A2 6.4198e-19 $X=3.53 $Y=1.35 $X2=0 $Y2=0
cc_103 N_A1_c_100_n A2 0.00744928f $X=1.825 $Y=1.295 $X2=0 $Y2=0
cc_104 N_A1_M1013_g N_A2_c_203_n 0.0272915f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A1_M1020_g N_A2_c_203_n 0.0410659f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A1_c_94_n N_A2_c_203_n 0.00798889f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A1_c_100_n N_A2_c_203_n 0.0144204f $X=1.825 $Y=1.295 $X2=0 $Y2=0
cc_108 N_A1_c_95_n N_B1_c_284_n 0.0023336f $X=3.57 $Y=1.16 $X2=-0.19 $Y2=-0.245
cc_109 N_A1_c_98_n N_B1_c_284_n 0.0143828f $X=3.53 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_110 N_A1_M1020_g N_B1_M1002_g 0.0371529f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A1_c_95_n B1 0.014723f $X=3.57 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A1_c_96_n B1 7.75083e-19 $X=3.53 $Y=1.35 $X2=0 $Y2=0
cc_113 N_A1_c_95_n N_B1_c_293_n 0.00110601f $X=3.57 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A1_c_96_n N_B1_c_293_n 0.0217296f $X=3.53 $Y=1.35 $X2=0 $Y2=0
cc_115 N_A1_M1006_g N_VPWR_c_355_n 0.00757423f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A1_c_97_n N_VPWR_c_355_n 0.00603039f $X=1.36 $Y=1.35 $X2=0 $Y2=0
cc_117 N_A1_c_99_n N_VPWR_c_355_n 0.0153409f $X=1.42 $Y=1.295 $X2=0 $Y2=0
cc_118 N_A1_M1006_g N_VPWR_c_356_n 7.45395e-19 $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A1_M1012_g N_VPWR_c_356_n 0.0143822f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A1_M1013_g N_VPWR_c_356_n 0.015452f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A1_M1020_g N_VPWR_c_357_n 0.013743f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A1_M1006_g N_VPWR_c_361_n 0.00585385f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A1_M1012_g N_VPWR_c_361_n 0.00486043f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A1_M1013_g N_VPWR_c_362_n 0.00486043f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A1_M1020_g N_VPWR_c_362_n 0.00564095f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A1_M1006_g N_VPWR_c_353_n 0.0115052f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A1_M1012_g N_VPWR_c_353_n 0.00824727f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A1_M1013_g N_VPWR_c_353_n 0.0082726f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A1_M1020_g N_VPWR_c_353_n 0.00950825f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A1_M1012_g N_A_115_367#_c_441_n 0.0135574f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A1_M1013_g N_A_115_367#_c_441_n 0.0133703f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A1_c_97_n N_A_115_367#_c_441_n 0.00299406f $X=1.36 $Y=1.35 $X2=0 $Y2=0
cc_133 N_A1_c_99_n N_A_115_367#_c_441_n 0.037557f $X=1.42 $Y=1.295 $X2=0 $Y2=0
cc_134 N_A1_c_100_n N_A_115_367#_c_441_n 0.0134746f $X=1.825 $Y=1.295 $X2=0
+ $Y2=0
cc_135 N_A1_M1006_g N_A_115_367#_c_442_n 0.00221438f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A1_c_97_n N_A_115_367#_c_442_n 0.00224327f $X=1.36 $Y=1.35 $X2=0 $Y2=0
cc_137 N_A1_c_99_n N_A_115_367#_c_442_n 0.015242f $X=1.42 $Y=1.295 $X2=0 $Y2=0
cc_138 N_A1_M1020_g N_Y_c_488_n 0.00289854f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A1_c_96_n N_Y_c_488_n 0.00126677f $X=3.53 $Y=1.35 $X2=0 $Y2=0
cc_140 N_A1_M1020_g N_Y_c_483_n 0.0220793f $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A1_c_95_n N_Y_c_483_n 0.0150675f $X=3.57 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A1_c_96_n N_Y_c_483_n 7.62844e-19 $X=3.53 $Y=1.35 $X2=0 $Y2=0
cc_143 N_A1_M1020_g N_Y_c_493_n 8.92984e-19 $X=3.51 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A1_c_95_n N_A_32_47#_M1022_s 7.53634e-19 $X=3.57 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A1_c_87_n N_A_32_47#_c_564_n 0.0122129f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_146 N_A1_c_89_n N_A_32_47#_c_564_n 0.0126062f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_147 N_A1_c_97_n N_A_32_47#_c_564_n 0.00230884f $X=1.36 $Y=1.35 $X2=0 $Y2=0
cc_148 N_A1_c_99_n N_A_32_47#_c_564_n 0.0410001f $X=1.42 $Y=1.295 $X2=0 $Y2=0
cc_149 N_A1_c_97_n N_A_32_47#_c_561_n 0.00608363f $X=1.36 $Y=1.35 $X2=0 $Y2=0
cc_150 N_A1_c_99_n N_A_32_47#_c_561_n 0.0204654f $X=1.42 $Y=1.295 $X2=0 $Y2=0
cc_151 N_A1_c_91_n N_A_32_47#_c_570_n 0.0105376f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_152 N_A1_c_99_n N_A_32_47#_c_570_n 0.00677081f $X=1.42 $Y=1.295 $X2=0 $Y2=0
cc_153 N_A1_c_100_n N_A_32_47#_c_570_n 0.0316798f $X=1.825 $Y=1.295 $X2=0 $Y2=0
cc_154 N_A1_c_94_n N_A_32_47#_c_573_n 0.0402256f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A1_c_94_n N_A_32_47#_c_574_n 0.0302273f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A1_c_95_n N_A_32_47#_c_574_n 0.0124178f $X=3.57 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A1_c_96_n N_A_32_47#_c_574_n 3.779e-19 $X=3.53 $Y=1.35 $X2=0 $Y2=0
cc_158 N_A1_c_98_n N_A_32_47#_c_574_n 0.0103867f $X=3.53 $Y=1.185 $X2=0 $Y2=0
cc_159 N_A1_c_95_n N_A_32_47#_c_578_n 0.00324214f $X=3.57 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A1_c_96_n N_A_32_47#_c_578_n 2.56976e-19 $X=3.53 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A1_c_97_n N_A_32_47#_c_580_n 0.00240082f $X=1.36 $Y=1.35 $X2=0 $Y2=0
cc_162 N_A1_c_99_n N_A_32_47#_c_580_n 0.0148254f $X=1.42 $Y=1.295 $X2=0 $Y2=0
cc_163 N_A1_c_94_n N_A_32_47#_c_582_n 0.0145842f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A1_c_94_n N_A_32_47#_c_583_n 0.0145842f $X=3.445 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A1_c_95_n N_VGND_M1018_d 3.17466e-19 $X=3.57 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A1_c_87_n N_VGND_c_639_n 0.0120167f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_167 N_A1_c_89_n N_VGND_c_639_n 0.0103296f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_168 N_A1_c_91_n N_VGND_c_639_n 5.75816e-19 $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A1_c_89_n N_VGND_c_640_n 5.37623e-19 $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_170 N_A1_c_91_n N_VGND_c_640_n 0.00754158f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_171 N_A1_c_98_n N_VGND_c_642_n 0.00325355f $X=3.53 $Y=1.185 $X2=0 $Y2=0
cc_172 N_A1_c_89_n N_VGND_c_643_n 0.00486043f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_173 N_A1_c_91_n N_VGND_c_643_n 0.00365202f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_174 N_A1_c_87_n N_VGND_c_649_n 0.00486043f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_175 N_A1_c_98_n N_VGND_c_650_n 0.00439206f $X=3.53 $Y=1.185 $X2=0 $Y2=0
cc_176 N_A1_c_87_n N_VGND_c_651_n 0.00920269f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_177 N_A1_c_89_n N_VGND_c_651_n 0.00824727f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_178 N_A1_c_91_n N_VGND_c_651_n 0.00432244f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_179 N_A1_c_98_n N_VGND_c_651_n 0.0061038f $X=3.53 $Y=1.185 $X2=0 $Y2=0
cc_180 N_A2_M1001_g N_VPWR_c_356_n 0.00109252f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A2_M1021_g N_VPWR_c_357_n 0.00105138f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A2_M1001_g N_VPWR_c_362_n 0.00357877f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A2_M1005_g N_VPWR_c_362_n 0.00357877f $X=2.22 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A2_M1010_g N_VPWR_c_362_n 0.00357877f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A2_M1021_g N_VPWR_c_362_n 0.00357877f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A2_M1001_g N_VPWR_c_353_n 0.00537654f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A2_M1005_g N_VPWR_c_353_n 0.0053512f $X=2.22 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A2_M1010_g N_VPWR_c_353_n 0.0053512f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A2_M1021_g N_VPWR_c_353_n 0.00537654f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A2_M1001_g N_A_115_367#_c_441_n 0.00253514f $X=1.79 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A2_M1001_g N_A_115_367#_c_452_n 0.0115031f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A2_M1005_g N_A_115_367#_c_452_n 0.0114565f $X=2.22 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A2_M1010_g N_A_115_367#_c_454_n 0.0114565f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A2_M1021_g N_A_115_367#_c_454_n 0.0115031f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A2_M1005_g N_Y_c_494_n 0.01115f $X=2.22 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A2_M1010_g N_Y_c_494_n 0.01115f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_197 A2 N_Y_c_494_n 0.0355198f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_198 N_A2_c_203_n N_Y_c_494_n 5.64665e-19 $X=3.08 $Y=1.51 $X2=0 $Y2=0
cc_199 N_A2_M1021_g N_Y_c_488_n 0.0111034f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_200 A2 N_Y_c_488_n 0.016199f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_201 N_A2_M1021_g N_Y_c_483_n 0.00103938f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_202 A2 N_Y_c_483_n 0.00582801f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A2_M1001_g N_Y_c_502_n 0.0112111f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A2_M1005_g N_Y_c_502_n 0.0102126f $X=2.22 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A2_M1010_g N_Y_c_502_n 5.66402e-19 $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_206 A2 N_Y_c_502_n 0.0124153f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_207 N_A2_c_203_n N_Y_c_502_n 0.00200545f $X=3.08 $Y=1.51 $X2=0 $Y2=0
cc_208 N_A2_M1005_g N_Y_c_493_n 5.66402e-19 $X=2.22 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A2_M1010_g N_Y_c_493_n 0.0102126f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A2_M1021_g N_Y_c_493_n 0.0103514f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_211 A2 N_Y_c_493_n 0.0230948f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_212 N_A2_c_203_n N_Y_c_493_n 6.37898e-19 $X=3.08 $Y=1.51 $X2=0 $Y2=0
cc_213 N_A2_M1004_g N_A_32_47#_c_570_n 0.0098539f $X=1.79 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A2_M1008_g N_A_32_47#_c_573_n 0.00990046f $X=2.22 $Y=0.655 $X2=0 $Y2=0
cc_215 N_A2_M1016_g N_A_32_47#_c_573_n 0.00990046f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_216 N_A2_M1018_g N_A_32_47#_c_574_n 0.010079f $X=3.08 $Y=0.655 $X2=0 $Y2=0
cc_217 N_A2_M1004_g N_VGND_c_640_n 0.00754158f $X=1.79 $Y=0.655 $X2=0 $Y2=0
cc_218 N_A2_M1008_g N_VGND_c_640_n 5.37623e-19 $X=2.22 $Y=0.655 $X2=0 $Y2=0
cc_219 N_A2_M1004_g N_VGND_c_641_n 5.37623e-19 $X=1.79 $Y=0.655 $X2=0 $Y2=0
cc_220 N_A2_M1008_g N_VGND_c_641_n 0.00758038f $X=2.22 $Y=0.655 $X2=0 $Y2=0
cc_221 N_A2_M1016_g N_VGND_c_641_n 0.00758038f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A2_M1018_g N_VGND_c_641_n 5.37623e-19 $X=3.08 $Y=0.655 $X2=0 $Y2=0
cc_223 N_A2_M1016_g N_VGND_c_642_n 5.37623e-19 $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_224 N_A2_M1018_g N_VGND_c_642_n 0.00750039f $X=3.08 $Y=0.655 $X2=0 $Y2=0
cc_225 N_A2_M1004_g N_VGND_c_645_n 0.00365202f $X=1.79 $Y=0.655 $X2=0 $Y2=0
cc_226 N_A2_M1008_g N_VGND_c_645_n 0.00365202f $X=2.22 $Y=0.655 $X2=0 $Y2=0
cc_227 N_A2_M1016_g N_VGND_c_647_n 0.00365202f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_228 N_A2_M1018_g N_VGND_c_647_n 0.00365202f $X=3.08 $Y=0.655 $X2=0 $Y2=0
cc_229 N_A2_M1004_g N_VGND_c_651_n 0.00432244f $X=1.79 $Y=0.655 $X2=0 $Y2=0
cc_230 N_A2_M1008_g N_VGND_c_651_n 0.00432244f $X=2.22 $Y=0.655 $X2=0 $Y2=0
cc_231 N_A2_M1016_g N_VGND_c_651_n 0.00432244f $X=2.65 $Y=0.655 $X2=0 $Y2=0
cc_232 N_A2_M1018_g N_VGND_c_651_n 0.00432244f $X=3.08 $Y=0.655 $X2=0 $Y2=0
cc_233 N_B1_M1002_g N_VPWR_c_357_n 0.0126366f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_234 N_B1_M1007_g N_VPWR_c_357_n 6.51893e-19 $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_235 N_B1_M1002_g N_VPWR_c_358_n 7.33921e-19 $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_236 N_B1_M1007_g N_VPWR_c_358_n 0.0142652f $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B1_M1017_g N_VPWR_c_358_n 0.0142189f $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B1_M1023_g N_VPWR_c_358_n 7.27171e-19 $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B1_M1017_g N_VPWR_c_360_n 7.24342e-19 $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B1_M1023_g N_VPWR_c_360_n 0.0151914f $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B1_M1002_g N_VPWR_c_363_n 0.00564095f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B1_M1007_g N_VPWR_c_363_n 0.00486043f $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B1_M1017_g N_VPWR_c_364_n 0.00486043f $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B1_M1023_g N_VPWR_c_364_n 0.00486043f $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B1_M1002_g N_VPWR_c_353_n 0.00948291f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B1_M1007_g N_VPWR_c_353_n 0.00824727f $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B1_M1017_g N_VPWR_c_353_n 0.00824727f $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B1_M1023_g N_VPWR_c_353_n 0.00824727f $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_249 N_B1_c_286_n N_Y_c_481_n 0.0127649f $X=4.41 $Y=1.185 $X2=0 $Y2=0
cc_250 N_B1_c_288_n N_Y_c_481_n 0.012674f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_251 N_B1_c_290_n N_Y_c_481_n 0.0166105f $X=5.27 $Y=1.185 $X2=0 $Y2=0
cc_252 B1 N_Y_c_481_n 0.0709722f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_253 N_B1_c_293_n N_Y_c_481_n 0.007f $X=5.27 $Y=1.35 $X2=0 $Y2=0
cc_254 N_B1_M1007_g N_Y_c_482_n 0.0193587f $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_255 N_B1_M1017_g N_Y_c_482_n 0.0194f $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_256 B1 N_Y_c_482_n 0.0725729f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_257 N_B1_c_293_n N_Y_c_482_n 0.00250517f $X=5.27 $Y=1.35 $X2=0 $Y2=0
cc_258 N_B1_M1002_g N_Y_c_483_n 0.024311f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_259 B1 N_Y_c_483_n 0.0306136f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_260 N_B1_c_293_n N_Y_c_483_n 0.00256759f $X=5.27 $Y=1.35 $X2=0 $Y2=0
cc_261 N_B1_M1023_g N_Y_c_484_n 0.0232098f $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_262 N_B1_c_293_n N_Y_c_484_n 0.00250517f $X=5.27 $Y=1.35 $X2=0 $Y2=0
cc_263 N_B1_c_290_n Y 0.0212627f $X=5.27 $Y=1.185 $X2=0 $Y2=0
cc_264 B1 Y 0.0183002f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_265 N_B1_c_284_n N_A_32_47#_c_588_n 8.27067e-19 $X=3.98 $Y=1.185 $X2=0 $Y2=0
cc_266 N_B1_c_284_n N_A_32_47#_c_578_n 0.00570825f $X=3.98 $Y=1.185 $X2=0 $Y2=0
cc_267 N_B1_c_286_n N_A_32_47#_c_578_n 7.65258e-19 $X=4.41 $Y=1.185 $X2=0 $Y2=0
cc_268 B1 N_A_32_47#_c_578_n 0.00118347f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_269 N_B1_c_284_n N_A_32_47#_c_562_n 0.0133145f $X=3.98 $Y=1.185 $X2=0 $Y2=0
cc_270 N_B1_c_286_n N_A_32_47#_c_562_n 0.0103812f $X=4.41 $Y=1.185 $X2=0 $Y2=0
cc_271 N_B1_c_288_n N_A_32_47#_c_562_n 0.0104569f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_272 N_B1_c_290_n N_A_32_47#_c_562_n 0.0104569f $X=5.27 $Y=1.185 $X2=0 $Y2=0
cc_273 N_B1_c_284_n N_VGND_c_650_n 0.00357842f $X=3.98 $Y=1.185 $X2=0 $Y2=0
cc_274 N_B1_c_286_n N_VGND_c_650_n 0.00357877f $X=4.41 $Y=1.185 $X2=0 $Y2=0
cc_275 N_B1_c_288_n N_VGND_c_650_n 0.00357877f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_276 N_B1_c_290_n N_VGND_c_650_n 0.00357877f $X=5.27 $Y=1.185 $X2=0 $Y2=0
cc_277 N_B1_c_284_n N_VGND_c_651_n 0.00537652f $X=3.98 $Y=1.185 $X2=0 $Y2=0
cc_278 N_B1_c_286_n N_VGND_c_651_n 0.0053512f $X=4.41 $Y=1.185 $X2=0 $Y2=0
cc_279 N_B1_c_288_n N_VGND_c_651_n 0.0053512f $X=4.84 $Y=1.185 $X2=0 $Y2=0
cc_280 N_B1_c_290_n N_VGND_c_651_n 0.00636493f $X=5.27 $Y=1.185 $X2=0 $Y2=0
cc_281 N_VPWR_c_353_n N_A_115_367#_M1006_s 0.00380103f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_282 N_VPWR_c_353_n N_A_115_367#_M1013_s 0.00376627f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_353_n N_A_115_367#_M1005_d 0.00223565f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_353_n N_A_115_367#_M1021_d 0.00307052f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_361_n N_A_115_367#_c_460_n 0.0140491f $X=0.98 $Y=3.33 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_353_n N_A_115_367#_c_460_n 0.0090585f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_287 N_VPWR_M1012_d N_A_115_367#_c_441_n 0.00176461f $X=1.005 $Y=1.835 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_356_n N_A_115_367#_c_441_n 0.0170777f $X=1.145 $Y=2.18 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_355_n N_A_115_367#_c_442_n 0.00581759f $X=0.285 $Y=1.98 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_362_n N_A_115_367#_c_465_n 0.0125234f $X=3.58 $Y=3.33 $X2=0
+ $Y2=0
cc_291 N_VPWR_c_353_n N_A_115_367#_c_465_n 0.00738676f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_362_n N_A_115_367#_c_452_n 0.0361172f $X=3.58 $Y=3.33 $X2=0
+ $Y2=0
cc_293 N_VPWR_c_353_n N_A_115_367#_c_452_n 0.023676f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_294 N_VPWR_c_362_n N_A_115_367#_c_454_n 0.0493502f $X=3.58 $Y=3.33 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_353_n N_A_115_367#_c_454_n 0.0318403f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_362_n N_A_115_367#_c_471_n 0.0125234f $X=3.58 $Y=3.33 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_353_n N_A_115_367#_c_471_n 0.00738676f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_353_n N_Y_M1001_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_299 N_VPWR_c_353_n N_Y_M1010_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_300 N_VPWR_c_353_n N_Y_M1002_d 0.00467071f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_301 N_VPWR_c_353_n N_Y_M1017_d 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_302 N_VPWR_c_363_n N_Y_c_532_n 0.0131621f $X=4.46 $Y=3.33 $X2=0 $Y2=0
cc_303 N_VPWR_c_353_n N_Y_c_532_n 0.00808656f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_304 N_VPWR_M1007_s N_Y_c_482_n 0.0017993f $X=4.485 $Y=1.835 $X2=0 $Y2=0
cc_305 N_VPWR_c_358_n N_Y_c_482_n 0.0178454f $X=4.625 $Y=2.19 $X2=0 $Y2=0
cc_306 N_VPWR_M1020_d N_Y_c_483_n 0.00223295f $X=3.585 $Y=1.835 $X2=0 $Y2=0
cc_307 N_VPWR_c_357_n N_Y_c_483_n 0.0182522f $X=3.745 $Y=2.4 $X2=0 $Y2=0
cc_308 N_VPWR_c_364_n N_Y_c_538_n 0.0124525f $X=5.32 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_c_353_n N_Y_c_538_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_310 N_VPWR_M1023_s N_Y_c_484_n 0.00272817f $X=5.345 $Y=1.835 $X2=0 $Y2=0
cc_311 N_VPWR_c_360_n N_Y_c_484_n 0.0220268f $X=5.485 $Y=2.19 $X2=0 $Y2=0
cc_312 N_A_115_367#_c_452_n N_Y_M1001_s 0.00332344f $X=2.34 $Y=2.99 $X2=0 $Y2=0
cc_313 N_A_115_367#_c_454_n N_Y_M1010_s 0.00332344f $X=3.2 $Y=2.99 $X2=0 $Y2=0
cc_314 N_A_115_367#_M1005_d N_Y_c_494_n 0.00333177f $X=2.295 $Y=1.835 $X2=0
+ $Y2=0
cc_315 N_A_115_367#_c_476_p N_Y_c_494_n 0.0135055f $X=2.435 $Y=2.435 $X2=0 $Y2=0
cc_316 N_A_115_367#_M1021_d N_Y_c_488_n 0.0060555f $X=3.155 $Y=1.835 $X2=0 $Y2=0
cc_317 N_A_115_367#_c_478_p N_Y_c_488_n 0.0135055f $X=3.295 $Y=2.435 $X2=0 $Y2=0
cc_318 N_A_115_367#_c_452_n N_Y_c_502_n 0.0159805f $X=2.34 $Y=2.99 $X2=0 $Y2=0
cc_319 N_A_115_367#_c_454_n N_Y_c_493_n 0.0159805f $X=3.2 $Y=2.99 $X2=0 $Y2=0
cc_320 N_Y_c_481_n N_A_32_47#_M1003_s 0.003358f $X=5.425 $Y=0.865 $X2=0 $Y2=0
cc_321 N_Y_c_481_n N_A_32_47#_M1014_s 0.00417968f $X=5.425 $Y=0.865 $X2=0 $Y2=0
cc_322 Y N_A_32_47#_M1014_s 7.1606e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_323 N_Y_M1000_d N_A_32_47#_c_562_n 0.00329779f $X=4.055 $Y=0.235 $X2=0 $Y2=0
cc_324 N_Y_M1009_d N_A_32_47#_c_562_n 0.00329779f $X=4.915 $Y=0.235 $X2=0 $Y2=0
cc_325 N_Y_c_481_n N_A_32_47#_c_562_n 0.0893572f $X=5.425 $Y=0.865 $X2=0 $Y2=0
cc_326 N_Y_c_481_n N_VGND_c_650_n 3.55955e-19 $X=5.425 $Y=0.865 $X2=0 $Y2=0
cc_327 N_Y_M1000_d N_VGND_c_651_n 0.00225186f $X=4.055 $Y=0.235 $X2=0 $Y2=0
cc_328 N_Y_M1009_d N_VGND_c_651_n 0.00225186f $X=4.915 $Y=0.235 $X2=0 $Y2=0
cc_329 N_Y_c_481_n N_VGND_c_651_n 0.00109701f $X=5.425 $Y=0.865 $X2=0 $Y2=0
cc_330 N_A_32_47#_c_564_n N_VGND_M1011_d 0.00329816f $X=1.05 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_331 N_A_32_47#_c_570_n N_VGND_M1019_d 0.00349176f $X=1.91 $Y=0.82 $X2=0 $Y2=0
cc_332 N_A_32_47#_c_573_n N_VGND_M1008_d 0.00335437f $X=2.77 $Y=0.82 $X2=0 $Y2=0
cc_333 N_A_32_47#_c_574_n N_VGND_M1018_d 0.00423083f $X=3.63 $Y=0.82 $X2=0 $Y2=0
cc_334 N_A_32_47#_c_564_n N_VGND_c_639_n 0.0170777f $X=1.05 $Y=0.955 $X2=0 $Y2=0
cc_335 N_A_32_47#_c_570_n N_VGND_c_640_n 0.016459f $X=1.91 $Y=0.82 $X2=0 $Y2=0
cc_336 N_A_32_47#_c_573_n N_VGND_c_641_n 0.016459f $X=2.77 $Y=0.82 $X2=0 $Y2=0
cc_337 N_A_32_47#_c_574_n N_VGND_c_642_n 0.0178756f $X=3.63 $Y=0.82 $X2=0 $Y2=0
cc_338 N_A_32_47#_c_610_p N_VGND_c_643_n 0.0124525f $X=1.145 $Y=0.43 $X2=0 $Y2=0
cc_339 N_A_32_47#_c_570_n N_VGND_c_643_n 0.00188649f $X=1.91 $Y=0.82 $X2=0 $Y2=0
cc_340 N_A_32_47#_c_570_n N_VGND_c_645_n 0.00196209f $X=1.91 $Y=0.82 $X2=0 $Y2=0
cc_341 N_A_32_47#_c_613_p N_VGND_c_645_n 0.0124139f $X=2.005 $Y=0.42 $X2=0 $Y2=0
cc_342 N_A_32_47#_c_573_n N_VGND_c_645_n 0.00196209f $X=2.77 $Y=0.82 $X2=0 $Y2=0
cc_343 N_A_32_47#_c_573_n N_VGND_c_647_n 0.00196209f $X=2.77 $Y=0.82 $X2=0 $Y2=0
cc_344 N_A_32_47#_c_616_p N_VGND_c_647_n 0.0124139f $X=2.865 $Y=0.42 $X2=0 $Y2=0
cc_345 N_A_32_47#_c_574_n N_VGND_c_647_n 0.00196209f $X=3.63 $Y=0.82 $X2=0 $Y2=0
cc_346 N_A_32_47#_c_560_n N_VGND_c_649_n 0.0178111f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_347 N_A_32_47#_c_574_n N_VGND_c_650_n 0.00210007f $X=3.63 $Y=0.82 $X2=0 $Y2=0
cc_348 N_A_32_47#_c_588_n N_VGND_c_650_n 0.017167f $X=3.78 $Y=0.53 $X2=0 $Y2=0
cc_349 N_A_32_47#_c_562_n N_VGND_c_650_n 0.0993812f $X=5.485 $Y=0.435 $X2=0
+ $Y2=0
cc_350 N_A_32_47#_M1011_s N_VGND_c_651_n 0.00371702f $X=0.16 $Y=0.235 $X2=0
+ $Y2=0
cc_351 N_A_32_47#_M1015_s N_VGND_c_651_n 0.00400238f $X=1.005 $Y=0.235 $X2=0
+ $Y2=0
cc_352 N_A_32_47#_M1004_s N_VGND_c_651_n 0.00266476f $X=1.865 $Y=0.235 $X2=0
+ $Y2=0
cc_353 N_A_32_47#_M1016_s N_VGND_c_651_n 0.00266476f $X=2.725 $Y=0.235 $X2=0
+ $Y2=0
cc_354 N_A_32_47#_M1022_s N_VGND_c_651_n 0.00220342f $X=3.625 $Y=0.235 $X2=0
+ $Y2=0
cc_355 N_A_32_47#_M1003_s N_VGND_c_651_n 0.00223577f $X=4.485 $Y=0.235 $X2=0
+ $Y2=0
cc_356 N_A_32_47#_M1014_s N_VGND_c_651_n 0.00215176f $X=5.345 $Y=0.235 $X2=0
+ $Y2=0
cc_357 N_A_32_47#_c_560_n N_VGND_c_651_n 0.0100304f $X=0.285 $Y=0.42 $X2=0 $Y2=0
cc_358 N_A_32_47#_c_610_p N_VGND_c_651_n 0.00730901f $X=1.145 $Y=0.43 $X2=0
+ $Y2=0
cc_359 N_A_32_47#_c_570_n N_VGND_c_651_n 0.00865724f $X=1.91 $Y=0.82 $X2=0 $Y2=0
cc_360 N_A_32_47#_c_613_p N_VGND_c_651_n 0.00730033f $X=2.005 $Y=0.42 $X2=0
+ $Y2=0
cc_361 N_A_32_47#_c_573_n N_VGND_c_651_n 0.00891615f $X=2.77 $Y=0.82 $X2=0 $Y2=0
cc_362 N_A_32_47#_c_616_p N_VGND_c_651_n 0.00730033f $X=2.865 $Y=0.42 $X2=0
+ $Y2=0
cc_363 N_A_32_47#_c_574_n N_VGND_c_651_n 0.0087269f $X=3.63 $Y=0.82 $X2=0 $Y2=0
cc_364 N_A_32_47#_c_588_n N_VGND_c_651_n 0.011462f $X=3.78 $Y=0.53 $X2=0 $Y2=0
cc_365 N_A_32_47#_c_562_n N_VGND_c_651_n 0.0625136f $X=5.485 $Y=0.435 $X2=0
+ $Y2=0
cc_366 N_A_32_47#_c_580_n N_VGND_c_651_n 2.38061e-19 $X=1.15 $Y=0.82 $X2=0 $Y2=0
