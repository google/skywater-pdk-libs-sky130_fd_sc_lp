* File: sky130_fd_sc_lp__clkbuf_2.pxi.spice
* Created: Fri Aug 28 10:14:55 2020
* 
x_PM_SKY130_FD_SC_LP__CLKBUF_2%A N_A_M1002_g N_A_M1005_g A N_A_c_41_n N_A_c_42_n
+ PM_SKY130_FD_SC_LP__CLKBUF_2%A
x_PM_SKY130_FD_SC_LP__CLKBUF_2%A_27_47# N_A_27_47#_M1002_s N_A_27_47#_M1005_s
+ N_A_27_47#_M1000_g N_A_27_47#_M1001_g N_A_27_47#_M1003_g N_A_27_47#_M1004_g
+ N_A_27_47#_c_74_n N_A_27_47#_c_75_n N_A_27_47#_c_76_n N_A_27_47#_c_77_n
+ N_A_27_47#_c_78_n N_A_27_47#_c_79_n PM_SKY130_FD_SC_LP__CLKBUF_2%A_27_47#
x_PM_SKY130_FD_SC_LP__CLKBUF_2%VPWR N_VPWR_M1005_d N_VPWR_M1003_d N_VPWR_c_134_n
+ N_VPWR_c_135_n N_VPWR_c_136_n VPWR N_VPWR_c_137_n N_VPWR_c_138_n
+ N_VPWR_c_139_n N_VPWR_c_133_n PM_SKY130_FD_SC_LP__CLKBUF_2%VPWR
x_PM_SKY130_FD_SC_LP__CLKBUF_2%X N_X_M1001_d N_X_M1000_s N_X_c_183_n X X X X X
+ N_X_c_161_n X PM_SKY130_FD_SC_LP__CLKBUF_2%X
x_PM_SKY130_FD_SC_LP__CLKBUF_2%VGND N_VGND_M1002_d N_VGND_M1004_s N_VGND_c_192_n
+ N_VGND_c_193_n N_VGND_c_194_n VGND N_VGND_c_195_n N_VGND_c_196_n
+ N_VGND_c_197_n N_VGND_c_198_n PM_SKY130_FD_SC_LP__CLKBUF_2%VGND
cc_1 VNB N_A_M1005_g 0.0324622f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB A 0.00618067f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_3 VNB N_A_c_41_n 0.0314602f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.94
cc_4 VNB N_A_c_42_n 0.0206597f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.775
cc_5 VNB N_A_27_47#_M1000_g 0.00591171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_M1001_g 0.0390592f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.775
cc_7 VNB N_A_27_47#_M1003_g 0.00676096f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.94
cc_8 VNB N_A_27_47#_M1004_g 0.0481464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_74_n 0.0313161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_75_n 0.00614616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_76_n 0.00732776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_77_n 0.0135923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_78_n 0.0137262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_79_n 0.0417084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_133_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB X 0.0266039f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.94
cc_17 VNB X 0.0256069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_X_c_161_n 0.00343837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_192_n 0.00475331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_193_n 0.0131412f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.94
cc_21 VNB N_VGND_c_194_n 0.00465501f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.775
cc_22 VNB N_VGND_c_195_n 0.0169874f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.94
cc_23 VNB N_VGND_c_196_n 0.0180813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_197_n 0.00526407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_198_n 0.129078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VPB N_A_M1005_g 0.0240578f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_27 VPB N_A_27_47#_M1000_g 0.0206827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_A_27_47#_M1003_g 0.0239324f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.94
cc_29 VPB N_A_27_47#_c_75_n 0.0573584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_134_n 0.0048939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_135_n 0.0131407f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.775
cc_32 VPB N_VPWR_c_136_n 0.0417147f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.94
cc_33 VPB N_VPWR_c_137_n 0.0173901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_138_n 0.0166894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_139_n 0.00593688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_133_n 0.0474653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB X 0.00414482f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB X 0.0157086f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.94
cc_39 N_A_M1005_g N_A_27_47#_M1001_g 0.00389195f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_40 A N_A_27_47#_M1001_g 0.00253307f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_41 N_A_c_41_n N_A_27_47#_M1001_g 0.0192761f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_42 N_A_c_42_n N_A_27_47#_M1001_g 0.0105633f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_43 N_A_M1005_g N_A_27_47#_c_74_n 0.00594476f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_44 A N_A_27_47#_c_74_n 0.0253686f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_45 N_A_c_41_n N_A_27_47#_c_74_n 0.00816168f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_46 N_A_c_42_n N_A_27_47#_c_74_n 0.00544175f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_47 N_A_M1005_g N_A_27_47#_c_75_n 0.013199f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_48 N_A_M1005_g N_A_27_47#_c_76_n 0.0222055f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_49 A N_A_27_47#_c_76_n 0.0352792f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_50 N_A_c_41_n N_A_27_47#_c_76_n 0.00300839f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_51 N_A_c_41_n N_A_27_47#_c_78_n 0.00165146f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_52 N_A_M1005_g N_A_27_47#_c_79_n 0.0318729f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_53 N_A_M1005_g N_VPWR_c_134_n 0.00361965f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_54 N_A_M1005_g N_VPWR_c_137_n 0.00585385f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_55 N_A_M1005_g N_VPWR_c_133_n 0.0119078f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_56 A X 0.0293323f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_57 A N_VGND_c_192_n 0.0201833f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_58 N_A_c_41_n N_VGND_c_192_n 0.00261478f $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_59 N_A_c_42_n N_VGND_c_192_n 0.00328447f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_60 N_A_c_41_n N_VGND_c_195_n 3.60471e-19 $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_61 N_A_c_42_n N_VGND_c_195_n 0.00585385f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_62 A N_VGND_c_198_n 0.00678453f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_63 N_A_c_41_n N_VGND_c_198_n 4.44682e-19 $X=0.51 $Y=0.94 $X2=0 $Y2=0
cc_64 N_A_c_42_n N_VGND_c_198_n 0.00798939f $X=0.51 $Y=0.775 $X2=0 $Y2=0
cc_65 N_A_27_47#_M1000_g N_VPWR_c_134_n 0.00218819f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_66 N_A_27_47#_c_76_n N_VPWR_c_134_n 0.013485f $X=1.05 $Y=1.38 $X2=0 $Y2=0
cc_67 N_A_27_47#_M1003_g N_VPWR_c_136_n 0.00338307f $X=1.385 $Y=2.465 $X2=0
+ $Y2=0
cc_68 N_A_27_47#_c_75_n N_VPWR_c_137_n 0.0167439f $X=0.26 $Y=2.04 $X2=0 $Y2=0
cc_69 N_A_27_47#_M1000_g N_VPWR_c_138_n 0.00585385f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_70 N_A_27_47#_M1003_g N_VPWR_c_138_n 0.00585385f $X=1.385 $Y=2.465 $X2=0
+ $Y2=0
cc_71 N_A_27_47#_M1005_s N_VPWR_c_133_n 0.00238045f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_72 N_A_27_47#_M1000_g N_VPWR_c_133_n 0.0108762f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_73 N_A_27_47#_M1003_g N_VPWR_c_133_n 0.0116285f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_74 N_A_27_47#_c_75_n N_VPWR_c_133_n 0.0117986f $X=0.26 $Y=2.04 $X2=0 $Y2=0
cc_75 N_A_27_47#_M1001_g X 0.00286296f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_76 N_A_27_47#_M1004_g X 0.0202469f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A_27_47#_c_76_n X 0.0132093f $X=1.05 $Y=1.38 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_79_n X 0.00257088f $X=1.385 $Y=1.375 $X2=0 $Y2=0
cc_79 N_A_27_47#_M1000_g X 9.57063e-19 $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A_27_47#_M1001_g X 5.34577e-19 $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_81 N_A_27_47#_M1003_g X 0.00801994f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A_27_47#_M1004_g X 0.004586f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_76_n X 0.0209967f $X=1.05 $Y=1.38 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_79_n X 0.0171711f $X=1.385 $Y=1.375 $X2=0 $Y2=0
cc_85 N_A_27_47#_M1000_g X 0.00194942f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A_27_47#_M1003_g X 0.0159432f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_75_n X 0.00364441f $X=0.26 $Y=2.04 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_76_n X 0.0115429f $X=1.05 $Y=1.38 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_79_n X 0.00231511f $X=1.385 $Y=1.375 $X2=0 $Y2=0
cc_90 N_A_27_47#_M1001_g N_X_c_161_n 0.00349558f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_27_47#_M1004_g N_X_c_161_n 0.00349558f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_27_47#_M1001_g N_VGND_c_192_n 0.00163339f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_27_47#_M1004_g N_VGND_c_194_n 0.00375674f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_77_n N_VGND_c_195_n 0.0175785f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_95 N_A_27_47#_M1001_g N_VGND_c_196_n 0.00585385f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_27_47#_M1004_g N_VGND_c_196_n 0.00585385f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_27_47#_M1002_s N_VGND_c_198_n 0.00231961f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_M1001_g N_VGND_c_198_n 0.0109324f $X=0.96 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_27_47#_M1004_g N_VGND_c_198_n 0.00718088f $X=1.39 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_77_n N_VGND_c_198_n 0.0113939f $X=0.26 $Y=0.44 $X2=0 $Y2=0
cc_101 N_VPWR_c_133_n N_X_M1000_s 0.00302905f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_102 N_VPWR_c_138_n N_X_c_183_n 0.012556f $X=1.475 $Y=3.33 $X2=0 $Y2=0
cc_103 N_VPWR_c_133_n N_X_c_183_n 0.00988321f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_104 N_VPWR_M1003_d X 0.00248866f $X=1.46 $Y=1.835 $X2=0 $Y2=0
cc_105 N_VPWR_c_136_n X 0.0172604f $X=1.6 $Y=2.23 $X2=0 $Y2=0
cc_106 X N_VGND_c_194_n 0.0192273f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_107 N_X_c_161_n N_VGND_c_196_n 0.0138306f $X=1.175 $Y=0.44 $X2=0 $Y2=0
cc_108 N_X_M1001_d N_VGND_c_198_n 0.00260039f $X=1.035 $Y=0.235 $X2=0 $Y2=0
cc_109 X N_VGND_c_198_n 0.00973077f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_110 N_X_c_161_n N_VGND_c_198_n 0.00990886f $X=1.175 $Y=0.44 $X2=0 $Y2=0
