* File: sky130_fd_sc_lp__a41oi_0.pxi.spice
* Created: Fri Aug 28 10:03:16 2020
* 
x_PM_SKY130_FD_SC_LP__A41OI_0%B1 N_B1_M1006_g N_B1_c_72_n N_B1_M1001_g
+ N_B1_c_77_n B1 B1 N_B1_c_74_n PM_SKY130_FD_SC_LP__A41OI_0%B1
x_PM_SKY130_FD_SC_LP__A41OI_0%A1 N_A1_c_108_n N_A1_M1007_g N_A1_M1009_g
+ N_A1_c_110_n N_A1_c_111_n N_A1_c_116_n A1 A1 A1 N_A1_c_113_n
+ PM_SKY130_FD_SC_LP__A41OI_0%A1
x_PM_SKY130_FD_SC_LP__A41OI_0%A2 N_A2_M1005_g N_A2_M1004_g N_A2_c_159_n
+ N_A2_c_160_n A2 A2 A2 N_A2_c_162_n PM_SKY130_FD_SC_LP__A41OI_0%A2
x_PM_SKY130_FD_SC_LP__A41OI_0%A3 N_A3_M1003_g N_A3_M1000_g N_A3_c_201_n
+ N_A3_c_202_n A3 A3 A3 N_A3_c_204_n PM_SKY130_FD_SC_LP__A41OI_0%A3
x_PM_SKY130_FD_SC_LP__A41OI_0%A4 N_A4_M1002_g N_A4_M1008_g N_A4_c_242_n
+ N_A4_c_249_n N_A4_c_243_n N_A4_c_244_n A4 A4 N_A4_c_246_n
+ PM_SKY130_FD_SC_LP__A41OI_0%A4
x_PM_SKY130_FD_SC_LP__A41OI_0%Y N_Y_M1006_d N_Y_M1001_s N_Y_c_278_n N_Y_c_282_n
+ N_Y_c_277_n N_Y_c_279_n Y Y Y Y PM_SKY130_FD_SC_LP__A41OI_0%Y
x_PM_SKY130_FD_SC_LP__A41OI_0%A_176_479# N_A_176_479#_M1001_d
+ N_A_176_479#_M1004_d N_A_176_479#_M1002_d N_A_176_479#_c_318_n
+ N_A_176_479#_c_319_n N_A_176_479#_c_320_n N_A_176_479#_c_321_n
+ N_A_176_479#_c_322_n N_A_176_479#_c_323_n N_A_176_479#_c_324_n
+ PM_SKY130_FD_SC_LP__A41OI_0%A_176_479#
x_PM_SKY130_FD_SC_LP__A41OI_0%VPWR N_VPWR_M1009_d N_VPWR_M1000_d N_VPWR_c_363_n
+ N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_368_n
+ VPWR N_VPWR_c_369_n N_VPWR_c_362_n PM_SKY130_FD_SC_LP__A41OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A41OI_0%VGND N_VGND_M1006_s N_VGND_M1008_d N_VGND_c_399_n
+ N_VGND_c_400_n N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n VGND
+ N_VGND_c_404_n N_VGND_c_405_n PM_SKY130_FD_SC_LP__A41OI_0%VGND
cc_1 VNB N_B1_M1006_g 0.0271356f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_2 VNB N_B1_c_72_n 0.013038f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.735
cc_3 VNB B1 0.0444968f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_4 VNB N_B1_c_74_n 0.0790488f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.99
cc_5 VNB N_A1_c_108_n 0.0203758f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_6 VNB N_A1_M1007_g 0.0209123f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.495
cc_7 VNB N_A1_c_110_n 0.0186724f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.81
cc_8 VNB N_A1_c_111_n 0.00809342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A1 0.0079775f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_A1_c_113_n 0.0176171f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.495
cc_11 VNB N_A2_M1005_g 0.0215667f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_12 VNB N_A2_M1004_g 0.00719763f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.885
cc_13 VNB N_A2_c_159_n 0.0213471f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.81
cc_14 VNB N_A2_c_160_n 0.0159874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A2 0.00832635f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.81
cc_16 VNB N_A2_c_162_n 0.0155581f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.99
cc_17 VNB N_A3_M1003_g 0.0227994f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.445
cc_18 VNB N_A3_M1000_g 0.00842589f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.885
cc_19 VNB N_A3_c_201_n 0.021772f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.81
cc_20 VNB N_A3_c_202_n 0.0157662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A3 0.00759993f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.81
cc_22 VNB N_A3_c_204_n 0.0157662f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.99
cc_23 VNB N_A4_M1008_g 0.0350944f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.885
cc_24 VNB N_A4_c_242_n 0.00432856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A4_c_243_n 0.025421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A4_c_244_n 0.0181362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A4 0.0489426f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.99
cc_28 VNB N_A4_c_246_n 0.0198547f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.295
cc_29 VNB N_Y_c_277_n 0.00657331f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.81
cc_30 VNB N_VPWR_c_362_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_399_n 0.0139338f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.885
cc_32 VNB N_VGND_c_400_n 0.00488208f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.715
cc_33 VNB N_VGND_c_401_n 0.0176306f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.81
cc_34 VNB N_VGND_c_402_n 0.0549127f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_35 VNB N_VGND_c_403_n 0.00510915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_404_n 0.0121672f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.295
cc_37 VNB N_VGND_c_405_n 0.198144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_B1_c_72_n 0.00555508f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.735
cc_39 VPB N_B1_M1001_g 0.042259f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.715
cc_40 VPB N_B1_c_77_n 0.028519f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=1.81
cc_41 VPB N_A1_M1009_g 0.0366921f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.81
cc_42 VPB N_A1_c_111_n 0.00402126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A1_c_116_n 0.0113866f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_44 VPB A1 0.00375002f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_45 VPB N_A2_M1004_g 0.0472938f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=1.885
cc_46 VPB A2 0.00395677f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=1.81
cc_47 VPB N_A3_M1000_g 0.0484807f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=1.885
cc_48 VPB A3 0.00289349f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=1.81
cc_49 VPB N_A4_M1002_g 0.0462564f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.445
cc_50 VPB N_A4_c_242_n 0.00495589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A4_c_249_n 0.0224078f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=1.81
cc_52 VPB A4 0.026384f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.99
cc_53 VPB N_Y_c_278_n 0.0545917f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.715
cc_54 VPB N_Y_c_279_n 0.00741745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_176_479#_c_318_n 0.00560371f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_176_479#_c_319_n 0.00874824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_176_479#_c_320_n 0.00431928f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_58 VPB N_A_176_479#_c_321_n 0.00541639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_176_479#_c_322_n 0.0192209f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.99
cc_60 VPB N_A_176_479#_c_323_n 0.0369828f $X=-0.19 $Y=1.655 $X2=0.267 $Y2=0.925
cc_61 VPB N_A_176_479#_c_324_n 0.00713048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_363_n 0.00883076f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.715
cc_63 VPB N_VPWR_c_364_n 0.00909568f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=1.81
cc_64 VPB N_VPWR_c_365_n 0.0391634f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_65 VPB N_VPWR_c_366_n 0.00487897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_367_n 0.0166442f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=0.99
cc_67 VPB N_VPWR_c_368_n 0.00516749f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.99
cc_68 VPB N_VPWR_c_369_n 0.0286036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_362_n 0.084992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 N_B1_M1006_g N_A1_M1007_g 0.0171057f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_71 N_B1_M1001_g N_A1_M1009_g 0.0262792f $X=0.805 $Y=2.715 $X2=0 $Y2=0
cc_72 N_B1_c_72_n N_A1_c_111_n 0.00547115f $X=0.565 $Y=1.735 $X2=0 $Y2=0
cc_73 N_B1_c_77_n N_A1_c_116_n 0.00964291f $X=0.805 $Y=1.81 $X2=0 $Y2=0
cc_74 N_B1_c_72_n A1 6.4097e-19 $X=0.565 $Y=1.735 $X2=0 $Y2=0
cc_75 N_B1_c_77_n A1 6.89987e-19 $X=0.805 $Y=1.81 $X2=0 $Y2=0
cc_76 N_B1_c_74_n A1 5.18877e-19 $X=0.335 $Y=0.99 $X2=0 $Y2=0
cc_77 N_B1_c_74_n N_A1_c_113_n 0.0350537f $X=0.335 $Y=0.99 $X2=0 $Y2=0
cc_78 N_B1_M1001_g N_Y_c_278_n 0.0152774f $X=0.805 $Y=2.715 $X2=0 $Y2=0
cc_79 N_B1_c_77_n N_Y_c_278_n 0.00719654f $X=0.805 $Y=1.81 $X2=0 $Y2=0
cc_80 N_B1_M1006_g N_Y_c_282_n 0.00591525f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_81 N_B1_M1006_g N_Y_c_277_n 0.00848624f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_82 N_B1_c_72_n N_Y_c_277_n 0.00980186f $X=0.565 $Y=1.735 $X2=0 $Y2=0
cc_83 B1 N_Y_c_277_n 0.0488122f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_84 N_B1_c_74_n N_Y_c_277_n 0.0152086f $X=0.335 $Y=0.99 $X2=0 $Y2=0
cc_85 N_B1_c_72_n N_Y_c_279_n 0.00875574f $X=0.565 $Y=1.735 $X2=0 $Y2=0
cc_86 N_B1_c_77_n N_Y_c_279_n 0.0158729f $X=0.805 $Y=1.81 $X2=0 $Y2=0
cc_87 B1 N_Y_c_279_n 0.00188258f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_88 N_B1_c_74_n N_Y_c_279_n 0.00210326f $X=0.335 $Y=0.99 $X2=0 $Y2=0
cc_89 N_B1_M1001_g N_A_176_479#_c_318_n 0.00166989f $X=0.805 $Y=2.715 $X2=0
+ $Y2=0
cc_90 N_B1_M1001_g N_A_176_479#_c_320_n 0.00159959f $X=0.805 $Y=2.715 $X2=0
+ $Y2=0
cc_91 N_B1_M1001_g N_VPWR_c_365_n 0.00526658f $X=0.805 $Y=2.715 $X2=0 $Y2=0
cc_92 N_B1_M1001_g N_VPWR_c_362_n 0.0111317f $X=0.805 $Y=2.715 $X2=0 $Y2=0
cc_93 N_B1_M1006_g N_VGND_c_400_n 0.00482802f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_94 B1 N_VGND_c_400_n 0.0135105f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_95 N_B1_c_74_n N_VGND_c_400_n 0.00148503f $X=0.335 $Y=0.99 $X2=0 $Y2=0
cc_96 N_B1_M1006_g N_VGND_c_402_n 0.00555714f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_97 N_B1_M1006_g N_VGND_c_405_n 0.0113859f $X=0.565 $Y=0.445 $X2=0 $Y2=0
cc_98 B1 N_VGND_c_405_n 0.00684346f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_99 N_B1_c_74_n N_VGND_c_405_n 0.00102157f $X=0.335 $Y=0.99 $X2=0 $Y2=0
cc_100 N_A1_M1007_g N_A2_M1005_g 0.0311396f $X=1.075 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A1_c_111_n N_A2_M1004_g 0.00799879f $X=1.2 $Y=1.735 $X2=0 $Y2=0
cc_102 N_A1_c_116_n N_A2_M1004_g 0.0357318f $X=1.2 $Y=1.885 $X2=0 $Y2=0
cc_103 A1 N_A2_M1004_g 0.00111202f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_104 N_A1_c_108_n N_A2_c_159_n 0.0137892f $X=1.06 $Y=1.315 $X2=0 $Y2=0
cc_105 N_A1_c_110_n N_A2_c_160_n 0.0137892f $X=1.06 $Y=1.495 $X2=0 $Y2=0
cc_106 N_A1_c_111_n A2 6.68657e-19 $X=1.2 $Y=1.735 $X2=0 $Y2=0
cc_107 N_A1_c_116_n A2 3.26005e-19 $X=1.2 $Y=1.885 $X2=0 $Y2=0
cc_108 A1 A2 0.0823092f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_109 N_A1_c_113_n A2 5.82925e-19 $X=1.075 $Y=0.99 $X2=0 $Y2=0
cc_110 A1 N_A2_c_162_n 0.00448642f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_111 N_A1_c_113_n N_A2_c_162_n 0.0137892f $X=1.075 $Y=0.99 $X2=0 $Y2=0
cc_112 N_A1_M1007_g N_Y_c_277_n 0.00370037f $X=1.075 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A1_c_111_n N_Y_c_277_n 7.07997e-19 $X=1.2 $Y=1.735 $X2=0 $Y2=0
cc_114 A1 N_Y_c_277_n 0.0794386f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_115 N_A1_c_113_n N_Y_c_277_n 0.00487435f $X=1.075 $Y=0.99 $X2=0 $Y2=0
cc_116 N_A1_M1007_g Y 0.018758f $X=1.075 $Y=0.445 $X2=0 $Y2=0
cc_117 A1 Y 0.0272149f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_118 N_A1_c_113_n Y 0.00446517f $X=1.075 $Y=0.99 $X2=0 $Y2=0
cc_119 N_A1_M1009_g N_A_176_479#_c_318_n 0.00274279f $X=1.235 $Y=2.715 $X2=0
+ $Y2=0
cc_120 N_A1_M1009_g N_A_176_479#_c_319_n 0.0151764f $X=1.235 $Y=2.715 $X2=0
+ $Y2=0
cc_121 N_A1_c_116_n N_A_176_479#_c_319_n 2.72501e-19 $X=1.2 $Y=1.885 $X2=0 $Y2=0
cc_122 A1 N_A_176_479#_c_319_n 0.0153452f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_123 N_A1_c_110_n N_A_176_479#_c_320_n 0.00370497f $X=1.06 $Y=1.495 $X2=0
+ $Y2=0
cc_124 N_A1_c_116_n N_A_176_479#_c_320_n 0.00170844f $X=1.2 $Y=1.885 $X2=0 $Y2=0
cc_125 A1 N_A_176_479#_c_320_n 0.0137496f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_126 N_A1_M1009_g N_VPWR_c_363_n 0.00298143f $X=1.235 $Y=2.715 $X2=0 $Y2=0
cc_127 N_A1_M1009_g N_VPWR_c_365_n 0.00526658f $X=1.235 $Y=2.715 $X2=0 $Y2=0
cc_128 N_A1_M1009_g N_VPWR_c_362_n 0.0101042f $X=1.235 $Y=2.715 $X2=0 $Y2=0
cc_129 N_A1_M1007_g N_VGND_c_402_n 0.00363059f $X=1.075 $Y=0.445 $X2=0 $Y2=0
cc_130 N_A1_M1007_g N_VGND_c_405_n 0.0057288f $X=1.075 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A2_M1005_g N_A3_M1003_g 0.021237f $X=1.525 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A2_M1004_g N_A3_M1000_g 0.0440282f $X=1.665 $Y=2.715 $X2=0 $Y2=0
cc_133 N_A2_c_159_n N_A3_c_201_n 0.0117221f $X=1.615 $Y=1.33 $X2=0 $Y2=0
cc_134 N_A2_c_160_n N_A3_c_202_n 0.0117221f $X=1.615 $Y=1.495 $X2=0 $Y2=0
cc_135 N_A2_M1004_g A3 3.60022e-19 $X=1.665 $Y=2.715 $X2=0 $Y2=0
cc_136 A2 A3 0.0801159f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_137 N_A2_c_162_n A3 7.26553e-19 $X=1.615 $Y=0.99 $X2=0 $Y2=0
cc_138 A2 N_A3_c_204_n 0.00611808f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_139 N_A2_c_162_n N_A3_c_204_n 0.0117221f $X=1.615 $Y=0.99 $X2=0 $Y2=0
cc_140 N_A2_M1005_g Y 0.0221323f $X=1.525 $Y=0.445 $X2=0 $Y2=0
cc_141 A2 Y 0.0239579f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_142 N_A2_c_162_n Y 0.00118149f $X=1.615 $Y=0.99 $X2=0 $Y2=0
cc_143 N_A2_M1004_g N_A_176_479#_c_319_n 0.0154903f $X=1.665 $Y=2.715 $X2=0
+ $Y2=0
cc_144 N_A2_c_160_n N_A_176_479#_c_319_n 0.0025341f $X=1.615 $Y=1.495 $X2=0
+ $Y2=0
cc_145 A2 N_A_176_479#_c_319_n 0.0157906f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_146 N_A2_M1004_g N_A_176_479#_c_321_n 0.00277089f $X=1.665 $Y=2.715 $X2=0
+ $Y2=0
cc_147 A2 N_A_176_479#_c_324_n 0.0096157f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_148 N_A2_M1004_g N_VPWR_c_363_n 0.00170437f $X=1.665 $Y=2.715 $X2=0 $Y2=0
cc_149 N_A2_M1004_g N_VPWR_c_367_n 0.00526658f $X=1.665 $Y=2.715 $X2=0 $Y2=0
cc_150 N_A2_M1004_g N_VPWR_c_362_n 0.0101178f $X=1.665 $Y=2.715 $X2=0 $Y2=0
cc_151 N_A2_M1005_g N_VGND_c_402_n 0.00363059f $X=1.525 $Y=0.445 $X2=0 $Y2=0
cc_152 N_A2_M1005_g N_VGND_c_405_n 0.00585737f $X=1.525 $Y=0.445 $X2=0 $Y2=0
cc_153 N_A3_M1003_g N_A4_M1008_g 0.0199888f $X=2.095 $Y=0.445 $X2=0 $Y2=0
cc_154 A3 N_A4_M1008_g 0.00369748f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_155 N_A3_c_204_n N_A4_M1008_g 0.0120575f $X=2.185 $Y=0.99 $X2=0 $Y2=0
cc_156 N_A3_M1000_g N_A4_c_249_n 0.0354784f $X=2.095 $Y=2.715 $X2=0 $Y2=0
cc_157 A3 N_A4_c_249_n 8.02993e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_158 N_A3_c_202_n N_A4_c_243_n 0.0120575f $X=2.185 $Y=1.495 $X2=0 $Y2=0
cc_159 N_A3_M1000_g N_A4_c_244_n 0.00613141f $X=2.095 $Y=2.715 $X2=0 $Y2=0
cc_160 N_A3_M1000_g A4 7.80528e-19 $X=2.095 $Y=2.715 $X2=0 $Y2=0
cc_161 N_A3_c_201_n A4 0.00191531f $X=2.185 $Y=1.33 $X2=0 $Y2=0
cc_162 A3 A4 0.0740806f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_163 N_A3_c_201_n N_A4_c_246_n 0.0120575f $X=2.185 $Y=1.33 $X2=0 $Y2=0
cc_164 A3 N_A4_c_246_n 0.00223331f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_165 N_A3_M1003_g Y 0.0195375f $X=2.095 $Y=0.445 $X2=0 $Y2=0
cc_166 A3 Y 0.0238665f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_167 N_A3_c_204_n Y 0.00118269f $X=2.185 $Y=0.99 $X2=0 $Y2=0
cc_168 N_A3_M1000_g N_A_176_479#_c_321_n 0.00274545f $X=2.095 $Y=2.715 $X2=0
+ $Y2=0
cc_169 N_A3_M1000_g N_A_176_479#_c_322_n 0.0156717f $X=2.095 $Y=2.715 $X2=0
+ $Y2=0
cc_170 N_A3_c_202_n N_A_176_479#_c_322_n 6.05309e-19 $X=2.185 $Y=1.495 $X2=0
+ $Y2=0
cc_171 A3 N_A_176_479#_c_322_n 0.0249812f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_172 N_A3_M1000_g N_VPWR_c_364_n 0.00175636f $X=2.095 $Y=2.715 $X2=0 $Y2=0
cc_173 N_A3_M1000_g N_VPWR_c_367_n 0.00526658f $X=2.095 $Y=2.715 $X2=0 $Y2=0
cc_174 N_A3_M1000_g N_VPWR_c_362_n 0.0100905f $X=2.095 $Y=2.715 $X2=0 $Y2=0
cc_175 N_A3_M1003_g N_VGND_c_401_n 0.00131895f $X=2.095 $Y=0.445 $X2=0 $Y2=0
cc_176 N_A3_M1003_g N_VGND_c_402_n 0.00363059f $X=2.095 $Y=0.445 $X2=0 $Y2=0
cc_177 N_A3_M1003_g N_VGND_c_405_n 0.00612932f $X=2.095 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A4_M1008_g Y 0.00448127f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_179 N_A4_M1002_g N_A_176_479#_c_322_n 0.0189564f $X=2.525 $Y=2.715 $X2=0
+ $Y2=0
cc_180 N_A4_c_249_n N_A_176_479#_c_322_n 0.00397164f $X=2.665 $Y=1.81 $X2=0
+ $Y2=0
cc_181 N_A4_c_244_n N_A_176_479#_c_322_n 7.40865e-19 $X=2.755 $Y=1.585 $X2=0
+ $Y2=0
cc_182 A4 N_A_176_479#_c_322_n 0.0313306f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A4_M1002_g N_A_176_479#_c_323_n 0.00603396f $X=2.525 $Y=2.715 $X2=0
+ $Y2=0
cc_184 N_A4_M1002_g N_VPWR_c_364_n 0.00302979f $X=2.525 $Y=2.715 $X2=0 $Y2=0
cc_185 N_A4_M1002_g N_VPWR_c_369_n 0.00526658f $X=2.525 $Y=2.715 $X2=0 $Y2=0
cc_186 N_A4_M1002_g N_VPWR_c_362_n 0.0108747f $X=2.525 $Y=2.715 $X2=0 $Y2=0
cc_187 N_A4_M1008_g N_VGND_c_401_n 0.0120362f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_188 A4 N_VGND_c_401_n 0.0143781f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A4_c_246_n N_VGND_c_401_n 0.00431014f $X=2.755 $Y=1.08 $X2=0 $Y2=0
cc_190 N_A4_M1008_g N_VGND_c_402_n 0.00486043f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_191 N_A4_M1008_g N_VGND_c_405_n 0.00870566f $X=2.665 $Y=0.445 $X2=0 $Y2=0
cc_192 N_Y_c_278_n N_A_176_479#_c_318_n 0.0168148f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_193 N_Y_c_278_n N_A_176_479#_c_320_n 0.0157849f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_194 N_Y_c_278_n N_VPWR_c_365_n 0.0186437f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_195 N_Y_c_278_n N_VPWR_c_362_n 0.0112813f $X=0.59 $Y=2.54 $X2=0 $Y2=0
cc_196 Y N_VGND_c_401_n 0.0175619f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_197 N_Y_c_282_n N_VGND_c_402_n 0.0103546f $X=0.72 $Y=0.655 $X2=0 $Y2=0
cc_198 Y N_VGND_c_402_n 0.0819475f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_199 N_Y_M1006_d N_VGND_c_405_n 0.00290803f $X=0.64 $Y=0.235 $X2=0 $Y2=0
cc_200 N_Y_c_282_n N_VGND_c_405_n 0.0075774f $X=0.72 $Y=0.655 $X2=0 $Y2=0
cc_201 Y N_VGND_c_405_n 0.0581304f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_202 Y A_230_47# 0.00489519f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_203 Y A_320_47# 0.0107514f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_204 Y A_434_47# 0.0110636f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_205 N_A_176_479#_c_318_n N_VPWR_c_363_n 0.00304534f $X=1.02 $Y=2.54 $X2=0
+ $Y2=0
cc_206 N_A_176_479#_c_319_n N_VPWR_c_363_n 0.021452f $X=1.745 $Y=2.115 $X2=0
+ $Y2=0
cc_207 N_A_176_479#_c_321_n N_VPWR_c_363_n 0.00304534f $X=1.88 $Y=2.54 $X2=0
+ $Y2=0
cc_208 N_A_176_479#_c_321_n N_VPWR_c_364_n 0.00305856f $X=1.88 $Y=2.54 $X2=0
+ $Y2=0
cc_209 N_A_176_479#_c_322_n N_VPWR_c_364_n 0.0227239f $X=2.615 $Y=2.115 $X2=0
+ $Y2=0
cc_210 N_A_176_479#_c_323_n N_VPWR_c_364_n 0.00308399f $X=2.74 $Y=2.54 $X2=0
+ $Y2=0
cc_211 N_A_176_479#_c_318_n N_VPWR_c_365_n 0.0164167f $X=1.02 $Y=2.54 $X2=0
+ $Y2=0
cc_212 N_A_176_479#_c_321_n N_VPWR_c_367_n 0.0164167f $X=1.88 $Y=2.54 $X2=0
+ $Y2=0
cc_213 N_A_176_479#_c_323_n N_VPWR_c_369_n 0.0183256f $X=2.74 $Y=2.54 $X2=0
+ $Y2=0
cc_214 N_A_176_479#_c_318_n N_VPWR_c_362_n 0.00993371f $X=1.02 $Y=2.54 $X2=0
+ $Y2=0
cc_215 N_A_176_479#_c_321_n N_VPWR_c_362_n 0.00993371f $X=1.88 $Y=2.54 $X2=0
+ $Y2=0
cc_216 N_A_176_479#_c_323_n N_VPWR_c_362_n 0.0110888f $X=2.74 $Y=2.54 $X2=0
+ $Y2=0
cc_217 N_VGND_c_405_n A_230_47# 0.00242369f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_218 N_VGND_c_405_n A_320_47# 0.00341334f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_219 N_VGND_c_405_n A_434_47# 0.00946231f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
