# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o211ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o211ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.210000 1.345000 1.560000 1.630000 ;
        RECT 1.115000 1.630000 1.560000 1.925000 ;
        RECT 1.115000 1.925000 3.780000 2.120000 ;
        RECT 3.500000 1.345000 3.780000 1.925000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.855000 1.425000 3.330000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.950000 1.345000 5.125000 1.760000 ;
        RECT 4.955000 1.760000 5.125000 1.930000 ;
        RECT 4.955000 1.930000 7.720000 2.100000 ;
        RECT 7.390000 1.425000 7.720000 1.930000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.355000 1.425000 7.045000 1.760000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  2.587200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 2.290000 8.070000 2.440000 ;
        RECT 2.025000 2.440000 4.415000 2.510000 ;
        RECT 2.025000 2.510000 2.235000 2.630000 ;
        RECT 4.205000 2.510000 4.415000 3.075000 ;
        RECT 4.215000 1.930000 4.425000 2.270000 ;
        RECT 4.215000 2.270000 8.070000 2.290000 ;
        RECT 5.085000 2.440000 5.310000 3.075000 ;
        RECT 5.675000 0.965000 7.025000 1.075000 ;
        RECT 5.675000 1.075000 8.070000 1.255000 ;
        RECT 5.900000 2.440000 8.070000 2.505000 ;
        RECT 5.900000 2.505000 6.135000 3.075000 ;
        RECT 7.145000 2.505000 7.335000 3.075000 ;
        RECT 7.890000 1.255000 8.070000 2.270000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.245000  1.815000 0.535000 3.245000 ;
      RECT 0.305000  0.255000 0.505000 0.995000 ;
      RECT 0.305000  0.995000 4.915000 1.175000 ;
      RECT 0.675000  0.085000 1.005000 0.825000 ;
      RECT 0.705000  1.815000 0.925000 2.290000 ;
      RECT 0.705000  2.290000 1.805000 2.520000 ;
      RECT 0.705000  2.520000 0.925000 3.075000 ;
      RECT 1.105000  2.690000 1.435000 3.245000 ;
      RECT 1.175000  0.255000 1.365000 0.995000 ;
      RECT 1.535000  0.085000 1.865000 0.805000 ;
      RECT 1.605000  2.520000 1.805000 2.810000 ;
      RECT 1.605000  2.810000 3.525000 3.075000 ;
      RECT 2.035000  0.255000 2.225000 0.995000 ;
      RECT 2.395000  0.085000 2.725000 0.825000 ;
      RECT 2.895000  0.255000 3.085000 0.995000 ;
      RECT 3.255000  0.085000 3.585000 0.825000 ;
      RECT 3.315000  2.680000 3.525000 2.810000 ;
      RECT 3.705000  2.680000 4.035000 3.245000 ;
      RECT 3.755000  0.255000 3.985000 0.995000 ;
      RECT 4.155000  0.265000 7.535000 0.455000 ;
      RECT 4.155000  0.455000 4.485000 0.825000 ;
      RECT 4.585000  2.610000 4.915000 3.245000 ;
      RECT 4.655000  0.625000 8.045000 0.795000 ;
      RECT 4.655000  0.795000 4.915000 0.995000 ;
      RECT 5.480000  2.610000 5.730000 3.245000 ;
      RECT 6.305000  2.675000 6.975000 3.245000 ;
      RECT 7.505000  2.675000 7.835000 3.245000 ;
      RECT 7.715000  0.365000 8.045000 0.625000 ;
      RECT 7.715000  0.795000 8.045000 0.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__o211ai_4
