* File: sky130_fd_sc_lp__o41ai_m.pxi.spice
* Created: Fri Aug 28 11:20:53 2020
* 
x_PM_SKY130_FD_SC_LP__O41AI_M%B1 N_B1_c_67_n N_B1_M1000_g N_B1_M1006_g
+ N_B1_c_69_n B1 B1 B1 N_B1_c_71_n N_B1_c_72_n PM_SKY130_FD_SC_LP__O41AI_M%B1
x_PM_SKY130_FD_SC_LP__O41AI_M%A4 N_A4_M1005_g N_A4_M1004_g N_A4_c_107_n
+ N_A4_c_108_n A4 A4 A4 N_A4_c_109_n N_A4_c_110_n PM_SKY130_FD_SC_LP__O41AI_M%A4
x_PM_SKY130_FD_SC_LP__O41AI_M%A3 N_A3_M1008_g N_A3_M1007_g N_A3_c_149_n
+ N_A3_c_150_n A3 A3 A3 N_A3_c_151_n N_A3_c_152_n PM_SKY130_FD_SC_LP__O41AI_M%A3
x_PM_SKY130_FD_SC_LP__O41AI_M%A2 N_A2_M1009_g N_A2_M1001_g A2 A2 A2 A2 A2
+ N_A2_c_188_n PM_SKY130_FD_SC_LP__O41AI_M%A2
x_PM_SKY130_FD_SC_LP__O41AI_M%A1 N_A1_M1003_g N_A1_M1002_g N_A1_c_224_n
+ N_A1_c_225_n A1 A1 A1 N_A1_c_227_n PM_SKY130_FD_SC_LP__O41AI_M%A1
x_PM_SKY130_FD_SC_LP__O41AI_M%VPWR N_VPWR_M1000_s N_VPWR_M1003_d N_VPWR_c_251_n
+ N_VPWR_c_252_n N_VPWR_c_253_n N_VPWR_c_254_n N_VPWR_c_255_n N_VPWR_c_256_n
+ N_VPWR_c_257_n VPWR N_VPWR_c_250_n PM_SKY130_FD_SC_LP__O41AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O41AI_M%Y N_Y_M1006_s N_Y_M1000_d N_Y_c_276_n N_Y_c_277_n
+ Y Y Y Y N_Y_c_279_n N_Y_c_280_n PM_SKY130_FD_SC_LP__O41AI_M%Y
x_PM_SKY130_FD_SC_LP__O41AI_M%A_175_47# N_A_175_47#_M1006_d N_A_175_47#_M1007_d
+ N_A_175_47#_M1002_d N_A_175_47#_c_310_n N_A_175_47#_c_305_n
+ N_A_175_47#_c_306_n N_A_175_47#_c_323_n N_A_175_47#_c_307_n
+ N_A_175_47#_c_308_n N_A_175_47#_c_309_n PM_SKY130_FD_SC_LP__O41AI_M%A_175_47#
x_PM_SKY130_FD_SC_LP__O41AI_M%VGND N_VGND_M1004_d N_VGND_M1009_d N_VGND_c_350_n
+ N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n N_VGND_c_354_n N_VGND_c_355_n
+ VGND N_VGND_c_356_n N_VGND_c_357_n PM_SKY130_FD_SC_LP__O41AI_M%VGND
cc_1 VNB N_B1_c_67_n 0.023068f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.238
cc_2 VNB N_B1_M1000_g 0.0137975f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.065
cc_3 VNB N_B1_c_69_n 0.0231921f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.435
cc_4 VNB B1 0.0029205f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB N_B1_c_71_n 0.0254706f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.93
cc_6 VNB N_B1_c_72_n 0.0207147f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.765
cc_7 VNB N_A4_M1004_g 0.0312673f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.765
cc_8 VNB N_A4_c_107_n 0.0239241f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_9 VNB N_A4_c_108_n 0.009614f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_10 VNB N_A4_c_109_n 0.0162095f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.765
cc_11 VNB N_A4_c_110_n 9.16675e-19 $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.555
cc_12 VNB N_A3_M1007_g 0.030509f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.765
cc_13 VNB N_A3_c_149_n 0.0208703f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_14 VNB N_A3_c_150_n 0.00771831f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_15 VNB N_A3_c_151_n 0.0151728f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.765
cc_16 VNB N_A3_c_152_n 0.00576325f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.555
cc_17 VNB N_A2_M1009_g 0.052075f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.435
cc_18 VNB N_A1_M1003_g 4.92816e-19 $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.435
cc_19 VNB N_A1_M1002_g 0.035285f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.765
cc_20 VNB N_A1_c_224_n 0.0249397f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=1.435
cc_21 VNB N_A1_c_225_n 0.0173121f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_22 VNB A1 0.0446085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_227_n 0.0191428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_250_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_276_n 0.00460268f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.765
cc_26 VNB N_Y_c_277_n 0.00529045f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.445
cc_27 VNB Y 0.0486309f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_28 VNB N_Y_c_279_n 0.00172504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_280_n 0.0138247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_175_47#_c_305_n 0.0131606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_175_47#_c_306_n 0.00578023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_175_47#_c_307_n 0.0162284f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.765
cc_33 VNB N_A_175_47#_c_308_n 4.08405e-19 $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.925
cc_34 VNB N_A_175_47#_c_309_n 0.0056261f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.295
cc_35 VNB N_VGND_c_350_n 0.00228545f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.445
cc_36 VNB N_VGND_c_351_n 4.17679e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_37 VNB N_VGND_c_352_n 0.0377193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_353_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.93
cc_39 VNB N_VGND_c_354_n 0.015936f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.93
cc_40 VNB N_VGND_c_355_n 0.00436274f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.765
cc_41 VNB N_VGND_c_356_n 0.0217632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_357_n 0.200948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_B1_M1000_g 0.0303416f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.065
cc_44 VPB N_A4_M1005_g 0.0207519f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.435
cc_45 VPB N_A4_c_108_n 0.00878886f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_46 VPB N_A4_c_110_n 0.00118194f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.555
cc_47 VPB N_A3_M1008_g 0.0193566f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.435
cc_48 VPB N_A3_c_150_n 0.00819179f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_49 VPB N_A3_c_152_n 0.0030652f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=0.555
cc_50 VPB N_A2_M1009_g 0.0179465f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.435
cc_51 VPB A2 0.0845967f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=0.93
cc_52 VPB N_A2_c_188_n 0.0798651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A1_M1003_g 0.0249905f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=1.435
cc_54 VPB A1 0.0186865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_251_n 0.0133258f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.765
cc_56 VPB N_VPWR_c_252_n 0.0482075f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.445
cc_57 VPB N_VPWR_c_253_n 0.0501425f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_58 VPB N_VPWR_c_254_n 0.0106904f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_255_n 0.0112126f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.93
cc_60 VPB N_VPWR_c_256_n 0.0610587f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=0.93
cc_61 VPB N_VPWR_c_257_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=0.765
cc_62 VPB N_VPWR_c_250_n 0.0878874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_Y_c_276_n 0.00214315f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.765
cc_64 VPB N_Y_c_277_n 0.00283986f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=0.445
cc_65 VPB N_Y_c_279_n 0.00984303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 B1 N_A4_M1004_g 0.00120635f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_67 N_B1_c_72_n N_A4_M1004_g 0.0218998f $X=0.677 $Y=0.765 $X2=0 $Y2=0
cc_68 N_B1_M1000_g N_A4_c_107_n 0.0185247f $X=0.555 $Y=2.065 $X2=0 $Y2=0
cc_69 N_B1_c_69_n N_A4_c_107_n 0.0128623f $X=0.677 $Y=1.435 $X2=0 $Y2=0
cc_70 N_B1_c_67_n N_A4_c_109_n 0.0128623f $X=0.677 $Y=1.238 $X2=0 $Y2=0
cc_71 B1 N_A4_c_109_n 0.00131255f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_72 N_B1_c_67_n N_A4_c_110_n 0.00147929f $X=0.677 $Y=1.238 $X2=0 $Y2=0
cc_73 N_B1_M1000_g N_A4_c_110_n 0.00120031f $X=0.555 $Y=2.065 $X2=0 $Y2=0
cc_74 B1 N_A4_c_110_n 0.0175641f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_75 N_B1_M1000_g A2 0.00102925f $X=0.555 $Y=2.065 $X2=0 $Y2=0
cc_76 N_B1_M1000_g N_VPWR_c_252_n 0.00368657f $X=0.555 $Y=2.065 $X2=0 $Y2=0
cc_77 B1 N_Y_M1006_s 0.00279625f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_78 N_B1_M1000_g N_Y_c_276_n 0.0156536f $X=0.555 $Y=2.065 $X2=0 $Y2=0
cc_79 N_B1_c_69_n N_Y_c_276_n 0.00456165f $X=0.677 $Y=1.435 $X2=0 $Y2=0
cc_80 B1 N_Y_c_276_n 0.0147925f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_81 N_B1_M1000_g N_Y_c_277_n 0.016787f $X=0.555 $Y=2.065 $X2=0 $Y2=0
cc_82 B1 Y 0.0399752f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_83 N_B1_c_71_n Y 0.0230652f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_84 N_B1_c_72_n Y 8.79971e-19 $X=0.677 $Y=0.765 $X2=0 $Y2=0
cc_85 B1 N_Y_c_280_n 0.00907033f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_86 N_B1_c_72_n N_Y_c_280_n 0.00585812f $X=0.677 $Y=0.765 $X2=0 $Y2=0
cc_87 B1 N_A_175_47#_c_310_n 0.0131321f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_88 N_B1_c_72_n N_A_175_47#_c_310_n 0.0013917f $X=0.677 $Y=0.765 $X2=0 $Y2=0
cc_89 B1 N_A_175_47#_c_306_n 0.0131547f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_90 N_B1_c_72_n N_A_175_47#_c_306_n 0.00143851f $X=0.677 $Y=0.765 $X2=0 $Y2=0
cc_91 N_B1_c_72_n N_VGND_c_350_n 0.00144595f $X=0.677 $Y=0.765 $X2=0 $Y2=0
cc_92 B1 N_VGND_c_352_n 0.00426263f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_93 N_B1_c_71_n N_VGND_c_352_n 0.00316469f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_94 N_B1_c_72_n N_VGND_c_352_n 0.0048701f $X=0.677 $Y=0.765 $X2=0 $Y2=0
cc_95 B1 N_VGND_c_357_n 0.00568396f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_96 N_B1_c_71_n N_VGND_c_357_n 0.0039016f $X=0.71 $Y=0.93 $X2=0 $Y2=0
cc_97 N_B1_c_72_n N_VGND_c_357_n 0.00974176f $X=0.677 $Y=0.765 $X2=0 $Y2=0
cc_98 N_A4_M1005_g N_A3_M1008_g 0.0221566f $X=1.16 $Y=2.065 $X2=0 $Y2=0
cc_99 N_A4_c_110_n N_A3_M1008_g 0.00151917f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_100 N_A4_M1004_g N_A3_M1007_g 0.0238137f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A4_c_107_n N_A3_c_149_n 0.0139409f $X=1.25 $Y=1.53 $X2=0 $Y2=0
cc_102 N_A4_c_108_n N_A3_c_150_n 0.0139409f $X=1.25 $Y=1.695 $X2=0 $Y2=0
cc_103 N_A4_c_109_n N_A3_c_151_n 0.0139409f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_104 N_A4_c_110_n N_A3_c_151_n 7.13759e-19 $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_105 N_A4_M1005_g N_A3_c_152_n 6.96255e-19 $X=1.16 $Y=2.065 $X2=0 $Y2=0
cc_106 N_A4_c_109_n N_A3_c_152_n 0.00439653f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_107 N_A4_c_110_n N_A3_c_152_n 0.0537724f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_108 N_A4_M1005_g A2 0.0107821f $X=1.16 $Y=2.065 $X2=0 $Y2=0
cc_109 N_A4_c_108_n A2 0.00275793f $X=1.25 $Y=1.695 $X2=0 $Y2=0
cc_110 N_A4_c_110_n A2 0.014627f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_111 N_A4_c_108_n N_Y_c_276_n 0.004039f $X=1.25 $Y=1.695 $X2=0 $Y2=0
cc_112 N_A4_c_110_n N_Y_c_276_n 0.0356712f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_113 N_A4_c_110_n A_247_371# 0.00327996f $X=1.25 $Y=1.19 $X2=-0.19 $Y2=-0.245
cc_114 N_A4_M1004_g N_A_175_47#_c_310_n 2.06449e-19 $X=1.285 $Y=0.445 $X2=0
+ $Y2=0
cc_115 N_A4_M1004_g N_A_175_47#_c_305_n 0.0127145f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A4_c_109_n N_A_175_47#_c_305_n 0.00258429f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_117 N_A4_c_110_n N_A_175_47#_c_305_n 0.0126404f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_118 N_A4_c_109_n N_A_175_47#_c_306_n 0.00169678f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_119 N_A4_c_110_n N_A_175_47#_c_306_n 0.00311656f $X=1.25 $Y=1.19 $X2=0 $Y2=0
cc_120 N_A4_M1004_g N_VGND_c_350_n 0.00877283f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_121 N_A4_M1004_g N_VGND_c_352_n 0.0035715f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A4_M1004_g N_VGND_c_357_n 0.00441734f $X=1.285 $Y=0.445 $X2=0 $Y2=0
cc_123 N_A3_M1008_g N_A2_M1009_g 0.0212597f $X=1.7 $Y=2.065 $X2=0 $Y2=0
cc_124 N_A3_M1007_g N_A2_M1009_g 0.0275898f $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A3_c_151_n N_A2_M1009_g 0.0414616f $X=1.79 $Y=1.19 $X2=0 $Y2=0
cc_126 N_A3_c_152_n N_A2_M1009_g 0.00861447f $X=1.79 $Y=1.19 $X2=0 $Y2=0
cc_127 N_A3_M1008_g A2 0.00959258f $X=1.7 $Y=2.065 $X2=0 $Y2=0
cc_128 N_A3_c_150_n A2 0.00275425f $X=1.79 $Y=1.695 $X2=0 $Y2=0
cc_129 N_A3_c_152_n A2 0.0181365f $X=1.79 $Y=1.19 $X2=0 $Y2=0
cc_130 N_A3_c_151_n A1 0.00467428f $X=1.79 $Y=1.19 $X2=0 $Y2=0
cc_131 N_A3_c_152_n A1 0.0513127f $X=1.79 $Y=1.19 $X2=0 $Y2=0
cc_132 N_A3_c_152_n A_355_371# 0.00408785f $X=1.79 $Y=1.19 $X2=-0.19 $Y2=-0.245
cc_133 N_A3_M1007_g N_A_175_47#_c_305_n 0.012846f $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A3_c_151_n N_A_175_47#_c_305_n 0.00213861f $X=1.79 $Y=1.19 $X2=0 $Y2=0
cc_135 N_A3_c_152_n N_A_175_47#_c_305_n 0.0200234f $X=1.79 $Y=1.19 $X2=0 $Y2=0
cc_136 N_A3_M1007_g N_A_175_47#_c_323_n 2.1266e-19 $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A3_c_151_n N_A_175_47#_c_309_n 0.00157619f $X=1.79 $Y=1.19 $X2=0 $Y2=0
cc_138 N_A3_M1007_g N_VGND_c_350_n 0.00455727f $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A3_M1007_g N_VGND_c_351_n 7.49917e-19 $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A3_M1007_g N_VGND_c_354_n 0.00429465f $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A3_M1007_g N_VGND_c_357_n 0.00630109f $X=1.81 $Y=0.445 $X2=0 $Y2=0
cc_142 A2 N_A1_M1003_g 0.0106299f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_143 N_A2_M1009_g N_A1_M1002_g 0.0225036f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A2_M1009_g A1 0.0256016f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_145 A2 A1 0.0206341f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_146 N_A2_c_188_n A1 4.77605e-19 $X=2.15 $Y=2.6 $X2=0 $Y2=0
cc_147 N_A2_M1009_g N_A1_c_227_n 0.0912461f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_148 A2 N_VPWR_c_252_n 0.0515442f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_149 N_A2_M1009_g N_VPWR_c_253_n 0.0018945f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_150 A2 N_VPWR_c_253_n 0.0570159f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_151 N_A2_c_188_n N_VPWR_c_253_n 0.00175279f $X=2.15 $Y=2.6 $X2=0 $Y2=0
cc_152 N_A2_M1009_g N_VPWR_c_254_n 0.00104116f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_153 A2 N_VPWR_c_254_n 0.00405123f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_154 A2 N_VPWR_c_256_n 0.112362f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_155 N_A2_c_188_n N_VPWR_c_256_n 0.00643118f $X=2.15 $Y=2.6 $X2=0 $Y2=0
cc_156 A2 N_VPWR_c_250_n 0.0776942f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_157 N_A2_c_188_n N_VPWR_c_250_n 0.00853149f $X=2.15 $Y=2.6 $X2=0 $Y2=0
cc_158 A2 N_Y_c_276_n 0.0207504f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_159 N_A2_M1009_g N_A_175_47#_c_323_n 2.1266e-19 $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A2_M1009_g N_A_175_47#_c_307_n 0.0121373f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A2_M1009_g N_VGND_c_351_n 0.0064925f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A2_M1009_g N_VGND_c_354_n 0.00414412f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A2_M1009_g N_VGND_c_357_n 0.00486498f $X=2.24 $Y=0.445 $X2=0 $Y2=0
cc_164 N_A1_M1003_g N_VPWR_c_253_n 0.00490279f $X=2.6 $Y=2.065 $X2=0 $Y2=0
cc_165 N_A1_M1003_g N_VPWR_c_254_n 0.00439117f $X=2.6 $Y=2.065 $X2=0 $Y2=0
cc_166 N_A1_c_225_n N_VPWR_c_254_n 8.60181e-19 $X=2.69 $Y=1.645 $X2=0 $Y2=0
cc_167 A1 N_VPWR_c_254_n 0.0322212f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_168 N_A1_M1002_g N_A_175_47#_c_307_n 0.0133279f $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_169 A1 N_A_175_47#_c_307_n 0.0595141f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A1_c_227_n N_A_175_47#_c_307_n 0.00501445f $X=2.69 $Y=1.14 $X2=0 $Y2=0
cc_171 N_A1_M1002_g N_A_175_47#_c_308_n 3.52891e-19 $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_172 A1 N_A_175_47#_c_309_n 0.00418564f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_173 N_A1_M1002_g N_VGND_c_351_n 0.0112481f $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_174 N_A1_M1002_g N_VGND_c_356_n 0.0035715f $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_175 N_A1_M1002_g N_VGND_c_357_n 0.00540777f $X=2.69 $Y=0.445 $X2=0 $Y2=0
cc_176 N_VPWR_c_252_n N_Y_c_277_n 0.00777231f $X=0.34 $Y=2.13 $X2=0 $Y2=0
cc_177 N_VPWR_c_252_n N_Y_c_279_n 0.00784616f $X=0.34 $Y=2.13 $X2=0 $Y2=0
cc_178 N_Y_c_280_n N_A_175_47#_c_310_n 0.0039986f $X=0.36 $Y=0.43 $X2=0 $Y2=0
cc_179 N_Y_c_280_n N_VGND_c_352_n 0.0181759f $X=0.36 $Y=0.43 $X2=0 $Y2=0
cc_180 N_Y_M1006_s N_VGND_c_357_n 0.00711772f $X=0.235 $Y=0.235 $X2=0 $Y2=0
cc_181 N_Y_c_280_n N_VGND_c_357_n 0.011006f $X=0.36 $Y=0.43 $X2=0 $Y2=0
cc_182 N_A_175_47#_c_305_n N_VGND_c_350_n 0.0218189f $X=1.92 $Y=0.75 $X2=0 $Y2=0
cc_183 N_A_175_47#_c_307_n N_VGND_c_351_n 0.0193674f $X=2.82 $Y=0.75 $X2=0 $Y2=0
cc_184 N_A_175_47#_c_310_n N_VGND_c_352_n 0.00725952f $X=1.07 $Y=0.51 $X2=0
+ $Y2=0
cc_185 N_A_175_47#_c_305_n N_VGND_c_352_n 0.00283061f $X=1.92 $Y=0.75 $X2=0
+ $Y2=0
cc_186 N_A_175_47#_c_305_n N_VGND_c_354_n 0.00406811f $X=1.92 $Y=0.75 $X2=0
+ $Y2=0
cc_187 N_A_175_47#_c_323_n N_VGND_c_354_n 0.0081737f $X=2.025 $Y=0.51 $X2=0
+ $Y2=0
cc_188 N_A_175_47#_c_307_n N_VGND_c_354_n 0.002793f $X=2.82 $Y=0.75 $X2=0 $Y2=0
cc_189 N_A_175_47#_c_307_n N_VGND_c_356_n 0.00283061f $X=2.82 $Y=0.75 $X2=0
+ $Y2=0
cc_190 N_A_175_47#_c_308_n N_VGND_c_356_n 0.00812612f $X=2.905 $Y=0.51 $X2=0
+ $Y2=0
cc_191 N_A_175_47#_M1006_d N_VGND_c_357_n 0.0068193f $X=0.875 $Y=0.235 $X2=0
+ $Y2=0
cc_192 N_A_175_47#_M1007_d N_VGND_c_357_n 0.00257997f $X=1.885 $Y=0.235 $X2=0
+ $Y2=0
cc_193 N_A_175_47#_M1002_d N_VGND_c_357_n 0.00316012f $X=2.765 $Y=0.235 $X2=0
+ $Y2=0
cc_194 N_A_175_47#_c_310_n N_VGND_c_357_n 0.00615038f $X=1.07 $Y=0.51 $X2=0
+ $Y2=0
cc_195 N_A_175_47#_c_305_n N_VGND_c_357_n 0.0122453f $X=1.92 $Y=0.75 $X2=0 $Y2=0
cc_196 N_A_175_47#_c_323_n N_VGND_c_357_n 0.00762225f $X=2.025 $Y=0.51 $X2=0
+ $Y2=0
cc_197 N_A_175_47#_c_307_n N_VGND_c_357_n 0.0101677f $X=2.82 $Y=0.75 $X2=0 $Y2=0
cc_198 N_A_175_47#_c_308_n N_VGND_c_357_n 0.00688329f $X=2.905 $Y=0.51 $X2=0
+ $Y2=0
