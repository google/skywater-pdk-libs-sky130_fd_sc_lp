* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o221a_lp A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_482_419# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_114_47# a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_84_21# a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND A1 a_272_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_272_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_270_419# A2 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VPWR C1 a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 VPWR A1 a_270_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_272_47# B1 a_490_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_490_141# B2 a_272_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_490_141# C1 a_84_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_84_21# B2 a_482_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
