* File: sky130_fd_sc_lp__maj3_1.spice
* Created: Fri Aug 28 10:42:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__maj3_1.pex.spice"
.subckt sky130_fd_sc_lp__maj3_1  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 A_117_57# N_C_M1004_g N_A_30_57#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1197 PD=0.78 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g A_117_57# VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0756 PD=0.75 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.7 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1006 A_315_57# N_A_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0693 PD=0.66 PS=0.75 NRD=18.564 NRS=14.28 M=1 R=2.8 SA=75001.2 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_30_57#_M1007_d N_B_M1007_g A_315_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1001 A_479_57# N_B_M1001_g N_A_30_57#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_C_M1012_g A_479_57# VNB NSHORT L=0.15 W=0.42 AD=0.1176
+ AS=0.0441 PD=0.876667 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8 SA=75002.4
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1011 N_X_M1011_d N_A_30_57#_M1011_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.2352 PD=2.25 PS=1.75333 NRD=0 NRS=11.424 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 A_117_391# N_C_M1005_g N_A_30_57#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_117_391# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1013 A_275_391# N_A_M1013_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_30_57#_M1000_d N_B_M1000_g A_275_391# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.10855 AS=0.0441 PD=0.94 PS=0.63 NRD=53.9386 NRS=23.443 M=1 R=2.8
+ SA=75001.4 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1008 A_479_389# N_B_M1008_g N_A_30_57#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.10855 PD=0.63 PS=0.94 NRD=23.443 NRS=53.9386 M=1 R=2.8 SA=75002
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_C_M1009_g A_479_389# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.113925 AS=0.0441 PD=0.8875 PS=0.63 NRD=112.566 NRS=23.443 M=1 R=2.8
+ SA=75002.3 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1010 N_X_M1010_d N_A_30_57#_M1010_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.341775 PD=3.09 PS=2.6625 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__maj3_1.pxi.spice"
*
.ends
*
*
