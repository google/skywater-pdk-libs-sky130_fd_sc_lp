* File: sky130_fd_sc_lp__buflp_2.pxi.spice
* Created: Wed Sep  2 09:36:34 2020
* 
x_PM_SKY130_FD_SC_LP__BUFLP_2%A_98_21# N_A_98_21#_M1010_d N_A_98_21#_M1011_d
+ N_A_98_21#_M1003_g N_A_98_21#_M1001_g N_A_98_21#_c_60_n N_A_98_21#_M1005_g
+ N_A_98_21#_M1000_g N_A_98_21#_c_63_n N_A_98_21#_M1004_g N_A_98_21#_M1006_g
+ N_A_98_21#_c_66_n N_A_98_21#_M1009_g N_A_98_21#_M1007_g N_A_98_21#_c_69_n
+ N_A_98_21#_c_70_n N_A_98_21#_c_71_n N_A_98_21#_c_72_n N_A_98_21#_c_73_n
+ N_A_98_21#_c_143_p N_A_98_21#_c_74_n N_A_98_21#_c_75_n N_A_98_21#_c_76_n
+ N_A_98_21#_c_77_n PM_SKY130_FD_SC_LP__BUFLP_2%A_98_21#
x_PM_SKY130_FD_SC_LP__BUFLP_2%A N_A_M1002_g N_A_M1008_g N_A_M1011_g N_A_M1010_g
+ N_A_c_177_n N_A_c_178_n A A A A A N_A_c_180_n PM_SKY130_FD_SC_LP__BUFLP_2%A
x_PM_SKY130_FD_SC_LP__BUFLP_2%VPWR N_VPWR_M1001_s N_VPWR_M1009_s N_VPWR_c_221_n
+ N_VPWR_c_222_n N_VPWR_c_223_n VPWR N_VPWR_c_224_n N_VPWR_c_225_n
+ N_VPWR_c_220_n N_VPWR_c_227_n PM_SKY130_FD_SC_LP__BUFLP_2%VPWR
x_PM_SKY130_FD_SC_LP__BUFLP_2%A_128_367# N_A_128_367#_M1001_d
+ N_A_128_367#_M1004_d N_A_128_367#_c_262_n N_A_128_367#_c_260_n
+ N_A_128_367#_c_266_n N_A_128_367#_c_268_n N_A_128_367#_c_261_n
+ PM_SKY130_FD_SC_LP__BUFLP_2%A_128_367#
x_PM_SKY130_FD_SC_LP__BUFLP_2%X N_X_M1005_s N_X_M1000_s N_X_c_289_n N_X_c_286_n
+ X X X N_X_c_288_n X PM_SKY130_FD_SC_LP__BUFLP_2%X
x_PM_SKY130_FD_SC_LP__BUFLP_2%VGND N_VGND_M1003_d N_VGND_M1007_d N_VGND_c_313_n
+ N_VGND_c_314_n N_VGND_c_315_n VGND N_VGND_c_316_n N_VGND_c_317_n
+ N_VGND_c_318_n N_VGND_c_319_n PM_SKY130_FD_SC_LP__BUFLP_2%VGND
x_PM_SKY130_FD_SC_LP__BUFLP_2%A_128_47# N_A_128_47#_M1003_s N_A_128_47#_M1006_d
+ N_A_128_47#_c_361_n N_A_128_47#_c_359_n N_A_128_47#_c_360_n
+ PM_SKY130_FD_SC_LP__BUFLP_2%A_128_47#
cc_1 VNB N_A_98_21#_M1003_g 0.0278948f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.655
cc_2 VNB N_A_98_21#_M1001_g 0.0192195f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.465
cc_3 VNB N_A_98_21#_c_60_n 0.00927676f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.34
cc_4 VNB N_A_98_21#_M1005_g 0.0209547f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.655
cc_5 VNB N_A_98_21#_M1000_g 0.0116729f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.465
cc_6 VNB N_A_98_21#_c_63_n 0.0121512f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.34
cc_7 VNB N_A_98_21#_M1004_g 0.0111209f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.465
cc_8 VNB N_A_98_21#_M1006_g 0.0218169f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.655
cc_9 VNB N_A_98_21#_c_66_n 0.0412804f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.34
cc_10 VNB N_A_98_21#_M1009_g 0.00345975f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.465
cc_11 VNB N_A_98_21#_M1007_g 0.0220228f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.655
cc_12 VNB N_A_98_21#_c_69_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.34
cc_13 VNB N_A_98_21#_c_70_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.34
cc_14 VNB N_A_98_21#_c_71_n 0.00350226f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=1.34
cc_15 VNB N_A_98_21#_c_72_n 0.00323667f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=1.265
cc_16 VNB N_A_98_21#_c_73_n 0.00863674f $X=-0.19 $Y=-0.245 $X2=2.915 $Y2=0.8
cc_17 VNB N_A_98_21#_c_74_n 0.0177963f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.465
cc_18 VNB N_A_98_21#_c_75_n 0.0393057f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=2.03
cc_19 VNB N_A_98_21#_c_76_n 0.00371266f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=1.43
cc_20 VNB N_A_98_21#_c_77_n 0.00972716f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.8
cc_21 VNB N_A_M1002_g 0.0125743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_M1008_g 0.029574f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.265
cc_23 VNB N_A_M1010_g 0.0343787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_c_177_n 0.011631f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.655
cc_25 VNB N_A_c_178_n 0.00162136f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.655
cc_26 VNB A 2.81715e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_c_180_n 0.037314f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=1.34
cc_28 VNB N_VPWR_c_220_n 0.143779f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.655
cc_29 VNB N_X_c_286_n 0.00191926f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.465
cc_30 VNB X 0.00183274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_288_n 0.00450593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_313_n 0.0122131f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.265
cc_33 VNB N_VGND_c_314_n 0.0516846f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.655
cc_34 VNB N_VGND_c_315_n 0.00283848f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.465
cc_35 VNB N_VGND_c_316_n 0.0400467f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.265
cc_36 VNB N_VGND_c_317_n 0.0252107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_318_n 0.189363f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.34
cc_38 VNB N_VGND_c_319_n 0.00516132f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.265
cc_39 VNB N_A_128_47#_c_359_n 0.00846803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_128_47#_c_360_n 0.00470919f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.34
cc_41 VPB N_A_98_21#_M1001_g 0.0271666f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=2.465
cc_42 VPB N_A_98_21#_M1000_g 0.019028f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=2.465
cc_43 VPB N_A_98_21#_M1004_g 0.019028f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=2.465
cc_44 VPB N_A_98_21#_M1009_g 0.0237501f $X=-0.19 $Y=1.655 $X2=1.855 $Y2=2.465
cc_45 VPB N_A_98_21#_c_75_n 0.0414398f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=2.03
cc_46 VPB N_A_M1002_g 0.0236413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_c_178_n 0.0257988f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.655
cc_48 VPB A 0.0144345f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_221_n 0.0121872f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.265
cc_50 VPB N_VPWR_c_222_n 0.0676326f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.655
cc_51 VPB N_VPWR_c_223_n 0.0203377f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.34
cc_52 VPB N_VPWR_c_224_n 0.0369619f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=1.415
cc_53 VPB N_VPWR_c_225_n 0.0335683f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=1.265
cc_54 VPB N_VPWR_c_220_n 0.0617451f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=0.655
cc_55 VPB N_VPWR_c_227_n 0.00631788f $X=-0.19 $Y=1.655 $X2=1.855 $Y2=2.465
cc_56 VPB N_A_128_367#_c_260_n 0.00658097f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.655
cc_57 VPB N_A_128_367#_c_261_n 0.00658097f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.34
cc_58 N_A_98_21#_M1009_g N_A_M1002_g 0.0195085f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_59 N_A_98_21#_M1007_g N_A_M1008_g 0.0228336f $X=1.995 $Y=0.655 $X2=0 $Y2=0
cc_60 N_A_98_21#_c_72_n N_A_M1008_g 0.00374987f $X=2.2 $Y=1.265 $X2=0 $Y2=0
cc_61 N_A_98_21#_c_73_n N_A_M1008_g 0.0129847f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_62 N_A_98_21#_c_74_n N_A_M1008_g 0.00164334f $X=3.08 $Y=0.465 $X2=0 $Y2=0
cc_63 N_A_98_21#_c_73_n N_A_M1010_g 0.0116312f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_64 N_A_98_21#_c_74_n N_A_M1010_g 0.00927499f $X=3.08 $Y=0.465 $X2=0 $Y2=0
cc_65 N_A_98_21#_c_75_n N_A_M1010_g 0.0253462f $X=3.075 $Y=2.03 $X2=0 $Y2=0
cc_66 N_A_98_21#_c_77_n N_A_M1010_g 0.00506989f $X=3.08 $Y=0.8 $X2=0 $Y2=0
cc_67 N_A_98_21#_c_75_n N_A_c_178_n 0.0028928f $X=3.075 $Y=2.03 $X2=0 $Y2=0
cc_68 N_A_98_21#_c_66_n A 2.89866e-19 $X=1.78 $Y=1.34 $X2=0 $Y2=0
cc_69 N_A_98_21#_M1009_g A 0.00121877f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_98_21#_c_72_n A 0.014487f $X=2.2 $Y=1.265 $X2=0 $Y2=0
cc_71 N_A_98_21#_c_73_n A 0.0257739f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_72 N_A_98_21#_c_75_n A 0.0841047f $X=3.075 $Y=2.03 $X2=0 $Y2=0
cc_73 N_A_98_21#_c_76_n A 0.0245979f $X=2.2 $Y=1.43 $X2=0 $Y2=0
cc_74 N_A_98_21#_c_66_n N_A_c_180_n 0.0169314f $X=1.78 $Y=1.34 $X2=0 $Y2=0
cc_75 N_A_98_21#_M1007_g N_A_c_180_n 0.00657325f $X=1.995 $Y=0.655 $X2=0 $Y2=0
cc_76 N_A_98_21#_c_72_n N_A_c_180_n 0.00178471f $X=2.2 $Y=1.265 $X2=0 $Y2=0
cc_77 N_A_98_21#_c_73_n N_A_c_180_n 0.0016642f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_78 N_A_98_21#_c_76_n N_A_c_180_n 0.00233626f $X=2.2 $Y=1.43 $X2=0 $Y2=0
cc_79 N_A_98_21#_M1001_g N_VPWR_c_222_n 0.0294905f $X=0.565 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A_98_21#_c_66_n N_VPWR_c_223_n 0.00441317f $X=1.78 $Y=1.34 $X2=0 $Y2=0
cc_81 N_A_98_21#_M1009_g N_VPWR_c_223_n 0.018765f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A_98_21#_c_76_n N_VPWR_c_223_n 0.0220393f $X=2.2 $Y=1.43 $X2=0 $Y2=0
cc_83 N_A_98_21#_M1001_g N_VPWR_c_224_n 0.00547432f $X=0.565 $Y=2.465 $X2=0
+ $Y2=0
cc_84 N_A_98_21#_M1000_g N_VPWR_c_224_n 0.00357877f $X=0.995 $Y=2.465 $X2=0
+ $Y2=0
cc_85 N_A_98_21#_M1004_g N_VPWR_c_224_n 0.00357877f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_86 N_A_98_21#_M1009_g N_VPWR_c_224_n 0.00547432f $X=1.855 $Y=2.465 $X2=0
+ $Y2=0
cc_87 N_A_98_21#_M1001_g N_VPWR_c_220_n 0.0109207f $X=0.565 $Y=2.465 $X2=0 $Y2=0
cc_88 N_A_98_21#_M1000_g N_VPWR_c_220_n 0.0053512f $X=0.995 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_98_21#_M1004_g N_VPWR_c_220_n 0.0053512f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A_98_21#_M1009_g N_VPWR_c_220_n 0.0112356f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_91 N_A_98_21#_c_75_n N_VPWR_c_220_n 0.0104727f $X=3.075 $Y=2.03 $X2=0 $Y2=0
cc_92 N_A_98_21#_M1001_g N_A_128_367#_c_262_n 0.00202381f $X=0.565 $Y=2.465
+ $X2=0 $Y2=0
cc_93 N_A_98_21#_M1001_g N_A_128_367#_c_260_n 0.0143929f $X=0.565 $Y=2.465 $X2=0
+ $Y2=0
cc_94 N_A_98_21#_c_60_n N_A_128_367#_c_260_n 0.00322225f $X=0.92 $Y=1.34 $X2=0
+ $Y2=0
cc_95 N_A_98_21#_M1000_g N_A_128_367#_c_260_n 7.76258e-19 $X=0.995 $Y=2.465
+ $X2=0 $Y2=0
cc_96 N_A_98_21#_M1000_g N_A_128_367#_c_266_n 0.0115031f $X=0.995 $Y=2.465 $X2=0
+ $Y2=0
cc_97 N_A_98_21#_M1004_g N_A_128_367#_c_266_n 0.0115031f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_98 N_A_98_21#_M1009_g N_A_128_367#_c_268_n 0.00202381f $X=1.855 $Y=2.465
+ $X2=0 $Y2=0
cc_99 N_A_98_21#_M1004_g N_A_128_367#_c_261_n 7.76258e-19 $X=1.425 $Y=2.465
+ $X2=0 $Y2=0
cc_100 N_A_98_21#_c_66_n N_A_128_367#_c_261_n 0.00362155f $X=1.78 $Y=1.34 $X2=0
+ $Y2=0
cc_101 N_A_98_21#_M1009_g N_A_128_367#_c_261_n 0.0140864f $X=1.855 $Y=2.465
+ $X2=0 $Y2=0
cc_102 N_A_98_21#_M1006_g N_X_c_289_n 0.00441637f $X=1.495 $Y=0.655 $X2=0 $Y2=0
cc_103 N_A_98_21#_M1005_g N_X_c_286_n 0.00725442f $X=0.995 $Y=0.655 $X2=0 $Y2=0
cc_104 N_A_98_21#_M1006_g N_X_c_286_n 0.00355424f $X=1.495 $Y=0.655 $X2=0 $Y2=0
cc_105 N_A_98_21#_M1001_g X 0.00164123f $X=0.565 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_98_21#_M1000_g X 0.0217197f $X=0.995 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_98_21#_M1004_g X 0.0203594f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_98_21#_M1009_g X 0.0011872f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_98_21#_M1000_g N_X_c_288_n 0.00351276f $X=0.995 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A_98_21#_c_63_n N_X_c_288_n 0.016421f $X=1.35 $Y=1.34 $X2=0 $Y2=0
cc_111 N_A_98_21#_M1004_g N_X_c_288_n 0.00337539f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_98_21#_M1006_g N_X_c_288_n 0.00458509f $X=1.495 $Y=0.655 $X2=0 $Y2=0
cc_113 N_A_98_21#_c_66_n N_X_c_288_n 8.35463e-19 $X=1.78 $Y=1.34 $X2=0 $Y2=0
cc_114 N_A_98_21#_c_71_n N_X_c_288_n 0.00388491f $X=1.46 $Y=1.34 $X2=0 $Y2=0
cc_115 N_A_98_21#_c_76_n N_X_c_288_n 0.0112946f $X=2.2 $Y=1.43 $X2=0 $Y2=0
cc_116 N_A_98_21#_c_72_n N_VGND_M1007_d 0.0034086f $X=2.2 $Y=1.265 $X2=0 $Y2=0
cc_117 N_A_98_21#_c_73_n N_VGND_M1007_d 0.00164924f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_118 N_A_98_21#_c_143_p N_VGND_M1007_d 0.00283821f $X=2.285 $Y=0.8 $X2=0 $Y2=0
cc_119 N_A_98_21#_M1003_g N_VGND_c_314_n 0.0213563f $X=0.565 $Y=0.655 $X2=0
+ $Y2=0
cc_120 N_A_98_21#_M1007_g N_VGND_c_315_n 0.0047325f $X=1.995 $Y=0.655 $X2=0
+ $Y2=0
cc_121 N_A_98_21#_c_73_n N_VGND_c_315_n 0.00986593f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_122 N_A_98_21#_c_143_p N_VGND_c_315_n 0.0134161f $X=2.285 $Y=0.8 $X2=0 $Y2=0
cc_123 N_A_98_21#_c_74_n N_VGND_c_315_n 0.00952477f $X=3.08 $Y=0.465 $X2=0 $Y2=0
cc_124 N_A_98_21#_M1003_g N_VGND_c_316_n 0.00547432f $X=0.565 $Y=0.655 $X2=0
+ $Y2=0
cc_125 N_A_98_21#_M1005_g N_VGND_c_316_n 0.00357842f $X=0.995 $Y=0.655 $X2=0
+ $Y2=0
cc_126 N_A_98_21#_M1006_g N_VGND_c_316_n 0.00357877f $X=1.495 $Y=0.655 $X2=0
+ $Y2=0
cc_127 N_A_98_21#_M1007_g N_VGND_c_316_n 0.00547432f $X=1.995 $Y=0.655 $X2=0
+ $Y2=0
cc_128 N_A_98_21#_c_73_n N_VGND_c_317_n 0.00679134f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_129 N_A_98_21#_c_74_n N_VGND_c_317_n 0.0210428f $X=3.08 $Y=0.465 $X2=0 $Y2=0
cc_130 N_A_98_21#_M1010_d N_VGND_c_318_n 0.00232718f $X=2.94 $Y=0.235 $X2=0
+ $Y2=0
cc_131 N_A_98_21#_M1003_g N_VGND_c_318_n 0.0109207f $X=0.565 $Y=0.655 $X2=0
+ $Y2=0
cc_132 N_A_98_21#_M1005_g N_VGND_c_318_n 0.00553547f $X=0.995 $Y=0.655 $X2=0
+ $Y2=0
cc_133 N_A_98_21#_M1006_g N_VGND_c_318_n 0.0057905f $X=1.495 $Y=0.655 $X2=0
+ $Y2=0
cc_134 N_A_98_21#_M1007_g N_VGND_c_318_n 0.0102291f $X=1.995 $Y=0.655 $X2=0
+ $Y2=0
cc_135 N_A_98_21#_c_73_n N_VGND_c_318_n 0.0119613f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_136 N_A_98_21#_c_143_p N_VGND_c_318_n 7.32637e-19 $X=2.285 $Y=0.8 $X2=0 $Y2=0
cc_137 N_A_98_21#_c_74_n N_VGND_c_318_n 0.0126363f $X=3.08 $Y=0.465 $X2=0 $Y2=0
cc_138 N_A_98_21#_M1005_g N_A_128_47#_c_361_n 0.0109138f $X=0.995 $Y=0.655 $X2=0
+ $Y2=0
cc_139 N_A_98_21#_M1006_g N_A_128_47#_c_361_n 0.0143648f $X=1.495 $Y=0.655 $X2=0
+ $Y2=0
cc_140 N_A_98_21#_M1003_g N_A_128_47#_c_359_n 0.0120698f $X=0.565 $Y=0.655 $X2=0
+ $Y2=0
cc_141 N_A_98_21#_c_60_n N_A_128_47#_c_359_n 0.00411081f $X=0.92 $Y=1.34 $X2=0
+ $Y2=0
cc_142 N_A_98_21#_M1005_g N_A_128_47#_c_359_n 0.011994f $X=0.995 $Y=0.655 $X2=0
+ $Y2=0
cc_143 N_A_98_21#_M1006_g N_A_128_47#_c_359_n 7.01971e-19 $X=1.495 $Y=0.655
+ $X2=0 $Y2=0
cc_144 N_A_98_21#_M1006_g N_A_128_47#_c_360_n 0.00355554f $X=1.495 $Y=0.655
+ $X2=0 $Y2=0
cc_145 N_A_98_21#_c_66_n N_A_128_47#_c_360_n 0.00787729f $X=1.78 $Y=1.34 $X2=0
+ $Y2=0
cc_146 N_A_98_21#_M1007_g N_A_128_47#_c_360_n 0.0123732f $X=1.995 $Y=0.655 $X2=0
+ $Y2=0
cc_147 N_A_98_21#_c_72_n N_A_128_47#_c_360_n 0.00859455f $X=2.2 $Y=1.265 $X2=0
+ $Y2=0
cc_148 N_A_98_21#_c_76_n N_A_128_47#_c_360_n 0.00992925f $X=2.2 $Y=1.43 $X2=0
+ $Y2=0
cc_149 N_A_M1002_g N_VPWR_c_223_n 0.00759697f $X=2.47 $Y=2.205 $X2=0 $Y2=0
cc_150 A N_VPWR_c_223_n 0.0850744f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_151 N_A_M1002_g N_VPWR_c_225_n 0.00200596f $X=2.47 $Y=2.205 $X2=0 $Y2=0
cc_152 N_A_c_178_n N_VPWR_c_225_n 0.00295778f $X=2.862 $Y=1.775 $X2=0 $Y2=0
cc_153 A N_VPWR_c_225_n 0.0107254f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A_M1002_g N_VPWR_c_220_n 0.00228107f $X=2.47 $Y=2.205 $X2=0 $Y2=0
cc_155 N_A_c_178_n N_VPWR_c_220_n 0.00368913f $X=2.862 $Y=1.775 $X2=0 $Y2=0
cc_156 A N_VPWR_c_220_n 0.0114362f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A_M1008_g N_VGND_c_315_n 0.00957891f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_M1010_g N_VGND_c_315_n 0.00198482f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_M1008_g N_VGND_c_317_n 0.00392053f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_M1010_g N_VGND_c_317_n 0.00424868f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_M1008_g N_VGND_c_318_n 0.00444666f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_M1010_g N_VGND_c_318_n 0.00689221f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_M1008_g N_A_128_47#_c_360_n 8.89399e-19 $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_164 N_VPWR_c_220_n N_A_128_367#_M1001_d 0.00223562f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_165 N_VPWR_c_220_n N_A_128_367#_M1004_d 0.00223562f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_166 N_VPWR_c_224_n N_A_128_367#_c_262_n 0.0154369f $X=1.975 $Y=3.33 $X2=0
+ $Y2=0
cc_167 N_VPWR_c_220_n N_A_128_367#_c_262_n 0.00952129f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_168 N_VPWR_c_222_n N_A_128_367#_c_260_n 0.0399503f $X=0.28 $Y=1.98 $X2=0
+ $Y2=0
cc_169 N_VPWR_c_224_n N_A_128_367#_c_266_n 0.0368226f $X=1.975 $Y=3.33 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_220_n N_A_128_367#_c_266_n 0.024428f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_171 N_VPWR_c_224_n N_A_128_367#_c_268_n 0.0154369f $X=1.975 $Y=3.33 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_220_n N_A_128_367#_c_268_n 0.00952129f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_223_n N_A_128_367#_c_261_n 0.0399503f $X=2.14 $Y=1.98 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_220_n N_X_M1000_s 0.00225186f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_175 N_A_128_367#_c_266_n N_X_M1000_s 0.00332344f $X=1.555 $Y=2.99 $X2=0 $Y2=0
cc_176 N_A_128_367#_c_260_n X 0.033702f $X=0.78 $Y=1.98 $X2=0 $Y2=0
cc_177 N_A_128_367#_c_266_n X 0.0159805f $X=1.555 $Y=2.99 $X2=0 $Y2=0
cc_178 N_A_128_367#_c_261_n X 0.033702f $X=1.64 $Y=1.98 $X2=0 $Y2=0
cc_179 N_X_M1005_s N_VGND_c_318_n 0.00281482f $X=1.07 $Y=0.235 $X2=0 $Y2=0
cc_180 N_X_M1005_s N_A_128_47#_c_361_n 0.00472489f $X=1.07 $Y=0.235 $X2=0 $Y2=0
cc_181 N_X_c_289_n N_A_128_47#_c_361_n 0.0196319f $X=1.28 $Y=0.845 $X2=0 $Y2=0
cc_182 N_X_c_286_n N_A_128_47#_c_359_n 0.0195517f $X=1.28 $Y=1.095 $X2=0 $Y2=0
cc_183 N_X_c_289_n N_A_128_47#_c_360_n 0.0195142f $X=1.28 $Y=0.845 $X2=0 $Y2=0
cc_184 N_VGND_c_318_n N_A_128_47#_M1003_s 0.00223559f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_185 N_VGND_c_318_n N_A_128_47#_M1006_d 0.00280658f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_186 N_VGND_c_316_n N_A_128_47#_c_361_n 0.0374555f $X=2.115 $Y=0 $X2=0 $Y2=0
cc_187 N_VGND_c_318_n N_A_128_47#_c_361_n 0.0239316f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_188 N_VGND_c_314_n N_A_128_47#_c_359_n 0.025893f $X=0.28 $Y=0.38 $X2=0 $Y2=0
cc_189 N_VGND_c_316_n N_A_128_47#_c_359_n 0.01906f $X=2.115 $Y=0 $X2=0 $Y2=0
cc_190 N_VGND_c_318_n N_A_128_47#_c_359_n 0.0124545f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_191 N_VGND_c_316_n N_A_128_47#_c_360_n 0.0207136f $X=2.115 $Y=0 $X2=0 $Y2=0
cc_192 N_VGND_c_318_n N_A_128_47#_c_360_n 0.0126421f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_193 N_VGND_c_318_n A_516_47# 0.00268865f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
