* File: sky130_fd_sc_lp__buf_8.pxi.spice
* Created: Wed Sep  2 09:35:09 2020
* 
x_PM_SKY130_FD_SC_LP__BUF_8%A N_A_M1006_g N_A_M1000_g N_A_M1012_g N_A_M1007_g
+ N_A_M1021_g N_A_M1020_g N_A_c_126_p A A N_A_c_116_n N_A_c_117_n A N_A_c_118_n
+ PM_SKY130_FD_SC_LP__BUF_8%A
x_PM_SKY130_FD_SC_LP__BUF_8%A_27_47# N_A_27_47#_M1006_s N_A_27_47#_M1012_s
+ N_A_27_47#_M1000_s N_A_27_47#_M1007_s N_A_27_47#_M1002_g N_A_27_47#_M1001_g
+ N_A_27_47#_M1004_g N_A_27_47#_M1003_g N_A_27_47#_M1009_g N_A_27_47#_M1005_g
+ N_A_27_47#_M1010_g N_A_27_47#_M1008_g N_A_27_47#_M1011_g N_A_27_47#_M1013_g
+ N_A_27_47#_M1016_g N_A_27_47#_M1014_g N_A_27_47#_M1017_g N_A_27_47#_M1015_g
+ N_A_27_47#_M1019_g N_A_27_47#_M1018_g N_A_27_47#_c_188_n N_A_27_47#_c_204_n
+ N_A_27_47#_c_212_n N_A_27_47#_c_189_n N_A_27_47#_c_205_n N_A_27_47#_c_206_n
+ N_A_27_47#_c_343_p N_A_27_47#_c_257_p N_A_27_47#_c_190_n N_A_27_47#_c_207_n
+ N_A_27_47#_c_191_n N_A_27_47#_c_192_n N_A_27_47#_c_279_p N_A_27_47#_c_193_n
+ N_A_27_47#_c_209_n N_A_27_47#_c_194_n N_A_27_47#_c_195_n
+ PM_SKY130_FD_SC_LP__BUF_8%A_27_47#
x_PM_SKY130_FD_SC_LP__BUF_8%VPWR N_VPWR_M1000_d N_VPWR_M1020_d N_VPWR_M1003_s
+ N_VPWR_M1008_s N_VPWR_M1014_s N_VPWR_M1018_s N_VPWR_c_365_n N_VPWR_c_366_n
+ N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_371_n
+ N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_375_n N_VPWR_c_376_n
+ N_VPWR_c_377_n N_VPWR_c_378_n VPWR N_VPWR_c_379_n N_VPWR_c_380_n
+ N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_364_n PM_SKY130_FD_SC_LP__BUF_8%VPWR
x_PM_SKY130_FD_SC_LP__BUF_8%X N_X_M1002_s N_X_M1009_s N_X_M1011_s N_X_M1017_s
+ N_X_M1001_d N_X_M1005_d N_X_M1013_d N_X_M1015_d N_X_c_548_p N_X_c_523_n
+ N_X_c_458_n N_X_c_459_n N_X_c_448_n N_X_c_449_n N_X_c_527_n N_X_c_549_p
+ N_X_c_450_n N_X_c_460_n N_X_c_545_p N_X_c_531_n N_X_c_451_n N_X_c_461_n
+ N_X_c_550_p N_X_c_535_n N_X_c_452_n N_X_c_462_n N_X_c_463_n N_X_c_453_n
+ N_X_c_454_n N_X_c_464_n N_X_c_455_n N_X_c_465_n X X N_X_c_456_n N_X_c_466_n X
+ X PM_SKY130_FD_SC_LP__BUF_8%X
x_PM_SKY130_FD_SC_LP__BUF_8%VGND N_VGND_M1006_d N_VGND_M1021_d N_VGND_M1004_d
+ N_VGND_M1010_d N_VGND_M1016_d N_VGND_M1019_d N_VGND_c_559_n N_VGND_c_560_n
+ N_VGND_c_561_n N_VGND_c_562_n N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n
+ N_VGND_c_566_n N_VGND_c_567_n N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n
+ N_VGND_c_571_n N_VGND_c_572_n VGND N_VGND_c_573_n N_VGND_c_574_n
+ N_VGND_c_575_n N_VGND_c_576_n N_VGND_c_577_n PM_SKY130_FD_SC_LP__BUF_8%VGND
cc_1 VNB N_A_M1006_g 0.0295294f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A_M1000_g 7.24268e-19 $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_A_M1012_g 0.0222145f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_4 VNB N_A_M1007_g 4.57454e-19 $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_5 VNB N_A_M1021_g 0.0217865f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_6 VNB N_A_M1020_g 4.70211e-19 $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_7 VNB N_A_c_116_n 0.0686914f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.48
cc_8 VNB N_A_c_117_n 0.0231787f $X=-0.19 $Y=-0.245 $X2=0.683 $Y2=1.377
cc_9 VNB N_A_c_118_n 0.00137021f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.377
cc_10 VNB N_A_27_47#_M1002_g 0.0215666f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_11 VNB N_A_27_47#_M1001_g 4.20731e-19 $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.655
cc_12 VNB N_A_27_47#_M1004_g 0.0215225f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=2.465
cc_13 VNB N_A_27_47#_M1003_g 4.57127e-19 $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.48
cc_14 VNB N_A_27_47#_M1009_g 0.0215283f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_15 VNB N_A_27_47#_M1005_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.48
cc_16 VNB N_A_27_47#_M1010_g 0.0215283f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.48
cc_17 VNB N_A_27_47#_M1008_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_M1011_g 0.0215283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_M1013_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=0.744 $Y2=1.377
cc_20 VNB N_A_27_47#_M1016_g 0.0215283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_M1014_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_M1017_g 0.0215072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_M1015_g 4.57333e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_M1019_g 0.0267714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_M1018_g 4.92178e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_188_n 0.0207101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_189_n 0.00754163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_190_n 0.00157401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_191_n 0.00165721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_192_n 7.33997e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_193_n 0.00288935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_194_n 0.0010924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_c_195_n 0.155925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_364_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_448_n 0.00236792f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.48
cc_36 VNB N_X_c_449_n 0.0031671f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.48
cc_37 VNB N_X_c_450_n 0.00245068f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.377
cc_38 VNB N_X_c_451_n 0.0024047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_452_n 8.54366e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_453_n 0.00205183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_454_n 0.00209878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_455_n 0.00205183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_456_n 0.00992391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB X 0.0223168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_559_n 0.00461568f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=1.645
cc_46 VNB N_VGND_c_560_n 0.0019485f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.48
cc_47 VNB N_VGND_c_561_n 0.0039852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_562_n 0.00403119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_563_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.48
cc_50 VNB N_VGND_c_564_n 0.00400382f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.48
cc_51 VNB N_VGND_c_565_n 0.0119587f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.48
cc_52 VNB N_VGND_c_566_n 0.0288096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_567_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_568_n 0.00419476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_569_n 0.0154323f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.377
cc_56 VNB N_VGND_c_570_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_57 VNB N_VGND_c_571_n 0.0166607f $X=-0.19 $Y=-0.245 $X2=0.744 $Y2=1.377
cc_58 VNB N_VGND_c_572_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.377
cc_59 VNB N_VGND_c_573_n 0.0174638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_574_n 0.0166607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_575_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_576_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_577_n 0.268956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VPB N_A_M1000_g 0.0257233f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_65 VPB N_A_M1007_g 0.0190095f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_66 VPB N_A_M1020_g 0.0191965f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.465
cc_67 VPB N_A_27_47#_M1001_g 0.018828f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.655
cc_68 VPB N_A_27_47#_M1003_g 0.0190063f $X=-0.19 $Y=1.655 $X2=1.18 $Y2=1.48
cc_69 VPB N_A_27_47#_M1005_g 0.0190295f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.48
cc_70 VPB N_A_27_47#_M1008_g 0.0190295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_M1013_g 0.0190295f $X=-0.19 $Y=1.655 $X2=0.744 $Y2=1.377
cc_72 VPB N_A_27_47#_M1014_g 0.0190295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_M1015_g 0.0190083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_M1018_g 0.0233553f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_204_n 0.0406001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_205_n 0.00237632f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_206_n 0.0104412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_207_n 0.00157409f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_192_n 8.26908e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_209_n 0.00210048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_365_n 0.00461568f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=1.645
cc_82 VPB N_VPWR_c_366_n 0.00194769f $X=-0.19 $Y=1.655 $X2=1.18 $Y2=1.48
cc_83 VPB N_VPWR_c_367_n 0.00399712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_368_n 0.0039947f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.48
cc_85 VPB N_VPWR_c_369_n 0.0170141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_370_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_371_n 0.0125965f $X=-0.19 $Y=1.655 $X2=0.744 $Y2=1.377
cc_88 VPB N_VPWR_c_372_n 0.0044909f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=1.377
cc_89 VPB N_VPWR_c_373_n 0.0170141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_374_n 0.00416886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_375_n 0.0154359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_376_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_377_n 0.0172542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_378_n 0.00487897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_379_n 0.0176747f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_380_n 0.0170141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_381_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_382_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_364_n 0.0464292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_X_c_458_n 0.00233281f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.48
cc_101 VPB N_X_c_459_n 0.00262442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_X_c_460_n 0.00232361f $X=-0.19 $Y=1.655 $X2=0.744 $Y2=1.377
cc_103 VPB N_X_c_461_n 0.00240637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_X_c_462_n 8.4517e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_X_c_463_n 0.00219438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_X_c_464_n 0.00210048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_X_c_465_n 0.00210048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_X_c_466_n 0.0102459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB X 0.00463472f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 N_A_M1021_g N_A_27_47#_M1002_g 0.0208815f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_111 N_A_M1020_g N_A_27_47#_M1001_g 0.0208815f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_M1006_g N_A_27_47#_c_212_n 0.00994158f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_113 N_A_M1012_g N_A_27_47#_c_212_n 0.0107228f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_114 N_A_c_126_p N_A_27_47#_c_212_n 0.00376606f $X=1.18 $Y=1.48 $X2=0 $Y2=0
cc_115 N_A_c_116_n N_A_27_47#_c_212_n 5.18639e-19 $X=1.335 $Y=1.48 $X2=0 $Y2=0
cc_116 N_A_c_117_n N_A_27_47#_c_212_n 0.0328506f $X=0.683 $Y=1.377 $X2=0 $Y2=0
cc_117 N_A_c_116_n N_A_27_47#_c_189_n 2.03585e-19 $X=1.335 $Y=1.48 $X2=0 $Y2=0
cc_118 N_A_c_117_n N_A_27_47#_c_189_n 0.0239351f $X=0.683 $Y=1.377 $X2=0 $Y2=0
cc_119 N_A_M1000_g N_A_27_47#_c_205_n 0.0160357f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A_M1007_g N_A_27_47#_c_205_n 0.0149289f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_c_116_n N_A_27_47#_c_205_n 0.00268009f $X=1.335 $Y=1.48 $X2=0 $Y2=0
cc_122 N_A_c_117_n N_A_27_47#_c_205_n 0.0441902f $X=0.683 $Y=1.377 $X2=0 $Y2=0
cc_123 N_A_c_116_n N_A_27_47#_c_206_n 0.00139491f $X=1.335 $Y=1.48 $X2=0 $Y2=0
cc_124 N_A_c_117_n N_A_27_47#_c_206_n 0.026203f $X=0.683 $Y=1.377 $X2=0 $Y2=0
cc_125 N_A_M1021_g N_A_27_47#_c_190_n 0.0152177f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_126 N_A_c_126_p N_A_27_47#_c_190_n 0.00649467f $X=1.18 $Y=1.48 $X2=0 $Y2=0
cc_127 N_A_M1020_g N_A_27_47#_c_207_n 0.0156007f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_c_126_p N_A_27_47#_c_207_n 0.00652308f $X=1.18 $Y=1.48 $X2=0 $Y2=0
cc_129 N_A_M1021_g N_A_27_47#_c_191_n 0.0021261f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_130 N_A_c_126_p N_A_27_47#_c_191_n 6.52292e-19 $X=1.18 $Y=1.48 $X2=0 $Y2=0
cc_131 N_A_c_118_n N_A_27_47#_c_191_n 0.00480537f $X=0.88 $Y=1.377 $X2=0 $Y2=0
cc_132 N_A_c_116_n N_A_27_47#_c_192_n 0.00383378f $X=1.335 $Y=1.48 $X2=0 $Y2=0
cc_133 N_A_M1012_g N_A_27_47#_c_193_n 0.0051423f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_134 N_A_c_126_p N_A_27_47#_c_193_n 0.0176802f $X=1.18 $Y=1.48 $X2=0 $Y2=0
cc_135 N_A_c_116_n N_A_27_47#_c_193_n 0.00253619f $X=1.335 $Y=1.48 $X2=0 $Y2=0
cc_136 N_A_c_118_n N_A_27_47#_c_193_n 0.00301828f $X=0.88 $Y=1.377 $X2=0 $Y2=0
cc_137 N_A_c_126_p N_A_27_47#_c_209_n 0.021133f $X=1.18 $Y=1.48 $X2=0 $Y2=0
cc_138 N_A_c_116_n N_A_27_47#_c_209_n 0.00253619f $X=1.335 $Y=1.48 $X2=0 $Y2=0
cc_139 N_A_c_126_p N_A_27_47#_c_194_n 0.0152784f $X=1.18 $Y=1.48 $X2=0 $Y2=0
cc_140 N_A_c_116_n N_A_27_47#_c_194_n 0.00162571f $X=1.335 $Y=1.48 $X2=0 $Y2=0
cc_141 N_A_c_116_n N_A_27_47#_c_195_n 0.0208815f $X=1.335 $Y=1.48 $X2=0 $Y2=0
cc_142 N_A_M1000_g N_VPWR_c_365_n 0.00309734f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_M1007_g N_VPWR_c_365_n 0.0016342f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_M1020_g N_VPWR_c_366_n 0.00164187f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_M1007_g N_VPWR_c_373_n 0.00585385f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_M1020_g N_VPWR_c_373_n 0.00585385f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_M1000_g N_VPWR_c_379_n 0.00585385f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_M1000_g N_VPWR_c_364_n 0.0116345f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_M1007_g N_VPWR_c_364_n 0.0106302f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_M1020_g N_VPWR_c_364_n 0.0106555f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_M1006_g N_VGND_c_559_n 0.00343894f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_152 N_A_M1012_g N_VGND_c_559_n 0.00197579f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_153 N_A_M1021_g N_VGND_c_560_n 0.00164187f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_154 N_A_M1012_g N_VGND_c_567_n 0.00585385f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_155 N_A_M1021_g N_VGND_c_567_n 0.00585385f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_156 N_A_M1006_g N_VGND_c_573_n 0.00585385f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_157 N_A_M1006_g N_VGND_c_577_n 0.00729459f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_158 N_A_M1012_g N_VGND_c_577_n 0.00629024f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_159 N_A_M1021_g N_VGND_c_577_n 0.0106555f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_205_n N_VPWR_M1000_d 0.00176773f $X=0.99 $Y=1.835 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_27_47#_c_207_n N_VPWR_M1020_d 0.00180215f $X=1.525 $Y=1.835 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_205_n N_VPWR_c_365_n 0.0135577f $X=0.99 $Y=1.835 $X2=0 $Y2=0
cc_163 N_A_27_47#_M1001_g N_VPWR_c_366_n 0.0125052f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_M1003_g N_VPWR_c_366_n 9.28559e-19 $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_207_n N_VPWR_c_366_n 0.014734f $X=1.525 $Y=1.835 $X2=0 $Y2=0
cc_166 N_A_27_47#_M1003_g N_VPWR_c_367_n 0.00162836f $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_M1005_g N_VPWR_c_367_n 0.00162593f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_M1008_g N_VPWR_c_368_n 0.00162328f $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_M1013_g N_VPWR_c_368_n 0.00163155f $X=3.485 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_M1013_g N_VPWR_c_369_n 0.00585385f $X=3.485 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_M1014_g N_VPWR_c_369_n 0.00585385f $X=3.915 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_M1014_g N_VPWR_c_370_n 0.0016342f $X=3.915 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_M1015_g N_VPWR_c_370_n 0.0016342f $X=4.345 $Y=2.465 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_M1018_g N_VPWR_c_372_n 0.00340667f $X=4.775 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_257_p N_VPWR_c_373_n 0.00931637f $X=1.12 $Y=2.075 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1001_g N_VPWR_c_375_n 0.00564095f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_M1003_g N_VPWR_c_375_n 0.00585385f $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_M1005_g N_VPWR_c_377_n 0.00585385f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1008_g N_VPWR_c_377_n 0.00585385f $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_204_n N_VPWR_c_379_n 0.011826f $X=0.26 $Y=2.075 $X2=0 $Y2=0
cc_181 N_A_27_47#_M1015_g N_VPWR_c_380_n 0.00585385f $X=4.345 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_M1018_g N_VPWR_c_380_n 0.00585385f $X=4.775 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_M1000_s N_VPWR_c_364_n 0.00262668f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_M1007_s N_VPWR_c_364_n 0.00310272f $X=0.98 $Y=1.835 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_M1001_g N_VPWR_c_364_n 0.00959071f $X=1.765 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_M1003_g N_VPWR_c_364_n 0.0106165f $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_M1005_g N_VPWR_c_364_n 0.0106439f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_M1008_g N_VPWR_c_364_n 0.0106439f $X=3.055 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_M1013_g N_VPWR_c_364_n 0.0106302f $X=3.485 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_M1014_g N_VPWR_c_364_n 0.0106302f $X=3.915 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1015_g N_VPWR_c_364_n 0.0106302f $X=4.345 $Y=2.465 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1018_g N_VPWR_c_364_n 0.01159f $X=4.775 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_204_n N_VPWR_c_364_n 0.0108215f $X=0.26 $Y=2.075 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_257_p N_VPWR_c_364_n 0.0095288f $X=1.12 $Y=2.075 $X2=0 $Y2=0
cc_195 N_A_27_47#_M1003_g N_X_c_458_n 0.0146201f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A_27_47#_M1005_g N_X_c_458_n 0.0148796f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_279_p N_X_c_458_n 0.0420862f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_195_n N_X_c_458_n 0.00243878f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_199 N_A_27_47#_M1001_g N_X_c_459_n 9.70485e-19 $X=1.765 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_207_n N_X_c_459_n 0.0117851f $X=1.525 $Y=1.835 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_279_p N_X_c_459_n 0.0194383f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_195_n N_X_c_459_n 0.00253619f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_203 N_A_27_47#_M1004_g N_X_c_448_n 0.0150929f $X=2.195 $Y=0.655 $X2=0 $Y2=0
cc_204 N_A_27_47#_M1009_g N_X_c_448_n 0.0154538f $X=2.625 $Y=0.655 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_279_p N_X_c_448_n 0.0420861f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_195_n N_X_c_448_n 0.00246815f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_207 N_A_27_47#_M1002_g N_X_c_449_n 0.00141838f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_190_n N_X_c_449_n 0.013645f $X=1.525 $Y=1.13 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_191_n N_X_c_449_n 7.72648e-19 $X=1.61 $Y=1.395 $X2=0 $Y2=0
cc_210 N_A_27_47#_c_279_p N_X_c_449_n 0.0198432f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_195_n N_X_c_449_n 0.00256759f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_212 N_A_27_47#_M1010_g N_X_c_450_n 0.0155031f $X=3.055 $Y=0.655 $X2=0 $Y2=0
cc_213 N_A_27_47#_M1011_g N_X_c_450_n 0.0155031f $X=3.485 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_279_p N_X_c_450_n 0.042447f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_215 N_A_27_47#_c_195_n N_X_c_450_n 0.00246815f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_216 N_A_27_47#_M1008_g N_X_c_460_n 0.0149289f $X=3.055 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_27_47#_M1013_g N_X_c_460_n 0.0149289f $X=3.485 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_279_p N_X_c_460_n 0.0417254f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_195_n N_X_c_460_n 0.00243878f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_220 N_A_27_47#_M1016_g N_X_c_451_n 0.0155031f $X=3.915 $Y=0.655 $X2=0 $Y2=0
cc_221 N_A_27_47#_M1017_g N_X_c_451_n 0.0155031f $X=4.345 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_279_p N_X_c_451_n 0.0420861f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_195_n N_X_c_451_n 0.00246815f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_224 N_A_27_47#_M1014_g N_X_c_461_n 0.0149289f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A_27_47#_M1015_g N_X_c_461_n 0.0149289f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_279_p N_X_c_461_n 0.0420862f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_195_n N_X_c_461_n 0.00243878f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_228 N_A_27_47#_M1019_g N_X_c_452_n 0.0182536f $X=4.775 $Y=0.655 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_279_p N_X_c_452_n 0.00377973f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_230 N_A_27_47#_M1018_g N_X_c_462_n 0.0176794f $X=4.775 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_279_p N_X_c_462_n 0.00341888f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_279_p N_X_c_463_n 0.0218684f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_195_n N_X_c_463_n 0.00253619f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_279_p N_X_c_453_n 0.0206533f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_195_n N_X_c_453_n 0.00256759f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_279_p N_X_c_454_n 0.0210583f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_195_n N_X_c_454_n 0.00256759f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_279_p N_X_c_464_n 0.0210584f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_195_n N_X_c_464_n 0.00253619f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_279_p N_X_c_455_n 0.0206533f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_195_n N_X_c_455_n 0.00256759f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_279_p N_X_c_465_n 0.0210584f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_195_n N_X_c_465_n 0.00253619f $X=4.775 $Y=1.48 $X2=0 $Y2=0
cc_244 N_A_27_47#_M1019_g X 0.0205744f $X=4.775 $Y=0.655 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_279_p X 0.0147523f $X=4.575 $Y=1.48 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_212_n N_VGND_M1006_d 0.00332539f $X=0.99 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_247 N_A_27_47#_c_190_n N_VGND_M1021_d 0.00180108f $X=1.525 $Y=1.13 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_212_n N_VGND_c_559_n 0.0132096f $X=0.99 $Y=0.925 $X2=0 $Y2=0
cc_249 N_A_27_47#_M1002_g N_VGND_c_560_n 0.00901192f $X=1.765 $Y=0.655 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_M1004_g N_VGND_c_560_n 7.15732e-19 $X=2.195 $Y=0.655 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_190_n N_VGND_c_560_n 0.0147161f $X=1.525 $Y=1.13 $X2=0 $Y2=0
cc_252 N_A_27_47#_M1004_g N_VGND_c_561_n 0.00161359f $X=2.195 $Y=0.655 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_M1009_g N_VGND_c_561_n 0.00162736f $X=2.625 $Y=0.655 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_M1010_g N_VGND_c_562_n 0.00165192f $X=3.055 $Y=0.655 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_M1011_g N_VGND_c_562_n 0.0016368f $X=3.485 $Y=0.655 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_M1011_g N_VGND_c_563_n 0.00585385f $X=3.485 $Y=0.655 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1016_g N_VGND_c_563_n 0.00585385f $X=3.915 $Y=0.655 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1016_g N_VGND_c_564_n 0.0016342f $X=3.915 $Y=0.655 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1017_g N_VGND_c_564_n 0.00162736f $X=4.345 $Y=0.655 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1019_g N_VGND_c_566_n 0.00346837f $X=4.775 $Y=0.655 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_343_p N_VGND_c_567_n 0.0113494f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_262 N_A_27_47#_M1002_g N_VGND_c_569_n 0.00564095f $X=1.765 $Y=0.655 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1004_g N_VGND_c_569_n 0.00585385f $X=2.195 $Y=0.655 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_M1009_g N_VGND_c_571_n 0.00585385f $X=2.625 $Y=0.655 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_M1010_g N_VGND_c_571_n 0.00585385f $X=3.055 $Y=0.655 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_188_n N_VGND_c_573_n 0.0144694f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_267 N_A_27_47#_M1017_g N_VGND_c_574_n 0.00585385f $X=4.345 $Y=0.655 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_M1019_g N_VGND_c_574_n 0.00585385f $X=4.775 $Y=0.655 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_M1006_s N_VGND_c_577_n 0.00224546f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_M1012_s N_VGND_c_577_n 0.0027206f $X=0.98 $Y=0.235 $X2=0 $Y2=0
cc_271 N_A_27_47#_M1002_g N_VGND_c_577_n 0.00959071f $X=1.765 $Y=0.655 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1004_g N_VGND_c_577_n 0.0106302f $X=2.195 $Y=0.655 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1009_g N_VGND_c_577_n 0.0106302f $X=2.625 $Y=0.655 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_M1010_g N_VGND_c_577_n 0.0106165f $X=3.055 $Y=0.655 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1011_g N_VGND_c_577_n 0.0106302f $X=3.485 $Y=0.655 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1016_g N_VGND_c_577_n 0.0106302f $X=3.915 $Y=0.655 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_M1017_g N_VGND_c_577_n 0.0106302f $X=4.345 $Y=0.655 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_M1019_g N_VGND_c_577_n 0.0115763f $X=4.775 $Y=0.655 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_c_188_n N_VGND_c_577_n 0.0111175f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_212_n N_VGND_c_577_n 0.0103332f $X=0.99 $Y=0.925 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_343_p N_VGND_c_577_n 0.00978101f $X=1.12 $Y=0.47 $X2=0 $Y2=0
cc_282 N_VPWR_c_364_n N_X_M1001_d 0.00379183f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_283 N_VPWR_c_364_n N_X_M1005_d 0.00275817f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_284 N_VPWR_c_364_n N_X_M1013_d 0.00310272f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_285 N_VPWR_c_364_n N_X_M1015_d 0.00310272f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_286 N_VPWR_c_375_n N_X_c_523_n 0.008858f $X=2.275 $Y=3.33 $X2=0 $Y2=0
cc_287 N_VPWR_c_364_n N_X_c_523_n 0.00879013f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_288 N_VPWR_M1003_s N_X_c_458_n 0.00176773f $X=2.27 $Y=1.835 $X2=0 $Y2=0
cc_289 N_VPWR_c_367_n N_X_c_458_n 0.0135577f $X=2.41 $Y=2.26 $X2=0 $Y2=0
cc_290 N_VPWR_c_377_n N_X_c_527_n 0.00954555f $X=3.145 $Y=3.33 $X2=0 $Y2=0
cc_291 N_VPWR_c_364_n N_X_c_527_n 0.00989813f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_292 N_VPWR_M1008_s N_X_c_460_n 0.00176773f $X=3.13 $Y=1.835 $X2=0 $Y2=0
cc_293 N_VPWR_c_368_n N_X_c_460_n 0.0135577f $X=3.27 $Y=2.26 $X2=0 $Y2=0
cc_294 N_VPWR_c_369_n N_X_c_531_n 0.00931637f $X=4 $Y=3.33 $X2=0 $Y2=0
cc_295 N_VPWR_c_364_n N_X_c_531_n 0.0095288f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_296 N_VPWR_M1014_s N_X_c_461_n 0.00176773f $X=3.99 $Y=1.835 $X2=0 $Y2=0
cc_297 N_VPWR_c_370_n N_X_c_461_n 0.0135577f $X=4.13 $Y=2.26 $X2=0 $Y2=0
cc_298 N_VPWR_c_380_n N_X_c_535_n 0.00931637f $X=4.86 $Y=3.33 $X2=0 $Y2=0
cc_299 N_VPWR_c_364_n N_X_c_535_n 0.0095288f $X=5.04 $Y=3.33 $X2=0 $Y2=0
cc_300 N_VPWR_M1018_s N_X_c_466_n 0.00440878f $X=4.85 $Y=1.835 $X2=0 $Y2=0
cc_301 N_VPWR_c_372_n N_X_c_466_n 0.0165898f $X=4.99 $Y=2.26 $X2=0 $Y2=0
cc_302 N_X_c_448_n N_VGND_M1004_d 0.00176773f $X=2.71 $Y=1.135 $X2=0 $Y2=0
cc_303 N_X_c_450_n N_VGND_M1010_d 0.00176773f $X=3.57 $Y=1.135 $X2=0 $Y2=0
cc_304 N_X_c_451_n N_VGND_M1016_d 0.00176773f $X=4.43 $Y=1.135 $X2=0 $Y2=0
cc_305 N_X_c_456_n N_VGND_M1019_d 0.00266426f $X=5.05 $Y=1.225 $X2=0 $Y2=0
cc_306 N_X_c_448_n N_VGND_c_561_n 0.0135577f $X=2.71 $Y=1.135 $X2=0 $Y2=0
cc_307 N_X_c_450_n N_VGND_c_562_n 0.0135577f $X=3.57 $Y=1.135 $X2=0 $Y2=0
cc_308 N_X_c_545_p N_VGND_c_563_n 0.0113476f $X=3.7 $Y=0.47 $X2=0 $Y2=0
cc_309 N_X_c_451_n N_VGND_c_564_n 0.0135577f $X=4.43 $Y=1.135 $X2=0 $Y2=0
cc_310 N_X_c_456_n N_VGND_c_566_n 0.0220667f $X=5.05 $Y=1.225 $X2=0 $Y2=0
cc_311 N_X_c_548_p N_VGND_c_569_n 0.0109351f $X=1.98 $Y=0.47 $X2=0 $Y2=0
cc_312 N_X_c_549_p N_VGND_c_571_n 0.0112101f $X=2.84 $Y=0.47 $X2=0 $Y2=0
cc_313 N_X_c_550_p N_VGND_c_574_n 0.0112101f $X=4.56 $Y=0.47 $X2=0 $Y2=0
cc_314 N_X_M1002_s N_VGND_c_577_n 0.00356516f $X=1.84 $Y=0.235 $X2=0 $Y2=0
cc_315 N_X_M1009_s N_VGND_c_577_n 0.00321837f $X=2.7 $Y=0.235 $X2=0 $Y2=0
cc_316 N_X_M1011_s N_VGND_c_577_n 0.00304497f $X=3.56 $Y=0.235 $X2=0 $Y2=0
cc_317 N_X_M1017_s N_VGND_c_577_n 0.00321837f $X=4.42 $Y=0.235 $X2=0 $Y2=0
cc_318 N_X_c_548_p N_VGND_c_577_n 0.00920999f $X=1.98 $Y=0.47 $X2=0 $Y2=0
cc_319 N_X_c_549_p N_VGND_c_577_n 0.00958901f $X=2.84 $Y=0.47 $X2=0 $Y2=0
cc_320 N_X_c_545_p N_VGND_c_577_n 0.00977851f $X=3.7 $Y=0.47 $X2=0 $Y2=0
cc_321 N_X_c_550_p N_VGND_c_577_n 0.00958901f $X=4.56 $Y=0.47 $X2=0 $Y2=0
