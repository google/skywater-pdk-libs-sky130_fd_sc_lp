* NGSPICE file created from sky130_fd_sc_lp__o2111a_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o2111a_m A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_348_47# D1 a_80_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.1e+11p ps=1.84e+06u
M1001 VPWR a_80_21# X VPB phighvt w=420000u l=150000u
+  ad=4.746e+11p pd=4.78e+06u as=1.113e+11p ps=1.37e+06u
M1002 VGND A2 a_492_47# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.289e+11p ps=2.77e+06u
M1003 a_564_535# A2 a_80_21# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.352e+11p ps=2.8e+06u
M1004 VGND a_80_21# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VPWR A1 a_564_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_492_47# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_420_47# C1 a_348_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 VPWR C1 a_80_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_492_47# B1 a_420_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_80_21# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_80_21# D1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

