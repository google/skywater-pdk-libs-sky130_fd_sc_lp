* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux4_m A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 a_345_126# S0 a_273_463# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_273_126# A2 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=5.208e+11p ps=5.84e+06u
M1002 X a_1184_171# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=7.371e+11p ps=6.87e+06u
M1003 VGND A3 a_453_126# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 a_688_126# a_59_463# a_647_463# VPB phighvt w=420000u l=150000u
+  ad=3.423e+11p pd=3.31e+06u as=8.82e+10p ps=1.26e+06u
M1005 a_345_126# a_1118_37# a_1184_171# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1006 a_453_126# S0 a_345_126# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.751e+11p ps=2.99e+06u
M1007 VPWR A3 a_431_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1008 X a_1184_171# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1009 VGND A0 a_774_126# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 VPWR S1 a_1118_37# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 a_647_463# A1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1184_171# S1 a_688_126# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_431_463# a_59_463# a_345_126# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND S0 a_59_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1015 a_688_126# S0 a_616_126# VNB nshort w=420000u l=150000u
+  ad=3.423e+11p pd=3.31e+06u as=8.82e+10p ps=1.26e+06u
M1016 a_774_126# a_59_463# a_688_126# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_805_463# S0 a_688_126# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1018 a_1184_171# a_1118_37# a_688_126# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1019 VPWR A0 a_805_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_345_126# a_59_463# a_273_126# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_345_126# S1 a_1184_171# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_616_126# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR S0 a_59_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1024 a_273_463# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND S1 a_1118_37# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends
