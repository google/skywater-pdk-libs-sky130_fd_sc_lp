* File: sky130_fd_sc_lp__sdfxtp_1.pxi.spice
* Created: Wed Sep  2 10:36:32 2020
* 
x_PM_SKY130_FD_SC_LP__SDFXTP_1%A_78_123# N_A_78_123#_M1017_s N_A_78_123#_M1020_s
+ N_A_78_123#_c_219_n N_A_78_123#_M1010_g N_A_78_123#_M1011_g
+ N_A_78_123#_c_221_n N_A_78_123#_c_227_n N_A_78_123#_c_228_n
+ N_A_78_123#_c_222_n N_A_78_123#_c_230_n N_A_78_123#_c_231_n
+ N_A_78_123#_c_223_n N_A_78_123#_c_224_n N_A_78_123#_c_225_n
+ PM_SKY130_FD_SC_LP__SDFXTP_1%A_78_123#
x_PM_SKY130_FD_SC_LP__SDFXTP_1%D N_D_M1006_g N_D_M1028_g N_D_c_310_n N_D_c_315_n
+ D D D D D N_D_c_312_n PM_SKY130_FD_SC_LP__SDFXTP_1%D
x_PM_SKY130_FD_SC_LP__SDFXTP_1%SCE N_SCE_c_359_n N_SCE_M1017_g N_SCE_c_367_n
+ N_SCE_M1020_g N_SCE_c_361_n N_SCE_c_362_n N_SCE_c_368_n N_SCE_c_369_n
+ N_SCE_c_370_n N_SCE_M1023_g N_SCE_M1031_g SCE SCE N_SCE_c_365_n
+ PM_SKY130_FD_SC_LP__SDFXTP_1%SCE
x_PM_SKY130_FD_SC_LP__SDFXTP_1%SCD N_SCD_M1007_g N_SCD_M1016_g SCD SCD
+ N_SCD_c_429_n PM_SKY130_FD_SC_LP__SDFXTP_1%SCD
x_PM_SKY130_FD_SC_LP__SDFXTP_1%CLK N_CLK_M1009_g N_CLK_M1027_g CLK CLK CLK
+ N_CLK_c_478_n PM_SKY130_FD_SC_LP__SDFXTP_1%CLK
x_PM_SKY130_FD_SC_LP__SDFXTP_1%A_628_123# N_A_628_123#_M1009_d
+ N_A_628_123#_M1027_d N_A_628_123#_M1004_g N_A_628_123#_M1024_g
+ N_A_628_123#_M1018_g N_A_628_123#_M1029_g N_A_628_123#_M1008_g
+ N_A_628_123#_M1025_g N_A_628_123#_c_526_n N_A_628_123#_c_527_n
+ N_A_628_123#_c_528_n N_A_628_123#_c_529_n N_A_628_123#_c_530_n
+ N_A_628_123#_c_531_n N_A_628_123#_c_546_n N_A_628_123#_c_547_n
+ N_A_628_123#_c_548_n N_A_628_123#_c_532_n N_A_628_123#_c_533_n
+ N_A_628_123#_c_577_p N_A_628_123#_c_550_n N_A_628_123#_c_551_n
+ N_A_628_123#_c_534_n N_A_628_123#_c_553_n N_A_628_123#_c_554_n
+ N_A_628_123#_c_555_n N_A_628_123#_c_535_n N_A_628_123#_c_586_p
+ N_A_628_123#_c_536_n N_A_628_123#_c_537_n N_A_628_123#_c_538_n
+ N_A_628_123#_c_579_p N_A_628_123#_c_556_n N_A_628_123#_c_557_n
+ N_A_628_123#_c_558_n N_A_628_123#_c_539_n N_A_628_123#_c_540_n
+ PM_SKY130_FD_SC_LP__SDFXTP_1%A_628_123#
x_PM_SKY130_FD_SC_LP__SDFXTP_1%A_823_47# N_A_823_47#_M1004_d N_A_823_47#_M1024_d
+ N_A_823_47#_c_768_n N_A_823_47#_c_769_n N_A_823_47#_c_770_n
+ N_A_823_47#_M1002_g N_A_823_47#_M1012_g N_A_823_47#_M1014_g
+ N_A_823_47#_c_751_n N_A_823_47#_c_752_n N_A_823_47#_c_753_n
+ N_A_823_47#_M1021_g N_A_823_47#_c_755_n N_A_823_47#_c_756_n
+ N_A_823_47#_c_757_n N_A_823_47#_c_758_n N_A_823_47#_c_759_n
+ N_A_823_47#_c_760_n N_A_823_47#_c_827_p N_A_823_47#_c_852_p
+ N_A_823_47#_c_831_p N_A_823_47#_c_761_n N_A_823_47#_c_762_n
+ N_A_823_47#_c_763_n N_A_823_47#_c_764_n N_A_823_47#_c_765_n
+ N_A_823_47#_c_766_n N_A_823_47#_c_767_n PM_SKY130_FD_SC_LP__SDFXTP_1%A_823_47#
x_PM_SKY130_FD_SC_LP__SDFXTP_1%A_1201_99# N_A_1201_99#_M1003_d
+ N_A_1201_99#_M1013_d N_A_1201_99#_M1030_g N_A_1201_99#_M1015_g
+ N_A_1201_99#_c_921_n N_A_1201_99#_c_922_n N_A_1201_99#_c_916_n
+ N_A_1201_99#_c_917_n N_A_1201_99#_c_918_n
+ PM_SKY130_FD_SC_LP__SDFXTP_1%A_1201_99#
x_PM_SKY130_FD_SC_LP__SDFXTP_1%A_1051_125# N_A_1051_125#_M1018_d
+ N_A_1051_125#_M1002_d N_A_1051_125#_M1013_g N_A_1051_125#_M1003_g
+ N_A_1051_125#_c_982_n N_A_1051_125#_c_983_n N_A_1051_125#_c_990_n
+ N_A_1051_125#_c_991_n N_A_1051_125#_c_984_n N_A_1051_125#_c_985_n
+ N_A_1051_125#_c_986_n N_A_1051_125#_c_987_n
+ PM_SKY130_FD_SC_LP__SDFXTP_1%A_1051_125#
x_PM_SKY130_FD_SC_LP__SDFXTP_1%A_1657_383# N_A_1657_383#_M1000_d
+ N_A_1657_383#_M1001_d N_A_1657_383#_M1022_g N_A_1657_383#_M1026_g
+ N_A_1657_383#_c_1068_n N_A_1657_383#_c_1069_n N_A_1657_383#_M1019_g
+ N_A_1657_383#_M1005_g N_A_1657_383#_c_1071_n N_A_1657_383#_c_1081_n
+ N_A_1657_383#_c_1082_n N_A_1657_383#_c_1072_n N_A_1657_383#_c_1083_n
+ N_A_1657_383#_c_1073_n N_A_1657_383#_c_1074_n N_A_1657_383#_c_1075_n
+ N_A_1657_383#_c_1085_n N_A_1657_383#_c_1076_n N_A_1657_383#_c_1077_n
+ PM_SKY130_FD_SC_LP__SDFXTP_1%A_1657_383#
x_PM_SKY130_FD_SC_LP__SDFXTP_1%A_1459_449# N_A_1459_449#_M1014_d
+ N_A_1459_449#_M1008_d N_A_1459_449#_M1000_g N_A_1459_449#_M1001_g
+ N_A_1459_449#_c_1162_n N_A_1459_449#_c_1171_n N_A_1459_449#_c_1172_n
+ N_A_1459_449#_c_1182_n N_A_1459_449#_c_1163_n N_A_1459_449#_c_1164_n
+ N_A_1459_449#_c_1165_n N_A_1459_449#_c_1166_n N_A_1459_449#_c_1167_n
+ N_A_1459_449#_c_1194_n N_A_1459_449#_c_1168_n
+ PM_SKY130_FD_SC_LP__SDFXTP_1%A_1459_449#
x_PM_SKY130_FD_SC_LP__SDFXTP_1%VPWR N_VPWR_M1020_d N_VPWR_M1007_d N_VPWR_M1024_s
+ N_VPWR_M1015_d N_VPWR_M1022_d N_VPWR_M1005_s N_VPWR_c_1265_n N_VPWR_c_1266_n
+ N_VPWR_c_1267_n N_VPWR_c_1268_n N_VPWR_c_1269_n N_VPWR_c_1270_n
+ N_VPWR_c_1271_n N_VPWR_c_1272_n N_VPWR_c_1273_n VPWR N_VPWR_c_1274_n
+ N_VPWR_c_1275_n N_VPWR_c_1276_n N_VPWR_c_1277_n N_VPWR_c_1278_n
+ N_VPWR_c_1264_n N_VPWR_c_1280_n N_VPWR_c_1281_n N_VPWR_c_1282_n
+ N_VPWR_c_1283_n PM_SKY130_FD_SC_LP__SDFXTP_1%VPWR
x_PM_SKY130_FD_SC_LP__SDFXTP_1%A_319_123# N_A_319_123#_M1006_d
+ N_A_319_123#_M1018_s N_A_319_123#_M1028_d N_A_319_123#_M1002_s
+ N_A_319_123#_c_1405_n N_A_319_123#_c_1391_n N_A_319_123#_c_1392_n
+ N_A_319_123#_c_1393_n N_A_319_123#_c_1432_n N_A_319_123#_c_1397_n
+ N_A_319_123#_c_1394_n N_A_319_123#_c_1395_n N_A_319_123#_c_1396_n
+ N_A_319_123#_c_1400_n N_A_319_123#_c_1401_n N_A_319_123#_c_1469_n
+ N_A_319_123#_c_1402_n N_A_319_123#_c_1403_n
+ PM_SKY130_FD_SC_LP__SDFXTP_1%A_319_123#
x_PM_SKY130_FD_SC_LP__SDFXTP_1%Q N_Q_M1019_d N_Q_M1005_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__SDFXTP_1%Q
x_PM_SKY130_FD_SC_LP__SDFXTP_1%VGND N_VGND_M1017_d N_VGND_M1016_d N_VGND_M1004_s
+ N_VGND_M1030_d N_VGND_M1026_d N_VGND_M1019_s N_VGND_c_1533_n N_VGND_c_1534_n
+ N_VGND_c_1535_n N_VGND_c_1536_n N_VGND_c_1537_n N_VGND_c_1538_n
+ N_VGND_c_1539_n N_VGND_c_1540_n N_VGND_c_1541_n N_VGND_c_1542_n
+ N_VGND_c_1543_n N_VGND_c_1544_n N_VGND_c_1545_n VGND N_VGND_c_1546_n
+ N_VGND_c_1547_n N_VGND_c_1548_n N_VGND_c_1549_n N_VGND_c_1550_n
+ N_VGND_c_1551_n N_VGND_c_1552_n PM_SKY130_FD_SC_LP__SDFXTP_1%VGND
cc_1 VNB N_A_78_123#_c_219_n 0.00534261f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.505
cc_2 VNB N_A_78_123#_M1010_g 0.0259309f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=0.825
cc_3 VNB N_A_78_123#_c_221_n 0.0342924f $X=-0.19 $Y=-0.245 $X2=0.18 $Y2=1.655
cc_4 VNB N_A_78_123#_c_222_n 0.00835044f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.385
cc_5 VNB N_A_78_123#_c_223_n 0.024877f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.8
cc_6 VNB N_A_78_123#_c_224_n 0.00428832f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.82
cc_7 VNB N_A_78_123#_c_225_n 0.00867913f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.655
cc_8 VNB N_D_M1006_g 0.0228068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_D_c_310_n 0.0163433f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=0.825
cc_10 VNB D 0.00776366f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=2.295
cc_11 VNB N_D_c_312_n 0.0204224f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=2.385
cc_12 VNB N_SCE_c_359_n 0.0111846f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.455
cc_13 VNB N_SCE_M1017_g 0.034898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_SCE_c_361_n 0.11548f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=0.825
cc_15 VNB N_SCE_c_362_n 0.0132311f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=0.825
cc_16 VNB N_SCE_M1031_g 0.0353074f $X=-0.19 $Y=-0.245 $X2=0.18 $Y2=1.655
cc_17 VNB SCE 0.0134468f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.385
cc_18 VNB N_SCE_c_365_n 0.0421515f $X=-0.19 $Y=-0.245 $X2=0.18 $Y2=0.8
cc_19 VNB N_SCD_M1016_g 0.034992f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.505
cc_20 VNB SCD 0.00666246f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=0.825
cc_21 VNB N_SCD_c_429_n 0.0215545f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=2.775
cc_22 VNB N_CLK_M1009_g 0.0254881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB CLK 0.0074805f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.415
cc_24 VNB N_CLK_c_478_n 0.0482602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_628_123#_M1024_g 0.0105264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_628_123#_M1018_g 0.0372858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_628_123#_c_526_n 0.0247742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_628_123#_c_527_n 0.0319918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_628_123#_c_528_n 0.0204347f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.8
cc_30 VNB N_A_628_123#_c_529_n 0.00864035f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.8
cc_31 VNB N_A_628_123#_c_530_n 0.0268519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_628_123#_c_531_n 0.0131172f $X=-0.19 $Y=-0.245 $X2=0.18 $Y2=1.655
cc_33 VNB N_A_628_123#_c_532_n 0.00480796f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=2.295
cc_34 VNB N_A_628_123#_c_533_n 0.00706032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_628_123#_c_534_n 0.00270469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_628_123#_c_535_n 0.0096533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_628_123#_c_536_n 0.00347595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_628_123#_c_537_n 0.0360127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_628_123#_c_538_n 0.0193654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_628_123#_c_539_n 0.00209904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_628_123#_c_540_n 0.0192221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_823_47#_c_751_n 0.030134f $X=-0.19 $Y=-0.245 $X2=0.18 $Y2=1.655
cc_43 VNB N_A_823_47#_c_752_n 0.0194162f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.47
cc_44 VNB N_A_823_47#_c_753_n 0.0207456f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.6
cc_45 VNB N_A_823_47#_M1021_g 0.0070935f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=2.385
cc_46 VNB N_A_823_47#_c_755_n 0.00121923f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.13
cc_47 VNB N_A_823_47#_c_756_n 0.0210253f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.8
cc_48 VNB N_A_823_47#_c_757_n 0.0276023f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.8
cc_49 VNB N_A_823_47#_c_758_n 0.0282008f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=2.062
cc_50 VNB N_A_823_47#_c_759_n 0.0474029f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.655
cc_51 VNB N_A_823_47#_c_760_n 0.00113394f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=2.13
cc_52 VNB N_A_823_47#_c_761_n 9.76731e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_823_47#_c_762_n 6.35912e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_823_47#_c_763_n 0.00133218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_823_47#_c_764_n 0.0205279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_823_47#_c_765_n 0.00295376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_823_47#_c_766_n 0.0155309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_823_47#_c_767_n 0.0225492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1201_99#_M1030_g 0.0532765f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.415
cc_60 VNB N_A_1201_99#_c_916_n 0.0064692f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.6
cc_61 VNB N_A_1201_99#_c_917_n 0.00273486f $X=-0.19 $Y=-0.245 $X2=1.995
+ $Y2=2.385
cc_62 VNB N_A_1201_99#_c_918_n 0.00669967f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.13
cc_63 VNB N_A_1051_125#_M1013_g 0.0100047f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.415
cc_64 VNB N_A_1051_125#_M1003_g 0.0214165f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=2.295
cc_65 VNB N_A_1051_125#_c_982_n 0.003401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1051_125#_c_983_n 0.00245038f $X=-0.19 $Y=-0.245 $X2=0.18
+ $Y2=1.655
cc_67 VNB N_A_1051_125#_c_984_n 0.020443f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.385
cc_68 VNB N_A_1051_125#_c_985_n 0.00242816f $X=-0.19 $Y=-0.245 $X2=2.115
+ $Y2=2.13
cc_69 VNB N_A_1051_125#_c_986_n 0.0018958f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.8
cc_70 VNB N_A_1051_125#_c_987_n 0.0395603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1657_383#_M1026_g 0.0571689f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=2.295
cc_72 VNB N_A_1657_383#_c_1068_n 0.0149758f $X=-0.19 $Y=-0.245 $X2=2.13
+ $Y2=2.775
cc_73 VNB N_A_1657_383#_c_1069_n 0.0222934f $X=-0.19 $Y=-0.245 $X2=1.145
+ $Y2=1.415
cc_74 VNB N_A_1657_383#_M1005_g 0.00882801f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.6
cc_75 VNB N_A_1657_383#_c_1071_n 0.00611505f $X=-0.19 $Y=-0.245 $X2=1.995
+ $Y2=2.385
cc_76 VNB N_A_1657_383#_c_1072_n 0.00817933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1657_383#_c_1073_n 0.00779647f $X=-0.19 $Y=-0.245 $X2=1.07
+ $Y2=1.82
cc_78 VNB N_A_1657_383#_c_1074_n 2.01195e-19 $X=-0.19 $Y=-0.245 $X2=1.07
+ $Y2=1.82
cc_79 VNB N_A_1657_383#_c_1075_n 0.00854883f $X=-0.19 $Y=-0.245 $X2=1.07
+ $Y2=1.655
cc_80 VNB N_A_1657_383#_c_1076_n 0.00306277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1657_383#_c_1077_n 0.0297569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1459_449#_M1000_g 0.0294906f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.415
cc_83 VNB N_A_1459_449#_c_1162_n 0.0148499f $X=-0.19 $Y=-0.245 $X2=1.145
+ $Y2=1.415
cc_84 VNB N_A_1459_449#_c_1163_n 0.00553998f $X=-0.19 $Y=-0.245 $X2=1.235
+ $Y2=2.385
cc_85 VNB N_A_1459_449#_c_1164_n 9.4756e-19 $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.3
cc_86 VNB N_A_1459_449#_c_1165_n 0.003884f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=2.13
cc_87 VNB N_A_1459_449#_c_1166_n 0.00842365f $X=-0.19 $Y=-0.245 $X2=0.18 $Y2=0.8
cc_88 VNB N_A_1459_449#_c_1167_n 0.0177024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1459_449#_c_1168_n 0.00354405f $X=-0.19 $Y=-0.245 $X2=1.07
+ $Y2=1.82
cc_90 VNB N_VPWR_c_1264_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_319_123#_c_1391_n 9.71559e-19 $X=-0.19 $Y=-0.245 $X2=0.18
+ $Y2=1.655
cc_92 VNB N_A_319_123#_c_1392_n 0.0203331f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.6
cc_93 VNB N_A_319_123#_c_1393_n 0.00455365f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.6
cc_94 VNB N_A_319_123#_c_1394_n 0.00267922f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=2.13
cc_95 VNB N_A_319_123#_c_1395_n 0.012642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_319_123#_c_1396_n 0.00429803f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.8
cc_97 VNB Q 0.0585854f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.505
cc_98 VNB N_VGND_c_1533_n 0.0115803f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.6
cc_99 VNB N_VGND_c_1534_n 0.0202325f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.385
cc_100 VNB N_VGND_c_1535_n 0.0156419f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=2.13
cc_101 VNB N_VGND_c_1536_n 0.0141227f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.8
cc_102 VNB N_VGND_c_1537_n 0.0591092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1538_n 0.00959172f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=1.82
cc_104 VNB N_VGND_c_1539_n 0.0158356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1540_n 0.0256261f $X=-0.19 $Y=-0.245 $X2=2.15 $Y2=2.295
cc_106 VNB N_VGND_c_1541_n 0.00295189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1542_n 0.0467768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1543_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1544_n 0.0206284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1545_n 0.00497312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1546_n 0.0564327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1547_n 0.0201041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1548_n 0.0170759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1549_n 0.574567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1550_n 0.0063235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1551_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1552_n 0.00540978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VPB N_A_78_123#_M1011_g 0.0178384f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.775
cc_119 VPB N_A_78_123#_c_227_n 0.0224415f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.6
cc_120 VPB N_A_78_123#_c_228_n 0.010422f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.385
cc_121 VPB N_A_78_123#_c_222_n 0.0611058f $X=-0.19 $Y=1.655 $X2=1.235 $Y2=2.385
cc_122 VPB N_A_78_123#_c_230_n 0.00222359f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=2.13
cc_123 VPB N_A_78_123#_c_231_n 0.0364876f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=2.13
cc_124 VPB N_A_78_123#_c_224_n 0.026597f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.82
cc_125 VPB N_D_M1028_g 0.0358493f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.505
cc_126 VPB N_D_c_310_n 0.010572f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=0.825
cc_127 VPB N_D_c_315_n 0.021883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB D 0.00326334f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.295
cc_129 VPB N_SCE_c_359_n 0.0338391f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.455
cc_130 VPB N_SCE_c_367_n 0.0202824f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.505
cc_131 VPB N_SCE_c_368_n 0.0287255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_SCE_c_369_n 0.0240684f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.295
cc_133 VPB N_SCE_c_370_n 0.0153071f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.775
cc_134 VPB N_SCD_M1007_g 0.0491484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB SCD 0.0104865f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=0.825
cc_136 VPB N_SCD_c_429_n 0.012275f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.775
cc_137 VPB N_CLK_M1027_g 0.0484179f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.505
cc_138 VPB CLK 0.0115712f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.415
cc_139 VPB N_CLK_c_478_n 0.0308941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_628_123#_M1024_g 0.059423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_628_123#_M1029_g 0.0319409f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.47
cc_142 VPB N_A_628_123#_M1008_g 0.0224766f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.385
cc_143 VPB N_A_628_123#_c_529_n 0.00652564f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.8
cc_144 VPB N_A_628_123#_c_530_n 0.0175193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_628_123#_c_546_n 0.0052442f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.655
cc_146 VPB N_A_628_123#_c_547_n 0.0079471f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=2.13
cc_147 VPB N_A_628_123#_c_548_n 0.00261185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_628_123#_c_533_n 0.0146695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_628_123#_c_550_n 0.0321381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_628_123#_c_551_n 8.07584e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_628_123#_c_534_n 4.26531e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_628_123#_c_553_n 0.00312712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_628_123#_c_554_n 0.00492875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_628_123#_c_555_n 0.0021863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_628_123#_c_556_n 0.0130684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_628_123#_c_557_n 0.00800701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_628_123#_c_558_n 0.0458726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_628_123#_c_539_n 0.00149687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_823_47#_c_768_n 0.0476981f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.505
cc_160 VPB N_A_823_47#_c_769_n 0.0186869f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.655
cc_161 VPB N_A_823_47#_c_770_n 0.0191645f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.415
cc_162 VPB N_A_823_47#_M1021_g 0.0586423f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.385
cc_163 VPB N_A_823_47#_c_756_n 0.00383046f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.8
cc_164 VPB N_A_823_47#_c_757_n 0.0247609f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.8
cc_165 VPB N_A_1201_99#_M1030_g 0.00174663f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.415
cc_166 VPB N_A_1201_99#_M1015_g 0.0228055f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.295
cc_167 VPB N_A_1201_99#_c_921_n 0.00741282f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.775
cc_168 VPB N_A_1201_99#_c_922_n 0.0347364f $X=-0.19 $Y=1.655 $X2=0.18 $Y2=0.965
cc_169 VPB N_A_1201_99#_c_916_n 0.00136379f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.6
cc_170 VPB N_A_1051_125#_M1013_g 0.0429892f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.415
cc_171 VPB N_A_1051_125#_c_982_n 0.00198069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_1051_125#_c_990_n 0.00514897f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.6
cc_173 VPB N_A_1051_125#_c_991_n 0.00197387f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_1657_383#_M1022_g 0.0266993f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.415
cc_175 VPB N_A_1657_383#_M1026_g 0.0130427f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.295
cc_176 VPB N_A_1657_383#_M1005_g 0.0272715f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.6
cc_177 VPB N_A_1657_383#_c_1081_n 0.00886411f $X=-0.19 $Y=1.655 $X2=1.235
+ $Y2=2.385
cc_178 VPB N_A_1657_383#_c_1082_n 0.0434203f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=2.13
cc_179 VPB N_A_1657_383#_c_1083_n 0.0108268f $X=-0.19 $Y=1.655 $X2=0.18
+ $Y2=1.655
cc_180 VPB N_A_1657_383#_c_1074_n 0.00636307f $X=-0.19 $Y=1.655 $X2=1.07
+ $Y2=1.82
cc_181 VPB N_A_1657_383#_c_1085_n 0.00773185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_1657_383#_c_1077_n 0.0137266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_1459_449#_M1001_g 0.0219657f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=2.295
cc_184 VPB N_A_1459_449#_c_1162_n 0.00528566f $X=-0.19 $Y=1.655 $X2=1.145
+ $Y2=1.415
cc_185 VPB N_A_1459_449#_c_1171_n 0.016842f $X=-0.19 $Y=1.655 $X2=0.18 $Y2=0.965
cc_186 VPB N_A_1459_449#_c_1172_n 0.00488504f $X=-0.19 $Y=1.655 $X2=0.615
+ $Y2=2.47
cc_187 VPB N_A_1459_449#_c_1163_n 0.00852879f $X=-0.19 $Y=1.655 $X2=1.235
+ $Y2=2.385
cc_188 VPB N_A_1459_449#_c_1164_n 0.00133499f $X=-0.19 $Y=1.655 $X2=2.115
+ $Y2=2.3
cc_189 VPB N_A_1459_449#_c_1166_n 0.00344759f $X=-0.19 $Y=1.655 $X2=0.18 $Y2=0.8
cc_190 VPB N_A_1459_449#_c_1168_n 6.57797e-19 $X=-0.19 $Y=1.655 $X2=1.07
+ $Y2=1.82
cc_191 VPB N_VPWR_c_1265_n 0.00538161f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.6
cc_192 VPB N_VPWR_c_1266_n 0.00478541f $X=-0.19 $Y=1.655 $X2=1.235 $Y2=2.385
cc_193 VPB N_VPWR_c_1267_n 0.00992298f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=2.13
cc_194 VPB N_VPWR_c_1268_n 0.011508f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.8
cc_195 VPB N_VPWR_c_1269_n 0.0174692f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.062
cc_196 VPB N_VPWR_c_1270_n 0.0416012f $X=-0.19 $Y=1.655 $X2=1.07 $Y2=1.655
cc_197 VPB N_VPWR_c_1271_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1272_n 0.0189835f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1273_n 0.00497553f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=2.295
cc_200 VPB N_VPWR_c_1274_n 0.0294642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1275_n 0.0580555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1276_n 0.0602972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1277_n 0.0187166f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1278_n 0.0182379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1264_n 0.133085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1280_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1281_n 0.0133608f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1282_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1283_n 0.00449427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_319_123#_c_1397_n 0.00904862f $X=-0.19 $Y=1.655 $X2=1.235
+ $Y2=2.385
cc_211 VPB N_A_319_123#_c_1394_n 0.00327935f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=2.13
cc_212 VPB N_A_319_123#_c_1395_n 0.00736068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_319_123#_c_1400_n 0.0203462f $X=-0.19 $Y=1.655 $X2=0.18 $Y2=1.655
cc_214 VPB N_A_319_123#_c_1401_n 0.00107993f $X=-0.19 $Y=1.655 $X2=0.615
+ $Y2=2.062
cc_215 VPB N_A_319_123#_c_1402_n 0.00801464f $X=-0.19 $Y=1.655 $X2=2.15 $Y2=2.13
cc_216 VPB N_A_319_123#_c_1403_n 0.00681549f $X=-0.19 $Y=1.655 $X2=2.15
+ $Y2=2.295
cc_217 VPB Q 0.0571044f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.505
cc_218 N_A_78_123#_M1010_g N_D_M1006_g 0.0220853f $X=1.16 $Y=0.825 $X2=0 $Y2=0
cc_219 N_A_78_123#_M1011_g N_D_M1028_g 0.0258661f $X=2.13 $Y=2.775 $X2=0 $Y2=0
cc_220 N_A_78_123#_c_228_n N_D_M1028_g 0.0112562f $X=1.995 $Y=2.385 $X2=0 $Y2=0
cc_221 N_A_78_123#_c_222_n N_D_M1028_g 0.00339837f $X=1.235 $Y=2.385 $X2=0 $Y2=0
cc_222 N_A_78_123#_c_230_n N_D_M1028_g 0.00165533f $X=2.15 $Y=2.13 $X2=0 $Y2=0
cc_223 N_A_78_123#_c_231_n N_D_M1028_g 0.0201142f $X=2.15 $Y=2.13 $X2=0 $Y2=0
cc_224 N_A_78_123#_c_224_n N_D_M1028_g 8.50836e-19 $X=1.07 $Y=1.82 $X2=0 $Y2=0
cc_225 N_A_78_123#_c_222_n N_D_c_310_n 0.001048f $X=1.235 $Y=2.385 $X2=0 $Y2=0
cc_226 N_A_78_123#_c_225_n N_D_c_310_n 0.0220853f $X=1.07 $Y=1.655 $X2=0 $Y2=0
cc_227 N_A_78_123#_c_228_n N_D_c_315_n 0.00115172f $X=1.995 $Y=2.385 $X2=0 $Y2=0
cc_228 N_A_78_123#_c_224_n N_D_c_315_n 0.0220853f $X=1.07 $Y=1.82 $X2=0 $Y2=0
cc_229 N_A_78_123#_c_219_n D 0.00118992f $X=1.145 $Y=1.505 $X2=0 $Y2=0
cc_230 N_A_78_123#_M1010_g D 0.00331164f $X=1.16 $Y=0.825 $X2=0 $Y2=0
cc_231 N_A_78_123#_c_228_n D 0.0256233f $X=1.995 $Y=2.385 $X2=0 $Y2=0
cc_232 N_A_78_123#_c_222_n D 0.0321341f $X=1.235 $Y=2.385 $X2=0 $Y2=0
cc_233 N_A_78_123#_c_230_n D 0.00981204f $X=2.15 $Y=2.13 $X2=0 $Y2=0
cc_234 N_A_78_123#_c_231_n D 5.79309e-19 $X=2.15 $Y=2.13 $X2=0 $Y2=0
cc_235 N_A_78_123#_c_224_n D 4.91173e-19 $X=1.07 $Y=1.82 $X2=0 $Y2=0
cc_236 N_A_78_123#_c_219_n N_D_c_312_n 0.0220853f $X=1.145 $Y=1.505 $X2=0 $Y2=0
cc_237 N_A_78_123#_c_219_n N_SCE_c_359_n 0.00681208f $X=1.145 $Y=1.505 $X2=0
+ $Y2=0
cc_238 N_A_78_123#_c_221_n N_SCE_c_359_n 0.00562418f $X=0.18 $Y=1.655 $X2=0
+ $Y2=0
cc_239 N_A_78_123#_c_222_n N_SCE_c_359_n 0.0284216f $X=1.235 $Y=2.385 $X2=0
+ $Y2=0
cc_240 N_A_78_123#_c_224_n N_SCE_c_359_n 0.018078f $X=1.07 $Y=1.82 $X2=0 $Y2=0
cc_241 N_A_78_123#_M1010_g N_SCE_M1017_g 0.0203237f $X=1.16 $Y=0.825 $X2=0 $Y2=0
cc_242 N_A_78_123#_c_221_n N_SCE_M1017_g 0.00446622f $X=0.18 $Y=1.655 $X2=0
+ $Y2=0
cc_243 N_A_78_123#_c_227_n N_SCE_c_367_n 0.00765967f $X=0.615 $Y=2.6 $X2=0 $Y2=0
cc_244 N_A_78_123#_c_222_n N_SCE_c_367_n 0.00932616f $X=1.235 $Y=2.385 $X2=0
+ $Y2=0
cc_245 N_A_78_123#_M1010_g N_SCE_c_361_n 0.010454f $X=1.16 $Y=0.825 $X2=0 $Y2=0
cc_246 N_A_78_123#_c_228_n N_SCE_c_368_n 0.00787904f $X=1.995 $Y=2.385 $X2=0
+ $Y2=0
cc_247 N_A_78_123#_c_222_n N_SCE_c_368_n 0.0124974f $X=1.235 $Y=2.385 $X2=0
+ $Y2=0
cc_248 N_A_78_123#_c_224_n N_SCE_c_368_n 0.0214165f $X=1.07 $Y=1.82 $X2=0 $Y2=0
cc_249 N_A_78_123#_c_222_n N_SCE_c_369_n 0.0189218f $X=1.235 $Y=2.385 $X2=0
+ $Y2=0
cc_250 N_A_78_123#_c_227_n N_SCE_c_370_n 8.19448e-19 $X=0.615 $Y=2.6 $X2=0 $Y2=0
cc_251 N_A_78_123#_c_228_n N_SCE_c_370_n 0.00830175f $X=1.995 $Y=2.385 $X2=0
+ $Y2=0
cc_252 N_A_78_123#_c_219_n SCE 0.00520086f $X=1.145 $Y=1.505 $X2=0 $Y2=0
cc_253 N_A_78_123#_M1010_g SCE 0.01498f $X=1.16 $Y=0.825 $X2=0 $Y2=0
cc_254 N_A_78_123#_c_221_n SCE 0.0250942f $X=0.18 $Y=1.655 $X2=0 $Y2=0
cc_255 N_A_78_123#_c_222_n SCE 0.0631019f $X=1.235 $Y=2.385 $X2=0 $Y2=0
cc_256 N_A_78_123#_c_223_n SCE 0.0121528f $X=0.515 $Y=0.8 $X2=0 $Y2=0
cc_257 N_A_78_123#_c_224_n SCE 0.00110013f $X=1.07 $Y=1.82 $X2=0 $Y2=0
cc_258 N_A_78_123#_c_219_n N_SCE_c_365_n 0.00195542f $X=1.145 $Y=1.505 $X2=0
+ $Y2=0
cc_259 N_A_78_123#_M1010_g N_SCE_c_365_n 0.00344643f $X=1.16 $Y=0.825 $X2=0
+ $Y2=0
cc_260 N_A_78_123#_c_221_n N_SCE_c_365_n 0.00833148f $X=0.18 $Y=1.655 $X2=0
+ $Y2=0
cc_261 N_A_78_123#_c_222_n N_SCE_c_365_n 0.00579559f $X=1.235 $Y=2.385 $X2=0
+ $Y2=0
cc_262 N_A_78_123#_c_223_n N_SCE_c_365_n 0.00751427f $X=0.515 $Y=0.8 $X2=0 $Y2=0
cc_263 N_A_78_123#_M1011_g N_SCD_M1007_g 0.0356706f $X=2.13 $Y=2.775 $X2=0 $Y2=0
cc_264 N_A_78_123#_c_228_n N_SCD_M1007_g 5.14196e-19 $X=1.995 $Y=2.385 $X2=0
+ $Y2=0
cc_265 N_A_78_123#_c_230_n N_SCD_M1007_g 4.82958e-19 $X=2.15 $Y=2.13 $X2=0 $Y2=0
cc_266 N_A_78_123#_c_231_n N_SCD_M1007_g 0.020401f $X=2.15 $Y=2.13 $X2=0 $Y2=0
cc_267 N_A_78_123#_c_228_n SCD 3.49453e-19 $X=1.995 $Y=2.385 $X2=0 $Y2=0
cc_268 N_A_78_123#_c_230_n SCD 0.0193856f $X=2.15 $Y=2.13 $X2=0 $Y2=0
cc_269 N_A_78_123#_c_231_n SCD 0.00528247f $X=2.15 $Y=2.13 $X2=0 $Y2=0
cc_270 N_A_78_123#_c_222_n N_VPWR_M1020_d 0.00268916f $X=1.235 $Y=2.385
+ $X2=-0.19 $Y2=-0.245
cc_271 N_A_78_123#_c_222_n N_VPWR_c_1265_n 0.0216849f $X=1.235 $Y=2.385 $X2=0
+ $Y2=0
cc_272 N_A_78_123#_M1011_g N_VPWR_c_1270_n 0.0037886f $X=2.13 $Y=2.775 $X2=0
+ $Y2=0
cc_273 N_A_78_123#_c_227_n N_VPWR_c_1274_n 0.0176612f $X=0.615 $Y=2.6 $X2=0
+ $Y2=0
cc_274 N_A_78_123#_M1020_s N_VPWR_c_1264_n 0.00216391f $X=0.49 $Y=2.455 $X2=0
+ $Y2=0
cc_275 N_A_78_123#_M1011_g N_VPWR_c_1264_n 0.00564534f $X=2.13 $Y=2.775 $X2=0
+ $Y2=0
cc_276 N_A_78_123#_c_227_n N_VPWR_c_1264_n 0.0123808f $X=0.615 $Y=2.6 $X2=0
+ $Y2=0
cc_277 N_A_78_123#_c_228_n N_VPWR_c_1264_n 0.0155374f $X=1.995 $Y=2.385 $X2=0
+ $Y2=0
cc_278 N_A_78_123#_c_222_n N_VPWR_c_1264_n 0.00663315f $X=1.235 $Y=2.385 $X2=0
+ $Y2=0
cc_279 N_A_78_123#_c_228_n A_283_491# 0.00196273f $X=1.995 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_280 N_A_78_123#_c_228_n N_A_319_123#_M1028_d 0.00170524f $X=1.995 $Y=2.385
+ $X2=0 $Y2=0
cc_281 N_A_78_123#_M1011_g N_A_319_123#_c_1405_n 0.0129223f $X=2.13 $Y=2.775
+ $X2=0 $Y2=0
cc_282 N_A_78_123#_c_228_n N_A_319_123#_c_1405_n 0.0254534f $X=1.995 $Y=2.385
+ $X2=0 $Y2=0
cc_283 N_A_78_123#_c_231_n N_A_319_123#_c_1405_n 0.00247025f $X=2.15 $Y=2.13
+ $X2=0 $Y2=0
cc_284 N_A_78_123#_c_230_n N_A_319_123#_c_1394_n 0.00177573f $X=2.15 $Y=2.13
+ $X2=0 $Y2=0
cc_285 N_A_78_123#_c_228_n N_A_319_123#_c_1401_n 0.00114996f $X=1.995 $Y=2.385
+ $X2=0 $Y2=0
cc_286 N_A_78_123#_M1011_g N_A_319_123#_c_1403_n 0.00402491f $X=2.13 $Y=2.775
+ $X2=0 $Y2=0
cc_287 N_A_78_123#_c_228_n N_A_319_123#_c_1403_n 0.0124689f $X=1.995 $Y=2.385
+ $X2=0 $Y2=0
cc_288 N_A_78_123#_c_230_n N_A_319_123#_c_1403_n 0.0194629f $X=2.15 $Y=2.13
+ $X2=0 $Y2=0
cc_289 N_A_78_123#_c_231_n N_A_319_123#_c_1403_n 0.0017175f $X=2.15 $Y=2.13
+ $X2=0 $Y2=0
cc_290 N_A_78_123#_M1010_g N_VGND_c_1533_n 0.00140973f $X=1.16 $Y=0.825 $X2=0
+ $Y2=0
cc_291 N_A_78_123#_c_223_n N_VGND_c_1540_n 0.0096573f $X=0.515 $Y=0.8 $X2=0
+ $Y2=0
cc_292 N_A_78_123#_M1010_g N_VGND_c_1549_n 9.15321e-19 $X=1.16 $Y=0.825 $X2=0
+ $Y2=0
cc_293 N_A_78_123#_c_223_n N_VGND_c_1549_n 0.0154096f $X=0.515 $Y=0.8 $X2=0
+ $Y2=0
cc_294 N_D_M1006_g N_SCE_c_361_n 0.00896132f $X=1.52 $Y=0.825 $X2=0 $Y2=0
cc_295 D N_SCE_c_361_n 0.00546336f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_296 N_D_M1028_g N_SCE_c_368_n 0.064877f $X=1.7 $Y=2.775 $X2=0 $Y2=0
cc_297 N_D_M1006_g N_SCE_M1031_g 0.00717696f $X=1.52 $Y=0.825 $X2=0 $Y2=0
cc_298 D N_SCE_M1031_g 0.00768673f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_299 N_D_M1006_g SCE 0.00197417f $X=1.52 $Y=0.825 $X2=0 $Y2=0
cc_300 D SCE 0.0275277f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_301 N_D_c_310_n SCD 0.00353105f $X=1.61 $Y=1.79 $X2=0 $Y2=0
cc_302 D SCD 0.0213749f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_303 D N_SCD_c_429_n 6.03645e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_304 N_D_c_312_n N_SCD_c_429_n 0.005387f $X=1.61 $Y=1.45 $X2=0 $Y2=0
cc_305 N_D_M1028_g N_VPWR_c_1270_n 0.00550964f $X=1.7 $Y=2.775 $X2=0 $Y2=0
cc_306 N_D_M1028_g N_VPWR_c_1264_n 0.00626038f $X=1.7 $Y=2.775 $X2=0 $Y2=0
cc_307 D N_A_319_123#_M1006_d 0.00431772f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_308 N_D_M1028_g N_A_319_123#_c_1405_n 0.00614187f $X=1.7 $Y=2.775 $X2=0 $Y2=0
cc_309 N_D_M1006_g N_A_319_123#_c_1391_n 0.00126227f $X=1.52 $Y=0.825 $X2=0
+ $Y2=0
cc_310 D N_A_319_123#_c_1391_n 0.037162f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_311 N_D_M1006_g N_A_319_123#_c_1393_n 6.60134e-19 $X=1.52 $Y=0.825 $X2=0
+ $Y2=0
cc_312 D N_A_319_123#_c_1393_n 0.0148404f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_313 N_D_c_312_n N_A_319_123#_c_1393_n 9.31826e-19 $X=1.61 $Y=1.45 $X2=0 $Y2=0
cc_314 D N_VGND_c_1533_n 0.0153043f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_315 D N_VGND_c_1542_n 0.0124231f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_316 D N_VGND_c_1549_n 0.0102181f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_317 N_SCE_M1031_g N_SCD_M1016_g 0.0405382f $X=2.245 $Y=0.825 $X2=0 $Y2=0
cc_318 N_SCE_M1031_g SCD 7.59348e-19 $X=2.245 $Y=0.825 $X2=0 $Y2=0
cc_319 N_SCE_c_367_n N_VPWR_c_1265_n 0.00355035f $X=0.83 $Y=2.345 $X2=0 $Y2=0
cc_320 N_SCE_c_368_n N_VPWR_c_1265_n 0.00106002f $X=1.265 $Y=2.27 $X2=0 $Y2=0
cc_321 N_SCE_c_370_n N_VPWR_c_1265_n 0.0037301f $X=1.34 $Y=2.345 $X2=0 $Y2=0
cc_322 N_SCE_c_370_n N_VPWR_c_1270_n 0.00585385f $X=1.34 $Y=2.345 $X2=0 $Y2=0
cc_323 N_SCE_c_367_n N_VPWR_c_1274_n 0.00549943f $X=0.83 $Y=2.345 $X2=0 $Y2=0
cc_324 N_SCE_c_367_n N_VPWR_c_1264_n 0.00766972f $X=0.83 $Y=2.345 $X2=0 $Y2=0
cc_325 N_SCE_c_370_n N_VPWR_c_1264_n 0.00640801f $X=1.34 $Y=2.345 $X2=0 $Y2=0
cc_326 N_SCE_c_370_n N_A_319_123#_c_1405_n 9.11007e-19 $X=1.34 $Y=2.345 $X2=0
+ $Y2=0
cc_327 N_SCE_c_361_n N_A_319_123#_c_1391_n 0.00253772f $X=2.17 $Y=0.2 $X2=0
+ $Y2=0
cc_328 N_SCE_M1031_g N_A_319_123#_c_1391_n 0.009902f $X=2.245 $Y=0.825 $X2=0
+ $Y2=0
cc_329 N_SCE_M1031_g N_A_319_123#_c_1392_n 0.00784684f $X=2.245 $Y=0.825 $X2=0
+ $Y2=0
cc_330 N_SCE_M1031_g N_A_319_123#_c_1393_n 6.05142e-19 $X=2.245 $Y=0.825 $X2=0
+ $Y2=0
cc_331 N_SCE_M1017_g N_VGND_c_1533_n 0.0118153f $X=0.73 $Y=0.825 $X2=0 $Y2=0
cc_332 N_SCE_c_361_n N_VGND_c_1533_n 0.0182907f $X=2.17 $Y=0.2 $X2=0 $Y2=0
cc_333 SCE N_VGND_c_1533_n 0.013405f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_334 N_SCE_c_361_n N_VGND_c_1534_n 0.0102903f $X=2.17 $Y=0.2 $X2=0 $Y2=0
cc_335 N_SCE_M1031_g N_VGND_c_1534_n 0.00168632f $X=2.245 $Y=0.825 $X2=0 $Y2=0
cc_336 N_SCE_c_362_n N_VGND_c_1540_n 0.00693208f $X=0.805 $Y=0.2 $X2=0 $Y2=0
cc_337 N_SCE_c_361_n N_VGND_c_1542_n 0.037467f $X=2.17 $Y=0.2 $X2=0 $Y2=0
cc_338 N_SCE_c_361_n N_VGND_c_1549_n 0.0545129f $X=2.17 $Y=0.2 $X2=0 $Y2=0
cc_339 N_SCE_c_362_n N_VGND_c_1549_n 0.0108676f $X=0.805 $Y=0.2 $X2=0 $Y2=0
cc_340 N_SCD_M1016_g N_CLK_M1009_g 0.0182944f $X=2.605 $Y=0.825 $X2=0 $Y2=0
cc_341 N_SCD_M1007_g N_CLK_c_478_n 0.0405651f $X=2.6 $Y=2.775 $X2=0 $Y2=0
cc_342 SCD N_CLK_c_478_n 9.95358e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_343 N_SCD_c_429_n N_CLK_c_478_n 0.0182944f $X=2.515 $Y=1.59 $X2=0 $Y2=0
cc_344 N_SCD_M1007_g N_A_628_123#_c_546_n 3.43378e-19 $X=2.6 $Y=2.775 $X2=0
+ $Y2=0
cc_345 N_SCD_M1007_g N_A_628_123#_c_548_n 3.49442e-19 $X=2.6 $Y=2.775 $X2=0
+ $Y2=0
cc_346 N_SCD_M1007_g N_VPWR_c_1266_n 0.00617328f $X=2.6 $Y=2.775 $X2=0 $Y2=0
cc_347 N_SCD_M1007_g N_VPWR_c_1270_n 0.00502699f $X=2.6 $Y=2.775 $X2=0 $Y2=0
cc_348 N_SCD_M1007_g N_VPWR_c_1264_n 0.00630632f $X=2.6 $Y=2.775 $X2=0 $Y2=0
cc_349 N_SCD_M1007_g N_A_319_123#_c_1405_n 0.00940795f $X=2.6 $Y=2.775 $X2=0
+ $Y2=0
cc_350 N_SCD_M1016_g N_A_319_123#_c_1391_n 0.00178706f $X=2.605 $Y=0.825 $X2=0
+ $Y2=0
cc_351 N_SCD_M1016_g N_A_319_123#_c_1392_n 0.0161018f $X=2.605 $Y=0.825 $X2=0
+ $Y2=0
cc_352 SCD N_A_319_123#_c_1392_n 0.0405459f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_353 N_SCD_c_429_n N_A_319_123#_c_1392_n 0.00440502f $X=2.515 $Y=1.59 $X2=0
+ $Y2=0
cc_354 SCD N_A_319_123#_c_1393_n 0.0183626f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_355 N_SCD_M1007_g N_A_319_123#_c_1432_n 0.00390891f $X=2.6 $Y=2.775 $X2=0
+ $Y2=0
cc_356 N_SCD_M1007_g N_A_319_123#_c_1397_n 3.91988e-19 $X=2.6 $Y=2.775 $X2=0
+ $Y2=0
cc_357 SCD N_A_319_123#_c_1397_n 5.68901e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_358 N_SCD_M1007_g N_A_319_123#_c_1394_n 0.00412569f $X=2.6 $Y=2.775 $X2=0
+ $Y2=0
cc_359 N_SCD_M1016_g N_A_319_123#_c_1394_n 0.00338371f $X=2.605 $Y=0.825 $X2=0
+ $Y2=0
cc_360 SCD N_A_319_123#_c_1394_n 0.0251628f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_361 N_SCD_c_429_n N_A_319_123#_c_1394_n 7.26895e-19 $X=2.515 $Y=1.59 $X2=0
+ $Y2=0
cc_362 N_SCD_M1007_g N_A_319_123#_c_1401_n 0.00396622f $X=2.6 $Y=2.775 $X2=0
+ $Y2=0
cc_363 SCD N_A_319_123#_c_1401_n 0.0010755f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_364 N_SCD_M1007_g N_A_319_123#_c_1403_n 0.0161925f $X=2.6 $Y=2.775 $X2=0
+ $Y2=0
cc_365 SCD N_A_319_123#_c_1403_n 0.0186001f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_366 N_SCD_c_429_n N_A_319_123#_c_1403_n 7.90547e-19 $X=2.515 $Y=1.59 $X2=0
+ $Y2=0
cc_367 N_SCD_M1016_g N_VGND_c_1534_n 0.00969346f $X=2.605 $Y=0.825 $X2=0 $Y2=0
cc_368 N_SCD_M1016_g N_VGND_c_1542_n 0.00349617f $X=2.605 $Y=0.825 $X2=0 $Y2=0
cc_369 N_SCD_M1016_g N_VGND_c_1549_n 0.00396651f $X=2.605 $Y=0.825 $X2=0 $Y2=0
cc_370 CLK N_A_628_123#_M1024_g 0.00339315f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_371 N_CLK_c_478_n N_A_628_123#_M1024_g 0.00956896f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_372 CLK N_A_628_123#_c_527_n 0.00221723f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_373 N_CLK_c_478_n N_A_628_123#_c_527_n 0.0095844f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_374 N_CLK_M1009_g N_A_628_123#_c_531_n 0.00484488f $X=3.065 $Y=0.825 $X2=0
+ $Y2=0
cc_375 CLK N_A_628_123#_c_531_n 0.0350806f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_376 N_CLK_c_478_n N_A_628_123#_c_531_n 0.00527802f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_377 N_CLK_M1027_g N_A_628_123#_c_546_n 0.00597339f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_378 CLK N_A_628_123#_c_547_n 0.0180379f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_379 N_CLK_M1027_g N_A_628_123#_c_548_n 0.00454828f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_380 CLK N_A_628_123#_c_548_n 0.0140992f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_381 N_CLK_c_478_n N_A_628_123#_c_548_n 0.00356541f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_382 CLK N_A_628_123#_c_533_n 0.0881418f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_383 N_CLK_c_478_n N_A_628_123#_c_533_n 0.00134726f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_384 N_CLK_M1009_g N_A_628_123#_c_538_n 0.00579926f $X=3.065 $Y=0.825 $X2=0
+ $Y2=0
cc_385 N_CLK_M1027_g N_VPWR_c_1266_n 0.00320608f $X=3.065 $Y=2.775 $X2=0 $Y2=0
cc_386 N_CLK_M1027_g N_VPWR_c_1267_n 0.00266635f $X=3.065 $Y=2.775 $X2=0 $Y2=0
cc_387 N_CLK_M1027_g N_VPWR_c_1272_n 0.00549943f $X=3.065 $Y=2.775 $X2=0 $Y2=0
cc_388 N_CLK_M1027_g N_VPWR_c_1264_n 0.0112899f $X=3.065 $Y=2.775 $X2=0 $Y2=0
cc_389 N_CLK_M1009_g N_A_319_123#_c_1392_n 0.00648423f $X=3.065 $Y=0.825 $X2=0
+ $Y2=0
cc_390 CLK N_A_319_123#_c_1392_n 0.0117868f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_391 N_CLK_c_478_n N_A_319_123#_c_1392_n 0.00412511f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_392 N_CLK_M1027_g N_A_319_123#_c_1432_n 4.80547e-19 $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_393 N_CLK_M1027_g N_A_319_123#_c_1397_n 0.00581246f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_394 CLK N_A_319_123#_c_1397_n 0.0133127f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_395 N_CLK_M1027_g N_A_319_123#_c_1394_n 0.00327874f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_396 CLK N_A_319_123#_c_1394_n 0.0501437f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_397 N_CLK_c_478_n N_A_319_123#_c_1394_n 0.0157036f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_398 N_CLK_M1027_g N_A_319_123#_c_1400_n 0.0104728f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_399 CLK N_A_319_123#_c_1400_n 0.0121302f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_400 N_CLK_c_478_n N_A_319_123#_c_1400_n 0.00269615f $X=3.34 $Y=1.375 $X2=0
+ $Y2=0
cc_401 N_CLK_M1027_g N_A_319_123#_c_1401_n 0.00135808f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_402 N_CLK_M1027_g N_A_319_123#_c_1403_n 0.0037681f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_403 CLK N_A_319_123#_c_1403_n 4.19579e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_404 N_CLK_M1009_g N_VGND_c_1534_n 0.00350978f $X=3.065 $Y=0.825 $X2=0 $Y2=0
cc_405 N_CLK_M1009_g N_VGND_c_1535_n 0.00149837f $X=3.065 $Y=0.825 $X2=0 $Y2=0
cc_406 N_CLK_M1009_g N_VGND_c_1544_n 0.00405474f $X=3.065 $Y=0.825 $X2=0 $Y2=0
cc_407 N_CLK_M1009_g N_VGND_c_1549_n 0.00472204f $X=3.065 $Y=0.825 $X2=0 $Y2=0
cc_408 N_A_628_123#_c_577_p N_A_823_47#_M1024_d 0.00824917f $X=4.15 $Y=2.895
+ $X2=0 $Y2=0
cc_409 N_A_628_123#_c_550_n N_A_823_47#_M1024_d 0.00798963f $X=5.76 $Y=2.98
+ $X2=0 $Y2=0
cc_410 N_A_628_123#_c_579_p N_A_823_47#_M1024_d 0.00120743f $X=4.05 $Y=2.47
+ $X2=0 $Y2=0
cc_411 N_A_628_123#_M1029_g N_A_823_47#_c_768_n 0.0176811f $X=5.71 $Y=2.455
+ $X2=0 $Y2=0
cc_412 N_A_628_123#_c_529_n N_A_823_47#_c_768_n 0.01606f $X=5.255 $Y=1.61 $X2=0
+ $Y2=0
cc_413 N_A_628_123#_c_553_n N_A_823_47#_c_768_n 2.99951e-19 $X=5.845 $Y=2.635
+ $X2=0 $Y2=0
cc_414 N_A_628_123#_c_550_n N_A_823_47#_c_770_n 0.00651141f $X=5.76 $Y=2.98
+ $X2=0 $Y2=0
cc_415 N_A_628_123#_c_553_n N_A_823_47#_c_770_n 8.18406e-19 $X=5.845 $Y=2.635
+ $X2=0 $Y2=0
cc_416 N_A_628_123#_c_535_n N_A_823_47#_c_751_n 0.00581732f $X=7.99 $Y=1.38
+ $X2=0 $Y2=0
cc_417 N_A_628_123#_c_586_p N_A_823_47#_c_751_n 0.00470006f $X=7.605 $Y=1.38
+ $X2=0 $Y2=0
cc_418 N_A_628_123#_c_536_n N_A_823_47#_c_751_n 0.0041038f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_419 N_A_628_123#_c_535_n N_A_823_47#_c_752_n 0.0110904f $X=7.99 $Y=1.38 $X2=0
+ $Y2=0
cc_420 N_A_628_123#_c_537_n N_A_823_47#_c_752_n 0.00554227f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_421 N_A_628_123#_c_535_n N_A_823_47#_c_753_n 0.00700034f $X=7.99 $Y=1.38
+ $X2=0 $Y2=0
cc_422 N_A_628_123#_c_586_p N_A_823_47#_c_753_n 0.00166088f $X=7.605 $Y=1.38
+ $X2=0 $Y2=0
cc_423 N_A_628_123#_c_557_n N_A_823_47#_c_753_n 2.28767e-19 $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_424 N_A_628_123#_c_558_n N_A_823_47#_c_753_n 0.0127591f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_425 N_A_628_123#_c_539_n N_A_823_47#_c_753_n 0.00665478f $X=7.477 $Y=1.755
+ $X2=0 $Y2=0
cc_426 N_A_628_123#_M1008_g N_A_823_47#_M1021_g 0.0103687f $X=7.22 $Y=2.665
+ $X2=0 $Y2=0
cc_427 N_A_628_123#_c_555_n N_A_823_47#_M1021_g 0.00127806f $X=7.435 $Y=2.635
+ $X2=0 $Y2=0
cc_428 N_A_628_123#_c_558_n N_A_823_47#_M1021_g 0.0123101f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_429 N_A_628_123#_c_539_n N_A_823_47#_M1021_g 0.0043028f $X=7.477 $Y=1.755
+ $X2=0 $Y2=0
cc_430 N_A_628_123#_c_526_n N_A_823_47#_c_755_n 0.00293824f $X=3.95 $Y=0.765
+ $X2=0 $Y2=0
cc_431 N_A_628_123#_c_532_n N_A_823_47#_c_755_n 0.00711951f $X=4.05 $Y=0.985
+ $X2=0 $Y2=0
cc_432 N_A_628_123#_M1024_g N_A_823_47#_c_756_n 0.00377871f $X=4.05 $Y=2.725
+ $X2=0 $Y2=0
cc_433 N_A_628_123#_M1018_g N_A_823_47#_c_756_n 0.00465711f $X=5.18 $Y=0.835
+ $X2=0 $Y2=0
cc_434 N_A_628_123#_c_526_n N_A_823_47#_c_756_n 0.00801051f $X=3.95 $Y=0.765
+ $X2=0 $Y2=0
cc_435 N_A_628_123#_c_528_n N_A_823_47#_c_756_n 9.65879e-19 $X=3.955 $Y=1.435
+ $X2=0 $Y2=0
cc_436 N_A_628_123#_c_532_n N_A_823_47#_c_756_n 0.0229767f $X=4.05 $Y=0.985
+ $X2=0 $Y2=0
cc_437 N_A_628_123#_c_533_n N_A_823_47#_c_756_n 0.109768f $X=4.05 $Y=2.385 $X2=0
+ $Y2=0
cc_438 N_A_628_123#_c_577_p N_A_823_47#_c_756_n 0.0124151f $X=4.15 $Y=2.895
+ $X2=0 $Y2=0
cc_439 N_A_628_123#_c_550_n N_A_823_47#_c_756_n 0.0137058f $X=5.76 $Y=2.98 $X2=0
+ $Y2=0
cc_440 N_A_628_123#_c_579_p N_A_823_47#_c_756_n 0.0129302f $X=4.05 $Y=2.47 $X2=0
+ $Y2=0
cc_441 N_A_628_123#_M1024_g N_A_823_47#_c_757_n 0.0418615f $X=4.05 $Y=2.725
+ $X2=0 $Y2=0
cc_442 N_A_628_123#_c_529_n N_A_823_47#_c_757_n 0.00671722f $X=5.255 $Y=1.61
+ $X2=0 $Y2=0
cc_443 N_A_628_123#_c_533_n N_A_823_47#_c_757_n 0.00450189f $X=4.05 $Y=2.385
+ $X2=0 $Y2=0
cc_444 N_A_628_123#_M1018_g N_A_823_47#_c_758_n 0.00760724f $X=5.18 $Y=0.835
+ $X2=0 $Y2=0
cc_445 N_A_628_123#_M1018_g N_A_823_47#_c_759_n 0.00132716f $X=5.18 $Y=0.835
+ $X2=0 $Y2=0
cc_446 N_A_628_123#_M1018_g N_A_823_47#_c_760_n 7.27288e-19 $X=5.18 $Y=0.835
+ $X2=0 $Y2=0
cc_447 N_A_628_123#_c_535_n N_A_823_47#_c_763_n 0.0120778f $X=7.99 $Y=1.38 $X2=0
+ $Y2=0
cc_448 N_A_628_123#_c_586_p N_A_823_47#_c_763_n 0.014306f $X=7.605 $Y=1.38 $X2=0
+ $Y2=0
cc_449 N_A_628_123#_c_536_n N_A_823_47#_c_763_n 0.0159164f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_450 N_A_628_123#_c_537_n N_A_823_47#_c_763_n 0.00101459f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_451 N_A_628_123#_c_540_n N_A_823_47#_c_763_n 0.00162702f $X=8.155 $Y=0.855
+ $X2=0 $Y2=0
cc_452 N_A_628_123#_c_536_n N_A_823_47#_c_764_n 0.00137437f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_453 N_A_628_123#_c_537_n N_A_823_47#_c_764_n 0.0184306f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_454 N_A_628_123#_M1018_g N_A_823_47#_c_766_n 0.0105839f $X=5.18 $Y=0.835
+ $X2=0 $Y2=0
cc_455 N_A_628_123#_c_530_n N_A_823_47#_c_766_n 0.00673494f $X=5.635 $Y=1.61
+ $X2=0 $Y2=0
cc_456 N_A_628_123#_c_537_n N_A_823_47#_c_767_n 2.18342e-19 $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_457 N_A_628_123#_c_540_n N_A_823_47#_c_767_n 0.00736704f $X=8.155 $Y=0.855
+ $X2=0 $Y2=0
cc_458 N_A_628_123#_c_554_n N_A_1201_99#_M1013_d 0.00427673f $X=7.35 $Y=2.72
+ $X2=0 $Y2=0
cc_459 N_A_628_123#_c_530_n N_A_1201_99#_M1030_g 0.020797f $X=5.635 $Y=1.61
+ $X2=0 $Y2=0
cc_460 N_A_628_123#_c_534_n N_A_1201_99#_M1030_g 0.0048229f $X=5.76 $Y=1.61
+ $X2=0 $Y2=0
cc_461 N_A_628_123#_c_554_n N_A_1201_99#_M1015_g 0.0128803f $X=7.35 $Y=2.72
+ $X2=0 $Y2=0
cc_462 N_A_628_123#_c_556_n N_A_1201_99#_M1015_g 0.00448001f $X=5.845 $Y=2.72
+ $X2=0 $Y2=0
cc_463 N_A_628_123#_M1029_g N_A_1201_99#_c_921_n 5.71018e-19 $X=5.71 $Y=2.455
+ $X2=0 $Y2=0
cc_464 N_A_628_123#_c_534_n N_A_1201_99#_c_921_n 0.00164692f $X=5.76 $Y=1.61
+ $X2=0 $Y2=0
cc_465 N_A_628_123#_c_553_n N_A_1201_99#_c_921_n 0.0602829f $X=5.845 $Y=2.635
+ $X2=0 $Y2=0
cc_466 N_A_628_123#_c_554_n N_A_1201_99#_c_921_n 0.0579004f $X=7.35 $Y=2.72
+ $X2=0 $Y2=0
cc_467 N_A_628_123#_M1029_g N_A_1201_99#_c_922_n 0.0576764f $X=5.71 $Y=2.455
+ $X2=0 $Y2=0
cc_468 N_A_628_123#_c_553_n N_A_1201_99#_c_922_n 0.00426513f $X=5.845 $Y=2.635
+ $X2=0 $Y2=0
cc_469 N_A_628_123#_c_554_n N_A_1201_99#_c_922_n 5.27217e-19 $X=7.35 $Y=2.72
+ $X2=0 $Y2=0
cc_470 N_A_628_123#_M1008_g N_A_1201_99#_c_916_n 0.00635692f $X=7.22 $Y=2.665
+ $X2=0 $Y2=0
cc_471 N_A_628_123#_c_554_n N_A_1201_99#_c_916_n 0.00880073f $X=7.35 $Y=2.72
+ $X2=0 $Y2=0
cc_472 N_A_628_123#_c_586_p N_A_1201_99#_c_916_n 0.00737783f $X=7.605 $Y=1.38
+ $X2=0 $Y2=0
cc_473 N_A_628_123#_c_557_n N_A_1201_99#_c_916_n 0.0456723f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_474 N_A_628_123#_c_558_n N_A_1201_99#_c_916_n 0.0102508f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_475 N_A_628_123#_c_539_n N_A_1201_99#_c_916_n 0.0161092f $X=7.477 $Y=1.755
+ $X2=0 $Y2=0
cc_476 N_A_628_123#_c_586_p N_A_1201_99#_c_918_n 0.00330189f $X=7.605 $Y=1.38
+ $X2=0 $Y2=0
cc_477 N_A_628_123#_c_558_n N_A_1201_99#_c_918_n 0.00342102f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_478 N_A_628_123#_c_554_n N_A_1051_125#_M1013_g 0.01246f $X=7.35 $Y=2.72 $X2=0
+ $Y2=0
cc_479 N_A_628_123#_c_557_n N_A_1051_125#_M1013_g 2.02219e-19 $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_480 N_A_628_123#_c_558_n N_A_1051_125#_M1013_g 0.0528451f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_481 N_A_628_123#_c_539_n N_A_1051_125#_M1013_g 4.88046e-19 $X=7.477 $Y=1.755
+ $X2=0 $Y2=0
cc_482 N_A_628_123#_M1018_g N_A_1051_125#_c_982_n 0.00322844f $X=5.18 $Y=0.835
+ $X2=0 $Y2=0
cc_483 N_A_628_123#_M1029_g N_A_1051_125#_c_982_n 0.00177245f $X=5.71 $Y=2.455
+ $X2=0 $Y2=0
cc_484 N_A_628_123#_c_529_n N_A_1051_125#_c_982_n 0.00659904f $X=5.255 $Y=1.61
+ $X2=0 $Y2=0
cc_485 N_A_628_123#_c_530_n N_A_1051_125#_c_982_n 0.0088935f $X=5.635 $Y=1.61
+ $X2=0 $Y2=0
cc_486 N_A_628_123#_c_534_n N_A_1051_125#_c_982_n 0.0132506f $X=5.76 $Y=1.61
+ $X2=0 $Y2=0
cc_487 N_A_628_123#_c_553_n N_A_1051_125#_c_982_n 0.00534525f $X=5.845 $Y=2.635
+ $X2=0 $Y2=0
cc_488 N_A_628_123#_M1018_g N_A_1051_125#_c_983_n 0.00150568f $X=5.18 $Y=0.835
+ $X2=0 $Y2=0
cc_489 N_A_628_123#_M1029_g N_A_1051_125#_c_990_n 0.00296985f $X=5.71 $Y=2.455
+ $X2=0 $Y2=0
cc_490 N_A_628_123#_c_530_n N_A_1051_125#_c_990_n 0.00693225f $X=5.635 $Y=1.61
+ $X2=0 $Y2=0
cc_491 N_A_628_123#_c_534_n N_A_1051_125#_c_990_n 0.00901284f $X=5.76 $Y=1.61
+ $X2=0 $Y2=0
cc_492 N_A_628_123#_c_553_n N_A_1051_125#_c_990_n 0.0131414f $X=5.845 $Y=2.635
+ $X2=0 $Y2=0
cc_493 N_A_628_123#_M1029_g N_A_1051_125#_c_991_n 0.00151965f $X=5.71 $Y=2.455
+ $X2=0 $Y2=0
cc_494 N_A_628_123#_c_550_n N_A_1051_125#_c_991_n 0.0108566f $X=5.76 $Y=2.98
+ $X2=0 $Y2=0
cc_495 N_A_628_123#_c_553_n N_A_1051_125#_c_991_n 0.0268379f $X=5.845 $Y=2.635
+ $X2=0 $Y2=0
cc_496 N_A_628_123#_c_530_n N_A_1051_125#_c_984_n 0.00479544f $X=5.635 $Y=1.61
+ $X2=0 $Y2=0
cc_497 N_A_628_123#_c_534_n N_A_1051_125#_c_984_n 0.0321181f $X=5.76 $Y=1.61
+ $X2=0 $Y2=0
cc_498 N_A_628_123#_M1018_g N_A_1051_125#_c_985_n 0.0144786f $X=5.18 $Y=0.835
+ $X2=0 $Y2=0
cc_499 N_A_628_123#_c_530_n N_A_1051_125#_c_985_n 0.00675528f $X=5.635 $Y=1.61
+ $X2=0 $Y2=0
cc_500 N_A_628_123#_c_534_n N_A_1051_125#_c_985_n 0.00366136f $X=5.76 $Y=1.61
+ $X2=0 $Y2=0
cc_501 N_A_628_123#_c_535_n N_A_1657_383#_M1026_g 8.618e-19 $X=7.99 $Y=1.38
+ $X2=0 $Y2=0
cc_502 N_A_628_123#_c_536_n N_A_1657_383#_M1026_g 9.14012e-19 $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_503 N_A_628_123#_c_540_n N_A_1657_383#_M1026_g 0.0618155f $X=8.155 $Y=0.855
+ $X2=0 $Y2=0
cc_504 N_A_628_123#_c_554_n N_A_1459_449#_M1008_d 0.00468341f $X=7.35 $Y=2.72
+ $X2=0 $Y2=0
cc_505 N_A_628_123#_c_555_n N_A_1459_449#_M1008_d 0.00624962f $X=7.435 $Y=2.635
+ $X2=0 $Y2=0
cc_506 N_A_628_123#_c_555_n N_A_1459_449#_c_1172_n 0.0232968f $X=7.435 $Y=2.635
+ $X2=0 $Y2=0
cc_507 N_A_628_123#_c_557_n N_A_1459_449#_c_1172_n 0.0201064f $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_508 N_A_628_123#_c_558_n N_A_1459_449#_c_1172_n 8.80045e-19 $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_509 N_A_628_123#_c_535_n N_A_1459_449#_c_1182_n 0.00135772f $X=7.99 $Y=1.38
+ $X2=0 $Y2=0
cc_510 N_A_628_123#_c_536_n N_A_1459_449#_c_1182_n 0.0171645f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_511 N_A_628_123#_c_537_n N_A_1459_449#_c_1182_n 0.00116306f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_512 N_A_628_123#_c_540_n N_A_1459_449#_c_1182_n 0.0134661f $X=8.155 $Y=0.855
+ $X2=0 $Y2=0
cc_513 N_A_628_123#_c_535_n N_A_1459_449#_c_1163_n 0.0223959f $X=7.99 $Y=1.38
+ $X2=0 $Y2=0
cc_514 N_A_628_123#_c_537_n N_A_1459_449#_c_1163_n 0.00286261f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_515 N_A_628_123#_c_535_n N_A_1459_449#_c_1164_n 0.0129697f $X=7.99 $Y=1.38
+ $X2=0 $Y2=0
cc_516 N_A_628_123#_c_558_n N_A_1459_449#_c_1164_n 2.48753e-19 $X=7.435 $Y=1.92
+ $X2=0 $Y2=0
cc_517 N_A_628_123#_c_539_n N_A_1459_449#_c_1164_n 0.0138878f $X=7.477 $Y=1.755
+ $X2=0 $Y2=0
cc_518 N_A_628_123#_c_535_n N_A_1459_449#_c_1165_n 8.06711e-19 $X=7.99 $Y=1.38
+ $X2=0 $Y2=0
cc_519 N_A_628_123#_c_536_n N_A_1459_449#_c_1165_n 0.0328733f $X=8.155 $Y=1.02
+ $X2=0 $Y2=0
cc_520 N_A_628_123#_c_540_n N_A_1459_449#_c_1165_n 0.00396065f $X=8.155 $Y=0.855
+ $X2=0 $Y2=0
cc_521 N_A_628_123#_M1008_g N_A_1459_449#_c_1194_n 0.00138985f $X=7.22 $Y=2.665
+ $X2=0 $Y2=0
cc_522 N_A_628_123#_c_554_n N_A_1459_449#_c_1194_n 0.0143278f $X=7.35 $Y=2.72
+ $X2=0 $Y2=0
cc_523 N_A_628_123#_c_555_n N_A_1459_449#_c_1194_n 0.0089485f $X=7.435 $Y=2.635
+ $X2=0 $Y2=0
cc_524 N_A_628_123#_c_535_n N_A_1459_449#_c_1168_n 0.01499f $X=7.99 $Y=1.38
+ $X2=0 $Y2=0
cc_525 N_A_628_123#_c_547_n N_VPWR_M1024_s 0.00296017f $X=3.865 $Y=2.47 $X2=0
+ $Y2=0
cc_526 N_A_628_123#_c_579_p N_VPWR_M1024_s 8.52667e-19 $X=4.05 $Y=2.47 $X2=0
+ $Y2=0
cc_527 N_A_628_123#_c_554_n N_VPWR_M1015_d 0.00943699f $X=7.35 $Y=2.72 $X2=0
+ $Y2=0
cc_528 N_A_628_123#_M1024_g N_VPWR_c_1267_n 0.00508913f $X=4.05 $Y=2.725 $X2=0
+ $Y2=0
cc_529 N_A_628_123#_c_546_n N_VPWR_c_1267_n 0.0242041f $X=3.28 $Y=2.6 $X2=0
+ $Y2=0
cc_530 N_A_628_123#_c_547_n N_VPWR_c_1267_n 0.0165959f $X=3.865 $Y=2.47 $X2=0
+ $Y2=0
cc_531 N_A_628_123#_c_577_p N_VPWR_c_1267_n 0.0123064f $X=4.15 $Y=2.895 $X2=0
+ $Y2=0
cc_532 N_A_628_123#_c_551_n N_VPWR_c_1267_n 0.0137976f $X=4.235 $Y=2.98 $X2=0
+ $Y2=0
cc_533 N_A_628_123#_c_579_p N_VPWR_c_1267_n 0.00233451f $X=4.05 $Y=2.47 $X2=0
+ $Y2=0
cc_534 N_A_628_123#_c_546_n N_VPWR_c_1272_n 0.0176268f $X=3.28 $Y=2.6 $X2=0
+ $Y2=0
cc_535 N_A_628_123#_M1024_g N_VPWR_c_1275_n 0.00452629f $X=4.05 $Y=2.725 $X2=0
+ $Y2=0
cc_536 N_A_628_123#_M1029_g N_VPWR_c_1275_n 2.16845e-19 $X=5.71 $Y=2.455 $X2=0
+ $Y2=0
cc_537 N_A_628_123#_c_550_n N_VPWR_c_1275_n 0.0924404f $X=5.76 $Y=2.98 $X2=0
+ $Y2=0
cc_538 N_A_628_123#_c_551_n N_VPWR_c_1275_n 0.0112205f $X=4.235 $Y=2.98 $X2=0
+ $Y2=0
cc_539 N_A_628_123#_c_554_n N_VPWR_c_1275_n 0.00939221f $X=7.35 $Y=2.72 $X2=0
+ $Y2=0
cc_540 N_A_628_123#_c_556_n N_VPWR_c_1275_n 0.0113273f $X=5.845 $Y=2.72 $X2=0
+ $Y2=0
cc_541 N_A_628_123#_M1008_g N_VPWR_c_1276_n 0.00400062f $X=7.22 $Y=2.665 $X2=0
+ $Y2=0
cc_542 N_A_628_123#_c_554_n N_VPWR_c_1276_n 0.0173604f $X=7.35 $Y=2.72 $X2=0
+ $Y2=0
cc_543 N_A_628_123#_M1027_d N_VPWR_c_1264_n 0.00216391f $X=3.14 $Y=2.455 $X2=0
+ $Y2=0
cc_544 N_A_628_123#_M1024_g N_VPWR_c_1264_n 0.00718518f $X=4.05 $Y=2.725 $X2=0
+ $Y2=0
cc_545 N_A_628_123#_M1008_g N_VPWR_c_1264_n 0.00698731f $X=7.22 $Y=2.665 $X2=0
+ $Y2=0
cc_546 N_A_628_123#_c_546_n N_VPWR_c_1264_n 0.01237f $X=3.28 $Y=2.6 $X2=0 $Y2=0
cc_547 N_A_628_123#_c_547_n N_VPWR_c_1264_n 0.00778318f $X=3.865 $Y=2.47 $X2=0
+ $Y2=0
cc_548 N_A_628_123#_c_550_n N_VPWR_c_1264_n 0.0569899f $X=5.76 $Y=2.98 $X2=0
+ $Y2=0
cc_549 N_A_628_123#_c_551_n N_VPWR_c_1264_n 0.00629602f $X=4.235 $Y=2.98 $X2=0
+ $Y2=0
cc_550 N_A_628_123#_c_554_n N_VPWR_c_1264_n 0.0398421f $X=7.35 $Y=2.72 $X2=0
+ $Y2=0
cc_551 N_A_628_123#_c_579_p N_VPWR_c_1264_n 0.00655637f $X=4.05 $Y=2.47 $X2=0
+ $Y2=0
cc_552 N_A_628_123#_c_556_n N_VPWR_c_1264_n 0.00650045f $X=5.845 $Y=2.72 $X2=0
+ $Y2=0
cc_553 N_A_628_123#_c_554_n N_VPWR_c_1281_n 0.0240258f $X=7.35 $Y=2.72 $X2=0
+ $Y2=0
cc_554 N_A_628_123#_c_556_n N_VPWR_c_1281_n 0.00395126f $X=5.845 $Y=2.72 $X2=0
+ $Y2=0
cc_555 N_A_628_123#_c_546_n N_A_319_123#_c_1405_n 6.2717e-19 $X=3.28 $Y=2.6
+ $X2=0 $Y2=0
cc_556 N_A_628_123#_c_546_n N_A_319_123#_c_1432_n 0.00236376f $X=3.28 $Y=2.6
+ $X2=0 $Y2=0
cc_557 N_A_628_123#_c_548_n N_A_319_123#_c_1432_n 0.00149145f $X=3.445 $Y=2.47
+ $X2=0 $Y2=0
cc_558 N_A_628_123#_M1018_g N_A_319_123#_c_1395_n 0.0118316f $X=5.18 $Y=0.835
+ $X2=0 $Y2=0
cc_559 N_A_628_123#_c_547_n N_A_319_123#_c_1400_n 0.0194209f $X=3.865 $Y=2.47
+ $X2=0 $Y2=0
cc_560 N_A_628_123#_c_548_n N_A_319_123#_c_1400_n 0.0258965f $X=3.445 $Y=2.47
+ $X2=0 $Y2=0
cc_561 N_A_628_123#_c_533_n N_A_319_123#_c_1400_n 0.0238952f $X=4.05 $Y=2.385
+ $X2=0 $Y2=0
cc_562 N_A_628_123#_c_550_n N_A_319_123#_c_1400_n 0.0138044f $X=5.76 $Y=2.98
+ $X2=0 $Y2=0
cc_563 N_A_628_123#_c_579_p N_A_319_123#_c_1400_n 0.0214895f $X=4.05 $Y=2.47
+ $X2=0 $Y2=0
cc_564 N_A_628_123#_c_548_n N_A_319_123#_c_1401_n 0.00126481f $X=3.445 $Y=2.47
+ $X2=0 $Y2=0
cc_565 N_A_628_123#_c_550_n N_A_319_123#_c_1469_n 0.00236355f $X=5.76 $Y=2.98
+ $X2=0 $Y2=0
cc_566 N_A_628_123#_c_550_n N_A_319_123#_c_1402_n 0.0135414f $X=5.76 $Y=2.98
+ $X2=0 $Y2=0
cc_567 N_A_628_123#_c_548_n N_A_319_123#_c_1403_n 0.00261736f $X=3.445 $Y=2.47
+ $X2=0 $Y2=0
cc_568 N_A_628_123#_c_553_n A_1157_449# 0.00366202f $X=5.845 $Y=2.635 $X2=-0.19
+ $Y2=-0.245
cc_569 N_A_628_123#_c_554_n A_1157_449# 7.56375e-19 $X=7.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.245
cc_570 N_A_628_123#_c_526_n N_VGND_c_1535_n 0.00459147f $X=3.95 $Y=0.765 $X2=0
+ $Y2=0
cc_571 N_A_628_123#_c_531_n N_VGND_c_1535_n 0.0167147f $X=3.865 $Y=0.85 $X2=0
+ $Y2=0
cc_572 N_A_628_123#_c_532_n N_VGND_c_1535_n 0.00425222f $X=4.05 $Y=0.985 $X2=0
+ $Y2=0
cc_573 N_A_628_123#_c_538_n N_VGND_c_1535_n 8.97164e-19 $X=3.95 $Y=0.93 $X2=0
+ $Y2=0
cc_574 N_A_628_123#_c_540_n N_VGND_c_1537_n 0.00316774f $X=8.155 $Y=0.855 $X2=0
+ $Y2=0
cc_575 N_A_628_123#_c_531_n N_VGND_c_1544_n 0.0080519f $X=3.865 $Y=0.85 $X2=0
+ $Y2=0
cc_576 N_A_628_123#_c_526_n N_VGND_c_1546_n 0.00423618f $X=3.95 $Y=0.765 $X2=0
+ $Y2=0
cc_577 N_A_628_123#_c_532_n N_VGND_c_1546_n 0.00264988f $X=4.05 $Y=0.985 $X2=0
+ $Y2=0
cc_578 N_A_628_123#_c_526_n N_VGND_c_1549_n 0.00839159f $X=3.95 $Y=0.765 $X2=0
+ $Y2=0
cc_579 N_A_628_123#_c_531_n N_VGND_c_1549_n 0.0157476f $X=3.865 $Y=0.85 $X2=0
+ $Y2=0
cc_580 N_A_628_123#_c_532_n N_VGND_c_1549_n 0.00483864f $X=4.05 $Y=0.985 $X2=0
+ $Y2=0
cc_581 N_A_628_123#_c_540_n N_VGND_c_1549_n 0.00458257f $X=8.155 $Y=0.855 $X2=0
+ $Y2=0
cc_582 N_A_823_47#_c_761_n N_A_1201_99#_M1003_d 0.0117744f $X=7.435 $Y=0.47
+ $X2=-0.19 $Y2=-0.245
cc_583 N_A_823_47#_c_759_n N_A_1201_99#_M1030_g 0.00118025f $X=5.63 $Y=0.35
+ $X2=0 $Y2=0
cc_584 N_A_823_47#_c_760_n N_A_1201_99#_M1030_g 0.00501002f $X=5.765 $Y=0.815
+ $X2=0 $Y2=0
cc_585 N_A_823_47#_c_827_p N_A_1201_99#_M1030_g 0.0132669f $X=6.735 $Y=0.9 $X2=0
+ $Y2=0
cc_586 N_A_823_47#_c_766_n N_A_1201_99#_M1030_g 0.0241921f $X=5.63 $Y=0.515
+ $X2=0 $Y2=0
cc_587 N_A_823_47#_c_751_n N_A_1201_99#_c_916_n 0.00194546f $X=7.585 $Y=1.395
+ $X2=0 $Y2=0
cc_588 N_A_823_47#_c_827_p N_A_1201_99#_c_917_n 0.0134661f $X=6.735 $Y=0.9 $X2=0
+ $Y2=0
cc_589 N_A_823_47#_c_831_p N_A_1201_99#_c_917_n 0.00563137f $X=6.82 $Y=0.815
+ $X2=0 $Y2=0
cc_590 N_A_823_47#_c_761_n N_A_1201_99#_c_917_n 0.0139093f $X=7.435 $Y=0.47
+ $X2=0 $Y2=0
cc_591 N_A_823_47#_c_763_n N_A_1201_99#_c_917_n 0.0290675f $X=7.6 $Y=1.03 $X2=0
+ $Y2=0
cc_592 N_A_823_47#_c_767_n N_A_1201_99#_c_917_n 0.00410492f $X=7.585 $Y=0.865
+ $X2=0 $Y2=0
cc_593 N_A_823_47#_c_761_n N_A_1201_99#_c_918_n 0.00244963f $X=7.435 $Y=0.47
+ $X2=0 $Y2=0
cc_594 N_A_823_47#_c_764_n N_A_1201_99#_c_918_n 0.00410492f $X=7.6 $Y=1.03 $X2=0
+ $Y2=0
cc_595 N_A_823_47#_c_753_n N_A_1051_125#_M1013_g 5.99421e-19 $X=7.765 $Y=1.47
+ $X2=0 $Y2=0
cc_596 N_A_823_47#_c_827_p N_A_1051_125#_M1003_g 0.0110071f $X=6.735 $Y=0.9
+ $X2=0 $Y2=0
cc_597 N_A_823_47#_c_831_p N_A_1051_125#_M1003_g 0.00842196f $X=6.82 $Y=0.815
+ $X2=0 $Y2=0
cc_598 N_A_823_47#_c_761_n N_A_1051_125#_M1003_g 0.00490063f $X=7.435 $Y=0.47
+ $X2=0 $Y2=0
cc_599 N_A_823_47#_c_762_n N_A_1051_125#_M1003_g 0.00548744f $X=6.905 $Y=0.47
+ $X2=0 $Y2=0
cc_600 N_A_823_47#_c_763_n N_A_1051_125#_M1003_g 7.2135e-19 $X=7.6 $Y=1.03 $X2=0
+ $Y2=0
cc_601 N_A_823_47#_c_767_n N_A_1051_125#_M1003_g 0.0123302f $X=7.585 $Y=0.865
+ $X2=0 $Y2=0
cc_602 N_A_823_47#_c_758_n N_A_1051_125#_c_983_n 0.0161328f $X=5.68 $Y=0.375
+ $X2=0 $Y2=0
cc_603 N_A_823_47#_c_759_n N_A_1051_125#_c_983_n 9.62037e-19 $X=5.63 $Y=0.35
+ $X2=0 $Y2=0
cc_604 N_A_823_47#_c_766_n N_A_1051_125#_c_983_n 0.00354606f $X=5.63 $Y=0.515
+ $X2=0 $Y2=0
cc_605 N_A_823_47#_c_768_n N_A_1051_125#_c_990_n 0.011239f $X=5.205 $Y=2.06
+ $X2=0 $Y2=0
cc_606 N_A_823_47#_c_768_n N_A_1051_125#_c_991_n 0.00301071f $X=5.205 $Y=2.06
+ $X2=0 $Y2=0
cc_607 N_A_823_47#_c_770_n N_A_1051_125#_c_991_n 0.00838538f $X=5.28 $Y=2.135
+ $X2=0 $Y2=0
cc_608 N_A_823_47#_c_759_n N_A_1051_125#_c_984_n 8.60196e-19 $X=5.63 $Y=0.35
+ $X2=0 $Y2=0
cc_609 N_A_823_47#_c_827_p N_A_1051_125#_c_984_n 0.0495162f $X=6.735 $Y=0.9
+ $X2=0 $Y2=0
cc_610 N_A_823_47#_c_852_p N_A_1051_125#_c_984_n 0.0105534f $X=5.85 $Y=0.9 $X2=0
+ $Y2=0
cc_611 N_A_823_47#_c_766_n N_A_1051_125#_c_984_n 0.0040278f $X=5.63 $Y=0.515
+ $X2=0 $Y2=0
cc_612 N_A_823_47#_c_827_p N_A_1051_125#_c_986_n 0.00968339f $X=6.735 $Y=0.9
+ $X2=0 $Y2=0
cc_613 N_A_823_47#_c_751_n N_A_1051_125#_c_987_n 0.0123302f $X=7.585 $Y=1.395
+ $X2=0 $Y2=0
cc_614 N_A_823_47#_c_827_p N_A_1051_125#_c_987_n 0.00236732f $X=6.735 $Y=0.9
+ $X2=0 $Y2=0
cc_615 N_A_823_47#_M1021_g N_A_1657_383#_M1022_g 0.0258528f $X=8 $Y=2.685 $X2=0
+ $Y2=0
cc_616 N_A_823_47#_c_752_n N_A_1657_383#_M1026_g 0.0121813f $X=7.925 $Y=1.47
+ $X2=0 $Y2=0
cc_617 N_A_823_47#_M1021_g N_A_1657_383#_c_1081_n 6.2387e-19 $X=8 $Y=2.685 $X2=0
+ $Y2=0
cc_618 N_A_823_47#_M1021_g N_A_1657_383#_c_1082_n 0.0205211f $X=8 $Y=2.685 $X2=0
+ $Y2=0
cc_619 N_A_823_47#_c_761_n N_A_1459_449#_M1014_d 0.00387183f $X=7.435 $Y=0.47
+ $X2=-0.19 $Y2=-0.245
cc_620 N_A_823_47#_c_763_n N_A_1459_449#_M1014_d 0.00251037f $X=7.6 $Y=1.03
+ $X2=-0.19 $Y2=-0.245
cc_621 N_A_823_47#_M1021_g N_A_1459_449#_c_1172_n 0.0195419f $X=8 $Y=2.685 $X2=0
+ $Y2=0
cc_622 N_A_823_47#_c_761_n N_A_1459_449#_c_1182_n 0.0146248f $X=7.435 $Y=0.47
+ $X2=0 $Y2=0
cc_623 N_A_823_47#_c_763_n N_A_1459_449#_c_1182_n 0.00963175f $X=7.6 $Y=1.03
+ $X2=0 $Y2=0
cc_624 N_A_823_47#_c_767_n N_A_1459_449#_c_1182_n 0.00177107f $X=7.585 $Y=0.865
+ $X2=0 $Y2=0
cc_625 N_A_823_47#_M1021_g N_A_1459_449#_c_1163_n 0.0115334f $X=8 $Y=2.685 $X2=0
+ $Y2=0
cc_626 N_A_823_47#_c_752_n N_A_1459_449#_c_1164_n 0.0030555f $X=7.925 $Y=1.47
+ $X2=0 $Y2=0
cc_627 N_A_823_47#_M1021_g N_A_1459_449#_c_1164_n 0.00330494f $X=8 $Y=2.685
+ $X2=0 $Y2=0
cc_628 N_A_823_47#_c_763_n N_A_1459_449#_c_1165_n 0.0052781f $X=7.6 $Y=1.03
+ $X2=0 $Y2=0
cc_629 N_A_823_47#_M1021_g N_A_1459_449#_c_1194_n 0.00690222f $X=8 $Y=2.685
+ $X2=0 $Y2=0
cc_630 N_A_823_47#_c_751_n N_A_1459_449#_c_1168_n 2.71776e-19 $X=7.585 $Y=1.395
+ $X2=0 $Y2=0
cc_631 N_A_823_47#_c_752_n N_A_1459_449#_c_1168_n 0.00460491f $X=7.925 $Y=1.47
+ $X2=0 $Y2=0
cc_632 N_A_823_47#_M1021_g N_VPWR_c_1276_n 0.00503195f $X=8 $Y=2.685 $X2=0 $Y2=0
cc_633 N_A_823_47#_M1021_g N_VPWR_c_1264_n 0.00525227f $X=8 $Y=2.685 $X2=0 $Y2=0
cc_634 N_A_823_47#_c_768_n N_A_319_123#_c_1395_n 0.0139181f $X=5.205 $Y=2.06
+ $X2=0 $Y2=0
cc_635 N_A_823_47#_c_770_n N_A_319_123#_c_1395_n 0.00170569f $X=5.28 $Y=2.135
+ $X2=0 $Y2=0
cc_636 N_A_823_47#_c_756_n N_A_319_123#_c_1395_n 0.0902416f $X=4.5 $Y=1.63 $X2=0
+ $Y2=0
cc_637 N_A_823_47#_c_757_n N_A_319_123#_c_1395_n 0.00797576f $X=4.5 $Y=1.63
+ $X2=0 $Y2=0
cc_638 N_A_823_47#_c_756_n N_A_319_123#_c_1396_n 0.0263381f $X=4.5 $Y=1.63 $X2=0
+ $Y2=0
cc_639 N_A_823_47#_c_758_n N_A_319_123#_c_1396_n 0.0222308f $X=5.68 $Y=0.375
+ $X2=0 $Y2=0
cc_640 N_A_823_47#_M1024_d N_A_319_123#_c_1400_n 0.00216422f $X=4.125 $Y=2.405
+ $X2=0 $Y2=0
cc_641 N_A_823_47#_c_769_n N_A_319_123#_c_1400_n 0.00591425f $X=4.665 $Y=2.06
+ $X2=0 $Y2=0
cc_642 N_A_823_47#_c_756_n N_A_319_123#_c_1400_n 0.0135484f $X=4.5 $Y=1.63 $X2=0
+ $Y2=0
cc_643 N_A_823_47#_c_768_n N_A_319_123#_c_1469_n 3.34556e-19 $X=5.205 $Y=2.06
+ $X2=0 $Y2=0
cc_644 N_A_823_47#_c_756_n N_A_319_123#_c_1469_n 4.9596e-19 $X=4.5 $Y=1.63 $X2=0
+ $Y2=0
cc_645 N_A_823_47#_c_768_n N_A_319_123#_c_1402_n 0.00969419f $X=5.205 $Y=2.06
+ $X2=0 $Y2=0
cc_646 N_A_823_47#_c_770_n N_A_319_123#_c_1402_n 7.55263e-19 $X=5.28 $Y=2.135
+ $X2=0 $Y2=0
cc_647 N_A_823_47#_c_756_n N_A_319_123#_c_1402_n 0.024803f $X=4.5 $Y=1.63 $X2=0
+ $Y2=0
cc_648 N_A_823_47#_c_827_p N_VGND_M1030_d 0.0151014f $X=6.735 $Y=0.9 $X2=0 $Y2=0
cc_649 N_A_823_47#_c_758_n N_VGND_c_1536_n 0.0112365f $X=5.68 $Y=0.375 $X2=0
+ $Y2=0
cc_650 N_A_823_47#_c_759_n N_VGND_c_1536_n 0.00309533f $X=5.63 $Y=0.35 $X2=0
+ $Y2=0
cc_651 N_A_823_47#_c_760_n N_VGND_c_1536_n 0.00680473f $X=5.765 $Y=0.815 $X2=0
+ $Y2=0
cc_652 N_A_823_47#_c_827_p N_VGND_c_1536_n 0.0249648f $X=6.735 $Y=0.9 $X2=0
+ $Y2=0
cc_653 N_A_823_47#_c_762_n N_VGND_c_1536_n 0.00744311f $X=6.905 $Y=0.47 $X2=0
+ $Y2=0
cc_654 N_A_823_47#_c_761_n N_VGND_c_1537_n 0.0287785f $X=7.435 $Y=0.47 $X2=0
+ $Y2=0
cc_655 N_A_823_47#_c_762_n N_VGND_c_1537_n 0.00625485f $X=6.905 $Y=0.47 $X2=0
+ $Y2=0
cc_656 N_A_823_47#_c_767_n N_VGND_c_1537_n 0.00322662f $X=7.585 $Y=0.865 $X2=0
+ $Y2=0
cc_657 N_A_823_47#_c_755_n N_VGND_c_1546_n 0.0174714f $X=4.405 $Y=0.375 $X2=0
+ $Y2=0
cc_658 N_A_823_47#_c_758_n N_VGND_c_1546_n 0.0773915f $X=5.68 $Y=0.375 $X2=0
+ $Y2=0
cc_659 N_A_823_47#_c_759_n N_VGND_c_1546_n 0.0065119f $X=5.63 $Y=0.35 $X2=0
+ $Y2=0
cc_660 N_A_823_47#_c_765_n N_VGND_c_1546_n 0.0128106f $X=4.5 $Y=0.375 $X2=0
+ $Y2=0
cc_661 N_A_823_47#_M1004_d N_VGND_c_1549_n 0.00215439f $X=4.115 $Y=0.235 $X2=0
+ $Y2=0
cc_662 N_A_823_47#_c_755_n N_VGND_c_1549_n 0.0116511f $X=4.405 $Y=0.375 $X2=0
+ $Y2=0
cc_663 N_A_823_47#_c_758_n N_VGND_c_1549_n 0.0458489f $X=5.68 $Y=0.375 $X2=0
+ $Y2=0
cc_664 N_A_823_47#_c_759_n N_VGND_c_1549_n 0.010104f $X=5.63 $Y=0.35 $X2=0 $Y2=0
cc_665 N_A_823_47#_c_827_p N_VGND_c_1549_n 0.0202513f $X=6.735 $Y=0.9 $X2=0
+ $Y2=0
cc_666 N_A_823_47#_c_761_n N_VGND_c_1549_n 0.0294499f $X=7.435 $Y=0.47 $X2=0
+ $Y2=0
cc_667 N_A_823_47#_c_762_n N_VGND_c_1549_n 0.00601145f $X=6.905 $Y=0.47 $X2=0
+ $Y2=0
cc_668 N_A_823_47#_c_765_n N_VGND_c_1549_n 0.0073517f $X=4.5 $Y=0.375 $X2=0
+ $Y2=0
cc_669 N_A_823_47#_c_767_n N_VGND_c_1549_n 0.00518872f $X=7.585 $Y=0.865 $X2=0
+ $Y2=0
cc_670 N_A_823_47#_c_760_n A_1137_125# 0.00217171f $X=5.765 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_671 N_A_823_47#_c_827_p A_1137_125# 0.00299188f $X=6.735 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_672 N_A_823_47#_c_852_p A_1137_125# 0.00116918f $X=5.85 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_673 N_A_1201_99#_M1030_g N_A_1051_125#_M1013_g 0.00481978f $X=6.08 $Y=0.835
+ $X2=0 $Y2=0
cc_674 N_A_1201_99#_M1015_g N_A_1051_125#_M1013_g 0.0140877f $X=6.08 $Y=2.455
+ $X2=0 $Y2=0
cc_675 N_A_1201_99#_c_921_n N_A_1051_125#_M1013_g 0.0371874f $X=7 $Y=2.075 $X2=0
+ $Y2=0
cc_676 N_A_1201_99#_c_922_n N_A_1051_125#_M1013_g 0.01091f $X=6.195 $Y=1.85
+ $X2=0 $Y2=0
cc_677 N_A_1201_99#_c_916_n N_A_1051_125#_M1013_g 0.00592433f $X=7.085 $Y=1.685
+ $X2=0 $Y2=0
cc_678 N_A_1201_99#_M1030_g N_A_1051_125#_M1003_g 0.0105442f $X=6.08 $Y=0.835
+ $X2=0 $Y2=0
cc_679 N_A_1201_99#_c_917_n N_A_1051_125#_M1003_g 0.00626211f $X=7.16 $Y=0.9
+ $X2=0 $Y2=0
cc_680 N_A_1201_99#_c_918_n N_A_1051_125#_M1003_g 0.00192541f $X=7.132 $Y=1.335
+ $X2=0 $Y2=0
cc_681 N_A_1201_99#_M1030_g N_A_1051_125#_c_984_n 0.0165299f $X=6.08 $Y=0.835
+ $X2=0 $Y2=0
cc_682 N_A_1201_99#_c_921_n N_A_1051_125#_c_984_n 0.026884f $X=7 $Y=2.075 $X2=0
+ $Y2=0
cc_683 N_A_1201_99#_c_922_n N_A_1051_125#_c_984_n 0.00407103f $X=6.195 $Y=1.85
+ $X2=0 $Y2=0
cc_684 N_A_1201_99#_M1030_g N_A_1051_125#_c_986_n 8.87573e-19 $X=6.08 $Y=0.835
+ $X2=0 $Y2=0
cc_685 N_A_1201_99#_c_921_n N_A_1051_125#_c_986_n 0.0131032f $X=7 $Y=2.075 $X2=0
+ $Y2=0
cc_686 N_A_1201_99#_c_918_n N_A_1051_125#_c_986_n 0.0229744f $X=7.132 $Y=1.335
+ $X2=0 $Y2=0
cc_687 N_A_1201_99#_M1030_g N_A_1051_125#_c_987_n 0.00971833f $X=6.08 $Y=0.835
+ $X2=0 $Y2=0
cc_688 N_A_1201_99#_c_921_n N_A_1051_125#_c_987_n 0.00594134f $X=7 $Y=2.075
+ $X2=0 $Y2=0
cc_689 N_A_1201_99#_c_916_n N_A_1051_125#_c_987_n 0.00192541f $X=7.085 $Y=1.685
+ $X2=0 $Y2=0
cc_690 N_A_1201_99#_c_921_n N_VPWR_M1015_d 0.00738417f $X=7 $Y=2.075 $X2=0 $Y2=0
cc_691 N_A_1201_99#_M1015_g N_VPWR_c_1275_n 6.65218e-19 $X=6.08 $Y=2.455 $X2=0
+ $Y2=0
cc_692 N_A_1201_99#_M1013_d N_VPWR_c_1264_n 0.00283464f $X=6.865 $Y=2.245 $X2=0
+ $Y2=0
cc_693 N_A_1201_99#_M1030_g N_VGND_c_1536_n 0.00199781f $X=6.08 $Y=0.835 $X2=0
+ $Y2=0
cc_694 N_A_1201_99#_M1030_g N_VGND_c_1546_n 0.00415323f $X=6.08 $Y=0.835 $X2=0
+ $Y2=0
cc_695 N_A_1201_99#_M1030_g N_VGND_c_1549_n 0.00469432f $X=6.08 $Y=0.835 $X2=0
+ $Y2=0
cc_696 N_A_1051_125#_M1013_g N_VPWR_c_1276_n 0.00400062f $X=6.79 $Y=2.665 $X2=0
+ $Y2=0
cc_697 N_A_1051_125#_M1013_g N_VPWR_c_1264_n 0.00686705f $X=6.79 $Y=2.665 $X2=0
+ $Y2=0
cc_698 N_A_1051_125#_M1013_g N_VPWR_c_1281_n 0.00659856f $X=6.79 $Y=2.665 $X2=0
+ $Y2=0
cc_699 N_A_1051_125#_c_982_n N_A_319_123#_c_1395_n 0.0366306f $X=5.2 $Y=1.875
+ $X2=0 $Y2=0
cc_700 N_A_1051_125#_c_983_n N_A_319_123#_c_1395_n 0.00740707f $X=5.395 $Y=0.82
+ $X2=0 $Y2=0
cc_701 N_A_1051_125#_c_990_n N_A_319_123#_c_1395_n 0.0127496f $X=5.465 $Y=2.045
+ $X2=0 $Y2=0
cc_702 N_A_1051_125#_c_991_n N_A_319_123#_c_1395_n 0.00656779f $X=5.495 $Y=2.45
+ $X2=0 $Y2=0
cc_703 N_A_1051_125#_c_985_n N_A_319_123#_c_1395_n 0.0130074f $X=5.312 $Y=1.26
+ $X2=0 $Y2=0
cc_704 N_A_1051_125#_c_990_n N_A_319_123#_c_1469_n 9.11993e-19 $X=5.465 $Y=2.045
+ $X2=0 $Y2=0
cc_705 N_A_1051_125#_c_991_n N_A_319_123#_c_1469_n 0.00728872f $X=5.495 $Y=2.45
+ $X2=0 $Y2=0
cc_706 N_A_1051_125#_c_990_n N_A_319_123#_c_1402_n 0.00366418f $X=5.465 $Y=2.045
+ $X2=0 $Y2=0
cc_707 N_A_1051_125#_c_991_n N_A_319_123#_c_1402_n 0.0152181f $X=5.495 $Y=2.45
+ $X2=0 $Y2=0
cc_708 N_A_1051_125#_M1003_g N_VGND_c_1536_n 0.00509716f $X=6.86 $Y=0.725 $X2=0
+ $Y2=0
cc_709 N_A_1051_125#_M1003_g N_VGND_c_1537_n 0.00395727f $X=6.86 $Y=0.725 $X2=0
+ $Y2=0
cc_710 N_A_1051_125#_M1003_g N_VGND_c_1549_n 0.00534666f $X=6.86 $Y=0.725 $X2=0
+ $Y2=0
cc_711 N_A_1657_383#_M1026_g N_A_1459_449#_M1000_g 0.0196057f $X=8.605 $Y=0.535
+ $X2=0 $Y2=0
cc_712 N_A_1657_383#_c_1072_n N_A_1459_449#_M1000_g 7.68644e-19 $X=9.345 $Y=0.48
+ $X2=0 $Y2=0
cc_713 N_A_1657_383#_c_1073_n N_A_1459_449#_M1000_g 0.00796494f $X=9.485
+ $Y=1.415 $X2=0 $Y2=0
cc_714 N_A_1657_383#_M1022_g N_A_1459_449#_M1001_g 0.00803367f $X=8.51 $Y=2.685
+ $X2=0 $Y2=0
cc_715 N_A_1657_383#_M1026_g N_A_1459_449#_M1001_g 0.0117108f $X=8.605 $Y=0.535
+ $X2=0 $Y2=0
cc_716 N_A_1657_383#_c_1081_n N_A_1459_449#_M1001_g 0.0148412f $X=9.265 $Y=2.08
+ $X2=0 $Y2=0
cc_717 N_A_1657_383#_c_1083_n N_A_1459_449#_M1001_g 0.00330324f $X=9.35 $Y=2.2
+ $X2=0 $Y2=0
cc_718 N_A_1657_383#_c_1074_n N_A_1459_449#_M1001_g 0.00298203f $X=9.485
+ $Y=1.985 $X2=0 $Y2=0
cc_719 N_A_1657_383#_c_1074_n N_A_1459_449#_c_1162_n 0.00109322f $X=9.485
+ $Y=1.985 $X2=0 $Y2=0
cc_720 N_A_1657_383#_c_1076_n N_A_1459_449#_c_1162_n 7.94271e-19 $X=9.615 $Y=1.5
+ $X2=0 $Y2=0
cc_721 N_A_1657_383#_c_1081_n N_A_1459_449#_c_1171_n 0.0051471f $X=9.265 $Y=2.08
+ $X2=0 $Y2=0
cc_722 N_A_1657_383#_c_1074_n N_A_1459_449#_c_1171_n 0.00301019f $X=9.485
+ $Y=1.985 $X2=0 $Y2=0
cc_723 N_A_1657_383#_M1022_g N_A_1459_449#_c_1172_n 0.0012893f $X=8.51 $Y=2.685
+ $X2=0 $Y2=0
cc_724 N_A_1657_383#_M1026_g N_A_1459_449#_c_1172_n 4.50336e-19 $X=8.605
+ $Y=0.535 $X2=0 $Y2=0
cc_725 N_A_1657_383#_c_1081_n N_A_1459_449#_c_1172_n 0.00839867f $X=9.265
+ $Y=2.08 $X2=0 $Y2=0
cc_726 N_A_1657_383#_c_1082_n N_A_1459_449#_c_1172_n 9.9492e-19 $X=8.45 $Y=2.08
+ $X2=0 $Y2=0
cc_727 N_A_1657_383#_M1026_g N_A_1459_449#_c_1182_n 0.00815958f $X=8.605
+ $Y=0.535 $X2=0 $Y2=0
cc_728 N_A_1657_383#_c_1081_n N_A_1459_449#_c_1163_n 0.00969624f $X=9.265
+ $Y=2.08 $X2=0 $Y2=0
cc_729 N_A_1657_383#_c_1082_n N_A_1459_449#_c_1163_n 0.00328529f $X=8.45 $Y=2.08
+ $X2=0 $Y2=0
cc_730 N_A_1657_383#_M1026_g N_A_1459_449#_c_1165_n 0.015233f $X=8.605 $Y=0.535
+ $X2=0 $Y2=0
cc_731 N_A_1657_383#_c_1075_n N_A_1459_449#_c_1165_n 2.70793e-19 $X=9.405
+ $Y=0.985 $X2=0 $Y2=0
cc_732 N_A_1657_383#_M1026_g N_A_1459_449#_c_1166_n 0.0145542f $X=8.605 $Y=0.535
+ $X2=0 $Y2=0
cc_733 N_A_1657_383#_c_1081_n N_A_1459_449#_c_1166_n 0.0493457f $X=9.265 $Y=2.08
+ $X2=0 $Y2=0
cc_734 N_A_1657_383#_c_1073_n N_A_1459_449#_c_1166_n 0.00829992f $X=9.485
+ $Y=1.415 $X2=0 $Y2=0
cc_735 N_A_1657_383#_c_1074_n N_A_1459_449#_c_1166_n 0.0128908f $X=9.485
+ $Y=1.985 $X2=0 $Y2=0
cc_736 N_A_1657_383#_c_1076_n N_A_1459_449#_c_1166_n 0.018604f $X=9.615 $Y=1.5
+ $X2=0 $Y2=0
cc_737 N_A_1657_383#_c_1077_n N_A_1459_449#_c_1166_n 3.70993e-19 $X=9.615
+ $Y=1.41 $X2=0 $Y2=0
cc_738 N_A_1657_383#_M1026_g N_A_1459_449#_c_1167_n 0.0436695f $X=8.605 $Y=0.535
+ $X2=0 $Y2=0
cc_739 N_A_1657_383#_c_1073_n N_A_1459_449#_c_1167_n 0.00345352f $X=9.485
+ $Y=1.415 $X2=0 $Y2=0
cc_740 N_A_1657_383#_c_1077_n N_A_1459_449#_c_1167_n 0.0191506f $X=9.615 $Y=1.41
+ $X2=0 $Y2=0
cc_741 N_A_1657_383#_M1022_g N_A_1459_449#_c_1194_n 0.00156293f $X=8.51 $Y=2.685
+ $X2=0 $Y2=0
cc_742 N_A_1657_383#_M1026_g N_A_1459_449#_c_1168_n 0.0105145f $X=8.605 $Y=0.535
+ $X2=0 $Y2=0
cc_743 N_A_1657_383#_c_1081_n N_A_1459_449#_c_1168_n 0.0135448f $X=9.265 $Y=2.08
+ $X2=0 $Y2=0
cc_744 N_A_1657_383#_c_1082_n N_A_1459_449#_c_1168_n 0.00319413f $X=8.45 $Y=2.08
+ $X2=0 $Y2=0
cc_745 N_A_1657_383#_c_1081_n N_VPWR_M1022_d 0.00256375f $X=9.265 $Y=2.08 $X2=0
+ $Y2=0
cc_746 N_A_1657_383#_M1022_g N_VPWR_c_1268_n 0.0173169f $X=8.51 $Y=2.685 $X2=0
+ $Y2=0
cc_747 N_A_1657_383#_c_1081_n N_VPWR_c_1268_n 0.0221068f $X=9.265 $Y=2.08 $X2=0
+ $Y2=0
cc_748 N_A_1657_383#_c_1083_n N_VPWR_c_1268_n 0.0208031f $X=9.35 $Y=2.2 $X2=0
+ $Y2=0
cc_749 N_A_1657_383#_c_1068_n N_VPWR_c_1269_n 0.00402558f $X=10.01 $Y=1.41 $X2=0
+ $Y2=0
cc_750 N_A_1657_383#_M1005_g N_VPWR_c_1269_n 0.0088297f $X=10.085 $Y=2.465 $X2=0
+ $Y2=0
cc_751 N_A_1657_383#_c_1083_n N_VPWR_c_1269_n 0.0592646f $X=9.35 $Y=2.2 $X2=0
+ $Y2=0
cc_752 N_A_1657_383#_c_1074_n N_VPWR_c_1269_n 0.0130859f $X=9.485 $Y=1.985 $X2=0
+ $Y2=0
cc_753 N_A_1657_383#_c_1085_n N_VPWR_c_1269_n 0.0164092f $X=9.417 $Y=2.08 $X2=0
+ $Y2=0
cc_754 N_A_1657_383#_c_1076_n N_VPWR_c_1269_n 0.00320974f $X=9.615 $Y=1.5 $X2=0
+ $Y2=0
cc_755 N_A_1657_383#_c_1077_n N_VPWR_c_1269_n 9.30675e-19 $X=9.615 $Y=1.41 $X2=0
+ $Y2=0
cc_756 N_A_1657_383#_M1022_g N_VPWR_c_1276_n 0.00530923f $X=8.51 $Y=2.685 $X2=0
+ $Y2=0
cc_757 N_A_1657_383#_c_1083_n N_VPWR_c_1277_n 0.0105393f $X=9.35 $Y=2.2 $X2=0
+ $Y2=0
cc_758 N_A_1657_383#_M1005_g N_VPWR_c_1278_n 0.00585385f $X=10.085 $Y=2.465
+ $X2=0 $Y2=0
cc_759 N_A_1657_383#_M1022_g N_VPWR_c_1264_n 0.00525227f $X=8.51 $Y=2.685 $X2=0
+ $Y2=0
cc_760 N_A_1657_383#_M1005_g N_VPWR_c_1264_n 0.012823f $X=10.085 $Y=2.465 $X2=0
+ $Y2=0
cc_761 N_A_1657_383#_c_1083_n N_VPWR_c_1264_n 0.0107063f $X=9.35 $Y=2.2 $X2=0
+ $Y2=0
cc_762 N_A_1657_383#_c_1069_n Q 0.0247571f $X=10.085 $Y=1.335 $X2=0 $Y2=0
cc_763 N_A_1657_383#_c_1073_n Q 0.00500588f $X=9.485 $Y=1.415 $X2=0 $Y2=0
cc_764 N_A_1657_383#_c_1074_n Q 0.0052251f $X=9.485 $Y=1.985 $X2=0 $Y2=0
cc_765 N_A_1657_383#_c_1076_n Q 0.00921212f $X=9.615 $Y=1.5 $X2=0 $Y2=0
cc_766 N_A_1657_383#_M1026_g N_VGND_c_1537_n 0.00426374f $X=8.605 $Y=0.535 $X2=0
+ $Y2=0
cc_767 N_A_1657_383#_M1026_g N_VGND_c_1538_n 0.00823385f $X=8.605 $Y=0.535 $X2=0
+ $Y2=0
cc_768 N_A_1657_383#_c_1072_n N_VGND_c_1538_n 0.00120849f $X=9.345 $Y=0.48 $X2=0
+ $Y2=0
cc_769 N_A_1657_383#_c_1069_n N_VGND_c_1539_n 0.0204601f $X=10.085 $Y=1.335
+ $X2=0 $Y2=0
cc_770 N_A_1657_383#_c_1072_n N_VGND_c_1539_n 0.0754745f $X=9.345 $Y=0.48 $X2=0
+ $Y2=0
cc_771 N_A_1657_383#_c_1076_n N_VGND_c_1539_n 0.00320947f $X=9.615 $Y=1.5 $X2=0
+ $Y2=0
cc_772 N_A_1657_383#_c_1077_n N_VGND_c_1539_n 0.00813228f $X=9.615 $Y=1.41 $X2=0
+ $Y2=0
cc_773 N_A_1657_383#_c_1072_n N_VGND_c_1547_n 0.0170085f $X=9.345 $Y=0.48 $X2=0
+ $Y2=0
cc_774 N_A_1657_383#_c_1069_n N_VGND_c_1548_n 0.00509087f $X=10.085 $Y=1.335
+ $X2=0 $Y2=0
cc_775 N_A_1657_383#_M1026_g N_VGND_c_1549_n 0.00773363f $X=8.605 $Y=0.535 $X2=0
+ $Y2=0
cc_776 N_A_1657_383#_c_1069_n N_VGND_c_1549_n 0.00490561f $X=10.085 $Y=1.335
+ $X2=0 $Y2=0
cc_777 N_A_1657_383#_c_1072_n N_VGND_c_1549_n 0.0123602f $X=9.345 $Y=0.48 $X2=0
+ $Y2=0
cc_778 N_A_1459_449#_M1001_g N_VPWR_c_1268_n 0.0113938f $X=9.135 $Y=2.475 $X2=0
+ $Y2=0
cc_779 N_A_1459_449#_M1001_g N_VPWR_c_1269_n 0.00320417f $X=9.135 $Y=2.475 $X2=0
+ $Y2=0
cc_780 N_A_1459_449#_c_1194_n N_VPWR_c_1276_n 0.0062685f $X=7.87 $Y=2.68 $X2=0
+ $Y2=0
cc_781 N_A_1459_449#_M1001_g N_VPWR_c_1277_n 0.00441186f $X=9.135 $Y=2.475 $X2=0
+ $Y2=0
cc_782 N_A_1459_449#_M1008_d N_VPWR_c_1264_n 0.0033464f $X=7.295 $Y=2.245 $X2=0
+ $Y2=0
cc_783 N_A_1459_449#_M1001_g N_VPWR_c_1264_n 0.0044119f $X=9.135 $Y=2.475 $X2=0
+ $Y2=0
cc_784 N_A_1459_449#_c_1194_n N_VPWR_c_1264_n 0.0086577f $X=7.87 $Y=2.68 $X2=0
+ $Y2=0
cc_785 N_A_1459_449#_c_1182_n N_VGND_c_1537_n 0.0237609f $X=8.42 $Y=0.51 $X2=0
+ $Y2=0
cc_786 N_A_1459_449#_M1000_g N_VGND_c_1538_n 0.00318802f $X=9.13 $Y=0.645 $X2=0
+ $Y2=0
cc_787 N_A_1459_449#_c_1182_n N_VGND_c_1538_n 0.0214657f $X=8.42 $Y=0.51 $X2=0
+ $Y2=0
cc_788 N_A_1459_449#_c_1165_n N_VGND_c_1538_n 0.0175531f $X=8.505 $Y=1.305 $X2=0
+ $Y2=0
cc_789 N_A_1459_449#_c_1166_n N_VGND_c_1538_n 0.0113863f $X=9.055 $Y=1.39 $X2=0
+ $Y2=0
cc_790 N_A_1459_449#_c_1167_n N_VGND_c_1538_n 0.00343229f $X=9.055 $Y=1.39 $X2=0
+ $Y2=0
cc_791 N_A_1459_449#_M1000_g N_VGND_c_1539_n 0.00362914f $X=9.13 $Y=0.645 $X2=0
+ $Y2=0
cc_792 N_A_1459_449#_M1000_g N_VGND_c_1547_n 0.00499542f $X=9.13 $Y=0.645 $X2=0
+ $Y2=0
cc_793 N_A_1459_449#_M1000_g N_VGND_c_1549_n 0.0103534f $X=9.13 $Y=0.645 $X2=0
+ $Y2=0
cc_794 N_A_1459_449#_c_1182_n N_VGND_c_1549_n 0.0224537f $X=8.42 $Y=0.51 $X2=0
+ $Y2=0
cc_795 N_A_1459_449#_c_1182_n A_1664_65# 0.00284253f $X=8.42 $Y=0.51 $X2=-0.19
+ $Y2=-0.245
cc_796 N_A_1459_449#_c_1165_n A_1664_65# 9.86239e-19 $X=8.505 $Y=1.305 $X2=-0.19
+ $Y2=-0.245
cc_797 N_VPWR_c_1264_n A_283_491# 0.00314438f $X=10.32 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_798 N_VPWR_c_1264_n N_A_319_123#_M1028_d 0.00236474f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_799 N_VPWR_c_1266_n N_A_319_123#_c_1405_n 0.0245556f $X=2.84 $Y=2.825 $X2=0
+ $Y2=0
cc_800 N_VPWR_c_1270_n N_A_319_123#_c_1405_n 0.0288157f $X=2.755 $Y=3.33 $X2=0
+ $Y2=0
cc_801 N_VPWR_c_1264_n N_A_319_123#_c_1405_n 0.0288908f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_802 N_VPWR_c_1266_n N_A_319_123#_c_1397_n 0.00347353f $X=2.84 $Y=2.825 $X2=0
+ $Y2=0
cc_803 N_VPWR_M1007_d N_A_319_123#_c_1400_n 0.00301601f $X=2.675 $Y=2.455 $X2=0
+ $Y2=0
cc_804 N_VPWR_c_1266_n N_A_319_123#_c_1400_n 0.00489105f $X=2.84 $Y=2.825 $X2=0
+ $Y2=0
cc_805 N_VPWR_c_1267_n N_A_319_123#_c_1400_n 0.00182959f $X=3.8 $Y=2.89 $X2=0
+ $Y2=0
cc_806 N_VPWR_M1007_d N_A_319_123#_c_1401_n 0.00392321f $X=2.675 $Y=2.455 $X2=0
+ $Y2=0
cc_807 N_VPWR_c_1266_n N_A_319_123#_c_1401_n 0.00101567f $X=2.84 $Y=2.825 $X2=0
+ $Y2=0
cc_808 N_VPWR_c_1264_n N_A_319_123#_c_1403_n 0.00316001f $X=10.32 $Y=3.33 $X2=0
+ $Y2=0
cc_809 N_VPWR_c_1264_n A_441_491# 0.00270181f $X=10.32 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_810 N_VPWR_c_1264_n N_Q_M1005_d 0.00336915f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_811 N_VPWR_c_1269_n Q 0.0012665f $X=9.87 $Y=1.98 $X2=0 $Y2=0
cc_812 N_VPWR_c_1278_n Q 0.0181659f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_813 N_VPWR_c_1264_n Q 0.0104192f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_814 N_VPWR_c_1269_n N_VGND_c_1539_n 0.00773234f $X=9.87 $Y=1.98 $X2=0 $Y2=0
cc_815 N_A_319_123#_c_1405_n A_441_491# 0.00728855f $X=2.415 $Y=2.805 $X2=-0.19
+ $Y2=-0.245
cc_816 N_A_319_123#_c_1432_n A_441_491# 0.0017662f $X=2.5 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_817 N_A_319_123#_c_1403_n A_441_491# 3.80108e-19 $X=2.57 $Y=2.12 $X2=-0.19
+ $Y2=-0.245
cc_818 N_A_319_123#_c_1391_n N_VGND_c_1534_n 0.00810818f $X=2.03 $Y=0.85 $X2=0
+ $Y2=0
cc_819 N_A_319_123#_c_1392_n N_VGND_c_1534_n 0.0173048f $X=2.905 $Y=1.24 $X2=0
+ $Y2=0
cc_820 N_A_319_123#_c_1391_n N_VGND_c_1542_n 0.00375018f $X=2.03 $Y=0.85 $X2=0
+ $Y2=0
cc_821 N_A_319_123#_c_1391_n N_VGND_c_1549_n 0.00620257f $X=2.03 $Y=0.85 $X2=0
+ $Y2=0
cc_822 Q N_VGND_c_1539_n 0.0338201f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_823 Q N_VGND_c_1548_n 0.0112788f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_824 Q N_VGND_c_1549_n 0.00980826f $X=10.235 $Y=0.47 $X2=0 $Y2=0
