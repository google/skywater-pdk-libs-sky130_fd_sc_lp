* File: sky130_fd_sc_lp__dfsbp_lp.pex.spice
* Created: Fri Aug 28 10:23:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%D 1 3 8 10 12 16 18 19 23 24 25
c35 16 0 1.42388e-19 $X=0.835 $Y=0.855
c36 10 0 1.1902e-19 $X=0.835 $Y=0.78
r37 23 26 67.1496 $w=5.05e-07 $l=5.05e-07 $layer=POLY_cond $X=0.472 $Y=1.275
+ $X2=0.472 $Y2=1.78
r38 23 25 24.2607 $w=5.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.472 $Y=1.275
+ $X2=0.472 $Y2=1.11
r39 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.275 $X2=0.385 $Y2=1.275
r40 18 19 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r41 18 24 0.542326 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.275
r42 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.835 $Y=0.78
+ $X2=0.835 $Y2=0.855
r43 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.835 $Y=0.78
+ $X2=0.835 $Y2=0.495
r44 8 26 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.6 $Y=2.545 $X2=0.6
+ $Y2=1.78
r45 4 16 139.985 $w=1.5e-07 $l=2.73e-07 $layer=POLY_cond $X=0.562 $Y=0.855
+ $X2=0.835 $Y2=0.855
r46 4 13 44.6106 $w=1.5e-07 $l=8.7e-08 $layer=POLY_cond $X=0.562 $Y=0.855
+ $X2=0.475 $Y2=0.855
r47 4 25 31.9593 $w=3.25e-07 $l=1.8e-07 $layer=POLY_cond $X=0.562 $Y=0.93
+ $X2=0.562 $Y2=1.11
r48 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=0.78
+ $X2=0.475 $Y2=0.855
r49 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.475 $Y=0.78 $X2=0.475
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%CLK 3 5 7 10 12 14 15 16 19 21
c57 10 0 1.08548e-19 $X=2.075 $Y=1.135
c58 3 0 2.10375e-19 $X=1.725 $Y=2.545
r59 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.615
+ $X2=1.725 $Y2=1.45
r60 16 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.615 $X2=1.725 $Y2=1.615
r61 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.15 $Y=1.06 $X2=2.15
+ $Y2=0.775
r62 11 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.865 $Y=1.135
+ $X2=1.79 $Y2=1.135
r63 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.075 $Y=1.135
+ $X2=2.15 $Y2=1.06
r64 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.075 $Y=1.135
+ $X2=1.865 $Y2=1.135
r65 8 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.79 $Y=1.21 $X2=1.79
+ $Y2=1.135
r66 8 21 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.79 $Y=1.21 $X2=1.79
+ $Y2=1.45
r67 5 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.79 $Y=1.06 $X2=1.79
+ $Y2=1.135
r68 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.79 $Y=1.06 $X2=1.79
+ $Y2=0.775
r69 1 19 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.78
+ $X2=1.725 $Y2=1.615
r70 1 3 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.725 $Y=1.78
+ $X2=1.725 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%A_476_409# 1 2 9 13 17 21 25 27 28 31 34 35
+ 37 38 40 43 44 45 47 48 52 53 59 61 66 67
c209 67 0 1.43583e-19 $X=7.745 $Y=1.465
c210 66 0 1.422e-19 $X=7.58 $Y=1.465
c211 38 0 3.91296e-21 $X=4.355 $Y=1.495
c212 28 0 4.93603e-20 $X=2.685 $Y=2.98
c213 25 0 1.61015e-19 $X=2.52 $Y=2.475
c214 13 0 1.24203e-19 $X=4.445 $Y=0.835
r215 66 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.58 $Y=1.465
+ $X2=7.58 $Y2=1.3
r216 65 67 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.58 $Y=1.465
+ $X2=7.745 $Y2=1.465
r217 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.58
+ $Y=1.465 $X2=7.58 $Y2=1.465
r218 62 65 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.5 $Y=1.465 $X2=7.58
+ $Y2=1.465
r219 59 70 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.615
+ $X2=3.395 $Y2=1.78
r220 58 60 5.4488 $w=4.48e-07 $l=2.05e-07 $layer=LI1_cond $X=3.395 $Y=1.555
+ $X2=3.6 $Y2=1.555
r221 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.395
+ $Y=1.615 $X2=3.395 $Y2=1.615
r222 55 58 6.37908 $w=4.48e-07 $l=2.4e-07 $layer=LI1_cond $X=3.155 $Y=1.555
+ $X2=3.395 $Y2=1.555
r223 53 79 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.48 $Y=1.77
+ $X2=8.48 $Y2=1.935
r224 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.48
+ $Y=1.77 $X2=8.48 $Y2=1.77
r225 50 52 6.08838 $w=2.63e-07 $l=1.4e-07 $layer=LI1_cond $X=8.447 $Y=1.63
+ $X2=8.447 $Y2=1.77
r226 48 50 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=8.315 $Y=1.545
+ $X2=8.447 $Y2=1.63
r227 48 67 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.315 $Y=1.545
+ $X2=7.745 $Y2=1.545
r228 46 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.5 $Y=1.63 $X2=7.5
+ $Y2=1.465
r229 46 47 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=7.5 $Y=1.63
+ $X2=7.5 $Y2=2.505
r230 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.415 $Y=2.59
+ $X2=7.5 $Y2=2.505
r231 44 45 187.241 $w=1.68e-07 $l=2.87e-06 $layer=LI1_cond $X=7.415 $Y=2.59
+ $X2=4.545 $Y2=2.59
r232 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.46 $Y=2.675
+ $X2=4.545 $Y2=2.59
r233 42 43 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.46 $Y=2.675
+ $X2=4.46 $Y2=2.895
r234 41 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=2.98
+ $X2=3.6 $Y2=2.98
r235 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.375 $Y=2.98
+ $X2=4.46 $Y2=2.895
r236 40 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.375 $Y=2.98
+ $X2=3.685 $Y2=2.98
r237 38 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.495
+ $X2=4.355 $Y2=1.33
r238 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.355
+ $Y=1.495 $X2=4.355 $Y2=1.495
r239 35 60 2.25926 $w=4.48e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=1.555
+ $X2=3.6 $Y2=1.555
r240 35 37 17.8083 $w=4.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.685 $Y=1.555
+ $X2=4.355 $Y2=1.555
r241 34 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.895 $X2=3.6
+ $Y2=2.98
r242 33 60 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=3.6 $Y=1.78 $X2=3.6
+ $Y2=1.555
r243 33 34 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=3.6 $Y=1.78
+ $X2=3.6 $Y2=2.895
r244 29 55 2.55512 $w=3.3e-07 $l=2.25e-07 $layer=LI1_cond $X=3.155 $Y=1.33
+ $X2=3.155 $Y2=1.555
r245 29 31 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.155 $Y=1.33
+ $X2=3.155 $Y2=0.81
r246 27 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=2.98
+ $X2=3.6 $Y2=2.98
r247 27 28 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.515 $Y=2.98
+ $X2=2.685 $Y2=2.98
r248 23 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.52 $Y=2.895
+ $X2=2.685 $Y2=2.98
r249 23 25 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.52 $Y=2.895
+ $X2=2.52 $Y2=2.475
r250 21 79 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.47 $Y=2.595
+ $X2=8.47 $Y2=1.935
r251 17 75 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.52 $Y=0.835
+ $X2=7.52 $Y2=1.3
r252 13 72 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.445 $Y=0.835
+ $X2=4.445 $Y2=1.33
r253 9 70 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=3.435 $Y=2.595
+ $X2=3.435 $Y2=1.78
r254 2 25 300 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=2 $X=2.38
+ $Y=2.045 $X2=2.52 $Y2=2.475
r255 1 31 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.565 $X2=3.155 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%A_946_99# 1 2 9 11 13 15 16 17 19 21 24 31
c78 17 0 7.61133e-20 $X=5.695 $Y=1.3
c79 13 0 1.23194e-19 $X=4.885 $Y=2.595
c80 11 0 5.92729e-20 $X=4.885 $Y=1.885
r81 28 31 4.65142 $w=4.48e-07 $l=1.75e-07 $layer=LI1_cond $X=5.78 $Y=0.84
+ $X2=5.955 $Y2=0.84
r82 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.215
+ $Y=1.38 $X2=5.215 $Y2=1.38
r83 23 28 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=5.78 $Y=1.065
+ $X2=5.78 $Y2=0.84
r84 23 24 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.78 $Y=1.065
+ $X2=5.78 $Y2=1.215
r85 19 21 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=5.38 $Y=2.2 $X2=6.05
+ $Y2=2.2
r86 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.38 $Y=1.3
+ $X2=5.215 $Y2=1.3
r87 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.695 $Y=1.3
+ $X2=5.78 $Y2=1.215
r88 17 18 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.695 $Y=1.3
+ $X2=5.38 $Y2=1.3
r89 16 19 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=5.215 $Y=2.075
+ $X2=5.38 $Y2=2.2
r90 15 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=1.385
+ $X2=5.215 $Y2=1.3
r91 15 16 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.215 $Y=1.385
+ $X2=5.215 $Y2=2.075
r92 11 27 56.854 $w=6.26e-07 $l=5.83845e-07 $layer=POLY_cond $X=4.885 $Y=1.885
+ $X2=5.055 $Y2=1.38
r93 11 13 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.885 $Y=1.885
+ $X2=4.885 $Y2=2.595
r94 7 27 45.2819 $w=6.26e-07 $l=3.22102e-07 $layer=POLY_cond $X=4.805 $Y=1.215
+ $X2=5.055 $Y2=1.38
r95 7 9 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4.805 $Y=1.215
+ $X2=4.805 $Y2=0.835
r96 2 21 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.91
+ $Y=2.095 $X2=6.05 $Y2=2.24
r97 1 31 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=5.81
+ $Y=0.625 $X2=5.955 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%A_712_419# 1 2 9 15 19 23 27 31 32 35 37 40
+ 41 42 43 45 46 49 50 51 52 55 58 60 61 62 65 70 71 74
c189 71 0 1.43583e-19 $X=7.04 $Y=1.41
c190 70 0 1.96053e-19 $X=7.04 $Y=1.41
c191 62 0 5.92729e-20 $X=6.47 $Y=1.33
c192 61 0 1.99585e-19 $X=6.875 $Y=1.33
c193 55 0 3.013e-19 $X=5.785 $Y=1.73
c194 41 0 3.91296e-21 $X=4.195 $Y=2.16
c195 32 0 2.94985e-20 $X=7.04 $Y=1.915
r196 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.04
+ $Y=1.41 $X2=7.04 $Y2=1.41
r197 66 68 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.13 $Y=1.33
+ $X2=6.385 $Y2=1.33
r198 62 68 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=1.33
+ $X2=6.385 $Y2=1.33
r199 61 70 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.875 $Y=1.33
+ $X2=7.04 $Y2=1.33
r200 61 62 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.875 $Y=1.33
+ $X2=6.47 $Y2=1.33
r201 60 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=1.245
+ $X2=6.385 $Y2=1.33
r202 59 60 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=6.385 $Y=0.435
+ $X2=6.385 $Y2=1.245
r203 57 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=1.415
+ $X2=6.13 $Y2=1.33
r204 57 58 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.13 $Y=1.415
+ $X2=6.13 $Y2=1.565
r205 55 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.785 $Y=1.73
+ $X2=5.785 $Y2=1.565
r206 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.785
+ $Y=1.73 $X2=5.785 $Y2=1.73
r207 52 58 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.045 $Y=1.73
+ $X2=6.13 $Y2=1.565
r208 52 54 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=6.045 $Y=1.73
+ $X2=5.785 $Y2=1.73
r209 50 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.3 $Y=0.35
+ $X2=6.385 $Y2=0.435
r210 50 51 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.3 $Y=0.35
+ $X2=5.515 $Y2=0.35
r211 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.43 $Y=0.435
+ $X2=5.515 $Y2=0.35
r212 48 49 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.43 $Y=0.435
+ $X2=5.43 $Y2=0.865
r213 47 65 4.81226 $w=1.85e-07 $l=9.21954e-08 $layer=LI1_cond $X=4.87 $Y=0.95
+ $X2=4.785 $Y2=0.965
r214 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.345 $Y=0.95
+ $X2=5.43 $Y2=0.865
r215 46 47 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.345 $Y=0.95
+ $X2=4.87 $Y2=0.95
r216 44 65 1.64875 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.785 $Y=1.065
+ $X2=4.785 $Y2=0.965
r217 44 45 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.785 $Y=1.065
+ $X2=4.785 $Y2=2.075
r218 42 65 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.7 $Y=0.965
+ $X2=4.785 $Y2=0.965
r219 42 43 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=4.7 $Y=0.965
+ $X2=4.335 $Y2=0.965
r220 40 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.7 $Y=2.16
+ $X2=4.785 $Y2=2.075
r221 40 41 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.7 $Y=2.16
+ $X2=4.195 $Y2=2.16
r222 37 43 6.92652 $w=2e-07 $l=1.67705e-07 $layer=LI1_cond $X=4.21 $Y=0.865
+ $X2=4.335 $Y2=0.965
r223 37 39 5.856 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=4.21 $Y=0.865 $X2=4.21
+ $Y2=0.745
r224 33 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.03 $Y=2.245
+ $X2=4.195 $Y2=2.16
r225 33 35 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.03 $Y=2.245
+ $X2=4.03 $Y2=2.395
r226 31 71 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.04 $Y=1.75
+ $X2=7.04 $Y2=1.41
r227 31 32 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.04 $Y=1.75
+ $X2=7.04 $Y2=1.915
r228 30 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.04 $Y=1.245
+ $X2=7.04 $Y2=1.41
r229 25 27 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.875 $Y=1.29
+ $X2=6.17 $Y2=1.29
r230 23 30 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.13 $Y=0.835
+ $X2=7.13 $Y2=1.245
r231 19 32 168.948 $w=2.5e-07 $l=6.8e-07 $layer=POLY_cond $X=7.08 $Y=2.595
+ $X2=7.08 $Y2=1.915
r232 13 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.17 $Y=1.215
+ $X2=6.17 $Y2=1.29
r233 13 15 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=6.17 $Y=1.215
+ $X2=6.17 $Y2=0.835
r234 11 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.875 $Y=1.365
+ $X2=5.875 $Y2=1.29
r235 11 74 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.875 $Y=1.365
+ $X2=5.875 $Y2=1.565
r236 7 55 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.785 $Y=1.895
+ $X2=5.785 $Y2=1.73
r237 7 9 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=5.785 $Y=1.895
+ $X2=5.785 $Y2=2.595
r238 2 35 600 $w=1.7e-07 $l=6.01581e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=2.095 $X2=4.03 $Y2=2.395
r239 1 39 182 $w=1.7e-07 $l=3.8923e-07 $layer=licon1_NDIFF $count=1 $X=3.965
+ $Y=0.445 $X2=4.17 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%SET_B 3 7 9 11 12 13 16 21 22 23 24 25 30
+ 33 34 39 40
c139 40 0 1.99585e-19 $X=6.56 $Y=1.77
c140 39 0 1.78105e-19 $X=6.5 $Y=1.77
c141 33 0 9.2472e-20 $X=9.75 $Y=1.43
c142 24 0 5.84766e-20 $X=9.695 $Y=2.035
c143 7 0 7.61133e-20 $X=6.56 $Y=0.835
r144 38 40 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.5 $Y=1.77 $X2=6.56
+ $Y2=1.77
r145 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.5
+ $Y=1.77 $X2=6.5 $Y2=1.77
r146 35 38 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=6.315 $Y=1.77
+ $X2=6.5 $Y2=1.77
r147 34 49 18.844 $w=3.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.77 $Y=1.43
+ $X2=9.77 $Y2=2.035
r148 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.75
+ $Y=1.43 $X2=9.75 $Y2=1.43
r149 30 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=2.035
+ $X2=9.84 $Y2=2.035
r150 28 39 11.311 $w=2.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.53 $Y=2.035
+ $X2=6.53 $Y2=1.77
r151 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=2.035
+ $X2=6.48 $Y2=2.035
r152 25 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=2.035
+ $X2=6.48 $Y2=2.035
r153 24 30 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=2.035
+ $X2=9.84 $Y2=2.035
r154 24 25 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=9.695 $Y=2.035
+ $X2=6.625 $Y2=2.035
r155 22 33 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.75 $Y=1.77
+ $X2=9.75 $Y2=1.43
r156 22 23 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.75 $Y=1.77
+ $X2=9.75 $Y2=1.935
r157 21 33 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.75 $Y=1.265
+ $X2=9.75 $Y2=1.43
r158 18 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.69 $Y=0.975
+ $X2=9.69 $Y2=1.265
r159 16 23 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.71 $Y=2.595
+ $X2=9.71 $Y2=1.935
r160 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.615 $Y=0.9
+ $X2=9.69 $Y2=0.975
r161 12 13 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=9.615 $Y=0.9
+ $X2=8.97 $Y2=0.9
r162 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.895 $Y=0.825
+ $X2=8.97 $Y2=0.9
r163 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.895 $Y=0.825
+ $X2=8.895 $Y2=0.54
r164 5 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.56 $Y=1.605
+ $X2=6.56 $Y2=1.77
r165 5 7 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=6.56 $Y=1.605 $X2=6.56
+ $Y2=0.835
r166 1 35 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.935
+ $X2=6.315 $Y2=1.77
r167 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.315 $Y=1.935
+ $X2=6.315 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%A_263_409# 1 2 9 11 13 15 16 18 20 21 23 24
+ 28 29 30 31 32 33 35 36 38 39 40 44 45 46 48 49 52 56 60 66 70
c203 60 0 1.08548e-19 $X=2.295 $Y=1.72
c204 48 0 1.42388e-19 $X=1.295 $Y=1.075
c205 45 0 1.55371e-19 $X=2.58 $Y=1.135
c206 40 0 5.38522e-20 $X=7.695 $Y=1.945
r207 61 70 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.295 $Y=1.72
+ $X2=2.58 $Y2=1.72
r208 61 67 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=2.295 $Y=1.72
+ $X2=2.255 $Y2=1.72
r209 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=1.72 $X2=2.295 $Y2=1.72
r210 58 60 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=2.295 $Y=1.96
+ $X2=2.295 $Y2=1.72
r211 57 66 3.35233 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=1.625 $Y=2.045
+ $X2=1.417 $Y2=2.045
r212 56 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.13 $Y=2.045
+ $X2=2.295 $Y2=1.96
r213 56 57 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.13 $Y=2.045
+ $X2=1.625 $Y2=2.045
r214 52 54 19.7165 $w=4.13e-07 $l=7.1e-07 $layer=LI1_cond $X=1.417 $Y=2.19
+ $X2=1.417 $Y2=2.9
r215 50 66 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=1.417 $Y=2.13
+ $X2=1.417 $Y2=2.045
r216 50 52 1.66618 $w=4.13e-07 $l=6e-08 $layer=LI1_cond $X=1.417 $Y=2.13
+ $X2=1.417 $Y2=2.19
r217 49 66 3.22182 $w=2.92e-07 $l=1.58915e-07 $layer=LI1_cond $X=1.295 $Y=1.96
+ $X2=1.417 $Y2=2.045
r218 48 65 9.76 $w=3.5e-07 $l=3.77889e-07 $layer=LI1_cond $X=1.295 $Y=1.075
+ $X2=1.575 $Y2=0.845
r219 48 49 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.295 $Y=1.075
+ $X2=1.295 $Y2=1.96
r220 42 44 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=8.03 $Y=1.87
+ $X2=8.03 $Y2=0.835
r221 41 44 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.03 $Y=0.255
+ $X2=8.03 $Y2=0.835
r222 39 42 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.955 $Y=1.945
+ $X2=8.03 $Y2=1.87
r223 39 40 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=7.955 $Y=1.945
+ $X2=7.695 $Y2=1.945
r224 36 40 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=7.57 $Y=2.02
+ $X2=7.695 $Y2=1.945
r225 36 38 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.57 $Y=2.02
+ $X2=7.57 $Y2=2.595
r226 33 35 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.295 $Y=2.02
+ $X2=4.295 $Y2=2.595
r227 31 41 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.955 $Y=0.18
+ $X2=8.03 $Y2=0.255
r228 31 32 2045.94 $w=1.5e-07 $l=3.99e-06 $layer=POLY_cond $X=7.955 $Y=0.18
+ $X2=3.965 $Y2=0.18
r229 29 33 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=4.17 $Y=1.945
+ $X2=4.295 $Y2=2.02
r230 29 30 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=4.17 $Y=1.945
+ $X2=3.95 $Y2=1.945
r231 26 47 59.6593 $w=1.58e-07 $l=1.9896e-07 $layer=POLY_cond $X=3.89 $Y=0.94
+ $X2=3.882 $Y2=1.135
r232 26 28 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.89 $Y=0.94
+ $X2=3.89 $Y2=0.655
r233 25 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.89 $Y=0.255
+ $X2=3.965 $Y2=0.18
r234 25 28 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.89 $Y=0.255
+ $X2=3.89 $Y2=0.655
r235 24 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.875 $Y=1.87
+ $X2=3.95 $Y2=1.945
r236 23 47 23.0517 $w=1.58e-07 $l=7.84219e-08 $layer=POLY_cond $X=3.875 $Y=1.21
+ $X2=3.882 $Y2=1.135
r237 23 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.875 $Y=1.21
+ $X2=3.875 $Y2=1.87
r238 22 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.015 $Y=1.135
+ $X2=2.94 $Y2=1.135
r239 21 47 4.07462 $w=1.5e-07 $l=8.2e-08 $layer=POLY_cond $X=3.8 $Y=1.135
+ $X2=3.882 $Y2=1.135
r240 21 22 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=3.8 $Y=1.135
+ $X2=3.015 $Y2=1.135
r241 18 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.94 $Y=1.06
+ $X2=2.94 $Y2=1.135
r242 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.94 $Y=1.06
+ $X2=2.94 $Y2=0.775
r243 17 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.135
+ $X2=2.58 $Y2=1.135
r244 16 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=1.135
+ $X2=2.94 $Y2=1.135
r245 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.865 $Y=1.135
+ $X2=2.655 $Y2=1.135
r246 15 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.555
+ $X2=2.58 $Y2=1.72
r247 14 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.21
+ $X2=2.58 $Y2=1.135
r248 14 15 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.58 $Y=1.21
+ $X2=2.58 $Y2=1.555
r249 11 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.06
+ $X2=2.58 $Y2=1.135
r250 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.58 $Y=1.06
+ $X2=2.58 $Y2=0.775
r251 7 67 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.885
+ $X2=2.255 $Y2=1.72
r252 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.255 $Y=1.885
+ $X2=2.255 $Y2=2.545
r253 2 54 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=2.045 $X2=1.46 $Y2=2.9
r254 2 52 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=2.045 $X2=1.46 $Y2=2.19
r255 1 65 182 $w=1.7e-07 $l=3.03109e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.565 $X2=1.575 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%A_1686_40# 1 2 9 11 12 15 19 22 23 25 26 29
+ 31 35 37
c97 25 0 9.2472e-20 $X=9.755 $Y=1
c98 19 0 2.89781e-20 $X=9.13 $Y=1.885
c99 11 0 1.1224e-19 $X=8.885 $Y=1.29
r100 33 35 48.8636 $w=2.48e-07 $l=1.06e-06 $layer=LI1_cond $X=10.49 $Y=1.085
+ $X2=10.49 $Y2=2.145
r101 32 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.085 $Y=1
+ $X2=9.92 $Y2=1
r102 31 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.365 $Y=1
+ $X2=10.49 $Y2=1.085
r103 31 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.365 $Y=1
+ $X2=10.085 $Y2=1
r104 27 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.92 $Y=0.915
+ $X2=9.92 $Y2=1
r105 27 29 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=9.92 $Y=0.915
+ $X2=9.92 $Y2=0.495
r106 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.755 $Y=1 $X2=9.92
+ $Y2=1
r107 25 26 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.755 $Y=1
+ $X2=9.375 $Y2=1
r108 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.21
+ $Y=1.38 $X2=9.21 $Y2=1.38
r109 20 26 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=9.242 $Y=1.085
+ $X2=9.375 $Y2=1
r110 20 22 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=9.242 $Y=1.085
+ $X2=9.242 $Y2=1.38
r111 18 23 28.3893 $w=4.9e-07 $l=2.6e-07 $layer=POLY_cond $X=9.13 $Y=1.64
+ $X2=9.13 $Y2=1.38
r112 18 19 39.5539 $w=4.9e-07 $l=2.45e-07 $layer=POLY_cond $X=9.13 $Y=1.64
+ $X2=9.13 $Y2=1.885
r113 17 23 1.63785 $w=4.9e-07 $l=1.5e-08 $layer=POLY_cond $X=9.13 $Y=1.365
+ $X2=9.13 $Y2=1.38
r114 15 19 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=9.01 $Y=2.595
+ $X2=9.01 $Y2=1.885
r115 11 17 38.2759 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=8.885 $Y=1.29
+ $X2=9.13 $Y2=1.365
r116 11 12 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=8.885 $Y=1.29
+ $X2=8.58 $Y2=1.29
r117 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.505 $Y=1.215
+ $X2=8.58 $Y2=1.29
r118 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=8.505 $Y=1.215
+ $X2=8.505 $Y2=0.54
r119 2 35 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=10.385
+ $Y=2 $X2=10.53 $Y2=2.145
r120 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=9.775
+ $Y=0.285 $X2=9.92 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%A_1519_125# 1 2 3 10 12 13 14 15 17 19 22
+ 24 26 27 28 29 31 33 36 39 40 41 42 44 47 49 51 52 55 58 62 64 65 66 69 70 72
+ 73 74 75 78 82 86 89 92 97
c220 97 0 1.8111e-19 $X=11.125 $Y=1.505
r221 93 95 23.9565 $w=6.7e-07 $l=3e-07 $layer=POLY_cond $X=10.495 $Y=1.505
+ $X2=10.795 $Y2=1.505
r222 86 88 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.97 $Y=2.24
+ $X2=7.97 $Y2=2.415
r223 82 92 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=10.88 $Y=2.895
+ $X2=10.88 $Y2=1.84
r224 79 97 51.5677 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.96 $Y=1.505
+ $X2=11.125 $Y2=1.505
r225 79 95 13.1761 $w=6.7e-07 $l=1.65e-07 $layer=POLY_cond $X=10.96 $Y=1.505
+ $X2=10.795 $Y2=1.505
r226 78 79 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.96
+ $Y=1.335 $X2=10.96 $Y2=1.335
r227 76 92 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.96 $Y=1.675
+ $X2=10.96 $Y2=1.84
r228 76 78 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=10.96 $Y=1.675
+ $X2=10.96 $Y2=1.335
r229 74 82 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.795 $Y=2.98
+ $X2=10.88 $Y2=2.895
r230 74 75 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=10.795 $Y=2.98
+ $X2=10.14 $Y2=2.98
r231 73 75 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.975 $Y=2.895
+ $X2=10.14 $Y2=2.98
r232 72 91 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.975 $Y=2.5
+ $X2=9.975 $Y2=2.415
r233 72 73 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=9.975 $Y=2.5
+ $X2=9.975 $Y2=2.895
r234 71 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.93 $Y=2.415
+ $X2=8.845 $Y2=2.415
r235 70 91 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.81 $Y=2.415
+ $X2=9.975 $Y2=2.415
r236 70 71 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=9.81 $Y=2.415
+ $X2=8.93 $Y2=2.415
r237 69 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.845 $Y=2.33
+ $X2=8.845 $Y2=2.415
r238 68 69 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=8.845 $Y=1.085
+ $X2=8.845 $Y2=2.33
r239 67 88 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.135 $Y=2.415
+ $X2=7.97 $Y2=2.415
r240 66 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=2.415
+ $X2=8.845 $Y2=2.415
r241 66 67 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=8.76 $Y=2.415
+ $X2=8.135 $Y2=2.415
r242 65 84 12.5109 $w=4.67e-07 $l=3.48999e-07 $layer=LI1_cond $X=8.095 $Y=1
+ $X2=7.815 $Y2=0.845
r243 64 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.76 $Y=1
+ $X2=8.845 $Y2=1.085
r244 64 65 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=8.76 $Y=1 $X2=8.095
+ $Y2=1
r245 60 88 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=2.5
+ $X2=7.97 $Y2=2.415
r246 60 62 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=7.97 $Y=2.5 $X2=7.97
+ $Y2=2.9
r247 53 54 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=11.285 $Y=0.855
+ $X2=11.545 $Y2=0.855
r248 49 58 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.635 $Y=0.78
+ $X2=12.635 $Y2=0.855
r249 49 51 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.635 $Y=0.78
+ $X2=12.635 $Y2=0.495
r250 45 58 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=12.585 $Y=0.855
+ $X2=12.635 $Y2=0.855
r251 45 56 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=12.585 $Y=0.855
+ $X2=12.275 $Y2=0.855
r252 45 47 357.773 $w=2.5e-07 $l=1.44e-06 $layer=POLY_cond $X=12.585 $Y=0.93
+ $X2=12.585 $Y2=2.37
r253 42 56 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.275 $Y=0.78
+ $X2=12.275 $Y2=0.855
r254 42 44 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.275 $Y=0.78
+ $X2=12.275 $Y2=0.495
r255 41 54 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.62 $Y=0.855
+ $X2=11.545 $Y2=0.855
r256 40 56 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.2 $Y=0.855
+ $X2=12.275 $Y2=0.855
r257 40 41 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=12.2 $Y=0.855
+ $X2=11.62 $Y2=0.855
r258 39 55 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=11.545 $Y=1.17
+ $X2=11.495 $Y2=1.245
r259 38 54 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.545 $Y=0.93
+ $X2=11.545 $Y2=0.855
r260 38 39 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.545 $Y=0.93
+ $X2=11.545 $Y2=1.17
r261 34 55 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=11.495 $Y=1.32
+ $X2=11.495 $Y2=1.245
r262 34 36 293.175 $w=2.5e-07 $l=1.18e-06 $layer=POLY_cond $X=11.495 $Y=1.32
+ $X2=11.495 $Y2=2.5
r263 31 53 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.285 $Y=0.78
+ $X2=11.285 $Y2=0.855
r264 31 33 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.285 $Y=0.78
+ $X2=11.285 $Y2=0.495
r265 29 55 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=11.37 $Y=1.245
+ $X2=11.495 $Y2=1.245
r266 29 97 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=11.37 $Y=1.245
+ $X2=11.125 $Y2=1.245
r267 27 53 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.21 $Y=0.855
+ $X2=11.285 $Y2=0.855
r268 27 28 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=11.21 $Y=0.855
+ $X2=11 $Y2=0.855
r269 24 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.925 $Y=0.78
+ $X2=11 $Y2=0.855
r270 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.925 $Y=0.78
+ $X2=10.925 $Y2=0.495
r271 20 95 25.9839 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.795 $Y=1.84
+ $X2=10.795 $Y2=1.505
r272 20 22 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.795 $Y=1.84
+ $X2=10.795 $Y2=2.5
r273 19 93 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.495 $Y=1.17
+ $X2=10.495 $Y2=1.505
r274 18 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.495 $Y=0.93
+ $X2=10.495 $Y2=0.855
r275 18 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.495 $Y=0.93
+ $X2=10.495 $Y2=1.17
r276 15 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.495 $Y=0.78
+ $X2=10.495 $Y2=0.855
r277 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.495 $Y=0.78
+ $X2=10.495 $Y2=0.495
r278 13 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.42 $Y=0.855
+ $X2=10.495 $Y2=0.855
r279 13 14 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.42 $Y=0.855
+ $X2=10.21 $Y2=0.855
r280 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.135 $Y=0.78
+ $X2=10.21 $Y2=0.855
r281 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.135 $Y=0.78
+ $X2=10.135 $Y2=0.495
r282 3 91 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=9.835
+ $Y=2.095 $X2=9.975 $Y2=2.495
r283 2 86 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=7.695
+ $Y=2.095 $X2=7.97 $Y2=2.24
r284 2 62 600 $w=1.7e-07 $l=9.32416e-07 $layer=licon1_PDIFF $count=1 $X=7.695
+ $Y=2.095 $X2=7.97 $Y2=2.9
r285 1 84 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=7.595
+ $Y=0.625 $X2=7.815 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%A_2383_57# 1 2 9 13 17 23 26 28 31 35 39 40
+ 43 46
c67 46 0 6.93588e-20 $X=12.295 $Y=1.575
r68 43 45 10.5425 $w=3.78e-07 $l=2.3e-07 $layer=LI1_cond $X=12.085 $Y=0.495
+ $X2=12.085 $Y2=0.725
r69 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.155
+ $Y=1.155 $X2=13.155 $Y2=1.155
r70 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=13.155 $Y=1.49
+ $X2=13.155 $Y2=1.155
r71 36 46 3.11956 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=12.485 $Y=1.575
+ $X2=12.295 $Y2=1.575
r72 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.99 $Y=1.575
+ $X2=13.155 $Y2=1.49
r73 35 36 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=12.99 $Y=1.575
+ $X2=12.485 $Y2=1.575
r74 31 33 21.5325 $w=3.78e-07 $l=7.1e-07 $layer=LI1_cond $X=12.295 $Y=2.015
+ $X2=12.295 $Y2=2.725
r75 29 46 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=12.295 $Y=1.66
+ $X2=12.295 $Y2=1.575
r76 29 31 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=12.295 $Y=1.66
+ $X2=12.295 $Y2=2.015
r77 28 46 3.40559 $w=2.75e-07 $l=1.41244e-07 $layer=LI1_cond $X=12.19 $Y=1.49
+ $X2=12.295 $Y2=1.575
r78 28 45 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=12.19 $Y=1.49
+ $X2=12.19 $Y2=0.725
r79 25 40 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=13.155 $Y=1.495
+ $X2=13.155 $Y2=1.155
r80 25 26 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.155 $Y=1.495
+ $X2=13.155 $Y2=1.66
r81 22 40 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=13.155 $Y=1.14
+ $X2=13.155 $Y2=1.155
r82 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=13.155 $Y=1.065
+ $X2=13.425 $Y2=1.065
r83 19 22 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=13.065 $Y=1.065
+ $X2=13.155 $Y2=1.065
r84 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.425 $Y=0.99
+ $X2=13.425 $Y2=1.065
r85 15 17 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=13.425 $Y=0.99
+ $X2=13.425 $Y2=0.495
r86 13 26 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=13.115 $Y=2.37
+ $X2=13.115 $Y2=1.66
r87 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.065 $Y=0.99
+ $X2=13.065 $Y2=1.065
r88 7 9 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=13.065 $Y=0.99
+ $X2=13.065 $Y2=0.495
r89 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.175
+ $Y=1.87 $X2=12.32 $Y2=2.725
r90 2 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.175
+ $Y=1.87 $X2=12.32 $Y2=2.015
r91 1 43 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=11.915
+ $Y=0.285 $X2=12.06 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 42 46 50
+ 55 56 58 59 60 69 80 87 92 99 100 106 109 112 115
r141 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r142 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r143 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r144 106 107 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r145 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r146 100 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=12.72 $Y2=3.33
r147 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r148 97 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.015 $Y=3.33
+ $X2=12.85 $Y2=3.33
r149 97 99 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=13.015 $Y=3.33
+ $X2=13.68 $Y2=3.33
r150 96 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r151 96 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r152 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r153 93 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.395 $Y=3.33
+ $X2=11.27 $Y2=3.33
r154 93 95 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.395 $Y=3.33
+ $X2=11.76 $Y2=3.33
r155 92 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.685 $Y=3.33
+ $X2=12.85 $Y2=3.33
r156 92 95 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=12.685 $Y=3.33
+ $X2=11.76 $Y2=3.33
r157 91 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r158 91 110 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=9.36 $Y2=3.33
r159 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r160 88 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.44 $Y=3.33
+ $X2=9.275 $Y2=3.33
r161 88 90 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=9.44 $Y=3.33
+ $X2=10.8 $Y2=3.33
r162 87 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.145 $Y=3.33
+ $X2=11.27 $Y2=3.33
r163 87 90 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.145 $Y=3.33
+ $X2=10.8 $Y2=3.33
r164 86 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r165 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r166 82 85 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 80 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.11 $Y=3.33
+ $X2=9.275 $Y2=3.33
r168 80 85 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.11 $Y=3.33
+ $X2=8.88 $Y2=3.33
r169 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r170 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r171 76 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r172 75 78 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r173 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r174 73 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.15 $Y2=3.33
r175 73 75 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.52 $Y2=3.33
r176 72 107 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=5.04 $Y2=3.33
r177 71 72 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r178 69 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=5.15 $Y2=3.33
r179 69 71 184.305 $w=1.68e-07 $l=2.825e-06 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=2.16 $Y2=3.33
r180 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r181 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r182 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r183 65 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r184 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r185 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r186 62 103 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=3.33
+ $X2=0.25 $Y2=3.33
r187 62 64 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.5 $Y=3.33
+ $X2=0.72 $Y2=3.33
r188 60 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r189 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r190 60 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r191 58 78 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.48 $Y2=3.33
r192 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.66 $Y2=3.33
r193 57 82 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.96 $Y2=3.33
r194 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.66 $Y2=3.33
r195 55 67 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.68 $Y2=3.33
r196 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.99 $Y2=3.33
r197 54 71 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=2.16 $Y2=3.33
r198 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=1.99 $Y2=3.33
r199 50 53 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=12.85 $Y=2.015
+ $X2=12.85 $Y2=2.725
r200 48 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.85 $Y=3.245
+ $X2=12.85 $Y2=3.33
r201 48 53 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=12.85 $Y=3.245
+ $X2=12.85 $Y2=2.725
r202 44 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.27 $Y=3.245
+ $X2=11.27 $Y2=3.33
r203 44 46 48.8636 $w=2.48e-07 $l=1.06e-06 $layer=LI1_cond $X=11.27 $Y=3.245
+ $X2=11.27 $Y2=2.185
r204 40 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.275 $Y=3.245
+ $X2=9.275 $Y2=3.33
r205 40 42 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=9.275 $Y=3.245
+ $X2=9.275 $Y2=2.895
r206 36 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.66 $Y=3.245
+ $X2=6.66 $Y2=3.33
r207 36 38 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=6.66 $Y=3.245
+ $X2=6.66 $Y2=3.02
r208 32 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=3.33
r209 32 34 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=2.945
r210 28 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=3.33
r211 28 30 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=2.475
r212 24 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.335 $Y=2.19
+ $X2=0.335 $Y2=2.9
r213 22 103 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=3.245
+ $X2=0.25 $Y2=3.33
r214 22 27 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.335 $Y=3.245
+ $X2=0.335 $Y2=2.9
r215 7 53 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=12.71
+ $Y=1.87 $X2=12.85 $Y2=2.725
r216 7 50 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.71
+ $Y=1.87 $X2=12.85 $Y2=2.015
r217 6 46 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=10.92
+ $Y=2 $X2=11.23 $Y2=2.185
r218 5 42 600 $w=1.7e-07 $l=8.67179e-07 $layer=licon1_PDIFF $count=1 $X=9.135
+ $Y=2.095 $X2=9.275 $Y2=2.895
r219 4 38 600 $w=1.7e-07 $l=1.02914e-06 $layer=licon1_PDIFF $count=1 $X=6.44
+ $Y=2.095 $X2=6.66 $Y2=3.02
r220 3 34 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=5.01
+ $Y=2.095 $X2=5.15 $Y2=2.945
r221 2 30 300 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=2 $X=1.85
+ $Y=2.045 $X2=1.99 $Y2=2.475
r222 1 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=2.045 $X2=0.335 $Y2=2.9
r223 1 24 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=2.045 $X2=0.335 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%A_145_409# 1 2 3 4 15 17 21 24 25 26 28 30
+ 31 32 33 34 37 41 43 44 49
c115 49 0 1.55371e-19 $X=2.725 $Y=1.185
c116 41 0 1.24203e-19 $X=3.675 $Y=0.655
c117 21 0 1.1902e-19 $X=1.92 $Y=0.35
r118 47 48 10.6092 $w=3.53e-07 $l=2.3e-07 $layer=LI1_cond $X=1.037 $Y=0.495
+ $X2=1.037 $Y2=0.725
r119 44 47 4.70716 $w=3.53e-07 $l=1.45e-07 $layer=LI1_cond $X=1.037 $Y=0.35
+ $X2=1.037 $Y2=0.495
r120 43 48 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=0.945 $Y=2.025
+ $X2=0.945 $Y2=0.725
r121 39 41 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.675 $Y=0.435
+ $X2=3.675 $Y2=0.655
r122 35 37 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.17 $Y=2.13
+ $X2=3.17 $Y2=2.395
r123 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.005 $Y=2.045
+ $X2=3.17 $Y2=2.13
r124 33 34 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.005 $Y=2.045
+ $X2=2.81 $Y2=2.045
r125 31 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.51 $Y=0.35
+ $X2=3.675 $Y2=0.435
r126 31 32 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.51 $Y=0.35 $X2=2.81
+ $Y2=0.35
r127 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.725 $Y=1.96
+ $X2=2.81 $Y2=2.045
r128 29 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=1.27
+ $X2=2.725 $Y2=1.185
r129 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.725 $Y=1.27
+ $X2=2.725 $Y2=1.96
r130 28 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=1.1
+ $X2=2.725 $Y2=1.185
r131 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.725 $Y=0.435
+ $X2=2.81 $Y2=0.35
r132 27 28 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.725 $Y=0.435
+ $X2=2.725 $Y2=1.1
r133 25 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.185
+ $X2=2.725 $Y2=1.185
r134 25 26 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.64 $Y=1.185
+ $X2=2.09 $Y2=1.185
r135 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.005 $Y=1.1
+ $X2=2.09 $Y2=1.185
r136 23 24 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.005 $Y=0.435
+ $X2=2.005 $Y2=1.1
r137 22 44 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.215 $Y=0.35
+ $X2=1.037 $Y2=0.35
r138 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.92 $Y=0.35
+ $X2=2.005 $Y2=0.435
r139 21 22 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.92 $Y=0.35
+ $X2=1.215 $Y2=0.35
r140 15 43 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=2.19
+ $X2=0.865 $Y2=2.025
r141 15 17 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.865 $Y=2.19
+ $X2=0.865 $Y2=2.9
r142 4 37 600 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=1 $X=3.025
+ $Y=2.095 $X2=3.17 $Y2=2.395
r143 3 17 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.725
+ $Y=2.045 $X2=0.865 $Y2=2.9
r144 3 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.725
+ $Y=2.045 $X2=0.865 $Y2=2.19
r145 2 41 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.55
+ $Y=0.445 $X2=3.675 $Y2=0.655
r146 1 47 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.285 $X2=1.05 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%Q_N 1 2 11 16 19 20 24
c39 11 0 1.8111e-19 $X=11.76 $Y=2.145
r40 20 28 3.73456 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.71 $Y=1.665
+ $X2=11.71 $Y2=1.78
r41 19 20 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.71 $Y=1.295
+ $X2=11.71 $Y2=1.665
r42 19 24 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.71 $Y=1.295
+ $X2=11.71 $Y2=1.18
r43 18 24 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=11.58 $Y=0.725
+ $X2=11.58 $Y2=1.18
r44 16 18 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=11.5 $Y=0.495
+ $X2=11.5 $Y2=0.725
r45 11 13 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=11.76 $Y=2.145
+ $X2=11.76 $Y2=2.855
r46 11 28 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=11.76 $Y=2.145
+ $X2=11.76 $Y2=1.78
r47 2 13 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=11.62
+ $Y=2 $X2=11.76 $Y2=2.855
r48 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.62
+ $Y=2 $X2=11.76 $Y2=2.145
r49 1 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.36
+ $Y=0.285 $X2=11.5 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%Q 1 2 10 13 14 15 28 29
r23 28 29 10.0909 $w=5.88e-07 $l=1.65e-07 $layer=LI1_cond $X=13.51 $Y=2.015
+ $X2=13.51 $Y2=1.85
r24 15 23 1.01363 $w=5.88e-07 $l=5e-08 $layer=LI1_cond $X=13.51 $Y=2.775
+ $X2=13.51 $Y2=2.725
r25 14 23 6.48721 $w=5.88e-07 $l=3.2e-07 $layer=LI1_cond $X=13.51 $Y=2.405
+ $X2=13.51 $Y2=2.725
r26 14 19 5.27085 $w=5.88e-07 $l=2.6e-07 $layer=LI1_cond $X=13.51 $Y=2.405
+ $X2=13.51 $Y2=2.145
r27 13 19 2.22998 $w=5.88e-07 $l=1.1e-07 $layer=LI1_cond $X=13.51 $Y=2.035
+ $X2=13.51 $Y2=2.145
r28 13 28 0.40545 $w=5.88e-07 $l=2e-08 $layer=LI1_cond $X=13.51 $Y=2.035
+ $X2=13.51 $Y2=2.015
r29 12 29 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=13.72 $Y=0.725
+ $X2=13.72 $Y2=1.85
r30 10 12 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=13.64 $Y=0.495
+ $X2=13.64 $Y2=0.725
r31 2 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.24
+ $Y=1.87 $X2=13.38 $Y2=2.015
r32 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=13.24
+ $Y=1.87 $X2=13.38 $Y2=2.725
r33 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.5
+ $Y=0.285 $X2=13.64 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFSBP_LP%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46
+ 50 53 54 56 57 58 67 74 89 98 99 105 108 111 114
c147 40 0 1.1224e-19 $X=9.11 $Y=0.52
r148 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r149 112 115 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=12.72 $Y2=0
r150 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r151 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r152 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r153 99 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=12.72 $Y2=0
r154 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r155 96 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.015 $Y=0
+ $X2=12.85 $Y2=0
r156 96 98 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=13.015 $Y=0
+ $X2=13.68 $Y2=0
r157 95 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r158 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r159 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.32 $Y2=0
r160 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=0 $X2=10.32
+ $Y2=0
r161 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r162 89 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.545 $Y=0
+ $X2=10.71 $Y2=0
r163 89 94 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=10.545 $Y=0
+ $X2=10.32 $Y2=0
r164 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r165 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r166 85 88 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.88 $Y2=0
r167 84 87 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=7.44 $Y=0 $X2=8.88
+ $Y2=0
r168 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r169 82 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.08 $Y=0
+ $X2=6.915 $Y2=0
r170 82 84 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.08 $Y=0 $X2=7.44
+ $Y2=0
r171 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r172 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r173 78 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r174 77 80 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r175 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r176 75 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.04 $Y2=0
r177 75 77 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.52 $Y2=0
r178 74 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.75 $Y=0
+ $X2=6.915 $Y2=0
r179 74 80 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.75 $Y=0 $X2=6.48
+ $Y2=0
r180 73 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r181 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r182 70 73 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r183 69 72 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r184 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r185 67 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=5.04 $Y2=0
r186 67 72 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=4.56 $Y2=0
r187 66 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r188 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r189 63 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=2.16 $Y2=0
r190 63 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r191 62 65 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r192 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r193 60 102 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r194 60 62 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r195 58 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r196 58 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r197 58 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r198 56 87 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=8.945 $Y=0 $X2=8.88
+ $Y2=0
r199 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.945 $Y=0 $X2=9.11
+ $Y2=0
r200 55 91 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.275 $Y=0 $X2=9.36
+ $Y2=0
r201 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.275 $Y=0 $X2=9.11
+ $Y2=0
r202 53 65 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.16
+ $Y2=0
r203 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.365
+ $Y2=0
r204 52 69 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.64
+ $Y2=0
r205 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.365
+ $Y2=0
r206 48 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.85 $Y=0.085
+ $X2=12.85 $Y2=0
r207 48 50 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=12.85 $Y=0.085
+ $X2=12.85 $Y2=0.495
r208 47 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.875 $Y=0
+ $X2=10.71 $Y2=0
r209 46 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.685 $Y=0
+ $X2=12.85 $Y2=0
r210 46 47 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=12.685 $Y=0
+ $X2=10.875 $Y2=0
r211 42 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.71 $Y=0.085
+ $X2=10.71 $Y2=0
r212 42 44 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.71 $Y=0.085
+ $X2=10.71 $Y2=0.495
r213 38 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.11 $Y=0.085
+ $X2=9.11 $Y2=0
r214 38 40 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=9.11 $Y=0.085
+ $X2=9.11 $Y2=0.52
r215 34 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=0.085
+ $X2=6.915 $Y2=0
r216 34 36 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=6.915 $Y=0.085
+ $X2=6.915 $Y2=0.835
r217 30 105 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0
r218 30 32 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0.52
r219 26 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.365 $Y=0.085
+ $X2=2.365 $Y2=0
r220 26 28 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.365 $Y=0.085
+ $X2=2.365 $Y2=0.73
r221 22 102 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r222 22 24 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.495
r223 7 50 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.71
+ $Y=0.285 $X2=12.85 $Y2=0.495
r224 6 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.57
+ $Y=0.285 $X2=10.71 $Y2=0.495
r225 5 40 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=8.97
+ $Y=0.33 $X2=9.11 $Y2=0.52
r226 4 36 182 $w=1.7e-07 $l=3.70405e-07 $layer=licon1_NDIFF $count=1 $X=6.635
+ $Y=0.625 $X2=6.915 $Y2=0.835
r227 3 32 182 $w=1.7e-07 $l=2.46982e-07 $layer=licon1_NDIFF $count=1 $X=4.88
+ $Y=0.625 $X2=5.08 $Y2=0.52
r228 2 28 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.565 $X2=2.365 $Y2=0.73
r229 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.26 $Y2=0.495
.ends

