# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a221oi_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a221oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.960000 1.210000 5.165000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.540000 1.345000 3.790000 1.615000 ;
        RECT 3.540000 1.615000 5.675000 1.785000 ;
        RECT 5.335000 1.210000 5.675000 1.615000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.425000 1.210000 2.815000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 1.425000 2.255000 1.615000 ;
        RECT 1.025000 1.615000 3.330000 1.785000 ;
        RECT 3.000000 1.375000 3.330000 1.615000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.465000 1.750000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.058400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.920000 0.855000 2.735000 ;
        RECT 0.635000 0.255000 0.895000 0.785000 ;
        RECT 0.635000 0.785000 4.465000 1.040000 ;
        RECT 0.635000 1.040000 0.855000 1.920000 ;
        RECT 4.205000 0.665000 4.465000 0.785000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.095000  1.925000 0.355000 2.905000 ;
      RECT 0.095000  2.905000 1.285000 3.075000 ;
      RECT 0.205000  0.085000 0.465000 1.040000 ;
      RECT 1.025000  1.955000 3.095000 2.125000 ;
      RECT 1.025000  2.125000 1.285000 2.905000 ;
      RECT 1.065000  0.085000 1.775000 0.615000 ;
      RECT 1.475000  2.295000 1.735000 2.905000 ;
      RECT 1.475000  2.905000 3.550000 3.075000 ;
      RECT 1.905000  2.125000 2.235000 2.735000 ;
      RECT 1.955000  0.285000 3.085000 0.615000 ;
      RECT 2.405000  2.295000 2.595000 2.905000 ;
      RECT 2.765000  2.125000 3.095000 2.735000 ;
      RECT 3.260000  0.085000 3.590000 0.615000 ;
      RECT 3.265000  1.955000 5.395000 2.125000 ;
      RECT 3.265000  2.125000 3.550000 2.905000 ;
      RECT 3.720000  2.295000 4.050000 3.245000 ;
      RECT 3.775000  0.255000 4.965000 0.485000 ;
      RECT 4.220000  2.125000 4.455000 3.075000 ;
      RECT 4.635000  0.485000 4.965000 1.040000 ;
      RECT 4.635000  2.295000 4.965000 3.245000 ;
      RECT 5.135000  0.085000 5.395000 1.040000 ;
      RECT 5.145000  2.125000 5.395000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__a221oi_2
