* File: sky130_fd_sc_lp__a221oi_1.pxi.spice
* Created: Fri Aug 28 09:53:18 2020
* 
x_PM_SKY130_FD_SC_LP__A221OI_1%C1 N_C1_M1009_g N_C1_M1007_g C1 C1 N_C1_c_55_n
+ PM_SKY130_FD_SC_LP__A221OI_1%C1
x_PM_SKY130_FD_SC_LP__A221OI_1%B2 N_B2_M1001_g N_B2_M1004_g B2 N_B2_c_86_n
+ N_B2_c_87_n N_B2_c_88_n PM_SKY130_FD_SC_LP__A221OI_1%B2
x_PM_SKY130_FD_SC_LP__A221OI_1%B1 N_B1_M1003_g N_B1_M1006_g B1 N_B1_c_123_n
+ N_B1_c_124_n N_B1_c_125_n PM_SKY130_FD_SC_LP__A221OI_1%B1
x_PM_SKY130_FD_SC_LP__A221OI_1%A1 N_A1_M1005_g N_A1_M1000_g A1 A1 A1
+ N_A1_c_157_n N_A1_c_158_n PM_SKY130_FD_SC_LP__A221OI_1%A1
x_PM_SKY130_FD_SC_LP__A221OI_1%A2 N_A2_M1008_g N_A2_M1002_g A2 N_A2_c_188_n
+ N_A2_c_189_n PM_SKY130_FD_SC_LP__A221OI_1%A2
x_PM_SKY130_FD_SC_LP__A221OI_1%Y N_Y_M1007_s N_Y_M1003_d N_Y_M1009_s N_Y_c_213_n
+ N_Y_c_234_p Y Y Y Y Y Y Y N_Y_c_211_n PM_SKY130_FD_SC_LP__A221OI_1%Y
x_PM_SKY130_FD_SC_LP__A221OI_1%A_110_367# N_A_110_367#_M1009_d
+ N_A_110_367#_M1004_d N_A_110_367#_c_241_n N_A_110_367#_c_242_n
+ N_A_110_367#_c_243_n N_A_110_367#_c_254_p
+ PM_SKY130_FD_SC_LP__A221OI_1%A_110_367#
x_PM_SKY130_FD_SC_LP__A221OI_1%A_217_367# N_A_217_367#_M1004_s
+ N_A_217_367#_M1006_d N_A_217_367#_M1002_d N_A_217_367#_c_261_n
+ N_A_217_367#_c_262_n N_A_217_367#_c_263_n N_A_217_367#_c_298_p
+ N_A_217_367#_c_264_n N_A_217_367#_c_265_n N_A_217_367#_c_266_n
+ PM_SKY130_FD_SC_LP__A221OI_1%A_217_367#
x_PM_SKY130_FD_SC_LP__A221OI_1%VPWR N_VPWR_M1000_d N_VPWR_c_306_n VPWR
+ N_VPWR_c_307_n N_VPWR_c_308_n N_VPWR_c_305_n N_VPWR_c_310_n
+ PM_SKY130_FD_SC_LP__A221OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A221OI_1%VGND N_VGND_M1007_d N_VGND_M1008_d N_VGND_c_341_n
+ N_VGND_c_342_n N_VGND_c_343_n VGND N_VGND_c_344_n N_VGND_c_345_n
+ PM_SKY130_FD_SC_LP__A221OI_1%VGND
cc_1 VNB N_C1_M1009_g 0.00749333f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB N_C1_M1007_g 0.0233518f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.655
cc_3 VNB C1 0.00317638f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_C1_c_55_n 0.0493633f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.375
cc_5 VNB N_B2_M1004_g 0.00881992f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.655
cc_6 VNB N_B2_c_86_n 0.0325701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B2_c_87_n 0.00459177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B2_c_88_n 0.0181519f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.375
cc_9 VNB N_B1_M1006_g 0.00790407f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.655
cc_10 VNB N_B1_c_123_n 0.0276838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_c_124_n 0.00688498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_125_n 0.016922f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.375
cc_13 VNB N_A1_M1000_g 0.00820307f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.655
cc_14 VNB A1 0.00208896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A1 0.00675466f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_16 VNB N_A1_c_157_n 0.0305866f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.375
cc_17 VNB N_A1_c_158_n 0.018491f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.375
cc_18 VNB N_A2_M1002_g 0.0118262f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.655
cc_19 VNB A2 0.0163708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_c_188_n 0.0380744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_c_189_n 0.0223217f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.375
cc_22 VNB Y 0.00824409f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.375
cc_23 VNB Y 0.033727f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.375
cc_24 VNB N_Y_c_211_n 0.0283132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_305_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.702 $Y2=1.665
cc_26 VNB N_VGND_c_341_n 0.0319236f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.655
cc_27 VNB N_VGND_c_342_n 0.0110036f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_28 VNB N_VGND_c_343_n 0.0331498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_344_n 0.0414671f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.375
cc_30 VNB N_VGND_c_345_n 0.189996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_C1_M1009_g 0.0277444f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_32 VPB C1 0.0041971f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_33 VPB N_B2_M1004_g 0.0242392f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.655
cc_34 VPB N_B1_M1006_g 0.0198184f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.655
cc_35 VPB N_A1_M1000_g 0.0204935f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.655
cc_36 VPB N_A2_M1002_g 0.0258794f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.655
cc_37 VPB Y 0.0575045f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.375
cc_38 VPB N_A_110_367#_c_241_n 5.42696e-19 $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.655
cc_39 VPB N_A_110_367#_c_242_n 0.0101065f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_40 VPB N_A_110_367#_c_243_n 0.00981378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_217_367#_c_261_n 0.0082033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_217_367#_c_262_n 0.00405719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_217_367#_c_263_n 0.00482627f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.375
cc_44 VPB N_A_217_367#_c_264_n 0.0142475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_217_367#_c_265_n 0.0456129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_217_367#_c_266_n 0.00936055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_306_n 0.00561478f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.655
cc_48 VPB N_VPWR_c_307_n 0.0622309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_308_n 0.018397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_305_n 0.0478867f $X=-0.19 $Y=1.655 $X2=0.702 $Y2=1.665
cc_51 VPB N_VPWR_c_310_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 C1 N_B2_M1004_g 0.00465343f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_53 N_C1_c_55_n N_B2_M1004_g 7.10275e-19 $X=0.71 $Y=1.375 $X2=0 $Y2=0
cc_54 N_C1_M1007_g N_B2_c_86_n 5.86767e-19 $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_55 C1 N_B2_c_86_n 3.09009e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_56 N_C1_c_55_n N_B2_c_86_n 0.0144832f $X=0.71 $Y=1.375 $X2=0 $Y2=0
cc_57 N_C1_M1007_g N_B2_c_87_n 2.39145e-19 $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_58 C1 N_B2_c_87_n 0.0242626f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_59 N_C1_c_55_n N_B2_c_87_n 0.00211217f $X=0.71 $Y=1.375 $X2=0 $Y2=0
cc_60 N_C1_M1007_g N_B2_c_88_n 0.0115045f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_61 N_C1_M1007_g N_Y_c_213_n 0.011219f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_62 C1 N_Y_c_213_n 0.0188061f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_63 N_C1_c_55_n N_Y_c_213_n 0.00143628f $X=0.71 $Y=1.375 $X2=0 $Y2=0
cc_64 N_C1_c_55_n Y 0.00536922f $X=0.71 $Y=1.375 $X2=0 $Y2=0
cc_65 N_C1_M1007_g Y 0.00572998f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_66 C1 Y 0.0420544f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_C1_c_55_n Y 0.0199747f $X=0.71 $Y=1.375 $X2=0 $Y2=0
cc_68 N_C1_M1009_g N_A_110_367#_c_241_n 0.00158305f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_69 N_C1_M1009_g N_A_110_367#_c_242_n 0.0100324f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_70 C1 N_A_110_367#_c_242_n 0.0252511f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_C1_c_55_n N_A_110_367#_c_242_n 0.0013635f $X=0.71 $Y=1.375 $X2=0 $Y2=0
cc_72 N_C1_M1009_g N_A_217_367#_c_261_n 0.00176212f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_73 N_C1_M1009_g N_A_217_367#_c_263_n 0.00240065f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_74 C1 N_A_217_367#_c_263_n 0.00373682f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_75 N_C1_M1009_g N_VPWR_c_307_n 0.00577794f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_76 N_C1_M1009_g N_VPWR_c_305_n 0.0128129f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_77 N_C1_M1007_g N_VGND_c_341_n 0.0189419f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_78 N_C1_M1007_g N_VGND_c_345_n 0.00560729f $X=0.64 $Y=0.655 $X2=0 $Y2=0
cc_79 N_B2_M1004_g N_B1_M1006_g 0.0273523f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_80 N_B2_c_86_n N_B1_c_123_n 0.0438154f $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_81 N_B2_c_87_n N_B1_c_123_n 3.79323e-19 $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_82 N_B2_c_86_n N_B1_c_124_n 0.00224248f $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_83 N_B2_c_87_n N_B1_c_124_n 0.0251034f $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_84 N_B2_c_88_n N_B1_c_125_n 0.0438154f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_85 N_B2_c_86_n N_Y_c_213_n 0.00458327f $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_86 N_B2_c_87_n N_Y_c_213_n 0.0248671f $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_87 N_B2_c_88_n N_Y_c_213_n 0.0159922f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_88 N_B2_c_87_n Y 7.68718e-19 $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_89 N_B2_M1004_g N_A_110_367#_c_242_n 0.00501976f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_90 N_B2_M1004_g N_A_110_367#_c_243_n 0.0135436f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B2_M1004_g N_A_217_367#_c_261_n 0.016092f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_92 N_B2_M1004_g N_A_217_367#_c_262_n 0.0145899f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_93 N_B2_c_87_n N_A_217_367#_c_262_n 9.48869e-19 $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_94 N_B2_M1004_g N_A_217_367#_c_263_n 0.00338675f $X=1.425 $Y=2.465 $X2=0
+ $Y2=0
cc_95 N_B2_c_86_n N_A_217_367#_c_263_n 0.00484319f $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_96 N_B2_c_87_n N_A_217_367#_c_263_n 0.025882f $X=1.305 $Y=1.35 $X2=0 $Y2=0
cc_97 N_B2_M1004_g N_VPWR_c_307_n 0.00357877f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_98 N_B2_M1004_g N_VPWR_c_305_n 0.00682391f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_99 N_B2_c_88_n N_VGND_c_341_n 0.016016f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_100 N_B2_c_88_n N_VGND_c_344_n 0.00487821f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_101 N_B2_c_88_n N_VGND_c_345_n 0.00446189f $X=1.32 $Y=1.185 $X2=0 $Y2=0
cc_102 N_B1_M1006_g N_A1_M1000_g 0.0225583f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_103 N_B1_c_123_n A1 5.08372e-19 $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_104 N_B1_c_124_n A1 0.0165393f $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_105 N_B1_c_123_n N_A1_c_157_n 0.0209094f $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_106 N_B1_c_124_n N_A1_c_157_n 0.00110396f $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_107 N_B1_c_125_n N_A1_c_158_n 0.0104861f $X=1.875 $Y=1.185 $X2=0 $Y2=0
cc_108 N_B1_c_123_n N_Y_c_213_n 0.00369942f $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_109 N_B1_c_124_n N_Y_c_213_n 0.0291437f $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_110 N_B1_c_125_n N_Y_c_213_n 0.00965217f $X=1.875 $Y=1.185 $X2=0 $Y2=0
cc_111 N_B1_M1006_g N_A_217_367#_c_261_n 6.30568e-19 $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_112 N_B1_M1006_g N_A_217_367#_c_262_n 0.0131834f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_B1_c_123_n N_A_217_367#_c_262_n 0.00233882f $X=1.875 $Y=1.35 $X2=0
+ $Y2=0
cc_114 N_B1_c_124_n N_A_217_367#_c_262_n 0.0268196f $X=1.875 $Y=1.35 $X2=0 $Y2=0
cc_115 N_B1_M1006_g N_A_217_367#_c_266_n 0.00171833f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_B1_c_123_n N_A_217_367#_c_266_n 0.00207565f $X=1.875 $Y=1.35 $X2=0
+ $Y2=0
cc_117 N_B1_c_124_n N_A_217_367#_c_266_n 0.00694405f $X=1.875 $Y=1.35 $X2=0
+ $Y2=0
cc_118 N_B1_M1006_g N_VPWR_c_307_n 0.00585385f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B1_M1006_g N_VPWR_c_305_n 0.0109797f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B1_c_125_n N_VGND_c_341_n 0.00247173f $X=1.875 $Y=1.185 $X2=0 $Y2=0
cc_121 N_B1_c_125_n N_VGND_c_344_n 0.00585385f $X=1.875 $Y=1.185 $X2=0 $Y2=0
cc_122 N_B1_c_125_n N_VGND_c_345_n 0.00656731f $X=1.875 $Y=1.185 $X2=0 $Y2=0
cc_123 N_A1_M1000_g N_A2_M1002_g 0.0208882f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_124 A1 A2 0.0268327f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A1_c_157_n A2 2.56847e-19 $X=2.415 $Y=1.35 $X2=0 $Y2=0
cc_126 A1 N_A2_c_188_n 0.0048404f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A1_c_157_n N_A2_c_188_n 0.0205208f $X=2.415 $Y=1.35 $X2=0 $Y2=0
cc_128 A1 N_A2_c_189_n 0.0048404f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_129 N_A1_c_158_n N_A2_c_189_n 0.0254131f $X=2.415 $Y=1.185 $X2=0 $Y2=0
cc_130 N_A1_M1000_g N_A_217_367#_c_264_n 0.0161443f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_131 A1 N_A_217_367#_c_264_n 0.0307689f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A1_c_157_n N_A_217_367#_c_264_n 0.00142157f $X=2.415 $Y=1.35 $X2=0
+ $Y2=0
cc_133 N_A1_c_157_n N_A_217_367#_c_266_n 9.47052e-19 $X=2.415 $Y=1.35 $X2=0
+ $Y2=0
cc_134 N_A1_M1000_g N_VPWR_c_306_n 0.00353208f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A1_M1000_g N_VPWR_c_307_n 0.00585385f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A1_M1000_g N_VPWR_c_305_n 0.01087f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A1_c_158_n N_VGND_c_343_n 0.00145663f $X=2.415 $Y=1.185 $X2=0 $Y2=0
cc_138 A1 N_VGND_c_344_n 0.0135178f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_139 N_A1_c_158_n N_VGND_c_344_n 0.00585385f $X=2.415 $Y=1.185 $X2=0 $Y2=0
cc_140 A1 N_VGND_c_345_n 0.0106004f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_141 N_A1_c_158_n N_VGND_c_345_n 0.0114286f $X=2.415 $Y=1.185 $X2=0 $Y2=0
cc_142 A1 A_480_47# 0.0135102f $X=2.555 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_143 N_A2_M1002_g N_A_217_367#_c_264_n 0.0195273f $X=2.865 $Y=2.465 $X2=0
+ $Y2=0
cc_144 A2 N_A_217_367#_c_264_n 0.0259924f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_145 N_A2_c_188_n N_A_217_367#_c_264_n 0.00492355f $X=2.99 $Y=1.35 $X2=0 $Y2=0
cc_146 N_A2_M1002_g N_VPWR_c_306_n 0.00346341f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A2_M1002_g N_VPWR_c_308_n 0.00585385f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A2_M1002_g N_VPWR_c_305_n 0.0117069f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_149 A2 N_VGND_c_343_n 0.0248549f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_150 N_A2_c_188_n N_VGND_c_343_n 0.00483488f $X=2.99 $Y=1.35 $X2=0 $Y2=0
cc_151 N_A2_c_189_n N_VGND_c_343_n 0.0181765f $X=2.972 $Y=1.185 $X2=0 $Y2=0
cc_152 N_A2_c_189_n N_VGND_c_344_n 0.00486043f $X=2.972 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A2_c_189_n N_VGND_c_345_n 0.00864313f $X=2.972 $Y=1.185 $X2=0 $Y2=0
cc_154 Y N_A_217_367#_c_263_n 0.00350867f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_155 Y N_VPWR_c_307_n 0.0188791f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_156 N_Y_M1009_s N_VPWR_c_305_n 0.00302127f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_157 Y N_VPWR_c_305_n 0.0110024f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_158 N_Y_c_213_n N_VGND_M1007_d 0.0172577f $X=1.89 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_159 N_Y_c_213_n N_VGND_c_341_n 0.0449705f $X=1.89 $Y=0.93 $X2=0 $Y2=0
cc_160 N_Y_c_211_n N_VGND_c_341_n 0.0282017f $X=0.425 $Y=0.43 $X2=0 $Y2=0
cc_161 N_Y_c_234_p N_VGND_c_344_n 0.0212513f $X=2.055 $Y=0.38 $X2=0 $Y2=0
cc_162 N_Y_M1007_s N_VGND_c_345_n 0.00244073f $X=0.3 $Y=0.235 $X2=0 $Y2=0
cc_163 N_Y_M1003_d N_VGND_c_345_n 0.00436037f $X=1.86 $Y=0.235 $X2=0 $Y2=0
cc_164 N_Y_c_213_n N_VGND_c_345_n 0.0227645f $X=1.89 $Y=0.93 $X2=0 $Y2=0
cc_165 N_Y_c_234_p N_VGND_c_345_n 0.0127519f $X=2.055 $Y=0.38 $X2=0 $Y2=0
cc_166 N_Y_c_211_n N_VGND_c_345_n 0.0165607f $X=0.425 $Y=0.43 $X2=0 $Y2=0
cc_167 N_Y_c_213_n A_300_47# 0.00298885f $X=1.89 $Y=0.93 $X2=-0.19 $Y2=-0.245
cc_168 N_A_110_367#_c_243_n N_A_217_367#_M1004_s 0.00495471f $X=1.545 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_169 N_A_110_367#_c_242_n N_A_217_367#_c_261_n 0.0624615f $X=0.69 $Y=2.085
+ $X2=0 $Y2=0
cc_170 N_A_110_367#_c_243_n N_A_217_367#_c_261_n 0.0205857f $X=1.545 $Y=2.99
+ $X2=0 $Y2=0
cc_171 N_A_110_367#_M1004_d N_A_217_367#_c_262_n 0.00197722f $X=1.5 $Y=1.835
+ $X2=0 $Y2=0
cc_172 N_A_110_367#_c_254_p N_A_217_367#_c_262_n 0.0151327f $X=1.64 $Y=2.21
+ $X2=0 $Y2=0
cc_173 N_A_110_367#_c_241_n N_VPWR_c_307_n 0.0197904f $X=0.7 $Y=2.905 $X2=0
+ $Y2=0
cc_174 N_A_110_367#_c_243_n N_VPWR_c_307_n 0.0555856f $X=1.545 $Y=2.99 $X2=0
+ $Y2=0
cc_175 N_A_110_367#_M1009_d N_VPWR_c_305_n 0.00215158f $X=0.55 $Y=1.835 $X2=0
+ $Y2=0
cc_176 N_A_110_367#_M1004_d N_VPWR_c_305_n 0.00305741f $X=1.5 $Y=1.835 $X2=0
+ $Y2=0
cc_177 N_A_110_367#_c_241_n N_VPWR_c_305_n 0.0119513f $X=0.7 $Y=2.905 $X2=0
+ $Y2=0
cc_178 N_A_110_367#_c_243_n N_VPWR_c_305_n 0.0343175f $X=1.545 $Y=2.99 $X2=0
+ $Y2=0
cc_179 N_A_217_367#_c_264_n N_VPWR_M1000_d 0.00261503f $X=2.975 $Y=1.79
+ $X2=-0.19 $Y2=1.655
cc_180 N_A_217_367#_c_264_n N_VPWR_c_306_n 0.0200142f $X=2.975 $Y=1.79 $X2=0
+ $Y2=0
cc_181 N_A_217_367#_c_298_p N_VPWR_c_307_n 0.0188066f $X=2.09 $Y=1.98 $X2=0
+ $Y2=0
cc_182 N_A_217_367#_c_265_n N_VPWR_c_308_n 0.0181659f $X=3.08 $Y=1.98 $X2=0
+ $Y2=0
cc_183 N_A_217_367#_M1004_s N_VPWR_c_305_n 0.0021598f $X=1.085 $Y=1.835 $X2=0
+ $Y2=0
cc_184 N_A_217_367#_M1006_d N_VPWR_c_305_n 0.00298555f $X=1.95 $Y=1.835 $X2=0
+ $Y2=0
cc_185 N_A_217_367#_M1002_d N_VPWR_c_305_n 0.00336915f $X=2.94 $Y=1.835 $X2=0
+ $Y2=0
cc_186 N_A_217_367#_c_298_p N_VPWR_c_305_n 0.0123631f $X=2.09 $Y=1.98 $X2=0
+ $Y2=0
cc_187 N_A_217_367#_c_265_n N_VPWR_c_305_n 0.0104192f $X=3.08 $Y=1.98 $X2=0
+ $Y2=0
cc_188 N_VGND_c_345_n A_300_47# 0.00309736f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_189 N_VGND_c_345_n A_480_47# 0.00692346f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
