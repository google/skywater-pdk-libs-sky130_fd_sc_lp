* File: sky130_fd_sc_lp__a21boi_m.pxi.spice
* Created: Fri Aug 28 09:50:29 2020
* 
x_PM_SKY130_FD_SC_LP__A21BOI_M%B1_N N_B1_N_M1005_g N_B1_N_M1002_g N_B1_N_c_64_n
+ N_B1_N_c_65_n B1_N B1_N B1_N B1_N N_B1_N_c_67_n
+ PM_SKY130_FD_SC_LP__A21BOI_M%B1_N
x_PM_SKY130_FD_SC_LP__A21BOI_M%A_27_535# N_A_27_535#_M1002_s N_A_27_535#_M1005_s
+ N_A_27_535#_c_100_n N_A_27_535#_M1003_g N_A_27_535#_c_102_n
+ N_A_27_535#_c_103_n N_A_27_535#_M1004_g N_A_27_535#_c_104_n N_A_27_535#_c_98_n
+ N_A_27_535#_c_106_n N_A_27_535#_c_107_n N_A_27_535#_c_108_n
+ N_A_27_535#_c_109_n N_A_27_535#_c_99_n N_A_27_535#_c_110_n
+ PM_SKY130_FD_SC_LP__A21BOI_M%A_27_535#
x_PM_SKY130_FD_SC_LP__A21BOI_M%A1 N_A1_M1007_g N_A1_M1000_g N_A1_c_163_n
+ N_A1_c_164_n N_A1_c_165_n N_A1_c_170_n A1 A1 A1 N_A1_c_167_n
+ PM_SKY130_FD_SC_LP__A21BOI_M%A1
x_PM_SKY130_FD_SC_LP__A21BOI_M%A2 N_A2_M1001_g N_A2_M1006_g N_A2_c_212_n
+ N_A2_c_213_n N_A2_c_214_n A2 A2 N_A2_c_216_n PM_SKY130_FD_SC_LP__A21BOI_M%A2
x_PM_SKY130_FD_SC_LP__A21BOI_M%VPWR N_VPWR_M1005_d N_VPWR_M1000_d N_VPWR_c_246_n
+ N_VPWR_c_247_n VPWR N_VPWR_c_248_n N_VPWR_c_249_n N_VPWR_c_250_n
+ N_VPWR_c_245_n N_VPWR_c_252_n N_VPWR_c_253_n PM_SKY130_FD_SC_LP__A21BOI_M%VPWR
x_PM_SKY130_FD_SC_LP__A21BOI_M%Y N_Y_M1003_d N_Y_M1004_s Y Y Y Y Y N_Y_c_278_n
+ PM_SKY130_FD_SC_LP__A21BOI_M%Y
x_PM_SKY130_FD_SC_LP__A21BOI_M%A_306_395# N_A_306_395#_M1004_d
+ N_A_306_395#_M1006_d N_A_306_395#_c_304_n N_A_306_395#_c_300_n
+ N_A_306_395#_c_301_n N_A_306_395#_c_302_n
+ PM_SKY130_FD_SC_LP__A21BOI_M%A_306_395#
x_PM_SKY130_FD_SC_LP__A21BOI_M%VGND N_VGND_M1002_d N_VGND_M1001_d N_VGND_c_318_n
+ N_VGND_c_319_n N_VGND_c_320_n N_VGND_c_321_n VGND N_VGND_c_322_n
+ N_VGND_c_323_n N_VGND_c_324_n N_VGND_c_325_n PM_SKY130_FD_SC_LP__A21BOI_M%VGND
cc_1 VNB N_B1_N_M1005_g 0.00996229f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_2 VNB N_B1_N_M1002_g 0.0220539f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.445
cc_3 VNB N_B1_N_c_64_n 0.0236573f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.31
cc_4 VNB N_B1_N_c_65_n 0.0166859f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.475
cc_5 VNB B1_N 0.00869537f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_B1_N_c_67_n 0.0165065f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.97
cc_7 VNB N_A_27_535#_M1003_g 0.0605319f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.31
cc_8 VNB N_A_27_535#_c_98_n 0.0487111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_535#_c_99_n 0.0157146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_M1007_g 0.0193875f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_11 VNB N_A1_c_163_n 0.0269299f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_12 VNB N_A1_c_164_n 0.0310206f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_A1_c_165_n 0.0118757f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_14 VNB A1 0.00542901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_167_n 0.0211758f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=0.925
cc_16 VNB N_A2_M1006_g 0.0183199f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.445
cc_17 VNB N_A2_c_212_n 0.022671f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.97
cc_18 VNB N_A2_c_213_n 0.0342966f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.805
cc_19 VNB N_A2_c_214_n 0.0214226f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.475
cc_20 VNB A2 0.00872245f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_21 VNB N_A2_c_216_n 0.0360713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_245_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.665
cc_23 VNB N_Y_c_278_n 0.0085167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_318_n 0.00494119f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.97
cc_25 VNB N_VGND_c_319_n 0.0127533f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_26 VNB N_VGND_c_320_n 0.0219539f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_27 VNB N_VGND_c_321_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_322_n 0.032694f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=0.925
cc_29 VNB N_VGND_c_323_n 0.016145f $X=-0.19 $Y=-0.245 $X2=0.642 $Y2=1.665
cc_30 VNB N_VGND_c_324_n 0.184179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_325_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_B1_N_M1005_g 0.0727613f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_33 VPB B1_N 0.00793107f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_34 VPB N_A_27_535#_c_100_n 0.0458526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_27_535#_M1003_g 0.00368347f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.31
cc_36 VPB N_A_27_535#_c_102_n 0.025683f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_37 VPB N_A_27_535#_c_103_n 0.0194964f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_38 VPB N_A_27_535#_c_104_n 0.0113524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_27_535#_c_98_n 0.0397337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_27_535#_c_106_n 0.0114303f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.97
cc_41 VPB N_A_27_535#_c_107_n 0.0217221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_27_535#_c_108_n 0.00450053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_27_535#_c_109_n 0.0514736f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.665
cc_44 VPB N_A_27_535#_c_110_n 0.0092115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A1_M1000_g 0.0187104f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.31
cc_46 VPB N_A1_c_165_n 0.00126055f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_47 VPB N_A1_c_170_n 0.0120679f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_48 VPB N_A2_M1006_g 0.0378274f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.445
cc_49 VPB N_VPWR_c_246_n 0.00580306f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.97
cc_50 VPB N_VPWR_c_247_n 0.0452113f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_51 VPB N_VPWR_c_248_n 0.0153607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_249_n 0.0319085f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=0.97
cc_53 VPB N_VPWR_c_250_n 0.0217138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_245_n 0.0889962f $X=-0.19 $Y=1.655 $X2=0.642 $Y2=1.665
cc_55 VPB N_VPWR_c_252_n 0.00510247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_253_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_278_n 0.00239236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_306_395#_c_300_n 0.0269913f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.31
cc_59 VPB N_A_306_395#_c_301_n 0.00279087f $X=-0.19 $Y=1.655 $X2=0.565 $Y2=1.475
cc_60 VPB N_A_306_395#_c_302_n 4.08405e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_61 N_B1_N_M1005_g N_A_27_535#_M1003_g 0.00542971f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_62 N_B1_N_M1002_g N_A_27_535#_M1003_g 0.0162922f $X=0.615 $Y=0.445 $X2=0
+ $Y2=0
cc_63 B1_N N_A_27_535#_M1003_g 0.00713803f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_64 N_B1_N_c_67_n N_A_27_535#_M1003_g 0.0333234f $X=0.565 $Y=0.97 $X2=0 $Y2=0
cc_65 N_B1_N_M1005_g N_A_27_535#_c_104_n 0.04127f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_66 B1_N N_A_27_535#_c_104_n 0.00443312f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_67 N_B1_N_M1002_g N_A_27_535#_c_98_n 0.00523038f $X=0.615 $Y=0.445 $X2=0
+ $Y2=0
cc_68 B1_N N_A_27_535#_c_98_n 0.0944364f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_69 N_B1_N_c_67_n N_A_27_535#_c_98_n 0.0436603f $X=0.565 $Y=0.97 $X2=0 $Y2=0
cc_70 N_B1_N_M1005_g N_A_27_535#_c_106_n 3.57552e-19 $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_71 N_B1_N_M1005_g N_A_27_535#_c_107_n 0.0162981f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_72 B1_N N_A_27_535#_c_107_n 0.0151654f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_73 N_B1_N_M1005_g N_A_27_535#_c_108_n 0.00129025f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_74 B1_N N_A_27_535#_c_99_n 9.79197e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_75 N_B1_N_c_67_n N_A_27_535#_c_99_n 0.00367103f $X=0.565 $Y=0.97 $X2=0 $Y2=0
cc_76 N_B1_N_M1005_g N_VPWR_c_246_n 0.0122587f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_77 N_B1_N_M1005_g N_VPWR_c_248_n 0.0035715f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_78 N_B1_N_M1005_g N_VPWR_c_245_n 0.00525749f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_79 N_B1_N_M1005_g N_Y_c_278_n 5.63317e-19 $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_80 N_B1_N_M1002_g N_Y_c_278_n 0.00110146f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_81 B1_N N_Y_c_278_n 0.0655899f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_82 N_B1_N_c_67_n N_Y_c_278_n 6.23168e-19 $X=0.565 $Y=0.97 $X2=0 $Y2=0
cc_83 N_B1_N_M1002_g N_VGND_c_318_n 0.00288714f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_84 B1_N N_VGND_c_318_n 0.00413949f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_85 N_B1_N_M1002_g N_VGND_c_320_n 0.00585385f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_86 N_B1_N_M1002_g N_VGND_c_324_n 0.00733776f $X=0.615 $Y=0.445 $X2=0 $Y2=0
cc_87 B1_N N_VGND_c_324_n 0.00787983f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A_27_535#_M1003_g N_A1_M1007_g 0.0423641f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_27_535#_c_102_n N_A1_M1000_g 0.0155406f $X=1.38 $Y=1.79 $X2=0 $Y2=0
cc_90 N_A_27_535#_c_102_n N_A1_c_164_n 0.00958878f $X=1.38 $Y=1.79 $X2=0 $Y2=0
cc_91 N_A_27_535#_M1003_g N_A1_c_165_n 0.00277151f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_27_535#_c_102_n N_A1_c_170_n 0.00659532f $X=1.38 $Y=1.79 $X2=0 $Y2=0
cc_93 N_A_27_535#_M1003_g A1 6.87401e-19 $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_27_535#_c_107_n N_VPWR_c_246_n 0.0218865f $X=1.055 $Y=2.58 $X2=0 $Y2=0
cc_95 N_A_27_535#_c_108_n N_VPWR_c_246_n 0.01471f $X=1.14 $Y=2.9 $X2=0 $Y2=0
cc_96 N_A_27_535#_c_109_n N_VPWR_c_246_n 0.00230183f $X=1.14 $Y=2.9 $X2=0 $Y2=0
cc_97 N_A_27_535#_c_103_n N_VPWR_c_247_n 0.00114726f $X=1.455 $Y=1.865 $X2=0
+ $Y2=0
cc_98 N_A_27_535#_c_109_n N_VPWR_c_247_n 0.00851036f $X=1.14 $Y=2.9 $X2=0 $Y2=0
cc_99 N_A_27_535#_c_106_n N_VPWR_c_248_n 0.00938235f $X=0.26 $Y=2.82 $X2=0 $Y2=0
cc_100 N_A_27_535#_c_107_n N_VPWR_c_248_n 0.00283061f $X=1.055 $Y=2.58 $X2=0
+ $Y2=0
cc_101 N_A_27_535#_c_107_n N_VPWR_c_249_n 0.00312446f $X=1.055 $Y=2.58 $X2=0
+ $Y2=0
cc_102 N_A_27_535#_c_108_n N_VPWR_c_249_n 0.0106099f $X=1.14 $Y=2.9 $X2=0 $Y2=0
cc_103 N_A_27_535#_c_109_n N_VPWR_c_249_n 0.00851942f $X=1.14 $Y=2.9 $X2=0 $Y2=0
cc_104 N_A_27_535#_M1005_s N_VPWR_c_245_n 0.00243592f $X=0.135 $Y=2.675 $X2=0
+ $Y2=0
cc_105 N_A_27_535#_c_103_n N_VPWR_c_245_n 0.00391649f $X=1.455 $Y=1.865 $X2=0
+ $Y2=0
cc_106 N_A_27_535#_c_106_n N_VPWR_c_245_n 0.00786677f $X=0.26 $Y=2.82 $X2=0
+ $Y2=0
cc_107 N_A_27_535#_c_107_n N_VPWR_c_245_n 0.0112972f $X=1.055 $Y=2.58 $X2=0
+ $Y2=0
cc_108 N_A_27_535#_c_108_n N_VPWR_c_245_n 0.00636614f $X=1.14 $Y=2.9 $X2=0 $Y2=0
cc_109 N_A_27_535#_c_109_n N_VPWR_c_245_n 0.00846221f $X=1.14 $Y=2.9 $X2=0 $Y2=0
cc_110 N_A_27_535#_c_100_n N_Y_c_278_n 0.00578666f $X=0.965 $Y=2.735 $X2=0 $Y2=0
cc_111 N_A_27_535#_M1003_g N_Y_c_278_n 0.029005f $X=1.045 $Y=0.445 $X2=0 $Y2=0
cc_112 N_A_27_535#_c_102_n N_Y_c_278_n 0.014068f $X=1.38 $Y=1.79 $X2=0 $Y2=0
cc_113 N_A_27_535#_c_103_n N_Y_c_278_n 0.00227289f $X=1.455 $Y=1.865 $X2=0 $Y2=0
cc_114 N_A_27_535#_c_104_n N_Y_c_278_n 0.00210135f $X=1.005 $Y=1.79 $X2=0 $Y2=0
cc_115 N_A_27_535#_c_107_n N_Y_c_278_n 0.00847719f $X=1.055 $Y=2.58 $X2=0 $Y2=0
cc_116 N_A_27_535#_c_109_n N_Y_c_278_n 0.00317058f $X=1.14 $Y=2.9 $X2=0 $Y2=0
cc_117 N_A_27_535#_c_102_n N_A_306_395#_c_301_n 0.00170609f $X=1.38 $Y=1.79
+ $X2=0 $Y2=0
cc_118 N_A_27_535#_M1003_g N_VGND_c_318_n 0.00288714f $X=1.045 $Y=0.445 $X2=0
+ $Y2=0
cc_119 N_A_27_535#_c_99_n N_VGND_c_320_n 0.0194396f $X=0.4 $Y=0.46 $X2=0 $Y2=0
cc_120 N_A_27_535#_M1003_g N_VGND_c_322_n 0.00579368f $X=1.045 $Y=0.445 $X2=0
+ $Y2=0
cc_121 N_A_27_535#_M1002_s N_VGND_c_324_n 0.00239077f $X=0.275 $Y=0.235 $X2=0
+ $Y2=0
cc_122 N_A_27_535#_M1003_g N_VGND_c_324_n 0.010503f $X=1.045 $Y=0.445 $X2=0
+ $Y2=0
cc_123 N_A_27_535#_c_99_n N_VGND_c_324_n 0.0139896f $X=0.4 $Y=0.46 $X2=0 $Y2=0
cc_124 N_A1_c_164_n N_A2_M1006_g 0.0107311f $X=1.66 $Y=1.475 $X2=0 $Y2=0
cc_125 N_A1_c_170_n N_A2_M1006_g 0.0234765f $X=1.865 $Y=1.825 $X2=0 $Y2=0
cc_126 N_A1_M1007_g N_A2_c_212_n 0.0171954f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_127 A1 N_A2_c_212_n 0.00673296f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_128 A1 N_A2_c_213_n 4.30154e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_129 N_A1_c_167_n N_A2_c_213_n 0.00708471f $X=1.61 $Y=0.97 $X2=0 $Y2=0
cc_130 N_A1_c_163_n N_A2_c_214_n 0.00660442f $X=1.66 $Y=1.325 $X2=0 $Y2=0
cc_131 N_A1_c_164_n N_A2_c_214_n 0.00709584f $X=1.66 $Y=1.475 $X2=0 $Y2=0
cc_132 N_A1_c_164_n A2 8.76006e-19 $X=1.66 $Y=1.475 $X2=0 $Y2=0
cc_133 A1 A2 0.0324539f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_134 N_A1_c_167_n A2 0.00335245f $X=1.61 $Y=0.97 $X2=0 $Y2=0
cc_135 A1 N_A2_c_216_n 5.79128e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 N_A1_c_167_n N_A2_c_216_n 0.00660442f $X=1.61 $Y=0.97 $X2=0 $Y2=0
cc_137 N_A1_M1000_g N_VPWR_c_247_n 0.00829547f $X=1.885 $Y=2.185 $X2=0 $Y2=0
cc_138 N_A1_M1000_g N_VPWR_c_245_n 0.00328986f $X=1.885 $Y=2.185 $X2=0 $Y2=0
cc_139 N_A1_M1007_g N_Y_c_278_n 0.00684912f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A1_c_165_n N_Y_c_278_n 0.00444961f $X=1.865 $Y=1.675 $X2=0 $Y2=0
cc_141 N_A1_c_170_n N_Y_c_278_n 3.86745e-19 $X=1.865 $Y=1.825 $X2=0 $Y2=0
cc_142 A1 N_Y_c_278_n 0.0651874f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A1_M1000_g N_A_306_395#_c_304_n 2.03427e-19 $X=1.885 $Y=2.185 $X2=0
+ $Y2=0
cc_144 N_A1_M1000_g N_A_306_395#_c_300_n 0.0105187f $X=1.885 $Y=2.185 $X2=0
+ $Y2=0
cc_145 N_A1_c_164_n N_A_306_395#_c_300_n 2.62232e-19 $X=1.66 $Y=1.475 $X2=0
+ $Y2=0
cc_146 N_A1_c_170_n N_A_306_395#_c_300_n 0.00953289f $X=1.865 $Y=1.825 $X2=0
+ $Y2=0
cc_147 A1 N_A_306_395#_c_300_n 4.2263e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_148 N_A1_c_164_n N_A_306_395#_c_301_n 0.00131472f $X=1.66 $Y=1.475 $X2=0
+ $Y2=0
cc_149 A1 N_A_306_395#_c_301_n 0.0102699f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_150 N_A1_M1007_g N_VGND_c_319_n 0.00190464f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_151 A1 N_VGND_c_319_n 6.59889e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_152 N_A1_M1007_g N_VGND_c_322_n 0.00555499f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_153 A1 N_VGND_c_322_n 0.00608199f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_154 N_A1_M1007_g N_VGND_c_324_n 0.0104275f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_155 A1 N_VGND_c_324_n 0.00800989f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_156 N_A1_c_167_n N_VGND_c_324_n 2.85386e-19 $X=1.61 $Y=0.97 $X2=0 $Y2=0
cc_157 A1 A_310_47# 0.00488416f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_158 N_A2_M1006_g N_VPWR_c_247_n 0.0143932f $X=2.315 $Y=2.185 $X2=0 $Y2=0
cc_159 N_A2_M1006_g N_VPWR_c_245_n 0.00328986f $X=2.315 $Y=2.185 $X2=0 $Y2=0
cc_160 N_A2_M1006_g N_A_306_395#_c_300_n 0.0165654f $X=2.315 $Y=2.185 $X2=0
+ $Y2=0
cc_161 N_A2_c_214_n N_A_306_395#_c_300_n 0.00305181f $X=2.295 $Y=1.435 $X2=0
+ $Y2=0
cc_162 A2 N_A_306_395#_c_300_n 0.0134753f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_163 N_A2_M1006_g N_A_306_395#_c_302_n 3.52891e-19 $X=2.315 $Y=2.185 $X2=0
+ $Y2=0
cc_164 N_A2_c_212_n N_VGND_c_319_n 0.0113371f $X=2.222 $Y=0.765 $X2=0 $Y2=0
cc_165 N_A2_c_213_n N_VGND_c_319_n 0.00403872f $X=2.222 $Y=0.915 $X2=0 $Y2=0
cc_166 A2 N_VGND_c_319_n 0.0124432f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_167 N_A2_c_212_n N_VGND_c_322_n 0.00486043f $X=2.222 $Y=0.765 $X2=0 $Y2=0
cc_168 N_A2_c_213_n N_VGND_c_323_n 3.8682e-19 $X=2.222 $Y=0.915 $X2=0 $Y2=0
cc_169 N_A2_c_212_n N_VGND_c_324_n 0.00765364f $X=2.222 $Y=0.765 $X2=0 $Y2=0
cc_170 N_A2_c_213_n N_VGND_c_324_n 5.54654e-19 $X=2.222 $Y=0.915 $X2=0 $Y2=0
cc_171 A2 N_VGND_c_324_n 0.00245938f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_172 N_VPWR_c_247_n N_A_306_395#_c_300_n 0.0207154f $X=2.1 $Y=2.25 $X2=0 $Y2=0
cc_173 N_Y_c_278_n N_A_306_395#_c_304_n 5.51287e-19 $X=1.26 $Y=0.43 $X2=0 $Y2=0
cc_174 N_Y_c_278_n N_A_306_395#_c_301_n 0.0119339f $X=1.26 $Y=0.43 $X2=0 $Y2=0
cc_175 N_Y_c_278_n N_VGND_c_322_n 0.0131352f $X=1.26 $Y=0.43 $X2=0 $Y2=0
cc_176 N_Y_M1003_d N_VGND_c_324_n 0.00415099f $X=1.12 $Y=0.235 $X2=0 $Y2=0
cc_177 N_Y_c_278_n N_VGND_c_324_n 0.00872539f $X=1.26 $Y=0.43 $X2=0 $Y2=0
cc_178 N_VGND_c_324_n A_310_47# 0.0112623f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
