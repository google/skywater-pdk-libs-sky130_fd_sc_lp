* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or2_4 A B VGND VNB VPB VPWR X
M1000 VPWR a_27_367# X VPB phighvt w=1.26e+06u l=150000u
+  ad=1.2222e+12p pd=9.5e+06u as=7.056e+11p ps=6.16e+06u
M1001 X a_27_367# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=9.66e+11p ps=9.02e+06u
M1002 X a_27_367# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_367# B VGND VNB nshort w=840000u l=150000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1004 VPWR a_27_367# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_27_367# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_27_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_27_367# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A a_27_367# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_110_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1010 X a_27_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_110_367# B a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends
