* File: sky130_fd_sc_lp__a21o_0.spice
* Created: Fri Aug 28 09:50:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21o_0.pex.spice"
.subckt sky130_fd_sc_lp__a21o_0  VNB VPB B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_80_275#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0714 AS=0.1113 PD=0.76 PS=1.37 NRD=9.996 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_80_275#_M1002_d N_B1_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07245 AS=0.0714 PD=0.765 PS=0.76 NRD=2.856 NRS=7.14 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 A_405_47# N_A1_M1004_g N_A_80_275#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.07245 PD=0.66 PS=0.765 NRD=18.564 NRS=15.708 M=1 R=2.8
+ SA=75001.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_405_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_80_275#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_A_319_473#_M1000_d N_B1_M1000_g N_A_80_275#_M1000_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_319_473#_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_319_473#_M1001_d N_A2_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
c_66 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a21o_0.pxi.spice"
*
.ends
*
*
