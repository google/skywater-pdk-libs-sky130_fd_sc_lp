* File: sky130_fd_sc_lp__a32oi_1.spice
* Created: Fri Aug 28 10:01:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a32oi_1  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1006 A_141_69# N_B2_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84 AD=0.0945
+ AS=0.2226 PD=1.065 PS=2.21 NRD=8.208 NRS=0 M=1 R=5.6 SA=75000.2 SB=75002.2
+ A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g A_141_69# VNB NSHORT L=0.15 W=0.84 AD=0.168
+ AS=0.0945 PD=1.24 PS=1.065 NRD=6.42 NRS=8.208 M=1 R=5.6 SA=75000.6 SB=75001.9
+ A=0.126 P=1.98 MULT=1
MM1001 A_326_69# N_A1_M1001_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.168 PD=1.23 PS=1.24 NRD=19.992 NRS=10.704 M=1 R=5.6 SA=75001.1 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1008 A_434_69# N_A2_M1008_g A_326_69# VNB NSHORT L=0.15 W=0.84 AD=0.1848
+ AS=0.1638 PD=1.28 PS=1.23 NRD=23.568 NRS=19.992 M=1 R=5.6 SA=75001.7
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A3_M1009_g A_434_69# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1848 PD=2.21 PS=1.28 NRD=0 NRS=23.568 M=1 R=5.6 SA=75002.2 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g N_A_58_367#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1002 N_A_58_367#_M1002_d N_B1_M1002_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.21735 AS=0.1764 PD=1.605 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_58_367#_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.21735 PD=1.88 PS=1.605 NRD=0 NRS=3.9006 M=1 R=8.4 SA=75001.1
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1007 N_A_58_367#_M1007_d N_A2_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3906 PD=1.54 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A3_M1003_g N_A_58_367#_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a32oi_1.pxi.spice"
*
.ends
*
*
