* File: sky130_fd_sc_lp__o32a_4.pxi.spice
* Created: Fri Aug 28 11:17:33 2020
* 
x_PM_SKY130_FD_SC_LP__O32A_4%A2 N_A2_M1012_g N_A2_M1013_g N_A2_M1018_g
+ N_A2_M1015_g N_A2_c_147_n N_A2_c_138_n N_A2_c_139_n N_A2_c_140_n A2 A2 A2
+ N_A2_c_141_n N_A2_c_142_n N_A2_c_143_n N_A2_c_144_n
+ PM_SKY130_FD_SC_LP__O32A_4%A2
x_PM_SKY130_FD_SC_LP__O32A_4%A1 N_A1_c_228_n N_A1_M1006_g N_A1_M1002_g
+ N_A1_c_230_n N_A1_M1019_g N_A1_M1024_g A1 N_A1_c_233_n
+ PM_SKY130_FD_SC_LP__O32A_4%A1
x_PM_SKY130_FD_SC_LP__O32A_4%A3 N_A3_c_281_n N_A3_M1017_g N_A3_M1005_g
+ N_A3_M1025_g N_A3_c_284_n N_A3_M1022_g A3 A3 A3 N_A3_c_286_n
+ PM_SKY130_FD_SC_LP__O32A_4%A3
x_PM_SKY130_FD_SC_LP__O32A_4%B2 N_B2_M1003_g N_B2_c_335_n N_B2_M1014_g
+ N_B2_M1026_g N_B2_M1023_g N_B2_c_337_n N_B2_c_345_n B2 B2 N_B2_c_339_n
+ N_B2_c_340_n N_B2_c_348_n PM_SKY130_FD_SC_LP__O32A_4%B2
x_PM_SKY130_FD_SC_LP__O32A_4%B1 N_B1_c_431_n N_B1_M1008_g N_B1_M1001_g
+ N_B1_c_433_n N_B1_M1021_g N_B1_M1010_g B1 N_B1_c_436_n
+ PM_SKY130_FD_SC_LP__O32A_4%B1
x_PM_SKY130_FD_SC_LP__O32A_4%A_547_367# N_A_547_367#_M1003_s
+ N_A_547_367#_M1021_d N_A_547_367#_M1005_d N_A_547_367#_M1014_d
+ N_A_547_367#_M1026_d N_A_547_367#_M1000_g N_A_547_367#_M1004_g
+ N_A_547_367#_M1007_g N_A_547_367#_M1011_g N_A_547_367#_M1009_g
+ N_A_547_367#_M1016_g N_A_547_367#_M1020_g N_A_547_367#_M1027_g
+ N_A_547_367#_c_504_n N_A_547_367#_c_503_n N_A_547_367#_c_497_n
+ N_A_547_367#_c_498_n N_A_547_367#_c_499_n N_A_547_367#_c_516_n
+ N_A_547_367#_c_521_n N_A_547_367#_c_488_n N_A_547_367#_c_500_n
+ N_A_547_367#_c_489_n N_A_547_367#_c_588_p N_A_547_367#_c_490_n
+ N_A_547_367#_c_491_n N_A_547_367#_c_492_n
+ PM_SKY130_FD_SC_LP__O32A_4%A_547_367#
x_PM_SKY130_FD_SC_LP__O32A_4%A_112_367# N_A_112_367#_M1013_s
+ N_A_112_367#_M1015_s N_A_112_367#_M1025_s N_A_112_367#_c_643_n
+ N_A_112_367#_c_644_n N_A_112_367#_c_651_n N_A_112_367#_c_682_p
+ N_A_112_367#_c_645_n N_A_112_367#_c_646_n N_A_112_367#_c_647_n
+ PM_SKY130_FD_SC_LP__O32A_4%A_112_367#
x_PM_SKY130_FD_SC_LP__O32A_4%A_195_367# N_A_195_367#_M1013_d
+ N_A_195_367#_M1024_s N_A_195_367#_c_693_n N_A_195_367#_c_694_n
+ N_A_195_367#_c_697_n N_A_195_367#_c_695_n N_A_195_367#_c_696_n
+ PM_SKY130_FD_SC_LP__O32A_4%A_195_367#
x_PM_SKY130_FD_SC_LP__O32A_4%VPWR N_VPWR_M1002_d N_VPWR_M1001_s N_VPWR_M1004_d
+ N_VPWR_M1011_d N_VPWR_M1027_d N_VPWR_c_714_n N_VPWR_c_715_n N_VPWR_c_716_n
+ N_VPWR_c_717_n N_VPWR_c_718_n N_VPWR_c_719_n N_VPWR_c_720_n VPWR
+ N_VPWR_c_721_n N_VPWR_c_722_n N_VPWR_c_723_n N_VPWR_c_724_n N_VPWR_c_725_n
+ N_VPWR_c_726_n N_VPWR_c_727_n N_VPWR_c_728_n N_VPWR_c_713_n VPWR
+ PM_SKY130_FD_SC_LP__O32A_4%VPWR
x_PM_SKY130_FD_SC_LP__O32A_4%A_823_367# N_A_823_367#_M1014_s
+ N_A_823_367#_M1010_d N_A_823_367#_c_830_n N_A_823_367#_c_831_n
+ N_A_823_367#_c_834_n N_A_823_367#_c_832_n N_A_823_367#_c_833_n
+ PM_SKY130_FD_SC_LP__O32A_4%A_823_367#
x_PM_SKY130_FD_SC_LP__O32A_4%X N_X_M1000_d N_X_M1009_d N_X_M1004_s N_X_M1016_s
+ N_X_c_903_p N_X_c_889_n N_X_c_850_n N_X_c_851_n N_X_c_856_n N_X_c_857_n
+ N_X_c_904_p N_X_c_893_n N_X_c_852_n N_X_c_858_n N_X_c_853_n N_X_c_859_n X X
+ N_X_c_854_n X PM_SKY130_FD_SC_LP__O32A_4%X
x_PM_SKY130_FD_SC_LP__O32A_4%A_44_65# N_A_44_65#_M1012_s N_A_44_65#_M1006_s
+ N_A_44_65#_M1018_s N_A_44_65#_M1022_s N_A_44_65#_M1008_s N_A_44_65#_M1023_d
+ N_A_44_65#_c_909_n N_A_44_65#_c_910_n N_A_44_65#_c_911_n N_A_44_65#_c_912_n
+ N_A_44_65#_c_925_n N_A_44_65#_c_913_n N_A_44_65#_c_914_n N_A_44_65#_c_942_n
+ N_A_44_65#_c_915_n N_A_44_65#_c_916_n N_A_44_65#_c_917_n N_A_44_65#_c_918_n
+ N_A_44_65#_c_932_n N_A_44_65#_c_919_n PM_SKY130_FD_SC_LP__O32A_4%A_44_65#
x_PM_SKY130_FD_SC_LP__O32A_4%VGND N_VGND_M1012_d N_VGND_M1019_d N_VGND_M1017_d
+ N_VGND_M1000_s N_VGND_M1007_s N_VGND_M1020_s N_VGND_c_996_n N_VGND_c_997_n
+ N_VGND_c_998_n N_VGND_c_999_n N_VGND_c_1000_n N_VGND_c_1001_n N_VGND_c_1002_n
+ N_VGND_c_1003_n N_VGND_c_1004_n N_VGND_c_1005_n VGND N_VGND_c_1006_n
+ N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n
+ N_VGND_c_1011_n N_VGND_c_1012_n N_VGND_c_1013_n VGND
+ PM_SKY130_FD_SC_LP__O32A_4%VGND
cc_1 VNB N_A2_M1012_g 0.0291361f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.745
cc_2 VNB N_A2_M1015_g 0.00245046f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=2.465
cc_3 VNB N_A2_c_138_n 0.00125274f $X=-0.19 $Y=-0.245 $X2=2.095 $Y2=1.695
cc_4 VNB N_A2_c_139_n 0.00559934f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.44
cc_5 VNB N_A2_c_140_n 0.0289083f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.44
cc_6 VNB N_A2_c_141_n 0.0398266f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.51
cc_7 VNB N_A2_c_142_n 0.0170694f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.275
cc_8 VNB N_A2_c_143_n 0.0189522f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.645
cc_9 VNB N_A2_c_144_n 0.00135233f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.645
cc_10 VNB N_A1_c_228_n 0.0188073f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.345
cc_11 VNB N_A1_M1002_g 0.00228976f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=2.465
cc_12 VNB N_A1_c_230_n 0.0161722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1024_g 0.00262668f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=2.465
cc_14 VNB A1 0.00216792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_233_n 0.037186f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.402
cc_16 VNB N_A3_c_281_n 0.0165829f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.345
cc_17 VNB N_A3_M1005_g 0.00257133f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=2.465
cc_18 VNB N_A3_M1025_g 0.00316601f $X=-0.19 $Y=-0.245 $X2=2.19 $Y2=0.745
cc_19 VNB N_A3_c_284_n 0.0178494f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=1.605
cc_20 VNB A3 0.0214869f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.78
cc_21 VNB N_A3_c_286_n 0.0621853f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_B2_M1003_g 0.0241088f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.745
cc_23 VNB N_B2_c_335_n 0.0274082f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.675
cc_24 VNB N_B2_M1023_g 0.0235626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B2_c_337_n 0.00258189f $X=-0.19 $Y=-0.245 $X2=2.095 $Y2=1.695
cc_26 VNB B2 0.00267707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B2_c_339_n 0.0294176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B2_c_340_n 0.00172422f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.51
cc_29 VNB N_B1_c_431_n 0.0167813f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.345
cc_30 VNB N_B1_M1001_g 0.00242759f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=2.465
cc_31 VNB N_B1_c_433_n 0.0159372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B1_M1010_g 0.00228995f $X=-0.19 $Y=-0.245 $X2=2.23 $Y2=2.465
cc_33 VNB B1 0.00253508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B1_c_436_n 0.0368743f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.402
cc_35 VNB N_A_547_367#_M1000_g 0.0271933f $X=-0.19 $Y=-0.245 $X2=2.095 $Y2=1.535
cc_36 VNB N_A_547_367#_M1007_g 0.0214062f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_37 VNB N_A_547_367#_M1009_g 0.0213918f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.51
cc_38 VNB N_A_547_367#_M1020_g 0.025885f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.645
cc_39 VNB N_A_547_367#_c_488_n 0.0259177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_547_367#_c_489_n 0.00120004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_547_367#_c_490_n 0.0022501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_547_367#_c_491_n 0.0026564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_547_367#_c_492_n 0.0734879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VPWR_c_713_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_850_n 0.00313892f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.44
cc_46 VNB N_X_c_851_n 0.00245786f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.44
cc_47 VNB N_X_c_852_n 0.00152954f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.51
cc_48 VNB N_X_c_853_n 0.00134924f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.605
cc_49 VNB N_X_c_854_n 0.00990216f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.645
cc_50 VNB X 0.0221686f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.645
cc_51 VNB N_A_44_65#_c_909_n 0.0316346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_44_65#_c_910_n 0.00485698f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.44
cc_53 VNB N_A_44_65#_c_911_n 0.00989965f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.44
cc_54 VNB N_A_44_65#_c_912_n 0.00307647f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_55 VNB N_A_44_65#_c_913_n 8.83459e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_44_65#_c_914_n 0.00236116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_44_65#_c_915_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.605
cc_58 VNB N_A_44_65#_c_916_n 0.00620266f $X=-0.19 $Y=-0.245 $X2=1.11 $Y2=1.645
cc_59 VNB N_A_44_65#_c_917_n 0.00726481f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.645
cc_60 VNB N_A_44_65#_c_918_n 0.00447203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_44_65#_c_919_n 0.00181812f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.645
cc_62 VNB N_VGND_c_996_n 0.00187549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_997_n 0.0023483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_998_n 0.00957225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_999_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1000_n 0.0113984f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=1.51
cc_67 VNB N_VGND_c_1001_n 0.0281524f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.51
cc_68 VNB N_VGND_c_1002_n 0.015575f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.275
cc_69 VNB N_VGND_c_1003_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.605
cc_70 VNB N_VGND_c_1004_n 0.015687f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.645
cc_71 VNB N_VGND_c_1005_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1006_n 0.0188967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1007_n 0.0678798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1008_n 0.0131655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1009_n 0.0131655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1010_n 0.0184917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1011_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1012_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1013_n 0.428881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VPB N_A2_M1013_g 0.0225139f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=2.465
cc_81 VPB N_A2_M1015_g 0.0198913f $X=-0.19 $Y=1.655 $X2=2.23 $Y2=2.465
cc_82 VPB N_A2_c_147_n 0.00581175f $X=-0.19 $Y=1.655 $X2=2.01 $Y2=1.78
cc_83 VPB N_A2_c_138_n 3.75592e-19 $X=-0.19 $Y=1.655 $X2=2.095 $Y2=1.695
cc_84 VPB N_A2_c_141_n 0.0115904f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.51
cc_85 VPB N_A2_c_143_n 0.0274631f $X=-0.19 $Y=1.655 $X2=1.11 $Y2=1.645
cc_86 VPB N_A1_M1002_g 0.0182888f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=2.465
cc_87 VPB N_A1_M1024_g 0.0189655f $X=-0.19 $Y=1.655 $X2=2.23 $Y2=2.465
cc_88 VPB N_A3_M1005_g 0.01884f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=2.465
cc_89 VPB N_A3_M1025_g 0.0240313f $X=-0.19 $Y=1.655 $X2=2.19 $Y2=0.745
cc_90 VPB N_B2_c_335_n 0.00666273f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=1.675
cc_91 VPB N_B2_M1014_g 0.0225298f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=2.465
cc_92 VPB N_B2_M1026_g 0.0225139f $X=-0.19 $Y=1.655 $X2=2.19 $Y2=0.745
cc_93 VPB N_B2_c_337_n 7.29158e-19 $X=-0.19 $Y=1.655 $X2=2.095 $Y2=1.695
cc_94 VPB N_B2_c_345_n 0.00157844f $X=-0.19 $Y=1.655 $X2=2.21 $Y2=1.44
cc_95 VPB B2 0.00141562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_B2_c_339_n 0.0076529f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_B2_c_348_n 0.00587864f $X=-0.19 $Y=1.655 $X2=2.21 $Y2=1.275
cc_98 VPB N_B1_M1001_g 0.0184996f $X=-0.19 $Y=1.655 $X2=0.9 $Y2=2.465
cc_99 VPB N_B1_M1010_g 0.0182889f $X=-0.19 $Y=1.655 $X2=2.23 $Y2=2.465
cc_100 VPB N_A_547_367#_M1004_g 0.0233894f $X=-0.19 $Y=1.655 $X2=2.21 $Y2=1.402
cc_101 VPB N_A_547_367#_M1011_g 0.0188565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_547_367#_M1016_g 0.0188421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_547_367#_M1027_g 0.0224142f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.645
cc_104 VPB N_A_547_367#_c_497_n 0.0104809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_547_367#_c_498_n 0.00239269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_547_367#_c_499_n 0.00671935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_547_367#_c_500_n 0.0102356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_547_367#_c_489_n 0.0248435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_547_367#_c_492_n 0.00700947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_112_367#_c_643_n 0.00744706f $X=-0.19 $Y=1.655 $X2=2.19 $Y2=0.745
cc_111 VPB N_A_112_367#_c_644_n 0.0326198f $X=-0.19 $Y=1.655 $X2=2.23 $Y2=1.605
cc_112 VPB N_A_112_367#_c_645_n 0.00698181f $X=-0.19 $Y=1.655 $X2=2.21 $Y2=1.44
cc_113 VPB N_A_112_367#_c_646_n 0.00396063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_112_367#_c_647_n 0.00890434f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_115 VPB N_VPWR_c_714_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=2.095 $Y2=1.535
cc_116 VPB N_VPWR_c_715_n 0.0684818f $X=-0.19 $Y=1.655 $X2=2.095 $Y2=1.402
cc_117 VPB N_VPWR_c_716_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=2.21 $Y2=1.44
cc_118 VPB N_VPWR_c_717_n 0.0105962f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_119 VPB N_VPWR_c_718_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.51
cc_120 VPB N_VPWR_c_719_n 0.0112967f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=1.51
cc_121 VPB N_VPWR_c_720_n 0.0415885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_721_n 0.040076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_722_n 0.0298666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_723_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_724_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_725_n 0.00436966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_726_n 0.00436966f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_727_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_728_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_713_n 0.0778481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_X_c_856_n 0.00304705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_X_c_857_n 0.00206601f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_133 VPB N_X_c_858_n 0.0111105f $X=-0.19 $Y=1.655 $X2=2.21 $Y2=1.44
cc_134 VPB N_X_c_859_n 0.00144314f $X=-0.19 $Y=1.655 $X2=1.11 $Y2=1.645
cc_135 VPB X 0.00514909f $X=-0.19 $Y=1.655 $X2=1.33 $Y2=1.645
cc_136 N_A2_M1012_g N_A1_c_228_n 0.0088679f $X=0.56 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_137 N_A2_M1013_g N_A1_M1002_g 0.0262268f $X=0.9 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A2_c_147_n N_A1_M1002_g 0.00630129f $X=2.01 $Y=1.78 $X2=0 $Y2=0
cc_139 N_A2_c_144_n N_A1_M1002_g 0.0073685f $X=1.33 $Y=1.645 $X2=0 $Y2=0
cc_140 N_A2_c_139_n N_A1_c_230_n 0.00167845f $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_141 N_A2_c_142_n N_A1_c_230_n 0.0317022f $X=2.21 $Y=1.275 $X2=0 $Y2=0
cc_142 N_A2_M1015_g N_A1_M1024_g 0.0328418f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A2_c_147_n N_A1_M1024_g 0.0107543f $X=2.01 $Y=1.78 $X2=0 $Y2=0
cc_144 N_A2_c_144_n N_A1_M1024_g 4.73352e-19 $X=1.33 $Y=1.645 $X2=0 $Y2=0
cc_145 N_A2_c_147_n A1 0.0241477f $X=2.01 $Y=1.78 $X2=0 $Y2=0
cc_146 N_A2_c_139_n A1 0.0194663f $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_147 N_A2_c_140_n A1 2.89248e-19 $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_148 N_A2_c_141_n A1 4.16167e-19 $X=0.9 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A2_c_142_n A1 3.78166e-19 $X=2.21 $Y=1.275 $X2=0 $Y2=0
cc_150 N_A2_c_144_n A1 0.00790265f $X=1.33 $Y=1.645 $X2=0 $Y2=0
cc_151 N_A2_c_147_n N_A1_c_233_n 0.00249657f $X=2.01 $Y=1.78 $X2=0 $Y2=0
cc_152 N_A2_c_138_n N_A1_c_233_n 0.00331626f $X=2.095 $Y=1.695 $X2=0 $Y2=0
cc_153 N_A2_c_140_n N_A1_c_233_n 0.0215394f $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_154 N_A2_c_141_n N_A1_c_233_n 0.0262268f $X=0.9 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A2_c_144_n N_A1_c_233_n 0.00960231f $X=1.33 $Y=1.645 $X2=0 $Y2=0
cc_156 N_A2_c_142_n N_A3_c_281_n 0.0160601f $X=2.21 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A2_M1015_g N_A3_M1005_g 0.0216345f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A2_c_139_n A3 0.0215073f $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_159 N_A2_c_140_n A3 9.96297e-19 $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_160 N_A2_c_142_n A3 0.0014569f $X=2.21 $Y=1.275 $X2=0 $Y2=0
cc_161 N_A2_c_138_n N_A3_c_286_n 7.94424e-19 $X=2.095 $Y=1.695 $X2=0 $Y2=0
cc_162 N_A2_c_139_n N_A3_c_286_n 3.02283e-19 $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_163 N_A2_c_140_n N_A3_c_286_n 0.0221274f $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_164 N_A2_M1015_g N_A_547_367#_c_503_n 2.58097e-19 $X=2.23 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A2_c_143_n N_A_112_367#_M1013_s 0.00231902f $X=1.11 $Y=1.645 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A2_c_141_n N_A_112_367#_c_643_n 0.00129419f $X=0.9 $Y=1.51 $X2=0 $Y2=0
cc_167 N_A2_c_143_n N_A_112_367#_c_643_n 0.0216939f $X=1.11 $Y=1.645 $X2=0 $Y2=0
cc_168 N_A2_M1013_g N_A_112_367#_c_651_n 0.0121823f $X=0.9 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A2_M1015_g N_A_112_367#_c_651_n 0.0140682f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A2_c_147_n N_A_112_367#_c_651_n 0.00851944f $X=2.01 $Y=1.78 $X2=0 $Y2=0
cc_171 N_A2_c_139_n N_A_112_367#_c_651_n 0.00433722f $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_172 N_A2_c_140_n N_A_112_367#_c_651_n 3.53691e-19 $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_173 N_A2_c_143_n N_A_112_367#_c_651_n 0.065158f $X=1.11 $Y=1.645 $X2=0 $Y2=0
cc_174 N_A2_M1015_g N_A_112_367#_c_646_n 0.00106565f $X=2.23 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A2_c_147_n N_A_112_367#_c_646_n 0.0128113f $X=2.01 $Y=1.78 $X2=0 $Y2=0
cc_176 N_A2_c_139_n N_A_112_367#_c_646_n 0.00207697f $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_177 N_A2_c_140_n N_A_112_367#_c_646_n 6.34049e-19 $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_178 N_A2_c_143_n N_A_195_367#_M1013_d 8.44873e-19 $X=1.11 $Y=1.645 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A2_c_144_n N_A_195_367#_M1013_d 9.65569e-19 $X=1.33 $Y=1.645 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A2_c_147_n N_A_195_367#_M1024_s 0.00219084f $X=2.01 $Y=1.78 $X2=0 $Y2=0
cc_181 N_A2_M1013_g N_A_195_367#_c_693_n 0.00215206f $X=0.9 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A2_M1013_g N_A_195_367#_c_694_n 0.0067084f $X=0.9 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A2_M1015_g N_A_195_367#_c_695_n 0.00205939f $X=2.23 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A2_M1015_g N_A_195_367#_c_696_n 0.0062009f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A2_c_147_n N_VPWR_M1002_d 0.00176891f $X=2.01 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_186 N_A2_M1013_g N_VPWR_c_714_n 0.00109224f $X=0.9 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A2_M1015_g N_VPWR_c_714_n 0.00103397f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A2_M1015_g N_VPWR_c_715_n 0.0054895f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A2_M1013_g N_VPWR_c_721_n 0.0054895f $X=0.9 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A2_M1013_g N_VPWR_c_713_n 0.0112379f $X=0.9 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A2_M1015_g N_VPWR_c_713_n 0.0100572f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A2_M1012_g N_A_44_65#_c_909_n 0.00354524f $X=0.56 $Y=0.745 $X2=0 $Y2=0
cc_193 N_A2_M1012_g N_A_44_65#_c_910_n 0.0153173f $X=0.56 $Y=0.745 $X2=0 $Y2=0
cc_194 N_A2_c_141_n N_A_44_65#_c_910_n 0.00902477f $X=0.9 $Y=1.51 $X2=0 $Y2=0
cc_195 N_A2_c_143_n N_A_44_65#_c_910_n 0.0556322f $X=1.11 $Y=1.645 $X2=0 $Y2=0
cc_196 N_A2_c_143_n N_A_44_65#_c_911_n 0.0234831f $X=1.11 $Y=1.645 $X2=0 $Y2=0
cc_197 N_A2_c_147_n N_A_44_65#_c_925_n 0.00424227f $X=2.01 $Y=1.78 $X2=0 $Y2=0
cc_198 N_A2_c_139_n N_A_44_65#_c_925_n 0.0145527f $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_199 N_A2_c_140_n N_A_44_65#_c_925_n 3.1276e-19 $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_200 N_A2_c_142_n N_A_44_65#_c_925_n 0.0128646f $X=2.21 $Y=1.275 $X2=0 $Y2=0
cc_201 N_A2_M1012_g N_A_44_65#_c_913_n 0.00283898f $X=0.56 $Y=0.745 $X2=0 $Y2=0
cc_202 N_A2_c_147_n N_A_44_65#_c_913_n 0.00368571f $X=2.01 $Y=1.78 $X2=0 $Y2=0
cc_203 N_A2_c_144_n N_A_44_65#_c_913_n 0.0140692f $X=1.33 $Y=1.645 $X2=0 $Y2=0
cc_204 N_A2_c_139_n N_A_44_65#_c_932_n 0.00402648f $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_205 N_A2_c_140_n N_A_44_65#_c_932_n 4.48278e-19 $X=2.21 $Y=1.44 $X2=0 $Y2=0
cc_206 N_A2_c_142_n N_VGND_c_996_n 0.00904966f $X=2.21 $Y=1.275 $X2=0 $Y2=0
cc_207 N_A2_c_142_n N_VGND_c_997_n 4.27755e-19 $X=2.21 $Y=1.275 $X2=0 $Y2=0
cc_208 N_A2_c_142_n N_VGND_c_1004_n 0.00414769f $X=2.21 $Y=1.275 $X2=0 $Y2=0
cc_209 N_A2_M1012_g N_VGND_c_1006_n 0.00414769f $X=0.56 $Y=0.745 $X2=0 $Y2=0
cc_210 N_A2_M1012_g N_VGND_c_1010_n 0.0137422f $X=0.56 $Y=0.745 $X2=0 $Y2=0
cc_211 N_A2_M1012_g N_VGND_c_1013_n 0.00821268f $X=0.56 $Y=0.745 $X2=0 $Y2=0
cc_212 N_A2_c_142_n N_VGND_c_1013_n 0.00792084f $X=2.21 $Y=1.275 $X2=0 $Y2=0
cc_213 N_A1_M1002_g N_A_112_367#_c_651_n 0.010446f $X=1.33 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A1_M1024_g N_A_112_367#_c_651_n 0.0106711f $X=1.76 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A1_M1002_g N_A_195_367#_c_697_n 0.00959697f $X=1.33 $Y=2.465 $X2=0
+ $Y2=0
cc_216 N_A1_M1024_g N_A_195_367#_c_697_n 0.00959697f $X=1.76 $Y=2.465 $X2=0
+ $Y2=0
cc_217 N_A1_M1002_g N_VPWR_c_714_n 0.00988124f $X=1.33 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A1_M1024_g N_VPWR_c_714_n 0.00991121f $X=1.76 $Y=2.465 $X2=0 $Y2=0
cc_219 N_A1_M1024_g N_VPWR_c_715_n 0.00486043f $X=1.76 $Y=2.465 $X2=0 $Y2=0
cc_220 N_A1_M1002_g N_VPWR_c_721_n 0.00486043f $X=1.33 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A1_M1002_g N_VPWR_c_713_n 0.00445201f $X=1.33 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A1_M1024_g N_VPWR_c_713_n 0.00454571f $X=1.76 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A1_c_228_n N_A_44_65#_c_912_n 5.57288e-19 $X=1.33 $Y=1.275 $X2=0 $Y2=0
cc_224 N_A1_c_230_n N_A_44_65#_c_912_n 5.11798e-19 $X=1.76 $Y=1.275 $X2=0 $Y2=0
cc_225 N_A1_c_230_n N_A_44_65#_c_925_n 0.012781f $X=1.76 $Y=1.275 $X2=0 $Y2=0
cc_226 A1 N_A_44_65#_c_925_n 0.0121689f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_227 N_A1_c_228_n N_A_44_65#_c_913_n 0.0233099f $X=1.33 $Y=1.275 $X2=0 $Y2=0
cc_228 N_A1_c_230_n N_A_44_65#_c_913_n 9.4689e-19 $X=1.76 $Y=1.275 $X2=0 $Y2=0
cc_229 A1 N_A_44_65#_c_913_n 0.0153015f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_230 N_A1_c_233_n N_A_44_65#_c_913_n 7.92618e-19 $X=1.76 $Y=1.44 $X2=0 $Y2=0
cc_231 N_A1_c_228_n N_VGND_c_996_n 3.2514e-19 $X=1.33 $Y=1.275 $X2=0 $Y2=0
cc_232 N_A1_c_230_n N_VGND_c_996_n 0.00858106f $X=1.76 $Y=1.275 $X2=0 $Y2=0
cc_233 N_A1_c_228_n N_VGND_c_1002_n 0.00499542f $X=1.33 $Y=1.275 $X2=0 $Y2=0
cc_234 N_A1_c_230_n N_VGND_c_1002_n 0.00414769f $X=1.76 $Y=1.275 $X2=0 $Y2=0
cc_235 N_A1_c_228_n N_VGND_c_1010_n 0.00370849f $X=1.33 $Y=1.275 $X2=0 $Y2=0
cc_236 N_A1_c_228_n N_VGND_c_1013_n 0.009973f $X=1.33 $Y=1.275 $X2=0 $Y2=0
cc_237 N_A1_c_230_n N_VGND_c_1013_n 0.00787505f $X=1.76 $Y=1.275 $X2=0 $Y2=0
cc_238 N_A3_c_284_n N_B2_M1003_g 0.00818819f $X=3.11 $Y=1.255 $X2=0 $Y2=0
cc_239 A3 N_B2_M1003_g 0.00396292f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_240 N_A3_c_286_n N_B2_M1003_g 0.00196794f $X=3.11 $Y=1.43 $X2=0 $Y2=0
cc_241 N_A3_M1025_g N_B2_c_335_n 0.00130433f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_242 A3 N_B2_c_335_n 0.00169418f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_243 N_A3_c_286_n N_B2_c_335_n 0.00713542f $X=3.11 $Y=1.43 $X2=0 $Y2=0
cc_244 N_A3_M1025_g N_B2_c_337_n 7.4406e-19 $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_245 A3 N_B2_c_337_n 0.0151112f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_246 N_A3_c_286_n N_B2_c_337_n 6.55039e-19 $X=3.11 $Y=1.43 $X2=0 $Y2=0
cc_247 N_A3_M1025_g N_B2_c_345_n 8.82997e-19 $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A3_M1005_g N_A_547_367#_c_504_n 0.00193114f $X=2.66 $Y=2.465 $X2=0
+ $Y2=0
cc_249 N_A3_M1025_g N_A_547_367#_c_504_n 5.89773e-19 $X=3.09 $Y=2.465 $X2=0
+ $Y2=0
cc_250 N_A3_M1005_g N_A_547_367#_c_503_n 0.00906203f $X=2.66 $Y=2.465 $X2=0
+ $Y2=0
cc_251 N_A3_M1025_g N_A_547_367#_c_503_n 0.0113541f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_252 N_A3_M1025_g N_A_547_367#_c_497_n 0.0125611f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_253 A3 N_A_547_367#_c_498_n 0.00125331f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_254 N_A3_M1025_g N_A_547_367#_c_499_n 0.00317379f $X=3.09 $Y=2.465 $X2=0
+ $Y2=0
cc_255 N_A3_M1005_g N_A_112_367#_c_645_n 0.0134716f $X=2.66 $Y=2.465 $X2=0 $Y2=0
cc_256 N_A3_M1025_g N_A_112_367#_c_645_n 0.0148248f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_257 A3 N_A_112_367#_c_645_n 0.0701191f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_258 N_A3_c_286_n N_A_112_367#_c_645_n 0.00977896f $X=3.11 $Y=1.43 $X2=0 $Y2=0
cc_259 N_A3_M1005_g N_VPWR_c_715_n 0.00547432f $X=2.66 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A3_M1025_g N_VPWR_c_715_n 0.00357842f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A3_M1005_g N_VPWR_c_713_n 0.00990114f $X=2.66 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A3_M1025_g N_VPWR_c_713_n 0.00675085f $X=3.09 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A3_c_281_n N_A_44_65#_c_942_n 0.0131507f $X=2.66 $Y=1.275 $X2=0 $Y2=0
cc_264 N_A3_c_284_n N_A_44_65#_c_942_n 0.0157518f $X=3.11 $Y=1.255 $X2=0 $Y2=0
cc_265 A3 N_A_44_65#_c_942_n 0.0828163f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_266 N_A3_c_286_n N_A_44_65#_c_942_n 0.00222047f $X=3.11 $Y=1.43 $X2=0 $Y2=0
cc_267 N_A3_c_284_n N_A_44_65#_c_916_n 0.00183238f $X=3.11 $Y=1.255 $X2=0 $Y2=0
cc_268 N_A3_c_281_n N_VGND_c_996_n 4.47393e-19 $X=2.66 $Y=1.275 $X2=0 $Y2=0
cc_269 N_A3_c_281_n N_VGND_c_997_n 0.00774532f $X=2.66 $Y=1.275 $X2=0 $Y2=0
cc_270 N_A3_c_284_n N_VGND_c_997_n 0.00966512f $X=3.11 $Y=1.255 $X2=0 $Y2=0
cc_271 N_A3_c_281_n N_VGND_c_1004_n 0.00481374f $X=2.66 $Y=1.275 $X2=0 $Y2=0
cc_272 N_A3_c_284_n N_VGND_c_1007_n 0.00414769f $X=3.11 $Y=1.255 $X2=0 $Y2=0
cc_273 N_A3_c_281_n N_VGND_c_1013_n 0.00915999f $X=2.66 $Y=1.275 $X2=0 $Y2=0
cc_274 N_A3_c_284_n N_VGND_c_1013_n 0.00816552f $X=3.11 $Y=1.255 $X2=0 $Y2=0
cc_275 N_B2_M1003_g N_B1_c_431_n 0.0264047f $X=3.975 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_276 N_B2_M1014_g N_B1_M1001_g 0.0357457f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_277 N_B2_c_340_n N_B1_M1001_g 4.38578e-19 $X=5.165 $Y=1.645 $X2=0 $Y2=0
cc_278 N_B2_c_348_n N_B1_M1001_g 0.0111548f $X=4.945 $Y=1.645 $X2=0 $Y2=0
cc_279 N_B2_M1023_g N_B1_c_433_n 0.0221743f $X=5.34 $Y=0.745 $X2=0 $Y2=0
cc_280 N_B2_M1026_g N_B1_M1010_g 0.0261571f $X=5.335 $Y=2.465 $X2=0 $Y2=0
cc_281 N_B2_c_340_n N_B1_M1010_g 0.0058995f $X=5.165 $Y=1.645 $X2=0 $Y2=0
cc_282 N_B2_c_348_n N_B1_M1010_g 0.00862526f $X=4.945 $Y=1.645 $X2=0 $Y2=0
cc_283 N_B2_M1003_g B1 7.31524e-19 $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_284 N_B2_c_335_n B1 2.62412e-19 $X=4.04 $Y=1.675 $X2=0 $Y2=0
cc_285 N_B2_M1023_g B1 2.93177e-19 $X=5.34 $Y=0.745 $X2=0 $Y2=0
cc_286 N_B2_c_337_n B1 0.010105f $X=4.025 $Y=1.51 $X2=0 $Y2=0
cc_287 N_B2_c_339_n B1 4.34648e-19 $X=5.46 $Y=1.51 $X2=0 $Y2=0
cc_288 N_B2_c_340_n B1 0.00790265f $X=5.165 $Y=1.645 $X2=0 $Y2=0
cc_289 N_B2_c_348_n B1 0.0242978f $X=4.945 $Y=1.645 $X2=0 $Y2=0
cc_290 N_B2_c_335_n N_B1_c_436_n 0.0212374f $X=4.04 $Y=1.675 $X2=0 $Y2=0
cc_291 N_B2_c_337_n N_B1_c_436_n 0.00492383f $X=4.025 $Y=1.51 $X2=0 $Y2=0
cc_292 N_B2_c_339_n N_B1_c_436_n 0.0261571f $X=5.46 $Y=1.51 $X2=0 $Y2=0
cc_293 N_B2_c_340_n N_B1_c_436_n 0.00865548f $X=5.165 $Y=1.645 $X2=0 $Y2=0
cc_294 N_B2_c_348_n N_B1_c_436_n 0.00246333f $X=4.945 $Y=1.645 $X2=0 $Y2=0
cc_295 N_B2_c_345_n N_A_547_367#_M1014_d 9.67538e-19 $X=4.195 $Y=1.78 $X2=0
+ $Y2=0
cc_296 B2 N_A_547_367#_M1026_d 0.00204972f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_297 B2 N_A_547_367#_M1004_g 5.73789e-19 $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_298 N_B2_c_335_n N_A_547_367#_c_498_n 2.73845e-19 $X=4.04 $Y=1.675 $X2=0
+ $Y2=0
cc_299 N_B2_c_345_n N_A_547_367#_c_498_n 0.00423925f $X=4.195 $Y=1.78 $X2=0
+ $Y2=0
cc_300 N_B2_c_335_n N_A_547_367#_c_516_n 2.50349e-19 $X=4.04 $Y=1.675 $X2=0
+ $Y2=0
cc_301 N_B2_M1014_g N_A_547_367#_c_516_n 0.0122056f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_302 N_B2_M1026_g N_A_547_367#_c_516_n 0.0121823f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_B2_c_345_n N_A_547_367#_c_516_n 0.0129516f $X=4.195 $Y=1.78 $X2=0 $Y2=0
cc_304 N_B2_c_348_n N_A_547_367#_c_516_n 0.0397382f $X=4.945 $Y=1.645 $X2=0
+ $Y2=0
cc_305 N_B2_c_340_n N_A_547_367#_c_521_n 3.78713e-19 $X=5.165 $Y=1.645 $X2=0
+ $Y2=0
cc_306 N_B2_c_348_n N_A_547_367#_c_521_n 0.00501581f $X=4.945 $Y=1.645 $X2=0
+ $Y2=0
cc_307 N_B2_M1023_g N_A_547_367#_c_488_n 0.0152966f $X=5.34 $Y=0.745 $X2=0 $Y2=0
cc_308 B2 N_A_547_367#_c_488_n 0.0644802f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_309 N_B2_c_339_n N_A_547_367#_c_488_n 0.00885689f $X=5.46 $Y=1.51 $X2=0 $Y2=0
cc_310 N_B2_M1026_g N_A_547_367#_c_489_n 0.00474649f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_B2_c_339_n N_A_547_367#_c_489_n 8.8037e-19 $X=5.46 $Y=1.51 $X2=0 $Y2=0
cc_312 N_B2_c_340_n N_A_547_367#_c_489_n 0.0397382f $X=5.165 $Y=1.645 $X2=0
+ $Y2=0
cc_313 N_B2_M1003_g N_A_547_367#_c_490_n 0.0117689f $X=3.975 $Y=0.745 $X2=0
+ $Y2=0
cc_314 N_B2_c_335_n N_A_547_367#_c_490_n 0.0035384f $X=4.04 $Y=1.675 $X2=0 $Y2=0
cc_315 N_B2_c_337_n N_A_547_367#_c_490_n 0.0145004f $X=4.025 $Y=1.51 $X2=0 $Y2=0
cc_316 N_B2_c_348_n N_A_547_367#_c_490_n 0.00530838f $X=4.945 $Y=1.645 $X2=0
+ $Y2=0
cc_317 N_B2_M1023_g N_A_547_367#_c_491_n 0.0131547f $X=5.34 $Y=0.745 $X2=0 $Y2=0
cc_318 N_B2_c_340_n N_A_547_367#_c_491_n 0.0290441f $X=5.165 $Y=1.645 $X2=0
+ $Y2=0
cc_319 N_B2_c_339_n N_A_547_367#_c_492_n 0.00360915f $X=5.46 $Y=1.51 $X2=0 $Y2=0
cc_320 N_B2_M1014_g N_A_112_367#_c_645_n 0.00124012f $X=4.04 $Y=2.465 $X2=0
+ $Y2=0
cc_321 N_B2_c_345_n N_A_112_367#_c_645_n 0.00834734f $X=4.195 $Y=1.78 $X2=0
+ $Y2=0
cc_322 N_B2_M1014_g N_A_112_367#_c_647_n 0.00276429f $X=4.04 $Y=2.465 $X2=0
+ $Y2=0
cc_323 N_B2_c_348_n N_VPWR_M1001_s 0.00176891f $X=4.945 $Y=1.645 $X2=0 $Y2=0
cc_324 N_B2_M1014_g N_VPWR_c_715_n 0.0054895f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_325 N_B2_M1014_g N_VPWR_c_716_n 0.00108483f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_326 N_B2_M1026_g N_VPWR_c_716_n 0.00109224f $X=5.335 $Y=2.465 $X2=0 $Y2=0
cc_327 N_B2_M1026_g N_VPWR_c_717_n 0.00332357f $X=5.335 $Y=2.465 $X2=0 $Y2=0
cc_328 N_B2_M1026_g N_VPWR_c_722_n 0.0054895f $X=5.335 $Y=2.465 $X2=0 $Y2=0
cc_329 N_B2_M1014_g N_VPWR_c_713_n 0.01125f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_330 N_B2_M1026_g N_VPWR_c_713_n 0.0112379f $X=5.335 $Y=2.465 $X2=0 $Y2=0
cc_331 N_B2_c_345_n N_A_823_367#_M1014_s 2.41924e-19 $X=4.195 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_332 N_B2_c_348_n N_A_823_367#_M1014_s 0.00156645f $X=4.945 $Y=1.645 $X2=-0.19
+ $Y2=-0.245
cc_333 B2 N_A_823_367#_M1010_d 4.05978e-19 $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_334 N_B2_c_340_n N_A_823_367#_M1010_d 0.00140446f $X=5.165 $Y=1.645 $X2=0
+ $Y2=0
cc_335 N_B2_M1014_g N_A_823_367#_c_830_n 0.00215206f $X=4.04 $Y=2.465 $X2=0
+ $Y2=0
cc_336 N_B2_M1014_g N_A_823_367#_c_831_n 0.00640122f $X=4.04 $Y=2.465 $X2=0
+ $Y2=0
cc_337 N_B2_M1026_g N_A_823_367#_c_832_n 0.00215206f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_338 N_B2_M1026_g N_A_823_367#_c_833_n 0.00639285f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_339 N_B2_M1003_g N_A_44_65#_c_915_n 0.0128794f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_340 N_B2_M1023_g N_A_44_65#_c_917_n 0.0132987f $X=5.34 $Y=0.745 $X2=0 $Y2=0
cc_341 N_B2_M1003_g N_A_44_65#_c_919_n 3.59852e-19 $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_342 N_B2_M1023_g N_VGND_c_998_n 0.00245321f $X=5.34 $Y=0.745 $X2=0 $Y2=0
cc_343 N_B2_M1003_g N_VGND_c_1007_n 0.00302501f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_344 N_B2_M1023_g N_VGND_c_1007_n 0.00302501f $X=5.34 $Y=0.745 $X2=0 $Y2=0
cc_345 N_B2_M1003_g N_VGND_c_1013_n 0.00470833f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_346 N_B2_M1023_g N_VGND_c_1013_n 0.00486099f $X=5.34 $Y=0.745 $X2=0 $Y2=0
cc_347 N_B1_M1001_g N_A_547_367#_c_516_n 0.0104754f $X=4.475 $Y=2.465 $X2=0
+ $Y2=0
cc_348 N_B1_M1010_g N_A_547_367#_c_516_n 0.010446f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_349 N_B1_c_431_n N_A_547_367#_c_521_n 0.0126823f $X=4.475 $Y=1.275 $X2=0
+ $Y2=0
cc_350 N_B1_c_433_n N_A_547_367#_c_521_n 0.0108471f $X=4.905 $Y=1.275 $X2=0
+ $Y2=0
cc_351 B1 N_A_547_367#_c_521_n 0.0228016f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_352 N_B1_c_436_n N_A_547_367#_c_521_n 5.91533e-19 $X=4.905 $Y=1.44 $X2=0
+ $Y2=0
cc_353 N_B1_c_431_n N_A_547_367#_c_490_n 0.00353861f $X=4.475 $Y=1.275 $X2=0
+ $Y2=0
cc_354 N_B1_c_431_n N_A_547_367#_c_491_n 0.00139898f $X=4.475 $Y=1.275 $X2=0
+ $Y2=0
cc_355 N_B1_c_433_n N_A_547_367#_c_491_n 0.0102072f $X=4.905 $Y=1.275 $X2=0
+ $Y2=0
cc_356 B1 N_A_547_367#_c_491_n 0.00341102f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_357 N_B1_M1001_g N_VPWR_c_715_n 0.00486043f $X=4.475 $Y=2.465 $X2=0 $Y2=0
cc_358 N_B1_M1001_g N_VPWR_c_716_n 0.00994527f $X=4.475 $Y=2.465 $X2=0 $Y2=0
cc_359 N_B1_M1010_g N_VPWR_c_716_n 0.00994143f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_360 N_B1_M1010_g N_VPWR_c_722_n 0.00486043f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_361 N_B1_M1001_g N_VPWR_c_713_n 0.0044641f $X=4.475 $Y=2.465 $X2=0 $Y2=0
cc_362 N_B1_M1010_g N_VPWR_c_713_n 0.00445201f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_363 N_B1_M1001_g N_A_823_367#_c_834_n 0.00959697f $X=4.475 $Y=2.465 $X2=0
+ $Y2=0
cc_364 N_B1_M1010_g N_A_823_367#_c_834_n 0.00959697f $X=4.905 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_B1_c_431_n N_A_44_65#_c_915_n 0.00850882f $X=4.475 $Y=1.275 $X2=0 $Y2=0
cc_366 N_B1_c_433_n N_A_44_65#_c_917_n 0.00912207f $X=4.905 $Y=1.275 $X2=0 $Y2=0
cc_367 N_B1_c_431_n N_A_44_65#_c_919_n 0.00660963f $X=4.475 $Y=1.275 $X2=0 $Y2=0
cc_368 N_B1_c_431_n N_VGND_c_1007_n 0.00303788f $X=4.475 $Y=1.275 $X2=0 $Y2=0
cc_369 N_B1_c_433_n N_VGND_c_1007_n 0.00302501f $X=4.905 $Y=1.275 $X2=0 $Y2=0
cc_370 N_B1_c_431_n N_VGND_c_1013_n 0.00440875f $X=4.475 $Y=1.275 $X2=0 $Y2=0
cc_371 N_B1_c_433_n N_VGND_c_1013_n 0.00436111f $X=4.905 $Y=1.275 $X2=0 $Y2=0
cc_372 N_A_547_367#_c_497_n N_A_112_367#_M1025_s 0.00495471f $X=3.66 $Y=2.99
+ $X2=0 $Y2=0
cc_373 N_A_547_367#_M1005_d N_A_112_367#_c_645_n 0.00176461f $X=2.735 $Y=1.835
+ $X2=0 $Y2=0
cc_374 N_A_547_367#_c_503_n N_A_112_367#_c_645_n 0.0170777f $X=2.875 $Y=2.13
+ $X2=0 $Y2=0
cc_375 N_A_547_367#_c_497_n N_A_112_367#_c_647_n 0.0189128f $X=3.66 $Y=2.99
+ $X2=0 $Y2=0
cc_376 N_A_547_367#_c_498_n N_A_112_367#_c_647_n 0.0136671f $X=3.79 $Y=2.205
+ $X2=0 $Y2=0
cc_377 N_A_547_367#_c_499_n N_A_112_367#_c_647_n 0.0393274f $X=3.825 $Y=2.52
+ $X2=0 $Y2=0
cc_378 N_A_547_367#_c_516_n N_VPWR_M1001_s 0.00339715f $X=5.455 $Y=2.12 $X2=0
+ $Y2=0
cc_379 N_A_547_367#_c_489_n N_VPWR_M1004_d 0.00517251f $X=6.047 $Y=2.035 $X2=0
+ $Y2=0
cc_380 N_A_547_367#_c_504_n N_VPWR_c_715_n 0.01906f $X=2.875 $Y=2.905 $X2=0
+ $Y2=0
cc_381 N_A_547_367#_c_497_n N_VPWR_c_715_n 0.0555622f $X=3.66 $Y=2.99 $X2=0
+ $Y2=0
cc_382 N_A_547_367#_M1004_g N_VPWR_c_717_n 0.0146864f $X=6.365 $Y=2.465 $X2=0
+ $Y2=0
cc_383 N_A_547_367#_M1011_g N_VPWR_c_717_n 6.47957e-19 $X=6.795 $Y=2.465 $X2=0
+ $Y2=0
cc_384 N_A_547_367#_c_500_n N_VPWR_c_717_n 0.0415095f $X=5.55 $Y=2.515 $X2=0
+ $Y2=0
cc_385 N_A_547_367#_c_489_n N_VPWR_c_717_n 0.0209021f $X=6.047 $Y=2.035 $X2=0
+ $Y2=0
cc_386 N_A_547_367#_M1004_g N_VPWR_c_718_n 7.27171e-19 $X=6.365 $Y=2.465 $X2=0
+ $Y2=0
cc_387 N_A_547_367#_M1011_g N_VPWR_c_718_n 0.0142791f $X=6.795 $Y=2.465 $X2=0
+ $Y2=0
cc_388 N_A_547_367#_M1016_g N_VPWR_c_718_n 0.0142791f $X=7.225 $Y=2.465 $X2=0
+ $Y2=0
cc_389 N_A_547_367#_M1027_g N_VPWR_c_718_n 7.27171e-19 $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_390 N_A_547_367#_M1016_g N_VPWR_c_720_n 7.27171e-19 $X=7.225 $Y=2.465 $X2=0
+ $Y2=0
cc_391 N_A_547_367#_M1027_g N_VPWR_c_720_n 0.0153838f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_392 N_A_547_367#_c_500_n N_VPWR_c_722_n 0.0178111f $X=5.55 $Y=2.515 $X2=0
+ $Y2=0
cc_393 N_A_547_367#_M1004_g N_VPWR_c_723_n 0.00486043f $X=6.365 $Y=2.465 $X2=0
+ $Y2=0
cc_394 N_A_547_367#_M1011_g N_VPWR_c_723_n 0.00486043f $X=6.795 $Y=2.465 $X2=0
+ $Y2=0
cc_395 N_A_547_367#_M1016_g N_VPWR_c_724_n 0.00486043f $X=7.225 $Y=2.465 $X2=0
+ $Y2=0
cc_396 N_A_547_367#_M1027_g N_VPWR_c_724_n 0.00486043f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_A_547_367#_M1005_d N_VPWR_c_713_n 0.00223559f $X=2.735 $Y=1.835 $X2=0
+ $Y2=0
cc_398 N_A_547_367#_M1014_d N_VPWR_c_713_n 0.00368223f $X=3.7 $Y=1.835 $X2=0
+ $Y2=0
cc_399 N_A_547_367#_M1026_d N_VPWR_c_713_n 0.00371702f $X=5.41 $Y=1.835 $X2=0
+ $Y2=0
cc_400 N_A_547_367#_M1004_g N_VPWR_c_713_n 0.00824727f $X=6.365 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_A_547_367#_M1011_g N_VPWR_c_713_n 0.00824727f $X=6.795 $Y=2.465 $X2=0
+ $Y2=0
cc_402 N_A_547_367#_M1016_g N_VPWR_c_713_n 0.00824727f $X=7.225 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A_547_367#_M1027_g N_VPWR_c_713_n 0.00824727f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_404 N_A_547_367#_c_504_n N_VPWR_c_713_n 0.0124545f $X=2.875 $Y=2.905 $X2=0
+ $Y2=0
cc_405 N_A_547_367#_c_497_n N_VPWR_c_713_n 0.0328425f $X=3.66 $Y=2.99 $X2=0
+ $Y2=0
cc_406 N_A_547_367#_c_500_n N_VPWR_c_713_n 0.0100304f $X=5.55 $Y=2.515 $X2=0
+ $Y2=0
cc_407 N_A_547_367#_c_516_n N_A_823_367#_M1014_s 0.00360982f $X=5.455 $Y=2.12
+ $X2=-0.19 $Y2=-0.245
cc_408 N_A_547_367#_c_516_n N_A_823_367#_M1010_d 0.00353353f $X=5.455 $Y=2.12
+ $X2=0 $Y2=0
cc_409 N_A_547_367#_c_516_n N_A_823_367#_c_830_n 0.0158119f $X=5.455 $Y=2.12
+ $X2=0 $Y2=0
cc_410 N_A_547_367#_c_516_n N_A_823_367#_c_834_n 0.0323235f $X=5.455 $Y=2.12
+ $X2=0 $Y2=0
cc_411 N_A_547_367#_c_516_n N_A_823_367#_c_832_n 0.0154042f $X=5.455 $Y=2.12
+ $X2=0 $Y2=0
cc_412 N_A_547_367#_M1007_g N_X_c_850_n 0.0135652f $X=6.795 $Y=0.665 $X2=0 $Y2=0
cc_413 N_A_547_367#_M1009_g N_X_c_850_n 0.0138879f $X=7.225 $Y=0.665 $X2=0 $Y2=0
cc_414 N_A_547_367#_c_588_p N_X_c_850_n 0.0478398f $X=7.475 $Y=1.49 $X2=0 $Y2=0
cc_415 N_A_547_367#_c_492_n N_X_c_850_n 0.00243542f $X=7.655 $Y=1.49 $X2=0 $Y2=0
cc_416 N_A_547_367#_M1000_g N_X_c_851_n 0.00119507f $X=6.365 $Y=0.665 $X2=0
+ $Y2=0
cc_417 N_A_547_367#_c_488_n N_X_c_851_n 0.01174f $X=5.795 $Y=1.165 $X2=0 $Y2=0
cc_418 N_A_547_367#_c_588_p N_X_c_851_n 0.0146297f $X=7.475 $Y=1.49 $X2=0 $Y2=0
cc_419 N_A_547_367#_c_492_n N_X_c_851_n 0.00253619f $X=7.655 $Y=1.49 $X2=0 $Y2=0
cc_420 N_A_547_367#_M1011_g N_X_c_856_n 0.0130035f $X=6.795 $Y=2.465 $X2=0 $Y2=0
cc_421 N_A_547_367#_M1016_g N_X_c_856_n 0.0131657f $X=7.225 $Y=2.465 $X2=0 $Y2=0
cc_422 N_A_547_367#_c_588_p N_X_c_856_n 0.0471185f $X=7.475 $Y=1.49 $X2=0 $Y2=0
cc_423 N_A_547_367#_c_492_n N_X_c_856_n 0.00243542f $X=7.655 $Y=1.49 $X2=0 $Y2=0
cc_424 N_A_547_367#_M1004_g N_X_c_857_n 6.81074e-19 $X=6.365 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_547_367#_c_489_n N_X_c_857_n 0.00985754f $X=6.047 $Y=2.035 $X2=0
+ $Y2=0
cc_426 N_A_547_367#_c_588_p N_X_c_857_n 0.0154426f $X=7.475 $Y=1.49 $X2=0 $Y2=0
cc_427 N_A_547_367#_c_492_n N_X_c_857_n 0.00253619f $X=7.655 $Y=1.49 $X2=0 $Y2=0
cc_428 N_A_547_367#_M1020_g N_X_c_852_n 0.0164214f $X=7.655 $Y=0.665 $X2=0 $Y2=0
cc_429 N_A_547_367#_c_588_p N_X_c_852_n 0.00803119f $X=7.475 $Y=1.49 $X2=0 $Y2=0
cc_430 N_A_547_367#_M1027_g N_X_c_858_n 0.0156991f $X=7.655 $Y=2.465 $X2=0 $Y2=0
cc_431 N_A_547_367#_c_588_p N_X_c_858_n 0.00730993f $X=7.475 $Y=1.49 $X2=0 $Y2=0
cc_432 N_A_547_367#_c_588_p N_X_c_853_n 0.0146297f $X=7.475 $Y=1.49 $X2=0 $Y2=0
cc_433 N_A_547_367#_c_492_n N_X_c_853_n 0.00253619f $X=7.655 $Y=1.49 $X2=0 $Y2=0
cc_434 N_A_547_367#_c_588_p N_X_c_859_n 0.0154426f $X=7.475 $Y=1.49 $X2=0 $Y2=0
cc_435 N_A_547_367#_c_492_n N_X_c_859_n 0.00253619f $X=7.655 $Y=1.49 $X2=0 $Y2=0
cc_436 N_A_547_367#_M1020_g X 0.020234f $X=7.655 $Y=0.665 $X2=0 $Y2=0
cc_437 N_A_547_367#_c_588_p X 0.0155178f $X=7.475 $Y=1.49 $X2=0 $Y2=0
cc_438 N_A_547_367#_c_521_n N_A_44_65#_M1008_s 0.00332139f $X=4.955 $Y=0.955
+ $X2=0 $Y2=0
cc_439 N_A_547_367#_c_488_n N_A_44_65#_M1023_d 0.00387504f $X=5.795 $Y=1.165
+ $X2=0 $Y2=0
cc_440 N_A_547_367#_M1003_s N_A_44_65#_c_915_n 0.00250873f $X=4.05 $Y=0.325
+ $X2=0 $Y2=0
cc_441 N_A_547_367#_c_521_n N_A_44_65#_c_915_n 0.00388708f $X=4.955 $Y=0.955
+ $X2=0 $Y2=0
cc_442 N_A_547_367#_c_490_n N_A_44_65#_c_915_n 0.0193847f $X=4.19 $Y=0.68 $X2=0
+ $Y2=0
cc_443 N_A_547_367#_M1021_d N_A_44_65#_c_917_n 0.0018652f $X=4.98 $Y=0.325 $X2=0
+ $Y2=0
cc_444 N_A_547_367#_c_521_n N_A_44_65#_c_917_n 0.00396432f $X=4.955 $Y=0.955
+ $X2=0 $Y2=0
cc_445 N_A_547_367#_c_488_n N_A_44_65#_c_917_n 0.00294998f $X=5.795 $Y=1.165
+ $X2=0 $Y2=0
cc_446 N_A_547_367#_c_491_n N_A_44_65#_c_917_n 0.0152552f $X=5.12 $Y=0.7 $X2=0
+ $Y2=0
cc_447 N_A_547_367#_M1000_g N_A_44_65#_c_918_n 8.07663e-19 $X=6.365 $Y=0.665
+ $X2=0 $Y2=0
cc_448 N_A_547_367#_c_488_n N_A_44_65#_c_918_n 0.0251967f $X=5.795 $Y=1.165
+ $X2=0 $Y2=0
cc_449 N_A_547_367#_c_521_n N_A_44_65#_c_919_n 0.0147769f $X=4.955 $Y=0.955
+ $X2=0 $Y2=0
cc_450 N_A_547_367#_c_488_n N_VGND_M1000_s 0.00234883f $X=5.795 $Y=1.165 $X2=0
+ $Y2=0
cc_451 N_A_547_367#_M1000_g N_VGND_c_998_n 0.012781f $X=6.365 $Y=0.665 $X2=0
+ $Y2=0
cc_452 N_A_547_367#_M1007_g N_VGND_c_998_n 6.15775e-19 $X=6.795 $Y=0.665 $X2=0
+ $Y2=0
cc_453 N_A_547_367#_c_488_n N_VGND_c_998_n 0.0231274f $X=5.795 $Y=1.165 $X2=0
+ $Y2=0
cc_454 N_A_547_367#_c_588_p N_VGND_c_998_n 4.5251e-19 $X=7.475 $Y=1.49 $X2=0
+ $Y2=0
cc_455 N_A_547_367#_M1000_g N_VGND_c_999_n 6.19888e-19 $X=6.365 $Y=0.665 $X2=0
+ $Y2=0
cc_456 N_A_547_367#_M1007_g N_VGND_c_999_n 0.0111833f $X=6.795 $Y=0.665 $X2=0
+ $Y2=0
cc_457 N_A_547_367#_M1009_g N_VGND_c_999_n 0.0110386f $X=7.225 $Y=0.665 $X2=0
+ $Y2=0
cc_458 N_A_547_367#_M1020_g N_VGND_c_999_n 6.10117e-19 $X=7.655 $Y=0.665 $X2=0
+ $Y2=0
cc_459 N_A_547_367#_M1009_g N_VGND_c_1001_n 6.19888e-19 $X=7.225 $Y=0.665 $X2=0
+ $Y2=0
cc_460 N_A_547_367#_M1020_g N_VGND_c_1001_n 0.0121709f $X=7.655 $Y=0.665 $X2=0
+ $Y2=0
cc_461 N_A_547_367#_M1000_g N_VGND_c_1008_n 0.00477554f $X=6.365 $Y=0.665 $X2=0
+ $Y2=0
cc_462 N_A_547_367#_M1007_g N_VGND_c_1008_n 0.00477554f $X=6.795 $Y=0.665 $X2=0
+ $Y2=0
cc_463 N_A_547_367#_M1009_g N_VGND_c_1009_n 0.00477554f $X=7.225 $Y=0.665 $X2=0
+ $Y2=0
cc_464 N_A_547_367#_M1020_g N_VGND_c_1009_n 0.00477554f $X=7.655 $Y=0.665 $X2=0
+ $Y2=0
cc_465 N_A_547_367#_M1000_g N_VGND_c_1013_n 0.00825815f $X=6.365 $Y=0.665 $X2=0
+ $Y2=0
cc_466 N_A_547_367#_M1007_g N_VGND_c_1013_n 0.00825815f $X=6.795 $Y=0.665 $X2=0
+ $Y2=0
cc_467 N_A_547_367#_M1009_g N_VGND_c_1013_n 0.00825815f $X=7.225 $Y=0.665 $X2=0
+ $Y2=0
cc_468 N_A_547_367#_M1020_g N_VGND_c_1013_n 0.00825815f $X=7.655 $Y=0.665 $X2=0
+ $Y2=0
cc_469 N_A_112_367#_c_651_n N_A_195_367#_M1013_d 0.00353353f $X=2.35 $Y=2.12
+ $X2=-0.19 $Y2=1.655
cc_470 N_A_112_367#_c_651_n N_A_195_367#_M1024_s 0.0043084f $X=2.35 $Y=2.12
+ $X2=0 $Y2=0
cc_471 N_A_112_367#_c_651_n N_A_195_367#_c_693_n 0.0154042f $X=2.35 $Y=2.12
+ $X2=0 $Y2=0
cc_472 N_A_112_367#_c_651_n N_A_195_367#_c_697_n 0.0323235f $X=2.35 $Y=2.12
+ $X2=0 $Y2=0
cc_473 N_A_112_367#_c_651_n N_A_195_367#_c_695_n 0.0186241f $X=2.35 $Y=2.12
+ $X2=0 $Y2=0
cc_474 N_A_112_367#_c_651_n N_VPWR_M1002_d 0.00339715f $X=2.35 $Y=2.12 $X2=-0.19
+ $Y2=1.655
cc_475 N_A_112_367#_c_682_p N_VPWR_c_715_n 0.0124525f $X=2.445 $Y=2.45 $X2=0
+ $Y2=0
cc_476 N_A_112_367#_c_644_n N_VPWR_c_721_n 0.0167395f $X=0.685 $Y=2.52 $X2=0
+ $Y2=0
cc_477 N_A_112_367#_M1013_s N_VPWR_c_713_n 0.00371907f $X=0.56 $Y=1.835 $X2=0
+ $Y2=0
cc_478 N_A_112_367#_M1015_s N_VPWR_c_713_n 0.00536646f $X=2.305 $Y=1.835 $X2=0
+ $Y2=0
cc_479 N_A_112_367#_M1025_s N_VPWR_c_713_n 0.0021598f $X=3.165 $Y=1.835 $X2=0
+ $Y2=0
cc_480 N_A_112_367#_c_644_n N_VPWR_c_713_n 0.00998284f $X=0.685 $Y=2.52 $X2=0
+ $Y2=0
cc_481 N_A_112_367#_c_682_p N_VPWR_c_713_n 0.00730901f $X=2.445 $Y=2.45 $X2=0
+ $Y2=0
cc_482 N_A_112_367#_c_646_n N_A_44_65#_c_932_n 0.00541874f $X=2.54 $Y=1.79 $X2=0
+ $Y2=0
cc_483 N_A_195_367#_c_697_n N_VPWR_M1002_d 0.00350137f $X=1.88 $Y=2.46 $X2=0.56
+ $Y2=1.345
cc_484 N_A_195_367#_c_697_n N_VPWR_c_714_n 0.0166559f $X=1.88 $Y=2.46 $X2=2.095
+ $Y2=1.535
cc_485 N_A_195_367#_c_696_n N_VPWR_c_715_n 0.0185348f $X=2.015 $Y=2.91 $X2=2.095
+ $Y2=1.402
cc_486 N_A_195_367#_c_694_n N_VPWR_c_721_n 0.0157163f $X=1.115 $Y=2.91 $X2=0
+ $Y2=0
cc_487 N_A_195_367#_M1013_d N_VPWR_c_713_n 0.00248313f $X=0.975 $Y=1.835 $X2=0
+ $Y2=0
cc_488 N_A_195_367#_M1024_s N_VPWR_c_713_n 0.0028048f $X=1.835 $Y=1.835 $X2=0
+ $Y2=0
cc_489 N_A_195_367#_c_694_n N_VPWR_c_713_n 0.00985509f $X=1.115 $Y=2.91 $X2=0
+ $Y2=0
cc_490 N_A_195_367#_c_697_n N_VPWR_c_713_n 0.0115403f $X=1.88 $Y=2.46 $X2=0
+ $Y2=0
cc_491 N_A_195_367#_c_696_n N_VPWR_c_713_n 0.0114114f $X=2.015 $Y=2.91 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_713_n N_A_823_367#_M1014_s 0.00252334f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_493 N_VPWR_c_713_n N_A_823_367#_M1010_d 0.00248313f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_715_n N_A_823_367#_c_831_n 0.0160686f $X=4.525 $Y=3.33 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_713_n N_A_823_367#_c_831_n 0.0100496f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_M1001_s N_A_823_367#_c_834_n 0.00350137f $X=4.55 $Y=1.835 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_716_n N_A_823_367#_c_834_n 0.0166559f $X=4.69 $Y=2.835 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_713_n N_A_823_367#_c_834_n 0.0115403f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_722_n N_A_823_367#_c_833_n 0.0157163f $X=5.985 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_713_n N_A_823_367#_c_833_n 0.00985509f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_713_n N_X_M1004_s 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_502 N_VPWR_c_713_n N_X_M1016_s 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_503 N_VPWR_c_723_n N_X_c_889_n 0.0124525f $X=6.845 $Y=3.33 $X2=0 $Y2=0
cc_504 N_VPWR_c_713_n N_X_c_889_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_505 N_VPWR_M1011_d N_X_c_856_n 0.00176461f $X=6.87 $Y=1.835 $X2=0 $Y2=0
cc_506 N_VPWR_c_718_n N_X_c_856_n 0.0170777f $X=7.01 $Y=2.18 $X2=0 $Y2=0
cc_507 N_VPWR_c_724_n N_X_c_893_n 0.0124525f $X=7.705 $Y=3.33 $X2=0 $Y2=0
cc_508 N_VPWR_c_713_n N_X_c_893_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_509 N_VPWR_M1027_d N_X_c_858_n 0.00270455f $X=7.73 $Y=1.835 $X2=0 $Y2=0
cc_510 N_VPWR_c_720_n N_X_c_858_n 0.023955f $X=7.87 $Y=2.18 $X2=0 $Y2=0
cc_511 N_X_c_850_n N_VGND_M1007_s 0.00176461f $X=7.345 $Y=1.14 $X2=0 $Y2=0
cc_512 N_X_c_852_n N_VGND_M1020_s 2.33864e-19 $X=7.81 $Y=1.14 $X2=0 $Y2=0
cc_513 N_X_c_854_n N_VGND_M1020_s 0.0021884f $X=7.942 $Y=1.225 $X2=0 $Y2=0
cc_514 N_X_c_850_n N_VGND_c_999_n 0.0170777f $X=7.345 $Y=1.14 $X2=0 $Y2=0
cc_515 N_X_c_852_n N_VGND_c_1001_n 0.00362085f $X=7.81 $Y=1.14 $X2=0 $Y2=0
cc_516 N_X_c_854_n N_VGND_c_1001_n 0.0203341f $X=7.942 $Y=1.225 $X2=0 $Y2=0
cc_517 N_X_c_903_p N_VGND_c_1008_n 0.0120977f $X=6.58 $Y=0.42 $X2=0 $Y2=0
cc_518 N_X_c_904_p N_VGND_c_1009_n 0.0120977f $X=7.44 $Y=0.42 $X2=0 $Y2=0
cc_519 N_X_M1000_d N_VGND_c_1013_n 0.00571434f $X=6.44 $Y=0.245 $X2=0 $Y2=0
cc_520 N_X_M1009_d N_VGND_c_1013_n 0.00571434f $X=7.3 $Y=0.245 $X2=0 $Y2=0
cc_521 N_X_c_903_p N_VGND_c_1013_n 0.00691495f $X=6.58 $Y=0.42 $X2=0 $Y2=0
cc_522 N_X_c_904_p N_VGND_c_1013_n 0.00691495f $X=7.44 $Y=0.42 $X2=0 $Y2=0
cc_523 N_A_44_65#_c_910_n N_VGND_M1012_d 0.00721225f $X=1.16 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_524 N_A_44_65#_c_913_n N_VGND_M1012_d 0.00394282f $X=1.64 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_525 N_A_44_65#_c_925_n N_VGND_M1019_d 0.00476476f $X=2.31 $Y=0.955 $X2=0
+ $Y2=0
cc_526 N_A_44_65#_c_942_n N_VGND_M1017_d 0.00370902f $X=3.23 $Y=0.955 $X2=0
+ $Y2=0
cc_527 N_A_44_65#_c_912_n N_VGND_c_996_n 0.0194243f $X=1.545 $Y=0.45 $X2=0 $Y2=0
cc_528 N_A_44_65#_c_925_n N_VGND_c_996_n 0.0170777f $X=2.31 $Y=0.955 $X2=0 $Y2=0
cc_529 N_A_44_65#_c_914_n N_VGND_c_996_n 0.0155793f $X=2.435 $Y=0.47 $X2=0 $Y2=0
cc_530 N_A_44_65#_c_914_n N_VGND_c_997_n 0.0155793f $X=2.435 $Y=0.47 $X2=0 $Y2=0
cc_531 N_A_44_65#_c_942_n N_VGND_c_997_n 0.0171813f $X=3.23 $Y=0.955 $X2=0 $Y2=0
cc_532 N_A_44_65#_c_916_n N_VGND_c_997_n 0.00962585f $X=3.855 $Y=0.34 $X2=0
+ $Y2=0
cc_533 N_A_44_65#_c_917_n N_VGND_c_998_n 0.0147177f $X=5.465 $Y=0.345 $X2=0
+ $Y2=0
cc_534 N_A_44_65#_c_918_n N_VGND_c_998_n 0.0353829f $X=5.63 $Y=0.47 $X2=0 $Y2=0
cc_535 N_A_44_65#_c_912_n N_VGND_c_1002_n 0.016703f $X=1.545 $Y=0.45 $X2=0 $Y2=0
cc_536 N_A_44_65#_c_914_n N_VGND_c_1004_n 0.0134916f $X=2.435 $Y=0.47 $X2=0
+ $Y2=0
cc_537 N_A_44_65#_c_909_n N_VGND_c_1006_n 0.0140356f $X=0.345 $Y=0.47 $X2=0
+ $Y2=0
cc_538 N_A_44_65#_c_915_n N_VGND_c_1007_n 0.0423306f $X=4.525 $Y=0.34 $X2=0
+ $Y2=0
cc_539 N_A_44_65#_c_916_n N_VGND_c_1007_n 0.0448042f $X=3.855 $Y=0.34 $X2=0
+ $Y2=0
cc_540 N_A_44_65#_c_917_n N_VGND_c_1007_n 0.0666169f $X=5.465 $Y=0.345 $X2=0
+ $Y2=0
cc_541 N_A_44_65#_c_919_n N_VGND_c_1007_n 0.0178385f $X=4.655 $Y=0.34 $X2=0
+ $Y2=0
cc_542 N_A_44_65#_c_909_n N_VGND_c_1010_n 0.0253056f $X=0.345 $Y=0.47 $X2=0
+ $Y2=0
cc_543 N_A_44_65#_c_910_n N_VGND_c_1010_n 0.0318053f $X=1.16 $Y=1.17 $X2=0 $Y2=0
cc_544 N_A_44_65#_c_912_n N_VGND_c_1010_n 0.0273527f $X=1.545 $Y=0.45 $X2=0
+ $Y2=0
cc_545 N_A_44_65#_c_913_n N_VGND_c_1010_n 0.00646361f $X=1.64 $Y=0.955 $X2=0
+ $Y2=0
cc_546 N_A_44_65#_c_909_n N_VGND_c_1013_n 0.00977851f $X=0.345 $Y=0.47 $X2=0
+ $Y2=0
cc_547 N_A_44_65#_c_912_n N_VGND_c_1013_n 0.0090585f $X=1.545 $Y=0.45 $X2=0
+ $Y2=0
cc_548 N_A_44_65#_c_914_n N_VGND_c_1013_n 0.0093995f $X=2.435 $Y=0.47 $X2=0
+ $Y2=0
cc_549 N_A_44_65#_c_915_n N_VGND_c_1013_n 0.0239351f $X=4.525 $Y=0.34 $X2=0
+ $Y2=0
cc_550 N_A_44_65#_c_916_n N_VGND_c_1013_n 0.0242986f $X=3.855 $Y=0.34 $X2=0
+ $Y2=0
cc_551 N_A_44_65#_c_917_n N_VGND_c_1013_n 0.0370371f $X=5.465 $Y=0.345 $X2=0
+ $Y2=0
cc_552 N_A_44_65#_c_919_n N_VGND_c_1013_n 0.00981287f $X=4.655 $Y=0.34 $X2=0
+ $Y2=0
