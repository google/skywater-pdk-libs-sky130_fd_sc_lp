* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VGND a_80_237# X VNB nshort w=840000u l=150000u
+  ad=7.602e+11p pd=5.17e+06u as=2.226e+11p ps=2.21e+06u
M1001 a_300_367# B1 a_80_237# VPB phighvt w=1.26e+06u l=150000u
+  ad=6.867e+11p pd=6.13e+06u as=3.339e+11p ps=3.05e+06u
M1002 a_378_47# A1 a_80_237# VNB nshort w=840000u l=150000u
+  ad=3.528e+11p pd=2.52e+06u as=3.318e+11p ps=2.47e+06u
M1003 a_80_237# B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_300_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=8.127e+11p ps=6.33e+06u
M1005 VGND A2 a_378_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_300_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_80_237# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends
