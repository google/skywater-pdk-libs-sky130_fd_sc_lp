# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__einvn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__einvn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.355000 1.185000 6.135000 1.515000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.827000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.210000 0.775000 1.645000 ;
        RECT 0.105000 1.645000 0.415000 2.960000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.355000 0.690000 6.475000 1.015000 ;
        RECT 5.355000 1.685000 8.265000 1.875000 ;
        RECT 5.355000 1.875000 5.685000 2.735000 ;
        RECT 6.215000 1.875000 6.545000 2.735000 ;
        RECT 6.305000 1.015000 6.475000 1.140000 ;
        RECT 6.305000 1.140000 8.225000 1.665000 ;
        RECT 6.305000 1.665000 8.265000 1.685000 ;
        RECT 7.075000 1.875000 7.405000 2.735000 ;
        RECT 7.145000 0.595000 7.335000 1.140000 ;
        RECT 7.935000 1.875000 8.265000 2.735000 ;
        RECT 8.005000 0.595000 8.225000 1.140000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 9.120000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 9.310000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.095000  0.085000 0.390000 1.040000 ;
      RECT 0.585000  0.265000 0.795000 0.665000 ;
      RECT 0.585000  0.665000 1.315000 1.040000 ;
      RECT 0.595000  1.815000 0.805000 3.245000 ;
      RECT 0.985000  1.040000 1.315000 3.075000 ;
      RECT 1.485000  0.255000 1.780000 1.285000 ;
      RECT 1.485000  1.285000 5.185000 1.505000 ;
      RECT 1.485000  1.675000 5.185000 1.925000 ;
      RECT 1.485000  1.925000 1.745000 3.075000 ;
      RECT 1.915000  2.095000 2.245000 3.245000 ;
      RECT 1.950000  0.085000 2.210000 1.115000 ;
      RECT 2.380000  0.255000 2.640000 1.285000 ;
      RECT 2.415000  1.925000 2.605000 3.075000 ;
      RECT 2.775000  2.095000 3.105000 3.245000 ;
      RECT 2.810000  0.085000 3.070000 1.115000 ;
      RECT 3.240000  0.255000 3.500000 1.285000 ;
      RECT 3.275000  1.925000 3.465000 3.075000 ;
      RECT 3.635000  2.095000 3.965000 3.245000 ;
      RECT 3.670000  0.085000 3.930000 1.115000 ;
      RECT 4.100000  0.255000 4.360000 1.285000 ;
      RECT 4.135000  1.925000 4.325000 3.075000 ;
      RECT 4.495000  2.095000 4.825000 3.245000 ;
      RECT 4.530000  0.085000 4.790000 1.115000 ;
      RECT 4.960000  0.255000 8.695000 0.425000 ;
      RECT 4.960000  0.425000 6.975000 0.520000 ;
      RECT 4.960000  0.520000 5.185000 1.285000 ;
      RECT 4.995000  1.925000 5.185000 2.905000 ;
      RECT 4.995000  2.905000 8.695000 3.075000 ;
      RECT 5.855000  2.055000 6.045000 2.905000 ;
      RECT 6.645000  0.520000 6.975000 0.970000 ;
      RECT 6.715000  2.055000 6.905000 2.905000 ;
      RECT 7.505000  0.425000 7.835000 0.970000 ;
      RECT 7.575000  2.055000 7.765000 2.905000 ;
      RECT 8.395000  0.425000 8.695000 1.095000 ;
      RECT 8.435000  1.825000 8.695000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_lp__einvn_8
END LIBRARY
