# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__isobufsrc_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__isobufsrc_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.345000 0.435000 1.760000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.965000 1.425000 1.295000 1.695000 ;
        RECT 0.965000 1.695000 4.305000 1.865000 ;
        RECT 2.065000 1.425000 3.205000 1.695000 ;
        RECT 4.045000 1.345000 4.305000 1.695000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  1.646400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.200000 0.255000 1.530000 0.745000 ;
        RECT 1.200000 0.745000 4.030000 0.915000 ;
        RECT 1.630000 2.035000 4.700000 2.205000 ;
        RECT 1.630000 2.205000 1.960000 2.255000 ;
        RECT 2.060000 0.255000 2.390000 0.745000 ;
        RECT 2.920000 0.255000 3.250000 0.745000 ;
        RECT 3.410000 2.205000 3.620000 2.715000 ;
        RECT 3.840000 0.915000 4.030000 1.005000 ;
        RECT 3.840000 1.005000 4.700000 1.175000 ;
        RECT 3.850000 0.255000 4.030000 0.745000 ;
        RECT 4.475000 1.175000 4.700000 2.035000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.260000  0.255000 0.520000 1.005000 ;
      RECT 0.260000  1.005000 0.785000 1.085000 ;
      RECT 0.260000  1.085000 3.635000 1.175000 ;
      RECT 0.260000  1.930000 0.785000 2.100000 ;
      RECT 0.260000  2.100000 0.530000 3.075000 ;
      RECT 0.615000  1.175000 3.635000 1.255000 ;
      RECT 0.615000  1.255000 0.785000 1.930000 ;
      RECT 0.690000  0.085000 1.020000 0.835000 ;
      RECT 0.750000  2.270000 1.080000 2.425000 ;
      RECT 0.750000  2.425000 2.820000 2.655000 ;
      RECT 0.750000  2.655000 1.030000 3.245000 ;
      RECT 1.200000  2.825000 3.190000 2.885000 ;
      RECT 1.200000  2.885000 4.040000 3.065000 ;
      RECT 1.565000  1.255000 1.895000 1.515000 ;
      RECT 1.700000  0.085000 1.890000 0.575000 ;
      RECT 2.560000  0.085000 2.750000 0.575000 ;
      RECT 2.990000  2.375000 3.190000 2.825000 ;
      RECT 3.375000  1.255000 3.635000 1.515000 ;
      RECT 3.420000  0.085000 3.680000 0.575000 ;
      RECT 3.840000  2.375000 4.040000 2.885000 ;
      RECT 4.210000  0.085000 4.540000 0.835000 ;
      RECT 4.210000  2.375000 4.540000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__isobufsrc_4
END LIBRARY
