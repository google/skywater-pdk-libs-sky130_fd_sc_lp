* File: sky130_fd_sc_lp__a22oi_lp.spice
* Created: Fri Aug 28 09:55:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22oi_lp.pex.spice"
.subckt sky130_fd_sc_lp__a22oi_lp  VNB VPB B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1005 A_171_47# N_B2_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g A_171_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0504 PD=0.81 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1000 A_357_47# N_A1_M1000_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0819 PD=0.84 PS=0.81 NRD=44.28 NRS=31.428 M=1 R=2.8 SA=75001.1 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g A_357_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0882 PD=1.41 PS=0.84 NRD=0 NRS=44.28 M=1 R=2.8 SA=75001.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_B2_M1004_g N_A_64_409#_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1002 N_A_64_409#_M1002_d N_B1_M1002_g N_Y_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_64_409#_M1002_d VPB PHIGHVT L=0.25 W=1
+ AD=0.145 AS=0.14 PD=1.29 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_A_64_409#_M1001_d N_A2_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.145 PD=2.57 PS=1.29 NRD=0 NRS=1.9503 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__a22oi_lp.pxi.spice"
*
.ends
*
*
