* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o211a_m A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_217_49# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND A2 a_217_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR C1 a_80_60# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_217_49# B1 a_488_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 X a_80_60# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_80_60# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR A1 a_300_371# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 X a_80_60# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_300_371# A2 a_80_60# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_488_49# C1 a_80_60# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
