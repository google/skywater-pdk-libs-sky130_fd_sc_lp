* File: sky130_fd_sc_lp__inputiso0n_lp.pex.spice
* Created: Wed Sep  2 09:54:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INPUTISO0N_LP%A 3 7 11 13 19 20
c35 19 0 1.16381e-19 $X=0.87 $Y=1.48
r36 18 20 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.87 $Y=1.48
+ $X2=1.03 $Y2=1.48
r37 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.87
+ $Y=1.48 $X2=0.87 $Y2=1.48
r38 15 18 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.67 $Y=1.48 $X2=0.87
+ $Y2=1.48
r39 13 19 2.97013 $w=7.43e-07 $l=1.85e-07 $layer=LI1_cond $X=0.717 $Y=1.665
+ $X2=0.717 $Y2=1.48
r40 9 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.645
+ $X2=1.03 $Y2=1.48
r41 9 11 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.03 $Y=1.645
+ $X2=1.03 $Y2=2.655
r42 5 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.315
+ $X2=1.03 $Y2=1.48
r43 5 7 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.03 $Y=1.315 $X2=1.03
+ $Y2=0.675
r44 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=1.645
+ $X2=0.67 $Y2=1.48
r45 1 3 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.67 $Y=1.645
+ $X2=0.67 $Y2=2.655
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0N_LP%SLEEP_B 3 7 11 13 19 20
c41 20 0 1.48936e-19 $X=1.82 $Y=1.48
c42 7 0 1.16381e-19 $X=1.46 $Y=2.655
r43 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.82
+ $Y=1.48 $X2=1.82 $Y2=1.48
r44 17 19 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.46 $Y=1.48
+ $X2=1.82 $Y2=1.48
r45 15 17 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.39 $Y=1.48 $X2=1.46
+ $Y2=1.48
r46 13 20 3.3026 $w=6.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.48
r47 9 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=1.645
+ $X2=1.82 $Y2=1.48
r48 9 11 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.82 $Y=1.645
+ $X2=1.82 $Y2=2.655
r49 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.46 $Y=1.645
+ $X2=1.46 $Y2=1.48
r50 5 7 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.46 $Y=1.645
+ $X2=1.46 $Y2=2.655
r51 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.315
+ $X2=1.39 $Y2=1.48
r52 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.39 $Y=1.315 $X2=1.39
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0N_LP%A_138_93# 1 2 7 9 12 14 16 19 23 25 26
+ 29 31 32 33 34 37
c69 37 0 9.55314e-20 $X=2.515 $Y=1.17
r70 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.515
+ $Y=1.17 $X2=2.515 $Y2=1.17
r71 33 36 2.47908 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=1.225
+ $X2=2.48 $Y2=1.14
r72 33 34 20.5191 $w=4.08e-07 $l=7.3e-07 $layer=LI1_cond $X=2.48 $Y=1.225
+ $X2=2.48 $Y2=1.955
r73 31 34 8.45803 $w=1.7e-07 $l=2.43824e-07 $layer=LI1_cond $X=2.275 $Y=2.04
+ $X2=2.48 $Y2=1.955
r74 31 32 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.275 $Y=2.04
+ $X2=1.41 $Y2=2.04
r75 27 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.245 $Y=2.125
+ $X2=1.41 $Y2=2.04
r76 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=1.245 $Y=2.125
+ $X2=1.245 $Y2=2.655
r77 25 36 5.97895 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.275 $Y=1.14
+ $X2=2.48 $Y2=1.14
r78 25 26 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=2.275 $Y=1.14
+ $X2=0.98 $Y2=1.14
r79 21 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.815 $Y=1.055
+ $X2=0.98 $Y2=1.14
r80 21 23 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.815 $Y=1.055
+ $X2=0.815 $Y2=0.675
r81 17 37 97.1997 $w=2.55e-07 $l=5.88154e-07 $layer=POLY_cond $X=2.75 $Y=1.675
+ $X2=2.57 $Y2=1.17
r82 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.75 $Y=1.675
+ $X2=2.75 $Y2=2.465
r83 14 37 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=2.75 $Y=1.005
+ $X2=2.57 $Y2=1.17
r84 14 16 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.75 $Y=1.005
+ $X2=2.75 $Y2=0.675
r85 10 37 97.1997 $w=2.55e-07 $l=5.88154e-07 $layer=POLY_cond $X=2.39 $Y=1.675
+ $X2=2.57 $Y2=1.17
r86 10 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.39 $Y=1.675
+ $X2=2.39 $Y2=2.465
r87 7 37 32.933 $w=2.55e-07 $l=1.8e-07 $layer=POLY_cond $X=2.39 $Y=1.17 $X2=2.57
+ $Y2=1.17
r88 7 9 106.04 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.39 $Y=1.17 $X2=2.39
+ $Y2=0.675
r89 2 29 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=2.445 $X2=1.245 $Y2=2.655
r90 1 23 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.465 $X2=0.815 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0N_LP%VPWR 1 2 9 13 16 17 18 23 32 33 36
c34 13 0 9.55314e-20 $X=2.175 $Y=2.38
r35 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 33 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 30 36 13.5049 $w=1.7e-07 $l=3.43e-07 $layer=LI1_cond $X=2.675 $Y=3.33
+ $X2=2.332 $Y2=3.33
r39 30 32 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.675 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r41 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 23 36 13.5049 $w=1.7e-07 $l=3.42e-07 $layer=LI1_cond $X=1.99 $Y=3.33
+ $X2=2.332 $Y2=3.33
r43 23 28 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.99 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 22 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 18 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 18 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 18 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 16 21 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=0.29 $Y=3.33 $X2=0.24
+ $Y2=3.33
r50 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.29 $Y=3.33
+ $X2=0.455 $Y2=3.33
r51 15 25 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.62 $Y=3.33 $X2=0.72
+ $Y2=3.33
r52 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.455 $Y2=3.33
r53 11 36 2.81621 $w=6.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.332 $Y=3.245
+ $X2=2.332 $Y2=3.33
r54 11 13 15.1038 $w=6.83e-07 $l=8.65e-07 $layer=LI1_cond $X=2.332 $Y=3.245
+ $X2=2.332 $Y2=2.38
r55 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.455 $Y=3.245
+ $X2=0.455 $Y2=3.33
r56 7 9 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.455 $Y=3.245
+ $X2=0.455 $Y2=2.655
r57 2 13 300 $w=1.7e-07 $l=3.10805e-07 $layer=licon1_PDIFF $count=2 $X=1.895
+ $Y=2.445 $X2=2.175 $Y2=2.38
r58 1 9 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.33
+ $Y=2.445 $X2=0.455 $Y2=2.655
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0N_LP%X 1 2 7 8 9 10 11 18 21 24 27 30 35
r10 33 35 7.54576 $w=4.18e-07 $l=2.75e-07 $layer=LI1_cond $X=3.065 $Y=2.125
+ $X2=3.065 $Y2=2.4
r11 18 21 5.48782 $w=4.18e-07 $l=2e-07 $layer=LI1_cond $X=3.065 $Y=0.72
+ $X2=3.065 $Y2=0.92
r12 11 38 13.5824 $w=4.18e-07 $l=4.95e-07 $layer=LI1_cond $X=3.065 $Y=2.405
+ $X2=3.065 $Y2=2.9
r13 11 35 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=2.405
+ $X2=3.065 $Y2=2.4
r14 10 33 2.46952 $w=4.18e-07 $l=9e-08 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=3.065 $Y2=2.125
r15 10 30 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=2.035
+ $X2=3.065 $Y2=2.03
r16 9 30 10.0153 $w=4.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.065 $Y=1.665
+ $X2=3.065 $Y2=2.03
r17 9 27 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=1.665
+ $X2=3.065 $Y2=1.66
r18 8 27 10.0153 $w=4.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.065 $Y=1.295
+ $X2=3.065 $Y2=1.66
r19 8 24 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=1.295
+ $X2=3.065 $Y2=1.29
r20 7 24 10.0153 $w=4.18e-07 $l=3.65e-07 $layer=LI1_cond $X=3.065 $Y=0.925
+ $X2=3.065 $Y2=1.29
r21 7 21 0.137196 $w=4.18e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=0.925
+ $X2=3.065 $Y2=0.92
r22 2 38 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.835 $X2=2.965 $Y2=2.9
r23 2 33 400 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=1.835 $X2=2.965 $Y2=2.125
r24 1 18 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=2.825
+ $Y=0.465 $X2=2.965 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__INPUTISO0N_LP%VGND 1 4 16 17 22 28
r23 27 28 12.4206 $w=9.23e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=0.377
+ $X2=2.335 $Y2=0.377
r24 24 27 0.131892 $w=9.23e-07 $l=1e-08 $layer=LI1_cond $X=2.16 $Y=0.377
+ $X2=2.17 $Y2=0.377
r25 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r26 20 24 6.33081 $w=9.23e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.377
+ $X2=2.16 $Y2=0.377
r27 20 22 13.4097 $w=9.23e-07 $l=2.4e-07 $layer=LI1_cond $X=1.68 $Y=0.377
+ $X2=1.44 $Y2=0.377
r28 17 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r29 16 28 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=2.335
+ $Y2=0
r30 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r31 12 22 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.44
+ $Y2=0
r32 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 9 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r34 8 12 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r35 8 9 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r36 4 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r37 4 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r38 4 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r39 1 27 91 $w=1.7e-07 $l=8.03166e-07 $layer=licon1_NDIFF $count=2 $X=1.465
+ $Y=0.465 $X2=2.17 $Y2=0.675
.ends

