* NGSPICE file created from sky130_fd_sc_lp__invkapwr_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__invkapwr_1 A KAPWR VGND VNB VPB VPWR Y
M1000 KAPWR A Y VPB phighvt w=840000u l=150000u
+  ad=4.452e+11p pd=4.42e+06u as=2.352e+11p ps=2.24e+06u
M1001 VGND A Y VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.113e+11p ps=1.37e+06u
M1002 Y A KAPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

