* NGSPICE file created from sky130_fd_sc_lp__nand3b_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand3b_lp A_N B C VGND VNB VPB VPWR Y
M1000 a_156_141# a_90_247# Y VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1001 VPWR C Y VPB phighvt w=1e+06u l=250000u
+  ad=6e+11p pd=5.2e+06u as=5.65e+11p ps=5.13e+06u
M1002 VGND C a_234_141# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.008e+11p ps=1.32e+06u
M1003 Y B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_90_247# A_N a_420_141# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1005 a_234_141# B a_156_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_420_141# A_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_90_247# Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_90_247# A_N VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends

