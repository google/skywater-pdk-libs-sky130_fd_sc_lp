* File: sky130_fd_sc_lp__xor3_1.spice
* Created: Fri Aug 28 11:37:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xor3_1.pex.spice"
.subckt sky130_fd_sc_lp__xor3_1  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_86_305#_M1007_g N_A_42_411#_M1007_s VNB NSHORT L=0.15
+ W=0.64 AD=0.23675 AS=0.1824 PD=1.615 PS=1.85 NRD=59.04 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75003 A=0.096 P=1.58 MULT=1
MM1004 N_A_86_305#_M1004_d N_A_M1004_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.64
+ AD=0.176 AS=0.23675 PD=1.19 PS=1.615 NRD=0 NRS=59.04 M=1 R=4.26667 SA=75000.9
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1018 N_A_425_117#_M1018_d N_B_M1018_g N_A_86_305#_M1004_d VNB NSHORT L=0.15
+ W=0.64 AD=0.138023 AS=0.176 PD=1.24981 PS=1.19 NRD=0 NRS=50.616 M=1 R=4.26667
+ SA=75001.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_42_411#_M1020_d N_A_474_313#_M1020_g N_A_425_117#_M1018_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.129883 AS=0.0905774 PD=0.943019 PS=0.820189 NRD=32.856
+ NRS=33.564 M=1 R=2.8 SA=75002.1 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_402_411#_M1010_d N_B_M1010_g N_A_42_411#_M1020_d VNB NSHORT L=0.15
+ W=0.64 AD=0.169 AS=0.197917 PD=1.19 PS=1.43698 NRD=21.552 NRS=29.052 M=1
+ R=4.26667 SA=75002 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1021 N_A_86_305#_M1021_d N_A_474_313#_M1021_g N_A_402_411#_M1010_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.3328 AS=0.169 PD=2.32 PS=1.19 NRD=44.052 NRS=21.552 M=1
+ R=4.26667 SA=75002.6 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_B_M1005_g N_A_474_313#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.4662 AS=0.2394 PD=2.79 PS=2.25 NRD=38.568 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.5 A=0.126 P=1.98 MULT=1
MM1001 N_A_1363_127#_M1001_d N_A_1263_295#_M1001_g N_A_402_411#_M1001_s VNB
+ NSHORT L=0.15 W=0.64 AD=0.0896 AS=0.3552 PD=0.92 PS=2.39 NRD=0 NRS=50.616 M=1
+ R=4.26667 SA=75000.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1014 N_A_425_117#_M1014_d N_C_M1014_g N_A_1363_127#_M1001_d VNB NSHORT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_C_M1015_g N_A_1263_295#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.1197 PD=0.876667 PS=1.41 NRD=32.856 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1012 N_X_M1012_d N_A_1363_127#_M1012_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.2352 PD=2.25 PS=1.75333 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A_86_305#_M1000_g N_A_42_411#_M1000_s VPB PHIGHVT L=0.15
+ W=1 AD=0.335 AS=0.285 PD=1.67 PS=2.57 NRD=0 NRS=0 M=1 R=6.66667 SA=75000.2
+ SB=75002.7 A=0.15 P=2.3 MULT=1
MM1016 N_A_86_305#_M1016_d N_A_M1016_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1
+ AD=0.205109 AS=0.335 PD=1.5163 PS=1.67 NRD=0 NRS=76.8103 M=1 R=6.66667
+ SA=75001 SB=75001.9 A=0.15 P=2.3 MULT=1
MM1002 N_A_402_411#_M1002_d N_B_M1002_g N_A_86_305#_M1016_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.159146 AS=0.172291 PD=1.36216 PS=1.2737 NRD=0 NRS=27.3436 M=1
+ R=5.6 SA=75001.6 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1003 N_A_42_411#_M1003_d N_A_474_313#_M1003_g N_A_402_411#_M1002_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.121254 PD=0.92 PS=1.03784 NRD=0 NRS=24.6053 M=1
+ R=4.26667 SA=75002.1 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1013 N_A_425_117#_M1013_d N_B_M1013_g N_A_42_411#_M1003_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.133514 AS=0.0896 PD=1.06811 PS=0.92 NRD=36.9375 NRS=0 M=1
+ R=4.26667 SA=75002.5 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1019 N_A_86_305#_M1019_d N_A_474_313#_M1019_g N_A_425_117#_M1013_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.5922 AS=0.175236 PD=3.09 PS=1.40189 NRD=98.5 NRS=0 M=1
+ R=5.6 SA=75002.4 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_A_474_313#_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.3591 PD=3.09 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1017 N_A_1363_127#_M1017_d N_A_1263_295#_M1017_g N_A_425_117#_M1017_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1176 AS=0.6678 PD=1.12 PS=3.27 NRD=0 NRS=119.599
+ M=1 R=5.6 SA=75000.7 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1011 N_A_402_411#_M1011_d N_C_M1011_g N_A_1363_127#_M1017_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_C_M1008_g N_A_1263_295#_M1008_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.280488 AS=0.1824 PD=1.33053 PS=1.85 NRD=36.1495 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_X_M1009_d N_A_1363_127#_M1009_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.552212 PD=3.09 PS=2.61947 NRD=0 NRS=50.0183 M=1 R=8.4
+ SA=75000.8 SB=75000.2 A=0.189 P=2.82 MULT=1
DX22_noxref VNB VPB NWDIODE A=18.6667 P=23.79
c_97 VNB 0 1.8437e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__xor3_1.pxi.spice"
*
.ends
*
*
