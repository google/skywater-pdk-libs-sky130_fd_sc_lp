* File: sky130_fd_sc_lp__xor2_m.pex.spice
* Created: Fri Aug 28 11:36:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XOR2_M%A 1 3 7 11 13 17 23 24 26 33
c50 26 0 3.95594e-20 $X=1.2 $Y=2.405
c51 1 0 2.13341e-19 $X=0.905 $Y=2.5
r52 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.065
+ $Y=1.995 $X2=1.065 $Y2=1.995
r53 26 34 2.78398 $w=5.78e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=2.2
+ $X2=1.065 $Y2=2.2
r54 24 34 7.1146 $w=5.78e-07 $l=3.45e-07 $layer=LI1_cond $X=0.72 $Y=2.2
+ $X2=1.065 $Y2=2.2
r55 22 33 14.6871 $w=5.1e-07 $l=1.4e-07 $layer=POLY_cond $X=1.155 $Y=1.855
+ $X2=1.155 $Y2=1.995
r56 22 23 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.155 $Y=1.855
+ $X2=1.155 $Y2=1.78
r57 20 33 37.2422 $w=5.1e-07 $l=3.55e-07 $layer=POLY_cond $X=1.155 $Y=2.35
+ $X2=1.155 $Y2=1.995
r58 15 17 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=1.71 $Y=1.705
+ $X2=1.71 $Y2=0.99
r59 14 23 16.9349 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.41 $Y=1.78
+ $X2=1.155 $Y2=1.78
r60 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.635 $Y=1.78
+ $X2=1.71 $Y2=1.705
r61 13 14 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.635 $Y=1.78
+ $X2=1.41 $Y2=1.78
r62 5 23 10.1687 $w=3.3e-07 $l=2.14243e-07 $layer=POLY_cond $X=0.975 $Y=1.705
+ $X2=1.155 $Y2=1.78
r63 5 7 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=0.975 $Y=1.705
+ $X2=0.975 $Y2=0.99
r64 1 20 24.7327 $w=5.1e-07 $l=1.5e-07 $layer=POLY_cond $X=1.12 $Y=2.5 $X2=1.12
+ $Y2=2.35
r65 1 11 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.335 $Y=2.5
+ $X2=1.335 $Y2=2.885
r66 1 3 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.905 $Y=2.5
+ $X2=0.905 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_M%B 3 5 7 8 11 13 14 18 19 20 21 31 35
c65 11 0 3.95594e-20 $X=1.765 $Y=2.885
r66 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=0.43
+ $X2=2.16 $Y2=0.595
r67 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=0.43 $X2=2.16 $Y2=0.43
r68 31 34 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.16 $Y=0.335
+ $X2=2.16 $Y2=0.43
r69 20 21 6.80845 $w=6.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=0.925
+ $X2=1.92 $Y2=1.295
r70 19 20 6.80845 $w=6.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=0.555
+ $X2=1.92 $Y2=0.925
r71 19 35 2.30015 $w=6.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.92 $Y=0.555
+ $X2=1.92 $Y2=0.43
r72 18 36 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.07 $Y=0.99
+ $X2=2.07 $Y2=0.595
r73 16 18 566.606 $w=1.5e-07 $l=1.105e-06 $layer=POLY_cond $X=2.07 $Y=2.095
+ $X2=2.07 $Y2=0.99
r74 13 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.995 $Y=2.17
+ $X2=2.07 $Y2=2.095
r75 13 14 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.995 $Y=2.17
+ $X2=1.84 $Y2=2.17
r76 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.765 $Y=2.245
+ $X2=1.84 $Y2=2.17
r77 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.765 $Y=2.245
+ $X2=1.765 $Y2=2.885
r78 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.995 $Y=0.335
+ $X2=2.16 $Y2=0.335
r79 7 8 705.053 $w=1.5e-07 $l=1.375e-06 $layer=POLY_cond $X=1.995 $Y=0.335
+ $X2=0.62 $Y2=0.335
r80 3 5 971.691 $w=1.5e-07 $l=1.895e-06 $layer=POLY_cond $X=0.545 $Y=0.99
+ $X2=0.545 $Y2=2.885
r81 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.545 $Y=0.41
+ $X2=0.62 $Y2=0.335
r82 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.545 $Y=0.41
+ $X2=0.545 $Y2=0.99
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_M%A_41_535# 1 2 9 13 17 18 21 23 24 27 29 33 35
+ 36
c65 33 0 1.14239e-19 $X=0.76 $Y=1.645
c66 29 0 9.91016e-20 $X=2.685 $Y=1.645
r67 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.77
+ $Y=1.725 $X2=2.77 $Y2=1.725
r68 30 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.865 $Y=1.645
+ $X2=0.76 $Y2=1.645
r69 29 35 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=1.645
+ $X2=2.77 $Y2=1.645
r70 29 30 118.738 $w=1.68e-07 $l=1.82e-06 $layer=LI1_cond $X=2.685 $Y=1.645
+ $X2=0.865 $Y2=1.645
r71 25 33 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=1.56
+ $X2=0.76 $Y2=1.645
r72 25 27 26.671 $w=2.08e-07 $l=5.05e-07 $layer=LI1_cond $X=0.76 $Y=1.56
+ $X2=0.76 $Y2=1.055
r73 23 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.655 $Y=1.645
+ $X2=0.76 $Y2=1.645
r74 23 24 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.655 $Y=1.645
+ $X2=0.435 $Y2=1.645
r75 19 24 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.33 $Y=1.73
+ $X2=0.435 $Y2=1.645
r76 19 21 58.3593 $w=2.08e-07 $l=1.105e-06 $layer=LI1_cond $X=0.33 $Y=1.73
+ $X2=0.33 $Y2=2.835
r77 17 36 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.77 $Y=2.065
+ $X2=2.77 $Y2=1.725
r78 17 18 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=2.065
+ $X2=2.77 $Y2=2.23
r79 16 36 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.56
+ $X2=2.77 $Y2=1.725
r80 13 16 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.725 $Y=0.99
+ $X2=2.725 $Y2=1.56
r81 9 18 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.715 $Y=2.665
+ $X2=2.715 $Y2=2.23
r82 2 21 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=2.675 $X2=0.33 $Y2=2.835
r83 1 27 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.78 $X2=0.76 $Y2=1.055
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_M%VPWR 1 2 9 13 16 17 18 20 33 34 37
r43 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 30 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r47 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.12 $Y2=3.33
r49 25 27 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.12 $Y2=3.33
r53 20 22 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 18 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 18 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 16 27 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.98 $Y2=3.33
r59 15 30 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.98 $Y2=3.33
r61 11 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=3.245
+ $X2=1.98 $Y2=3.33
r62 11 13 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.98 $Y=3.245
+ $X2=1.98 $Y2=2.95
r63 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=3.245 $X2=1.12
+ $Y2=3.33
r64 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.12 $Y=3.245
+ $X2=1.12 $Y2=2.95
r65 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.675 $X2=1.98 $Y2=2.95
r66 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.675 $X2=1.12 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_M%A_282_535# 1 2 9 11 12 13
r24 13 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.46 $Y=2.52 $X2=2.46
+ $Y2=2.6
r25 11 13 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.335 $Y=2.52
+ $X2=2.46 $Y2=2.52
r26 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.335 $Y=2.52
+ $X2=1.655 $Y2=2.52
r27 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.56 $Y=2.605
+ $X2=1.655 $Y2=2.52
r28 7 9 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=1.56 $Y=2.605
+ $X2=1.56 $Y2=2.82
r29 2 16 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.375
+ $Y=2.455 $X2=2.5 $Y2=2.6
r30 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.675 $X2=1.55 $Y2=2.82
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_M%X 1 2 9 11 12 13 14 15 16
c28 9 0 1.46329e-19 $X=2.51 $Y=1.055
r29 16 36 9.31762 $w=2.33e-07 $l=1.9e-07 $layer=LI1_cond $X=3.12 $Y=2.742
+ $X2=2.93 $Y2=2.742
r30 15 16 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.12 $Y=2.405
+ $X2=3.12 $Y2=2.625
r31 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=2.035
+ $X2=3.12 $Y2=2.405
r32 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=2.035
r33 12 13 12.5394 $w=3.38e-07 $l=2.85e-07 $layer=LI1_cond $X=3.12 $Y=1.38
+ $X2=3.12 $Y2=1.665
r34 11 12 15.6756 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=2.615 $Y=1.295
+ $X2=3.035 $Y2=1.295
r35 7 11 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.52 $Y=1.21
+ $X2=2.615 $Y2=1.295
r36 7 9 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.52 $Y=1.21 $X2=2.52
+ $Y2=1.055
r37 2 36 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=2.455 $X2=2.93 $Y2=2.73
r38 1 9 182 $w=1.7e-07 $l=4.83322e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.78 $X2=2.51 $Y2=1.055
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_M%VGND 1 2 3 10 12 16 18 20 22 24 29 41 45
r30 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r31 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r32 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 36 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r34 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r36 30 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r37 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r38 29 44 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=3.115
+ $Y2=0
r39 29 35 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.64
+ $Y2=0
r40 28 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r41 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r42 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 25 38 3.50623 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=0 $X2=0.207
+ $Y2=0
r44 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.415 $Y=0 $X2=0.72
+ $Y2=0
r45 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r46 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.72
+ $Y2=0
r47 22 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r48 22 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r49 22 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r50 18 44 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.035 $Y=0.085
+ $X2=3.115 $Y2=0
r51 18 20 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=3.035 $Y=0.085
+ $X2=3.035 $Y2=0.925
r52 14 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r53 14 16 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.925
r54 10 38 3.33766 $w=1.9e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.207 $Y2=0
r55 10 12 49.0335 $w=1.88e-07 $l=8.4e-07 $layer=LI1_cond $X=0.32 $Y=0.085
+ $X2=0.32 $Y2=0.925
r56 3 20 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.8
+ $Y=0.78 $X2=3.035 $Y2=0.925
r57 2 16 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.78 $X2=1.21 $Y2=0.925
r58 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.78 $X2=0.33 $Y2=0.925
.ends

