* File: sky130_fd_sc_lp__o311ai_0.pex.spice
* Created: Wed Sep  2 10:23:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311AI_0%A1 2 3 5 6 8 12 15 18 20 21 22 27
c40 20 0 2.12572e-19 $X=0.72 $Y=0.925
r41 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.62
+ $Y=0.935 $X2=0.62 $Y2=0.935
r42 21 22 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.687 $Y=1.295
+ $X2=0.687 $Y2=1.665
r43 21 28 13.6026 $w=3.03e-07 $l=3.6e-07 $layer=LI1_cond $X=0.687 $Y=1.295
+ $X2=0.687 $Y2=0.935
r44 20 28 0.37785 $w=3.03e-07 $l=1e-08 $layer=LI1_cond $X=0.687 $Y=0.925
+ $X2=0.687 $Y2=0.935
r45 16 18 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.71 $Y=2.145
+ $X2=0.89 $Y2=2.145
r46 14 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.62 $Y=1.275
+ $X2=0.62 $Y2=0.935
r47 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.62 $Y=1.275
+ $X2=0.62 $Y2=1.44
r48 10 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.62 $Y=0.92
+ $X2=0.62 $Y2=0.935
r49 10 12 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.62 $Y=0.845
+ $X2=0.89 $Y2=0.845
r50 6 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.89 $Y=2.22 $X2=0.89
+ $Y2=2.145
r51 6 8 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.89 $Y=2.22 $X2=0.89
+ $Y2=2.65
r52 3 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.89 $Y=0.77 $X2=0.89
+ $Y2=0.845
r53 3 5 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.89 $Y=0.77 $X2=0.89
+ $Y2=0.45
r54 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.71 $Y=2.07 $X2=0.71
+ $Y2=2.145
r55 2 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.71 $Y=2.07 $X2=0.71
+ $Y2=1.44
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_0%A2 5 9 11 12 13 14 15 16 17 21
c47 15 0 2.70619e-19 $X=1.285 $Y=0.92
c48 5 0 9.63597e-20 $X=1.25 $Y=2.65
r49 16 17 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.182 $Y=1.295
+ $X2=1.182 $Y2=1.665
r50 16 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.16
+ $Y=1.325 $X2=1.16 $Y2=1.325
r51 14 15 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.285 $Y=0.77
+ $X2=1.285 $Y2=0.92
r52 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.16 $Y=1.665
+ $X2=1.16 $Y2=1.325
r53 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.665
+ $X2=1.16 $Y2=1.83
r54 11 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.16
+ $X2=1.16 $Y2=1.325
r55 11 15 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.25 $Y=1.16
+ $X2=1.25 $Y2=0.92
r56 9 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.32 $Y=0.45 $X2=1.32
+ $Y2=0.77
r57 5 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.25 $Y=2.65 $X2=1.25
+ $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_0%A3 2 5 9 11 12 13 17
r39 17 19 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.325
+ $X2=1.73 $Y2=1.16
r40 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.7 $Y=1.295 $X2=1.7
+ $Y2=1.665
r41 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.7
+ $Y=1.325 $X2=1.7 $Y2=1.325
r42 9 19 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.81 $Y=0.45 $X2=1.81
+ $Y2=1.16
r43 5 11 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.61 $Y=2.65 $X2=1.61
+ $Y2=1.83
r44 2 11 49.7341 $w=3.9e-07 $l=1.95e-07 $layer=POLY_cond $X=1.73 $Y=1.635
+ $X2=1.73 $Y2=1.83
r45 1 17 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=1.73 $Y=1.355 $X2=1.73
+ $Y2=1.325
r46 1 2 39.929 $w=3.9e-07 $l=2.8e-07 $layer=POLY_cond $X=1.73 $Y=1.355 $X2=1.73
+ $Y2=1.635
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_0%B1 1 3 6 9 12 16 17 18 19 23
r49 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.33
+ $Y=1.325 $X2=2.33 $Y2=1.325
r50 19 24 8.84058 $w=4.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.265 $Y=1.665
+ $X2=2.265 $Y2=1.325
r51 18 24 0.780051 $w=4.58e-07 $l=3e-08 $layer=LI1_cond $X=2.265 $Y=1.295
+ $X2=2.265 $Y2=1.325
r52 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.33 $Y=1.665
+ $X2=2.33 $Y2=1.325
r53 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=1.665
+ $X2=2.33 $Y2=1.83
r54 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=1.16
+ $X2=2.33 $Y2=1.325
r55 10 12 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.1 $Y=2.145
+ $X2=2.24 $Y2=2.145
r56 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.24 $Y=2.07 $X2=2.24
+ $Y2=2.145
r57 9 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.24 $Y=2.07 $X2=2.24
+ $Y2=1.83
r58 6 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.24 $Y=0.45 $X2=2.24
+ $Y2=1.16
r59 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.1 $Y=2.22 $X2=2.1
+ $Y2=2.145
r60 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.1 $Y=2.22 $X2=2.1
+ $Y2=2.65
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_0%C1 1 3 4 6 7 8 9 10 12 15 16 17 18 23
r45 17 18 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=1.295
+ $X2=3.14 $Y2=1.665
r46 16 17 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=0.925
+ $X2=3.14 $Y2=1.295
r47 16 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.005 $X2=3.09 $Y2=1.005
r48 14 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.09 $Y=1.345
+ $X2=3.09 $Y2=1.005
r49 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.345
+ $X2=3.09 $Y2=1.51
r50 13 23 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=3.09 $Y=0.92
+ $X2=3.09 $Y2=1.005
r51 12 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3 $Y=2.07 $X2=3
+ $Y2=1.51
r52 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.925 $Y=2.145
+ $X2=3 $Y2=2.07
r53 9 10 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.925 $Y=2.145
+ $X2=2.705 $Y2=2.145
r54 7 13 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.925 $Y=0.845
+ $X2=3.09 $Y2=0.92
r55 7 8 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.925 $Y=0.845
+ $X2=2.705 $Y2=0.845
r56 4 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.63 $Y=2.22
+ $X2=2.705 $Y2=2.145
r57 4 6 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.63 $Y=2.22 $X2=2.63
+ $Y2=2.65
r58 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.63 $Y=0.77
+ $X2=2.705 $Y2=0.845
r59 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.63 $Y=0.77 $X2=2.63
+ $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_0%VPWR 1 2 9 13 16 17 18 20 33 34 37
r33 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r39 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.84 $Y=3.33
+ $X2=0.675 $Y2=3.33
r41 25 27 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.84 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.51 $Y=3.33
+ $X2=0.675 $Y2=3.33
r45 20 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.51 $Y=3.33 $X2=0.24
+ $Y2=3.33
r46 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 16 30 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.205 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=3.33
+ $X2=2.37 $Y2=3.33
r50 15 33 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=2.37 $Y2=3.33
r52 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=3.245
+ $X2=2.37 $Y2=3.33
r53 11 13 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.37 $Y=3.245
+ $X2=2.37 $Y2=2.485
r54 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=3.245
+ $X2=0.675 $Y2=3.33
r55 7 9 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.675 $Y=3.245
+ $X2=0.675 $Y2=2.485
r56 2 13 300 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=2 $X=2.175
+ $Y=2.33 $X2=2.37 $Y2=2.485
r57 1 9 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.33 $X2=0.675 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_0%Y 1 2 3 12 14 19 21 22 24 25 35 40
r52 35 40 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.665 $Y=2.035
+ $X2=2.64 $Y2=2.035
r53 25 46 6.29515 $w=5.68e-07 $l=3e-07 $layer=LI1_cond $X=2.99 $Y=2.775 $X2=2.99
+ $Y2=2.475
r54 24 46 1.46887 $w=5.68e-07 $l=7e-08 $layer=LI1_cond $X=2.99 $Y=2.405 $X2=2.99
+ $Y2=2.475
r55 22 35 4.24538 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=2.97 $Y=2.035
+ $X2=2.665 $Y2=2.035
r56 22 24 5.25968 $w=7.58e-07 $l=2.85e-07 $layer=LI1_cond $X=2.99 $Y=2.12
+ $X2=2.99 $Y2=2.405
r57 22 40 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.61 $Y=2.035 $X2=2.64
+ $Y2=2.035
r58 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.16 $Y=2.035
+ $X2=2.61 $Y2=2.035
r59 16 22 67.6995 $w=2.28e-07 $l=1.335e-06 $layer=LI1_cond $X=2.75 $Y=0.615
+ $X2=2.75 $Y2=1.95
r60 15 19 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.75 $Y=0.45
+ $X2=2.845 $Y2=0.45
r61 15 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0.45
+ $X2=2.75 $Y2=0.615
r62 14 21 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=2.035
+ $X2=2.16 $Y2=2.035
r63 10 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.87 $Y=2.12
+ $X2=2.035 $Y2=2.035
r64 10 12 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.87 $Y=2.12
+ $X2=1.87 $Y2=2.475
r65 3 46 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.705
+ $Y=2.33 $X2=2.845 $Y2=2.475
r66 2 12 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=1.685
+ $Y=2.33 $X2=1.87 $Y2=2.475
r67 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.705
+ $Y=0.24 $X2=2.845 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_0%VGND 1 2 9 13 15 17 22 29 30 33 36
c42 22 0 1.54406e-19 $X=1.43 $Y=0
r43 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 27 36 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.715 $Y=0 $X2=1.572
+ $Y2=0
r46 27 29 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=1.715 $Y=0
+ $X2=3.12 $Y2=0
r47 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.84 $Y=0 $X2=0.675
+ $Y2=0
r50 23 25 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.84 $Y=0 $X2=1.2
+ $Y2=0
r51 22 36 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.43 $Y=0 $X2=1.572
+ $Y2=0
r52 22 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.43 $Y=0 $X2=1.2
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.675
+ $Y2=0
r56 17 19 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.24
+ $Y2=0
r57 15 30 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r58 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 15 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 11 36 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.572 $Y=0.085
+ $X2=1.572 $Y2=0
r61 11 13 14.7594 $w=2.83e-07 $l=3.65e-07 $layer=LI1_cond $X=1.572 $Y=0.085
+ $X2=1.572 $Y2=0.45
r62 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=0.085
+ $X2=0.675 $Y2=0
r63 7 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.675 $Y=0.085
+ $X2=0.675 $Y2=0.435
r64 2 13 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=1.395
+ $Y=0.24 $X2=1.57 $Y2=0.45
r65 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.55 $Y=0.24
+ $X2=0.675 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_0%A_193_48# 1 2 9 11 12 15
r39 13 15 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=2.037 $Y=0.785
+ $X2=2.037 $Y2=0.45
r40 11 13 7.16299 $w=2.05e-07 $l=1.96489e-07 $layer=LI1_cond $X=1.885 $Y=0.887
+ $X2=2.037 $Y2=0.785
r41 11 12 33.8137 $w=2.03e-07 $l=6.25e-07 $layer=LI1_cond $X=1.885 $Y=0.887
+ $X2=1.26 $Y2=0.887
r42 7 12 6.90357 $w=2.05e-07 $l=1.68449e-07 $layer=LI1_cond $X=1.135 $Y=0.785
+ $X2=1.26 $Y2=0.887
r43 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.135 $Y=0.785
+ $X2=1.135 $Y2=0.45
r44 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.885
+ $Y=0.24 $X2=2.025 $Y2=0.45
r45 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.965
+ $Y=0.24 $X2=1.105 $Y2=0.45
.ends

