* File: sky130_fd_sc_lp__and3b_1.spice
* Created: Wed Sep  2 09:32:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and3b_1.pex.spice"
.subckt sky130_fd_sc_lp__and3b_1  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1003 N_A_110_47#_M1003_d N_A_N_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_304_47# N_A_110_47#_M1007_g N_A_185_367#_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1008 A_376_47# N_B_M1008_g A_304_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_C_M1009_g A_376_47# VNB NSHORT L=0.15 W=0.42 AD=0.1148
+ AS=0.0441 PD=0.93 PS=0.63 NRD=61.428 NRS=14.28 M=1 R=2.8 SA=75000.9 SB=75000.9
+ A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_185_367#_M1005_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2296 PD=2.21 PS=1.86 NRD=0 NRS=4.284 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_A_110_47#_M1006_d N_A_N_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_110_47#_M1004_g N_A_185_367#_M1004_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.07665 AS=0.1113 PD=0.785 PS=1.37 NRD=18.7544 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_185_367#_M1002_d N_B_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06615 AS=0.07665 PD=0.735 PS=0.785 NRD=9.3772 NRS=21.0987 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_C_M1001_g N_A_185_367#_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.06615 PD=0.8175 PS=0.735 NRD=0 NRS=7.0329 M=1 R=2.8
+ SA=75001.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_185_367#_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=4.9447 M=1 R=8.4 SA=75000.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__and3b_1.pxi.spice"
*
.ends
*
*
