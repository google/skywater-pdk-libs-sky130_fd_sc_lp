* File: sky130_fd_sc_lp__a311oi_m.pex.spice
* Created: Wed Sep  2 09:26:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311OI_M%A3 2 3 4 7 9 11 15 18 19 20 21 22 23 24 25
+ 34
r47 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=0.95 $X2=0.61 $Y2=0.95
r48 24 25 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.665 $Y=2.405
+ $X2=0.665 $Y2=2.775
r49 23 24 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.665 $Y=2.035
+ $X2=0.665 $Y2=2.405
r50 22 23 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.665 $Y=1.665
+ $X2=0.665 $Y2=2.035
r51 21 22 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.665 $Y=1.295
+ $X2=0.665 $Y2=1.665
r52 21 35 14.1997 $w=2.78e-07 $l=3.45e-07 $layer=LI1_cond $X=0.665 $Y=1.295
+ $X2=0.665 $Y2=0.95
r53 20 35 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.665 $Y=0.925
+ $X2=0.665 $Y2=0.95
r54 19 20 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.665 $Y=0.555
+ $X2=0.665 $Y2=0.925
r55 17 34 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.61 $Y=1.29
+ $X2=0.61 $Y2=0.95
r56 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.29
+ $X2=0.61 $Y2=1.455
r57 13 34 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.61 $Y=0.935
+ $X2=0.61 $Y2=0.95
r58 13 15 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.61 $Y=0.86
+ $X2=0.92 $Y2=0.86
r59 9 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.92 $Y=0.785
+ $X2=0.92 $Y2=0.86
r60 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.92 $Y=0.785
+ $X2=0.92 $Y2=0.465
r61 5 7 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=0.88 $Y=2.235 $X2=0.88
+ $Y2=2.885
r62 3 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.805 $Y=2.16
+ $X2=0.88 $Y2=2.235
r63 3 4 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.805 $Y=2.16
+ $X2=0.595 $Y2=2.16
r64 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.52 $Y=2.085
+ $X2=0.595 $Y2=2.16
r65 2 18 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.52 $Y=2.085
+ $X2=0.52 $Y2=1.455
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_M%A2 3 5 9 12 13 14 15 16 17 18 19 26
c55 14 0 1.02376e-19 $X=1.275 $Y=2.565
r56 18 19 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.665
+ $X2=1.175 $Y2=2.035
r57 17 18 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.295
+ $X2=1.175 $Y2=1.665
r58 17 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.34 $X2=1.15 $Y2=1.34
r59 16 17 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=0.925
+ $X2=1.175 $Y2=1.295
r60 15 16 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=0.555
+ $X2=1.175 $Y2=0.925
r61 13 14 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.275 $Y=2.415
+ $X2=1.275 $Y2=2.565
r62 12 13 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.24 $Y=1.845
+ $X2=1.24 $Y2=2.415
r63 11 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.15 $Y=1.68
+ $X2=1.15 $Y2=1.34
r64 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.68
+ $X2=1.15 $Y2=1.845
r65 10 26 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.34
r66 9 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.31 $Y=2.885
+ $X2=1.31 $Y2=2.565
r67 3 10 21.6467 $w=3.34e-07 $l=2.04939e-07 $layer=POLY_cond $X=1.28 $Y=1.145
+ $X2=1.15 $Y2=1.295
r68 3 5 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.28 $Y=1.145 $X2=1.28
+ $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_M%A1 3 7 11 12 13 14 15 20
c47 3 0 1.00777e-19 $X=1.64 $Y=0.465
r48 14 15 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=2.035
r49 14 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69 $Y=1.7
+ $X2=1.69 $Y2=1.7
r50 13 14 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.295
+ $X2=1.685 $Y2=1.665
r51 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.69 $Y=2.04
+ $X2=1.69 $Y2=1.7
r52 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=2.04
+ $X2=1.69 $Y2=2.205
r53 10 20 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.535
+ $X2=1.69 $Y2=1.7
r54 7 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.74 $Y=2.885
+ $X2=1.74 $Y2=2.205
r55 3 10 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.64 $Y=0.465
+ $X2=1.64 $Y2=1.535
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_M%B1 3 8 10 11 13 14 15 16 17 18 23
c51 8 0 1.023e-19 $X=2.17 $Y=2.885
r52 17 18 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=2.035
r53 16 17 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.195 $Y=1.295
+ $X2=2.195 $Y2=1.665
r54 16 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23
+ $Y=1.375 $X2=2.23 $Y2=1.375
r55 14 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.23 $Y=1.715
+ $X2=2.23 $Y2=1.375
r56 14 15 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.715
+ $X2=2.23 $Y2=1.88
r57 13 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.21
+ $X2=2.23 $Y2=1.375
r58 11 13 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=2.14 $Y=0.935
+ $X2=2.14 $Y2=1.21
r59 10 11 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.105 $Y=0.785
+ $X2=2.105 $Y2=0.935
r60 8 15 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=2.17 $Y=2.885
+ $X2=2.17 $Y2=1.88
r61 3 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.07 $Y=0.465
+ $X2=2.07 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_M%C1 1 3 6 8 9 13 14 16 17 18 19 20 26
c44 6 0 1.07821e-19 $X=2.53 $Y=2.885
r45 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.77
+ $Y=1.765 $X2=2.77 $Y2=1.765
r46 19 20 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.705 $Y=2.035
+ $X2=2.705 $Y2=2.405
r47 19 27 10.372 $w=2.98e-07 $l=2.7e-07 $layer=LI1_cond $X=2.705 $Y=2.035
+ $X2=2.705 $Y2=1.765
r48 18 27 3.84148 $w=2.98e-07 $l=1e-07 $layer=LI1_cond $X=2.705 $Y=1.665
+ $X2=2.705 $Y2=1.765
r49 17 18 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.705 $Y=1.295
+ $X2=2.705 $Y2=1.665
r50 16 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.6
+ $X2=2.77 $Y2=1.765
r51 13 26 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.77 $Y=2.12
+ $X2=2.77 $Y2=1.765
r52 13 14 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.695 $Y=2.12
+ $X2=2.695 $Y2=2.27
r53 10 16 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=2.86 $Y=0.935
+ $X2=2.86 $Y2=1.6
r54 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.785 $Y=0.86
+ $X2=2.86 $Y2=0.935
r55 8 9 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.785 $Y=0.86
+ $X2=2.575 $Y2=0.86
r56 6 14 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.53 $Y=2.885
+ $X2=2.53 $Y2=2.27
r57 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.5 $Y=0.785
+ $X2=2.575 $Y2=0.86
r58 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.5 $Y=0.785 $X2=2.5
+ $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_M%VPWR 1 2 7 9 13 16 17 18 28 29
c42 29 0 2.67233e-20 $X=3.12 $Y=3.33
r43 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 23 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 20 32 3.52379 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=3.33
+ $X2=0.172 $Y2=3.33
r49 20 22 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=0.345 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 18 29 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 18 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 18 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 16 22 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.42 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 16 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.42 $Y=3.33
+ $X2=1.515 $Y2=3.33
r55 15 25 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.61 $Y=3.33 $X2=1.68
+ $Y2=3.33
r56 15 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.515 $Y2=3.33
r57 11 17 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.515 $Y=3.245
+ $X2=1.515 $Y2=3.33
r58 11 13 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=1.515 $Y=3.245
+ $X2=1.515 $Y2=2.97
r59 7 32 3.3201 $w=1.9e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.25 $Y=3.245
+ $X2=0.172 $Y2=3.33
r60 7 9 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.25 $Y=3.245
+ $X2=0.25 $Y2=2.95
r61 2 13 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.385
+ $Y=2.675 $X2=1.525 $Y2=2.97
r62 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.675 $X2=0.26 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_M%A_191_535# 1 2 9 11 12 13
c36 13 0 7.56524e-20 $X=1.955 $Y=2.54
c37 11 0 1.023e-19 $X=1.79 $Y=2.54
r38 13 16 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.955 $Y=2.54
+ $X2=1.955 $Y2=2.82
r39 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=2.54
+ $X2=1.955 $Y2=2.54
r40 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.79 $Y=2.54 $X2=1.2
+ $Y2=2.54
r41 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.095 $Y=2.625
+ $X2=1.2 $Y2=2.54
r42 7 9 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=1.095 $Y=2.625
+ $X2=1.095 $Y2=2.8
r43 2 16 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.815
+ $Y=2.675 $X2=1.955 $Y2=2.82
r44 1 9 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.955
+ $Y=2.675 $X2=1.095 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_M%Y 1 2 3 12 15 16 18 19 20 21 22 33 35 52
c42 22 0 1.07821e-19 $X=3.12 $Y=2.775
c43 12 0 2.61001e-19 $X=1.855 $Y=0.53
r44 51 52 7.50345 $w=4.88e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.61
+ $X2=2.63 $Y2=0.61
r45 32 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.12 $Y=0.855 $X2=3.12
+ $Y2=0.925
r46 22 33 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=2.835
+ $X2=3.12 $Y2=2.67
r47 22 47 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=3.035 $Y=2.835
+ $X2=2.75 $Y2=2.835
r48 21 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.12 $Y=2.405
+ $X2=3.12 $Y2=2.67
r49 20 21 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=2.035
+ $X2=3.12 $Y2=2.405
r50 19 20 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=2.035
r51 18 19 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.665
r52 16 32 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=3.12 $Y=0.61
+ $X2=3.12 $Y2=0.855
r53 16 51 9.88595 $w=4.88e-07 $l=4.05e-07 $layer=LI1_cond $X=3.12 $Y=0.61
+ $X2=2.715 $Y2=0.61
r54 16 18 23.6824 $w=1.68e-07 $l=3.63e-07 $layer=LI1_cond $X=3.12 $Y=0.932
+ $X2=3.12 $Y2=1.295
r55 16 35 0.456684 $w=1.68e-07 $l=7e-09 $layer=LI1_cond $X=3.12 $Y=0.932
+ $X2=3.12 $Y2=0.925
r56 15 52 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.94 $Y=0.77 $X2=2.63
+ $Y2=0.77
r57 10 15 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.845 $Y=0.685
+ $X2=1.94 $Y2=0.77
r58 10 12 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.845 $Y=0.685
+ $X2=1.845 $Y2=0.53
r59 3 47 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=2.605
+ $Y=2.675 $X2=2.75 $Y2=2.835
r60 2 51 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.255 $X2=2.715 $Y2=0.53
r61 1 12 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.255 $X2=1.855 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_M%VGND 1 2 7 9 13 15 17 24 25 31
r37 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 25 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r40 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.285
+ $Y2=0
r42 22 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=3.12
+ $Y2=0
r43 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r44 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 18 28 3.52379 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r46 18 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.72
+ $Y2=0
r47 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.285
+ $Y2=0
r48 17 20 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.12 $Y=0 $X2=0.72
+ $Y2=0
r49 15 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r50 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r51 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.285 $Y=0.085
+ $X2=2.285 $Y2=0
r52 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.285 $Y=0.085
+ $X2=2.285 $Y2=0.4
r53 7 28 3.3201 $w=1.9e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.25 $Y=0.085
+ $X2=0.172 $Y2=0
r54 7 9 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=0.25 $Y=0.085
+ $X2=0.25 $Y2=0.4
r55 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.255 $X2=2.285 $Y2=0.4
r56 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.255 $X2=0.26 $Y2=0.4
.ends

