* NGSPICE file created from sky130_fd_sc_lp__nand4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
M1000 VPWR A_N a_27_51# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.1895e+12p pd=2.933e+07u as=3.339e+11p ps=3.05e+06u
M1001 a_217_51# a_27_51# Y VNB nshort w=840000u l=150000u
+  ad=1.1508e+12p pd=1.114e+07u as=4.704e+11p ps=4.48e+06u
M1002 a_644_51# B a_217_51# VNB nshort w=840000u l=150000u
+  ad=1.0752e+12p pd=9.28e+06u as=0p ps=0u
M1003 a_1025_65# C a_644_51# VNB nshort w=840000u l=150000u
+  ad=1.1844e+12p pd=1.122e+07u as=0p ps=0u
M1004 VPWR C Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=2.8224e+12p ps=2.464e+07u
M1005 a_217_51# a_27_51# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR D Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_27_51# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y a_27_51# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_217_51# B a_644_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D a_1025_65# VNB nshort w=840000u l=150000u
+  ad=6.93e+11p pd=6.69e+06u as=0p ps=0u
M1013 a_644_51# B a_217_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1025_65# C a_644_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND D a_1025_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y D VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y a_27_51# a_217_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y C VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y a_27_51# a_217_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y a_27_51# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y D VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_217_51# B a_644_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1025_65# D VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_644_51# C a_1025_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_27_51# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A_N a_27_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1028 a_644_51# C a_1025_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR D Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR C Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1025_65# D VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

