* File: sky130_fd_sc_lp__o221a_0.spice
* Created: Fri Aug 28 11:07:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221a_0.pex.spice"
.subckt sky130_fd_sc_lp__o221a_0  VNB VPB C1 B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1008 N_A_127_106#_M1008_d N_C1_M1008_g N_A_32_484#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_A_213_106#_M1007_d N_B1_M1007_g N_A_127_106#_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_127_106#_M1000_d N_B2_M1000_g N_A_213_106#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_213_106#_M1001_d N_A2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A1_M1009_g N_A_213_106#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07665 AS=0.0588 PD=0.785 PS=0.7 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1010 N_X_M1010_d N_A_32_484#_M1010_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.07665 PD=1.37 PS=0.785 NRD=0 NRS=11.424 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_C1_M1005_g N_A_32_484#_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1984 AS=0.1696 PD=1.26 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003 A=0.096 P=1.58 MULT=1
MM1003 A_269_484# N_B1_M1003_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1984 PD=0.85 PS=1.26 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1002 N_A_32_484#_M1002_d N_B2_M1002_g A_269_484# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=16.9223 NRS=15.3857 M=1 R=4.26667
+ SA=75001.3 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1011 A_449_484# N_A2_M1011_g N_A_32_484#_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1248 PD=0.85 PS=1.03 NRD=15.3857 NRS=16.9223 M=1 R=4.26667
+ SA=75001.9 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_449_484# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1984 AS=0.0672 PD=1.26 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75002.2
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1006 N_X_M1006_d N_A_32_484#_M1006_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1984 PD=1.81 PS=1.26 NRD=0 NRS=0 M=1 R=4.26667 SA=75003
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o221a_0.pxi.spice"
*
.ends
*
*
