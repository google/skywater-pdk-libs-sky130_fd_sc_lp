* File: sky130_fd_sc_lp__a311oi_1.pex.spice
* Created: Fri Aug 28 09:58:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311OI_1%A3 3 6 8 9 13 15
r23 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.74 $Y=1.355
+ $X2=0.74 $Y2=1.52
r24 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.74 $Y=1.355
+ $X2=0.74 $Y2=1.19
r25 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.74
+ $Y=1.355 $X2=0.74 $Y2=1.355
r26 8 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.355 $X2=0.72
+ $Y2=1.355
r27 6 16 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=0.83 $Y=2.465
+ $X2=0.83 $Y2=1.52
r28 3 15 171.913 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.83 $Y=0.655
+ $X2=0.83 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_1%A2 3 6 8 11 13
r34 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.28 $Y=1.355
+ $X2=1.28 $Y2=1.52
r35 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.28 $Y=1.355
+ $X2=1.28 $Y2=1.19
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.28
+ $Y=1.355 $X2=1.28 $Y2=1.355
r37 6 14 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.285 $Y=2.465
+ $X2=1.285 $Y2=1.52
r38 3 13 171.913 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.275 $Y=0.655
+ $X2=1.275 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_1%A1 1 3 6 8 14 15
r30 13 15 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.82 $Y=1.355
+ $X2=1.94 $Y2=1.355
r31 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.355 $X2=1.82 $Y2=1.355
r32 10 13 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.73 $Y=1.355 $X2=1.82
+ $Y2=1.355
r33 8 14 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=1.68 $Y=1.352
+ $X2=1.82 $Y2=1.352
r34 4 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.94 $Y=1.52
+ $X2=1.94 $Y2=1.355
r35 4 6 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.94 $Y=1.52 $X2=1.94
+ $Y2=2.465
r36 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.73 $Y=1.19
+ $X2=1.73 $Y2=1.355
r37 1 3 171.913 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.73 $Y=1.19 $X2=1.73
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_1%B1 1 3 6 8 14 15
r32 13 15 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.39 $Y=1.35
+ $X2=2.525 $Y2=1.35
r33 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.39
+ $Y=1.35 $X2=2.39 $Y2=1.35
r34 10 13 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.3 $Y=1.35 $X2=2.39
+ $Y2=1.35
r35 8 14 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=1.35 $X2=2.39
+ $Y2=1.35
r36 4 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.525 $Y=1.515
+ $X2=2.525 $Y2=1.35
r37 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.525 $Y=1.515
+ $X2=2.525 $Y2=2.465
r38 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.185 $X2=2.3
+ $Y2=1.35
r39 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.3 $Y=1.185 $X2=2.3
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_1%C1 1 3 6 8 13
r26 10 13 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.885 $Y=1.35
+ $X2=3.07 $Y2=1.35
r27 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.35 $X2=3.07 $Y2=1.35
r28 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.515
+ $X2=2.885 $Y2=1.35
r29 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.885 $Y=1.515
+ $X2=2.885 $Y2=2.465
r30 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.185
+ $X2=2.885 $Y2=1.35
r31 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.885 $Y=1.185
+ $X2=2.885 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_1%VPWR 1 2 9 15 20 21 22 28 37 38 41
r40 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r43 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 32 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=3.33
+ $X2=1.625 $Y2=3.33
r45 32 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.79 $Y=3.33 $X2=2.16
+ $Y2=3.33
r46 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 28 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=3.33
+ $X2=1.625 $Y2=3.33
r48 28 30 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.46 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 26 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 22 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 22 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 20 25 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.615 $Y2=3.33
r56 19 30 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.78 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=3.33
+ $X2=0.615 $Y2=3.33
r58 15 18 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=1.625 $Y=2.115
+ $X2=1.625 $Y2=2.95
r59 13 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=3.245
+ $X2=1.625 $Y2=3.33
r60 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.625 $Y=3.245
+ $X2=1.625 $Y2=2.95
r61 9 12 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=0.615 $Y=1.98
+ $X2=0.615 $Y2=2.95
r62 7 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.615 $Y=3.245
+ $X2=0.615 $Y2=3.33
r63 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.615 $Y=3.245
+ $X2=0.615 $Y2=2.95
r64 2 18 400 $w=1.7e-07 $l=1.24044e-06 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.625 $Y2=2.95
r65 2 15 400 $w=1.7e-07 $l=3.90641e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.625 $Y2=2.115
r66 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.49
+ $Y=1.835 $X2=0.615 $Y2=2.95
r67 1 9 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.49
+ $Y=1.835 $X2=0.615 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_1%A_181_367# 1 2 9 13 14 17
r33 17 19 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=2.24 $Y=1.98
+ $X2=2.24 $Y2=2.91
r34 15 17 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.24 $Y=1.86 $X2=2.24
+ $Y2=1.98
r35 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.075 $Y=1.775
+ $X2=2.24 $Y2=1.86
r36 13 14 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.075 $Y=1.775
+ $X2=1.235 $Y2=1.775
r37 9 11 37.606 $w=2.83e-07 $l=9.3e-07 $layer=LI1_cond $X=1.092 $Y=1.98
+ $X2=1.092 $Y2=2.91
r38 7 14 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=1.092 $Y=1.86
+ $X2=1.235 $Y2=1.775
r39 7 9 4.85239 $w=2.83e-07 $l=1.2e-07 $layer=LI1_cond $X=1.092 $Y=1.86
+ $X2=1.092 $Y2=1.98
r40 2 19 400 $w=1.7e-07 $l=1.18216e-06 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.835 $X2=2.24 $Y2=2.91
r41 2 17 400 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.835 $X2=2.24 $Y2=1.98
r42 1 11 400 $w=1.7e-07 $l=1.15456e-06 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.835 $X2=1.07 $Y2=2.91
r43 1 9 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=0.905
+ $Y=1.835 $X2=1.07 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_1%Y 1 2 3 11 12 14 22 23 24 25 26 35 41 46 49
r57 41 46 0.316883 $w=1.73e-07 $l=5e-09 $layer=LI1_cond $X=2.645 $Y=0.927
+ $X2=2.64 $Y2=0.927
r58 35 53 3.30495 $w=7.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.865 $Y=0.635
+ $X2=2.075 $Y2=0.635
r59 26 58 23.4494 $w=1.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.1 $Y=0.927
+ $X2=2.73 $Y2=0.927
r60 26 49 12.3876 $w=4.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.1 $Y=0.84 $X2=3.1
+ $Y2=0.38
r61 25 58 2.85195 $w=1.73e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=0.927
+ $X2=2.73 $Y2=0.927
r62 25 41 2.53506 $w=1.73e-07 $l=4e-08 $layer=LI1_cond $X=2.685 $Y=0.927
+ $X2=2.645 $Y2=0.927
r63 25 46 2.53506 $w=1.73e-07 $l=4e-08 $layer=LI1_cond $X=2.6 $Y=0.927 $X2=2.64
+ $Y2=0.927
r64 24 53 1.33772 $w=7.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.635
+ $X2=2.075 $Y2=0.635
r65 24 25 14.651 $w=3.43e-07 $l=3.55e-07 $layer=LI1_cond $X=2.245 $Y=0.927
+ $X2=2.6 $Y2=0.927
r66 23 35 2.91151 $w=7.58e-07 $l=1.85e-07 $layer=LI1_cond $X=1.68 $Y=0.635
+ $X2=1.865 $Y2=0.635
r67 22 23 7.55418 $w=7.58e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.635
+ $X2=1.68 $Y2=0.635
r68 14 16 36.3313 $w=2.93e-07 $l=9.3e-07 $layer=LI1_cond $X=3.117 $Y=1.98
+ $X2=3.117 $Y2=2.91
r69 12 18 25.2481 $w=1.68e-07 $l=3.87e-07 $layer=LI1_cond $X=3.117 $Y=1.79
+ $X2=2.73 $Y2=1.79
r70 12 14 4.10192 $w=2.93e-07 $l=1.05e-07 $layer=LI1_cond $X=3.117 $Y=1.875
+ $X2=3.117 $Y2=1.98
r71 11 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=1.705
+ $X2=2.73 $Y2=1.79
r72 10 58 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=2.73 $Y=1.015
+ $X2=2.73 $Y2=0.927
r73 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.73 $Y=1.015
+ $X2=2.73 $Y2=1.705
r74 3 16 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.91
r75 3 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=1.98
r76 2 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.38
r77 1 53 91 $w=1.7e-07 $l=3.81838e-07 $layer=licon1_NDIFF $count=2 $X=1.805
+ $Y=0.235 $X2=2.075 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_1%VGND 1 2 9 13 15 17 22 29 30 33 36
r39 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r42 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=2.59
+ $Y2=0
r44 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=3.12
+ $Y2=0
r45 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r46 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r47 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=0 $X2=0.615
+ $Y2=0
r48 23 25 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.78 $Y=0 $X2=2.16
+ $Y2=0
r49 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.59
+ $Y2=0
r50 22 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.16
+ $Y2=0
r51 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r52 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.615
+ $Y2=0
r54 17 19 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.24
+ $Y2=0
r55 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r56 15 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r57 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0
r58 11 13 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0.545
r59 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.615 $Y=0.085
+ $X2=0.615 $Y2=0
r60 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.615 $Y=0.085
+ $X2=0.615 $Y2=0.38
r61 2 13 182 $w=1.7e-07 $l=4.03423e-07 $layer=licon1_NDIFF $count=1 $X=2.375
+ $Y=0.235 $X2=2.59 $Y2=0.545
r62 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.49
+ $Y=0.235 $X2=0.615 $Y2=0.38
.ends

