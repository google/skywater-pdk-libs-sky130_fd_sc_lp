* File: sky130_fd_sc_lp__buflp_m.spice
* Created: Fri Aug 28 10:12:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__buflp_m.pex.spice"
.subckt sky130_fd_sc_lp__buflp_m  VNB VPB A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1004 A_120_120# N_A_90_94#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_90_94#_M1001_g A_120_120# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1000 A_278_120# N_A_M1000_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_90_94#_M1005_d N_A_M1005_g A_278_120# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_120_490# N_A_90_94#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_90_94#_M1007_g A_120_490# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0798 AS=0.0504 PD=0.8 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 A_304_490# N_A_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0504
+ AS=0.0798 PD=0.66 PS=0.8 NRD=30.4759 NRS=46.886 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_90_94#_M1006_d N_A_M1006_g A_304_490# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__buflp_m.pxi.spice"
*
.ends
*
*
