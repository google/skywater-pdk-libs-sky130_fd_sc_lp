* File: sky130_fd_sc_lp__o31ai_4.pex.spice
* Created: Wed Sep  2 10:25:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31AI_4%A2 3 6 10 14 18 22 26 30 36 39 43 45 48 57
+ 60 63
c115 39 0 1.13296e-19 $X=0.495 $Y=1.16
c116 30 0 1.49848e-19 $X=3.595 $Y=2.465
c117 26 0 1.73643e-19 $X=3.595 $Y=0.655
r118 54 63 8.27948 $w=4.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.825 $Y=1.29
+ $X2=2.985 $Y2=1.29
r119 53 55 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.825 $Y=1.42
+ $X2=3.165 $Y2=1.42
r120 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.825
+ $Y=1.42 $X2=2.825 $Y2=1.42
r121 50 53 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.735 $Y=1.42
+ $X2=2.825 $Y2=1.42
r122 45 54 4.95819 $w=4.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.64 $Y=1.29
+ $X2=2.825 $Y2=1.29
r123 45 60 9.18691 $w=4.28e-07 $l=1.8e-07 $layer=LI1_cond $X=2.64 $Y=1.29
+ $X2=2.46 $Y2=1.29
r124 43 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r125 43 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.185
r126 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.495
+ $Y=1.35 $X2=0.495 $Y2=1.35
r127 39 42 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.495 $Y=1.16
+ $X2=0.495 $Y2=1.35
r128 37 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.505 $Y=1.42
+ $X2=3.595 $Y2=1.42
r129 37 55 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.505 $Y=1.42
+ $X2=3.165 $Y2=1.42
r130 36 63 32.0404 $w=1.78e-07 $l=5.2e-07 $layer=LI1_cond $X=3.505 $Y=1.415
+ $X2=2.985 $Y2=1.415
r131 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.505
+ $Y=1.42 $X2=3.505 $Y2=1.42
r132 33 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.66 $Y=1.16
+ $X2=0.495 $Y2=1.16
r133 33 60 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=0.66 $Y=1.16
+ $X2=2.46 $Y2=1.16
r134 28 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.585
+ $X2=3.595 $Y2=1.42
r135 28 30 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.595 $Y=1.585
+ $X2=3.595 $Y2=2.465
r136 24 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.255
+ $X2=3.595 $Y2=1.42
r137 24 26 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.595 $Y=1.255
+ $X2=3.595 $Y2=0.655
r138 20 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.585
+ $X2=3.165 $Y2=1.42
r139 20 22 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.165 $Y=1.585
+ $X2=3.165 $Y2=2.465
r140 16 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.255
+ $X2=3.165 $Y2=1.42
r141 16 18 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.165 $Y=1.255
+ $X2=3.165 $Y2=0.655
r142 12 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.585
+ $X2=2.735 $Y2=1.42
r143 12 14 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=2.735 $Y=1.585
+ $X2=2.735 $Y2=2.465
r144 8 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.255
+ $X2=2.735 $Y2=1.42
r145 8 10 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.735 $Y=1.255
+ $X2=2.735 $Y2=0.655
r146 6 49 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.585 $Y=2.465
+ $X2=0.585 $Y2=1.515
r147 3 48 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.585 $Y=0.655
+ $X2=0.585 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_4%A1 3 7 11 15 19 23 27 31 40 43 53 56 59
c93 53 0 1.13296e-19 $X=2.305 $Y=1.51
r94 50 59 4.50999 $w=3.33e-07 $l=5e-08 $layer=LI1_cond $X=1.785 $Y=1.592
+ $X2=1.835 $Y2=1.592
r95 49 51 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.785 $Y=1.51
+ $X2=1.875 $Y2=1.51
r96 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.785
+ $Y=1.51 $X2=1.785 $Y2=1.51
r97 43 50 3.61213 $w=3.33e-07 $l=1.05e-07 $layer=LI1_cond $X=1.68 $Y=1.592
+ $X2=1.785 $Y2=1.592
r98 43 56 9.49817 $w=3.33e-07 $l=1.95e-07 $layer=LI1_cond $X=1.68 $Y=1.592
+ $X2=1.485 $Y2=1.592
r99 41 53 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.125 $Y=1.51
+ $X2=2.305 $Y2=1.51
r100 41 51 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.125 $Y=1.51
+ $X2=1.875 $Y2=1.51
r101 40 59 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.125 $Y=1.51
+ $X2=1.835 $Y2=1.51
r102 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.51 $X2=2.125 $Y2=1.51
r103 36 49 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.445 $Y=1.51
+ $X2=1.785 $Y2=1.51
r104 36 45 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.445 $Y=1.51
+ $X2=1.015 $Y2=1.51
r105 35 56 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.445 $Y=1.51
+ $X2=1.485 $Y2=1.51
r106 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.445
+ $Y=1.51 $X2=1.445 $Y2=1.51
r107 29 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.675
+ $X2=2.305 $Y2=1.51
r108 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.305 $Y=1.675
+ $X2=2.305 $Y2=2.465
r109 25 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.345
+ $X2=2.305 $Y2=1.51
r110 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.305 $Y=1.345
+ $X2=2.305 $Y2=0.655
r111 21 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.675
+ $X2=1.875 $Y2=1.51
r112 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.875 $Y=1.675
+ $X2=1.875 $Y2=2.465
r113 17 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.345
+ $X2=1.875 $Y2=1.51
r114 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.875 $Y=1.345
+ $X2=1.875 $Y2=0.655
r115 13 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=1.51
r116 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=2.465
r117 9 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.345
+ $X2=1.445 $Y2=1.51
r118 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.445 $Y=1.345
+ $X2=1.445 $Y2=0.655
r119 5 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=1.51
r120 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=2.465
r121 1 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.345
+ $X2=1.015 $Y2=1.51
r122 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.015 $Y=1.345
+ $X2=1.015 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_4%A3 1 3 4 6 7 9 10 12 13 15 16 18 21 25 27 30
+ 31 33 34 36 40 41 42 51
c132 40 0 1.98746e-19 $X=5.005 $Y=1.595
c133 36 0 1.49848e-19 $X=4.735 $Y=1.595
c134 34 0 1.11345e-19 $X=7.555 $Y=1.44
c135 4 0 2.93317e-20 $X=4.025 $Y=1.725
r136 51 52 6.29478 $w=5.36e-07 $l=7e-08 $layer=POLY_cond $X=4.885 $Y=1.455
+ $X2=4.955 $Y2=1.455
r137 47 49 26.528 $w=5.36e-07 $l=2.95e-07 $layer=POLY_cond $X=4.16 $Y=1.455
+ $X2=4.455 $Y2=1.455
r138 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.16
+ $Y=1.51 $X2=4.16 $Y2=1.51
r139 45 47 12.1399 $w=5.36e-07 $l=1.35e-07 $layer=POLY_cond $X=4.025 $Y=1.455
+ $X2=4.16 $Y2=1.455
r140 42 48 8.85984 $w=5.38e-07 $l=4e-07 $layer=LI1_cond $X=4.56 $Y=1.595
+ $X2=4.16 $Y2=1.595
r141 41 48 1.77197 $w=5.38e-07 $l=8e-08 $layer=LI1_cond $X=4.08 $Y=1.595
+ $X2=4.16 $Y2=1.595
r142 39 51 4.04664 $w=5.36e-07 $l=4.5e-08 $layer=POLY_cond $X=4.84 $Y=1.455
+ $X2=4.885 $Y2=1.455
r143 39 49 34.6213 $w=5.36e-07 $l=3.85e-07 $layer=POLY_cond $X=4.84 $Y=1.455
+ $X2=4.455 $Y2=1.455
r144 38 40 9.76796 $w=5.38e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=1.595
+ $X2=5.005 $Y2=1.595
r145 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.84
+ $Y=1.51 $X2=4.84 $Y2=1.51
r146 36 42 3.87618 $w=5.38e-07 $l=1.75e-07 $layer=LI1_cond $X=4.735 $Y=1.595
+ $X2=4.56 $Y2=1.595
r147 36 38 2.32571 $w=5.38e-07 $l=1.05e-07 $layer=LI1_cond $X=4.735 $Y=1.595
+ $X2=4.84 $Y2=1.595
r148 34 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.555 $Y=1.44
+ $X2=7.555 $Y2=1.605
r149 34 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.555 $Y=1.44
+ $X2=7.555 $Y2=1.275
r150 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.555
+ $Y=1.44 $X2=7.555 $Y2=1.44
r151 31 33 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=7.28 $Y=1.435
+ $X2=7.555 $Y2=1.435
r152 29 31 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=7.195 $Y=1.535
+ $X2=7.28 $Y2=1.435
r153 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.195 $Y=1.535
+ $X2=7.195 $Y2=1.695
r154 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.11 $Y=1.78
+ $X2=7.195 $Y2=1.695
r155 27 40 137.332 $w=1.68e-07 $l=2.105e-06 $layer=LI1_cond $X=7.11 $Y=1.78
+ $X2=5.005 $Y2=1.78
r156 25 55 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.635 $Y=2.465
+ $X2=7.635 $Y2=1.605
r157 21 54 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.475 $Y=0.655
+ $X2=7.475 $Y2=1.275
r158 16 52 33.1734 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.955 $Y=1.185
+ $X2=4.955 $Y2=1.455
r159 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.955 $Y=1.185
+ $X2=4.955 $Y2=0.655
r160 13 51 33.1734 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.885 $Y=1.725
+ $X2=4.885 $Y2=1.455
r161 13 15 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.885 $Y=1.725
+ $X2=4.885 $Y2=2.465
r162 10 49 33.1734 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.455 $Y=1.725
+ $X2=4.455 $Y2=1.455
r163 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.455 $Y=1.725
+ $X2=4.455 $Y2=2.465
r164 7 49 33.1734 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.455 $Y=1.185
+ $X2=4.455 $Y2=1.455
r165 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.455 $Y=1.185
+ $X2=4.455 $Y2=0.655
r166 4 45 33.1734 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.025 $Y=1.725
+ $X2=4.025 $Y2=1.455
r167 4 6 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.025 $Y=1.725
+ $X2=4.025 $Y2=2.465
r168 1 45 33.1734 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.025 $Y=1.185
+ $X2=4.025 $Y2=1.455
r169 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.025 $Y=1.185
+ $X2=4.025 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_4%B1 1 3 6 10 12 14 17 19 21 24 26 28 31 34 35
+ 36 58 60 61 70 73 75
c93 31 0 1.11345e-19 $X=6.765 $Y=1.43
r94 61 70 3.65789 $w=3.25e-07 $l=7.7e-08 $layer=LI1_cond $X=5.597 $Y=1.362
+ $X2=5.52 $Y2=1.362
r95 58 59 6.42667 $w=4.5e-07 $l=6e-08 $layer=POLY_cond $X=7.045 $Y=1.495
+ $X2=7.105 $Y2=1.495
r96 55 73 1.95029 $w=3.23e-07 $l=5.5e-08 $layer=LI1_cond $X=6.425 $Y=1.362
+ $X2=6.48 $Y2=1.362
r97 55 60 0.425517 $w=3.23e-07 $l=1.2e-08 $layer=LI1_cond $X=6.425 $Y=1.362
+ $X2=6.413 $Y2=1.362
r98 54 56 2.14222 $w=4.5e-07 $l=2e-08 $layer=POLY_cond $X=6.425 $Y=1.495
+ $X2=6.445 $Y2=1.495
r99 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.425
+ $Y=1.43 $X2=6.425 $Y2=1.43
r100 52 54 19.28 $w=4.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.245 $Y=1.495
+ $X2=6.425 $Y2=1.495
r101 50 52 17.1378 $w=4.5e-07 $l=1.6e-07 $layer=POLY_cond $X=6.085 $Y=1.495
+ $X2=6.245 $Y2=1.495
r102 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.085
+ $Y=1.43 $X2=6.085 $Y2=1.43
r103 48 50 7.49778 $w=4.5e-07 $l=7e-08 $layer=POLY_cond $X=6.015 $Y=1.495
+ $X2=6.085 $Y2=1.495
r104 47 48 21.4222 $w=4.5e-07 $l=2e-07 $layer=POLY_cond $X=5.815 $Y=1.495
+ $X2=6.015 $Y2=1.495
r105 45 47 7.49778 $w=4.5e-07 $l=7e-08 $layer=POLY_cond $X=5.745 $Y=1.495
+ $X2=5.815 $Y2=1.495
r106 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.745
+ $Y=1.43 $X2=5.745 $Y2=1.43
r107 43 45 38.56 $w=4.5e-07 $l=3.6e-07 $layer=POLY_cond $X=5.385 $Y=1.495
+ $X2=5.745 $Y2=1.495
r108 42 43 7.49778 $w=4.5e-07 $l=7e-08 $layer=POLY_cond $X=5.315 $Y=1.495
+ $X2=5.385 $Y2=1.495
r109 36 75 5.32593 $w=3.23e-07 $l=8.6e-08 $layer=LI1_cond $X=6.489 $Y=1.362
+ $X2=6.575 $Y2=1.362
r110 36 73 0.319138 $w=3.23e-07 $l=9e-09 $layer=LI1_cond $X=6.489 $Y=1.362
+ $X2=6.48 $Y2=1.362
r111 36 60 0.319138 $w=3.23e-07 $l=9e-09 $layer=LI1_cond $X=6.404 $Y=1.362
+ $X2=6.413 $Y2=1.362
r112 36 51 11.3117 $w=3.23e-07 $l=3.19e-07 $layer=LI1_cond $X=6.404 $Y=1.362
+ $X2=6.085 $Y2=1.362
r113 35 51 3.01408 $w=3.23e-07 $l=8.5e-08 $layer=LI1_cond $X=6 $Y=1.362
+ $X2=6.085 $Y2=1.362
r114 35 46 9.04224 $w=3.23e-07 $l=2.55e-07 $layer=LI1_cond $X=6 $Y=1.362
+ $X2=5.745 $Y2=1.362
r115 34 70 0.199184 $w=2.45e-07 $l=4e-09 $layer=LI1_cond $X=5.516 $Y=1.362
+ $X2=5.52 $Y2=1.362
r116 34 46 5.10621 $w=3.23e-07 $l=1.44e-07 $layer=LI1_cond $X=5.601 $Y=1.362
+ $X2=5.745 $Y2=1.362
r117 34 61 0.141839 $w=3.23e-07 $l=4e-09 $layer=LI1_cond $X=5.601 $Y=1.362
+ $X2=5.597 $Y2=1.362
r118 32 58 29.9911 $w=4.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.765 $Y=1.495
+ $X2=7.045 $Y2=1.495
r119 32 56 34.2756 $w=4.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.765 $Y=1.495
+ $X2=6.445 $Y2=1.495
r120 31 75 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=6.765 $Y=1.435
+ $X2=6.575 $Y2=1.435
r121 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.765
+ $Y=1.43 $X2=6.765 $Y2=1.43
r122 26 59 28.7666 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=7.105 $Y=1.725
+ $X2=7.105 $Y2=1.495
r123 26 28 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.105 $Y=1.725
+ $X2=7.105 $Y2=2.465
r124 22 58 28.7666 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=7.045 $Y=1.265
+ $X2=7.045 $Y2=1.495
r125 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.045 $Y=1.265
+ $X2=7.045 $Y2=0.655
r126 19 56 28.7666 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.445 $Y=1.725
+ $X2=6.445 $Y2=1.495
r127 19 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.445 $Y=1.725
+ $X2=6.445 $Y2=2.465
r128 15 52 28.7666 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.245 $Y=1.265
+ $X2=6.245 $Y2=1.495
r129 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.245 $Y=1.265
+ $X2=6.245 $Y2=0.655
r130 12 48 28.7666 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.015 $Y=1.725
+ $X2=6.015 $Y2=1.495
r131 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.015 $Y=1.725
+ $X2=6.015 $Y2=2.465
r132 8 47 28.7666 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.815 $Y=1.265
+ $X2=5.815 $Y2=1.495
r133 8 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.815 $Y=1.265
+ $X2=5.815 $Y2=0.655
r134 4 43 28.7666 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.385 $Y=1.265
+ $X2=5.385 $Y2=1.495
r135 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.385 $Y=1.265
+ $X2=5.385 $Y2=0.655
r136 1 42 28.7666 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.315 $Y=1.725
+ $X2=5.315 $Y2=1.495
r137 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.315 $Y=1.725
+ $X2=5.315 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_4%A_49_367# 1 2 3 4 5 16 18 20 22 24 28 33 35
+ 36 40 42 45 46 47 49 50 51 52 54 58 62 67 68 71
c149 71 0 2.93317e-20 $X=4.67 $Y=2.985
c150 4 0 1.98746e-19 $X=4.53 $Y=1.835
r151 62 64 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.09 $Y=1.9
+ $X2=2.09 $Y2=2.015
r152 58 60 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.23 $Y=1.9
+ $X2=1.23 $Y2=2.015
r153 52 73 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=2.895
+ $X2=7.93 $Y2=2.98
r154 52 54 30.3624 $w=2.58e-07 $l=6.85e-07 $layer=LI1_cond $X=7.93 $Y=2.895
+ $X2=7.93 $Y2=2.21
r155 50 73 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.8 $Y=2.98 $X2=7.93
+ $Y2=2.98
r156 50 51 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.8 $Y=2.98
+ $X2=7.165 $Y2=2.98
r157 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.08 $Y=2.895
+ $X2=7.165 $Y2=2.98
r158 48 49 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.08 $Y=2.58
+ $X2=7.08 $Y2=2.895
r159 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.995 $Y=2.495
+ $X2=7.08 $Y2=2.58
r160 46 47 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=6.995 $Y=2.495
+ $X2=5.525 $Y2=2.495
r161 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.44 $Y=2.58
+ $X2=5.525 $Y2=2.495
r162 44 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.44 $Y=2.58
+ $X2=5.44 $Y2=2.895
r163 43 71 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=2.985
+ $X2=4.67 $Y2=2.985
r164 42 45 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.355 $Y=2.985
+ $X2=5.44 $Y2=2.895
r165 42 43 32.0404 $w=1.78e-07 $l=5.2e-07 $layer=LI1_cond $X=5.355 $Y=2.985
+ $X2=4.835 $Y2=2.985
r166 38 71 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.67 $Y=2.895
+ $X2=4.67 $Y2=2.985
r167 38 40 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.67 $Y=2.895
+ $X2=4.67 $Y2=2.47
r168 37 70 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=2.99
+ $X2=3.81 $Y2=2.99
r169 36 71 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.505 $Y=2.99
+ $X2=4.67 $Y2=2.985
r170 36 37 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.505 $Y=2.99
+ $X2=3.975 $Y2=2.99
r171 35 68 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=2.2
+ $X2=3.81 $Y2=2.035
r172 33 70 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.81 $Y2=2.99
r173 33 35 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.81 $Y2=2.2
r174 30 68 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.73 $Y=1.875
+ $X2=3.73 $Y2=2.035
r175 29 67 6.36606 $w=1.7e-07 $l=2.32164e-07 $layer=LI1_cond $X=3.075 $Y=1.79
+ $X2=2.855 $Y2=1.815
r176 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.645 $Y=1.79
+ $X2=3.73 $Y2=1.875
r177 28 29 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.645 $Y=1.79
+ $X2=3.075 $Y2=1.79
r178 25 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=1.9
+ $X2=2.09 $Y2=1.9
r179 24 67 6.36606 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=1.9
+ $X2=2.855 $Y2=1.815
r180 24 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.855 $Y=1.9
+ $X2=2.175 $Y2=1.9
r181 23 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=2.015
+ $X2=1.23 $Y2=2.015
r182 22 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=2.015
+ $X2=2.09 $Y2=2.015
r183 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.005 $Y=2.015
+ $X2=1.315 $Y2=2.015
r184 21 57 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.465 $Y=1.9
+ $X2=0.335 $Y2=1.9
r185 20 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.9
+ $X2=1.23 $Y2=1.9
r186 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.145 $Y=1.9
+ $X2=0.465 $Y2=1.9
r187 16 57 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.335 $Y=1.985
+ $X2=0.335 $Y2=1.9
r188 16 18 41.0004 $w=2.58e-07 $l=9.25e-07 $layer=LI1_cond $X=0.335 $Y=1.985
+ $X2=0.335 $Y2=2.91
r189 5 73 400 $w=1.7e-07 $l=1.1538e-06 $layer=licon1_PDIFF $count=1 $X=7.71
+ $Y=1.835 $X2=7.895 $Y2=2.9
r190 5 54 400 $w=1.7e-07 $l=4.58258e-07 $layer=licon1_PDIFF $count=1 $X=7.71
+ $Y=1.835 $X2=7.895 $Y2=2.21
r191 4 40 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=4.53
+ $Y=1.835 $X2=4.67 $Y2=2.47
r192 3 70 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=1.835 $X2=3.81 $Y2=2.91
r193 3 35 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=1.835 $X2=3.81 $Y2=2.2
r194 2 67 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.81
+ $Y=1.835 $X2=2.95 $Y2=1.98
r195 1 57 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=1.98
r196 1 18 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_4%A_132_367# 1 2 3 4 15 17 21 24 25 27 29 32
+ 36 38
r55 38 40 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.52 $Y=2.24
+ $X2=2.52 $Y2=2.355
r56 32 34 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.8 $Y=2.24 $X2=0.8
+ $Y2=2.355
r57 27 44 3.12017 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.36 $Y=2.885
+ $X2=3.36 $Y2=2.98
r58 27 29 33.3206 $w=2.28e-07 $l=6.65e-07 $layer=LI1_cond $X=3.36 $Y=2.885
+ $X2=3.36 $Y2=2.22
r59 26 42 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=2.98
+ $X2=2.52 $Y2=2.98
r60 25 44 3.77705 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=3.245 $Y=2.98
+ $X2=3.36 $Y2=2.98
r61 25 26 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=3.245 $Y=2.98
+ $X2=2.685 $Y2=2.98
r62 24 42 2.73294 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.52 $Y=2.885
+ $X2=2.52 $Y2=2.98
r63 23 40 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.44
+ $X2=2.52 $Y2=2.355
r64 23 24 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.52 $Y=2.44
+ $X2=2.52 $Y2=2.885
r65 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=2.355
+ $X2=1.66 $Y2=2.355
r66 21 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=2.355
+ $X2=2.52 $Y2=2.355
r67 21 22 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.355 $Y=2.355
+ $X2=1.825 $Y2=2.355
r68 18 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=2.355
+ $X2=0.8 $Y2=2.355
r69 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=2.355
+ $X2=1.66 $Y2=2.355
r70 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.495 $Y=2.355
+ $X2=0.965 $Y2=2.355
r71 13 34 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=2.44 $X2=0.8
+ $Y2=2.355
r72 13 15 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.8 $Y=2.44 $X2=0.8
+ $Y2=2.95
r73 4 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=1.835 $X2=3.38 $Y2=2.91
r74 4 29 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=3.24
+ $Y=1.835 $X2=3.38 $Y2=2.22
r75 3 42 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.835 $X2=2.52 $Y2=2.97
r76 3 38 400 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.835 $X2=2.52 $Y2=2.24
r77 2 36 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=1.52
+ $Y=1.835 $X2=1.66 $Y2=2.435
r78 1 32 400 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=2.24
r79 1 15 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_4%VPWR 1 2 3 4 15 19 23 27 30 31 33 34 35 37
+ 42 58 59 62 65
r117 65 66 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r120 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r121 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r122 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r123 53 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r125 50 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r126 49 50 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r127 47 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=2.09 $Y2=3.33
r128 47 49 217.578 $w=1.68e-07 $l=3.335e-06 $layer=LI1_cond $X=2.185 $Y=3.33
+ $X2=5.52 $Y2=3.33
r129 46 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 46 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r131 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r132 43 62 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.23 $Y2=3.33
r133 43 45 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.325 $Y=3.33
+ $X2=1.68 $Y2=3.33
r134 42 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.09 $Y2=3.33
r135 42 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r136 40 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r137 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r138 37 62 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=1.23 $Y2=3.33
r139 37 39 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=0.24 $Y2=3.33
r140 35 50 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.52 $Y2=3.33
r141 35 66 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 33 52 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.555 $Y=3.33
+ $X2=6.48 $Y2=3.33
r143 33 34 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.555 $Y=3.33
+ $X2=6.69 $Y2=3.33
r144 32 55 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.96 $Y2=3.33
r145 32 34 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.825 $Y=3.33
+ $X2=6.69 $Y2=3.33
r146 30 49 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.695 $Y=3.33
+ $X2=5.52 $Y2=3.33
r147 30 31 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.695 $Y=3.33
+ $X2=5.8 $Y2=3.33
r148 29 52 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.905 $Y=3.33
+ $X2=6.48 $Y2=3.33
r149 29 31 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.905 $Y=3.33
+ $X2=5.8 $Y2=3.33
r150 25 34 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.69 $Y=3.245
+ $X2=6.69 $Y2=3.33
r151 25 27 14.0854 $w=2.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.69 $Y=3.245
+ $X2=6.69 $Y2=2.915
r152 21 31 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=3.245
+ $X2=5.8 $Y2=3.33
r153 21 23 17.4286 $w=2.08e-07 $l=3.3e-07 $layer=LI1_cond $X=5.8 $Y=3.245
+ $X2=5.8 $Y2=2.915
r154 17 65 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=3.245
+ $X2=2.09 $Y2=3.33
r155 17 19 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=2.09 $Y=3.245
+ $X2=2.09 $Y2=2.775
r156 13 62 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r157 13 15 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.775
r158 4 27 600 $w=1.7e-07 $l=1.17576e-06 $layer=licon1_PDIFF $count=1 $X=6.52
+ $Y=1.835 $X2=6.72 $Y2=2.915
r159 3 23 600 $w=1.7e-07 $l=1.26854e-06 $layer=licon1_PDIFF $count=1 $X=5.39
+ $Y=1.835 $X2=5.8 $Y2=2.915
r160 2 19 600 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=1.95
+ $Y=1.835 $X2=2.09 $Y2=2.775
r161 1 15 600 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.835 $X2=1.23 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_4%Y 1 2 3 4 5 6 21 25 35 38 39 40 42 44 46 49
+ 50 53 54
r98 51 54 6.44587 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=7.482 $Y=2.24
+ $X2=7.482 $Y2=2.405
r99 51 53 4.64645 $w=2.32e-07 $l=1.03e-07 $layer=LI1_cond $X=7.482 $Y=2.24
+ $X2=7.482 $Y2=2.137
r100 48 50 7.50811 $w=4.63e-07 $l=9.5e-08 $layer=LI1_cond $X=6.83 $Y=0.932
+ $X2=6.925 $Y2=0.932
r101 48 49 3.21092 $w=4.63e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=0.932
+ $X2=6.745 $Y2=0.932
r102 41 42 32.3735 $w=1.83e-07 $l=5.4e-07 $layer=LI1_cond $X=7.982 $Y=1.165
+ $X2=7.982 $Y2=1.705
r103 39 42 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.89 $Y=1.79
+ $X2=7.982 $Y2=1.705
r104 39 40 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.89 $Y=1.79
+ $X2=7.63 $Y2=1.79
r105 38 53 4.64645 $w=2.32e-07 $l=1.2973e-07 $layer=LI1_cond $X=7.545 $Y=2.035
+ $X2=7.482 $Y2=2.137
r106 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.545 $Y=1.875
+ $X2=7.63 $Y2=1.79
r107 37 38 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.545 $Y=1.875
+ $X2=7.545 $Y2=2.035
r108 35 41 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.89 $Y=1.08
+ $X2=7.982 $Y2=1.165
r109 35 50 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=7.89 $Y=1.08
+ $X2=6.925 $Y2=1.08
r110 34 49 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=6.46 $Y=0.865
+ $X2=6.745 $Y2=0.865
r111 31 34 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.6 $Y=0.865
+ $X2=6.46 $Y2=0.865
r112 26 46 4.88354 $w=1.92e-07 $l=9e-08 $layer=LI1_cond $X=5.185 $Y=2.137
+ $X2=5.095 $Y2=2.137
r113 26 28 56.5366 $w=2.03e-07 $l=1.045e-06 $layer=LI1_cond $X=5.185 $Y=2.137
+ $X2=6.23 $Y2=2.137
r114 25 53 1.79954 $w=2.05e-07 $l=1.47e-07 $layer=LI1_cond $X=7.335 $Y=2.137
+ $X2=7.482 $Y2=2.137
r115 25 28 59.7827 $w=2.03e-07 $l=1.105e-06 $layer=LI1_cond $X=7.335 $Y=2.137
+ $X2=6.23 $Y2=2.137
r116 22 44 3.50369 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.335 $Y=2.125
+ $X2=4.24 $Y2=2.125
r117 21 46 4.88354 $w=1.92e-07 $l=9.58123e-08 $layer=LI1_cond $X=5.005 $Y=2.125
+ $X2=5.095 $Y2=2.137
r118 21 22 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=5.005 $Y=2.125
+ $X2=4.335 $Y2=2.125
r119 6 53 300 $w=1.7e-07 $l=4.80234e-07 $layer=licon1_PDIFF $count=2 $X=7.18
+ $Y=1.835 $X2=7.42 $Y2=2.21
r120 5 28 600 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=6.09
+ $Y=1.835 $X2=6.23 $Y2=2.14
r121 4 46 300 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=2 $X=4.96
+ $Y=1.835 $X2=5.1 $Y2=2.2
r122 3 44 300 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=2 $X=4.1
+ $Y=1.835 $X2=4.24 $Y2=2.2
r123 2 48 182 $w=1.7e-07 $l=8.47467e-07 $layer=licon1_NDIFF $count=1 $X=6.32
+ $Y=0.235 $X2=6.83 $Y2=0.865
r124 2 34 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=6.32
+ $Y=0.235 $X2=6.46 $Y2=0.865
r125 1 31 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.235 $X2=5.6 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 42 46
+ 48 50 53 54 55 56 57 59 64 76 88 91 94 98
r124 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r125 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r126 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r127 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r128 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r129 83 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r130 82 83 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r131 80 83 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=7.44
+ $Y2=0
r132 80 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r133 79 82 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.44
+ $Y2=0
r134 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r135 77 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.88 $Y=0 $X2=4.715
+ $Y2=0
r136 77 79 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.88 $Y=0 $X2=5.04
+ $Y2=0
r137 76 97 4.53846 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=7.605 $Y=0
+ $X2=7.882 $Y2=0
r138 76 82 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=0
+ $X2=7.44 $Y2=0
r139 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r140 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r141 72 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r142 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r143 69 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.255 $Y=0 $X2=2.09
+ $Y2=0
r144 69 71 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.255 $Y=0
+ $X2=2.64 $Y2=0
r145 68 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r146 68 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r147 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r148 65 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=0 $X2=1.23
+ $Y2=0
r149 65 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=0
+ $X2=1.68 $Y2=0
r150 64 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=2.09
+ $Y2=0
r151 64 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=1.68
+ $Y2=0
r152 63 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r153 63 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r154 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r155 60 85 3.99156 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=0
+ $X2=0.232 $Y2=0
r156 60 62 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.465 $Y=0
+ $X2=0.72 $Y2=0
r157 59 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.23
+ $Y2=0
r158 59 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r159 57 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r160 57 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r161 55 74 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.6
+ $Y2=0
r162 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=0 $X2=3.81
+ $Y2=0
r163 53 71 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.785 $Y=0
+ $X2=2.64 $Y2=0
r164 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.785 $Y=0 $X2=2.95
+ $Y2=0
r165 52 74 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.6
+ $Y2=0
r166 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=2.95
+ $Y2=0
r167 48 97 3.22771 $w=3.3e-07 $l=1.4854e-07 $layer=LI1_cond $X=7.77 $Y=0.085
+ $X2=7.882 $Y2=0
r168 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.77 $Y=0.085
+ $X2=7.77 $Y2=0.38
r169 44 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.715 $Y=0.085
+ $X2=4.715 $Y2=0
r170 44 46 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.715 $Y=0.085
+ $X2=4.715 $Y2=0.36
r171 43 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=0 $X2=3.81
+ $Y2=0
r172 42 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.55 $Y=0 $X2=4.715
+ $Y2=0
r173 42 43 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.55 $Y=0
+ $X2=3.975 $Y2=0
r174 38 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=0.085
+ $X2=3.81 $Y2=0
r175 38 40 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.81 $Y=0.085
+ $X2=3.81 $Y2=0.36
r176 34 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=0.085
+ $X2=2.95 $Y2=0
r177 34 36 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.95 $Y=0.085
+ $X2=2.95 $Y2=0.44
r178 30 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=0.085
+ $X2=2.09 $Y2=0
r179 30 32 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.09 $Y=0.085
+ $X2=2.09 $Y2=0.44
r180 26 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0
r181 26 28 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0.44
r182 22 85 3.22066 $w=2.6e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.232 $Y2=0
r183 22 24 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.38
r184 7 50 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=7.55
+ $Y=0.235 $X2=7.77 $Y2=0.38
r185 6 46 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=4.53
+ $Y=0.235 $X2=4.715 $Y2=0.36
r186 5 40 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.67
+ $Y=0.235 $X2=3.81 $Y2=0.36
r187 4 36 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.235 $X2=2.95 $Y2=0.44
r188 3 32 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.235 $X2=2.09 $Y2=0.44
r189 2 28 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.44
r190 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_4%A_132_47# 1 2 3 4 5 6 7 8 25 27 29 33 35 39
+ 41 45 47 51 53 55 59 66 68 69 75 79
c99 69 0 1.73643e-19 $X=3.375 $Y=0.82
r100 79 81 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=7.26 $Y=0.37
+ $X2=7.26 $Y2=0.392
r101 72 73 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=3.375 $Y=0.93
+ $X2=3.375 $Y2=1.07
r102 69 72 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=3.375 $Y=0.82 $X2=3.375
+ $Y2=0.93
r103 69 70 4.75232 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=0.82
+ $X2=3.375 $Y2=0.735
r104 60 77 2.95793 $w=2.75e-07 $l=1e-07 $layer=LI1_cond $X=5.265 $Y=0.392
+ $X2=5.165 $Y2=0.392
r105 60 62 32.0589 $w=2.73e-07 $l=7.65e-07 $layer=LI1_cond $X=5.265 $Y=0.392
+ $X2=6.03 $Y2=0.392
r106 59 81 1.82517 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=0.392
+ $X2=7.26 $Y2=0.392
r107 59 62 44.631 $w=2.73e-07 $l=1.065e-06 $layer=LI1_cond $X=7.095 $Y=0.392
+ $X2=6.03 $Y2=0.392
r108 56 58 3.05 $w=1.98e-07 $l=5.5e-08 $layer=LI1_cond $X=5.165 $Y=0.985
+ $X2=5.165 $Y2=0.93
r109 55 77 4.08194 $w=2e-07 $l=1.38e-07 $layer=LI1_cond $X=5.165 $Y=0.53
+ $X2=5.165 $Y2=0.392
r110 55 58 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=5.165 $Y=0.53
+ $X2=5.165 $Y2=0.93
r111 54 75 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=4.38 $Y=1.07
+ $X2=4.267 $Y2=1.07
r112 53 56 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.065 $Y=1.07
+ $X2=5.165 $Y2=0.985
r113 53 54 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.065 $Y=1.07
+ $X2=4.38 $Y2=1.07
r114 49 75 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.267 $Y=0.985
+ $X2=4.267 $Y2=1.07
r115 49 51 20.2318 $w=2.23e-07 $l=3.95e-07 $layer=LI1_cond $X=4.267 $Y=0.985
+ $X2=4.267 $Y2=0.59
r116 48 73 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.475 $Y=1.07
+ $X2=3.375 $Y2=1.07
r117 47 75 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=4.155 $Y=1.07
+ $X2=4.267 $Y2=1.07
r118 47 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.155 $Y=1.07
+ $X2=3.475 $Y2=1.07
r119 45 70 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=3.38 $Y=0.42
+ $X2=3.38 $Y2=0.735
r120 42 68 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.615 $Y=0.82
+ $X2=2.52 $Y2=0.82
r121 41 69 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.275 $Y=0.82
+ $X2=3.375 $Y2=0.82
r122 41 42 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.275 $Y=0.82
+ $X2=2.615 $Y2=0.82
r123 37 68 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=0.735
+ $X2=2.52 $Y2=0.82
r124 37 39 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=2.52 $Y=0.735
+ $X2=2.52 $Y2=0.42
r125 36 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.755 $Y=0.82
+ $X2=1.66 $Y2=0.82
r126 35 68 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.425 $Y=0.82
+ $X2=2.52 $Y2=0.82
r127 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.425 $Y=0.82
+ $X2=1.755 $Y2=0.82
r128 31 66 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=0.735
+ $X2=1.66 $Y2=0.82
r129 31 33 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=1.66 $Y=0.735
+ $X2=1.66 $Y2=0.42
r130 30 64 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.895 $Y=0.82
+ $X2=0.765 $Y2=0.82
r131 29 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.565 $Y=0.82
+ $X2=1.66 $Y2=0.82
r132 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=0.82
+ $X2=0.895 $Y2=0.82
r133 25 64 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.735
+ $X2=0.765 $Y2=0.82
r134 25 27 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.765 $Y=0.735
+ $X2=0.765 $Y2=0.42
r135 8 79 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=7.12
+ $Y=0.235 $X2=7.26 $Y2=0.37
r136 7 62 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.89
+ $Y=0.235 $X2=6.03 $Y2=0.38
r137 6 77 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.235 $X2=5.17 $Y2=0.42
r138 6 58 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.235 $X2=5.17 $Y2=0.93
r139 5 51 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=4.1
+ $Y=0.235 $X2=4.24 $Y2=0.59
r140 4 72 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.235 $X2=3.38 $Y2=0.93
r141 4 45 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.235 $X2=3.38 $Y2=0.42
r142 3 68 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.52 $Y2=0.82
r143 3 39 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.235 $X2=2.52 $Y2=0.42
r144 2 66 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.235 $X2=1.66 $Y2=0.82
r145 2 33 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.235 $X2=1.66 $Y2=0.42
r146 1 64 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.235 $X2=0.8 $Y2=0.82
r147 1 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.235 $X2=0.8 $Y2=0.42
.ends

