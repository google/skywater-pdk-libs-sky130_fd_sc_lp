* File: sky130_fd_sc_lp__clkinvlp_8.pxi.spice
* Created: Wed Sep  2 09:41:26 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINVLP_8%A N_A_M1014_g N_A_M1000_g N_A_M1001_g
+ N_A_M1002_g N_A_M1004_g N_A_M1005_g N_A_M1003_g N_A_M1013_g N_A_M1006_g
+ N_A_M1007_g N_A_M1008_g N_A_M1009_g N_A_M1011_g N_A_M1010_g N_A_c_81_n
+ N_A_M1012_g N_A_M1015_g A A PM_SKY130_FD_SC_LP__CLKINVLP_8%A
x_PM_SKY130_FD_SC_LP__CLKINVLP_8%VPWR N_VPWR_M1000_s N_VPWR_M1002_s
+ N_VPWR_M1006_s N_VPWR_M1011_s N_VPWR_M1015_s N_VPWR_c_209_n N_VPWR_c_210_n
+ N_VPWR_c_211_n N_VPWR_c_212_n N_VPWR_c_213_n N_VPWR_c_214_n N_VPWR_c_215_n
+ N_VPWR_c_216_n N_VPWR_c_217_n N_VPWR_c_218_n N_VPWR_c_219_n N_VPWR_c_220_n
+ VPWR N_VPWR_c_221_n N_VPWR_c_222_n N_VPWR_c_208_n
+ PM_SKY130_FD_SC_LP__CLKINVLP_8%VPWR
x_PM_SKY130_FD_SC_LP__CLKINVLP_8%Y N_Y_M1001_s N_Y_M1007_s N_Y_M1000_d
+ N_Y_M1005_d N_Y_M1008_d N_Y_M1012_d N_Y_c_280_n N_Y_c_289_n N_Y_c_281_n
+ N_Y_c_282_n N_Y_c_290_n N_Y_c_283_n N_Y_c_284_n N_Y_c_291_n N_Y_c_285_n
+ N_Y_c_286_n Y Y Y Y Y Y PM_SKY130_FD_SC_LP__CLKINVLP_8%Y
x_PM_SKY130_FD_SC_LP__CLKINVLP_8%VGND N_VGND_M1014_d N_VGND_M1003_d
+ N_VGND_M1010_d N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n N_VGND_c_377_n
+ N_VGND_c_378_n N_VGND_c_379_n VGND N_VGND_c_380_n N_VGND_c_381_n
+ N_VGND_c_382_n N_VGND_c_383_n PM_SKY130_FD_SC_LP__CLKINVLP_8%VGND
cc_1 VNB N_A_M1014_g 0.0369914f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.61
cc_2 VNB N_A_M1000_g 0.00506355f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.48
cc_3 VNB N_A_M1001_g 0.0244252f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.61
cc_4 VNB N_A_M1002_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.48
cc_5 VNB N_A_M1004_g 0.0271804f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=0.61
cc_6 VNB N_A_M1005_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.48
cc_7 VNB N_A_M1003_g 0.0267708f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=0.61
cc_8 VNB N_A_M1013_g 0.0267565f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=0.61
cc_9 VNB N_A_M1006_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.48
cc_10 VNB N_A_M1007_g 0.0260215f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=0.61
cc_11 VNB N_A_M1008_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.48
cc_12 VNB N_A_M1009_g 0.0260215f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=0.61
cc_13 VNB N_A_M1011_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.48
cc_14 VNB N_A_M1010_g 0.0385356f $X=-0.19 $Y=-0.245 $X2=3.205 $Y2=0.61
cc_15 VNB N_A_c_81_n 0.259149f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=1.565
cc_16 VNB N_A_M1012_g 0.00509532f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=2.48
cc_17 VNB N_A_M1015_g 0.00795919f $X=-0.19 $Y=-0.245 $X2=4.235 $Y2=2.48
cc_18 VNB A 0.0243288f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_VPWR_c_208_n 0.203486f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.407
cc_20 VNB N_Y_c_280_n 0.0105522f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=0.61
cc_21 VNB N_Y_c_281_n 0.0079368f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=0.61
cc_22 VNB N_Y_c_282_n 7.00526e-19 $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=0.61
cc_23 VNB N_Y_c_283_n 0.0295329f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=0.61
cc_24 VNB N_Y_c_284_n 0.00665756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_285_n 0.00345438f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.48
cc_26 VNB N_Y_c_286_n 0.00382697f $X=-0.19 $Y=-0.245 $X2=3.205 $Y2=1.235
cc_27 VNB Y 0.00607165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 2.3763e-19 $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=1.565
cc_29 VNB N_VGND_c_374_n 0.0111239f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.61
cc_30 VNB N_VGND_c_375_n 0.0257259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_376_n 0.00306361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_377_n 0.0254984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_378_n 0.0368108f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.48
cc_34 VNB N_VGND_c_379_n 0.00589254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_380_n 0.0340106f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=0.61
cc_36 VNB N_VGND_c_381_n 0.040807f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.48
cc_37 VNB N_VGND_c_382_n 0.327199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_383_n 0.00561514f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.48
cc_39 VPB N_A_M1000_g 0.0435143f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.48
cc_40 VPB N_A_M1002_g 0.0340581f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.48
cc_41 VPB N_A_M1005_g 0.0340581f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.48
cc_42 VPB N_A_M1006_g 0.0340581f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.48
cc_43 VPB N_A_M1008_g 0.0340581f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.48
cc_44 VPB N_A_M1011_g 0.0340581f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=2.48
cc_45 VPB N_A_M1012_g 0.0340581f $X=-0.19 $Y=1.655 $X2=3.705 $Y2=2.48
cc_46 VPB N_A_M1015_g 0.0461397f $X=-0.19 $Y=1.655 $X2=4.235 $Y2=2.48
cc_47 VPB A 0.00764565f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_48 VPB N_VPWR_c_209_n 0.0112117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_210_n 0.0508745f $X=-0.19 $Y=1.655 $X2=1.265 $Y2=0.61
cc_50 VPB N_VPWR_c_211_n 0.0199224f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.48
cc_51 VPB N_VPWR_c_212_n 0.00678226f $X=-0.19 $Y=1.655 $X2=1.625 $Y2=0.61
cc_52 VPB N_VPWR_c_213_n 0.00678226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_214_n 0.00678226f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=0.61
cc_54 VPB N_VPWR_c_215_n 0.0124877f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.48
cc_55 VPB N_VPWR_c_216_n 0.0608249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_217_n 0.0199224f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=1.565
cc_57 VPB N_VPWR_c_218_n 0.00577233f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=2.48
cc_58 VPB N_VPWR_c_219_n 0.0199224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_220_n 0.00577233f $X=-0.19 $Y=1.655 $X2=3.205 $Y2=1.235
cc_60 VPB N_VPWR_c_221_n 0.0199224f $X=-0.19 $Y=1.655 $X2=4.235 $Y2=2.48
cc_61 VPB N_VPWR_c_222_n 0.00577233f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.415
cc_62 VPB N_VPWR_c_208_n 0.0533656f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=1.407
cc_63 VPB N_Y_c_289_n 0.00232136f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.48
cc_64 VPB N_Y_c_290_n 0.00232136f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.48
cc_65 VPB N_Y_c_291_n 0.00232136f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.48
cc_66 VPB Y 0.00232136f $X=-0.19 $Y=1.655 $X2=3.705 $Y2=2.48
cc_67 N_A_M1000_g N_VPWR_c_210_n 0.0235557f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_68 N_A_M1002_g N_VPWR_c_210_n 8.05893e-19 $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_69 N_A_c_81_n N_VPWR_c_210_n 0.00122665f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_70 A N_VPWR_c_210_n 0.0288185f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_M1000_g N_VPWR_c_211_n 0.00687065f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_72 N_A_M1002_g N_VPWR_c_211_n 0.00687065f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_73 N_A_M1000_g N_VPWR_c_212_n 8.05893e-19 $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_74 N_A_M1002_g N_VPWR_c_212_n 0.0225326f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_75 N_A_M1005_g N_VPWR_c_212_n 0.0225326f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_76 N_A_M1006_g N_VPWR_c_212_n 8.05893e-19 $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_77 N_A_c_81_n N_VPWR_c_212_n 0.00233601f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_78 N_A_M1005_g N_VPWR_c_213_n 8.05893e-19 $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_79 N_A_M1006_g N_VPWR_c_213_n 0.0225326f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_80 N_A_M1008_g N_VPWR_c_213_n 0.0225326f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_81 N_A_M1011_g N_VPWR_c_213_n 8.05893e-19 $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_82 N_A_c_81_n N_VPWR_c_213_n 0.00233601f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_83 N_A_M1008_g N_VPWR_c_214_n 8.05893e-19 $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_84 N_A_M1011_g N_VPWR_c_214_n 0.0225326f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_85 N_A_c_81_n N_VPWR_c_214_n 0.00202524f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_86 N_A_M1012_g N_VPWR_c_214_n 0.0225326f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_87 N_A_M1015_g N_VPWR_c_214_n 8.05893e-19 $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_88 N_A_M1012_g N_VPWR_c_216_n 8.05893e-19 $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_89 N_A_M1015_g N_VPWR_c_216_n 0.0244443f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_90 N_A_M1005_g N_VPWR_c_217_n 0.00687065f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_91 N_A_M1006_g N_VPWR_c_217_n 0.00687065f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_92 N_A_M1008_g N_VPWR_c_219_n 0.00687065f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_93 N_A_M1011_g N_VPWR_c_219_n 0.00687065f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_94 N_A_M1012_g N_VPWR_c_221_n 0.00687065f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_95 N_A_M1015_g N_VPWR_c_221_n 0.00687065f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_96 N_A_M1000_g N_VPWR_c_208_n 0.0129282f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_97 N_A_M1002_g N_VPWR_c_208_n 0.0129282f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_98 N_A_M1005_g N_VPWR_c_208_n 0.0129282f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_99 N_A_M1006_g N_VPWR_c_208_n 0.0129282f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_100 N_A_M1008_g N_VPWR_c_208_n 0.0129282f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_101 N_A_M1011_g N_VPWR_c_208_n 0.0129282f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_102 N_A_M1012_g N_VPWR_c_208_n 0.0129282f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_103 N_A_M1015_g N_VPWR_c_208_n 0.0129282f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_104 N_A_M1004_g N_Y_c_280_n 0.00790787f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_105 N_A_M1003_g N_Y_c_280_n 0.00710902f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_106 N_A_c_81_n N_Y_c_280_n 0.0500081f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_107 N_A_M1002_g N_Y_c_289_n 0.00197414f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_108 N_A_M1005_g N_Y_c_289_n 0.0308281f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_109 N_A_M1006_g N_Y_c_289_n 0.0308281f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_110 N_A_M1008_g N_Y_c_289_n 0.00197414f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_111 N_A_M1013_g N_Y_c_281_n 0.00627067f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_112 N_A_M1007_g N_Y_c_281_n 0.00679033f $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_113 N_A_c_81_n N_Y_c_281_n 0.0283833f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_114 N_A_M1013_g N_Y_c_282_n 0.00300477f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_115 N_A_M1007_g N_Y_c_282_n 0.0176278f $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_116 N_A_M1009_g N_Y_c_282_n 0.0176278f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_117 N_A_M1010_g N_Y_c_282_n 0.00300477f $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_118 N_A_c_81_n N_Y_c_282_n 0.00101183f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_119 N_A_M1006_g N_Y_c_290_n 0.00197414f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_120 N_A_M1008_g N_Y_c_290_n 0.0308281f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_121 N_A_M1011_g N_Y_c_290_n 0.0308281f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_122 N_A_c_81_n N_Y_c_290_n 0.0035478f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_123 N_A_M1012_g N_Y_c_290_n 0.00197414f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_124 N_A_M1010_g N_Y_c_283_n 0.00845395f $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_125 N_A_c_81_n N_Y_c_283_n 0.0886231f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_126 N_A_M1007_g N_Y_c_284_n 6.18991e-19 $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_127 N_A_M1009_g N_Y_c_284_n 0.00750968f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_128 N_A_c_81_n N_Y_c_284_n 0.0336856f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_129 N_A_M1011_g N_Y_c_291_n 0.00197414f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_130 N_A_M1012_g N_Y_c_291_n 0.0308281f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_131 N_A_M1015_g N_Y_c_291_n 0.0411856f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_132 N_A_M1014_g N_Y_c_285_n 0.0034335f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_133 N_A_M1001_g N_Y_c_285_n 0.0116329f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_134 N_A_M1004_g N_Y_c_285_n 0.00895713f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_135 N_A_M1003_g N_Y_c_285_n 0.00126558f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_136 N_A_c_81_n N_Y_c_285_n 6.81418e-19 $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_137 N_A_M1003_g N_Y_c_286_n 8.7915e-19 $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_138 N_A_M1013_g N_Y_c_286_n 0.00173861f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_139 N_A_c_81_n N_Y_c_286_n 0.0141982f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_140 N_A_M1014_g Y 0.00885061f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_141 N_A_M1001_g Y 0.0107605f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_142 N_A_M1004_g Y 0.00702452f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_143 A Y 0.00711802f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A_M1014_g Y 2.69915e-19 $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_145 N_A_M1001_g Y 0.00122275f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_146 N_A_c_81_n Y 0.0182148f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_147 A Y 0.0298337f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A_M1000_g Y 0.0347043f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_149 N_A_M1002_g Y 0.0308281f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_150 N_A_M1005_g Y 0.00197414f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_151 N_A_c_81_n Y 3.96106e-19 $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_152 A Y 0.0161123f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_153 N_A_M1014_g N_VGND_c_375_n 0.0121806f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_154 N_A_M1001_g N_VGND_c_375_n 0.0010716f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_155 N_A_c_81_n N_VGND_c_375_n 0.00118321f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_156 A N_VGND_c_375_n 0.016704f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A_M1004_g N_VGND_c_376_n 0.00194234f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_158 N_A_M1003_g N_VGND_c_376_n 0.0129414f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_159 N_A_M1013_g N_VGND_c_376_n 0.0131259f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_160 N_A_M1007_g N_VGND_c_376_n 0.00223895f $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_161 N_A_c_81_n N_VGND_c_376_n 6.49557e-19 $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_162 N_A_M1009_g N_VGND_c_377_n 0.00223895f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_163 N_A_M1010_g N_VGND_c_377_n 0.0148579f $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_164 N_A_c_81_n N_VGND_c_377_n 0.00173776f $X=3.705 $Y=1.565 $X2=0 $Y2=0
cc_165 N_A_M1013_g N_VGND_c_378_n 0.00407525f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_166 N_A_M1007_g N_VGND_c_378_n 0.00464284f $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_167 N_A_M1009_g N_VGND_c_378_n 0.00464284f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_168 N_A_M1010_g N_VGND_c_378_n 0.00407525f $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_169 N_A_M1014_g N_VGND_c_380_n 0.00407525f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_170 N_A_M1001_g N_VGND_c_380_n 0.00306316f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_171 N_A_M1004_g N_VGND_c_380_n 0.00460068f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_172 N_A_M1003_g N_VGND_c_380_n 0.00407525f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_173 N_A_M1014_g N_VGND_c_382_n 0.00774993f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_174 N_A_M1001_g N_VGND_c_382_n 0.00413202f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_175 N_A_M1004_g N_VGND_c_382_n 0.00874311f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_176 N_A_M1003_g N_VGND_c_382_n 0.00774993f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_177 N_A_M1013_g N_VGND_c_382_n 0.00774993f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_178 N_A_M1007_g N_VGND_c_382_n 0.0088065f $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_179 N_A_M1009_g N_VGND_c_382_n 0.0088065f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_180 N_A_M1010_g N_VGND_c_382_n 0.00774993f $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_181 N_VPWR_c_212_n N_Y_c_280_n 0.0146643f $X=1.32 $Y=2.125 $X2=0 $Y2=0
cc_182 N_VPWR_c_212_n N_Y_c_289_n 0.0685263f $X=1.32 $Y=2.125 $X2=0 $Y2=0
cc_183 N_VPWR_c_213_n N_Y_c_289_n 0.0685263f $X=2.38 $Y=2.125 $X2=0 $Y2=0
cc_184 N_VPWR_c_217_n N_Y_c_289_n 0.0157615f $X=2.215 $Y=3.33 $X2=0 $Y2=0
cc_185 N_VPWR_c_208_n N_Y_c_289_n 0.0120285f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_186 N_VPWR_c_213_n N_Y_c_281_n 0.0146449f $X=2.38 $Y=2.125 $X2=0 $Y2=0
cc_187 N_VPWR_c_213_n N_Y_c_290_n 0.0685263f $X=2.38 $Y=2.125 $X2=0 $Y2=0
cc_188 N_VPWR_c_214_n N_Y_c_290_n 0.0685263f $X=3.44 $Y=2.125 $X2=0 $Y2=0
cc_189 N_VPWR_c_219_n N_Y_c_290_n 0.0157615f $X=3.275 $Y=3.33 $X2=0 $Y2=0
cc_190 N_VPWR_c_208_n N_Y_c_290_n 0.0120285f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_191 N_VPWR_c_214_n N_Y_c_283_n 0.0146643f $X=3.44 $Y=2.125 $X2=0 $Y2=0
cc_192 N_VPWR_c_214_n N_Y_c_291_n 0.0685263f $X=3.44 $Y=2.125 $X2=0 $Y2=0
cc_193 N_VPWR_c_216_n N_Y_c_291_n 0.0685263f $X=4.5 $Y=2.125 $X2=0 $Y2=0
cc_194 N_VPWR_c_221_n N_Y_c_291_n 0.0157615f $X=4.335 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_208_n N_Y_c_291_n 0.0120285f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_210_n Y 0.0685263f $X=0.26 $Y=2.125 $X2=0 $Y2=0
cc_197 N_VPWR_c_211_n Y 0.0157615f $X=1.155 $Y=3.33 $X2=0 $Y2=0
cc_198 N_VPWR_c_212_n Y 0.0685263f $X=1.32 $Y=2.125 $X2=0 $Y2=0
cc_199 N_VPWR_c_208_n Y 0.0120285f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_200 N_Y_c_285_n N_VGND_c_375_n 0.0330838f $X=1.05 $Y=0.545 $X2=0 $Y2=0
cc_201 N_Y_c_280_n N_VGND_c_376_n 3.29624e-19 $X=1.685 $Y=1.38 $X2=0 $Y2=0
cc_202 N_Y_c_282_n N_VGND_c_376_n 0.0110409f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_203 N_Y_c_285_n N_VGND_c_376_n 0.0161046f $X=1.05 $Y=0.545 $X2=0 $Y2=0
cc_204 N_Y_c_286_n N_VGND_c_376_n 0.0123519f $X=1.85 $Y=1.38 $X2=0 $Y2=0
cc_205 N_Y_c_282_n N_VGND_c_377_n 0.0110409f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_206 N_Y_c_283_n N_VGND_c_377_n 0.0135664f $X=3.805 $Y=1.38 $X2=0 $Y2=0
cc_207 N_Y_c_282_n N_VGND_c_378_n 0.00846545f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_208 N_Y_c_285_n N_VGND_c_380_n 0.0291015f $X=1.05 $Y=0.545 $X2=0 $Y2=0
cc_209 N_Y_c_282_n N_VGND_c_382_n 0.0111318f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_210 N_Y_c_285_n N_VGND_c_382_n 0.0211357f $X=1.05 $Y=0.545 $X2=0 $Y2=0
cc_211 N_Y_c_285_n A_268_67# 0.00418236f $X=1.05 $Y=0.545 $X2=-0.19 $Y2=-0.245
cc_212 Y A_268_67# 0.00148246f $X=0.635 $Y=0.84 $X2=-0.19 $Y2=-0.245
