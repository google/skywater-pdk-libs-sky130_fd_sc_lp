* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxtp_1 D GATE VGND VNB VPB VPWR Q
X0 VPWR GATE a_196_425# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 VPWR a_596_419# a_733_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR a_733_99# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_27_425# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_317_461# a_196_425# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_27_425# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_596_419# a_317_461# a_701_419# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_701_419# a_733_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND a_596_419# a_733_99# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_691_125# a_733_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_317_461# a_196_425# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VGND a_733_99# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VPWR a_27_425# a_524_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_524_419# a_196_425# a_596_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 VGND a_27_425# a_530_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_596_419# a_196_425# a_691_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND GATE a_196_425# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_530_125# a_317_461# a_596_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
