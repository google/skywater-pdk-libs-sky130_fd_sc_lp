* File: sky130_fd_sc_lp__a311o_m.pxi.spice
* Created: Wed Sep  2 09:25:27 2020
* 
x_PM_SKY130_FD_SC_LP__A311O_M%A3 N_A3_M1011_g N_A3_c_78_n N_A3_M1006_g
+ N_A3_c_79_n A3 A3 A3 N_A3_c_81_n N_A3_c_82_n PM_SKY130_FD_SC_LP__A311O_M%A3
x_PM_SKY130_FD_SC_LP__A311O_M%A2 N_A2_M1003_g N_A2_M1008_g N_A2_c_125_n
+ N_A2_c_130_n A2 A2 A2 A2 N_A2_c_127_n PM_SKY130_FD_SC_LP__A311O_M%A2
x_PM_SKY130_FD_SC_LP__A311O_M%A_54_154# N_A_54_154#_M1009_d N_A_54_154#_M1005_d
+ N_A_54_154#_M1007_d N_A_54_154#_c_170_n N_A_54_154#_M1002_g
+ N_A_54_154#_c_171_n N_A_54_154#_M1001_g N_A_54_154#_c_179_n
+ N_A_54_154#_c_180_n N_A_54_154#_c_172_n N_A_54_154#_c_181_n
+ N_A_54_154#_c_253_p N_A_54_154#_c_182_n N_A_54_154#_c_183_n
+ N_A_54_154#_c_173_n N_A_54_154#_c_174_n N_A_54_154#_c_175_n
+ N_A_54_154#_c_185_n N_A_54_154#_c_186_n N_A_54_154#_c_176_n
+ N_A_54_154#_c_221_p N_A_54_154#_c_217_p PM_SKY130_FD_SC_LP__A311O_M%A_54_154#
x_PM_SKY130_FD_SC_LP__A311O_M%A1 N_A1_M1009_g N_A1_M1010_g N_A1_c_266_n
+ N_A1_c_267_n A1 N_A1_c_269_n N_A1_c_270_n PM_SKY130_FD_SC_LP__A311O_M%A1
x_PM_SKY130_FD_SC_LP__A311O_M%B1 N_B1_M1000_g N_B1_M1004_g B1 N_B1_c_315_n
+ N_B1_c_316_n PM_SKY130_FD_SC_LP__A311O_M%B1
x_PM_SKY130_FD_SC_LP__A311O_M%C1 N_C1_c_345_n N_C1_M1005_g N_C1_M1007_g
+ N_C1_c_346_n N_C1_c_347_n C1 C1 N_C1_c_349_n PM_SKY130_FD_SC_LP__A311O_M%C1
x_PM_SKY130_FD_SC_LP__A311O_M%X N_X_M1001_s N_X_M1002_s X X X X X X X
+ N_X_c_377_n PM_SKY130_FD_SC_LP__A311O_M%X
x_PM_SKY130_FD_SC_LP__A311O_M%VPWR N_VPWR_M1002_d N_VPWR_M1003_d N_VPWR_c_397_n
+ N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n VPWR N_VPWR_c_401_n
+ N_VPWR_c_402_n N_VPWR_c_396_n N_VPWR_c_404_n PM_SKY130_FD_SC_LP__A311O_M%VPWR
x_PM_SKY130_FD_SC_LP__A311O_M%A_196_403# N_A_196_403#_M1011_d
+ N_A_196_403#_M1010_d N_A_196_403#_c_433_n N_A_196_403#_c_434_n
+ N_A_196_403#_c_435_n PM_SKY130_FD_SC_LP__A311O_M%A_196_403#
x_PM_SKY130_FD_SC_LP__A311O_M%VGND N_VGND_M1001_d N_VGND_M1000_d N_VGND_c_457_n
+ N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n VGND N_VGND_c_461_n
+ N_VGND_c_462_n N_VGND_c_463_n N_VGND_c_464_n PM_SKY130_FD_SC_LP__A311O_M%VGND
cc_1 VNB N_A3_M1011_g 0.00826568f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.225
cc_2 VNB N_A3_c_78_n 0.016321f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.77
cc_3 VNB N_A3_c_79_n 0.0178591f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.845
cc_4 VNB A3 0.00787142f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_5 VNB N_A3_c_81_n 0.0314055f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.325
cc_6 VNB N_A3_c_82_n 0.0129372f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.16
cc_7 VNB N_A2_M1008_g 0.0299598f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.77
cc_8 VNB N_A2_c_125_n 0.0204448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A2 0.0117985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_c_127_n 0.0153251f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.325
cc_11 VNB N_A_54_154#_c_170_n 0.0438372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_54_154#_c_171_n 0.0196201f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_13 VNB N_A_54_154#_c_172_n 0.0295026f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.16
cc_14 VNB N_A_54_154#_c_173_n 0.00784514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_54_154#_c_174_n 0.00374527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_54_154#_c_175_n 0.015448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_54_154#_c_176_n 0.00456282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_266_n 0.0159305f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.845
cc_19 VNB N_A1_c_267_n 0.014266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A1 0.00248824f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.845
cc_21 VNB N_A1_c_269_n 0.0161222f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_22 VNB N_A1_c_270_n 0.0302024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_M1000_g 0.0242967f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.225
cc_24 VNB N_B1_M1004_g 0.0219513f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.77
cc_25 VNB N_B1_c_315_n 0.0335356f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.845
cc_26 VNB N_B1_c_316_n 0.00667366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_C1_c_345_n 0.0205557f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.49
cc_28 VNB N_C1_c_346_n 0.0274469f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.45
cc_29 VNB N_C1_c_347_n 0.032924f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.845
cc_30 VNB C1 0.00706972f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_31 VNB N_C1_c_349_n 0.0721809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_377_n 0.0547246f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.325
cc_33 VNB N_VPWR_c_396_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_457_n 0.00298318f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.45
cc_35 VNB N_VGND_c_458_n 0.00311149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_459_n 0.0356383f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_37 VNB N_VGND_c_460_n 0.00525414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_461_n 0.0182881f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.325
cc_39 VNB N_VGND_c_462_n 0.0244078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_463_n 0.199068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_464_n 0.00514068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_A3_M1011_g 0.0294387f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.225
cc_43 VPB A3 0.00417425f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_44 VPB N_A2_M1003_g 0.0212393f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.225
cc_45 VPB N_A2_c_125_n 5.60561e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A2_c_130_n 0.0153139f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=0.845
cc_47 VPB A2 0.00140821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_54_154#_c_170_n 0.00462091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_54_154#_M1002_g 0.0440355f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_50 VPB N_A_54_154#_c_179_n 0.111851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_54_154#_c_180_n 0.0153564f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=1.325
cc_52 VPB N_A_54_154#_c_181_n 0.0223422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_54_154#_c_182_n 0.0208829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_54_154#_c_183_n 0.0485238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_54_154#_c_175_n 0.00313933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_54_154#_c_185_n 0.0199126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_54_154#_c_186_n 0.0101823f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A1_M1010_g 0.0210635f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=0.45
cc_59 VPB A1 0.00297171f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=0.845
cc_60 VPB N_A1_c_269_n 0.0151477f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_61 VPB N_B1_M1004_g 0.028546f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=0.77
cc_62 VPB N_C1_M1007_g 0.03789f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.16
cc_63 VPB C1 0.00933024f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_64 VPB N_X_c_377_n 0.0326541f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=1.325
cc_65 VPB N_VPWR_c_397_n 0.0158483f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=0.45
cc_66 VPB N_VPWR_c_398_n 0.0242156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_399_n 0.019485f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_68 VPB N_VPWR_c_400_n 0.00334761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_401_n 0.0207436f $X=-0.19 $Y=1.655 $X2=0.825 $Y2=1.49
cc_70 VPB N_VPWR_c_402_n 0.0448221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_396_n 0.0721382f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_404_n 0.00583335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_196_403#_c_433_n 0.00957398f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=0.77
cc_74 VPB N_A_196_403#_c_434_n 0.0058693f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=0.45
cc_75 VPB N_A_196_403#_c_435_n 0.0026221f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_76 N_A3_M1011_g N_A2_M1003_g 0.0172167f $X=0.905 $Y=2.225 $X2=0 $Y2=0
cc_77 N_A3_c_78_n N_A2_M1008_g 0.0496798f $X=1.025 $Y=0.77 $X2=0 $Y2=0
cc_78 A3 N_A2_M1008_g 2.61429e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_79 N_A3_c_82_n N_A2_M1008_g 0.00801504f $X=0.825 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A3_M1011_g N_A2_c_125_n 0.0197437f $X=0.905 $Y=2.225 $X2=0 $Y2=0
cc_81 N_A3_M1011_g A2 0.00163739f $X=0.905 $Y=2.225 $X2=0 $Y2=0
cc_82 N_A3_c_78_n A2 0.0065281f $X=1.025 $Y=0.77 $X2=0 $Y2=0
cc_83 A3 A2 0.0628587f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A3_c_82_n A2 0.00408437f $X=0.825 $Y=1.16 $X2=0 $Y2=0
cc_85 A3 N_A2_c_127_n 5.64874e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_86 N_A3_c_81_n N_A2_c_127_n 0.0204708f $X=0.825 $Y=1.325 $X2=0 $Y2=0
cc_87 N_A3_M1011_g N_A_54_154#_c_170_n 0.0063672f $X=0.905 $Y=2.225 $X2=0 $Y2=0
cc_88 A3 N_A_54_154#_c_170_n 0.0029948f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_89 N_A3_c_81_n N_A_54_154#_c_170_n 0.018078f $X=0.825 $Y=1.325 $X2=0 $Y2=0
cc_90 N_A3_c_82_n N_A_54_154#_c_170_n 0.00612201f $X=0.825 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A3_c_78_n N_A_54_154#_c_171_n 0.0120052f $X=1.025 $Y=0.77 $X2=0 $Y2=0
cc_92 N_A3_M1011_g N_A_54_154#_c_179_n 0.00564446f $X=0.905 $Y=2.225 $X2=0 $Y2=0
cc_93 N_A3_c_79_n N_A_54_154#_c_172_n 0.00954687f $X=1.025 $Y=0.845 $X2=0 $Y2=0
cc_94 A3 N_A_54_154#_c_172_n 6.88108e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_95 N_A3_M1011_g N_A_54_154#_c_181_n 0.0206502f $X=0.905 $Y=2.225 $X2=0 $Y2=0
cc_96 N_A3_M1011_g N_X_c_377_n 0.00216016f $X=0.905 $Y=2.225 $X2=0 $Y2=0
cc_97 N_A3_c_79_n N_X_c_377_n 3.70204e-19 $X=1.025 $Y=0.845 $X2=0 $Y2=0
cc_98 A3 N_X_c_377_n 0.0630437f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_99 N_A3_c_81_n N_X_c_377_n 0.00107569f $X=0.825 $Y=1.325 $X2=0 $Y2=0
cc_100 N_A3_c_82_n N_X_c_377_n 6.00969e-19 $X=0.825 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A3_M1011_g N_VPWR_c_397_n 0.0017832f $X=0.905 $Y=2.225 $X2=0 $Y2=0
cc_102 A3 N_VPWR_c_397_n 0.00769989f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_103 N_A3_c_81_n N_VPWR_c_397_n 5.55141e-19 $X=0.825 $Y=1.325 $X2=0 $Y2=0
cc_104 N_A3_M1011_g N_VPWR_c_396_n 8.50146e-19 $X=0.905 $Y=2.225 $X2=0 $Y2=0
cc_105 N_A3_M1011_g N_A_196_403#_c_434_n 0.00110864f $X=0.905 $Y=2.225 $X2=0
+ $Y2=0
cc_106 N_A3_c_78_n N_VGND_c_457_n 0.00315951f $X=1.025 $Y=0.77 $X2=0 $Y2=0
cc_107 N_A3_c_79_n N_VGND_c_457_n 0.00225996f $X=1.025 $Y=0.845 $X2=0 $Y2=0
cc_108 A3 N_VGND_c_457_n 0.011009f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_109 N_A3_c_81_n N_VGND_c_457_n 6.6595e-19 $X=0.825 $Y=1.325 $X2=0 $Y2=0
cc_110 N_A3_c_78_n N_VGND_c_459_n 0.0058025f $X=1.025 $Y=0.77 $X2=0 $Y2=0
cc_111 N_A3_c_79_n N_VGND_c_459_n 2.90496e-19 $X=1.025 $Y=0.845 $X2=0 $Y2=0
cc_112 N_A3_c_78_n N_VGND_c_463_n 0.0105767f $X=1.025 $Y=0.77 $X2=0 $Y2=0
cc_113 N_A3_c_79_n N_VGND_c_463_n 3.88736e-19 $X=1.025 $Y=0.845 $X2=0 $Y2=0
cc_114 A3 N_VGND_c_463_n 0.00142707f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_115 N_A2_M1003_g N_A_54_154#_c_179_n 0.00564446f $X=1.335 $Y=2.225 $X2=0
+ $Y2=0
cc_116 A2 N_A_54_154#_c_174_n 0.00913939f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_117 N_A2_M1003_g N_A1_M1010_g 0.0168423f $X=1.335 $Y=2.225 $X2=0 $Y2=0
cc_118 N_A2_M1008_g N_A1_c_266_n 0.0502935f $X=1.385 $Y=0.45 $X2=0 $Y2=0
cc_119 A2 N_A1_c_266_n 0.00525206f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_120 N_A2_c_125_n A1 5.82e-19 $X=1.365 $Y=1.665 $X2=0 $Y2=0
cc_121 A2 A1 0.0112078f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_122 N_A2_c_125_n N_A1_c_269_n 0.021561f $X=1.365 $Y=1.665 $X2=0 $Y2=0
cc_123 A2 N_A1_c_269_n 2.10958e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_124 N_A2_M1008_g N_A1_c_270_n 0.00977375f $X=1.385 $Y=0.45 $X2=0 $Y2=0
cc_125 A2 N_A1_c_270_n 0.00582135f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_126 N_A2_c_127_n N_A1_c_270_n 0.021561f $X=1.365 $Y=1.325 $X2=0 $Y2=0
cc_127 A2 N_B1_c_316_n 0.013009f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A2_M1003_g N_VPWR_c_398_n 0.0030878f $X=1.335 $Y=2.225 $X2=0 $Y2=0
cc_129 N_A2_M1003_g N_VPWR_c_396_n 8.50146e-19 $X=1.335 $Y=2.225 $X2=0 $Y2=0
cc_130 N_A2_M1003_g N_A_196_403#_c_433_n 0.0137304f $X=1.335 $Y=2.225 $X2=0
+ $Y2=0
cc_131 N_A2_c_130_n N_A_196_403#_c_433_n 0.00442432f $X=1.365 $Y=1.83 $X2=0
+ $Y2=0
cc_132 A2 N_A_196_403#_c_433_n 0.0226934f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_133 N_A2_M1003_g N_A_196_403#_c_434_n 2.0918e-19 $X=1.335 $Y=2.225 $X2=0
+ $Y2=0
cc_134 N_A2_c_130_n N_A_196_403#_c_434_n 6.9342e-19 $X=1.365 $Y=1.83 $X2=0 $Y2=0
cc_135 A2 N_A_196_403#_c_434_n 0.00922358f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_136 N_A2_M1008_g N_VGND_c_459_n 0.00394727f $X=1.385 $Y=0.45 $X2=0 $Y2=0
cc_137 A2 N_VGND_c_459_n 0.00963484f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_138 N_A2_M1008_g N_VGND_c_463_n 0.00528002f $X=1.385 $Y=0.45 $X2=0 $Y2=0
cc_139 A2 N_VGND_c_463_n 0.0133553f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_140 A2 A_220_48# 0.00139886f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_141 A2 A_292_48# 0.00227604f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_142 N_A_54_154#_c_179_n N_A1_M1010_g 0.0046849f $X=1.975 $Y=3.03 $X2=0 $Y2=0
cc_143 N_A_54_154#_c_183_n N_A1_M1010_g 0.00175853f $X=2.14 $Y=2.94 $X2=0 $Y2=0
cc_144 N_A_54_154#_c_174_n N_A1_c_266_n 0.00126155f $X=2.065 $Y=0.735 $X2=0
+ $Y2=0
cc_145 N_A_54_154#_c_174_n N_A1_c_267_n 0.00367717f $X=2.065 $Y=0.735 $X2=0
+ $Y2=0
cc_146 N_A_54_154#_c_175_n A1 0.00811499f $X=2.695 $Y=2.055 $X2=0 $Y2=0
cc_147 N_A_54_154#_c_174_n N_A1_c_269_n 0.00462608f $X=2.065 $Y=0.735 $X2=0
+ $Y2=0
cc_148 N_A_54_154#_c_173_n N_B1_M1000_g 0.0118284f $X=2.61 $Y=0.735 $X2=0 $Y2=0
cc_149 N_A_54_154#_c_175_n N_B1_M1000_g 0.00199766f $X=2.695 $Y=2.055 $X2=0
+ $Y2=0
cc_150 N_A_54_154#_c_182_n N_B1_M1004_g 0.00472478f $X=2.61 $Y=2.94 $X2=0 $Y2=0
cc_151 N_A_54_154#_c_183_n N_B1_M1004_g 0.0018112f $X=2.14 $Y=2.94 $X2=0 $Y2=0
cc_152 N_A_54_154#_c_185_n N_B1_M1004_g 0.00296944f $X=2.695 $Y=2.855 $X2=0
+ $Y2=0
cc_153 N_A_54_154#_c_173_n N_B1_c_315_n 0.00502379f $X=2.61 $Y=0.735 $X2=0 $Y2=0
cc_154 N_A_54_154#_c_175_n N_B1_c_315_n 0.0167388f $X=2.695 $Y=2.055 $X2=0 $Y2=0
cc_155 N_A_54_154#_c_173_n N_B1_c_316_n 0.0242537f $X=2.61 $Y=0.735 $X2=0 $Y2=0
cc_156 N_A_54_154#_c_175_n N_B1_c_316_n 0.0267485f $X=2.695 $Y=2.055 $X2=0 $Y2=0
cc_157 N_A_54_154#_c_176_n N_C1_c_345_n 0.00898095f $X=2.93 $Y=0.65 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A_54_154#_c_175_n N_C1_M1007_g 0.0178825f $X=2.695 $Y=2.055 $X2=0 $Y2=0
cc_159 N_A_54_154#_c_185_n N_C1_M1007_g 0.0185595f $X=2.695 $Y=2.855 $X2=0 $Y2=0
cc_160 N_A_54_154#_c_186_n N_C1_M1007_g 8.30205e-19 $X=2.93 $Y=2.16 $X2=0 $Y2=0
cc_161 N_A_54_154#_c_217_p N_C1_M1007_g 0.00321945f $X=2.695 $Y=2.16 $X2=0 $Y2=0
cc_162 N_A_54_154#_c_175_n N_C1_c_346_n 0.00660707f $X=2.695 $Y=2.055 $X2=0
+ $Y2=0
cc_163 N_A_54_154#_c_175_n N_C1_c_347_n 0.00907361f $X=2.695 $Y=2.055 $X2=0
+ $Y2=0
cc_164 N_A_54_154#_c_176_n N_C1_c_347_n 0.0161269f $X=2.93 $Y=0.65 $X2=0 $Y2=0
cc_165 N_A_54_154#_c_221_p N_C1_c_347_n 0.00123818f $X=2.93 $Y=0.515 $X2=0 $Y2=0
cc_166 N_A_54_154#_c_175_n C1 0.0310775f $X=2.695 $Y=2.055 $X2=0 $Y2=0
cc_167 N_A_54_154#_c_186_n C1 0.00490673f $X=2.93 $Y=2.16 $X2=0 $Y2=0
cc_168 N_A_54_154#_c_176_n C1 0.0011078f $X=2.93 $Y=0.65 $X2=0 $Y2=0
cc_169 N_A_54_154#_c_175_n N_C1_c_349_n 0.00737186f $X=2.695 $Y=2.055 $X2=0
+ $Y2=0
cc_170 N_A_54_154#_c_186_n N_C1_c_349_n 0.00602517f $X=2.93 $Y=2.16 $X2=0 $Y2=0
cc_171 N_A_54_154#_c_176_n N_C1_c_349_n 7.09129e-19 $X=2.93 $Y=0.65 $X2=0 $Y2=0
cc_172 N_A_54_154#_c_170_n N_X_c_377_n 0.0281896f $X=0.345 $Y=1.73 $X2=0 $Y2=0
cc_173 N_A_54_154#_M1002_g N_X_c_377_n 0.0249129f $X=0.475 $Y=2.225 $X2=0 $Y2=0
cc_174 N_A_54_154#_c_171_n N_X_c_377_n 0.00447135f $X=0.555 $Y=0.77 $X2=0 $Y2=0
cc_175 N_A_54_154#_c_172_n N_X_c_377_n 0.00990536f $X=0.555 $Y=0.845 $X2=0 $Y2=0
cc_176 N_A_54_154#_c_181_n N_X_c_377_n 0.0101502f $X=0.475 $Y=1.805 $X2=0 $Y2=0
cc_177 N_A_54_154#_M1002_g N_VPWR_c_397_n 0.0111879f $X=0.475 $Y=2.225 $X2=0
+ $Y2=0
cc_178 N_A_54_154#_c_179_n N_VPWR_c_397_n 0.0206468f $X=1.975 $Y=3.03 $X2=0
+ $Y2=0
cc_179 N_A_54_154#_c_179_n N_VPWR_c_398_n 0.0273571f $X=1.975 $Y=3.03 $X2=0
+ $Y2=0
cc_180 N_A_54_154#_c_182_n N_VPWR_c_398_n 0.0132149f $X=2.61 $Y=2.94 $X2=0 $Y2=0
cc_181 N_A_54_154#_c_183_n N_VPWR_c_398_n 0.00396537f $X=2.14 $Y=2.94 $X2=0
+ $Y2=0
cc_182 N_A_54_154#_c_180_n N_VPWR_c_399_n 0.00602857f $X=0.55 $Y=3.03 $X2=0
+ $Y2=0
cc_183 N_A_54_154#_c_179_n N_VPWR_c_401_n 0.0191142f $X=1.975 $Y=3.03 $X2=0
+ $Y2=0
cc_184 N_A_54_154#_c_179_n N_VPWR_c_402_n 0.0110537f $X=1.975 $Y=3.03 $X2=0
+ $Y2=0
cc_185 N_A_54_154#_c_182_n N_VPWR_c_402_n 0.039478f $X=2.61 $Y=2.94 $X2=0 $Y2=0
cc_186 N_A_54_154#_c_179_n N_VPWR_c_396_n 0.0400575f $X=1.975 $Y=3.03 $X2=0
+ $Y2=0
cc_187 N_A_54_154#_c_180_n N_VPWR_c_396_n 0.00849474f $X=0.55 $Y=3.03 $X2=0
+ $Y2=0
cc_188 N_A_54_154#_c_182_n N_VPWR_c_396_n 0.0280314f $X=2.61 $Y=2.94 $X2=0 $Y2=0
cc_189 N_A_54_154#_c_183_n N_VPWR_c_396_n 0.00783059f $X=2.14 $Y=2.94 $X2=0
+ $Y2=0
cc_190 N_A_54_154#_c_179_n N_A_196_403#_c_434_n 0.00436104f $X=1.975 $Y=3.03
+ $X2=0 $Y2=0
cc_191 N_A_54_154#_c_182_n N_A_196_403#_c_435_n 0.00572775f $X=2.61 $Y=2.94
+ $X2=0 $Y2=0
cc_192 N_A_54_154#_c_183_n N_A_196_403#_c_435_n 0.00386482f $X=2.14 $Y=2.94
+ $X2=0 $Y2=0
cc_193 N_A_54_154#_c_175_n N_A_196_403#_c_435_n 0.00377628f $X=2.695 $Y=2.055
+ $X2=0 $Y2=0
cc_194 N_A_54_154#_c_173_n N_VGND_M1000_d 0.00295582f $X=2.61 $Y=0.735 $X2=0
+ $Y2=0
cc_195 N_A_54_154#_c_171_n N_VGND_c_457_n 0.0119807f $X=0.555 $Y=0.77 $X2=0
+ $Y2=0
cc_196 N_A_54_154#_c_173_n N_VGND_c_458_n 0.0196725f $X=2.61 $Y=0.735 $X2=0
+ $Y2=0
cc_197 N_A_54_154#_c_253_p N_VGND_c_459_n 0.00798902f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_198 N_A_54_154#_c_173_n N_VGND_c_459_n 0.00260089f $X=2.61 $Y=0.735 $X2=0
+ $Y2=0
cc_199 N_A_54_154#_c_171_n N_VGND_c_461_n 0.0048178f $X=0.555 $Y=0.77 $X2=0
+ $Y2=0
cc_200 N_A_54_154#_c_172_n N_VGND_c_461_n 0.0012309f $X=0.555 $Y=0.845 $X2=0
+ $Y2=0
cc_201 N_A_54_154#_c_173_n N_VGND_c_462_n 0.00337753f $X=2.61 $Y=0.735 $X2=0
+ $Y2=0
cc_202 N_A_54_154#_c_221_p N_VGND_c_462_n 0.00816281f $X=2.93 $Y=0.515 $X2=0
+ $Y2=0
cc_203 N_A_54_154#_M1009_d N_VGND_c_463_n 0.0028698f $X=1.82 $Y=0.24 $X2=0 $Y2=0
cc_204 N_A_54_154#_M1005_d N_VGND_c_463_n 0.00257886f $X=2.79 $Y=0.24 $X2=0
+ $Y2=0
cc_205 N_A_54_154#_c_171_n N_VGND_c_463_n 0.00936814f $X=0.555 $Y=0.77 $X2=0
+ $Y2=0
cc_206 N_A_54_154#_c_172_n N_VGND_c_463_n 0.0011887f $X=0.555 $Y=0.845 $X2=0
+ $Y2=0
cc_207 N_A_54_154#_c_253_p N_VGND_c_463_n 0.00758842f $X=1.96 $Y=0.515 $X2=0
+ $Y2=0
cc_208 N_A_54_154#_c_173_n N_VGND_c_463_n 0.012232f $X=2.61 $Y=0.735 $X2=0 $Y2=0
cc_209 N_A_54_154#_c_221_p N_VGND_c_463_n 0.00748321f $X=2.93 $Y=0.515 $X2=0
+ $Y2=0
cc_210 N_A1_c_266_n N_B1_M1000_g 0.0146045f $X=1.78 $Y=0.77 $X2=0 $Y2=0
cc_211 N_A1_c_267_n N_B1_M1000_g 0.0152635f $X=1.78 $Y=0.92 $X2=0 $Y2=0
cc_212 N_A1_M1010_g N_B1_M1004_g 0.0171299f $X=1.925 $Y=2.225 $X2=0 $Y2=0
cc_213 A1 N_B1_M1004_g 0.00179839f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_214 N_A1_c_269_n N_B1_M1004_g 0.0206638f $X=1.905 $Y=1.665 $X2=0 $Y2=0
cc_215 N_A1_c_270_n N_B1_M1004_g 0.00755018f $X=1.905 $Y=1.5 $X2=0 $Y2=0
cc_216 A1 N_B1_c_315_n 7.36876e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_217 N_A1_c_270_n N_B1_c_315_n 0.0152635f $X=1.905 $Y=1.5 $X2=0 $Y2=0
cc_218 A1 N_B1_c_316_n 0.0121107f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A1_c_270_n N_B1_c_316_n 0.00372892f $X=1.905 $Y=1.5 $X2=0 $Y2=0
cc_220 N_A1_M1010_g N_VPWR_c_398_n 0.00471632f $X=1.925 $Y=2.225 $X2=0 $Y2=0
cc_221 N_A1_M1010_g N_VPWR_c_396_n 7.05681e-19 $X=1.925 $Y=2.225 $X2=0 $Y2=0
cc_222 N_A1_M1010_g N_A_196_403#_c_433_n 0.0132278f $X=1.925 $Y=2.225 $X2=0
+ $Y2=0
cc_223 A1 N_A_196_403#_c_433_n 0.0196456f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A1_c_269_n N_A_196_403#_c_433_n 0.00401873f $X=1.905 $Y=1.665 $X2=0
+ $Y2=0
cc_225 N_A1_M1010_g N_A_196_403#_c_435_n 2.0918e-19 $X=1.925 $Y=2.225 $X2=0
+ $Y2=0
cc_226 A1 N_A_196_403#_c_435_n 0.0160093f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_227 N_A1_c_269_n N_A_196_403#_c_435_n 8.52657e-19 $X=1.905 $Y=1.665 $X2=0
+ $Y2=0
cc_228 N_A1_c_266_n N_VGND_c_458_n 0.00146653f $X=1.78 $Y=0.77 $X2=0 $Y2=0
cc_229 N_A1_c_266_n N_VGND_c_459_n 0.0058025f $X=1.78 $Y=0.77 $X2=0 $Y2=0
cc_230 N_A1_c_267_n N_VGND_c_459_n 7.78467e-19 $X=1.78 $Y=0.92 $X2=0 $Y2=0
cc_231 N_A1_c_266_n N_VGND_c_463_n 0.0107903f $X=1.78 $Y=0.77 $X2=0 $Y2=0
cc_232 N_A1_c_267_n N_VGND_c_463_n 9.45133e-19 $X=1.78 $Y=0.92 $X2=0 $Y2=0
cc_233 N_B1_M1000_g N_C1_c_345_n 0.0180068f $X=2.175 $Y=0.45 $X2=-0.19
+ $Y2=-0.245
cc_234 N_B1_c_315_n N_C1_c_346_n 0.00322754f $X=2.265 $Y=1.095 $X2=0 $Y2=0
cc_235 N_B1_M1004_g N_C1_c_349_n 0.0660463f $X=2.355 $Y=2.225 $X2=0 $Y2=0
cc_236 N_B1_M1004_g N_A_196_403#_c_435_n 8.74262e-19 $X=2.355 $Y=2.225 $X2=0
+ $Y2=0
cc_237 N_B1_M1000_g N_VGND_c_458_n 0.00722433f $X=2.175 $Y=0.45 $X2=0 $Y2=0
cc_238 N_B1_M1000_g N_VGND_c_459_n 0.00408264f $X=2.175 $Y=0.45 $X2=0 $Y2=0
cc_239 N_B1_M1000_g N_VGND_c_463_n 0.00480387f $X=2.175 $Y=0.45 $X2=0 $Y2=0
cc_240 N_C1_M1007_g N_VPWR_c_402_n 5.2995e-19 $X=2.715 $Y=2.225 $X2=0 $Y2=0
cc_241 N_C1_M1007_g N_VPWR_c_396_n 2.81387e-19 $X=2.715 $Y=2.225 $X2=0 $Y2=0
cc_242 N_C1_c_345_n N_VGND_c_458_n 0.00718975f $X=2.715 $Y=0.77 $X2=0 $Y2=0
cc_243 N_C1_c_345_n N_VGND_c_462_n 0.0042308f $X=2.715 $Y=0.77 $X2=0 $Y2=0
cc_244 N_C1_c_347_n N_VGND_c_462_n 0.0010541f $X=3 $Y=0.845 $X2=0 $Y2=0
cc_245 N_C1_c_345_n N_VGND_c_463_n 0.00729017f $X=2.715 $Y=0.77 $X2=0 $Y2=0
cc_246 N_C1_c_347_n N_VGND_c_463_n 0.00106583f $X=3 $Y=0.845 $X2=0 $Y2=0
cc_247 N_X_c_377_n N_VPWR_c_397_n 0.0411284f $X=0.34 $Y=0.515 $X2=0 $Y2=0
cc_248 N_X_c_377_n N_VPWR_c_399_n 0.00797353f $X=0.34 $Y=0.515 $X2=0 $Y2=0
cc_249 N_X_c_377_n N_VPWR_c_396_n 0.00903473f $X=0.34 $Y=0.515 $X2=0 $Y2=0
cc_250 N_X_c_377_n N_A_196_403#_c_434_n 0.00389092f $X=0.34 $Y=0.515 $X2=0 $Y2=0
cc_251 N_X_c_377_n N_VGND_c_461_n 0.0116871f $X=0.34 $Y=0.515 $X2=0 $Y2=0
cc_252 N_X_M1001_s N_VGND_c_463_n 0.0028742f $X=0.215 $Y=0.24 $X2=0 $Y2=0
cc_253 N_X_c_377_n N_VGND_c_463_n 0.00989163f $X=0.34 $Y=0.515 $X2=0 $Y2=0
cc_254 N_VPWR_M1003_d N_A_196_403#_c_433_n 0.00392154f $X=1.41 $Y=2.015 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_398_n N_A_196_403#_c_433_n 0.0254128f $X=1.63 $Y=2.365 $X2=0
+ $Y2=0
cc_256 N_VGND_c_463_n A_220_48# 0.00251844f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_257 N_VGND_c_463_n A_292_48# 0.00669092f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
