* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
X0 VPWR a_395_398# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_782_119# CIN a_84_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A a_710_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 VGND a_84_21# SUM VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_710_419# B a_782_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_782_419# CIN a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VPWR A a_1653_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_309_131# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR B a_309_398# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_710_119# B a_782_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_84_21# a_395_398# a_940_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1653_137# B a_395_398# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR B a_941_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VGND A a_710_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_84_21# a_395_398# a_941_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 SUM a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_309_131# CIN a_395_398# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_309_398# CIN a_395_398# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_309_398# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_940_119# CIN VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_84_21# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_1653_367# B a_395_398# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_941_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 VGND B a_940_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 SUM a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VGND a_395_398# COUT VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_941_419# CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 COUT a_395_398# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 VGND B a_309_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_940_119# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VGND A a_1653_137# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 COUT a_395_398# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
