* File: sky130_fd_sc_lp__dfxbp_lp.pxi.spice
* Created: Wed Sep  2 09:45:00 2020
* 
x_PM_SKY130_FD_SC_LP__DFXBP_LP%CLK N_CLK_M1013_g N_CLK_c_221_n N_CLK_M1018_g
+ N_CLK_c_222_n N_CLK_M1006_g CLK CLK N_CLK_c_224_n
+ PM_SKY130_FD_SC_LP__DFXBP_LP%CLK
x_PM_SKY130_FD_SC_LP__DFXBP_LP%D N_D_M1028_g N_D_M1000_g N_D_c_257_n N_D_c_258_n
+ N_D_M1002_g N_D_c_260_n D N_D_c_261_n PM_SKY130_FD_SC_LP__DFXBP_LP%D
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_615_93# N_A_615_93#_M1020_d N_A_615_93#_M1031_d
+ N_A_615_93#_M1027_d N_A_615_93#_M1023_s N_A_615_93#_c_305_n
+ N_A_615_93#_M1019_g N_A_615_93#_c_306_n N_A_615_93#_c_323_n
+ N_A_615_93#_M1004_g N_A_615_93#_c_307_n N_A_615_93#_c_308_n
+ N_A_615_93#_c_309_n N_A_615_93#_c_310_n N_A_615_93#_c_324_n
+ N_A_615_93#_c_311_n N_A_615_93#_c_312_n N_A_615_93#_c_313_n
+ N_A_615_93#_c_314_n N_A_615_93#_c_315_n N_A_615_93#_c_316_n
+ N_A_615_93#_c_317_n N_A_615_93#_c_318_n N_A_615_93#_c_319_n
+ N_A_615_93#_c_327_n N_A_615_93#_c_320_n N_A_615_93#_c_329_n
+ N_A_615_93#_c_330_n N_A_615_93#_c_321_n PM_SKY130_FD_SC_LP__DFXBP_LP%A_615_93#
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_455_85# N_A_455_85#_M1016_d N_A_455_85#_M1026_d
+ N_A_455_85#_c_482_n N_A_455_85#_M1030_g N_A_455_85#_c_483_n
+ N_A_455_85#_c_484_n N_A_455_85#_c_485_n N_A_455_85#_M1020_g
+ N_A_455_85#_c_486_n N_A_455_85#_M1027_g N_A_455_85#_c_491_n
+ N_A_455_85#_c_487_n N_A_455_85#_c_493_n N_A_455_85#_c_488_n
+ PM_SKY130_FD_SC_LP__DFXBP_LP%A_455_85#
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_27_403# N_A_27_403#_M1018_s N_A_27_403#_M1013_s
+ N_A_27_403#_c_588_n N_A_27_403#_M1026_g N_A_27_403#_M1016_g
+ N_A_27_403#_c_591_n N_A_27_403#_c_573_n N_A_27_403#_M1034_g
+ N_A_27_403#_c_574_n N_A_27_403#_c_575_n N_A_27_403#_c_592_n
+ N_A_27_403#_M1033_g N_A_27_403#_c_576_n N_A_27_403#_M1009_g
+ N_A_27_403#_c_577_n N_A_27_403#_c_578_n N_A_27_403#_c_579_n
+ N_A_27_403#_c_580_n N_A_27_403#_M1023_g N_A_27_403#_M1022_g
+ N_A_27_403#_c_583_n N_A_27_403#_c_584_n N_A_27_403#_c_585_n
+ N_A_27_403#_c_586_n N_A_27_403#_c_587_n N_A_27_403#_c_599_n
+ N_A_27_403#_c_600_n N_A_27_403#_c_601_n N_A_27_403#_c_613_n
+ N_A_27_403#_c_614_n N_A_27_403#_c_602_n N_A_27_403#_c_603_n
+ N_A_27_403#_c_604_n N_A_27_403#_c_605_n PM_SKY130_FD_SC_LP__DFXBP_LP%A_27_403#
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_511_218# N_A_511_218#_M1034_s
+ N_A_511_218#_M1033_s N_A_511_218#_M1008_g N_A_511_218#_M1029_g
+ N_A_511_218#_c_748_n N_A_511_218#_c_749_n N_A_511_218#_M1005_g
+ N_A_511_218#_M1031_g N_A_511_218#_c_751_n N_A_511_218#_c_752_n
+ N_A_511_218#_c_753_n N_A_511_218#_c_759_n N_A_511_218#_c_754_n
+ N_A_511_218#_c_755_n N_A_511_218#_c_762_n
+ PM_SKY130_FD_SC_LP__DFXBP_LP%A_511_218#
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_1507_321# N_A_1507_321#_M1015_d
+ N_A_1507_321#_M1035_d N_A_1507_321#_M1021_g N_A_1507_321#_c_867_n
+ N_A_1507_321#_c_868_n N_A_1507_321#_M1010_g N_A_1507_321#_M1007_g
+ N_A_1507_321#_M1011_g N_A_1507_321#_M1014_g N_A_1507_321#_M1017_g
+ N_A_1507_321#_M1003_g N_A_1507_321#_M1012_g N_A_1507_321#_c_875_n
+ N_A_1507_321#_c_887_n N_A_1507_321#_c_888_n N_A_1507_321#_c_889_n
+ N_A_1507_321#_c_890_n N_A_1507_321#_c_876_n N_A_1507_321#_c_877_n
+ N_A_1507_321#_c_878_n N_A_1507_321#_c_879_n N_A_1507_321#_c_880_n
+ N_A_1507_321#_c_892_n N_A_1507_321#_c_881_n N_A_1507_321#_c_964_p
+ N_A_1507_321#_c_882_n N_A_1507_321#_c_883_n
+ PM_SKY130_FD_SC_LP__DFXBP_LP%A_1507_321#
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_1339_153# N_A_1339_153#_M1022_d
+ N_A_1339_153#_M1023_d N_A_1339_153#_M1035_g N_A_1339_153#_M1024_g
+ N_A_1339_153#_c_1017_n N_A_1339_153#_M1015_g N_A_1339_153#_c_1019_n
+ N_A_1339_153#_c_1028_n N_A_1339_153#_c_1033_n N_A_1339_153#_c_1046_n
+ N_A_1339_153#_c_1020_n N_A_1339_153#_c_1021_n N_A_1339_153#_c_1022_n
+ N_A_1339_153#_c_1023_n N_A_1339_153#_c_1040_n N_A_1339_153#_c_1024_n
+ N_A_1339_153#_c_1025_n N_A_1339_153#_c_1026_n
+ PM_SKY130_FD_SC_LP__DFXBP_LP%A_1339_153#
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_2062_367# N_A_2062_367#_M1012_d
+ N_A_2062_367#_M1014_d N_A_2062_367#_M1032_g N_A_2062_367#_c_1127_n
+ N_A_2062_367#_M1001_g N_A_2062_367#_M1025_g N_A_2062_367#_c_1121_n
+ N_A_2062_367#_c_1128_n N_A_2062_367#_c_1129_n N_A_2062_367#_c_1130_n
+ N_A_2062_367#_c_1131_n N_A_2062_367#_c_1122_n N_A_2062_367#_c_1123_n
+ N_A_2062_367#_c_1124_n N_A_2062_367#_c_1125_n N_A_2062_367#_c_1126_n
+ PM_SKY130_FD_SC_LP__DFXBP_LP%A_2062_367#
x_PM_SKY130_FD_SC_LP__DFXBP_LP%VPWR N_VPWR_M1013_d N_VPWR_M1004_d N_VPWR_M1033_d
+ N_VPWR_M1021_d N_VPWR_M1007_d N_VPWR_M1001_s N_VPWR_c_1182_n N_VPWR_c_1183_n
+ N_VPWR_c_1184_n N_VPWR_c_1185_n N_VPWR_c_1186_n N_VPWR_c_1187_n
+ N_VPWR_c_1188_n N_VPWR_c_1189_n VPWR N_VPWR_c_1190_n N_VPWR_c_1191_n
+ N_VPWR_c_1192_n N_VPWR_c_1193_n N_VPWR_c_1194_n N_VPWR_c_1181_n
+ N_VPWR_c_1196_n N_VPWR_c_1197_n N_VPWR_c_1198_n N_VPWR_c_1199_n
+ N_VPWR_c_1200_n PM_SKY130_FD_SC_LP__DFXBP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_239_403# N_A_239_403#_M1002_d
+ N_A_239_403#_M1028_d N_A_239_403#_M1008_d N_A_239_403#_c_1303_n
+ N_A_239_403#_c_1301_n N_A_239_403#_c_1305_n N_A_239_403#_c_1302_n
+ N_A_239_403#_c_1343_p N_A_239_403#_c_1306_n N_A_239_403#_c_1323_n
+ PM_SKY130_FD_SC_LP__DFXBP_LP%A_239_403#
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_349_323# N_A_349_323#_M1026_s
+ N_A_349_323#_M1004_s N_A_349_323#_c_1354_n N_A_349_323#_c_1355_n
+ N_A_349_323#_c_1356_n PM_SKY130_FD_SC_LP__DFXBP_LP%A_349_323#
x_PM_SKY130_FD_SC_LP__DFXBP_LP%Q N_Q_M1011_s N_Q_M1007_s N_Q_c_1390_n Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DFXBP_LP%Q
x_PM_SKY130_FD_SC_LP__DFXBP_LP%Q_N N_Q_N_M1025_d N_Q_N_M1001_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N PM_SKY130_FD_SC_LP__DFXBP_LP%Q_N
x_PM_SKY130_FD_SC_LP__DFXBP_LP%VGND N_VGND_M1006_d N_VGND_M1019_d N_VGND_M1009_d
+ N_VGND_M1010_d N_VGND_M1017_d N_VGND_M1032_s N_VGND_c_1435_n N_VGND_c_1436_n
+ N_VGND_c_1437_n N_VGND_c_1438_n N_VGND_c_1439_n N_VGND_c_1440_n
+ N_VGND_c_1441_n N_VGND_c_1442_n N_VGND_c_1443_n N_VGND_c_1444_n VGND
+ N_VGND_c_1445_n N_VGND_c_1446_n N_VGND_c_1447_n N_VGND_c_1448_n
+ N_VGND_c_1449_n N_VGND_c_1450_n N_VGND_c_1451_n N_VGND_c_1452_n
+ N_VGND_c_1453_n N_VGND_c_1454_n PM_SKY130_FD_SC_LP__DFXBP_LP%VGND
x_PM_SKY130_FD_SC_LP__DFXBP_LP%A_1232_153# N_A_1232_153#_M1022_s
+ N_A_1232_153#_M1010_s N_A_1232_153#_c_1567_n N_A_1232_153#_c_1568_n
+ N_A_1232_153#_c_1569_n N_A_1232_153#_c_1570_n
+ PM_SKY130_FD_SC_LP__DFXBP_LP%A_1232_153#
cc_1 VNB N_CLK_M1013_g 0.0195214f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.515
cc_2 VNB N_CLK_c_221_n 0.0187083f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.955
cc_3 VNB N_CLK_c_222_n 0.0159008f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.955
cc_4 VNB CLK 0.0107521f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB N_CLK_c_224_n 0.0571711f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.12
cc_6 VNB N_D_M1000_g 0.0228302f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.635
cc_7 VNB N_D_c_257_n 0.0206923f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.635
cc_8 VNB N_D_c_258_n 0.028009f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_9 VNB N_D_M1002_g 0.0211214f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.182
cc_10 VNB N_D_c_260_n 0.00574428f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.182
cc_11 VNB N_D_c_261_n 0.0292176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_615_93#_c_305_n 0.0153544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_615_93#_c_306_n 0.0139475f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.182
cc_14 VNB N_A_615_93#_c_307_n 0.00280422f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.555
cc_15 VNB N_A_615_93#_c_308_n 0.00898161f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.12
cc_16 VNB N_A_615_93#_c_309_n 0.0215255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_615_93#_c_310_n 0.00509676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_615_93#_c_311_n 0.00477616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_615_93#_c_312_n 0.0223821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_615_93#_c_313_n 0.00138846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_615_93#_c_314_n 0.00101942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_615_93#_c_315_n 0.0052749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_615_93#_c_316_n 0.00122679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_615_93#_c_317_n 2.22702e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_615_93#_c_318_n 0.0336498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_615_93#_c_319_n 0.00784233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_615_93#_c_320_n 0.00965539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_615_93#_c_321_n 0.00950819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_455_85#_c_482_n 0.0141997f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.635
cc_30 VNB N_A_455_85#_c_483_n 0.00941408f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.635
cc_31 VNB N_A_455_85#_c_484_n 0.00793581f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_32 VNB N_A_455_85#_c_485_n 0.0156505f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_33 VNB N_A_455_85#_c_486_n 0.0446123f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.182
cc_34 VNB N_A_455_85#_c_487_n 0.0110385f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.555
cc_35 VNB N_A_455_85#_c_488_n 0.00577389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_403#_M1016_g 0.0462139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_403#_c_573_n 0.0148742f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.182
cc_38 VNB N_A_27_403#_c_574_n 0.00686244f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.182
cc_39 VNB N_A_27_403#_c_575_n 0.0104369f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.555
cc_40 VNB N_A_27_403#_c_576_n 0.012615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_403#_c_577_n 0.0118471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_403#_c_578_n 0.00639742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_403#_c_579_n 6.60698e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_403#_c_580_n 0.0237135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_403#_M1023_g 0.00160781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_403#_M1022_g 0.0314971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_403#_c_583_n 0.00488725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_403#_c_584_n 0.00967135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_403#_c_585_n 0.00549867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_403#_c_586_n 0.0104327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_27_403#_c_587_n 0.0588655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_511_218#_M1008_g 0.0113481f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.635
cc_53 VNB N_A_511_218#_M1029_g 0.026293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_511_218#_c_748_n 0.329186f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.182
cc_55 VNB N_A_511_218#_c_749_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.182
cc_56 VNB N_A_511_218#_M1031_g 0.0618253f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.925
cc_57 VNB N_A_511_218#_c_751_n 0.0173256f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.12
cc_58 VNB N_A_511_218#_c_752_n 0.00634607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_511_218#_c_753_n 0.00225453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_511_218#_c_754_n 4.28188e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_511_218#_c_755_n 0.00886599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1507_321#_c_867_n 0.0424665f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_63 VNB N_A_1507_321#_c_868_n 0.0183331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1507_321#_M1007_g 0.0050099f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.12
cc_65 VNB N_A_1507_321#_M1011_g 0.0224345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1507_321#_M1014_g 0.00645651f $X=-0.19 $Y=-0.245 $X2=0.765
+ $Y2=1.12
cc_67 VNB N_A_1507_321#_M1017_g 0.0188742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1507_321#_M1003_g 0.0196394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1507_321#_M1012_g 0.0273115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1507_321#_c_875_n 0.020799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1507_321#_c_876_n 0.00980509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1507_321#_c_877_n 0.0220665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1507_321#_c_878_n 0.00582946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1507_321#_c_879_n 0.00233324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1507_321#_c_880_n 0.0509388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1507_321#_c_881_n 0.0162418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1507_321#_c_882_n 0.107631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1507_321#_c_883_n 0.0159125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1339_153#_M1024_g 0.0342795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1339_153#_c_1017_n 0.0231569f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.182
cc_81 VNB N_A_1339_153#_M1015_g 0.0366736f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=1.12
cc_82 VNB N_A_1339_153#_c_1019_n 0.0127933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1339_153#_c_1020_n 0.00544871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1339_153#_c_1021_n 0.00239867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1339_153#_c_1022_n 0.00384581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1339_153#_c_1023_n 0.0210988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1339_153#_c_1024_n 0.00167252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1339_153#_c_1025_n 0.00377004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1339_153#_c_1026_n 0.0255952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2062_367#_M1032_g 0.0420972f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.635
cc_91 VNB N_A_2062_367#_M1025_g 0.0431575f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.182
cc_92 VNB N_A_2062_367#_c_1121_n 0.0209288f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=1.182
cc_93 VNB N_A_2062_367#_c_1122_n 0.0226938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2062_367#_c_1123_n 0.00123036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2062_367#_c_1124_n 0.0278279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2062_367#_c_1125_n 0.0101689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2062_367#_c_1126_n 0.00474079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VPWR_c_1181_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_239_403#_c_1301_n 0.00642025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_239_403#_c_1302_n 0.00559202f $X=-0.19 $Y=-0.245 $X2=0.765
+ $Y2=0.555
cc_101 VNB N_Q_c_1390_n 0.0170062f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.955
cc_102 VNB Q 0.00849022f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_103 VNB Q_N 0.0613638f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.635
cc_104 VNB N_VGND_c_1435_n 0.0129758f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=0.555
cc_105 VNB N_VGND_c_1436_n 0.0095342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1437_n 0.0160629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1438_n 0.00612745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1439_n 0.0219093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1440_n 0.0192162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1441_n 0.0508155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1442_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1443_n 0.0461432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1444_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1445_n 0.0331586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1446_n 0.0553875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1447_n 0.0574961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1448_n 0.0305572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1449_n 0.0271986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1450_n 0.697454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1451_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1452_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1453_n 0.00397464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1454_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_1232_153#_c_1567_n 0.0171898f $X=-0.19 $Y=-0.245 $X2=0.91
+ $Y2=0.635
cc_125 VNB N_A_1232_153#_c_1568_n 0.0347201f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=0.47
cc_126 VNB N_A_1232_153#_c_1569_n 0.00451329f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=0.84
cc_127 VNB N_A_1232_153#_c_1570_n 0.0102503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VPB N_CLK_M1013_g 0.0453251f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.515
cc_129 VPB N_D_M1028_g 0.0303689f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.515
cc_130 VPB N_D_c_261_n 0.0284041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_615_93#_c_306_n 0.0138935f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.182
cc_132 VPB N_A_615_93#_c_323_n 0.0202448f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=1.12
cc_133 VPB N_A_615_93#_c_324_n 0.0228225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_615_93#_c_317_n 0.00170437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_615_93#_c_318_n 0.017098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_615_93#_c_327_n 0.00569126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_615_93#_c_320_n 0.00402704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_615_93#_c_329_n 0.0108438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_615_93#_c_330_n 0.00982852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_455_85#_c_486_n 0.00375913f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.182
cc_141 VPB N_A_455_85#_M1027_g 0.0253231f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=1.182
cc_142 VPB N_A_455_85#_c_491_n 0.00199261f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=1.12
cc_143 VPB N_A_455_85#_c_487_n 0.0011796f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=0.555
cc_144 VPB N_A_455_85#_c_493_n 0.00658077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_455_85#_c_488_n 0.0010645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_27_403#_c_588_n 0.0125411f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.635
cc_147 VPB N_A_27_403#_M1026_g 0.0161773f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.635
cc_148 VPB N_A_27_403#_M1016_g 0.00309979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_27_403#_c_591_n 0.274605f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.182
cc_150 VPB N_A_27_403#_c_592_n 0.0217439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_27_403#_c_578_n 0.00712374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_27_403#_c_579_n 0.0776591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_27_403#_M1023_g 0.0439505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_27_403#_c_583_n 0.00648663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_27_403#_c_585_n 0.00117007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_27_403#_c_587_n 0.0140924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_27_403#_c_599_n 0.0100351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_27_403#_c_600_n 0.00636976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_27_403#_c_601_n 0.0191977f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_27_403#_c_602_n 9.25161e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_27_403#_c_603_n 0.0266003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_27_403#_c_604_n 0.0518933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_27_403#_c_605_n 0.00708086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_511_218#_M1008_g 0.0269865f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.635
cc_165 VPB N_A_511_218#_M1005_g 0.0262401f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=1.12
cc_166 VPB N_A_511_218#_c_752_n 0.00390377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_511_218#_c_759_n 0.00446262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_511_218#_c_754_n 0.00119673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_511_218#_c_755_n 0.0217388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_511_218#_c_762_n 0.0206444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_1507_321#_M1021_g 0.0277645f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.635
cc_172 VPB N_A_1507_321#_M1007_g 0.0288665f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=1.12
cc_173 VPB N_A_1507_321#_M1014_g 0.033421f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=1.12
cc_174 VPB N_A_1507_321#_c_887_n 0.00142027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_1507_321#_c_888_n 0.00374712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_1507_321#_c_889_n 4.43442e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_1507_321#_c_890_n 0.0158167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_1507_321#_c_876_n 0.00786757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_1507_321#_c_892_n 0.00610304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_1507_321#_c_883_n 0.035789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_1339_153#_M1035_g 0.0382689f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.635
cc_182 VPB N_A_1339_153#_c_1028_n 0.0162107f $X=-0.19 $Y=1.655 $X2=0.765
+ $Y2=0.925
cc_183 VPB N_A_1339_153#_c_1022_n 0.00328096f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1339_153#_c_1025_n 7.54819e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1339_153#_c_1026_n 9.44314e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_2062_367#_c_1127_n 0.0235865f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=0.47
cc_187 VPB N_A_2062_367#_c_1128_n 0.0463594f $X=-0.19 $Y=1.655 $X2=0.765
+ $Y2=0.555
cc_188 VPB N_A_2062_367#_c_1129_n 0.0381773f $X=-0.19 $Y=1.655 $X2=0.765
+ $Y2=0.925
cc_189 VPB N_A_2062_367#_c_1130_n 0.0727349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_2062_367#_c_1131_n 0.00231174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_2062_367#_c_1124_n 0.00147005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1182_n 0.00254872f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1183_n 0.0161419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1184_n 0.0153497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1185_n 0.00562899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1186_n 0.0168231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1187_n 0.0408336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1188_n 0.058394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1189_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1190_n 0.0737311f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1191_n 0.0371316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1192_n 0.055686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1193_n 0.0454798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1194_n 0.0189248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1181_n 0.141292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1196_n 0.0237416f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1197_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1198_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1199_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1200_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_239_403#_c_1303_n 0.0135214f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.635
cc_212 VPB N_A_239_403#_c_1301_n 0.00429127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_239_403#_c_1305_n 0.00175011f $X=-0.19 $Y=1.655 $X2=0.765
+ $Y2=1.12
cc_214 VPB N_A_239_403#_c_1306_n 0.00262251f $X=-0.19 $Y=1.655 $X2=0.765
+ $Y2=1.12
cc_215 VPB N_A_349_323#_c_1354_n 0.0132081f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.635
cc_216 VPB N_A_349_323#_c_1355_n 0.00520258f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=0.47
cc_217 VPB N_A_349_323#_c_1356_n 0.00291659f $X=-0.19 $Y=1.655 $X2=0.55
+ $Y2=1.182
cc_218 VPB Q 0.0143264f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_219 VPB Q_N 0.0591357f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.635
cc_220 N_CLK_c_222_n N_D_M1000_g 0.0135624f $X=0.91 $Y=0.955 $X2=0 $Y2=0
cc_221 CLK N_D_M1000_g 0.00251655f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_222 N_CLK_c_224_n N_D_c_257_n 0.0056311f $X=0.765 $Y=1.12 $X2=0 $Y2=0
cc_223 N_CLK_c_224_n N_D_c_260_n 0.0135624f $X=0.765 $Y=1.12 $X2=0 $Y2=0
cc_224 N_CLK_M1013_g D 0.00127209f $X=0.54 $Y=2.515 $X2=0 $Y2=0
cc_225 N_CLK_M1013_g N_D_c_261_n 0.0601604f $X=0.54 $Y=2.515 $X2=0 $Y2=0
cc_226 N_CLK_c_224_n N_D_c_261_n 0.00296184f $X=0.765 $Y=1.12 $X2=0 $Y2=0
cc_227 N_CLK_M1013_g N_A_27_403#_c_587_n 0.0255218f $X=0.54 $Y=2.515 $X2=0 $Y2=0
cc_228 N_CLK_c_221_n N_A_27_403#_c_587_n 0.013307f $X=0.55 $Y=0.955 $X2=0 $Y2=0
cc_229 CLK N_A_27_403#_c_587_n 0.047627f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_230 N_CLK_c_224_n N_A_27_403#_c_587_n 0.00785944f $X=0.765 $Y=1.12 $X2=0
+ $Y2=0
cc_231 N_CLK_M1013_g N_A_27_403#_c_599_n 0.00533154f $X=0.54 $Y=2.515 $X2=0
+ $Y2=0
cc_232 N_CLK_M1013_g N_A_27_403#_c_600_n 0.00471673f $X=0.54 $Y=2.515 $X2=0
+ $Y2=0
cc_233 N_CLK_M1013_g N_A_27_403#_c_601_n 0.00853882f $X=0.54 $Y=2.515 $X2=0
+ $Y2=0
cc_234 N_CLK_M1013_g N_A_27_403#_c_613_n 0.0207463f $X=0.54 $Y=2.515 $X2=0 $Y2=0
cc_235 N_CLK_M1013_g N_A_27_403#_c_614_n 5.82128e-19 $X=0.54 $Y=2.515 $X2=0
+ $Y2=0
cc_236 N_CLK_M1013_g N_A_27_403#_c_605_n 3.84191e-19 $X=0.54 $Y=2.515 $X2=0
+ $Y2=0
cc_237 N_CLK_M1013_g N_VPWR_c_1182_n 0.0104977f $X=0.54 $Y=2.515 $X2=0 $Y2=0
cc_238 N_CLK_M1013_g N_VPWR_c_1181_n 0.00736586f $X=0.54 $Y=2.515 $X2=0 $Y2=0
cc_239 N_CLK_M1013_g N_VPWR_c_1196_n 0.00552944f $X=0.54 $Y=2.515 $X2=0 $Y2=0
cc_240 N_CLK_M1013_g N_A_239_403#_c_1305_n 8.88977e-19 $X=0.54 $Y=2.515 $X2=0
+ $Y2=0
cc_241 CLK A_125_85# 0.00133334f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_242 N_CLK_c_222_n N_VGND_c_1435_n 0.00659136f $X=0.91 $Y=0.955 $X2=0 $Y2=0
cc_243 CLK N_VGND_c_1435_n 0.0309325f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_244 N_CLK_c_221_n N_VGND_c_1445_n 0.00514647f $X=0.55 $Y=0.955 $X2=0 $Y2=0
cc_245 N_CLK_c_222_n N_VGND_c_1445_n 0.0044666f $X=0.91 $Y=0.955 $X2=0 $Y2=0
cc_246 CLK N_VGND_c_1445_n 0.00851294f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_247 N_CLK_c_221_n N_VGND_c_1450_n 0.00528353f $X=0.55 $Y=0.955 $X2=0 $Y2=0
cc_248 N_CLK_c_222_n N_VGND_c_1450_n 0.00528353f $X=0.91 $Y=0.955 $X2=0 $Y2=0
cc_249 CLK N_VGND_c_1450_n 0.011321f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_250 N_D_c_257_n N_A_27_403#_c_588_n 0.00288482f $X=1.41 $Y=1.525 $X2=0 $Y2=0
cc_251 N_D_c_261_n N_A_27_403#_M1026_g 0.00288482f $X=1.41 $Y=1.69 $X2=0 $Y2=0
cc_252 N_D_c_257_n N_A_27_403#_M1016_g 0.0025047f $X=1.41 $Y=1.525 $X2=0 $Y2=0
cc_253 N_D_M1002_g N_A_27_403#_M1016_g 0.0240898f $X=1.77 $Y=0.635 $X2=0 $Y2=0
cc_254 D N_A_27_403#_c_587_n 0.0091317f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_255 N_D_c_261_n N_A_27_403#_c_587_n 0.00156172f $X=1.41 $Y=1.69 $X2=0 $Y2=0
cc_256 N_D_M1028_g N_A_27_403#_c_600_n 0.00184553f $X=1.07 $Y=2.515 $X2=0 $Y2=0
cc_257 N_D_M1028_g N_A_27_403#_c_601_n 6.30887e-19 $X=1.07 $Y=2.515 $X2=0 $Y2=0
cc_258 N_D_M1028_g N_A_27_403#_c_613_n 0.0206468f $X=1.07 $Y=2.515 $X2=0 $Y2=0
cc_259 D N_A_27_403#_c_613_n 0.00492371f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_260 N_D_M1028_g N_A_27_403#_c_614_n 0.00664428f $X=1.07 $Y=2.515 $X2=0 $Y2=0
cc_261 N_D_M1028_g N_A_27_403#_c_602_n 0.0127412f $X=1.07 $Y=2.515 $X2=0 $Y2=0
cc_262 N_D_M1028_g N_VPWR_c_1182_n 0.00943405f $X=1.07 $Y=2.515 $X2=0 $Y2=0
cc_263 N_D_M1028_g N_VPWR_c_1190_n 0.00542131f $X=1.07 $Y=2.515 $X2=0 $Y2=0
cc_264 N_D_M1028_g N_VPWR_c_1181_n 0.00743427f $X=1.07 $Y=2.515 $X2=0 $Y2=0
cc_265 N_D_M1028_g N_A_239_403#_c_1301_n 0.00382241f $X=1.07 $Y=2.515 $X2=0
+ $Y2=0
cc_266 N_D_c_257_n N_A_239_403#_c_1301_n 0.00876579f $X=1.41 $Y=1.525 $X2=0
+ $Y2=0
cc_267 N_D_c_258_n N_A_239_403#_c_1301_n 0.00828213f $X=1.695 $Y=1.17 $X2=0
+ $Y2=0
cc_268 N_D_M1002_g N_A_239_403#_c_1301_n 0.00533548f $X=1.77 $Y=0.635 $X2=0
+ $Y2=0
cc_269 D N_A_239_403#_c_1301_n 0.0105259f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_270 N_D_M1028_g N_A_239_403#_c_1305_n 0.00518274f $X=1.07 $Y=2.515 $X2=0
+ $Y2=0
cc_271 D N_A_239_403#_c_1305_n 0.0082628f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_272 N_D_c_261_n N_A_239_403#_c_1305_n 0.00959902f $X=1.41 $Y=1.69 $X2=0 $Y2=0
cc_273 N_D_M1000_g N_A_239_403#_c_1302_n 0.00240956f $X=1.41 $Y=0.635 $X2=0
+ $Y2=0
cc_274 N_D_M1002_g N_A_239_403#_c_1302_n 0.00841438f $X=1.77 $Y=0.635 $X2=0
+ $Y2=0
cc_275 N_D_M1028_g N_A_349_323#_c_1356_n 0.00201586f $X=1.07 $Y=2.515 $X2=0
+ $Y2=0
cc_276 N_D_M1000_g N_VGND_c_1435_n 0.0128494f $X=1.41 $Y=0.635 $X2=0 $Y2=0
cc_277 N_D_M1002_g N_VGND_c_1435_n 0.00180891f $X=1.77 $Y=0.635 $X2=0 $Y2=0
cc_278 D N_VGND_c_1435_n 0.00614893f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_279 N_D_c_261_n N_VGND_c_1435_n 0.00411025f $X=1.41 $Y=1.69 $X2=0 $Y2=0
cc_280 N_D_M1000_g N_VGND_c_1446_n 0.00447026f $X=1.41 $Y=0.635 $X2=0 $Y2=0
cc_281 N_D_M1002_g N_VGND_c_1446_n 0.00514022f $X=1.77 $Y=0.635 $X2=0 $Y2=0
cc_282 N_D_M1000_g N_VGND_c_1450_n 0.00443817f $X=1.41 $Y=0.635 $X2=0 $Y2=0
cc_283 N_D_M1002_g N_VGND_c_1450_n 0.00528353f $X=1.77 $Y=0.635 $X2=0 $Y2=0
cc_284 N_A_615_93#_c_305_n N_A_455_85#_c_482_n 0.0155121f $X=3.15 $Y=1.125 $X2=0
+ $Y2=0
cc_285 N_A_615_93#_c_307_n N_A_455_85#_c_482_n 0.0117984f $X=4.15 $Y=1.05 $X2=0
+ $Y2=0
cc_286 N_A_615_93#_c_308_n N_A_455_85#_c_482_n 0.00181251f $X=4.315 $Y=0.805
+ $X2=0 $Y2=0
cc_287 N_A_615_93#_c_307_n N_A_455_85#_c_483_n 0.0041604f $X=4.15 $Y=1.05 $X2=0
+ $Y2=0
cc_288 N_A_615_93#_c_306_n N_A_455_85#_c_484_n 0.0138198f $X=3.64 $Y=1.585 $X2=0
+ $Y2=0
cc_289 N_A_615_93#_c_307_n N_A_455_85#_c_484_n 0.00258976f $X=4.15 $Y=1.05 $X2=0
+ $Y2=0
cc_290 N_A_615_93#_c_317_n N_A_455_85#_c_484_n 0.00102573f $X=3.24 $Y=1.05 $X2=0
+ $Y2=0
cc_291 N_A_615_93#_c_318_n N_A_455_85#_c_484_n 0.00820192f $X=3.24 $Y=1.29 $X2=0
+ $Y2=0
cc_292 N_A_615_93#_c_307_n N_A_455_85#_c_485_n 0.0083367f $X=4.15 $Y=1.05 $X2=0
+ $Y2=0
cc_293 N_A_615_93#_c_308_n N_A_455_85#_c_485_n 0.0118049f $X=4.315 $Y=0.805
+ $X2=0 $Y2=0
cc_294 N_A_615_93#_c_319_n N_A_455_85#_c_485_n 0.00320228f $X=4.695 $Y=1.05
+ $X2=0 $Y2=0
cc_295 N_A_615_93#_c_306_n N_A_455_85#_c_486_n 0.00425629f $X=3.64 $Y=1.585
+ $X2=0 $Y2=0
cc_296 N_A_615_93#_c_307_n N_A_455_85#_c_486_n 0.00168365f $X=4.15 $Y=1.05 $X2=0
+ $Y2=0
cc_297 N_A_615_93#_c_308_n N_A_455_85#_c_486_n 0.00129294f $X=4.315 $Y=0.805
+ $X2=0 $Y2=0
cc_298 N_A_615_93#_c_317_n N_A_455_85#_c_486_n 3.72382e-19 $X=3.24 $Y=1.05 $X2=0
+ $Y2=0
cc_299 N_A_615_93#_c_318_n N_A_455_85#_c_486_n 0.00315749f $X=3.24 $Y=1.29 $X2=0
+ $Y2=0
cc_300 N_A_615_93#_c_319_n N_A_455_85#_c_486_n 0.00899608f $X=4.695 $Y=1.05
+ $X2=0 $Y2=0
cc_301 N_A_615_93#_c_320_n N_A_455_85#_c_486_n 0.00710296f $X=4.587 $Y=1.755
+ $X2=0 $Y2=0
cc_302 N_A_615_93#_c_306_n N_A_455_85#_M1027_g 0.0260472f $X=3.64 $Y=1.585 $X2=0
+ $Y2=0
cc_303 N_A_615_93#_c_324_n N_A_455_85#_M1027_g 5.06259e-19 $X=6.14 $Y=2.2 $X2=0
+ $Y2=0
cc_304 N_A_615_93#_c_327_n N_A_455_85#_M1027_g 0.0134315f $X=4.56 $Y=1.92 $X2=0
+ $Y2=0
cc_305 N_A_615_93#_c_320_n N_A_455_85#_M1027_g 0.00375381f $X=4.587 $Y=1.755
+ $X2=0 $Y2=0
cc_306 N_A_615_93#_c_329_n N_A_455_85#_M1027_g 0.0109119f $X=4.587 $Y=2.2 $X2=0
+ $Y2=0
cc_307 N_A_615_93#_c_318_n N_A_455_85#_c_491_n 2.11318e-19 $X=3.24 $Y=1.29 $X2=0
+ $Y2=0
cc_308 N_A_615_93#_c_305_n N_A_455_85#_c_487_n 0.00103319f $X=3.15 $Y=1.125
+ $X2=0 $Y2=0
cc_309 N_A_615_93#_c_317_n N_A_455_85#_c_487_n 0.0172243f $X=3.24 $Y=1.05 $X2=0
+ $Y2=0
cc_310 N_A_615_93#_c_318_n N_A_455_85#_c_487_n 6.86452e-19 $X=3.24 $Y=1.29 $X2=0
+ $Y2=0
cc_311 N_A_615_93#_c_306_n N_A_455_85#_c_493_n 0.0129719f $X=3.64 $Y=1.585 $X2=0
+ $Y2=0
cc_312 N_A_615_93#_c_323_n N_A_455_85#_c_493_n 0.0181502f $X=3.765 $Y=1.66 $X2=0
+ $Y2=0
cc_313 N_A_615_93#_c_307_n N_A_455_85#_c_493_n 0.0194765f $X=4.15 $Y=1.05 $X2=0
+ $Y2=0
cc_314 N_A_615_93#_c_317_n N_A_455_85#_c_493_n 0.0238743f $X=3.24 $Y=1.05 $X2=0
+ $Y2=0
cc_315 N_A_615_93#_c_318_n N_A_455_85#_c_493_n 0.00665667f $X=3.24 $Y=1.29 $X2=0
+ $Y2=0
cc_316 N_A_615_93#_c_306_n N_A_455_85#_c_488_n 0.00297425f $X=3.64 $Y=1.585
+ $X2=0 $Y2=0
cc_317 N_A_615_93#_c_307_n N_A_455_85#_c_488_n 0.0267025f $X=4.15 $Y=1.05 $X2=0
+ $Y2=0
cc_318 N_A_615_93#_c_317_n N_A_455_85#_c_488_n 0.00411632f $X=3.24 $Y=1.05 $X2=0
+ $Y2=0
cc_319 N_A_615_93#_c_318_n N_A_455_85#_c_488_n 0.00196137f $X=3.24 $Y=1.29 $X2=0
+ $Y2=0
cc_320 N_A_615_93#_c_327_n N_A_455_85#_c_488_n 0.00597056f $X=4.56 $Y=1.92 $X2=0
+ $Y2=0
cc_321 N_A_615_93#_c_320_n N_A_455_85#_c_488_n 0.0263315f $X=4.587 $Y=1.755
+ $X2=0 $Y2=0
cc_322 N_A_615_93#_c_323_n N_A_27_403#_c_591_n 0.017134f $X=3.765 $Y=1.66 $X2=0
+ $Y2=0
cc_323 N_A_615_93#_c_329_n N_A_27_403#_c_591_n 0.00736082f $X=4.587 $Y=2.2 $X2=0
+ $Y2=0
cc_324 N_A_615_93#_c_308_n N_A_27_403#_c_573_n 0.00428494f $X=4.315 $Y=0.805
+ $X2=0 $Y2=0
cc_325 N_A_615_93#_c_309_n N_A_27_403#_c_573_n 0.00312855f $X=5.31 $Y=0.35 $X2=0
+ $Y2=0
cc_326 N_A_615_93#_c_311_n N_A_27_403#_c_573_n 0.00579854f $X=5.395 $Y=1.335
+ $X2=0 $Y2=0
cc_327 N_A_615_93#_c_319_n N_A_27_403#_c_573_n 9.37929e-19 $X=4.695 $Y=1.05
+ $X2=0 $Y2=0
cc_328 N_A_615_93#_c_311_n N_A_27_403#_c_574_n 0.00614703f $X=5.395 $Y=1.335
+ $X2=0 $Y2=0
cc_329 N_A_615_93#_c_320_n N_A_27_403#_c_575_n 3.97175e-19 $X=4.587 $Y=1.755
+ $X2=0 $Y2=0
cc_330 N_A_615_93#_c_324_n N_A_27_403#_c_592_n 0.0242444f $X=6.14 $Y=2.2 $X2=0
+ $Y2=0
cc_331 N_A_615_93#_c_327_n N_A_27_403#_c_592_n 0.0175905f $X=4.56 $Y=1.92 $X2=0
+ $Y2=0
cc_332 N_A_615_93#_c_320_n N_A_27_403#_c_592_n 7.00449e-19 $X=4.587 $Y=1.755
+ $X2=0 $Y2=0
cc_333 N_A_615_93#_c_311_n N_A_27_403#_c_576_n 0.0111033f $X=5.395 $Y=1.335
+ $X2=0 $Y2=0
cc_334 N_A_615_93#_c_311_n N_A_27_403#_c_577_n 0.00254286f $X=5.395 $Y=1.335
+ $X2=0 $Y2=0
cc_335 N_A_615_93#_c_312_n N_A_27_403#_c_577_n 0.0107174f $X=6.57 $Y=1.42 $X2=0
+ $Y2=0
cc_336 N_A_615_93#_c_313_n N_A_27_403#_c_577_n 8.5665e-19 $X=5.48 $Y=1.42 $X2=0
+ $Y2=0
cc_337 N_A_615_93#_c_312_n N_A_27_403#_c_578_n 0.00651055f $X=6.57 $Y=1.42 $X2=0
+ $Y2=0
cc_338 N_A_615_93#_c_324_n N_A_27_403#_c_579_n 0.0167613f $X=6.14 $Y=2.2 $X2=0
+ $Y2=0
cc_339 N_A_615_93#_c_330_n N_A_27_403#_c_579_n 0.0122348f $X=6.305 $Y=2.24 $X2=0
+ $Y2=0
cc_340 N_A_615_93#_c_312_n N_A_27_403#_c_580_n 0.0127565f $X=6.57 $Y=1.42 $X2=0
+ $Y2=0
cc_341 N_A_615_93#_c_330_n N_A_27_403#_M1023_g 0.0212879f $X=6.305 $Y=2.24 $X2=0
+ $Y2=0
cc_342 N_A_615_93#_c_312_n N_A_27_403#_M1022_g 0.00764441f $X=6.57 $Y=1.42 $X2=0
+ $Y2=0
cc_343 N_A_615_93#_c_314_n N_A_27_403#_M1022_g 0.0193892f $X=6.655 $Y=1.335
+ $X2=0 $Y2=0
cc_344 N_A_615_93#_c_316_n N_A_27_403#_M1022_g 0.00581373f $X=6.74 $Y=0.7 $X2=0
+ $Y2=0
cc_345 N_A_615_93#_c_321_n N_A_27_403#_M1022_g 2.72633e-19 $X=7.435 $Y=0.7 $X2=0
+ $Y2=0
cc_346 N_A_615_93#_c_312_n N_A_27_403#_c_583_n 0.00202826f $X=6.57 $Y=1.42 $X2=0
+ $Y2=0
cc_347 N_A_615_93#_c_313_n N_A_27_403#_c_583_n 0.00442186f $X=5.48 $Y=1.42 $X2=0
+ $Y2=0
cc_348 N_A_615_93#_c_311_n N_A_27_403#_c_584_n 0.00542036f $X=5.395 $Y=1.335
+ $X2=0 $Y2=0
cc_349 N_A_615_93#_c_312_n N_A_27_403#_c_585_n 0.00503859f $X=6.57 $Y=1.42 $X2=0
+ $Y2=0
cc_350 N_A_615_93#_c_312_n N_A_27_403#_c_586_n 0.00455582f $X=6.57 $Y=1.42 $X2=0
+ $Y2=0
cc_351 N_A_615_93#_c_319_n N_A_511_218#_M1034_s 0.00150826f $X=4.695 $Y=1.05
+ $X2=-0.19 $Y2=-0.245
cc_352 N_A_615_93#_c_324_n N_A_511_218#_M1033_s 0.0121642f $X=6.14 $Y=2.2 $X2=0
+ $Y2=0
cc_353 N_A_615_93#_c_317_n N_A_511_218#_M1008_g 8.44532e-19 $X=3.24 $Y=1.05
+ $X2=0 $Y2=0
cc_354 N_A_615_93#_c_318_n N_A_511_218#_M1008_g 0.0160171f $X=3.24 $Y=1.29 $X2=0
+ $Y2=0
cc_355 N_A_615_93#_c_305_n N_A_511_218#_M1029_g 0.0230432f $X=3.15 $Y=1.125
+ $X2=0 $Y2=0
cc_356 N_A_615_93#_c_317_n N_A_511_218#_M1029_g 0.00103399f $X=3.24 $Y=1.05
+ $X2=0 $Y2=0
cc_357 N_A_615_93#_c_305_n N_A_511_218#_c_748_n 0.0104164f $X=3.15 $Y=1.125
+ $X2=0 $Y2=0
cc_358 N_A_615_93#_c_309_n N_A_511_218#_c_748_n 0.0207487f $X=5.31 $Y=0.35 $X2=0
+ $Y2=0
cc_359 N_A_615_93#_c_310_n N_A_511_218#_c_748_n 0.00770546f $X=4.48 $Y=0.35
+ $X2=0 $Y2=0
cc_360 N_A_615_93#_c_330_n N_A_511_218#_M1005_g 2.78528e-19 $X=6.305 $Y=2.24
+ $X2=0 $Y2=0
cc_361 N_A_615_93#_c_312_n N_A_511_218#_M1031_g 0.00182904f $X=6.57 $Y=1.42
+ $X2=0 $Y2=0
cc_362 N_A_615_93#_c_314_n N_A_511_218#_M1031_g 7.55274e-19 $X=6.655 $Y=1.335
+ $X2=0 $Y2=0
cc_363 N_A_615_93#_c_315_n N_A_511_218#_M1031_g 0.0101704f $X=7.27 $Y=0.7 $X2=0
+ $Y2=0
cc_364 N_A_615_93#_c_321_n N_A_511_218#_M1031_g 0.0107148f $X=7.435 $Y=0.7 $X2=0
+ $Y2=0
cc_365 N_A_615_93#_c_318_n N_A_511_218#_c_751_n 0.0230432f $X=3.24 $Y=1.29 $X2=0
+ $Y2=0
cc_366 N_A_615_93#_c_308_n N_A_511_218#_c_752_n 0.00668935f $X=4.315 $Y=0.805
+ $X2=0 $Y2=0
cc_367 N_A_615_93#_c_311_n N_A_511_218#_c_752_n 0.0369477f $X=5.395 $Y=1.335
+ $X2=0 $Y2=0
cc_368 N_A_615_93#_c_313_n N_A_511_218#_c_752_n 0.0136729f $X=5.48 $Y=1.42 $X2=0
+ $Y2=0
cc_369 N_A_615_93#_c_319_n N_A_511_218#_c_752_n 0.013376f $X=4.695 $Y=1.05 $X2=0
+ $Y2=0
cc_370 N_A_615_93#_c_320_n N_A_511_218#_c_752_n 0.0397791f $X=4.587 $Y=1.755
+ $X2=0 $Y2=0
cc_371 N_A_615_93#_c_308_n N_A_511_218#_c_753_n 0.0115757f $X=4.315 $Y=0.805
+ $X2=0 $Y2=0
cc_372 N_A_615_93#_c_309_n N_A_511_218#_c_753_n 0.0280181f $X=5.31 $Y=0.35 $X2=0
+ $Y2=0
cc_373 N_A_615_93#_c_311_n N_A_511_218#_c_753_n 0.0121632f $X=5.395 $Y=1.335
+ $X2=0 $Y2=0
cc_374 N_A_615_93#_c_319_n N_A_511_218#_c_753_n 0.00492713f $X=4.695 $Y=1.05
+ $X2=0 $Y2=0
cc_375 N_A_615_93#_c_324_n N_A_511_218#_c_759_n 0.0194288f $X=6.14 $Y=2.2 $X2=0
+ $Y2=0
cc_376 N_A_615_93#_c_320_n N_A_511_218#_c_759_n 0.0205701f $X=4.587 $Y=1.755
+ $X2=0 $Y2=0
cc_377 N_A_615_93#_c_324_n N_A_511_218#_c_762_n 0.0408052f $X=6.14 $Y=2.2 $X2=0
+ $Y2=0
cc_378 N_A_615_93#_c_312_n N_A_511_218#_c_762_n 0.0860646f $X=6.57 $Y=1.42 $X2=0
+ $Y2=0
cc_379 N_A_615_93#_c_313_n N_A_511_218#_c_762_n 0.0123662f $X=5.48 $Y=1.42 $X2=0
+ $Y2=0
cc_380 N_A_615_93#_c_330_n N_A_511_218#_c_762_n 0.0230347f $X=6.305 $Y=2.24
+ $X2=0 $Y2=0
cc_381 N_A_615_93#_c_321_n N_A_1507_321#_c_868_n 0.00165468f $X=7.435 $Y=0.7
+ $X2=0 $Y2=0
cc_382 N_A_615_93#_c_321_n N_A_1507_321#_c_875_n 0.00657075f $X=7.435 $Y=0.7
+ $X2=0 $Y2=0
cc_383 N_A_615_93#_c_321_n N_A_1507_321#_c_883_n 2.35962e-19 $X=7.435 $Y=0.7
+ $X2=0 $Y2=0
cc_384 N_A_615_93#_c_315_n N_A_1339_153#_M1022_d 0.00674507f $X=7.27 $Y=0.7
+ $X2=-0.19 $Y2=-0.245
cc_385 N_A_615_93#_c_314_n N_A_1339_153#_c_1033_n 0.0132634f $X=6.655 $Y=1.335
+ $X2=0 $Y2=0
cc_386 N_A_615_93#_c_315_n N_A_1339_153#_c_1033_n 0.0128656f $X=7.27 $Y=0.7
+ $X2=0 $Y2=0
cc_387 N_A_615_93#_M1031_d N_A_1339_153#_c_1020_n 0.00100172f $X=7.295 $Y=0.855
+ $X2=0 $Y2=0
cc_388 N_A_615_93#_c_315_n N_A_1339_153#_c_1020_n 0.00463836f $X=7.27 $Y=0.7
+ $X2=0 $Y2=0
cc_389 N_A_615_93#_c_321_n N_A_1339_153#_c_1020_n 0.00865655f $X=7.435 $Y=0.7
+ $X2=0 $Y2=0
cc_390 N_A_615_93#_c_312_n N_A_1339_153#_c_1021_n 0.00899352f $X=6.57 $Y=1.42
+ $X2=0 $Y2=0
cc_391 N_A_615_93#_c_314_n N_A_1339_153#_c_1021_n 0.00562204f $X=6.655 $Y=1.335
+ $X2=0 $Y2=0
cc_392 N_A_615_93#_c_330_n N_A_1339_153#_c_1040_n 0.0639454f $X=6.305 $Y=2.24
+ $X2=0 $Y2=0
cc_393 N_A_615_93#_M1031_d N_A_1339_153#_c_1024_n 0.00152922f $X=7.295 $Y=0.855
+ $X2=0 $Y2=0
cc_394 N_A_615_93#_c_321_n N_A_1339_153#_c_1024_n 0.0130288f $X=7.435 $Y=0.7
+ $X2=0 $Y2=0
cc_395 N_A_615_93#_c_324_n N_VPWR_M1033_d 0.00512565f $X=6.14 $Y=2.2 $X2=0 $Y2=0
cc_396 N_A_615_93#_c_323_n N_VPWR_c_1183_n 0.0210517f $X=3.765 $Y=1.66 $X2=0
+ $Y2=0
cc_397 N_A_615_93#_c_327_n N_VPWR_c_1183_n 0.0513076f $X=4.56 $Y=1.92 $X2=0
+ $Y2=0
cc_398 N_A_615_93#_c_324_n N_VPWR_c_1184_n 0.02102f $X=6.14 $Y=2.2 $X2=0 $Y2=0
cc_399 N_A_615_93#_c_330_n N_VPWR_c_1184_n 0.0321522f $X=6.305 $Y=2.24 $X2=0
+ $Y2=0
cc_400 N_A_615_93#_c_329_n N_VPWR_c_1191_n 0.00876084f $X=4.587 $Y=2.2 $X2=0
+ $Y2=0
cc_401 N_A_615_93#_c_330_n N_VPWR_c_1192_n 0.019758f $X=6.305 $Y=2.24 $X2=0
+ $Y2=0
cc_402 N_A_615_93#_M1023_s N_VPWR_c_1181_n 0.00230667f $X=6.16 $Y=2.095 $X2=0
+ $Y2=0
cc_403 N_A_615_93#_c_323_n N_VPWR_c_1181_n 0.00141512f $X=3.765 $Y=1.66 $X2=0
+ $Y2=0
cc_404 N_A_615_93#_c_329_n N_VPWR_c_1181_n 0.0105985f $X=4.587 $Y=2.2 $X2=0
+ $Y2=0
cc_405 N_A_615_93#_c_330_n N_VPWR_c_1181_n 0.012508f $X=6.305 $Y=2.24 $X2=0
+ $Y2=0
cc_406 N_A_615_93#_c_323_n N_A_349_323#_c_1354_n 0.00633805f $X=3.765 $Y=1.66
+ $X2=0 $Y2=0
cc_407 N_A_615_93#_c_323_n N_A_349_323#_c_1355_n 0.00870881f $X=3.765 $Y=1.66
+ $X2=0 $Y2=0
cc_408 N_A_615_93#_c_318_n N_A_349_323#_c_1355_n 0.00157204f $X=3.24 $Y=1.29
+ $X2=0 $Y2=0
cc_409 N_A_615_93#_c_307_n N_VGND_M1019_d 0.0023291f $X=4.15 $Y=1.05 $X2=0 $Y2=0
cc_410 N_A_615_93#_c_317_n N_VGND_M1019_d 0.00149145f $X=3.24 $Y=1.05 $X2=0
+ $Y2=0
cc_411 N_A_615_93#_c_305_n N_VGND_c_1436_n 0.00323048f $X=3.15 $Y=1.125 $X2=0
+ $Y2=0
cc_412 N_A_615_93#_c_307_n N_VGND_c_1436_n 0.0158246f $X=4.15 $Y=1.05 $X2=0
+ $Y2=0
cc_413 N_A_615_93#_c_308_n N_VGND_c_1436_n 0.00813467f $X=4.315 $Y=0.805 $X2=0
+ $Y2=0
cc_414 N_A_615_93#_c_310_n N_VGND_c_1436_n 0.00673184f $X=4.48 $Y=0.35 $X2=0
+ $Y2=0
cc_415 N_A_615_93#_c_317_n N_VGND_c_1436_n 0.0102866f $X=3.24 $Y=1.05 $X2=0
+ $Y2=0
cc_416 N_A_615_93#_c_318_n N_VGND_c_1436_n 6.5957e-19 $X=3.24 $Y=1.29 $X2=0
+ $Y2=0
cc_417 N_A_615_93#_c_309_n N_VGND_c_1437_n 0.0141601f $X=5.31 $Y=0.35 $X2=0
+ $Y2=0
cc_418 N_A_615_93#_c_311_n N_VGND_c_1437_n 0.0285568f $X=5.395 $Y=1.335 $X2=0
+ $Y2=0
cc_419 N_A_615_93#_c_312_n N_VGND_c_1437_n 0.0151601f $X=6.57 $Y=1.42 $X2=0
+ $Y2=0
cc_420 N_A_615_93#_c_309_n N_VGND_c_1441_n 0.0617104f $X=5.31 $Y=0.35 $X2=0
+ $Y2=0
cc_421 N_A_615_93#_c_310_n N_VGND_c_1441_n 0.0222893f $X=4.48 $Y=0.35 $X2=0
+ $Y2=0
cc_422 N_A_615_93#_c_305_n N_VGND_c_1450_n 9.39239e-19 $X=3.15 $Y=1.125 $X2=0
+ $Y2=0
cc_423 N_A_615_93#_c_309_n N_VGND_c_1450_n 0.0336003f $X=5.31 $Y=0.35 $X2=0
+ $Y2=0
cc_424 N_A_615_93#_c_310_n N_VGND_c_1450_n 0.0114626f $X=4.48 $Y=0.35 $X2=0
+ $Y2=0
cc_425 N_A_615_93#_c_307_n A_763_119# 0.00366293f $X=4.15 $Y=1.05 $X2=-0.19
+ $Y2=-0.245
cc_426 N_A_615_93#_c_311_n A_1049_125# 0.00348527f $X=5.395 $Y=1.335 $X2=-0.19
+ $Y2=-0.245
cc_427 N_A_615_93#_c_311_n N_A_1232_153#_c_1567_n 0.00236321f $X=5.395 $Y=1.335
+ $X2=0 $Y2=0
cc_428 N_A_615_93#_c_312_n N_A_1232_153#_c_1567_n 0.0197026f $X=6.57 $Y=1.42
+ $X2=0 $Y2=0
cc_429 N_A_615_93#_c_314_n N_A_1232_153#_c_1567_n 0.0255883f $X=6.655 $Y=1.335
+ $X2=0 $Y2=0
cc_430 N_A_615_93#_c_316_n N_A_1232_153#_c_1567_n 0.0134723f $X=6.74 $Y=0.7
+ $X2=0 $Y2=0
cc_431 N_A_615_93#_c_315_n N_A_1232_153#_c_1568_n 0.0350179f $X=7.27 $Y=0.7
+ $X2=0 $Y2=0
cc_432 N_A_615_93#_c_316_n N_A_1232_153#_c_1568_n 0.012842f $X=6.74 $Y=0.7 $X2=0
+ $Y2=0
cc_433 N_A_615_93#_c_321_n N_A_1232_153#_c_1568_n 0.0239044f $X=7.435 $Y=0.7
+ $X2=0 $Y2=0
cc_434 N_A_615_93#_c_321_n N_A_1232_153#_c_1570_n 0.00752967f $X=7.435 $Y=0.7
+ $X2=0 $Y2=0
cc_435 N_A_455_85#_c_491_n N_A_27_403#_c_588_n 0.00156995f $X=2.495 $Y=1.595
+ $X2=0 $Y2=0
cc_436 N_A_455_85#_c_491_n N_A_27_403#_M1026_g 0.00407956f $X=2.495 $Y=1.595
+ $X2=0 $Y2=0
cc_437 N_A_455_85#_c_487_n N_A_27_403#_M1016_g 0.010908f $X=2.495 $Y=0.72 $X2=0
+ $Y2=0
cc_438 N_A_455_85#_M1027_g N_A_27_403#_c_591_n 0.0171388f $X=4.295 $Y=2.235
+ $X2=0 $Y2=0
cc_439 N_A_455_85#_c_486_n N_A_27_403#_c_575_n 0.0017096f $X=4.295 $Y=1.575
+ $X2=0 $Y2=0
cc_440 N_A_455_85#_c_491_n N_A_511_218#_M1008_g 0.00700125f $X=2.495 $Y=1.595
+ $X2=0 $Y2=0
cc_441 N_A_455_85#_c_487_n N_A_511_218#_M1008_g 0.0122009f $X=2.495 $Y=0.72
+ $X2=0 $Y2=0
cc_442 N_A_455_85#_c_493_n N_A_511_218#_M1008_g 0.0147129f $X=4.045 $Y=1.72
+ $X2=0 $Y2=0
cc_443 N_A_455_85#_c_487_n N_A_511_218#_M1029_g 0.00658707f $X=2.495 $Y=0.72
+ $X2=0 $Y2=0
cc_444 N_A_455_85#_c_482_n N_A_511_218#_c_748_n 0.0104164f $X=3.74 $Y=1.12 $X2=0
+ $Y2=0
cc_445 N_A_455_85#_c_485_n N_A_511_218#_c_748_n 0.0101494f $X=4.1 $Y=1.12 $X2=0
+ $Y2=0
cc_446 N_A_455_85#_c_487_n N_A_511_218#_c_751_n 0.00753066f $X=2.495 $Y=0.72
+ $X2=0 $Y2=0
cc_447 N_A_455_85#_c_493_n N_A_511_218#_c_751_n 0.00118352f $X=4.045 $Y=1.72
+ $X2=0 $Y2=0
cc_448 N_A_455_85#_c_486_n N_A_511_218#_c_752_n 2.58645e-19 $X=4.295 $Y=1.575
+ $X2=0 $Y2=0
cc_449 N_A_455_85#_c_493_n N_VPWR_M1004_d 0.00105617f $X=4.045 $Y=1.72 $X2=0
+ $Y2=0
cc_450 N_A_455_85#_c_488_n N_VPWR_M1004_d 7.63256e-19 $X=4.265 $Y=1.41 $X2=0
+ $Y2=0
cc_451 N_A_455_85#_c_486_n N_VPWR_c_1183_n 2.114e-19 $X=4.295 $Y=1.575 $X2=0
+ $Y2=0
cc_452 N_A_455_85#_M1027_g N_VPWR_c_1183_n 0.0210642f $X=4.295 $Y=2.235 $X2=0
+ $Y2=0
cc_453 N_A_455_85#_c_493_n N_VPWR_c_1183_n 0.00931009f $X=4.045 $Y=1.72 $X2=0
+ $Y2=0
cc_454 N_A_455_85#_c_488_n N_VPWR_c_1183_n 0.0075855f $X=4.265 $Y=1.41 $X2=0
+ $Y2=0
cc_455 N_A_455_85#_M1027_g N_VPWR_c_1181_n 0.00141512f $X=4.295 $Y=2.235 $X2=0
+ $Y2=0
cc_456 N_A_455_85#_c_493_n N_A_239_403#_M1008_d 0.011496f $X=4.045 $Y=1.72 $X2=0
+ $Y2=0
cc_457 N_A_455_85#_c_491_n N_A_239_403#_c_1301_n 0.00804704f $X=2.495 $Y=1.595
+ $X2=0 $Y2=0
cc_458 N_A_455_85#_c_487_n N_A_239_403#_c_1301_n 0.0356584f $X=2.495 $Y=0.72
+ $X2=0 $Y2=0
cc_459 N_A_455_85#_c_487_n N_A_239_403#_c_1302_n 0.0180055f $X=2.495 $Y=0.72
+ $X2=0 $Y2=0
cc_460 N_A_455_85#_c_493_n N_A_239_403#_c_1306_n 0.0195261f $X=4.045 $Y=1.72
+ $X2=0 $Y2=0
cc_461 N_A_455_85#_M1026_d N_A_239_403#_c_1323_n 0.00378666f $X=2.275 $Y=1.615
+ $X2=0 $Y2=0
cc_462 N_A_455_85#_c_491_n N_A_239_403#_c_1323_n 0.0211126f $X=2.495 $Y=1.595
+ $X2=0 $Y2=0
cc_463 N_A_455_85#_c_493_n N_A_239_403#_c_1323_n 0.00633479f $X=4.045 $Y=1.72
+ $X2=0 $Y2=0
cc_464 N_A_455_85#_c_493_n N_A_349_323#_M1004_s 0.00242809f $X=4.045 $Y=1.72
+ $X2=0 $Y2=0
cc_465 N_A_455_85#_M1026_d N_A_349_323#_c_1354_n 0.00486181f $X=2.275 $Y=1.615
+ $X2=0 $Y2=0
cc_466 N_A_455_85#_c_493_n N_A_349_323#_c_1354_n 0.00686828f $X=4.045 $Y=1.72
+ $X2=0 $Y2=0
cc_467 N_A_455_85#_c_493_n N_A_349_323#_c_1355_n 0.0210355f $X=4.045 $Y=1.72
+ $X2=0 $Y2=0
cc_468 N_A_455_85#_c_482_n N_VGND_c_1436_n 0.00310544f $X=3.74 $Y=1.12 $X2=0
+ $Y2=0
cc_469 N_A_455_85#_c_487_n N_VGND_c_1436_n 0.00629449f $X=2.495 $Y=0.72 $X2=0
+ $Y2=0
cc_470 N_A_455_85#_c_487_n N_VGND_c_1446_n 0.0119784f $X=2.495 $Y=0.72 $X2=0
+ $Y2=0
cc_471 N_A_455_85#_c_482_n N_VGND_c_1450_n 9.39239e-19 $X=3.74 $Y=1.12 $X2=0
+ $Y2=0
cc_472 N_A_455_85#_c_485_n N_VGND_c_1450_n 7.85159e-19 $X=4.1 $Y=1.12 $X2=0
+ $Y2=0
cc_473 N_A_455_85#_c_487_n N_VGND_c_1450_n 0.011704f $X=2.495 $Y=0.72 $X2=0
+ $Y2=0
cc_474 N_A_27_403#_c_588_n N_A_511_218#_M1008_g 0.0301068f $X=2.15 $Y=1.61 $X2=0
+ $Y2=0
cc_475 N_A_27_403#_c_591_n N_A_511_218#_M1008_g 0.00961497f $X=5.875 $Y=3.15
+ $X2=0 $Y2=0
cc_476 N_A_27_403#_M1016_g N_A_511_218#_M1029_g 0.0157866f $X=2.2 $Y=0.635 $X2=0
+ $Y2=0
cc_477 N_A_27_403#_c_573_n N_A_511_218#_c_748_n 0.00737233f $X=5.17 $Y=1.12
+ $X2=0 $Y2=0
cc_478 N_A_27_403#_c_576_n N_A_511_218#_c_748_n 0.00879826f $X=5.53 $Y=1.12
+ $X2=0 $Y2=0
cc_479 N_A_27_403#_M1022_g N_A_511_218#_c_748_n 0.00392393f $X=6.62 $Y=0.975
+ $X2=0 $Y2=0
cc_480 N_A_27_403#_M1023_g N_A_511_218#_M1005_g 0.0257151f $X=6.57 $Y=2.595
+ $X2=0 $Y2=0
cc_481 N_A_27_403#_M1022_g N_A_511_218#_M1031_g 0.0162159f $X=6.62 $Y=0.975
+ $X2=0 $Y2=0
cc_482 N_A_27_403#_M1016_g N_A_511_218#_c_751_n 0.0301068f $X=2.2 $Y=0.635 $X2=0
+ $Y2=0
cc_483 N_A_27_403#_c_573_n N_A_511_218#_c_752_n 0.00953708f $X=5.17 $Y=1.12
+ $X2=0 $Y2=0
cc_484 N_A_27_403#_c_575_n N_A_511_218#_c_752_n 0.00530963f $X=5.245 $Y=1.195
+ $X2=0 $Y2=0
cc_485 N_A_27_403#_c_576_n N_A_511_218#_c_752_n 2.73212e-19 $X=5.53 $Y=1.12
+ $X2=0 $Y2=0
cc_486 N_A_27_403#_c_583_n N_A_511_218#_c_752_n 0.00813344f $X=5.435 $Y=1.555
+ $X2=0 $Y2=0
cc_487 N_A_27_403#_c_573_n N_A_511_218#_c_753_n 0.00581406f $X=5.17 $Y=1.12
+ $X2=0 $Y2=0
cc_488 N_A_27_403#_c_574_n N_A_511_218#_c_759_n 2.25854e-19 $X=5.455 $Y=1.195
+ $X2=0 $Y2=0
cc_489 N_A_27_403#_c_575_n N_A_511_218#_c_759_n 0.00459634f $X=5.245 $Y=1.195
+ $X2=0 $Y2=0
cc_490 N_A_27_403#_c_592_n N_A_511_218#_c_759_n 0.00320109f $X=5.39 $Y=1.63
+ $X2=0 $Y2=0
cc_491 N_A_27_403#_c_579_n N_A_511_218#_c_759_n 3.14743e-19 $X=5.95 $Y=3.075
+ $X2=0 $Y2=0
cc_492 N_A_27_403#_M1023_g N_A_511_218#_c_754_n 5.37894e-19 $X=6.57 $Y=2.595
+ $X2=0 $Y2=0
cc_493 N_A_27_403#_c_586_n N_A_511_218#_c_754_n 4.77865e-19 $X=6.57 $Y=1.555
+ $X2=0 $Y2=0
cc_494 N_A_27_403#_c_586_n N_A_511_218#_c_755_n 0.0179697f $X=6.57 $Y=1.555
+ $X2=0 $Y2=0
cc_495 N_A_27_403#_c_592_n N_A_511_218#_c_762_n 0.0132109f $X=5.39 $Y=1.63 $X2=0
+ $Y2=0
cc_496 N_A_27_403#_c_578_n N_A_511_218#_c_762_n 0.00468915f $X=5.875 $Y=1.555
+ $X2=0 $Y2=0
cc_497 N_A_27_403#_c_579_n N_A_511_218#_c_762_n 0.0117455f $X=5.95 $Y=3.075
+ $X2=0 $Y2=0
cc_498 N_A_27_403#_c_580_n N_A_511_218#_c_762_n 0.00529981f $X=6.445 $Y=1.555
+ $X2=0 $Y2=0
cc_499 N_A_27_403#_M1023_g N_A_511_218#_c_762_n 0.0215893f $X=6.57 $Y=2.595
+ $X2=0 $Y2=0
cc_500 N_A_27_403#_M1022_g N_A_1339_153#_c_1033_n 9.79166e-19 $X=6.62 $Y=0.975
+ $X2=0 $Y2=0
cc_501 N_A_27_403#_M1022_g N_A_1339_153#_c_1021_n 6.96004e-19 $X=6.62 $Y=0.975
+ $X2=0 $Y2=0
cc_502 N_A_27_403#_M1023_g N_A_1339_153#_c_1040_n 0.0196024f $X=6.57 $Y=2.595
+ $X2=0 $Y2=0
cc_503 N_A_27_403#_c_613_n N_VPWR_M1013_d 0.00809719f $X=1.15 $Y=2.51 $X2=-0.19
+ $Y2=-0.245
cc_504 N_A_27_403#_c_601_n N_VPWR_c_1182_n 0.0171316f $X=0.275 $Y=2.87 $X2=0
+ $Y2=0
cc_505 N_A_27_403#_c_613_n N_VPWR_c_1182_n 0.0156554f $X=1.15 $Y=2.51 $X2=0
+ $Y2=0
cc_506 N_A_27_403#_c_602_n N_VPWR_c_1182_n 0.022106f $X=1.32 $Y=2.92 $X2=0 $Y2=0
cc_507 N_A_27_403#_c_591_n N_VPWR_c_1183_n 0.0254328f $X=5.875 $Y=3.15 $X2=0
+ $Y2=0
cc_508 N_A_27_403#_c_591_n N_VPWR_c_1184_n 0.024046f $X=5.875 $Y=3.15 $X2=0
+ $Y2=0
cc_509 N_A_27_403#_c_592_n N_VPWR_c_1184_n 0.018667f $X=5.39 $Y=1.63 $X2=0 $Y2=0
cc_510 N_A_27_403#_c_579_n N_VPWR_c_1184_n 0.00776438f $X=5.95 $Y=3.075 $X2=0
+ $Y2=0
cc_511 N_A_27_403#_M1023_g N_VPWR_c_1184_n 0.00103792f $X=6.57 $Y=2.595 $X2=0
+ $Y2=0
cc_512 N_A_27_403#_c_613_n N_VPWR_c_1190_n 0.00234125f $X=1.15 $Y=2.51 $X2=0
+ $Y2=0
cc_513 N_A_27_403#_c_602_n N_VPWR_c_1190_n 0.0112553f $X=1.32 $Y=2.92 $X2=0
+ $Y2=0
cc_514 N_A_27_403#_c_603_n N_VPWR_c_1190_n 0.0615798f $X=2.15 $Y=2.94 $X2=0
+ $Y2=0
cc_515 N_A_27_403#_c_604_n N_VPWR_c_1190_n 0.0491628f $X=2.15 $Y=2.94 $X2=0
+ $Y2=0
cc_516 N_A_27_403#_c_591_n N_VPWR_c_1191_n 0.0413469f $X=5.875 $Y=3.15 $X2=0
+ $Y2=0
cc_517 N_A_27_403#_c_591_n N_VPWR_c_1192_n 0.00796123f $X=5.875 $Y=3.15 $X2=0
+ $Y2=0
cc_518 N_A_27_403#_M1023_g N_VPWR_c_1192_n 0.0090344f $X=6.57 $Y=2.595 $X2=0
+ $Y2=0
cc_519 N_A_27_403#_c_591_n N_VPWR_c_1181_n 0.107135f $X=5.875 $Y=3.15 $X2=0
+ $Y2=0
cc_520 N_A_27_403#_c_592_n N_VPWR_c_1181_n 0.00143131f $X=5.39 $Y=1.63 $X2=0
+ $Y2=0
cc_521 N_A_27_403#_M1023_g N_VPWR_c_1181_n 0.0155898f $X=6.57 $Y=2.595 $X2=0
+ $Y2=0
cc_522 N_A_27_403#_c_601_n N_VPWR_c_1181_n 0.0123863f $X=0.275 $Y=2.87 $X2=0
+ $Y2=0
cc_523 N_A_27_403#_c_613_n N_VPWR_c_1181_n 0.00945186f $X=1.15 $Y=2.51 $X2=0
+ $Y2=0
cc_524 N_A_27_403#_c_602_n N_VPWR_c_1181_n 0.00635973f $X=1.32 $Y=2.92 $X2=0
+ $Y2=0
cc_525 N_A_27_403#_c_603_n N_VPWR_c_1181_n 0.0361236f $X=2.15 $Y=2.94 $X2=0
+ $Y2=0
cc_526 N_A_27_403#_c_604_n N_VPWR_c_1181_n 0.0104084f $X=2.15 $Y=2.94 $X2=0
+ $Y2=0
cc_527 N_A_27_403#_c_601_n N_VPWR_c_1196_n 0.0186734f $X=0.275 $Y=2.87 $X2=0
+ $Y2=0
cc_528 N_A_27_403#_c_613_n N_VPWR_c_1196_n 0.00260284f $X=1.15 $Y=2.51 $X2=0
+ $Y2=0
cc_529 N_A_27_403#_c_613_n N_A_239_403#_M1028_d 0.00353026f $X=1.15 $Y=2.51
+ $X2=0 $Y2=0
cc_530 N_A_27_403#_c_614_n N_A_239_403#_M1028_d 0.00679169f $X=1.235 $Y=2.775
+ $X2=0 $Y2=0
cc_531 N_A_27_403#_c_603_n N_A_239_403#_M1028_d 0.00424594f $X=2.15 $Y=2.94
+ $X2=0 $Y2=0
cc_532 N_A_27_403#_c_603_n N_A_239_403#_c_1303_n 0.00744001f $X=2.15 $Y=2.94
+ $X2=0 $Y2=0
cc_533 N_A_27_403#_c_588_n N_A_239_403#_c_1301_n 0.00777098f $X=2.15 $Y=1.61
+ $X2=0 $Y2=0
cc_534 N_A_27_403#_M1016_g N_A_239_403#_c_1301_n 0.00577335f $X=2.2 $Y=0.635
+ $X2=0 $Y2=0
cc_535 N_A_27_403#_M1026_g N_A_239_403#_c_1305_n 0.001056f $X=2.15 $Y=2.115
+ $X2=0 $Y2=0
cc_536 N_A_27_403#_c_613_n N_A_239_403#_c_1305_n 0.00715374f $X=1.15 $Y=2.51
+ $X2=0 $Y2=0
cc_537 N_A_27_403#_c_603_n N_A_239_403#_c_1305_n 0.00600853f $X=2.15 $Y=2.94
+ $X2=0 $Y2=0
cc_538 N_A_27_403#_c_588_n N_A_239_403#_c_1302_n 0.00288804f $X=2.15 $Y=1.61
+ $X2=0 $Y2=0
cc_539 N_A_27_403#_M1016_g N_A_239_403#_c_1302_n 0.00714892f $X=2.2 $Y=0.635
+ $X2=0 $Y2=0
cc_540 N_A_27_403#_M1026_g N_A_239_403#_c_1306_n 3.79235e-19 $X=2.15 $Y=2.115
+ $X2=0 $Y2=0
cc_541 N_A_27_403#_M1026_g N_A_239_403#_c_1323_n 0.0240083f $X=2.15 $Y=2.115
+ $X2=0 $Y2=0
cc_542 N_A_27_403#_M1026_g N_A_349_323#_c_1354_n 0.0121697f $X=2.15 $Y=2.115
+ $X2=0 $Y2=0
cc_543 N_A_27_403#_c_591_n N_A_349_323#_c_1354_n 0.0176105f $X=5.875 $Y=3.15
+ $X2=0 $Y2=0
cc_544 N_A_27_403#_M1026_g N_A_349_323#_c_1356_n 0.00185667f $X=2.15 $Y=2.115
+ $X2=0 $Y2=0
cc_545 N_A_27_403#_c_613_n N_A_349_323#_c_1356_n 0.00839927f $X=1.15 $Y=2.51
+ $X2=0 $Y2=0
cc_546 N_A_27_403#_c_603_n N_A_349_323#_c_1356_n 0.0375473f $X=2.15 $Y=2.94
+ $X2=0 $Y2=0
cc_547 N_A_27_403#_c_576_n N_VGND_c_1437_n 0.00392143f $X=5.53 $Y=1.12 $X2=0
+ $Y2=0
cc_548 N_A_27_403#_c_578_n N_VGND_c_1437_n 0.00119851f $X=5.875 $Y=1.555 $X2=0
+ $Y2=0
cc_549 N_A_27_403#_c_587_n N_VGND_c_1445_n 0.011248f $X=0.335 $Y=0.635 $X2=0
+ $Y2=0
cc_550 N_A_27_403#_M1016_g N_VGND_c_1446_n 0.00514022f $X=2.2 $Y=0.635 $X2=0
+ $Y2=0
cc_551 N_A_27_403#_M1016_g N_VGND_c_1450_n 0.00528353f $X=2.2 $Y=0.635 $X2=0
+ $Y2=0
cc_552 N_A_27_403#_c_576_n N_VGND_c_1450_n 7.94319e-19 $X=5.53 $Y=1.12 $X2=0
+ $Y2=0
cc_553 N_A_27_403#_c_587_n N_VGND_c_1450_n 0.0109904f $X=0.335 $Y=0.635 $X2=0
+ $Y2=0
cc_554 N_A_27_403#_c_576_n N_A_1232_153#_c_1567_n 0.00245654f $X=5.53 $Y=1.12
+ $X2=0 $Y2=0
cc_555 N_A_27_403#_c_580_n N_A_1232_153#_c_1567_n 0.00140028f $X=6.445 $Y=1.555
+ $X2=0 $Y2=0
cc_556 N_A_27_403#_M1022_g N_A_1232_153#_c_1567_n 0.0102824f $X=6.62 $Y=0.975
+ $X2=0 $Y2=0
cc_557 N_A_27_403#_M1022_g N_A_1232_153#_c_1568_n 9.74623e-19 $X=6.62 $Y=0.975
+ $X2=0 $Y2=0
cc_558 N_A_511_218#_M1005_g N_A_1507_321#_M1021_g 0.053006f $X=7.1 $Y=2.595
+ $X2=0 $Y2=0
cc_559 N_A_511_218#_M1031_g N_A_1507_321#_c_875_n 0.00835696f $X=7.22 $Y=1.065
+ $X2=0 $Y2=0
cc_560 N_A_511_218#_c_754_n N_A_1507_321#_c_883_n 3.21212e-19 $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_561 N_A_511_218#_c_755_n N_A_1507_321#_c_883_n 0.0174944f $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_562 N_A_511_218#_M1005_g N_A_1339_153#_c_1046_n 0.018757f $X=7.1 $Y=2.595
+ $X2=0 $Y2=0
cc_563 N_A_511_218#_c_754_n N_A_1339_153#_c_1046_n 0.0167046f $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_564 N_A_511_218#_c_755_n N_A_1339_153#_c_1046_n 0.00189649f $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_565 N_A_511_218#_M1031_g N_A_1339_153#_c_1020_n 0.0140502f $X=7.22 $Y=1.065
+ $X2=0 $Y2=0
cc_566 N_A_511_218#_c_754_n N_A_1339_153#_c_1020_n 0.0120793f $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_567 N_A_511_218#_c_755_n N_A_1339_153#_c_1020_n 0.00145404f $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_568 N_A_511_218#_c_754_n N_A_1339_153#_c_1021_n 0.012122f $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_569 N_A_511_218#_c_755_n N_A_1339_153#_c_1021_n 0.00404423f $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_570 N_A_511_218#_c_762_n N_A_1339_153#_c_1021_n 9.11266e-19 $X=6.935 $Y=1.775
+ $X2=0 $Y2=0
cc_571 N_A_511_218#_M1005_g N_A_1339_153#_c_1022_n 0.00360917f $X=7.1 $Y=2.595
+ $X2=0 $Y2=0
cc_572 N_A_511_218#_M1031_g N_A_1339_153#_c_1022_n 0.00669185f $X=7.22 $Y=1.065
+ $X2=0 $Y2=0
cc_573 N_A_511_218#_c_754_n N_A_1339_153#_c_1022_n 0.0237105f $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_574 N_A_511_218#_M1005_g N_A_1339_153#_c_1040_n 0.0198323f $X=7.1 $Y=2.595
+ $X2=0 $Y2=0
cc_575 N_A_511_218#_c_754_n N_A_1339_153#_c_1040_n 0.00329453f $X=7.1 $Y=1.77
+ $X2=0 $Y2=0
cc_576 N_A_511_218#_c_762_n N_A_1339_153#_c_1040_n 0.013477f $X=6.935 $Y=1.775
+ $X2=0 $Y2=0
cc_577 N_A_511_218#_c_762_n N_VPWR_M1033_d 0.00294042f $X=6.935 $Y=1.775 $X2=0
+ $Y2=0
cc_578 N_A_511_218#_M1005_g N_VPWR_c_1192_n 0.00939541f $X=7.1 $Y=2.595 $X2=0
+ $Y2=0
cc_579 N_A_511_218#_M1008_g N_VPWR_c_1181_n 0.00161547f $X=2.68 $Y=2.115 $X2=0
+ $Y2=0
cc_580 N_A_511_218#_M1005_g N_VPWR_c_1181_n 0.0163381f $X=7.1 $Y=2.595 $X2=0
+ $Y2=0
cc_581 N_A_511_218#_M1008_g N_A_239_403#_c_1306_n 0.00286506f $X=2.68 $Y=2.115
+ $X2=0 $Y2=0
cc_582 N_A_511_218#_M1008_g N_A_239_403#_c_1323_n 0.0125613f $X=2.68 $Y=2.115
+ $X2=0 $Y2=0
cc_583 N_A_511_218#_M1008_g N_A_349_323#_c_1354_n 0.0222936f $X=2.68 $Y=2.115
+ $X2=0 $Y2=0
cc_584 N_A_511_218#_M1008_g N_A_349_323#_c_1355_n 0.0045152f $X=2.68 $Y=2.115
+ $X2=0 $Y2=0
cc_585 N_A_511_218#_M1029_g N_VGND_c_1436_n 0.00588979f $X=2.79 $Y=0.805 $X2=0
+ $Y2=0
cc_586 N_A_511_218#_c_748_n N_VGND_c_1436_n 0.0256012f $X=7.145 $Y=0.18 $X2=0
+ $Y2=0
cc_587 N_A_511_218#_c_748_n N_VGND_c_1437_n 0.0216291f $X=7.145 $Y=0.18 $X2=0
+ $Y2=0
cc_588 N_A_511_218#_c_748_n N_VGND_c_1441_n 0.0523327f $X=7.145 $Y=0.18 $X2=0
+ $Y2=0
cc_589 N_A_511_218#_c_749_n N_VGND_c_1446_n 0.0207992f $X=2.865 $Y=0.18 $X2=0
+ $Y2=0
cc_590 N_A_511_218#_c_748_n N_VGND_c_1447_n 0.0323834f $X=7.145 $Y=0.18 $X2=0
+ $Y2=0
cc_591 N_A_511_218#_c_748_n N_VGND_c_1450_n 0.122719f $X=7.145 $Y=0.18 $X2=0
+ $Y2=0
cc_592 N_A_511_218#_c_749_n N_VGND_c_1450_n 0.0116041f $X=2.865 $Y=0.18 $X2=0
+ $Y2=0
cc_593 N_A_511_218#_c_748_n N_A_1232_153#_c_1568_n 0.0134088f $X=7.145 $Y=0.18
+ $X2=0 $Y2=0
cc_594 N_A_511_218#_M1031_g N_A_1232_153#_c_1568_n 0.0118022f $X=7.22 $Y=1.065
+ $X2=0 $Y2=0
cc_595 N_A_511_218#_c_748_n N_A_1232_153#_c_1569_n 0.00615835f $X=7.145 $Y=0.18
+ $X2=0 $Y2=0
cc_596 N_A_511_218#_M1031_g N_A_1232_153#_c_1570_n 0.00540533f $X=7.22 $Y=1.065
+ $X2=0 $Y2=0
cc_597 N_A_1507_321#_M1021_g N_A_1339_153#_M1035_g 0.0156712f $X=7.66 $Y=2.595
+ $X2=0 $Y2=0
cc_598 N_A_1507_321#_c_887_n N_A_1339_153#_M1035_g 0.00209397f $X=7.96 $Y=1.77
+ $X2=0 $Y2=0
cc_599 N_A_1507_321#_c_888_n N_A_1339_153#_M1035_g 0.0197127f $X=8.59 $Y=2.105
+ $X2=0 $Y2=0
cc_600 N_A_1507_321#_c_890_n N_A_1339_153#_M1035_g 0.0284428f $X=8.755 $Y=2.24
+ $X2=0 $Y2=0
cc_601 N_A_1507_321#_c_876_n N_A_1339_153#_M1035_g 0.00590404f $X=8.96 $Y=2.02
+ $X2=0 $Y2=0
cc_602 N_A_1507_321#_c_892_n N_A_1339_153#_M1035_g 0.00237914f $X=8.817 $Y=2.105
+ $X2=0 $Y2=0
cc_603 N_A_1507_321#_c_867_n N_A_1339_153#_M1024_g 0.00814151f $X=8.05 $Y=1.605
+ $X2=0 $Y2=0
cc_604 N_A_1507_321#_c_868_n N_A_1339_153#_M1024_g 0.0179302f $X=8.205 $Y=0.78
+ $X2=0 $Y2=0
cc_605 N_A_1507_321#_c_876_n N_A_1339_153#_M1024_g 0.00891148f $X=8.96 $Y=2.02
+ $X2=0 $Y2=0
cc_606 N_A_1507_321#_c_881_n N_A_1339_153#_M1024_g 0.00136516f $X=9.375 $Y=0.495
+ $X2=0 $Y2=0
cc_607 N_A_1507_321#_c_876_n N_A_1339_153#_c_1017_n 0.00952491f $X=8.96 $Y=2.02
+ $X2=0 $Y2=0
cc_608 N_A_1507_321#_c_892_n N_A_1339_153#_c_1017_n 0.00449085f $X=8.817
+ $Y=2.105 $X2=0 $Y2=0
cc_609 N_A_1507_321#_c_882_n N_A_1339_153#_c_1017_n 0.0014323f $X=11.2 $Y=1.42
+ $X2=0 $Y2=0
cc_610 N_A_1507_321#_c_876_n N_A_1339_153#_M1015_g 0.0113574f $X=8.96 $Y=2.02
+ $X2=0 $Y2=0
cc_611 N_A_1507_321#_c_881_n N_A_1339_153#_M1015_g 0.0119616f $X=9.375 $Y=0.495
+ $X2=0 $Y2=0
cc_612 N_A_1507_321#_c_867_n N_A_1339_153#_c_1019_n 0.0210932f $X=8.05 $Y=1.605
+ $X2=0 $Y2=0
cc_613 N_A_1507_321#_c_892_n N_A_1339_153#_c_1028_n 0.00137925f $X=8.817
+ $Y=2.105 $X2=0 $Y2=0
cc_614 N_A_1507_321#_c_883_n N_A_1339_153#_c_1028_n 0.0210932f $X=8.05 $Y=1.77
+ $X2=0 $Y2=0
cc_615 N_A_1507_321#_M1021_g N_A_1339_153#_c_1046_n 0.0126024f $X=7.66 $Y=2.595
+ $X2=0 $Y2=0
cc_616 N_A_1507_321#_M1021_g N_A_1339_153#_c_1022_n 0.00422249f $X=7.66 $Y=2.595
+ $X2=0 $Y2=0
cc_617 N_A_1507_321#_c_867_n N_A_1339_153#_c_1022_n 0.00324183f $X=8.05 $Y=1.605
+ $X2=0 $Y2=0
cc_618 N_A_1507_321#_c_887_n N_A_1339_153#_c_1022_n 0.0279039f $X=7.96 $Y=1.77
+ $X2=0 $Y2=0
cc_619 N_A_1507_321#_c_889_n N_A_1339_153#_c_1022_n 0.00636896f $X=8.125
+ $Y=2.105 $X2=0 $Y2=0
cc_620 N_A_1507_321#_c_883_n N_A_1339_153#_c_1022_n 0.0106041f $X=8.05 $Y=1.77
+ $X2=0 $Y2=0
cc_621 N_A_1507_321#_c_867_n N_A_1339_153#_c_1023_n 0.0131012f $X=8.05 $Y=1.605
+ $X2=0 $Y2=0
cc_622 N_A_1507_321#_c_875_n N_A_1339_153#_c_1023_n 0.00507375f $X=8.205
+ $Y=0.855 $X2=0 $Y2=0
cc_623 N_A_1507_321#_c_887_n N_A_1339_153#_c_1023_n 0.0242022f $X=7.96 $Y=1.77
+ $X2=0 $Y2=0
cc_624 N_A_1507_321#_c_888_n N_A_1339_153#_c_1023_n 0.00762782f $X=8.59 $Y=2.105
+ $X2=0 $Y2=0
cc_625 N_A_1507_321#_c_883_n N_A_1339_153#_c_1023_n 0.0114843f $X=8.05 $Y=1.77
+ $X2=0 $Y2=0
cc_626 N_A_1507_321#_M1021_g N_A_1339_153#_c_1040_n 0.00333521f $X=7.66 $Y=2.595
+ $X2=0 $Y2=0
cc_627 N_A_1507_321#_c_867_n N_A_1339_153#_c_1025_n 0.00271072f $X=8.05 $Y=1.605
+ $X2=0 $Y2=0
cc_628 N_A_1507_321#_c_887_n N_A_1339_153#_c_1025_n 0.0127899f $X=7.96 $Y=1.77
+ $X2=0 $Y2=0
cc_629 N_A_1507_321#_c_888_n N_A_1339_153#_c_1025_n 0.0162415f $X=8.59 $Y=2.105
+ $X2=0 $Y2=0
cc_630 N_A_1507_321#_c_876_n N_A_1339_153#_c_1025_n 0.0483551f $X=8.96 $Y=2.02
+ $X2=0 $Y2=0
cc_631 N_A_1507_321#_c_892_n N_A_1339_153#_c_1025_n 0.00875454f $X=8.817
+ $Y=2.105 $X2=0 $Y2=0
cc_632 N_A_1507_321#_c_887_n N_A_1339_153#_c_1026_n 0.00147474f $X=7.96 $Y=1.77
+ $X2=0 $Y2=0
cc_633 N_A_1507_321#_c_876_n N_A_1339_153#_c_1026_n 0.0118547f $X=8.96 $Y=2.02
+ $X2=0 $Y2=0
cc_634 N_A_1507_321#_c_879_n N_A_2062_367#_c_1121_n 0.00128405f $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_635 N_A_1507_321#_c_880_n N_A_2062_367#_c_1121_n 0.0181517f $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_636 N_A_1507_321#_M1007_g N_A_2062_367#_c_1129_n 2.4118e-19 $X=9.655 $Y=2.335
+ $X2=0 $Y2=0
cc_637 N_A_1507_321#_M1014_g N_A_2062_367#_c_1129_n 0.0160832f $X=10.185
+ $Y=2.335 $X2=0 $Y2=0
cc_638 N_A_1507_321#_c_879_n N_A_2062_367#_c_1130_n 0.0827147f $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_639 N_A_1507_321#_c_882_n N_A_2062_367#_c_1130_n 0.027759f $X=11.2 $Y=1.42
+ $X2=0 $Y2=0
cc_640 N_A_1507_321#_M1007_g N_A_2062_367#_c_1131_n 2.50179e-19 $X=9.655
+ $Y=2.335 $X2=0 $Y2=0
cc_641 N_A_1507_321#_M1014_g N_A_2062_367#_c_1131_n 0.00523404f $X=10.185
+ $Y=2.335 $X2=0 $Y2=0
cc_642 N_A_1507_321#_c_879_n N_A_2062_367#_c_1131_n 0.0265437f $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_643 N_A_1507_321#_c_882_n N_A_2062_367#_c_1131_n 0.00787003f $X=11.2 $Y=1.42
+ $X2=0 $Y2=0
cc_644 N_A_1507_321#_c_879_n N_A_2062_367#_c_1122_n 0.018717f $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_645 N_A_1507_321#_c_880_n N_A_2062_367#_c_1122_n 0.00579191f $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_646 N_A_1507_321#_c_879_n N_A_2062_367#_c_1123_n 0.0197915f $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_647 N_A_1507_321#_c_880_n N_A_2062_367#_c_1123_n 4.14154e-19 $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_648 N_A_1507_321#_M1003_g N_A_2062_367#_c_1125_n 0.00125204f $X=10.765
+ $Y=0.845 $X2=0 $Y2=0
cc_649 N_A_1507_321#_M1012_g N_A_2062_367#_c_1125_n 0.00946161f $X=11.125
+ $Y=0.845 $X2=0 $Y2=0
cc_650 N_A_1507_321#_c_879_n N_A_2062_367#_c_1125_n 0.025518f $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_651 N_A_1507_321#_c_880_n N_A_2062_367#_c_1125_n 0.00693392f $X=11.6 $Y=1.42
+ $X2=0 $Y2=0
cc_652 N_A_1507_321#_c_888_n N_VPWR_M1021_d 0.00718597f $X=8.59 $Y=2.105 $X2=0
+ $Y2=0
cc_653 N_A_1507_321#_c_889_n N_VPWR_M1021_d 0.00435561f $X=8.125 $Y=2.105 $X2=0
+ $Y2=0
cc_654 N_A_1507_321#_M1021_g N_VPWR_c_1185_n 0.00390885f $X=7.66 $Y=2.595 $X2=0
+ $Y2=0
cc_655 N_A_1507_321#_c_889_n N_VPWR_c_1185_n 0.0240558f $X=8.125 $Y=2.105 $X2=0
+ $Y2=0
cc_656 N_A_1507_321#_c_890_n N_VPWR_c_1185_n 0.0253356f $X=8.755 $Y=2.24 $X2=0
+ $Y2=0
cc_657 N_A_1507_321#_c_883_n N_VPWR_c_1185_n 0.00138403f $X=8.05 $Y=1.77 $X2=0
+ $Y2=0
cc_658 N_A_1507_321#_M1007_g N_VPWR_c_1186_n 0.0248782f $X=9.655 $Y=2.335 $X2=0
+ $Y2=0
cc_659 N_A_1507_321#_M1014_g N_VPWR_c_1186_n 0.0258202f $X=10.185 $Y=2.335 $X2=0
+ $Y2=0
cc_660 N_A_1507_321#_c_964_p N_VPWR_c_1186_n 0.0218475f $X=10.24 $Y=1.42 $X2=0
+ $Y2=0
cc_661 N_A_1507_321#_c_882_n N_VPWR_c_1186_n 0.00251517f $X=11.2 $Y=1.42 $X2=0
+ $Y2=0
cc_662 N_A_1507_321#_M1014_g N_VPWR_c_1188_n 0.00714707f $X=10.185 $Y=2.335
+ $X2=0 $Y2=0
cc_663 N_A_1507_321#_M1021_g N_VPWR_c_1192_n 0.00975641f $X=7.66 $Y=2.595 $X2=0
+ $Y2=0
cc_664 N_A_1507_321#_M1007_g N_VPWR_c_1193_n 0.00714193f $X=9.655 $Y=2.335 $X2=0
+ $Y2=0
cc_665 N_A_1507_321#_c_890_n N_VPWR_c_1193_n 0.0281861f $X=8.755 $Y=2.24 $X2=0
+ $Y2=0
cc_666 N_A_1507_321#_M1035_d N_VPWR_c_1181_n 0.0023218f $X=8.615 $Y=2.095 $X2=0
+ $Y2=0
cc_667 N_A_1507_321#_M1021_g N_VPWR_c_1181_n 0.0175132f $X=7.66 $Y=2.595 $X2=0
+ $Y2=0
cc_668 N_A_1507_321#_M1007_g N_VPWR_c_1181_n 0.00763694f $X=9.655 $Y=2.335 $X2=0
+ $Y2=0
cc_669 N_A_1507_321#_M1014_g N_VPWR_c_1181_n 0.00763694f $X=10.185 $Y=2.335
+ $X2=0 $Y2=0
cc_670 N_A_1507_321#_c_890_n N_VPWR_c_1181_n 0.0173447f $X=8.755 $Y=2.24 $X2=0
+ $Y2=0
cc_671 N_A_1507_321#_M1011_g N_Q_c_1390_n 0.0068274f $X=9.975 $Y=0.845 $X2=0
+ $Y2=0
cc_672 N_A_1507_321#_M1017_g N_Q_c_1390_n 3.61416e-19 $X=10.335 $Y=0.845 $X2=0
+ $Y2=0
cc_673 N_A_1507_321#_c_876_n N_Q_c_1390_n 0.0188273f $X=8.96 $Y=2.02 $X2=0 $Y2=0
cc_674 N_A_1507_321#_c_877_n N_Q_c_1390_n 0.0330818f $X=10.105 $Y=0.35 $X2=0
+ $Y2=0
cc_675 N_A_1507_321#_c_878_n N_Q_c_1390_n 0.0186973f $X=10.19 $Y=1.255 $X2=0
+ $Y2=0
cc_676 N_A_1507_321#_c_881_n N_Q_c_1390_n 0.0209316f $X=9.375 $Y=0.495 $X2=0
+ $Y2=0
cc_677 N_A_1507_321#_c_964_p N_Q_c_1390_n 0.0147547f $X=10.24 $Y=1.42 $X2=0
+ $Y2=0
cc_678 N_A_1507_321#_c_882_n N_Q_c_1390_n 0.0123228f $X=11.2 $Y=1.42 $X2=0 $Y2=0
cc_679 N_A_1507_321#_M1007_g Q 0.0290362f $X=9.655 $Y=2.335 $X2=0 $Y2=0
cc_680 N_A_1507_321#_M1011_g Q 0.00344039f $X=9.975 $Y=0.845 $X2=0 $Y2=0
cc_681 N_A_1507_321#_M1014_g Q 0.00128533f $X=10.185 $Y=2.335 $X2=0 $Y2=0
cc_682 N_A_1507_321#_c_890_n Q 0.0573372f $X=8.755 $Y=2.24 $X2=0 $Y2=0
cc_683 N_A_1507_321#_c_876_n Q 0.0709226f $X=8.96 $Y=2.02 $X2=0 $Y2=0
cc_684 N_A_1507_321#_c_878_n Q 0.00623541f $X=10.19 $Y=1.255 $X2=0 $Y2=0
cc_685 N_A_1507_321#_c_892_n Q 0.0144409f $X=8.817 $Y=2.105 $X2=0 $Y2=0
cc_686 N_A_1507_321#_c_964_p Q 0.0250026f $X=10.24 $Y=1.42 $X2=0 $Y2=0
cc_687 N_A_1507_321#_c_882_n Q 0.0122509f $X=11.2 $Y=1.42 $X2=0 $Y2=0
cc_688 N_A_1507_321#_c_868_n N_VGND_c_1438_n 0.00283345f $X=8.205 $Y=0.78 $X2=0
+ $Y2=0
cc_689 N_A_1507_321#_c_881_n N_VGND_c_1438_n 0.0119053f $X=9.375 $Y=0.495 $X2=0
+ $Y2=0
cc_690 N_A_1507_321#_M1017_g N_VGND_c_1439_n 0.00125495f $X=10.335 $Y=0.845
+ $X2=0 $Y2=0
cc_691 N_A_1507_321#_M1003_g N_VGND_c_1439_n 0.0117336f $X=10.765 $Y=0.845 $X2=0
+ $Y2=0
cc_692 N_A_1507_321#_M1012_g N_VGND_c_1439_n 0.00180891f $X=11.125 $Y=0.845
+ $X2=0 $Y2=0
cc_693 N_A_1507_321#_c_877_n N_VGND_c_1439_n 0.0136299f $X=10.105 $Y=0.35 $X2=0
+ $Y2=0
cc_694 N_A_1507_321#_c_878_n N_VGND_c_1439_n 0.028116f $X=10.19 $Y=1.255 $X2=0
+ $Y2=0
cc_695 N_A_1507_321#_c_879_n N_VGND_c_1439_n 0.0199268f $X=11.6 $Y=1.42 $X2=0
+ $Y2=0
cc_696 N_A_1507_321#_c_882_n N_VGND_c_1439_n 0.00231808f $X=11.2 $Y=1.42 $X2=0
+ $Y2=0
cc_697 N_A_1507_321#_M1012_g N_VGND_c_1440_n 0.00307912f $X=11.125 $Y=0.845
+ $X2=0 $Y2=0
cc_698 N_A_1507_321#_M1017_g N_VGND_c_1443_n 0.00375984f $X=10.335 $Y=0.845
+ $X2=0 $Y2=0
cc_699 N_A_1507_321#_c_877_n N_VGND_c_1443_n 0.0114622f $X=10.105 $Y=0.35 $X2=0
+ $Y2=0
cc_700 N_A_1507_321#_c_881_n N_VGND_c_1443_n 0.0762571f $X=9.375 $Y=0.495 $X2=0
+ $Y2=0
cc_701 N_A_1507_321#_c_868_n N_VGND_c_1447_n 0.00502664f $X=8.205 $Y=0.78 $X2=0
+ $Y2=0
cc_702 N_A_1507_321#_M1003_g N_VGND_c_1448_n 0.00340865f $X=10.765 $Y=0.845
+ $X2=0 $Y2=0
cc_703 N_A_1507_321#_M1012_g N_VGND_c_1448_n 0.00395022f $X=11.125 $Y=0.845
+ $X2=0 $Y2=0
cc_704 N_A_1507_321#_c_868_n N_VGND_c_1450_n 0.0103357f $X=8.205 $Y=0.78 $X2=0
+ $Y2=0
cc_705 N_A_1507_321#_M1017_g N_VGND_c_1450_n 0.00421657f $X=10.335 $Y=0.845
+ $X2=0 $Y2=0
cc_706 N_A_1507_321#_M1003_g N_VGND_c_1450_n 0.00392009f $X=10.765 $Y=0.845
+ $X2=0 $Y2=0
cc_707 N_A_1507_321#_M1012_g N_VGND_c_1450_n 0.00466677f $X=11.125 $Y=0.845
+ $X2=0 $Y2=0
cc_708 N_A_1507_321#_c_877_n N_VGND_c_1450_n 0.00657784f $X=10.105 $Y=0.35 $X2=0
+ $Y2=0
cc_709 N_A_1507_321#_c_881_n N_VGND_c_1450_n 0.0457185f $X=9.375 $Y=0.495 $X2=0
+ $Y2=0
cc_710 N_A_1507_321#_c_868_n N_A_1232_153#_c_1570_n 0.00680366f $X=8.205 $Y=0.78
+ $X2=0 $Y2=0
cc_711 N_A_1507_321#_c_875_n N_A_1232_153#_c_1570_n 0.00567266f $X=8.205
+ $Y=0.855 $X2=0 $Y2=0
cc_712 N_A_1339_153#_M1035_g N_VPWR_c_1185_n 0.0109878f $X=8.49 $Y=2.595 $X2=0
+ $Y2=0
cc_713 N_A_1339_153#_c_1040_n N_VPWR_c_1192_n 0.0177952f $X=6.835 $Y=2.28 $X2=0
+ $Y2=0
cc_714 N_A_1339_153#_M1035_g N_VPWR_c_1193_n 0.00939541f $X=8.49 $Y=2.595 $X2=0
+ $Y2=0
cc_715 N_A_1339_153#_M1023_d N_VPWR_c_1181_n 0.00223819f $X=6.695 $Y=2.095 $X2=0
+ $Y2=0
cc_716 N_A_1339_153#_M1035_g N_VPWR_c_1181_n 0.0181643f $X=8.49 $Y=2.595 $X2=0
+ $Y2=0
cc_717 N_A_1339_153#_c_1040_n N_VPWR_c_1181_n 0.0123247f $X=6.835 $Y=2.28 $X2=0
+ $Y2=0
cc_718 N_A_1339_153#_c_1046_n A_1445_419# 0.0134617f $X=7.445 $Y=2.2 $X2=-0.19
+ $Y2=-0.245
cc_719 N_A_1339_153#_c_1022_n A_1445_419# 2.2849e-19 $X=7.53 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_720 N_A_1339_153#_M1015_g N_Q_c_1390_n 0.00655925f $X=8.995 $Y=0.495 $X2=0
+ $Y2=0
cc_721 N_A_1339_153#_M1035_g Q 0.00171868f $X=8.49 $Y=2.595 $X2=0 $Y2=0
cc_722 N_A_1339_153#_M1015_g Q 0.00485762f $X=8.995 $Y=0.495 $X2=0 $Y2=0
cc_723 N_A_1339_153#_M1024_g N_VGND_c_1438_n 0.0107552f $X=8.635 $Y=0.495 $X2=0
+ $Y2=0
cc_724 N_A_1339_153#_M1015_g N_VGND_c_1438_n 0.00130258f $X=8.995 $Y=0.495 $X2=0
+ $Y2=0
cc_725 N_A_1339_153#_c_1019_n N_VGND_c_1438_n 0.00133367f $X=8.537 $Y=1.245
+ $X2=0 $Y2=0
cc_726 N_A_1339_153#_c_1023_n N_VGND_c_1438_n 0.00107951f $X=8.365 $Y=1.35 $X2=0
+ $Y2=0
cc_727 N_A_1339_153#_c_1025_n N_VGND_c_1438_n 0.00935245f $X=8.53 $Y=1.335 $X2=0
+ $Y2=0
cc_728 N_A_1339_153#_M1024_g N_VGND_c_1443_n 0.00445056f $X=8.635 $Y=0.495 $X2=0
+ $Y2=0
cc_729 N_A_1339_153#_M1015_g N_VGND_c_1443_n 0.00327726f $X=8.995 $Y=0.495 $X2=0
+ $Y2=0
cc_730 N_A_1339_153#_M1024_g N_VGND_c_1450_n 0.00796275f $X=8.635 $Y=0.495 $X2=0
+ $Y2=0
cc_731 N_A_1339_153#_M1015_g N_VGND_c_1450_n 0.00563495f $X=8.995 $Y=0.495 $X2=0
+ $Y2=0
cc_732 N_A_1339_153#_c_1023_n N_A_1232_153#_c_1570_n 0.0113008f $X=8.365 $Y=1.35
+ $X2=0 $Y2=0
cc_733 N_A_2062_367#_c_1129_n N_VPWR_c_1186_n 0.0605865f $X=10.45 $Y=1.98 $X2=0
+ $Y2=0
cc_734 N_A_2062_367#_c_1131_n N_VPWR_c_1186_n 0.00840433f $X=10.615 $Y=1.85
+ $X2=0 $Y2=0
cc_735 N_A_2062_367#_c_1127_n N_VPWR_c_1187_n 0.0276659f $X=12.415 $Y=2.01 $X2=0
+ $Y2=0
cc_736 N_A_2062_367#_c_1128_n N_VPWR_c_1187_n 0.00178319f $X=12.222 $Y=1.668
+ $X2=0 $Y2=0
cc_737 N_A_2062_367#_c_1130_n N_VPWR_c_1187_n 0.0261206f $X=12.005 $Y=1.85 $X2=0
+ $Y2=0
cc_738 N_A_2062_367#_c_1129_n N_VPWR_c_1188_n 0.00963752f $X=10.45 $Y=1.98 $X2=0
+ $Y2=0
cc_739 N_A_2062_367#_c_1127_n N_VPWR_c_1194_n 0.00769046f $X=12.415 $Y=2.01
+ $X2=0 $Y2=0
cc_740 N_A_2062_367#_c_1127_n N_VPWR_c_1181_n 0.014085f $X=12.415 $Y=2.01 $X2=0
+ $Y2=0
cc_741 N_A_2062_367#_c_1129_n N_VPWR_c_1181_n 0.0111417f $X=10.45 $Y=1.98 $X2=0
+ $Y2=0
cc_742 N_A_2062_367#_M1032_g Q_N 0.0029356f $X=12.105 $Y=0.495 $X2=0 $Y2=0
cc_743 N_A_2062_367#_c_1127_n Q_N 0.0225057f $X=12.415 $Y=2.01 $X2=0 $Y2=0
cc_744 N_A_2062_367#_M1025_g Q_N 0.0261786f $X=12.465 $Y=0.495 $X2=0 $Y2=0
cc_745 N_A_2062_367#_c_1121_n Q_N 0.00598623f $X=12.272 $Y=1.365 $X2=0 $Y2=0
cc_746 N_A_2062_367#_c_1128_n Q_N 0.00715128f $X=12.222 $Y=1.668 $X2=0 $Y2=0
cc_747 N_A_2062_367#_c_1130_n Q_N 0.0134526f $X=12.005 $Y=1.85 $X2=0 $Y2=0
cc_748 N_A_2062_367#_c_1122_n Q_N 0.00775774f $X=12.005 $Y=0.99 $X2=0 $Y2=0
cc_749 N_A_2062_367#_c_1123_n Q_N 0.0409299f $X=12.17 $Y=1.38 $X2=0 $Y2=0
cc_750 N_A_2062_367#_c_1124_n Q_N 0.0140734f $X=12.17 $Y=1.38 $X2=0 $Y2=0
cc_751 N_A_2062_367#_c_1126_n Q_N 0.00567519f $X=12.17 $Y=1.215 $X2=0 $Y2=0
cc_752 N_A_2062_367#_c_1125_n N_VGND_c_1439_n 0.0150699f $X=11.34 $Y=0.845 $X2=0
+ $Y2=0
cc_753 N_A_2062_367#_M1032_g N_VGND_c_1440_n 0.0140665f $X=12.105 $Y=0.495 $X2=0
+ $Y2=0
cc_754 N_A_2062_367#_M1025_g N_VGND_c_1440_n 0.002112f $X=12.465 $Y=0.495 $X2=0
+ $Y2=0
cc_755 N_A_2062_367#_c_1122_n N_VGND_c_1440_n 0.0267804f $X=12.005 $Y=0.99 $X2=0
+ $Y2=0
cc_756 N_A_2062_367#_c_1125_n N_VGND_c_1440_n 0.00764783f $X=11.34 $Y=0.845
+ $X2=0 $Y2=0
cc_757 N_A_2062_367#_c_1125_n N_VGND_c_1448_n 0.00667264f $X=11.34 $Y=0.845
+ $X2=0 $Y2=0
cc_758 N_A_2062_367#_M1032_g N_VGND_c_1449_n 0.00445056f $X=12.105 $Y=0.495
+ $X2=0 $Y2=0
cc_759 N_A_2062_367#_M1025_g N_VGND_c_1449_n 0.00502664f $X=12.465 $Y=0.495
+ $X2=0 $Y2=0
cc_760 N_A_2062_367#_M1032_g N_VGND_c_1450_n 0.00796275f $X=12.105 $Y=0.495
+ $X2=0 $Y2=0
cc_761 N_A_2062_367#_M1025_g N_VGND_c_1450_n 0.0100616f $X=12.465 $Y=0.495 $X2=0
+ $Y2=0
cc_762 N_A_2062_367#_c_1125_n N_VGND_c_1450_n 0.00989637f $X=11.34 $Y=0.845
+ $X2=0 $Y2=0
cc_763 N_VPWR_c_1183_n N_A_349_323#_c_1354_n 0.0224958f $X=4.03 $Y=2.15 $X2=0
+ $Y2=0
cc_764 N_VPWR_c_1190_n N_A_349_323#_c_1354_n 0.0210163f $X=3.865 $Y=3.33 $X2=0
+ $Y2=0
cc_765 N_VPWR_c_1181_n N_A_349_323#_c_1354_n 0.00912687f $X=12.72 $Y=3.33 $X2=0
+ $Y2=0
cc_766 N_VPWR_c_1183_n N_A_349_323#_c_1355_n 0.028959f $X=4.03 $Y=2.15 $X2=0
+ $Y2=0
cc_767 N_VPWR_c_1181_n N_A_349_323#_c_1356_n 0.0236949f $X=12.72 $Y=3.33 $X2=0
+ $Y2=0
cc_768 N_VPWR_c_1181_n A_1445_419# 0.0132771f $X=12.72 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_769 N_VPWR_c_1186_n Q 0.0708325f $X=9.92 $Y=1.98 $X2=0 $Y2=0
cc_770 N_VPWR_c_1193_n Q 0.0106618f $X=9.755 $Y=3.33 $X2=0 $Y2=0
cc_771 N_VPWR_c_1181_n Q 0.0114128f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_772 N_VPWR_c_1187_n Q_N 0.0625962f $X=12.15 $Y=2.28 $X2=0 $Y2=0
cc_773 N_VPWR_c_1194_n Q_N 0.0220321f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_774 N_VPWR_c_1181_n Q_N 0.0125808f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_775 N_A_239_403#_c_1303_n N_A_349_323#_M1026_s 0.00431926f $X=1.82 $Y=2.12
+ $X2=-0.19 $Y2=-0.245
cc_776 N_A_239_403#_c_1301_n N_A_349_323#_M1026_s 0.008656f $X=1.905 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_777 N_A_239_403#_c_1343_p N_A_349_323#_M1026_s 0.00190582f $X=1.905 $Y=2.12
+ $X2=-0.19 $Y2=-0.245
cc_778 N_A_239_403#_M1008_d N_A_349_323#_c_1354_n 0.00706692f $X=2.805 $Y=1.615
+ $X2=0 $Y2=0
cc_779 N_A_239_403#_c_1306_n N_A_349_323#_c_1354_n 0.0195261f $X=2.945 $Y=2.075
+ $X2=0 $Y2=0
cc_780 N_A_239_403#_c_1323_n N_A_349_323#_c_1354_n 0.0347295f $X=2.78 $Y=2.115
+ $X2=0 $Y2=0
cc_781 N_A_239_403#_c_1306_n N_A_349_323#_c_1355_n 0.018394f $X=2.945 $Y=2.075
+ $X2=0 $Y2=0
cc_782 N_A_239_403#_c_1303_n N_A_349_323#_c_1356_n 0.00710777f $X=1.82 $Y=2.12
+ $X2=0 $Y2=0
cc_783 N_A_239_403#_c_1343_p N_A_349_323#_c_1356_n 0.0116606f $X=1.905 $Y=2.12
+ $X2=0 $Y2=0
cc_784 N_A_239_403#_c_1323_n N_A_349_323#_c_1356_n 0.00161189f $X=2.78 $Y=2.115
+ $X2=0 $Y2=0
cc_785 N_A_239_403#_c_1302_n N_VGND_c_1435_n 0.0150699f $X=1.985 $Y=0.635 $X2=0
+ $Y2=0
cc_786 N_A_239_403#_c_1302_n N_VGND_c_1446_n 0.0116898f $X=1.985 $Y=0.635 $X2=0
+ $Y2=0
cc_787 N_A_239_403#_c_1302_n N_VGND_c_1450_n 0.01158f $X=1.985 $Y=0.635 $X2=0
+ $Y2=0
cc_788 Q_N N_VGND_c_1440_n 0.0153904f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_789 Q_N N_VGND_c_1449_n 0.0220321f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_790 Q_N N_VGND_c_1450_n 0.0125808f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_791 N_VGND_c_1437_n N_A_1232_153#_c_1567_n 0.0406934f $X=5.745 $Y=0.835 $X2=0
+ $Y2=0
cc_792 N_VGND_c_1447_n N_A_1232_153#_c_1568_n 0.0865384f $X=8.335 $Y=0 $X2=0
+ $Y2=0
cc_793 N_VGND_c_1450_n N_A_1232_153#_c_1568_n 0.0498987f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_794 N_VGND_c_1437_n N_A_1232_153#_c_1569_n 0.0119254f $X=5.745 $Y=0.835 $X2=0
+ $Y2=0
cc_795 N_VGND_c_1447_n N_A_1232_153#_c_1569_n 0.0168491f $X=8.335 $Y=0 $X2=0
+ $Y2=0
cc_796 N_VGND_c_1450_n N_A_1232_153#_c_1569_n 0.00867615f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_797 N_VGND_c_1438_n N_A_1232_153#_c_1570_n 0.0179429f $X=8.42 $Y=0.495 $X2=0
+ $Y2=0
cc_798 N_VGND_c_1447_n N_A_1232_153#_c_1570_n 0.0214013f $X=8.335 $Y=0 $X2=0
+ $Y2=0
cc_799 N_VGND_c_1450_n N_A_1232_153#_c_1570_n 0.0124501f $X=12.72 $Y=0 $X2=0
+ $Y2=0
