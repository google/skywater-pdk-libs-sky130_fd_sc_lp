* File: sky130_fd_sc_lp__or4_m.pxi.spice
* Created: Wed Sep  2 10:32:19 2020
* 
x_PM_SKY130_FD_SC_LP__OR4_M%D N_D_c_72_n N_D_M1006_g N_D_M1003_g N_D_c_68_n
+ N_D_c_69_n D D D D D N_D_c_71_n PM_SKY130_FD_SC_LP__OR4_M%D
x_PM_SKY130_FD_SC_LP__OR4_M%C N_C_M1009_g N_C_c_98_n N_C_M1002_g N_C_c_100_n C C
+ C N_C_c_102_n N_C_c_103_n PM_SKY130_FD_SC_LP__OR4_M%C
x_PM_SKY130_FD_SC_LP__OR4_M%B N_B_c_137_n N_B_M1005_g N_B_M1001_g N_B_c_139_n B
+ B N_B_c_140_n N_B_c_141_n PM_SKY130_FD_SC_LP__OR4_M%B
x_PM_SKY130_FD_SC_LP__OR4_M%A N_A_c_176_n N_A_M1000_g N_A_M1007_g N_A_c_178_n A
+ N_A_c_179_n N_A_c_180_n PM_SKY130_FD_SC_LP__OR4_M%A
x_PM_SKY130_FD_SC_LP__OR4_M%A_116_397# N_A_116_397#_M1006_d N_A_116_397#_M1001_d
+ N_A_116_397#_M1003_s N_A_116_397#_c_226_n N_A_116_397#_M1008_g
+ N_A_116_397#_M1004_g N_A_116_397#_c_229_n N_A_116_397#_c_222_n
+ N_A_116_397#_c_231_n N_A_116_397#_c_232_n N_A_116_397#_c_267_n
+ N_A_116_397#_c_233_n N_A_116_397#_c_223_n N_A_116_397#_c_224_n
+ N_A_116_397#_c_225_n N_A_116_397#_c_235_n N_A_116_397#_c_236_n
+ N_A_116_397#_c_237_n PM_SKY130_FD_SC_LP__OR4_M%A_116_397#
x_PM_SKY130_FD_SC_LP__OR4_M%VPWR N_VPWR_M1000_d N_VPWR_c_323_n N_VPWR_c_324_n
+ N_VPWR_c_325_n VPWR N_VPWR_c_326_n N_VPWR_c_322_n
+ PM_SKY130_FD_SC_LP__OR4_M%VPWR
x_PM_SKY130_FD_SC_LP__OR4_M%X N_X_M1004_d N_X_M1008_d X X X X X X X N_X_c_351_n
+ N_X_c_349_n PM_SKY130_FD_SC_LP__OR4_M%X
x_PM_SKY130_FD_SC_LP__OR4_M%VGND N_VGND_M1006_s N_VGND_M1009_d N_VGND_M1007_d
+ N_VGND_c_368_n N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n VGND
+ N_VGND_c_372_n N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n
+ N_VGND_c_377_n PM_SKY130_FD_SC_LP__OR4_M%VGND
cc_1 VNB N_D_M1006_g 0.0341706f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.445
cc_2 VNB N_D_c_68_n 0.042058f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.03
cc_3 VNB N_D_c_69_n 0.0254814f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_4 VNB D 0.00894729f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_D_c_71_n 0.0380391f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_6 VNB N_C_c_98_n 0.0230131f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.445
cc_7 VNB N_C_M1002_g 0.0123235f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.195
cc_8 VNB N_C_c_100_n 0.0220655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB C 0.00266071f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.03
cc_10 VNB N_C_c_102_n 0.0212163f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_11 VNB N_C_c_103_n 0.0183683f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_B_c_137_n 0.0222884f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.75
cc_13 VNB N_B_M1005_g 0.012284f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.445
cc_14 VNB N_B_c_139_n 0.0186715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_140_n 0.0187751f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_16 VNB N_B_c_141_n 0.0187895f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_17 VNB N_A_c_176_n 0.021425f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=1.75
cc_18 VNB N_A_M1007_g 0.0253617f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.825
cc_19 VNB N_A_c_178_n 0.0206698f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.03
cc_20 VNB N_A_c_179_n 0.0156217f $X=-0.19 $Y=-0.245 $X2=0.285 $Y2=1.75
cc_21 VNB N_A_c_180_n 0.0081988f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_22 VNB N_A_116_397#_M1004_g 0.0729245f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_23 VNB N_A_116_397#_c_222_n 0.0218527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_116_397#_c_223_n 0.00850046f $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=2.405
cc_25 VNB N_A_116_397#_c_224_n 0.00644118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_116_397#_c_225_n 0.0162019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_322_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_28 VNB X 0.0572869f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.825
cc_29 VNB N_X_c_349_n 0.00765173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_368_n 0.014599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_369_n 0.012755f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_32 VNB N_VGND_c_370_n 0.00277226f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_33 VNB N_VGND_c_371_n 0.00505305f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_34 VNB N_VGND_c_372_n 0.0252661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_373_n 0.0159754f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_36 VNB N_VGND_c_374_n 0.0182237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_375_n 0.191405f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_38 VNB N_VGND_c_376_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_377_n 0.00631443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_D_c_72_n 0.0427047f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.75
cc_41 VPB N_D_M1003_g 0.0238008f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.195
cc_42 VPB N_D_c_69_n 0.0140042f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_43 VPB D 0.043384f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_44 VPB N_C_M1002_g 0.0266933f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.195
cc_45 VPB N_B_M1005_g 0.0266783f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.445
cc_46 VPB N_A_c_176_n 0.0281613f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.75
cc_47 VPB N_A_M1000_g 0.0155585f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.955
cc_48 VPB N_A_116_397#_c_226_n 0.0573297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_116_397#_M1008_g 0.031848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_116_397#_M1004_g 0.00437116f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_51 VPB N_A_116_397#_c_229_n 0.0187684f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_52 VPB N_A_116_397#_c_222_n 4.66948e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_116_397#_c_231_n 0.0263163f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_54 VPB N_A_116_397#_c_232_n 0.0134867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_116_397#_c_233_n 0.0189889f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=2.035
cc_56 VPB N_A_116_397#_c_225_n 0.00200666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_116_397#_c_235_n 0.00341723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_116_397#_c_236_n 0.00166901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_116_397#_c_237_n 0.0512764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_323_n 0.0205886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_324_n 0.0720326f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.195
cc_62 VPB N_VPWR_c_325_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_326_n 0.0229627f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_64 VPB N_VPWR_c_322_n 0.108354f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_65 VPB X 0.0239087f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=1.825
cc_66 VPB N_X_c_351_n 0.0381681f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_67 N_D_c_71_n N_C_c_98_n 0.00363253f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_68 N_D_c_72_n N_C_M1002_g 0.0552013f $X=0.845 $Y=1.75 $X2=0 $Y2=0
cc_69 N_D_c_72_n N_C_c_100_n 0.00101511f $X=0.845 $Y=1.75 $X2=0 $Y2=0
cc_70 N_D_c_68_n N_C_c_102_n 0.0136966f $X=0.625 $Y=1.03 $X2=0 $Y2=0
cc_71 N_D_M1006_g N_C_c_103_n 0.0136966f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_72 N_D_c_72_n N_A_116_397#_c_222_n 0.010805f $X=0.845 $Y=1.75 $X2=0 $Y2=0
cc_73 N_D_M1006_g N_A_116_397#_c_222_n 0.00760501f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_74 D N_A_116_397#_c_222_n 0.0382329f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_75 N_D_c_71_n N_A_116_397#_c_222_n 0.00537249f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_76 N_D_c_72_n N_A_116_397#_c_231_n 0.00272308f $X=0.845 $Y=1.75 $X2=0 $Y2=0
cc_77 N_D_M1003_g N_A_116_397#_c_231_n 0.00504921f $X=0.92 $Y=2.195 $X2=0 $Y2=0
cc_78 N_D_c_72_n N_A_116_397#_c_235_n 0.00881941f $X=0.845 $Y=1.75 $X2=0 $Y2=0
cc_79 N_D_M1003_g N_A_116_397#_c_235_n 0.0139932f $X=0.92 $Y=2.195 $X2=0 $Y2=0
cc_80 D N_A_116_397#_c_235_n 0.0280099f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_81 N_D_M1003_g N_VPWR_c_322_n 0.00393927f $X=0.92 $Y=2.195 $X2=0 $Y2=0
cc_82 D N_VPWR_c_322_n 0.00780715f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_83 N_D_M1006_g N_VGND_c_369_n 0.00837342f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_84 N_D_c_68_n N_VGND_c_369_n 0.00589231f $X=0.625 $Y=1.03 $X2=0 $Y2=0
cc_85 D N_VGND_c_369_n 0.00607684f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_86 N_D_M1006_g N_VGND_c_372_n 0.00564095f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_87 N_D_M1006_g N_VGND_c_375_n 0.00961799f $X=0.625 $Y=0.445 $X2=0 $Y2=0
cc_88 D N_VGND_c_375_n 0.00345756f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_C_c_98_n N_B_c_137_n 0.0278477f $X=1.167 $Y=1.248 $X2=0 $Y2=0
cc_90 N_C_M1002_g N_B_M1005_g 0.0278477f $X=1.28 $Y=2.195 $X2=0 $Y2=0
cc_91 N_C_c_100_n N_B_c_139_n 0.0278477f $X=1.167 $Y=1.435 $X2=0 $Y2=0
cc_92 C B 0.0258924f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_93 N_C_c_102_n B 0.00202054f $X=1.19 $Y=0.93 $X2=0 $Y2=0
cc_94 C N_B_c_140_n 0.00251455f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_95 N_C_c_102_n N_B_c_140_n 0.0278477f $X=1.19 $Y=0.93 $X2=0 $Y2=0
cc_96 C N_B_c_141_n 0.00426692f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_97 N_C_c_103_n N_B_c_141_n 0.00617639f $X=1.167 $Y=0.765 $X2=0 $Y2=0
cc_98 N_C_M1002_g N_A_116_397#_c_222_n 0.00806445f $X=1.28 $Y=2.195 $X2=0 $Y2=0
cc_99 C N_A_116_397#_c_222_n 0.0600463f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_100 N_C_c_103_n N_A_116_397#_c_222_n 0.00884272f $X=1.167 $Y=0.765 $X2=0
+ $Y2=0
cc_101 N_C_M1002_g N_A_116_397#_c_231_n 0.0164902f $X=1.28 $Y=2.195 $X2=0 $Y2=0
cc_102 N_C_c_100_n N_A_116_397#_c_231_n 0.00444163f $X=1.167 $Y=1.435 $X2=0
+ $Y2=0
cc_103 C N_A_116_397#_c_231_n 0.00778616f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_104 N_C_M1002_g N_A_116_397#_c_235_n 0.00178724f $X=1.28 $Y=2.195 $X2=0 $Y2=0
cc_105 N_C_M1002_g N_VPWR_c_322_n 0.00393927f $X=1.28 $Y=2.195 $X2=0 $Y2=0
cc_106 C N_VGND_M1009_d 0.00416057f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_107 N_C_c_103_n N_VGND_c_369_n 0.00148579f $X=1.167 $Y=0.765 $X2=0 $Y2=0
cc_108 C N_VGND_c_370_n 0.00110313f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_109 N_C_c_103_n N_VGND_c_370_n 0.00555936f $X=1.167 $Y=0.765 $X2=0 $Y2=0
cc_110 C N_VGND_c_372_n 0.00434621f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_111 N_C_c_102_n N_VGND_c_372_n 0.00182358f $X=1.19 $Y=0.93 $X2=0 $Y2=0
cc_112 N_C_c_103_n N_VGND_c_372_n 0.00555499f $X=1.167 $Y=0.765 $X2=0 $Y2=0
cc_113 C N_VGND_c_375_n 0.0059602f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_114 N_C_c_102_n N_VGND_c_375_n 0.00189735f $X=1.19 $Y=0.93 $X2=0 $Y2=0
cc_115 N_C_c_103_n N_VGND_c_375_n 0.0108748f $X=1.167 $Y=0.765 $X2=0 $Y2=0
cc_116 N_B_M1005_g N_A_c_176_n 0.0604479f $X=1.64 $Y=2.195 $X2=-0.19 $Y2=-0.245
cc_117 N_B_c_139_n N_A_c_176_n 0.0108707f $X=1.742 $Y=1.435 $X2=-0.19 $Y2=-0.245
cc_118 B N_A_M1007_g 4.72661e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_119 N_B_c_141_n N_A_M1007_g 0.0210357f $X=1.742 $Y=0.765 $X2=0 $Y2=0
cc_120 N_B_c_137_n N_A_c_178_n 0.0108707f $X=1.742 $Y=1.258 $X2=0 $Y2=0
cc_121 B N_A_c_179_n 9.45757e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_122 N_B_c_140_n N_A_c_179_n 0.0108707f $X=1.73 $Y=0.93 $X2=0 $Y2=0
cc_123 N_B_c_137_n N_A_c_180_n 0.00365974f $X=1.742 $Y=1.258 $X2=0 $Y2=0
cc_124 N_B_M1005_g N_A_c_180_n 0.00151122f $X=1.64 $Y=2.195 $X2=0 $Y2=0
cc_125 B N_A_c_180_n 0.0291874f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_126 N_B_M1005_g N_A_116_397#_c_231_n 0.0150473f $X=1.64 $Y=2.195 $X2=0 $Y2=0
cc_127 N_B_c_139_n N_A_116_397#_c_231_n 0.00136881f $X=1.742 $Y=1.435 $X2=0
+ $Y2=0
cc_128 B N_A_116_397#_c_231_n 0.00778745f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_129 N_B_M1005_g N_A_116_397#_c_232_n 0.0147918f $X=1.64 $Y=2.195 $X2=0 $Y2=0
cc_130 N_B_c_141_n N_A_116_397#_c_224_n 0.00465408f $X=1.742 $Y=0.765 $X2=0
+ $Y2=0
cc_131 N_B_c_139_n N_A_116_397#_c_236_n 0.00394702f $X=1.742 $Y=1.435 $X2=0
+ $Y2=0
cc_132 B N_A_116_397#_c_236_n 0.00534404f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_133 N_B_M1005_g N_VPWR_c_322_n 0.00393927f $X=1.64 $Y=2.195 $X2=0 $Y2=0
cc_134 B N_VGND_c_370_n 0.0081944f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_135 N_B_c_140_n N_VGND_c_370_n 0.00507809f $X=1.73 $Y=0.93 $X2=0 $Y2=0
cc_136 N_B_c_141_n N_VGND_c_370_n 0.00829521f $X=1.742 $Y=0.765 $X2=0 $Y2=0
cc_137 N_B_c_141_n N_VGND_c_373_n 0.00486043f $X=1.742 $Y=0.765 $X2=0 $Y2=0
cc_138 B N_VGND_c_375_n 0.00414189f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_139 N_B_c_141_n N_VGND_c_375_n 0.00541582f $X=1.742 $Y=0.765 $X2=0 $Y2=0
cc_140 N_A_c_176_n N_A_116_397#_M1004_g 0.00197361f $X=2 $Y=1.825 $X2=0 $Y2=0
cc_141 N_A_M1007_g N_A_116_397#_M1004_g 0.0173131f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_c_179_n N_A_116_397#_M1004_g 0.0193418f $X=2.295 $Y=1.085 $X2=0 $Y2=0
cc_143 N_A_c_176_n N_A_116_397#_c_229_n 0.00288634f $X=2 $Y=1.825 $X2=0 $Y2=0
cc_144 N_A_M1000_g N_A_116_397#_c_229_n 0.00932369f $X=2 $Y=2.195 $X2=0 $Y2=0
cc_145 N_A_M1000_g N_A_116_397#_c_232_n 0.0181378f $X=2 $Y=2.195 $X2=0 $Y2=0
cc_146 N_A_M1007_g N_A_116_397#_c_267_n 0.00617227f $X=2.275 $Y=0.445 $X2=0
+ $Y2=0
cc_147 N_A_c_176_n N_A_116_397#_c_233_n 0.0116195f $X=2 $Y=1.825 $X2=0 $Y2=0
cc_148 N_A_c_180_n N_A_116_397#_c_233_n 0.0181627f $X=2.295 $Y=1.085 $X2=0 $Y2=0
cc_149 N_A_M1007_g N_A_116_397#_c_223_n 0.00834497f $X=2.275 $Y=0.445 $X2=0
+ $Y2=0
cc_150 N_A_c_179_n N_A_116_397#_c_223_n 0.00311486f $X=2.295 $Y=1.085 $X2=0
+ $Y2=0
cc_151 N_A_c_180_n N_A_116_397#_c_223_n 0.0155783f $X=2.295 $Y=1.085 $X2=0 $Y2=0
cc_152 N_A_M1007_g N_A_116_397#_c_224_n 0.00245333f $X=2.275 $Y=0.445 $X2=0
+ $Y2=0
cc_153 N_A_c_179_n N_A_116_397#_c_224_n 0.00206478f $X=2.295 $Y=1.085 $X2=0
+ $Y2=0
cc_154 N_A_c_180_n N_A_116_397#_c_224_n 0.0138362f $X=2.295 $Y=1.085 $X2=0 $Y2=0
cc_155 N_A_c_176_n N_A_116_397#_c_225_n 0.00553186f $X=2 $Y=1.825 $X2=0 $Y2=0
cc_156 N_A_M1007_g N_A_116_397#_c_225_n 0.00191687f $X=2.275 $Y=0.445 $X2=0
+ $Y2=0
cc_157 N_A_c_179_n N_A_116_397#_c_225_n 0.00349021f $X=2.295 $Y=1.085 $X2=0
+ $Y2=0
cc_158 N_A_c_180_n N_A_116_397#_c_225_n 0.0371014f $X=2.295 $Y=1.085 $X2=0 $Y2=0
cc_159 N_A_c_176_n N_A_116_397#_c_236_n 0.00855445f $X=2 $Y=1.825 $X2=0 $Y2=0
cc_160 N_A_M1000_g N_A_116_397#_c_236_n 0.0058826f $X=2 $Y=2.195 $X2=0 $Y2=0
cc_161 N_A_c_180_n N_A_116_397#_c_236_n 0.00176724f $X=2.295 $Y=1.085 $X2=0
+ $Y2=0
cc_162 N_A_M1000_g N_A_116_397#_c_237_n 0.00828381f $X=2 $Y=2.195 $X2=0 $Y2=0
cc_163 N_A_M1000_g N_VPWR_c_323_n 0.00154866f $X=2 $Y=2.195 $X2=0 $Y2=0
cc_164 N_A_M1007_g N_VGND_c_370_n 6.90856e-19 $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_M1007_g N_VGND_c_371_n 0.00436717f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A_M1007_g N_VGND_c_373_n 0.00412386f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A_M1007_g N_VGND_c_375_n 0.00626145f $X=2.275 $Y=0.445 $X2=0 $Y2=0
cc_168 N_A_116_397#_c_232_n A_343_397# 0.00500535f $X=1.94 $Y=2.94 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_116_397#_c_226_n N_VPWR_c_323_n 0.0258133f $X=2.67 $Y=2.85 $X2=0
+ $Y2=0
cc_170 N_A_116_397#_M1008_g N_VPWR_c_323_n 0.00881892f $X=2.745 $Y=2.195 $X2=0
+ $Y2=0
cc_171 N_A_116_397#_c_232_n N_VPWR_c_323_n 0.0574939f $X=1.94 $Y=2.94 $X2=0
+ $Y2=0
cc_172 N_A_116_397#_c_233_n N_VPWR_c_323_n 0.0249693f $X=2.64 $Y=1.88 $X2=0
+ $Y2=0
cc_173 N_A_116_397#_c_237_n N_VPWR_c_323_n 0.00524695f $X=1.94 $Y=2.85 $X2=0
+ $Y2=0
cc_174 N_A_116_397#_c_226_n N_VPWR_c_324_n 0.00445258f $X=2.67 $Y=2.85 $X2=0
+ $Y2=0
cc_175 N_A_116_397#_c_232_n N_VPWR_c_324_n 0.0167839f $X=1.94 $Y=2.94 $X2=0
+ $Y2=0
cc_176 N_A_116_397#_c_237_n N_VPWR_c_324_n 0.0059602f $X=1.94 $Y=2.85 $X2=0
+ $Y2=0
cc_177 N_A_116_397#_c_226_n N_VPWR_c_326_n 0.00581074f $X=2.67 $Y=2.85 $X2=0
+ $Y2=0
cc_178 N_A_116_397#_c_226_n N_VPWR_c_322_n 0.0111595f $X=2.67 $Y=2.85 $X2=0
+ $Y2=0
cc_179 N_A_116_397#_c_232_n N_VPWR_c_322_n 0.0108843f $X=1.94 $Y=2.94 $X2=0
+ $Y2=0
cc_180 N_A_116_397#_c_237_n N_VPWR_c_322_n 0.00813556f $X=1.94 $Y=2.85 $X2=0
+ $Y2=0
cc_181 N_A_116_397#_M1008_g X 0.00663958f $X=2.745 $Y=2.195 $X2=0 $Y2=0
cc_182 N_A_116_397#_M1004_g X 0.0329025f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_183 N_A_116_397#_c_233_n X 0.011204f $X=2.64 $Y=1.88 $X2=0 $Y2=0
cc_184 N_A_116_397#_c_223_n X 0.0112285f $X=2.64 $Y=0.735 $X2=0 $Y2=0
cc_185 N_A_116_397#_c_225_n X 0.0613643f $X=2.725 $Y=1.795 $X2=0 $Y2=0
cc_186 N_A_116_397#_c_226_n N_X_c_351_n 0.00359118f $X=2.67 $Y=2.85 $X2=0 $Y2=0
cc_187 N_A_116_397#_M1008_g N_X_c_351_n 0.0155624f $X=2.745 $Y=2.195 $X2=0 $Y2=0
cc_188 N_A_116_397#_c_229_n N_X_c_351_n 0.00478711f $X=2.885 $Y=1.8 $X2=0 $Y2=0
cc_189 N_A_116_397#_c_233_n N_X_c_351_n 0.00108594f $X=2.64 $Y=1.88 $X2=0 $Y2=0
cc_190 N_A_116_397#_M1004_g N_X_c_349_n 0.00332088f $X=2.885 $Y=0.445 $X2=0
+ $Y2=0
cc_191 N_A_116_397#_c_223_n N_VGND_M1007_d 0.00387987f $X=2.64 $Y=0.735 $X2=0
+ $Y2=0
cc_192 N_A_116_397#_M1004_g N_VGND_c_371_n 0.00462294f $X=2.885 $Y=0.445 $X2=0
+ $Y2=0
cc_193 N_A_116_397#_c_267_n N_VGND_c_371_n 0.00988056f $X=2.06 $Y=0.495 $X2=0
+ $Y2=0
cc_194 N_A_116_397#_c_223_n N_VGND_c_371_n 0.0240305f $X=2.64 $Y=0.735 $X2=0
+ $Y2=0
cc_195 N_A_116_397#_c_222_n N_VGND_c_372_n 0.00787177f $X=0.84 $Y=0.51 $X2=0
+ $Y2=0
cc_196 N_A_116_397#_c_267_n N_VGND_c_373_n 0.0109202f $X=2.06 $Y=0.495 $X2=0
+ $Y2=0
cc_197 N_A_116_397#_c_223_n N_VGND_c_373_n 0.00248107f $X=2.64 $Y=0.735 $X2=0
+ $Y2=0
cc_198 N_A_116_397#_M1004_g N_VGND_c_374_n 0.0054978f $X=2.885 $Y=0.445 $X2=0
+ $Y2=0
cc_199 N_A_116_397#_M1006_d N_VGND_c_375_n 0.00550887f $X=0.7 $Y=0.235 $X2=0
+ $Y2=0
cc_200 N_A_116_397#_M1001_d N_VGND_c_375_n 0.00424877f $X=1.92 $Y=0.235 $X2=0
+ $Y2=0
cc_201 N_A_116_397#_M1004_g N_VGND_c_375_n 0.0112627f $X=2.885 $Y=0.445 $X2=0
+ $Y2=0
cc_202 N_A_116_397#_c_222_n N_VGND_c_375_n 0.0069578f $X=0.84 $Y=0.51 $X2=0
+ $Y2=0
cc_203 N_A_116_397#_c_267_n N_VGND_c_375_n 0.00964148f $X=2.06 $Y=0.495 $X2=0
+ $Y2=0
cc_204 N_A_116_397#_c_223_n N_VGND_c_375_n 0.00779863f $X=2.64 $Y=0.735 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_323_n N_X_c_351_n 0.0444262f $X=2.45 $Y=2.26 $X2=0 $Y2=0
cc_206 N_VPWR_c_326_n N_X_c_351_n 0.0139886f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_207 N_VPWR_c_322_n N_X_c_351_n 0.0159751f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_208 N_X_c_349_n N_VGND_c_374_n 0.0179455f $X=3.1 $Y=0.385 $X2=0 $Y2=0
cc_209 N_X_M1004_d N_VGND_c_375_n 0.00216084f $X=2.96 $Y=0.235 $X2=0 $Y2=0
cc_210 N_X_c_349_n N_VGND_c_375_n 0.0122929f $X=3.1 $Y=0.385 $X2=0 $Y2=0
