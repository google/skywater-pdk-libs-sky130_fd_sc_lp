# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dfstp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.855000 1.835000 2.190000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.095000 0.255000 10.475000 1.095000 ;
        RECT 10.205000 1.095000 10.475000 3.075000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.090000 1.765000 7.605000 1.915000 ;
        RECT 4.090000 1.915000 6.055000 1.935000 ;
        RECT 4.090000 1.935000 4.300000 2.155000 ;
        RECT 4.270000 0.845000 4.805000 1.095000 ;
        RECT 4.270000 1.095000 4.440000 1.765000 ;
        RECT 5.885000 1.245000 7.605000 1.765000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.440000 0.840000 0.875000 1.390000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.245000 10.560000 3.415000 ;
      RECT 0.090000  0.390000  0.495000 0.670000 ;
      RECT 0.090000  0.670000  0.260000 1.560000 ;
      RECT 0.090000  1.560000  0.865000 1.810000 ;
      RECT 0.090000  1.810000  0.395000 2.965000 ;
      RECT 0.565000  2.305000  0.875000 3.245000 ;
      RECT 0.665000  0.085000  0.865000 0.670000 ;
      RECT 1.045000  0.410000  1.355000 1.515000 ;
      RECT 1.045000  1.515000  2.235000 1.685000 ;
      RECT 1.045000  1.685000  1.255000 2.965000 ;
      RECT 1.545000  0.085000  1.845000 0.970000 ;
      RECT 1.595000  2.360000  1.895000 3.245000 ;
      RECT 2.005000  1.685000  2.235000 1.845000 ;
      RECT 2.015000  0.640000  2.235000 1.175000 ;
      RECT 2.015000  1.175000  2.575000 1.345000 ;
      RECT 2.065000  2.015000  2.575000 2.185000 ;
      RECT 2.065000  2.185000  2.285000 2.690000 ;
      RECT 2.405000  0.645000  2.925000 0.975000 ;
      RECT 2.405000  1.345000  2.575000 2.015000 ;
      RECT 2.455000  2.355000  2.925000 2.685000 ;
      RECT 2.755000  0.975000  2.925000 1.555000 ;
      RECT 2.755000  1.555000  3.920000 1.725000 ;
      RECT 2.755000  1.725000  2.925000 2.355000 ;
      RECT 3.105000  0.935000  4.080000 1.105000 ;
      RECT 3.105000  1.105000  3.435000 1.385000 ;
      RECT 3.120000  1.895000  3.920000 2.155000 ;
      RECT 3.290000  0.085000  3.620000 0.765000 ;
      RECT 3.295000  2.360000  3.580000 3.245000 ;
      RECT 3.660000  1.285000  3.920000 1.555000 ;
      RECT 3.750000  2.155000  3.920000 2.360000 ;
      RECT 3.750000  2.360000  4.115000 2.690000 ;
      RECT 3.810000  0.280000  4.080000 0.935000 ;
      RECT 4.285000  2.355000  4.730000 3.245000 ;
      RECT 4.470000  2.105000  4.730000 2.355000 ;
      RECT 4.600000  0.085000  5.425000 0.610000 ;
      RECT 4.900000  2.105000  5.230000 2.835000 ;
      RECT 4.900000  2.835000  6.800000 3.075000 ;
      RECT 5.065000  0.610000  5.425000 0.885000 ;
      RECT 5.375000  1.380000  5.705000 1.595000 ;
      RECT 5.420000  2.125000  5.750000 2.495000 ;
      RECT 5.420000  2.495000  7.350000 2.665000 ;
      RECT 5.435000  1.210000  5.705000 1.380000 ;
      RECT 5.885000  0.285000  6.305000 0.905000 ;
      RECT 5.885000  0.905000  8.475000 1.075000 ;
      RECT 5.920000  2.105000  8.140000 2.265000 ;
      RECT 5.920000  2.265000  6.405000 2.325000 ;
      RECT 6.235000  2.095000  8.140000 2.105000 ;
      RECT 7.020000  2.435000  7.350000 2.495000 ;
      RECT 7.130000  0.085000  7.460000 0.735000 ;
      RECT 7.530000  2.435000  7.700000 3.245000 ;
      RECT 7.660000  0.315000  8.930000 0.485000 ;
      RECT 7.660000  0.485000  7.990000 0.735000 ;
      RECT 7.775000  1.075000  8.475000 1.335000 ;
      RECT 7.775000  1.335000  8.050000 2.095000 ;
      RECT 7.880000  2.265000  8.140000 2.690000 ;
      RECT 8.160000  0.665000  8.475000 0.905000 ;
      RECT 8.230000  1.585000  8.480000 1.925000 ;
      RECT 8.310000  1.925000  8.480000 3.245000 ;
      RECT 8.650000  0.485000  8.930000 3.065000 ;
      RECT 9.120000  0.700000  9.390000 1.315000 ;
      RECT 9.120000  1.315000 10.035000 1.645000 ;
      RECT 9.120000  1.645000  9.390000 2.485000 ;
      RECT 9.560000  1.825000 10.035000 3.245000 ;
      RECT 9.570000  0.085000  9.925000 1.095000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.210000  1.285000 1.380000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.210000  5.605000 1.380000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
    LAYER met1 ;
      RECT 1.055000 1.180000 1.345000 1.225000 ;
      RECT 1.055000 1.225000 5.665000 1.365000 ;
      RECT 1.055000 1.365000 1.345000 1.410000 ;
      RECT 5.375000 1.180000 5.665000 1.225000 ;
      RECT 5.375000 1.365000 5.665000 1.410000 ;
  END
END sky130_fd_sc_lp__dfstp_1
END LIBRARY
