* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_128_367# A3 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.1088e+12p pd=9.32e+06u as=1.3923e+12p ps=7.25e+06u
M1001 a_128_367# B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1002 a_390_47# A3 a_304_47# VNB nshort w=840000u l=150000u
+  ad=3.528e+11p pd=2.52e+06u as=2.352e+11p ps=2.24e+06u
M1003 Y A1 a_504_47# VNB nshort w=840000u l=150000u
+  ad=4.452e+11p pd=4.42e+06u as=2.436e+11p ps=2.26e+06u
M1004 VPWR A4 a_128_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_128_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_504_47# A2 a_390_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND B1 Y VNB nshort w=840000u l=150000u
+  ad=6.132e+11p pd=3.14e+06u as=0p ps=0u
M1008 VPWR A2 a_128_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_304_47# A4 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
