* File: sky130_fd_sc_lp__a41oi_4.pex.spice
* Created: Wed Sep  2 09:29:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 25 27 28 29
+ 30 31 48
c83 48 0 1.45437e-19 $X=1.765 $Y=1.455
r84 48 49 2.0896 $w=3.46e-07 $l=1.5e-08 $layer=POLY_cond $X=1.765 $Y=1.455
+ $X2=1.78 $Y2=1.455
r85 46 48 14.6272 $w=3.46e-07 $l=1.05e-07 $layer=POLY_cond $X=1.66 $Y=1.455
+ $X2=1.765 $Y2=1.455
r86 37 39 24.3786 $w=3.46e-07 $l=1.75e-07 $layer=POLY_cond $X=0.3 $Y=1.455
+ $X2=0.475 $Y2=1.455
r87 31 46 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.66
+ $Y=1.35 $X2=1.66 $Y2=1.35
r88 30 31 23.5611 $w=2.23e-07 $l=4.6e-07 $layer=LI1_cond $X=1.2 $Y=1.322
+ $X2=1.66 $Y2=1.322
r89 29 30 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.322
+ $X2=1.2 $Y2=1.322
r90 28 29 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.322
+ $X2=0.72 $Y2=1.322
r91 28 37 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.3
+ $Y=1.35 $X2=0.3 $Y2=1.35
r92 25 49 22.3532 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.78 $Y=1.725
+ $X2=1.78 $Y2=1.455
r93 25 27 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.78 $Y=1.725
+ $X2=1.78 $Y2=2.465
r94 22 48 22.3532 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=1.455
r95 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=0.655
r96 18 46 43.185 $w=3.46e-07 $l=3.1e-07 $layer=POLY_cond $X=1.35 $Y=1.455
+ $X2=1.66 $Y2=1.455
r97 18 43 2.0896 $w=3.46e-07 $l=1.5e-08 $layer=POLY_cond $X=1.35 $Y=1.455
+ $X2=1.335 $Y2=1.455
r98 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.35 $Y=1.515
+ $X2=1.35 $Y2=2.465
r99 15 43 22.3532 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.335 $Y=1.185
+ $X2=1.335 $Y2=1.455
r100 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.335 $Y=1.185
+ $X2=1.335 $Y2=0.655
r101 11 43 57.8121 $w=3.46e-07 $l=4.15e-07 $layer=POLY_cond $X=0.92 $Y=1.455
+ $X2=1.335 $Y2=1.455
r102 11 41 2.0896 $w=3.46e-07 $l=1.5e-08 $layer=POLY_cond $X=0.92 $Y=1.455
+ $X2=0.905 $Y2=1.455
r103 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.92 $Y=1.515
+ $X2=0.92 $Y2=2.465
r104 8 41 22.3532 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=1.455
r105 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=0.655
r106 4 41 57.8121 $w=3.46e-07 $l=4.15e-07 $layer=POLY_cond $X=0.49 $Y=1.455
+ $X2=0.905 $Y2=1.455
r107 4 39 2.0896 $w=3.46e-07 $l=1.5e-08 $layer=POLY_cond $X=0.49 $Y=1.455
+ $X2=0.475 $Y2=1.455
r108 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.49 $Y=1.515
+ $X2=0.49 $Y2=2.465
r109 1 39 22.3532 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=1.455
r110 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%A1 3 7 11 15 19 23 27 31 35 36 45 48 49 56
+ 66 74
c85 45 0 1.90297e-19 $X=3.93 $Y=1.49
c86 23 0 4.22466e-20 $X=3.59 $Y=0.745
r87 65 66 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.95 $Y=1.49 $X2=4.02
+ $Y2=1.49
r88 60 61 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.09 $Y=1.49 $X2=3.16
+ $Y2=1.49
r89 57 58 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.66 $Y=1.49 $X2=2.73
+ $Y2=1.49
r90 55 57 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.57 $Y=1.49 $X2=2.66
+ $Y2=1.49
r91 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.57
+ $Y=1.49 $X2=2.57 $Y2=1.49
r92 52 55 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.21 $Y=1.49
+ $X2=2.57 $Y2=1.49
r93 49 74 5.9984 $w=3.63e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=1.392
+ $X2=3.205 $Y2=1.392
r94 48 56 2.21016 $w=3.63e-07 $l=7e-08 $layer=LI1_cond $X=2.64 $Y=1.392 $X2=2.57
+ $Y2=1.392
r95 46 65 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.93 $Y=1.49 $X2=3.95
+ $Y2=1.49
r96 46 63 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.93 $Y=1.49
+ $X2=3.59 $Y2=1.49
r97 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=1.49 $X2=3.93 $Y2=1.49
r98 43 63 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.25 $Y=1.49
+ $X2=3.59 $Y2=1.49
r99 43 61 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.25 $Y=1.49 $X2=3.16
+ $Y2=1.49
r100 42 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.25 $Y=1.49
+ $X2=3.93 $Y2=1.49
r101 42 74 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.25 $Y=1.49
+ $X2=3.205 $Y2=1.49
r102 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.49 $X2=3.25 $Y2=1.49
r103 39 60 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.91 $Y=1.49
+ $X2=3.09 $Y2=1.49
r104 39 58 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.91 $Y=1.49
+ $X2=2.73 $Y2=1.49
r105 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.49 $X2=2.91 $Y2=1.49
r106 36 48 3.06266 $w=3.63e-07 $l=9.7e-08 $layer=LI1_cond $X=2.737 $Y=1.392
+ $X2=2.64 $Y2=1.392
r107 36 38 5.46226 $w=3.63e-07 $l=1.73e-07 $layer=LI1_cond $X=2.737 $Y=1.392
+ $X2=2.91 $Y2=1.392
r108 35 49 3.06266 $w=3.63e-07 $l=9.7e-08 $layer=LI1_cond $X=3.023 $Y=1.392
+ $X2=3.12 $Y2=1.392
r109 35 38 3.56784 $w=3.63e-07 $l=1.13e-07 $layer=LI1_cond $X=3.023 $Y=1.392
+ $X2=2.91 $Y2=1.392
r110 29 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.02 $Y=1.325
+ $X2=4.02 $Y2=1.49
r111 29 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.02 $Y=1.325
+ $X2=4.02 $Y2=0.745
r112 25 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.655
+ $X2=3.95 $Y2=1.49
r113 25 27 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.95 $Y=1.655
+ $X2=3.95 $Y2=2.465
r114 21 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.59 $Y=1.325
+ $X2=3.59 $Y2=1.49
r115 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.59 $Y=1.325
+ $X2=3.59 $Y2=0.745
r116 17 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.16 $Y=1.325
+ $X2=3.16 $Y2=1.49
r117 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.16 $Y=1.325
+ $X2=3.16 $Y2=0.745
r118 13 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.655
+ $X2=3.09 $Y2=1.49
r119 13 15 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.09 $Y=1.655
+ $X2=3.09 $Y2=2.465
r120 9 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=1.49
r121 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.73 $Y=1.325
+ $X2=2.73 $Y2=0.745
r122 5 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=1.655
+ $X2=2.66 $Y2=1.49
r123 5 7 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.66 $Y=1.655 $X2=2.66
+ $Y2=2.465
r124 1 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.655
+ $X2=2.21 $Y2=1.49
r125 1 3 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.21 $Y=1.655 $X2=2.21
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%A2 3 5 7 10 12 14 17 19 21 22 24 27 29 30 45
+ 47
c96 47 0 1.90297e-19 $X=5.83 $Y=1.44
c97 3 0 1.80978e-19 $X=4.38 $Y=2.465
r98 46 47 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.82 $Y=1.44 $X2=5.83
+ $Y2=1.44
r99 44 46 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.81 $Y=1.44 $X2=5.82
+ $Y2=1.44
r100 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.81
+ $Y=1.44 $X2=5.81 $Y2=1.44
r101 42 44 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=5.39 $Y=1.44
+ $X2=5.81 $Y2=1.44
r102 41 42 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.24 $Y=1.44
+ $X2=5.39 $Y2=1.44
r103 40 41 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=4.96 $Y=1.44
+ $X2=5.24 $Y2=1.44
r104 39 40 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.81 $Y=1.44
+ $X2=4.96 $Y2=1.44
r105 37 39 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.79 $Y=1.44 $X2=4.81
+ $Y2=1.44
r106 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.79
+ $Y=1.44 $X2=4.79 $Y2=1.44
r107 35 37 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=4.53 $Y=1.44
+ $X2=4.79 $Y2=1.44
r108 33 35 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.38 $Y=1.44
+ $X2=4.53 $Y2=1.44
r109 30 45 8.56945 $w=3.88e-07 $l=2.9e-07 $layer=LI1_cond $X=5.52 $Y=1.39
+ $X2=5.81 $Y2=1.39
r110 29 30 14.1839 $w=3.88e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.39
+ $X2=5.52 $Y2=1.39
r111 29 38 7.38745 $w=3.88e-07 $l=2.5e-07 $layer=LI1_cond $X=5.04 $Y=1.39
+ $X2=4.79 $Y2=1.39
r112 25 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.83 $Y=1.605
+ $X2=5.83 $Y2=1.44
r113 25 27 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.83 $Y=1.605
+ $X2=5.83 $Y2=2.465
r114 22 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.82 $Y=1.275
+ $X2=5.82 $Y2=1.44
r115 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.82 $Y=1.275
+ $X2=5.82 $Y2=0.745
r116 19 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.39 $Y=1.275
+ $X2=5.39 $Y2=1.44
r117 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.39 $Y=1.275
+ $X2=5.39 $Y2=0.745
r118 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=1.605
+ $X2=5.24 $Y2=1.44
r119 15 17 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.24 $Y=1.605
+ $X2=5.24 $Y2=2.465
r120 12 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.96 $Y=1.275
+ $X2=4.96 $Y2=1.44
r121 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.96 $Y=1.275
+ $X2=4.96 $Y2=0.745
r122 8 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.81 $Y=1.605
+ $X2=4.81 $Y2=1.44
r123 8 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.81 $Y=1.605
+ $X2=4.81 $Y2=2.465
r124 5 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.53 $Y=1.275
+ $X2=4.53 $Y2=1.44
r125 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.53 $Y=1.275
+ $X2=4.53 $Y2=0.745
r126 1 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.38 $Y=1.605
+ $X2=4.38 $Y2=1.44
r127 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.38 $Y=1.605
+ $X2=4.38 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%A3 3 7 9 11 14 16 18 19 21 24 26 28 36 39 50
+ 54
c91 19 0 1.51646e-19 $X=7.655 $Y=1.275
c92 16 0 1.51646e-19 $X=7.225 $Y=1.275
r93 53 54 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.07 $Y=1.44
+ $X2=8.085 $Y2=1.44
r94 49 51 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=7.37 $Y=1.44
+ $X2=7.655 $Y2=1.44
r95 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.37
+ $Y=1.44 $X2=7.37 $Y2=1.44
r96 47 49 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=7.225 $Y=1.44
+ $X2=7.37 $Y2=1.44
r97 46 47 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=7.12 $Y=1.44
+ $X2=7.225 $Y2=1.44
r98 45 46 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=6.795 $Y=1.44
+ $X2=7.12 $Y2=1.44
r99 44 45 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=6.69 $Y=1.44
+ $X2=6.795 $Y2=1.44
r100 39 50 8.46412 $w=1.88e-07 $l=1.45e-07 $layer=LI1_cond $X=7.44 $Y=1.295
+ $X2=7.44 $Y2=1.44
r101 37 53 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=8.05 $Y=1.44 $X2=8.07
+ $Y2=1.44
r102 37 51 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=8.05 $Y=1.44
+ $X2=7.655 $Y2=1.44
r103 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.05
+ $Y=1.44 $X2=8.05 $Y2=1.44
r104 34 50 1.7512 $w=1.88e-07 $l=3e-08 $layer=LI1_cond $X=7.44 $Y=1.47 $X2=7.44
+ $Y2=1.44
r105 34 36 25.8047 $w=2.28e-07 $l=5.15e-07 $layer=LI1_cond $X=7.535 $Y=1.47
+ $X2=8.05 $Y2=1.47
r106 32 44 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.35 $Y=1.44
+ $X2=6.69 $Y2=1.44
r107 32 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.35 $Y=1.44 $X2=6.26
+ $Y2=1.44
r108 31 50 42.4697 $w=2.68e-07 $l=9.95e-07 $layer=LI1_cond $X=6.35 $Y=1.45
+ $X2=7.345 $Y2=1.45
r109 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.35
+ $Y=1.44 $X2=6.35 $Y2=1.44
r110 26 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.085 $Y=1.275
+ $X2=8.085 $Y2=1.44
r111 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.085 $Y=1.275
+ $X2=8.085 $Y2=0.745
r112 22 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.07 $Y=1.605
+ $X2=8.07 $Y2=1.44
r113 22 24 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.07 $Y=1.605
+ $X2=8.07 $Y2=2.465
r114 19 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.275
+ $X2=7.655 $Y2=1.44
r115 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.655 $Y=1.275
+ $X2=7.655 $Y2=0.745
r116 16 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.225 $Y=1.275
+ $X2=7.225 $Y2=1.44
r117 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.225 $Y=1.275
+ $X2=7.225 $Y2=0.745
r118 12 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.12 $Y=1.605
+ $X2=7.12 $Y2=1.44
r119 12 14 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.12 $Y=1.605
+ $X2=7.12 $Y2=2.465
r120 9 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.275
+ $X2=6.795 $Y2=1.44
r121 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.795 $Y=1.275
+ $X2=6.795 $Y2=0.745
r122 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.605
+ $X2=6.69 $Y2=1.44
r123 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.69 $Y=1.605
+ $X2=6.69 $Y2=2.465
r124 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.26 $Y=1.605
+ $X2=6.26 $Y2=1.44
r125 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.26 $Y=1.605
+ $X2=6.26 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%A4 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 37 39
c76 19 0 9.06625e-20 $X=9.375 $Y=1.275
c77 12 0 9.06625e-20 $X=8.945 $Y=1.275
r78 55 56 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.79 $Y=1.44
+ $X2=9.805 $Y2=1.44
r79 53 55 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=9.61 $Y=1.44 $X2=9.79
+ $Y2=1.44
r80 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.61
+ $Y=1.44 $X2=9.61 $Y2=1.44
r81 51 53 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=9.375 $Y=1.44
+ $X2=9.61 $Y2=1.44
r82 50 51 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.36 $Y=1.44
+ $X2=9.375 $Y2=1.44
r83 49 50 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=8.945 $Y=1.44
+ $X2=9.36 $Y2=1.44
r84 48 49 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.93 $Y=1.44
+ $X2=8.945 $Y2=1.44
r85 46 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.59 $Y=1.44
+ $X2=8.93 $Y2=1.44
r86 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.59
+ $Y=1.44 $X2=8.59 $Y2=1.44
r87 44 46 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.515 $Y=1.44
+ $X2=8.59 $Y2=1.44
r88 42 44 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.5 $Y=1.44
+ $X2=8.515 $Y2=1.44
r89 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.29
+ $Y=1.44 $X2=10.29 $Y2=1.44
r90 37 56 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.88 $Y=1.44
+ $X2=9.805 $Y2=1.44
r91 37 39 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=9.88 $Y=1.44
+ $X2=10.29 $Y2=1.44
r92 32 40 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=10.32 $Y=1.392
+ $X2=10.29 $Y2=1.392
r93 31 40 13.4701 $w=3.83e-07 $l=4.5e-07 $layer=LI1_cond $X=9.84 $Y=1.392
+ $X2=10.29 $Y2=1.392
r94 31 54 6.88472 $w=3.83e-07 $l=2.3e-07 $layer=LI1_cond $X=9.84 $Y=1.392
+ $X2=9.61 $Y2=1.392
r95 30 54 7.4834 $w=3.83e-07 $l=2.5e-07 $layer=LI1_cond $X=9.36 $Y=1.392
+ $X2=9.61 $Y2=1.392
r96 29 30 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.392
+ $X2=9.36 $Y2=1.392
r97 29 47 8.68074 $w=3.83e-07 $l=2.9e-07 $layer=LI1_cond $X=8.88 $Y=1.392
+ $X2=8.59 $Y2=1.392
r98 26 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.805 $Y=1.275
+ $X2=9.805 $Y2=1.44
r99 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.805 $Y=1.275
+ $X2=9.805 $Y2=0.745
r100 22 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.79 $Y=1.605
+ $X2=9.79 $Y2=1.44
r101 22 24 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=9.79 $Y=1.605
+ $X2=9.79 $Y2=2.465
r102 19 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.375 $Y=1.275
+ $X2=9.375 $Y2=1.44
r103 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.375 $Y=1.275
+ $X2=9.375 $Y2=0.745
r104 15 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.36 $Y=1.605
+ $X2=9.36 $Y2=1.44
r105 15 17 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=9.36 $Y=1.605
+ $X2=9.36 $Y2=2.465
r106 12 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.945 $Y=1.275
+ $X2=8.945 $Y2=1.44
r107 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.945 $Y=1.275
+ $X2=8.945 $Y2=0.745
r108 8 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.93 $Y=1.605
+ $X2=8.93 $Y2=1.44
r109 8 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.93 $Y=1.605
+ $X2=8.93 $Y2=2.465
r110 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.515 $Y=1.275
+ $X2=8.515 $Y2=1.44
r111 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.515 $Y=1.275
+ $X2=8.515 $Y2=0.745
r112 1 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.5 $Y=1.605
+ $X2=8.5 $Y2=1.44
r113 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.5 $Y=1.605 $X2=8.5
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%A_30_367# 1 2 3 4 5 6 7 8 9 10 11 34 36 38
+ 42 44 46 48 52 56 58 63 66 68 69 72 76 80 84 88 92 96 100 104 111 115 117 118
+ 119 120 121 122
c141 69 0 1.80978e-19 $X=5.13 $Y=1.84
r142 104 106 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=10.04 $Y=1.98
+ $X2=10.04 $Y2=2.91
r143 102 104 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=10.04 $Y=1.925
+ $X2=10.04 $Y2=1.98
r144 101 122 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.24 $Y=1.84
+ $X2=9.145 $Y2=1.84
r145 100 102 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.91 $Y=1.84
+ $X2=10.04 $Y2=1.925
r146 100 101 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.91 $Y=1.84
+ $X2=9.24 $Y2=1.84
r147 96 98 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=9.145 $Y=1.98
+ $X2=9.145 $Y2=2.91
r148 94 122 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=1.925
+ $X2=9.145 $Y2=1.84
r149 94 96 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=9.145 $Y=1.925
+ $X2=9.145 $Y2=1.98
r150 93 121 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.38 $Y=1.84
+ $X2=8.285 $Y2=1.84
r151 92 122 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.05 $Y=1.84
+ $X2=9.145 $Y2=1.84
r152 92 93 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.05 $Y=1.84
+ $X2=8.38 $Y2=1.84
r153 88 90 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=8.285 $Y=1.98
+ $X2=8.285 $Y2=2.91
r154 86 121 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.285 $Y=1.925
+ $X2=8.285 $Y2=1.84
r155 86 88 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=8.285 $Y=1.925
+ $X2=8.285 $Y2=1.98
r156 85 120 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7 $Y=1.84 $X2=6.905
+ $Y2=1.84
r157 84 121 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.19 $Y=1.84
+ $X2=8.285 $Y2=1.84
r158 84 85 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=8.19 $Y=1.84 $X2=7
+ $Y2=1.84
r159 80 82 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.905 $Y=1.98
+ $X2=6.905 $Y2=2.91
r160 78 120 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=1.925
+ $X2=6.905 $Y2=1.84
r161 78 80 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.905 $Y=1.925
+ $X2=6.905 $Y2=1.98
r162 77 119 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.14 $Y=1.84
+ $X2=6.01 $Y2=1.84
r163 76 120 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.81 $Y=1.84
+ $X2=6.905 $Y2=1.84
r164 76 77 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.81 $Y=1.84
+ $X2=6.14 $Y2=1.84
r165 72 74 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=6.01 $Y=1.98
+ $X2=6.01 $Y2=2.91
r166 70 119 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=1.925
+ $X2=6.01 $Y2=1.84
r167 70 72 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=6.01 $Y=1.925
+ $X2=6.01 $Y2=1.98
r168 68 119 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.88 $Y=1.84
+ $X2=6.01 $Y2=1.84
r169 68 69 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.88 $Y=1.84
+ $X2=5.13 $Y2=1.84
r170 64 118 3.83171 $w=2.55e-07 $l=9.72111e-08 $layer=LI1_cond $X=5.01 $Y=2.285
+ $X2=4.995 $Y2=2.195
r171 64 66 6.96268 $w=2.38e-07 $l=1.45e-07 $layer=LI1_cond $X=5.01 $Y=2.285
+ $X2=5.01 $Y2=2.43
r172 61 118 3.83171 $w=2.55e-07 $l=9e-08 $layer=LI1_cond $X=4.995 $Y=2.105
+ $X2=4.995 $Y2=2.195
r173 61 63 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.995 $Y=2.105
+ $X2=4.995 $Y2=1.98
r174 60 69 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.995 $Y=1.925
+ $X2=5.13 $Y2=1.84
r175 60 63 2.34757 $w=2.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.995 $Y=1.925
+ $X2=4.995 $Y2=1.98
r176 59 117 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=2.195
+ $X2=4.165 $Y2=2.195
r177 58 118 2.62201 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=4.86 $Y=2.195
+ $X2=4.995 $Y2=2.195
r178 58 59 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=4.86 $Y=2.195
+ $X2=4.33 $Y2=2.195
r179 54 117 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.165 $Y=2.285
+ $X2=4.165 $Y2=2.195
r180 54 56 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=4.165 $Y=2.285
+ $X2=4.165 $Y2=2.97
r181 53 115 5.86152 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=2.195
+ $X2=2.885 $Y2=2.195
r182 52 117 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=2.195
+ $X2=4.165 $Y2=2.195
r183 52 53 62.2323 $w=1.78e-07 $l=1.01e-06 $layer=LI1_cond $X=4 $Y=2.195
+ $X2=2.99 $Y2=2.195
r184 49 113 3.69874 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=2.11 $Y=2.195
+ $X2=2.005 $Y2=2.195
r185 48 115 5.86152 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=2.78 $Y=2.195
+ $X2=2.885 $Y2=2.195
r186 48 49 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.78 $Y=2.195
+ $X2=2.11 $Y2=2.195
r187 46 113 3.17035 $w=2.1e-07 $l=9e-08 $layer=LI1_cond $X=2.005 $Y=2.285
+ $X2=2.005 $Y2=2.195
r188 46 47 32.7446 $w=2.08e-07 $l=6.2e-07 $layer=LI1_cond $X=2.005 $Y=2.285
+ $X2=2.005 $Y2=2.905
r189 45 111 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.23 $Y=2.99
+ $X2=1.135 $Y2=2.99
r190 44 47 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.9 $Y=2.99
+ $X2=2.005 $Y2=2.905
r191 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.9 $Y=2.99
+ $X2=1.23 $Y2=2.99
r192 40 111 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=2.905
+ $X2=1.135 $Y2=2.99
r193 40 42 45.5311 $w=1.88e-07 $l=7.8e-07 $layer=LI1_cond $X=1.135 $Y=2.905
+ $X2=1.135 $Y2=2.125
r194 39 109 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.37 $Y=2.99
+ $X2=0.24 $Y2=2.99
r195 38 111 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.04 $Y=2.99
+ $X2=1.135 $Y2=2.99
r196 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.04 $Y=2.99
+ $X2=0.37 $Y2=2.99
r197 34 109 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.905
+ $X2=0.24 $Y2=2.99
r198 34 36 40.5571 $w=2.58e-07 $l=9.15e-07 $layer=LI1_cond $X=0.24 $Y=2.905
+ $X2=0.24 $Y2=1.99
r199 11 106 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.865
+ $Y=1.835 $X2=10.005 $Y2=2.91
r200 11 104 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.865
+ $Y=1.835 $X2=10.005 $Y2=1.98
r201 10 98 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.005
+ $Y=1.835 $X2=9.145 $Y2=2.91
r202 10 96 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.005
+ $Y=1.835 $X2=9.145 $Y2=1.98
r203 9 90 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.145
+ $Y=1.835 $X2=8.285 $Y2=2.91
r204 9 88 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.145
+ $Y=1.835 $X2=8.285 $Y2=1.98
r205 8 82 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.765
+ $Y=1.835 $X2=6.905 $Y2=2.91
r206 8 80 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.765
+ $Y=1.835 $X2=6.905 $Y2=1.98
r207 7 74 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.905
+ $Y=1.835 $X2=6.045 $Y2=2.91
r208 7 72 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.905
+ $Y=1.835 $X2=6.045 $Y2=1.98
r209 6 66 300 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_PDIFF $count=2 $X=4.885
+ $Y=1.835 $X2=5.025 $Y2=2.43
r210 6 63 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.885
+ $Y=1.835 $X2=5.025 $Y2=1.98
r211 5 117 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.835 $X2=4.165 $Y2=2.22
r212 5 56 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.835 $X2=4.165 $Y2=2.97
r213 4 115 300 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=2 $X=2.735
+ $Y=1.835 $X2=2.875 $Y2=2.27
r214 3 113 300 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=2 $X=1.855
+ $Y=1.835 $X2=1.995 $Y2=2.27
r215 2 111 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.91
r216 2 42 400 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.125
r217 1 109 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.91
r218 1 36 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%Y 1 2 3 4 5 6 21 27 29 30 32 35 41 43 45 48
+ 50 51 52 53 54 55 56 64 67 79 82
c121 64 0 6.46567e-20 $X=3.64 $Y=0.927
c122 45 0 4.22466e-20 $X=4.265 $Y=1.15
c123 43 0 8.07799e-20 $X=4.265 $Y=1.84
r124 85 86 7.78772 $w=3.28e-07 $l=2.23e-07 $layer=LI1_cond $X=3.805 $Y=0.927
+ $X2=3.805 $Y2=1.15
r125 65 67 1.79269 $w=2.23e-07 $l=3.5e-08 $layer=LI1_cond $X=1.645 $Y=0.927
+ $X2=1.68 $Y2=0.927
r126 64 85 2.99809 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=0.927
+ $X2=3.805 $Y2=0.927
r127 64 79 2.04879 $w=2.23e-07 $l=4e-08 $layer=LI1_cond $X=3.64 $Y=0.927 $X2=3.6
+ $Y2=0.927
r128 56 85 0.069845 $w=3.28e-07 $l=2e-09 $layer=LI1_cond $X=3.805 $Y=0.925
+ $X2=3.805 $Y2=0.927
r129 56 82 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.805 $Y=0.925
+ $X2=3.805 $Y2=0.68
r130 56 79 1.17805 $w=2.23e-07 $l=2.3e-08 $layer=LI1_cond $X=3.577 $Y=0.927
+ $X2=3.6 $Y2=0.927
r131 55 56 23.4074 $w=2.23e-07 $l=4.57e-07 $layer=LI1_cond $X=3.12 $Y=0.927
+ $X2=3.577 $Y2=0.927
r132 55 74 8.96345 $w=2.23e-07 $l=1.75e-07 $layer=LI1_cond $X=3.12 $Y=0.927
+ $X2=2.945 $Y2=0.927
r133 54 74 15.622 $w=2.23e-07 $l=3.05e-07 $layer=LI1_cond $X=2.64 $Y=0.927
+ $X2=2.945 $Y2=0.927
r134 53 54 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0.927
+ $X2=2.64 $Y2=0.927
r135 52 65 4.84724 $w=2.05e-07 $l=9.5e-08 $layer=LI1_cond $X=1.55 $Y=0.927
+ $X2=1.645 $Y2=0.927
r136 52 53 23.305 $w=2.23e-07 $l=4.55e-07 $layer=LI1_cond $X=1.705 $Y=0.927
+ $X2=2.16 $Y2=0.927
r137 52 67 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=1.705 $Y=0.927
+ $X2=1.68 $Y2=0.927
r138 49 51 10.7874 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.565 $Y=1.77
+ $X2=1.815 $Y2=1.77
r139 49 50 7.96936 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=1.77
+ $X2=1.4 $Y2=1.77
r140 47 48 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=4.36 $Y=1.235
+ $X2=4.36 $Y2=1.745
r141 46 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.97 $Y=1.15
+ $X2=3.805 $Y2=1.15
r142 45 47 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.265 $Y=1.15
+ $X2=4.36 $Y2=1.235
r143 45 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.265 $Y=1.15
+ $X2=3.97 $Y2=1.15
r144 43 48 6.81649 $w=1.9e-07 $l=1.3435e-07 $layer=LI1_cond $X=4.265 $Y=1.84
+ $X2=4.36 $Y2=1.745
r145 43 51 143.014 $w=1.88e-07 $l=2.45e-06 $layer=LI1_cond $X=4.265 $Y=1.84
+ $X2=1.815 $Y2=1.84
r146 39 52 1.61756 $w=1.9e-07 $l=1.12e-07 $layer=LI1_cond $X=1.55 $Y=0.815
+ $X2=1.55 $Y2=0.927
r147 39 41 23.0574 $w=1.88e-07 $l=3.95e-07 $layer=LI1_cond $X=1.55 $Y=0.815
+ $X2=1.55 $Y2=0.42
r148 35 37 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.565 $Y=1.97
+ $X2=1.565 $Y2=2.65
r149 33 49 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=1.935
+ $X2=1.565 $Y2=1.77
r150 33 35 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.565 $Y=1.935
+ $X2=1.565 $Y2=1.97
r151 32 50 31.774 $w=1.83e-07 $l=5.3e-07 $layer=LI1_cond $X=0.87 $Y=1.697
+ $X2=1.4 $Y2=1.697
r152 29 52 4.84724 $w=2.05e-07 $l=1.04523e-07 $layer=LI1_cond $X=1.455 $Y=0.947
+ $X2=1.55 $Y2=0.927
r153 29 30 40.1671 $w=1.83e-07 $l=6.7e-07 $layer=LI1_cond $X=1.455 $Y=0.947
+ $X2=0.785 $Y2=0.947
r154 25 30 6.81807 $w=1.85e-07 $l=1.33285e-07 $layer=LI1_cond $X=0.69 $Y=0.855
+ $X2=0.785 $Y2=0.947
r155 25 27 25.3923 $w=1.88e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=0.855
+ $X2=0.69 $Y2=0.42
r156 21 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.705 $Y=1.97
+ $X2=0.705 $Y2=2.65
r157 19 32 7.54394 $w=1.85e-07 $l=2.06325e-07 $layer=LI1_cond $X=0.705 $Y=1.79
+ $X2=0.87 $Y2=1.697
r158 19 21 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.705 $Y=1.79
+ $X2=0.705 $Y2=1.97
r159 6 37 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=2.65
r160 6 35 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=1.97
r161 5 23 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.65
r162 5 21 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=1.97
r163 4 82 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=3.665
+ $Y=0.325 $X2=3.805 $Y2=0.68
r164 3 74 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.325 $X2=2.945 $Y2=0.92
r165 2 41 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.42
r166 1 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%VPWR 1 2 3 4 5 6 7 8 27 31 33 37 41 47 53 59
+ 65 70 71 73 74 76 77 78 87 91 96 101 114 115 118 121 124 127 130
r148 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r149 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r150 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r151 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r152 119 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r153 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r154 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r155 112 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r156 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r157 109 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r158 109 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r159 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r160 106 130 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=8.02 $Y=3.33
+ $X2=7.595 $Y2=3.33
r161 106 108 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.02 $Y=3.33
+ $X2=8.4 $Y2=3.33
r162 105 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r163 105 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r164 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r165 102 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.64 $Y=3.33
+ $X2=6.475 $Y2=3.33
r166 102 104 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.64 $Y=3.33
+ $X2=6.96 $Y2=3.33
r167 101 130 15.0812 $w=1.7e-07 $l=4.25e-07 $layer=LI1_cond $X=7.17 $Y=3.33
+ $X2=7.595 $Y2=3.33
r168 101 104 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.17 $Y=3.33
+ $X2=6.96 $Y2=3.33
r169 100 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r170 100 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r171 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r172 97 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.7 $Y=3.33
+ $X2=5.535 $Y2=3.33
r173 97 99 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=5.7 $Y=3.33 $X2=6
+ $Y2=3.33
r174 96 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.31 $Y=3.33
+ $X2=6.475 $Y2=3.33
r175 96 99 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.31 $Y=3.33 $X2=6
+ $Y2=3.33
r176 95 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r177 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r178 92 121 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.72 $Y=3.33
+ $X2=4.61 $Y2=3.33
r179 92 94 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.72 $Y=3.33
+ $X2=5.04 $Y2=3.33
r180 91 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=3.33
+ $X2=5.535 $Y2=3.33
r181 91 94 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.37 $Y=3.33
+ $X2=5.04 $Y2=3.33
r182 90 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r183 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r184 87 118 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.16 $Y=3.33
+ $X2=3.495 $Y2=3.33
r185 87 89 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r186 86 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r187 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r188 82 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r189 81 85 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r190 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r191 78 125 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r192 78 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r193 76 111 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=9.41 $Y=3.33
+ $X2=9.36 $Y2=3.33
r194 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.41 $Y=3.33
+ $X2=9.575 $Y2=3.33
r195 75 114 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=9.74 $Y=3.33
+ $X2=10.32 $Y2=3.33
r196 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.74 $Y=3.33
+ $X2=9.575 $Y2=3.33
r197 73 108 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.55 $Y=3.33
+ $X2=8.4 $Y2=3.33
r198 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.55 $Y=3.33
+ $X2=8.715 $Y2=3.33
r199 72 111 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r200 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=8.715 $Y2=3.33
r201 70 85 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.16 $Y2=3.33
r202 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=3.33
+ $X2=2.445 $Y2=3.33
r203 69 89 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=3.12 $Y2=3.33
r204 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=3.33
+ $X2=2.445 $Y2=3.33
r205 65 68 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=9.575 $Y=2.19
+ $X2=9.575 $Y2=2.95
r206 63 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.575 $Y=3.245
+ $X2=9.575 $Y2=3.33
r207 63 68 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.575 $Y=3.245
+ $X2=9.575 $Y2=2.95
r208 59 62 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=8.715 $Y=2.19
+ $X2=8.715 $Y2=2.95
r209 57 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.715 $Y=3.245
+ $X2=8.715 $Y2=3.33
r210 57 62 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.715 $Y=3.245
+ $X2=8.715 $Y2=2.95
r211 53 56 10.9082 $w=8.48e-07 $l=7.6e-07 $layer=LI1_cond $X=7.595 $Y=2.19
+ $X2=7.595 $Y2=2.95
r212 51 130 3.24638 $w=8.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.595 $Y=3.245
+ $X2=7.595 $Y2=3.33
r213 51 56 4.23412 $w=8.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.595 $Y=3.245
+ $X2=7.595 $Y2=2.95
r214 47 50 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=6.475 $Y=2.19
+ $X2=6.475 $Y2=2.95
r215 45 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.475 $Y=3.245
+ $X2=6.475 $Y2=3.33
r216 45 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.475 $Y=3.245
+ $X2=6.475 $Y2=2.95
r217 41 44 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.535 $Y=2.19
+ $X2=5.535 $Y2=2.95
r218 39 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=3.245
+ $X2=5.535 $Y2=3.33
r219 39 44 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.535 $Y=3.245
+ $X2=5.535 $Y2=2.95
r220 35 121 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=3.245
+ $X2=4.61 $Y2=3.33
r221 35 37 32.7399 $w=2.18e-07 $l=6.25e-07 $layer=LI1_cond $X=4.61 $Y=3.245
+ $X2=4.61 $Y2=2.62
r222 34 118 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.83 $Y=3.33
+ $X2=3.495 $Y2=3.33
r223 33 121 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.5 $Y=3.33
+ $X2=4.61 $Y2=3.33
r224 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.5 $Y=3.33
+ $X2=3.83 $Y2=3.33
r225 29 118 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=3.245
+ $X2=3.495 $Y2=3.33
r226 29 31 12.1393 $w=6.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.495 $Y=3.245
+ $X2=3.495 $Y2=2.565
r227 25 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=3.245
+ $X2=2.445 $Y2=3.33
r228 25 27 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=2.445 $Y=3.245
+ $X2=2.445 $Y2=2.62
r229 8 68 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.435
+ $Y=1.835 $X2=9.575 $Y2=2.95
r230 8 65 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=9.435
+ $Y=1.835 $X2=9.575 $Y2=2.19
r231 7 62 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.835 $X2=8.715 $Y2=2.95
r232 7 59 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=8.575
+ $Y=1.835 $X2=8.715 $Y2=2.19
r233 6 56 200 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=3 $X=7.195
+ $Y=1.835 $X2=7.335 $Y2=2.95
r234 6 53 200 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=3 $X=7.195
+ $Y=1.835 $X2=7.335 $Y2=2.19
r235 5 50 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.335
+ $Y=1.835 $X2=6.475 $Y2=2.95
r236 5 47 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=6.335
+ $Y=1.835 $X2=6.475 $Y2=2.19
r237 4 44 400 $w=1.7e-07 $l=1.22005e-06 $layer=licon1_PDIFF $count=1 $X=5.315
+ $Y=1.835 $X2=5.535 $Y2=2.95
r238 4 41 400 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_PDIFF $count=1 $X=5.315
+ $Y=1.835 $X2=5.535 $Y2=2.19
r239 3 37 300 $w=1.7e-07 $l=8.5213e-07 $layer=licon1_PDIFF $count=2 $X=4.455
+ $Y=1.835 $X2=4.595 $Y2=2.62
r240 2 31 150 $w=1.7e-07 $l=9.47576e-07 $layer=licon1_PDIFF $count=4 $X=3.165
+ $Y=1.835 $X2=3.665 $Y2=2.565
r241 1 27 300 $w=1.7e-07 $l=8.61293e-07 $layer=licon1_PDIFF $count=2 $X=2.285
+ $Y=1.835 $X2=2.445 $Y2=2.62
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 45 47 66 67 73
r117 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r118 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r119 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r120 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.32 $Y2=0
r121 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r122 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r123 60 61 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r124 57 60 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=8.4
+ $Y2=0
r125 57 58 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r126 55 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r127 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r128 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r129 52 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.12
+ $Y2=0
r130 52 54 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.68 $Y2=0
r131 51 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r132 51 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r133 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r134 48 70 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r135 48 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r136 47 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.12
+ $Y2=0
r137 47 50 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=0
+ $X2=0.72 $Y2=0
r138 45 61 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=8.4
+ $Y2=0
r139 45 58 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=2.16 $Y2=0
r140 43 63 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=9.425 $Y=0 $X2=9.36
+ $Y2=0
r141 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.425 $Y=0 $X2=9.59
+ $Y2=0
r142 42 66 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=9.755 $Y=0
+ $X2=10.32 $Y2=0
r143 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.755 $Y=0 $X2=9.59
+ $Y2=0
r144 40 60 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.565 $Y=0 $X2=8.4
+ $Y2=0
r145 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.565 $Y=0 $X2=8.73
+ $Y2=0
r146 39 63 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.895 $Y=0
+ $X2=9.36 $Y2=0
r147 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.895 $Y=0 $X2=8.73
+ $Y2=0
r148 37 54 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=0
+ $X2=1.68 $Y2=0
r149 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.98
+ $Y2=0
r150 36 57 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.16
+ $Y2=0
r151 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=1.98
+ $Y2=0
r152 32 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.59 $Y=0.085
+ $X2=9.59 $Y2=0
r153 32 34 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.59 $Y=0.085
+ $X2=9.59 $Y2=0.565
r154 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.73 $Y=0.085
+ $X2=8.73 $Y2=0
r155 28 30 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.73 $Y=0.085
+ $X2=8.73 $Y2=0.565
r156 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r157 24 26 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.505
r158 20 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r159 20 22 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.545
r160 16 70 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r161 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r162 5 34 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=9.45
+ $Y=0.325 $X2=9.59 $Y2=0.565
r163 4 30 182 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_NDIFF $count=1 $X=8.59
+ $Y=0.325 $X2=8.73 $Y2=0.565
r164 3 26 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.505
r165 2 22 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.545
r166 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%A_478_65# 1 2 3 4 5 16 20 24 28 30 34 35 38
r46 37 38 6.83464 $w=3.88e-07 $l=1.05e-07 $layer=LI1_cond $X=5.175 $Y=0.45
+ $X2=5.07 $Y2=0.45
r47 33 34 6.53914 $w=3.88e-07 $l=9.5e-08 $layer=LI1_cond $X=3.375 $Y=0.45
+ $X2=3.47 $Y2=0.45
r48 28 37 8.4217 $w=3.88e-07 $l=2.85e-07 $layer=LI1_cond $X=5.46 $Y=0.45
+ $X2=5.175 $Y2=0.45
r49 28 30 16.9911 $w=3.88e-07 $l=5.75e-07 $layer=LI1_cond $X=5.46 $Y=0.45
+ $X2=6.035 $Y2=0.45
r50 27 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.48 $Y=0.34
+ $X2=4.315 $Y2=0.34
r51 27 38 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.48 $Y=0.34 $X2=5.07
+ $Y2=0.34
r52 22 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=0.425
+ $X2=4.315 $Y2=0.34
r53 22 24 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=4.315 $Y=0.425
+ $X2=4.315 $Y2=0.45
r54 20 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.15 $Y=0.34
+ $X2=4.315 $Y2=0.34
r55 20 34 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.15 $Y=0.34
+ $X2=3.47 $Y2=0.34
r56 16 33 2.95498 $w=3.88e-07 $l=1e-07 $layer=LI1_cond $X=3.275 $Y=0.45
+ $X2=3.375 $Y2=0.45
r57 16 18 22.4579 $w=3.88e-07 $l=7.6e-07 $layer=LI1_cond $X=3.275 $Y=0.45
+ $X2=2.515 $Y2=0.45
r58 5 30 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.895
+ $Y=0.325 $X2=6.035 $Y2=0.47
r59 4 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.035
+ $Y=0.325 $X2=5.175 $Y2=0.47
r60 3 24 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=4.095
+ $Y=0.325 $X2=4.315 $Y2=0.45
r61 2 33 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.235
+ $Y=0.325 $X2=3.375 $Y2=0.47
r62 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.325 $X2=2.515 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%A_921_65# 1 2 3 4 13 17 20 25 31
r50 31 33 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=7.87 $Y=0.7 $X2=7.87
+ $Y2=0.9
r51 27 28 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=7.01 $Y=0.9 $X2=7.01
+ $Y2=0.92
r52 25 27 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=7.01 $Y=0.7 $X2=7.01
+ $Y2=0.9
r53 20 22 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=4.775 $Y=0.76
+ $X2=4.775 $Y2=0.92
r54 18 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=0.9
+ $X2=7.01 $Y2=0.9
r55 17 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.705 $Y=0.9
+ $X2=7.87 $Y2=0.9
r56 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.705 $Y=0.9
+ $X2=7.175 $Y2=0.9
r57 14 22 1.75975 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.9 $Y=0.92
+ $X2=4.775 $Y2=0.92
r58 14 16 37.2338 $w=2.08e-07 $l=7.05e-07 $layer=LI1_cond $X=4.9 $Y=0.92
+ $X2=5.605 $Y2=0.92
r59 13 28 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=6.845 $Y=0.92
+ $X2=7.01 $Y2=0.92
r60 13 16 65.4892 $w=2.08e-07 $l=1.24e-06 $layer=LI1_cond $X=6.845 $Y=0.92
+ $X2=5.605 $Y2=0.92
r61 4 31 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=7.73
+ $Y=0.325 $X2=7.87 $Y2=0.7
r62 3 25 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=6.87
+ $Y=0.325 $X2=7.01 $Y2=0.7
r63 2 16 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.465
+ $Y=0.325 $X2=5.605 $Y2=0.92
r64 1 20 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=4.605
+ $Y=0.325 $X2=4.745 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_4%A_1291_65# 1 2 3 4 5 16 18 24 28 30 34 36 41
+ 46
c61 41 0 3.03292e-19 $X=7.44 $Y=0.34
c62 28 0 1.81325e-19 $X=9.16 $Y=0.48
r63 41 44 8.17225 $w=1.88e-07 $l=1.4e-07 $layer=LI1_cond $X=7.44 $Y=0.34
+ $X2=7.44 $Y2=0.48
r64 36 39 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=6.575 $Y=0.34
+ $X2=6.575 $Y2=0.48
r65 32 34 16.8434 $w=2.58e-07 $l=3.8e-07 $layer=LI1_cond $X=10.055 $Y=0.86
+ $X2=10.055 $Y2=0.48
r66 31 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.255 $Y=0.945
+ $X2=9.16 $Y2=0.945
r67 30 32 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.925 $Y=0.945
+ $X2=10.055 $Y2=0.86
r68 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.925 $Y=0.945
+ $X2=9.255 $Y2=0.945
r69 26 46 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.16 $Y=0.86
+ $X2=9.16 $Y2=0.945
r70 26 28 22.1818 $w=1.88e-07 $l=3.8e-07 $layer=LI1_cond $X=9.16 $Y=0.86
+ $X2=9.16 $Y2=0.48
r71 24 46 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=9.065 $Y=0.945
+ $X2=9.16 $Y2=0.945
r72 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.065 $Y=0.945
+ $X2=8.395 $Y2=0.945
r73 21 25 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=8.305 $Y=0.86
+ $X2=8.395 $Y2=0.945
r74 21 23 24.0303 $w=1.78e-07 $l=3.9e-07 $layer=LI1_cond $X=8.305 $Y=0.86
+ $X2=8.305 $Y2=0.47
r75 20 23 2.77273 $w=1.78e-07 $l=4.5e-08 $layer=LI1_cond $X=8.305 $Y=0.425
+ $X2=8.305 $Y2=0.47
r76 19 41 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.535 $Y=0.34 $X2=7.44
+ $Y2=0.34
r77 18 20 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=8.215 $Y=0.34
+ $X2=8.305 $Y2=0.425
r78 18 19 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.215 $Y=0.34
+ $X2=7.535 $Y2=0.34
r79 17 36 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=6.675 $Y=0.34 $X2=6.575
+ $Y2=0.34
r80 16 41 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.345 $Y=0.34 $X2=7.44
+ $Y2=0.34
r81 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.345 $Y=0.34
+ $X2=6.675 $Y2=0.34
r82 5 34 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=9.88
+ $Y=0.325 $X2=10.02 $Y2=0.48
r83 4 28 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=9.02
+ $Y=0.325 $X2=9.16 $Y2=0.48
r84 3 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.16
+ $Y=0.325 $X2=8.3 $Y2=0.47
r85 2 44 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=7.3
+ $Y=0.325 $X2=7.44 $Y2=0.48
r86 1 39 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=6.455
+ $Y=0.325 $X2=6.58 $Y2=0.48
.ends

