* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor2_1 A B VGND VNB VPB VPWR Y
M1000 a_302_47# B VGND VNB nshort w=840000u l=150000u
+  ad=5.124e+11p pd=4.58e+06u as=5.502e+11p ps=4.67e+06u
M1001 Y B a_385_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.347e+11p pd=3.21e+06u as=4.914e+11p ps=3.3e+06u
M1002 a_33_47# B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.6317e+12p ps=1.015e+07u
M1003 Y a_33_47# a_302_47# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1004 a_116_47# B a_33_47# VNB nshort w=840000u l=150000u
+  ad=2.058e+11p pd=2.17e+06u as=2.226e+11p ps=2.21e+06u
M1005 VPWR a_33_47# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_33_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_116_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_385_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A a_302_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
