* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o22a_0 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 VGND a_80_313# X VNB nshort w=420000u l=150000u
+  ad=4.179e+11p pd=3.67e+06u as=1.113e+11p ps=1.37e+06u
M1001 a_80_313# B2 a_372_489# VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=1.536e+11p ps=1.76e+06u
M1002 a_286_125# A1 VGND VNB nshort w=420000u l=150000u
+  ad=2.688e+11p pd=2.96e+06u as=0p ps=0u
M1003 a_80_313# B1 a_286_125# VNB nshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1004 a_286_125# B2 a_80_313# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A1 a_536_489# VPB phighvt w=640000u l=150000u
+  ad=9.12e+11p pd=5.41e+06u as=2.432e+11p ps=2.04e+06u
M1006 VPWR a_80_313# X VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1007 a_372_489# B1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_286_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_536_489# A2 a_80_313# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
