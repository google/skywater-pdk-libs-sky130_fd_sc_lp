* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2111ai_lp A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 Y A2 a_483_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_483_409# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_167_57# C1 a_245_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_245_57# B1 a_347_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_347_57# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 Y D1 a_167_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VGND A1 a_347_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
