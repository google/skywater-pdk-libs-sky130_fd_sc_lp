* File: sky130_fd_sc_lp__mux2_8.pxi.spice
* Created: Wed Sep  2 10:00:26 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2_8%A_84_21# N_A_84_21#_M1016_s N_A_84_21#_M1008_s
+ N_A_84_21#_M1002_s N_A_84_21#_M1017_d N_A_84_21#_M1004_g N_A_84_21#_M1006_g
+ N_A_84_21#_M1005_g N_A_84_21#_M1012_g N_A_84_21#_M1009_g N_A_84_21#_M1015_g
+ N_A_84_21#_M1011_g N_A_84_21#_M1021_g N_A_84_21#_M1014_g N_A_84_21#_M1022_g
+ N_A_84_21#_M1025_g N_A_84_21#_M1024_g N_A_84_21#_M1031_g N_A_84_21#_M1027_g
+ N_A_84_21#_M1032_g N_A_84_21#_M1033_g N_A_84_21#_c_306_p N_A_84_21#_c_177_n
+ N_A_84_21#_c_178_n N_A_84_21#_c_179_n N_A_84_21#_c_255_p N_A_84_21#_c_180_n
+ N_A_84_21#_c_195_p N_A_84_21#_c_181_n N_A_84_21#_c_215_p N_A_84_21#_c_199_p
+ N_A_84_21#_c_222_p N_A_84_21#_c_201_p N_A_84_21#_c_210_p N_A_84_21#_c_200_p
+ N_A_84_21#_c_204_p N_A_84_21#_c_246_p N_A_84_21#_c_237_p N_A_84_21#_c_202_p
+ N_A_84_21#_c_226_p N_A_84_21#_c_218_p PM_SKY130_FD_SC_LP__MUX2_8%A_84_21#
x_PM_SKY130_FD_SC_LP__MUX2_8%S N_S_M1010_g N_S_M1007_g N_S_M1018_g N_S_M1023_g
+ N_S_M1030_g N_S_M1000_g N_S_c_452_n N_S_c_453_n N_S_c_463_n N_S_c_464_n
+ N_S_c_454_n N_S_c_455_n N_S_c_467_n N_S_c_499_n N_S_c_558_p N_S_c_559_p S
+ N_S_c_456_n N_S_c_457_n N_S_c_470_n PM_SKY130_FD_SC_LP__MUX2_8%S
x_PM_SKY130_FD_SC_LP__MUX2_8%A1 N_A1_M1016_g N_A1_c_631_n N_A1_M1019_g
+ N_A1_M1017_g N_A1_M1026_g N_A1_c_633_n N_A1_c_634_n N_A1_c_635_n N_A1_c_636_n
+ N_A1_c_637_n N_A1_c_638_n A1 N_A1_c_640_n N_A1_c_641_n
+ PM_SKY130_FD_SC_LP__MUX2_8%A1
x_PM_SKY130_FD_SC_LP__MUX2_8%A0 N_A0_M1002_g N_A0_M1028_g N_A0_M1008_g
+ N_A0_M1029_g N_A0_c_753_n N_A0_c_754_n N_A0_c_755_n N_A0_c_756_n N_A0_c_757_n
+ A0 N_A0_c_758_n N_A0_c_759_n PM_SKY130_FD_SC_LP__MUX2_8%A0
x_PM_SKY130_FD_SC_LP__MUX2_8%A_1179_311# N_A_1179_311#_M1030_d
+ N_A_1179_311#_M1000_d N_A_1179_311#_M1001_g N_A_1179_311#_M1003_g
+ N_A_1179_311#_M1020_g N_A_1179_311#_M1013_g N_A_1179_311#_c_856_n
+ N_A_1179_311#_c_857_n N_A_1179_311#_c_877_n N_A_1179_311#_c_879_n
+ N_A_1179_311#_c_858_n N_A_1179_311#_c_912_n N_A_1179_311#_c_859_n
+ N_A_1179_311#_c_860_n N_A_1179_311#_c_861_n N_A_1179_311#_c_869_n
+ N_A_1179_311#_c_924_n N_A_1179_311#_c_862_n N_A_1179_311#_c_863_n
+ N_A_1179_311#_c_880_n N_A_1179_311#_c_870_n
+ PM_SKY130_FD_SC_LP__MUX2_8%A_1179_311#
x_PM_SKY130_FD_SC_LP__MUX2_8%VPWR N_VPWR_M1006_s N_VPWR_M1012_s N_VPWR_M1021_s
+ N_VPWR_M1024_s N_VPWR_M1032_s N_VPWR_M1023_d N_VPWR_M1013_d N_VPWR_c_1006_n
+ N_VPWR_c_1007_n N_VPWR_c_1008_n N_VPWR_c_1009_n N_VPWR_c_1010_n
+ N_VPWR_c_1011_n N_VPWR_c_1012_n N_VPWR_c_1013_n N_VPWR_c_1014_n
+ N_VPWR_c_1015_n N_VPWR_c_1016_n N_VPWR_c_1017_n N_VPWR_c_1018_n
+ N_VPWR_c_1019_n N_VPWR_c_1020_n VPWR N_VPWR_c_1021_n N_VPWR_c_1022_n
+ N_VPWR_c_1023_n N_VPWR_c_1005_n N_VPWR_c_1025_n N_VPWR_c_1026_n
+ N_VPWR_c_1027_n PM_SKY130_FD_SC_LP__MUX2_8%VPWR
x_PM_SKY130_FD_SC_LP__MUX2_8%X N_X_M1004_s N_X_M1009_s N_X_M1014_s N_X_M1027_s
+ N_X_M1006_d N_X_M1015_d N_X_M1022_d N_X_M1031_d N_X_c_1159_n N_X_c_1162_n
+ N_X_c_1148_n N_X_c_1153_n N_X_c_1173_n N_X_c_1177_n N_X_c_1149_n N_X_c_1154_n
+ N_X_c_1189_n N_X_c_1193_n N_X_c_1150_n N_X_c_1155_n N_X_c_1156_n N_X_c_1210_n
+ N_X_c_1212_n N_X_c_1215_n N_X_c_1217_n N_X_c_1151_n N_X_c_1157_n N_X_c_1152_n
+ N_X_c_1158_n X X PM_SKY130_FD_SC_LP__MUX2_8%X
x_PM_SKY130_FD_SC_LP__MUX2_8%A_843_419# N_A_843_419#_M1007_s
+ N_A_843_419#_M1028_d N_A_843_419#_c_1286_n N_A_843_419#_c_1290_n
+ N_A_843_419#_c_1291_n PM_SKY130_FD_SC_LP__MUX2_8%A_843_419#
x_PM_SKY130_FD_SC_LP__MUX2_8%A_1243_419# N_A_1243_419#_M1003_s
+ N_A_1243_419#_M1026_s N_A_1243_419#_c_1308_n N_A_1243_419#_c_1311_n
+ N_A_1243_419#_c_1312_n PM_SKY130_FD_SC_LP__MUX2_8%A_1243_419#
x_PM_SKY130_FD_SC_LP__MUX2_8%VGND N_VGND_M1004_d N_VGND_M1005_d N_VGND_M1011_d
+ N_VGND_M1025_d N_VGND_M1033_d N_VGND_M1018_d N_VGND_M1020_d N_VGND_c_1334_n
+ N_VGND_c_1335_n N_VGND_c_1336_n N_VGND_c_1337_n N_VGND_c_1338_n
+ N_VGND_c_1339_n N_VGND_c_1340_n N_VGND_c_1341_n N_VGND_c_1342_n
+ N_VGND_c_1343_n N_VGND_c_1344_n N_VGND_c_1345_n N_VGND_c_1346_n
+ N_VGND_c_1347_n N_VGND_c_1348_n N_VGND_c_1349_n N_VGND_c_1350_n
+ N_VGND_c_1351_n VGND N_VGND_c_1352_n N_VGND_c_1353_n N_VGND_c_1354_n
+ N_VGND_c_1355_n PM_SKY130_FD_SC_LP__MUX2_8%VGND
x_PM_SKY130_FD_SC_LP__MUX2_8%A_839_47# N_A_839_47#_M1010_s N_A_839_47#_M1019_d
+ N_A_839_47#_c_1465_n N_A_839_47#_c_1469_n N_A_839_47#_c_1471_n
+ PM_SKY130_FD_SC_LP__MUX2_8%A_839_47#
x_PM_SKY130_FD_SC_LP__MUX2_8%A_1243_47# N_A_1243_47#_M1001_s
+ N_A_1243_47#_M1029_d N_A_1243_47#_c_1488_n N_A_1243_47#_c_1496_n
+ PM_SKY130_FD_SC_LP__MUX2_8%A_1243_47#
cc_1 VNB N_A_84_21#_M1004_g 0.0266656f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_2 VNB N_A_84_21#_M1006_g 0.0045013f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_3 VNB N_A_84_21#_M1005_g 0.0193485f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_4 VNB N_A_84_21#_M1012_g 0.00275385f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_5 VNB N_A_84_21#_M1009_g 0.0200385f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_6 VNB N_A_84_21#_M1015_g 0.0029962f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=2.465
cc_7 VNB N_A_84_21#_M1011_g 0.0200684f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.655
cc_8 VNB N_A_84_21#_M1021_g 0.00300052f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=2.465
cc_9 VNB N_A_84_21#_M1014_g 0.0200684f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.655
cc_10 VNB N_A_84_21#_M1022_g 0.00300052f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_11 VNB N_A_84_21#_M1025_g 0.0209398f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_12 VNB N_A_84_21#_M1024_g 0.00300052f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_13 VNB N_A_84_21#_M1031_g 0.0029978f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=2.465
cc_14 VNB N_A_84_21#_M1027_g 0.0209398f $X=-0.19 $Y=-0.245 $X2=3.145 $Y2=0.655
cc_15 VNB N_A_84_21#_M1032_g 0.00338868f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=2.465
cc_16 VNB N_A_84_21#_M1033_g 0.0218215f $X=-0.19 $Y=-0.245 $X2=3.575 $Y2=0.655
cc_17 VNB N_A_84_21#_c_177_n 0.185654f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.43
cc_18 VNB N_A_84_21#_c_178_n 9.35817e-19 $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=2.32
cc_19 VNB N_A_84_21#_c_179_n 0.0130477f $X=-0.19 $Y=-0.245 $X2=4.135 $Y2=1.35
cc_20 VNB N_A_84_21#_c_180_n 0.00287554f $X=-0.19 $Y=-0.245 $X2=4.22 $Y2=1.265
cc_21 VNB N_A_84_21#_c_181_n 0.00478382f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.43
cc_22 VNB N_S_M1010_g 0.0504336f $X=-0.19 $Y=-0.245 $X2=4.715 $Y2=2.095
cc_23 VNB N_S_M1018_g 0.0542323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_S_M1030_g 0.0347745f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_25 VNB N_S_c_452_n 0.00209806f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_26 VNB N_S_c_453_n 0.0102347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_S_c_454_n 0.0158916f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.655
cc_28 VNB N_S_c_455_n 0.0291197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_S_c_456_n 0.0112984f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_30 VNB N_S_c_457_n 0.00226315f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_31 VNB N_A1_M1016_g 0.0192718f $X=-0.19 $Y=-0.245 $X2=4.715 $Y2=2.095
cc_32 VNB N_A1_c_631_n 0.0157642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A1_M1019_g 0.0200288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A1_c_633_n 0.00372212f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.265
cc_35 VNB N_A1_c_634_n 0.0115843f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_36 VNB N_A1_c_635_n 0.0015019f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_37 VNB N_A1_c_636_n 0.00573365f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_38 VNB N_A1_c_637_n 0.00410544f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.655
cc_39 VNB N_A1_c_638_n 0.00545627f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=2.465
cc_40 VNB A1 0.00359107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A1_c_640_n 0.0325856f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.595
cc_42 VNB N_A1_c_641_n 0.00239171f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_43 VNB N_A0_M1008_g 0.0185461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A0_M1029_g 0.019262f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_45 VNB N_A0_c_753_n 0.0245687f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_46 VNB N_A0_c_754_n 3.10606e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A0_c_755_n 0.00199874f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_48 VNB N_A0_c_756_n 0.0122654f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_49 VNB N_A0_c_757_n 0.00758593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A0_c_758_n 0.0425087f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.595
cc_51 VNB N_A0_c_759_n 0.00372931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1179_311#_M1001_g 0.056247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1179_311#_M1020_g 0.0291228f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.595
cc_54 VNB N_A_1179_311#_M1013_g 0.00857867f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.265
cc_55 VNB N_A_1179_311#_c_856_n 0.0021491f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.595
cc_56 VNB N_A_1179_311#_c_857_n 0.012187f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_57 VNB N_A_1179_311#_c_858_n 0.00246339f $X=-0.19 $Y=-0.245 $X2=1.355
+ $Y2=1.595
cc_58 VNB N_A_1179_311#_c_859_n 0.0178024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1179_311#_c_860_n 0.00569276f $X=-0.19 $Y=-0.245 $X2=1.785
+ $Y2=1.265
cc_60 VNB N_A_1179_311#_c_861_n 0.0285788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1179_311#_c_862_n 0.0393299f $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=2.465
cc_62 VNB N_A_1179_311#_c_863_n 6.68563e-19 $X=-0.19 $Y=-0.245 $X2=2.215
+ $Y2=2.465
cc_63 VNB N_VPWR_c_1005_n 0.362705f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=2.405
cc_64 VNB N_X_c_1148_n 0.00462709f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.595
cc_65 VNB N_X_c_1149_n 0.00225436f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.265
cc_66 VNB N_X_c_1150_n 0.00497918f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.595
cc_67 VNB N_X_c_1151_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=3.575 $Y2=0.655
cc_68 VNB N_X_c_1152_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=3.625 $Y2=1.43
cc_69 VNB N_VGND_c_1334_n 0.0108703f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_70 VNB N_VGND_c_1335_n 0.0427456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1336_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1337_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1338_n 0.00513283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1339_n 0.00902567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1340_n 0.00529596f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.655
cc_76 VNB N_VGND_c_1341_n 0.00558649f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_77 VNB N_VGND_c_1342_n 0.0187217f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.265
cc_78 VNB N_VGND_c_1343_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.655
cc_79 VNB N_VGND_c_1344_n 0.0190399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1345_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.595
cc_81 VNB N_VGND_c_1346_n 0.0190399f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.465
cc_82 VNB N_VGND_c_1347_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1348_n 0.0187217f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=2.465
cc_84 VNB N_VGND_c_1349_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=2.465
cc_85 VNB N_VGND_c_1350_n 0.0409355f $X=-0.19 $Y=-0.245 $X2=3.145 $Y2=1.265
cc_86 VNB N_VGND_c_1351_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=3.145 $Y2=0.655
cc_87 VNB N_VGND_c_1352_n 0.0409333f $X=-0.19 $Y=-0.245 $X2=3.585 $Y2=1.43
cc_88 VNB N_VGND_c_1353_n 0.0194586f $X=-0.19 $Y=-0.245 $X2=4.225 $Y2=2.49
cc_89 VNB N_VGND_c_1354_n 0.4103f $X=-0.19 $Y=-0.245 $X2=4.67 $Y2=0.77
cc_90 VNB N_VGND_c_1355_n 0.00631736f $X=-0.19 $Y=-0.245 $X2=6.69 $Y2=2.52
cc_91 VPB N_A_84_21#_M1006_g 0.0259807f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_92 VPB N_A_84_21#_M1012_g 0.0189284f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_93 VPB N_A_84_21#_M1015_g 0.0195815f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_94 VPB N_A_84_21#_M1021_g 0.0196107f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_95 VPB N_A_84_21#_M1022_g 0.0196107f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.465
cc_96 VPB N_A_84_21#_M1024_g 0.0196107f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_97 VPB N_A_84_21#_M1031_g 0.0196033f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=2.465
cc_98 VPB N_A_84_21#_M1032_g 0.02163f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=2.465
cc_99 VPB N_A_84_21#_c_178_n 0.00305999f $X=-0.19 $Y=1.655 $X2=3.71 $Y2=2.32
cc_100 VPB N_S_M1007_g 0.0201295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_S_M1023_g 0.0221262f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.655
cc_102 VPB N_S_M1000_g 0.0272497f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_103 VPB N_S_c_452_n 0.00270499f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_104 VPB N_S_c_453_n 0.0253392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_S_c_463_n 0.00527619f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=0.655
cc_106 VPB N_S_c_464_n 0.00465461f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=0.655
cc_107 VPB N_S_c_454_n 0.00138909f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=0.655
cc_108 VPB N_S_c_455_n 0.00653614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_S_c_467_n 0.0164108f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_110 VPB N_S_c_456_n 0.0198547f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=0.655
cc_111 VPB N_S_c_457_n 0.00286907f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=0.655
cc_112 VPB N_S_c_470_n 0.00314257f $X=-0.19 $Y=1.655 $X2=3.145 $Y2=0.655
cc_113 VPB N_A1_M1017_g 0.01914f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.265
cc_114 VPB N_A1_M1026_g 0.02001f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.595
cc_115 VPB N_A1_c_634_n 0.0357456f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_116 VPB N_A1_c_636_n 0.005065f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=0.655
cc_117 VPB N_A1_c_637_n 0.00209101f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=0.655
cc_118 VPB N_A1_c_638_n 0.00108472f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_119 VPB A1 4.09789e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A1_c_641_n 0.00231119f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.465
cc_121 VPB N_A0_M1002_g 0.02095f $X=-0.19 $Y=1.655 $X2=4.715 $Y2=2.095
cc_122 VPB N_A0_M1028_g 0.0215829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A0_c_755_n 8.25483e-19 $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_124 VPB N_A0_c_756_n 0.0279903f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_125 VPB N_A_1179_311#_M1003_g 0.0217826f $X=-0.19 $Y=1.655 $X2=0.495
+ $Y2=1.265
cc_126 VPB N_A_1179_311#_M1013_g 0.0352167f $X=-0.19 $Y=1.655 $X2=0.925
+ $Y2=1.265
cc_127 VPB N_A_1179_311#_c_856_n 0.00101988f $X=-0.19 $Y=1.655 $X2=0.925
+ $Y2=1.595
cc_128 VPB N_A_1179_311#_c_857_n 0.0214125f $X=-0.19 $Y=1.655 $X2=0.925
+ $Y2=2.465
cc_129 VPB N_A_1179_311#_c_858_n 0.00398544f $X=-0.19 $Y=1.655 $X2=1.355
+ $Y2=1.595
cc_130 VPB N_A_1179_311#_c_869_n 0.0179193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_1179_311#_c_870_n 0.0286347f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_1006_n 0.0106521f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=0.655
cc_133 VPB N_VPWR_c_1007_n 0.0575933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_1008_n 0.0047158f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=0.655
cc_135 VPB N_VPWR_c_1009_n 0.0047158f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_136 VPB N_VPWR_c_1010_n 0.00412866f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=0.655
cc_137 VPB N_VPWR_c_1011_n 0.0158404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_1012_n 0.00276924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_1013_n 0.00552942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_1014_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_1015_n 0.0185788f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=0.655
cc_142 VPB N_VPWR_c_1016_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_1017_n 0.0185788f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_144 VPB N_VPWR_c_1018_n 0.00324402f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_145 VPB N_VPWR_c_1019_n 0.0185788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_1020_n 0.00324402f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=1.595
cc_147 VPB N_VPWR_c_1021_n 0.0432928f $X=-0.19 $Y=1.655 $X2=3.575 $Y2=0.655
cc_148 VPB N_VPWR_c_1022_n 0.0411748f $X=-0.19 $Y=1.655 $X2=3.585 $Y2=1.43
cc_149 VPB N_VPWR_c_1023_n 0.0167428f $X=-0.19 $Y=1.655 $X2=4.055 $Y2=2.405
cc_150 VPB N_VPWR_c_1005_n 0.0471789f $X=-0.19 $Y=1.655 $X2=3.795 $Y2=2.405
cc_151 VPB N_VPWR_c_1025_n 0.00510842f $X=-0.19 $Y=1.655 $X2=4.305 $Y2=0.77
cc_152 VPB N_VPWR_c_1026_n 0.00631288f $X=-0.19 $Y=1.655 $X2=5.69 $Y2=2.49
cc_153 VPB N_VPWR_c_1027_n 0.00510842f $X=-0.19 $Y=1.655 $X2=5.86 $Y2=2.52
cc_154 VPB N_X_c_1153_n 0.00476412f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_155 VPB N_X_c_1154_n 0.00248004f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=0.655
cc_156 VPB N_X_c_1155_n 0.00248004f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_157 VPB N_X_c_1156_n 0.00213175f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=1.595
cc_158 VPB N_X_c_1157_n 0.0025378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_X_c_1158_n 0.0025378f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=1.43
cc_160 N_A_84_21#_M1033_g N_S_M1010_g 0.0208288f $X=3.575 $Y=0.655 $X2=0 $Y2=0
cc_161 N_A_84_21#_c_177_n N_S_M1010_g 0.0134352f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_162 N_A_84_21#_c_179_n N_S_M1010_g 0.012326f $X=4.135 $Y=1.35 $X2=0 $Y2=0
cc_163 N_A_84_21#_c_180_n N_S_M1010_g 0.00930327f $X=4.22 $Y=1.265 $X2=0 $Y2=0
cc_164 N_A_84_21#_c_195_p N_S_M1010_g 0.00541266f $X=4.305 $Y=0.77 $X2=0 $Y2=0
cc_165 N_A_84_21#_c_181_n N_S_M1010_g 0.0040336f $X=3.71 $Y=1.43 $X2=0 $Y2=0
cc_166 N_A_84_21#_M1032_g N_S_M1007_g 0.0204173f $X=3.505 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A_84_21#_c_178_n N_S_M1007_g 0.00315303f $X=3.71 $Y=2.32 $X2=0 $Y2=0
cc_168 N_A_84_21#_c_199_p N_S_M1007_g 0.0153519f $X=4.225 $Y=2.447 $X2=0 $Y2=0
cc_169 N_A_84_21#_c_200_p N_S_M1007_g 7.08042e-19 $X=5.02 $Y=2.57 $X2=0 $Y2=0
cc_170 N_A_84_21#_c_201_p N_S_M1018_g 3.64956e-19 $X=5 $Y=0.725 $X2=0 $Y2=0
cc_171 N_A_84_21#_c_202_p N_S_M1018_g 0.0128833f $X=6.62 $Y=0.745 $X2=0 $Y2=0
cc_172 N_A_84_21#_c_200_p N_S_M1023_g 6.61941e-19 $X=5.02 $Y=2.57 $X2=0 $Y2=0
cc_173 N_A_84_21#_c_204_p N_S_M1023_g 0.0128531f $X=5.69 $Y=2.505 $X2=0 $Y2=0
cc_174 N_A_84_21#_c_178_n N_S_c_452_n 0.029564f $X=3.71 $Y=2.32 $X2=0 $Y2=0
cc_175 N_A_84_21#_c_179_n N_S_c_452_n 0.0277197f $X=4.135 $Y=1.35 $X2=0 $Y2=0
cc_176 N_A_84_21#_M1032_g N_S_c_453_n 0.00674947f $X=3.505 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A_84_21#_c_178_n N_S_c_453_n 0.00101973f $X=3.71 $Y=2.32 $X2=0 $Y2=0
cc_178 N_A_84_21#_c_179_n N_S_c_453_n 0.00100181f $X=4.135 $Y=1.35 $X2=0 $Y2=0
cc_179 N_A_84_21#_c_210_p N_S_c_453_n 3.56001e-19 $X=4.69 $Y=2.57 $X2=0 $Y2=0
cc_180 N_A_84_21#_M1002_s N_S_c_463_n 0.00176891f $X=4.715 $Y=2.095 $X2=0 $Y2=0
cc_181 N_A_84_21#_c_210_p N_S_c_463_n 0.0441016f $X=4.69 $Y=2.57 $X2=0 $Y2=0
cc_182 N_A_84_21#_c_204_p N_S_c_463_n 0.0170403f $X=5.69 $Y=2.505 $X2=0 $Y2=0
cc_183 N_A_84_21#_c_178_n N_S_c_464_n 0.0166323f $X=3.71 $Y=2.32 $X2=0 $Y2=0
cc_184 N_A_84_21#_c_215_p N_S_c_464_n 0.0149829f $X=4.055 $Y=2.447 $X2=0 $Y2=0
cc_185 N_A_84_21#_c_210_p N_S_c_464_n 0.0153281f $X=4.69 $Y=2.57 $X2=0 $Y2=0
cc_186 N_A_84_21#_c_204_p N_S_c_467_n 0.00717099f $X=5.69 $Y=2.505 $X2=0 $Y2=0
cc_187 N_A_84_21#_c_218_p N_S_c_467_n 0.00728987f $X=6.69 $Y=2.585 $X2=0 $Y2=0
cc_188 N_A_84_21#_c_204_p N_S_c_499_n 0.0017036f $X=5.69 $Y=2.505 $X2=0 $Y2=0
cc_189 N_A_84_21#_c_204_p N_S_c_456_n 3.99127e-19 $X=5.69 $Y=2.505 $X2=0 $Y2=0
cc_190 N_A_84_21#_c_180_n N_A1_M1016_g 0.00507892f $X=4.22 $Y=1.265 $X2=0 $Y2=0
cc_191 N_A_84_21#_c_222_p N_A1_M1016_g 0.0112111f $X=4.67 $Y=0.725 $X2=0 $Y2=0
cc_192 N_A_84_21#_c_201_p N_A1_M1019_g 0.00277056f $X=5 $Y=0.725 $X2=0 $Y2=0
cc_193 N_A_84_21#_c_202_p N_A1_M1019_g 0.00809622f $X=6.62 $Y=0.745 $X2=0 $Y2=0
cc_194 N_A_84_21#_c_218_p N_A1_M1017_g 0.0113748f $X=6.69 $Y=2.585 $X2=0 $Y2=0
cc_195 N_A_84_21#_c_226_p N_A1_M1026_g 0.00567885f $X=6.855 $Y=2.585 $X2=0 $Y2=0
cc_196 N_A_84_21#_c_179_n N_A1_c_635_n 0.0143085f $X=4.135 $Y=1.35 $X2=0 $Y2=0
cc_197 N_A_84_21#_c_180_n N_A1_c_635_n 0.018f $X=4.22 $Y=1.265 $X2=0 $Y2=0
cc_198 N_A_84_21#_c_222_p N_A1_c_635_n 0.0229349f $X=4.67 $Y=0.725 $X2=0 $Y2=0
cc_199 N_A_84_21#_c_181_n N_A1_c_637_n 0.00165463f $X=3.71 $Y=1.43 $X2=0 $Y2=0
cc_200 N_A_84_21#_c_179_n N_A1_c_640_n 6.34751e-19 $X=4.135 $Y=1.35 $X2=0 $Y2=0
cc_201 N_A_84_21#_c_201_p N_A1_c_640_n 0.00355137f $X=5 $Y=0.725 $X2=0 $Y2=0
cc_202 N_A_84_21#_c_210_p N_A0_M1002_g 0.00840566f $X=4.69 $Y=2.57 $X2=0 $Y2=0
cc_203 N_A_84_21#_c_200_p N_A0_M1002_g 0.00413557f $X=5.02 $Y=2.57 $X2=0 $Y2=0
cc_204 N_A_84_21#_c_200_p N_A0_M1028_g 0.00415376f $X=5.02 $Y=2.57 $X2=0 $Y2=0
cc_205 N_A_84_21#_c_204_p N_A0_M1028_g 0.00839198f $X=5.69 $Y=2.505 $X2=0 $Y2=0
cc_206 N_A_84_21#_c_237_p N_A0_M1008_g 0.00194187f $X=6.785 $Y=0.725 $X2=0 $Y2=0
cc_207 N_A_84_21#_c_202_p N_A0_M1008_g 0.00754223f $X=6.62 $Y=0.745 $X2=0 $Y2=0
cc_208 N_A_84_21#_c_237_p N_A0_M1029_g 0.0030989f $X=6.785 $Y=0.725 $X2=0 $Y2=0
cc_209 N_A_84_21#_c_202_p N_A0_c_753_n 0.102845f $X=6.62 $Y=0.745 $X2=0 $Y2=0
cc_210 N_A_84_21#_c_201_p N_A0_c_754_n 0.0123464f $X=5 $Y=0.725 $X2=0 $Y2=0
cc_211 N_A_84_21#_c_237_p N_A0_c_758_n 0.00111102f $X=6.785 $Y=0.725 $X2=0 $Y2=0
cc_212 N_A_84_21#_c_237_p N_A0_c_759_n 0.0117826f $X=6.785 $Y=0.725 $X2=0 $Y2=0
cc_213 N_A_84_21#_c_237_p N_A_1179_311#_M1001_g 2.39364e-19 $X=6.785 $Y=0.725
+ $X2=0 $Y2=0
cc_214 N_A_84_21#_c_202_p N_A_1179_311#_M1001_g 0.0125429f $X=6.62 $Y=0.745
+ $X2=0 $Y2=0
cc_215 N_A_84_21#_c_246_p N_A_1179_311#_M1003_g 8.04884e-19 $X=5.86 $Y=2.505
+ $X2=0 $Y2=0
cc_216 N_A_84_21#_c_218_p N_A_1179_311#_M1003_g 0.0124616f $X=6.69 $Y=2.585
+ $X2=0 $Y2=0
cc_217 N_A_84_21#_c_226_p N_A_1179_311#_M1013_g 8.6575e-19 $X=6.855 $Y=2.585
+ $X2=0 $Y2=0
cc_218 N_A_84_21#_c_218_p N_A_1179_311#_c_857_n 4.95835e-19 $X=6.69 $Y=2.585
+ $X2=0 $Y2=0
cc_219 N_A_84_21#_M1017_d N_A_1179_311#_c_877_n 0.0036337f $X=6.645 $Y=2.095
+ $X2=0 $Y2=0
cc_220 N_A_84_21#_c_218_p N_A_1179_311#_c_877_n 0.0410555f $X=6.69 $Y=2.585
+ $X2=0 $Y2=0
cc_221 N_A_84_21#_c_218_p N_A_1179_311#_c_879_n 0.0161517f $X=6.69 $Y=2.585
+ $X2=0 $Y2=0
cc_222 N_A_84_21#_c_226_p N_A_1179_311#_c_880_n 0.00245416f $X=6.855 $Y=2.585
+ $X2=0 $Y2=0
cc_223 N_A_84_21#_c_178_n N_VPWR_M1032_s 0.00923756f $X=3.71 $Y=2.32 $X2=0 $Y2=0
cc_224 N_A_84_21#_c_255_p N_VPWR_M1032_s 0.00313243f $X=3.795 $Y=2.405 $X2=0
+ $Y2=0
cc_225 N_A_84_21#_c_215_p N_VPWR_M1032_s 0.0111488f $X=4.055 $Y=2.447 $X2=0
+ $Y2=0
cc_226 N_A_84_21#_c_246_p N_VPWR_M1023_d 0.00483864f $X=5.86 $Y=2.505 $X2=0
+ $Y2=0
cc_227 N_A_84_21#_c_218_p N_VPWR_M1023_d 0.00335513f $X=6.69 $Y=2.585 $X2=0
+ $Y2=0
cc_228 N_A_84_21#_M1006_g N_VPWR_c_1007_n 0.00941302f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_229 N_A_84_21#_M1012_g N_VPWR_c_1008_n 0.00372815f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_230 N_A_84_21#_M1015_g N_VPWR_c_1008_n 0.00372815f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_231 N_A_84_21#_M1021_g N_VPWR_c_1009_n 0.00372815f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_232 N_A_84_21#_M1022_g N_VPWR_c_1009_n 0.00372815f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_233 N_A_84_21#_M1024_g N_VPWR_c_1010_n 0.00372815f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_234 N_A_84_21#_M1031_g N_VPWR_c_1010_n 0.00242144f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_235 N_A_84_21#_M1031_g N_VPWR_c_1011_n 0.0054895f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_236 N_A_84_21#_M1032_g N_VPWR_c_1011_n 0.00486043f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_237 N_A_84_21#_M1031_g N_VPWR_c_1012_n 6.3078e-19 $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_238 N_A_84_21#_M1032_g N_VPWR_c_1012_n 0.0106757f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A_84_21#_c_255_p N_VPWR_c_1012_n 0.0138594f $X=3.795 $Y=2.405 $X2=0
+ $Y2=0
cc_240 N_A_84_21#_c_215_p N_VPWR_c_1012_n 0.00704757f $X=4.055 $Y=2.447 $X2=0
+ $Y2=0
cc_241 N_A_84_21#_c_246_p N_VPWR_c_1013_n 0.0240343f $X=5.86 $Y=2.505 $X2=0
+ $Y2=0
cc_242 N_A_84_21#_M1006_g N_VPWR_c_1015_n 0.0054895f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_243 N_A_84_21#_M1012_g N_VPWR_c_1015_n 0.0054895f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_244 N_A_84_21#_M1015_g N_VPWR_c_1017_n 0.0054895f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_245 N_A_84_21#_M1021_g N_VPWR_c_1017_n 0.0054895f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_246 N_A_84_21#_M1022_g N_VPWR_c_1019_n 0.0054895f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_A_84_21#_M1024_g N_VPWR_c_1019_n 0.0054895f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_248 N_A_84_21#_c_199_p N_VPWR_c_1021_n 0.00170233f $X=4.225 $Y=2.447 $X2=0
+ $Y2=0
cc_249 N_A_84_21#_c_204_p N_VPWR_c_1021_n 0.00190334f $X=5.69 $Y=2.505 $X2=0
+ $Y2=0
cc_250 N_A_84_21#_c_218_p N_VPWR_c_1022_n 0.00203818f $X=6.69 $Y=2.585 $X2=0
+ $Y2=0
cc_251 N_A_84_21#_M1002_s N_VPWR_c_1005_n 0.00225186f $X=4.715 $Y=2.095 $X2=0
+ $Y2=0
cc_252 N_A_84_21#_M1017_d N_VPWR_c_1005_n 0.00281482f $X=6.645 $Y=2.095 $X2=0
+ $Y2=0
cc_253 N_A_84_21#_M1006_g N_VPWR_c_1005_n 0.010744f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_254 N_A_84_21#_M1012_g N_VPWR_c_1005_n 0.00979301f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_255 N_A_84_21#_M1015_g N_VPWR_c_1005_n 0.00979301f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_256 N_A_84_21#_M1021_g N_VPWR_c_1005_n 0.00979301f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_A_84_21#_M1022_g N_VPWR_c_1005_n 0.00979301f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_258 N_A_84_21#_M1024_g N_VPWR_c_1005_n 0.00979301f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_259 N_A_84_21#_M1031_g N_VPWR_c_1005_n 0.00979301f $X=3.075 $Y=2.465 $X2=0
+ $Y2=0
cc_260 N_A_84_21#_M1032_g N_VPWR_c_1005_n 0.00824727f $X=3.505 $Y=2.465 $X2=0
+ $Y2=0
cc_261 N_A_84_21#_c_255_p N_VPWR_c_1005_n 6.15054e-19 $X=3.795 $Y=2.405 $X2=0
+ $Y2=0
cc_262 N_A_84_21#_c_215_p N_VPWR_c_1005_n 0.00617756f $X=4.055 $Y=2.447 $X2=0
+ $Y2=0
cc_263 N_A_84_21#_c_199_p N_VPWR_c_1005_n 0.00394036f $X=4.225 $Y=2.447 $X2=0
+ $Y2=0
cc_264 N_A_84_21#_c_204_p N_VPWR_c_1005_n 0.00476757f $X=5.69 $Y=2.505 $X2=0
+ $Y2=0
cc_265 N_A_84_21#_c_246_p N_VPWR_c_1005_n 0.00126439f $X=5.86 $Y=2.505 $X2=0
+ $Y2=0
cc_266 N_A_84_21#_c_218_p N_VPWR_c_1005_n 0.00489094f $X=6.69 $Y=2.585 $X2=0
+ $Y2=0
cc_267 N_A_84_21#_M1004_g N_X_c_1159_n 0.00886489f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_268 N_A_84_21#_M1005_g N_X_c_1159_n 0.00986698f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_269 N_A_84_21#_M1009_g N_X_c_1159_n 6.3694e-19 $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_270 N_A_84_21#_M1006_g N_X_c_1162_n 0.013885f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_271 N_A_84_21#_M1012_g N_X_c_1162_n 0.0144592f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A_84_21#_M1015_g N_X_c_1162_n 7.09394e-19 $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A_84_21#_M1005_g N_X_c_1148_n 0.0149371f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_274 N_A_84_21#_M1009_g N_X_c_1148_n 0.01115f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_275 N_A_84_21#_c_306_p N_X_c_1148_n 0.0209192f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_276 N_A_84_21#_c_177_n N_X_c_1148_n 0.00269643f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_277 N_A_84_21#_M1012_g N_X_c_1153_n 0.0149371f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_278 N_A_84_21#_M1015_g N_X_c_1153_n 0.0113972f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_279 N_A_84_21#_c_306_p N_X_c_1153_n 0.01715f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_280 N_A_84_21#_c_177_n N_X_c_1153_n 0.00258605f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_281 N_A_84_21#_M1005_g N_X_c_1173_n 6.3694e-19 $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_282 N_A_84_21#_M1009_g N_X_c_1173_n 0.00986698f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_283 N_A_84_21#_M1011_g N_X_c_1173_n 0.00986698f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_284 N_A_84_21#_M1014_g N_X_c_1173_n 6.3694e-19 $X=2.215 $Y=0.655 $X2=0 $Y2=0
cc_285 N_A_84_21#_M1012_g N_X_c_1177_n 7.09394e-19 $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A_84_21#_M1015_g N_X_c_1177_n 0.0144592f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A_84_21#_M1021_g N_X_c_1177_n 0.0144592f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_288 N_A_84_21#_M1022_g N_X_c_1177_n 7.09394e-19 $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_289 N_A_84_21#_M1011_g N_X_c_1149_n 0.01115f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_290 N_A_84_21#_M1014_g N_X_c_1149_n 0.01115f $X=2.215 $Y=0.655 $X2=0 $Y2=0
cc_291 N_A_84_21#_c_306_p N_X_c_1149_n 0.0388321f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_292 N_A_84_21#_c_177_n N_X_c_1149_n 0.00224206f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_293 N_A_84_21#_M1021_g N_X_c_1154_n 0.0113972f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A_84_21#_M1022_g N_X_c_1154_n 0.0113972f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_295 N_A_84_21#_c_306_p N_X_c_1154_n 0.031822f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_296 N_A_84_21#_c_177_n N_X_c_1154_n 0.0021687f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_297 N_A_84_21#_M1011_g N_X_c_1189_n 6.3694e-19 $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_298 N_A_84_21#_M1014_g N_X_c_1189_n 0.00986698f $X=2.215 $Y=0.655 $X2=0 $Y2=0
cc_299 N_A_84_21#_M1025_g N_X_c_1189_n 0.0101725f $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_300 N_A_84_21#_M1027_g N_X_c_1189_n 6.35826e-19 $X=3.145 $Y=0.655 $X2=0 $Y2=0
cc_301 N_A_84_21#_M1021_g N_X_c_1193_n 7.09394e-19 $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A_84_21#_M1022_g N_X_c_1193_n 0.0144592f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A_84_21#_M1024_g N_X_c_1193_n 0.0144592f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A_84_21#_M1031_g N_X_c_1193_n 7.09394e-19 $X=3.075 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A_84_21#_M1025_g N_X_c_1150_n 0.0115433f $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_306 N_A_84_21#_M1027_g N_X_c_1150_n 0.0125187f $X=3.145 $Y=0.655 $X2=0 $Y2=0
cc_307 N_A_84_21#_M1033_g N_X_c_1150_n 0.00238712f $X=3.575 $Y=0.655 $X2=0 $Y2=0
cc_308 N_A_84_21#_c_306_p N_X_c_1150_n 0.0717012f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_309 N_A_84_21#_c_177_n N_X_c_1150_n 0.00669295f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_310 N_A_84_21#_M1024_g N_X_c_1155_n 0.0113506f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_311 N_A_84_21#_M1031_g N_X_c_1155_n 0.0113972f $X=3.075 $Y=2.465 $X2=0 $Y2=0
cc_312 N_A_84_21#_c_306_p N_X_c_1155_n 0.031822f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_313 N_A_84_21#_c_177_n N_X_c_1155_n 0.0021687f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_314 N_A_84_21#_M1031_g N_X_c_1156_n 9.74069e-19 $X=3.075 $Y=2.465 $X2=0 $Y2=0
cc_315 N_A_84_21#_c_306_p N_X_c_1156_n 0.0172704f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_316 N_A_84_21#_c_177_n N_X_c_1156_n 0.00253081f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_317 N_A_84_21#_c_178_n N_X_c_1156_n 0.00122282f $X=3.71 $Y=2.32 $X2=0 $Y2=0
cc_318 N_A_84_21#_M1024_g N_X_c_1210_n 7.12253e-19 $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_319 N_A_84_21#_M1031_g N_X_c_1210_n 0.0140258f $X=3.075 $Y=2.465 $X2=0 $Y2=0
cc_320 N_A_84_21#_M1025_g N_X_c_1212_n 6.29861e-19 $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_321 N_A_84_21#_M1027_g N_X_c_1212_n 0.0100645f $X=3.145 $Y=0.655 $X2=0 $Y2=0
cc_322 N_A_84_21#_M1033_g N_X_c_1212_n 0.00878119f $X=3.575 $Y=0.655 $X2=0 $Y2=0
cc_323 N_A_84_21#_M1004_g N_X_c_1215_n 0.00204705f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_324 N_A_84_21#_M1005_g N_X_c_1215_n 6.1301e-19 $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_325 N_A_84_21#_M1006_g N_X_c_1217_n 0.00209097f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_326 N_A_84_21#_M1012_g N_X_c_1217_n 6.1301e-19 $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_327 N_A_84_21#_M1009_g N_X_c_1151_n 9.7541e-19 $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_328 N_A_84_21#_M1011_g N_X_c_1151_n 9.7541e-19 $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_329 N_A_84_21#_c_306_p N_X_c_1151_n 0.0276081f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_330 N_A_84_21#_c_177_n N_X_c_1151_n 0.00232957f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_331 N_A_84_21#_M1015_g N_X_c_1157_n 0.0010286f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_332 N_A_84_21#_M1021_g N_X_c_1157_n 0.0010286f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_333 N_A_84_21#_c_306_p N_X_c_1157_n 0.0227182f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_334 N_A_84_21#_c_177_n N_X_c_1157_n 0.00226918f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_335 N_A_84_21#_M1014_g N_X_c_1152_n 9.7541e-19 $X=2.215 $Y=0.655 $X2=0 $Y2=0
cc_336 N_A_84_21#_M1025_g N_X_c_1152_n 9.7541e-19 $X=2.645 $Y=0.655 $X2=0 $Y2=0
cc_337 N_A_84_21#_c_306_p N_X_c_1152_n 0.0276081f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_338 N_A_84_21#_c_177_n N_X_c_1152_n 0.00232957f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_339 N_A_84_21#_M1022_g N_X_c_1158_n 0.0010286f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_340 N_A_84_21#_M1024_g N_X_c_1158_n 0.0010286f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_341 N_A_84_21#_c_306_p N_X_c_1158_n 0.0227182f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_342 N_A_84_21#_c_177_n N_X_c_1158_n 0.00226918f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_343 N_A_84_21#_M1004_g X 0.00868252f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_344 N_A_84_21#_M1006_g X 0.0114564f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_345 N_A_84_21#_M1005_g X 0.00509165f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_346 N_A_84_21#_M1012_g X 0.00660702f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_347 N_A_84_21#_M1009_g X 8.21373e-19 $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_348 N_A_84_21#_M1015_g X 0.00106519f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_349 N_A_84_21#_c_306_p X 0.0195238f $X=3.625 $Y=1.43 $X2=0 $Y2=0
cc_350 N_A_84_21#_c_177_n X 0.0343063f $X=3.585 $Y=1.43 $X2=0 $Y2=0
cc_351 N_A_84_21#_c_210_p N_A_843_419#_M1007_s 0.00508546f $X=4.69 $Y=2.57
+ $X2=-0.19 $Y2=-0.245
cc_352 N_A_84_21#_c_204_p N_A_843_419#_M1028_d 0.00482363f $X=5.69 $Y=2.505
+ $X2=0 $Y2=0
cc_353 N_A_84_21#_M1002_s N_A_843_419#_c_1286_n 0.00332774f $X=4.715 $Y=2.095
+ $X2=0 $Y2=0
cc_354 N_A_84_21#_c_210_p N_A_843_419#_c_1286_n 0.00434586f $X=4.69 $Y=2.57
+ $X2=0 $Y2=0
cc_355 N_A_84_21#_c_200_p N_A_843_419#_c_1286_n 0.0151837f $X=5.02 $Y=2.57 $X2=0
+ $Y2=0
cc_356 N_A_84_21#_c_204_p N_A_843_419#_c_1286_n 0.00434586f $X=5.69 $Y=2.505
+ $X2=0 $Y2=0
cc_357 N_A_84_21#_c_199_p N_A_843_419#_c_1290_n 0.0192244f $X=4.225 $Y=2.447
+ $X2=0 $Y2=0
cc_358 N_A_84_21#_c_204_p N_A_843_419#_c_1291_n 0.0190082f $X=5.69 $Y=2.505
+ $X2=0 $Y2=0
cc_359 N_A_84_21#_c_218_p N_A_1243_419#_M1003_s 0.00339898f $X=6.69 $Y=2.585
+ $X2=-0.19 $Y2=-0.245
cc_360 N_A_84_21#_M1017_d N_A_1243_419#_c_1308_n 0.004731f $X=6.645 $Y=2.095
+ $X2=0 $Y2=0
cc_361 N_A_84_21#_c_226_p N_A_1243_419#_c_1308_n 0.0184311f $X=6.855 $Y=2.585
+ $X2=0 $Y2=0
cc_362 N_A_84_21#_c_218_p N_A_1243_419#_c_1308_n 0.0047595f $X=6.69 $Y=2.585
+ $X2=0 $Y2=0
cc_363 N_A_84_21#_c_218_p N_A_1243_419#_c_1311_n 0.0154232f $X=6.69 $Y=2.585
+ $X2=0 $Y2=0
cc_364 N_A_84_21#_c_202_p N_VGND_M1018_d 0.00757759f $X=6.62 $Y=0.745 $X2=0
+ $Y2=0
cc_365 N_A_84_21#_M1004_g N_VGND_c_1335_n 0.00936134f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_366 N_A_84_21#_M1005_g N_VGND_c_1336_n 0.00325932f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_367 N_A_84_21#_M1009_g N_VGND_c_1336_n 0.00325932f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_368 N_A_84_21#_M1011_g N_VGND_c_1337_n 0.00325932f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_369 N_A_84_21#_M1014_g N_VGND_c_1337_n 0.00325932f $X=2.215 $Y=0.655 $X2=0
+ $Y2=0
cc_370 N_A_84_21#_M1025_g N_VGND_c_1338_n 0.00358565f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_371 N_A_84_21#_M1027_g N_VGND_c_1338_n 0.00569016f $X=3.145 $Y=0.655 $X2=0
+ $Y2=0
cc_372 N_A_84_21#_M1033_g N_VGND_c_1339_n 0.00406888f $X=3.575 $Y=0.655 $X2=0
+ $Y2=0
cc_373 N_A_84_21#_c_177_n N_VGND_c_1339_n 3.48248e-19 $X=3.585 $Y=1.43 $X2=0
+ $Y2=0
cc_374 N_A_84_21#_c_179_n N_VGND_c_1339_n 0.0133914f $X=4.135 $Y=1.35 $X2=0
+ $Y2=0
cc_375 N_A_84_21#_c_180_n N_VGND_c_1339_n 0.0169041f $X=4.22 $Y=1.265 $X2=0
+ $Y2=0
cc_376 N_A_84_21#_c_195_p N_VGND_c_1339_n 0.0131327f $X=4.305 $Y=0.77 $X2=0
+ $Y2=0
cc_377 N_A_84_21#_c_181_n N_VGND_c_1339_n 0.00813919f $X=3.71 $Y=1.43 $X2=0
+ $Y2=0
cc_378 N_A_84_21#_c_202_p N_VGND_c_1340_n 0.0252274f $X=6.62 $Y=0.745 $X2=0
+ $Y2=0
cc_379 N_A_84_21#_M1004_g N_VGND_c_1342_n 0.00550269f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_380 N_A_84_21#_M1005_g N_VGND_c_1342_n 0.00550269f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_381 N_A_84_21#_M1009_g N_VGND_c_1344_n 0.00550269f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_382 N_A_84_21#_M1011_g N_VGND_c_1344_n 0.00550269f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_383 N_A_84_21#_M1014_g N_VGND_c_1346_n 0.00550269f $X=2.215 $Y=0.655 $X2=0
+ $Y2=0
cc_384 N_A_84_21#_M1025_g N_VGND_c_1346_n 0.00550269f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_385 N_A_84_21#_M1027_g N_VGND_c_1348_n 0.00550269f $X=3.145 $Y=0.655 $X2=0
+ $Y2=0
cc_386 N_A_84_21#_M1033_g N_VGND_c_1348_n 0.00550269f $X=3.575 $Y=0.655 $X2=0
+ $Y2=0
cc_387 N_A_84_21#_c_202_p N_VGND_c_1350_n 0.00228632f $X=6.62 $Y=0.745 $X2=0
+ $Y2=0
cc_388 N_A_84_21#_c_195_p N_VGND_c_1352_n 5.77199e-19 $X=4.305 $Y=0.77 $X2=0
+ $Y2=0
cc_389 N_A_84_21#_c_202_p N_VGND_c_1352_n 0.00230949f $X=6.62 $Y=0.745 $X2=0
+ $Y2=0
cc_390 N_A_84_21#_M1016_s N_VGND_c_1354_n 0.00281482f $X=4.625 $Y=0.235 $X2=0
+ $Y2=0
cc_391 N_A_84_21#_M1008_s N_VGND_c_1354_n 0.00227342f $X=6.645 $Y=0.235 $X2=0
+ $Y2=0
cc_392 N_A_84_21#_M1004_g N_VGND_c_1354_n 0.0107186f $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_393 N_A_84_21#_M1005_g N_VGND_c_1354_n 0.00990228f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_394 N_A_84_21#_M1009_g N_VGND_c_1354_n 0.00990228f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_395 N_A_84_21#_M1011_g N_VGND_c_1354_n 0.00990228f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_396 N_A_84_21#_M1014_g N_VGND_c_1354_n 0.00990228f $X=2.215 $Y=0.655 $X2=0
+ $Y2=0
cc_397 N_A_84_21#_M1025_g N_VGND_c_1354_n 0.0100866f $X=2.645 $Y=0.655 $X2=0
+ $Y2=0
cc_398 N_A_84_21#_M1027_g N_VGND_c_1354_n 0.0100592f $X=3.145 $Y=0.655 $X2=0
+ $Y2=0
cc_399 N_A_84_21#_M1033_g N_VGND_c_1354_n 0.0100723f $X=3.575 $Y=0.655 $X2=0
+ $Y2=0
cc_400 N_A_84_21#_c_195_p N_VGND_c_1354_n 0.00117236f $X=4.305 $Y=0.77 $X2=0
+ $Y2=0
cc_401 N_A_84_21#_c_222_p N_VGND_c_1354_n 7.47138e-19 $X=4.67 $Y=0.725 $X2=0
+ $Y2=0
cc_402 N_A_84_21#_c_202_p N_VGND_c_1354_n 0.0119153f $X=6.62 $Y=0.745 $X2=0
+ $Y2=0
cc_403 N_A_84_21#_c_180_n N_A_839_47#_M1010_s 2.20368e-19 $X=4.22 $Y=1.265
+ $X2=-0.19 $Y2=-0.245
cc_404 N_A_84_21#_c_195_p N_A_839_47#_M1010_s 5.68593e-19 $X=4.305 $Y=0.77
+ $X2=-0.19 $Y2=-0.245
cc_405 N_A_84_21#_c_222_p N_A_839_47#_M1010_s 0.00542771f $X=4.67 $Y=0.725
+ $X2=-0.19 $Y2=-0.245
cc_406 N_A_84_21#_c_202_p N_A_839_47#_M1019_d 0.00494709f $X=6.62 $Y=0.745 $X2=0
+ $Y2=0
cc_407 N_A_84_21#_M1016_s N_A_839_47#_c_1465_n 0.0045759f $X=4.625 $Y=0.235
+ $X2=0 $Y2=0
cc_408 N_A_84_21#_c_222_p N_A_839_47#_c_1465_n 0.00542407f $X=4.67 $Y=0.725
+ $X2=0 $Y2=0
cc_409 N_A_84_21#_c_201_p N_A_839_47#_c_1465_n 0.01824f $X=5 $Y=0.725 $X2=0
+ $Y2=0
cc_410 N_A_84_21#_c_202_p N_A_839_47#_c_1465_n 0.00540481f $X=6.62 $Y=0.745
+ $X2=0 $Y2=0
cc_411 N_A_84_21#_c_195_p N_A_839_47#_c_1469_n 0.00602713f $X=4.305 $Y=0.77
+ $X2=0 $Y2=0
cc_412 N_A_84_21#_c_222_p N_A_839_47#_c_1469_n 0.0097141f $X=4.67 $Y=0.725 $X2=0
+ $Y2=0
cc_413 N_A_84_21#_c_202_p N_A_839_47#_c_1471_n 0.0186336f $X=6.62 $Y=0.745 $X2=0
+ $Y2=0
cc_414 N_A_84_21#_c_202_p N_A_1243_47#_M1001_s 0.00367877f $X=6.62 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_415 N_A_84_21#_M1008_s N_A_1243_47#_c_1488_n 0.00335484f $X=6.645 $Y=0.235
+ $X2=0 $Y2=0
cc_416 N_A_84_21#_c_237_p N_A_1243_47#_c_1488_n 0.0148564f $X=6.785 $Y=0.725
+ $X2=0 $Y2=0
cc_417 N_A_84_21#_c_202_p N_A_1243_47#_c_1488_n 0.0167779f $X=6.62 $Y=0.745
+ $X2=0 $Y2=0
cc_418 N_S_M1010_g N_A1_M1016_g 0.0382865f $X=4.12 $Y=0.555 $X2=0 $Y2=0
cc_419 N_S_M1018_g N_A1_M1019_g 0.0317965f $X=5.55 $Y=0.555 $X2=0 $Y2=0
cc_420 N_S_c_467_n N_A1_M1017_g 0.00284044f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_421 N_S_c_467_n N_A1_M1026_g 0.0047241f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_422 N_S_c_467_n N_A1_c_634_n 0.00433599f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_423 N_S_M1010_g N_A1_c_635_n 3.52838e-19 $X=4.12 $Y=0.555 $X2=0 $Y2=0
cc_424 N_S_c_463_n N_A1_c_636_n 0.0140528f $X=5.355 $Y=2.15 $X2=0 $Y2=0
cc_425 N_S_c_467_n N_A1_c_636_n 0.0493139f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_426 N_S_c_499_n N_A1_c_636_n 0.0229319f $X=5.665 $Y=2.035 $X2=0 $Y2=0
cc_427 N_S_c_456_n N_A1_c_636_n 0.0013891f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_428 N_S_c_457_n N_A1_c_636_n 0.0185381f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_429 N_S_M1010_g N_A1_c_637_n 0.0010488f $X=4.12 $Y=0.555 $X2=0 $Y2=0
cc_430 N_S_c_452_n N_A1_c_637_n 0.00598683f $X=4.19 $Y=1.77 $X2=0 $Y2=0
cc_431 N_S_c_453_n N_A1_c_637_n 0.00380825f $X=4.19 $Y=1.77 $X2=0 $Y2=0
cc_432 N_S_c_463_n N_A1_c_637_n 0.00264964f $X=5.355 $Y=2.15 $X2=0 $Y2=0
cc_433 N_S_c_464_n N_A1_c_637_n 0.00362881f $X=4.565 $Y=2.15 $X2=0 $Y2=0
cc_434 N_S_M1010_g N_A1_c_638_n 0.00498166f $X=4.12 $Y=0.555 $X2=0 $Y2=0
cc_435 N_S_c_452_n N_A1_c_638_n 0.0113888f $X=4.19 $Y=1.77 $X2=0 $Y2=0
cc_436 N_S_c_453_n N_A1_c_638_n 0.00141072f $X=4.19 $Y=1.77 $X2=0 $Y2=0
cc_437 N_S_c_463_n N_A1_c_638_n 0.00265275f $X=5.355 $Y=2.15 $X2=0 $Y2=0
cc_438 N_S_c_464_n N_A1_c_638_n 0.00529896f $X=4.565 $Y=2.15 $X2=0 $Y2=0
cc_439 N_S_c_467_n A1 0.0241667f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_440 N_S_M1018_g N_A1_c_640_n 0.00186526f $X=5.55 $Y=0.555 $X2=0 $Y2=0
cc_441 N_S_c_464_n N_A1_c_640_n 2.71463e-19 $X=4.565 $Y=2.15 $X2=0 $Y2=0
cc_442 N_S_c_467_n N_A1_c_641_n 0.0154228f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_443 N_S_M1007_g N_A0_M1002_g 0.0372117f $X=4.14 $Y=2.595 $X2=0 $Y2=0
cc_444 N_S_c_452_n N_A0_M1002_g 9.66873e-19 $X=4.19 $Y=1.77 $X2=0 $Y2=0
cc_445 N_S_c_463_n N_A0_M1002_g 0.00891024f $X=5.355 $Y=2.15 $X2=0 $Y2=0
cc_446 N_S_c_464_n N_A0_M1002_g 0.0046699f $X=4.565 $Y=2.15 $X2=0 $Y2=0
cc_447 N_S_c_463_n N_A0_M1028_g 0.0107472f $X=5.355 $Y=2.15 $X2=0 $Y2=0
cc_448 N_S_c_464_n N_A0_M1028_g 3.93205e-19 $X=4.565 $Y=2.15 $X2=0 $Y2=0
cc_449 N_S_M1018_g N_A0_c_753_n 0.0126113f $X=5.55 $Y=0.555 $X2=0 $Y2=0
cc_450 N_S_c_456_n N_A0_c_753_n 0.00106519f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_451 N_S_c_457_n N_A0_c_753_n 0.0120624f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_452 N_S_c_452_n N_A0_c_755_n 0.00352522f $X=4.19 $Y=1.77 $X2=0 $Y2=0
cc_453 N_S_c_453_n N_A0_c_755_n 3.67533e-19 $X=4.19 $Y=1.77 $X2=0 $Y2=0
cc_454 N_S_c_463_n N_A0_c_755_n 0.0234906f $X=5.355 $Y=2.15 $X2=0 $Y2=0
cc_455 N_S_c_456_n N_A0_c_755_n 0.00109896f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_456 N_S_M1010_g N_A0_c_756_n 4.9189e-19 $X=4.12 $Y=0.555 $X2=0 $Y2=0
cc_457 N_S_M1023_g N_A0_c_756_n 0.0397827f $X=5.57 $Y=2.595 $X2=0 $Y2=0
cc_458 N_S_c_452_n N_A0_c_756_n 7.38545e-19 $X=4.19 $Y=1.77 $X2=0 $Y2=0
cc_459 N_S_c_453_n N_A0_c_756_n 0.0157413f $X=4.19 $Y=1.77 $X2=0 $Y2=0
cc_460 N_S_c_463_n N_A0_c_756_n 0.00100734f $X=5.355 $Y=2.15 $X2=0 $Y2=0
cc_461 N_S_c_456_n N_A0_c_756_n 0.0212772f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_462 N_S_c_457_n N_A0_c_756_n 0.00513985f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_463 N_S_M1018_g N_A0_c_757_n 0.00891902f $X=5.55 $Y=0.555 $X2=0 $Y2=0
cc_464 N_S_c_456_n N_A0_c_757_n 2.15899e-19 $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_465 N_S_c_457_n N_A0_c_757_n 0.0199172f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_466 N_S_M1018_g N_A_1179_311#_M1001_g 0.0406403f $X=5.55 $Y=0.555 $X2=0 $Y2=0
cc_467 N_S_M1023_g N_A_1179_311#_M1003_g 0.0357121f $X=5.57 $Y=2.595 $X2=0 $Y2=0
cc_468 N_S_c_467_n N_A_1179_311#_M1003_g 0.00114504f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_469 N_S_c_457_n N_A_1179_311#_M1003_g 4.2286e-19 $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_470 N_S_M1030_g N_A_1179_311#_M1020_g 0.021964f $X=8.115 $Y=0.655 $X2=0 $Y2=0
cc_471 N_S_M1000_g N_A_1179_311#_M1013_g 0.0368799f $X=8.125 $Y=2.465 $X2=0
+ $Y2=0
cc_472 N_S_c_454_n N_A_1179_311#_M1013_g 0.00140132f $X=8.205 $Y=1.51 $X2=0
+ $Y2=0
cc_473 N_S_c_455_n N_A_1179_311#_M1013_g 0.00421405f $X=8.205 $Y=1.51 $X2=0
+ $Y2=0
cc_474 N_S_c_467_n N_A_1179_311#_M1013_g 0.00391839f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_475 N_S_c_558_p N_A_1179_311#_M1013_g 0.00149323f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_476 N_S_c_559_p N_A_1179_311#_M1013_g 0.00161355f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_477 N_S_c_470_n N_A_1179_311#_M1013_g 0.00192517f $X=7.92 $Y=1.92 $X2=0 $Y2=0
cc_478 N_S_M1023_g N_A_1179_311#_c_856_n 6.59012e-19 $X=5.57 $Y=2.595 $X2=0
+ $Y2=0
cc_479 N_S_c_463_n N_A_1179_311#_c_856_n 0.00173563f $X=5.355 $Y=2.15 $X2=0
+ $Y2=0
cc_480 N_S_c_467_n N_A_1179_311#_c_856_n 0.0140934f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_481 N_S_c_499_n N_A_1179_311#_c_856_n 3.30389e-19 $X=5.665 $Y=2.035 $X2=0
+ $Y2=0
cc_482 N_S_c_456_n N_A_1179_311#_c_856_n 0.00113205f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_483 N_S_c_457_n N_A_1179_311#_c_856_n 0.0302729f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_484 N_S_c_456_n N_A_1179_311#_c_857_n 0.0215068f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_485 N_S_c_457_n N_A_1179_311#_c_857_n 0.00113378f $X=5.52 $Y=1.72 $X2=0 $Y2=0
cc_486 N_S_c_467_n N_A_1179_311#_c_877_n 0.037832f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_487 N_S_M1023_g N_A_1179_311#_c_879_n 5.75556e-19 $X=5.57 $Y=2.595 $X2=0
+ $Y2=0
cc_488 N_S_c_463_n N_A_1179_311#_c_879_n 0.00504276f $X=5.355 $Y=2.15 $X2=0
+ $Y2=0
cc_489 N_S_c_467_n N_A_1179_311#_c_879_n 0.00433533f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_490 N_S_c_499_n N_A_1179_311#_c_879_n 3.58436e-19 $X=5.665 $Y=2.035 $X2=0
+ $Y2=0
cc_491 N_S_M1000_g N_A_1179_311#_c_858_n 0.00103129f $X=8.125 $Y=2.465 $X2=0
+ $Y2=0
cc_492 N_S_c_454_n N_A_1179_311#_c_858_n 0.00761961f $X=8.205 $Y=1.51 $X2=0
+ $Y2=0
cc_493 N_S_c_467_n N_A_1179_311#_c_858_n 0.0140414f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_494 N_S_c_558_p N_A_1179_311#_c_858_n 0.00122429f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_495 N_S_c_559_p N_A_1179_311#_c_858_n 0.00904353f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_496 N_S_c_470_n N_A_1179_311#_c_858_n 0.0105528f $X=7.92 $Y=1.92 $X2=0 $Y2=0
cc_497 N_S_M1000_g N_A_1179_311#_c_912_n 0.0124105f $X=8.125 $Y=2.465 $X2=0
+ $Y2=0
cc_498 N_S_c_454_n N_A_1179_311#_c_912_n 0.00407839f $X=8.205 $Y=1.51 $X2=0
+ $Y2=0
cc_499 N_S_c_467_n N_A_1179_311#_c_912_n 0.00951454f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_500 N_S_c_558_p N_A_1179_311#_c_912_n 0.00414239f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_501 N_S_c_559_p N_A_1179_311#_c_912_n 0.0128708f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_502 N_S_M1030_g N_A_1179_311#_c_859_n 0.014729f $X=8.115 $Y=0.655 $X2=0 $Y2=0
cc_503 N_S_c_454_n N_A_1179_311#_c_859_n 0.0399432f $X=8.205 $Y=1.51 $X2=0 $Y2=0
cc_504 N_S_c_455_n N_A_1179_311#_c_859_n 0.00423266f $X=8.205 $Y=1.51 $X2=0
+ $Y2=0
cc_505 N_S_M1030_g N_A_1179_311#_c_861_n 0.0121985f $X=8.115 $Y=0.655 $X2=0
+ $Y2=0
cc_506 N_S_c_454_n N_A_1179_311#_c_869_n 0.00936931f $X=8.205 $Y=1.51 $X2=0
+ $Y2=0
cc_507 N_S_c_455_n N_A_1179_311#_c_869_n 0.00265266f $X=8.205 $Y=1.51 $X2=0
+ $Y2=0
cc_508 N_S_c_558_p N_A_1179_311#_c_869_n 0.00639305f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_509 N_S_M1030_g N_A_1179_311#_c_924_n 0.00114744f $X=8.115 $Y=0.655 $X2=0
+ $Y2=0
cc_510 N_S_c_454_n N_A_1179_311#_c_924_n 0.0138698f $X=8.205 $Y=1.51 $X2=0 $Y2=0
cc_511 N_S_M1030_g N_A_1179_311#_c_862_n 0.0116298f $X=8.115 $Y=0.655 $X2=0
+ $Y2=0
cc_512 N_S_c_454_n N_A_1179_311#_c_862_n 0.00128883f $X=8.205 $Y=1.51 $X2=0
+ $Y2=0
cc_513 N_S_c_467_n N_A_1179_311#_c_863_n 0.00515758f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_514 N_S_c_467_n N_A_1179_311#_c_880_n 0.00389533f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_515 N_S_c_558_p N_A_1179_311#_c_880_n 0.00122429f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_516 N_S_c_464_n N_VPWR_M1032_s 9.83534e-19 $X=4.565 $Y=2.15 $X2=0 $Y2=0
cc_517 N_S_c_467_n N_VPWR_M1023_d 0.00193959f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_518 N_S_c_467_n N_VPWR_M1013_d 0.00133034f $X=7.775 $Y=2.035 $X2=0 $Y2=0
cc_519 N_S_c_558_p N_VPWR_M1013_d 0.00642328f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_520 N_S_c_559_p N_VPWR_M1013_d 0.00585447f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_521 N_S_c_470_n N_VPWR_M1013_d 0.001394f $X=7.92 $Y=1.92 $X2=0 $Y2=0
cc_522 N_S_M1007_g N_VPWR_c_1012_n 0.00815564f $X=4.14 $Y=2.595 $X2=0 $Y2=0
cc_523 N_S_M1023_g N_VPWR_c_1013_n 0.00510249f $X=5.57 $Y=2.595 $X2=0 $Y2=0
cc_524 N_S_M1000_g N_VPWR_c_1014_n 0.0110173f $X=8.125 $Y=2.465 $X2=0 $Y2=0
cc_525 N_S_M1007_g N_VPWR_c_1021_n 0.00428402f $X=4.14 $Y=2.595 $X2=0 $Y2=0
cc_526 N_S_M1023_g N_VPWR_c_1021_n 0.00428402f $X=5.57 $Y=2.595 $X2=0 $Y2=0
cc_527 N_S_M1000_g N_VPWR_c_1023_n 0.00486043f $X=8.125 $Y=2.465 $X2=0 $Y2=0
cc_528 N_S_M1007_g N_VPWR_c_1005_n 0.00676634f $X=4.14 $Y=2.595 $X2=0 $Y2=0
cc_529 N_S_M1023_g N_VPWR_c_1005_n 0.00649438f $X=5.57 $Y=2.595 $X2=0 $Y2=0
cc_530 N_S_M1000_g N_VPWR_c_1005_n 0.0055095f $X=8.125 $Y=2.465 $X2=0 $Y2=0
cc_531 N_S_c_464_n N_A_843_419#_M1007_s 0.0040556f $X=4.565 $Y=2.15 $X2=-0.19
+ $Y2=-0.245
cc_532 N_S_c_463_n N_A_843_419#_M1028_d 0.00252939f $X=5.355 $Y=2.15 $X2=0 $Y2=0
cc_533 N_S_M1007_g N_A_843_419#_c_1290_n 0.00501944f $X=4.14 $Y=2.595 $X2=0
+ $Y2=0
cc_534 N_S_M1023_g N_A_843_419#_c_1291_n 0.00422409f $X=5.57 $Y=2.595 $X2=0
+ $Y2=0
cc_535 N_S_c_467_n N_A_1243_419#_c_1312_n 0.00162491f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_536 N_S_M1010_g N_VGND_c_1339_n 0.0132565f $X=4.12 $Y=0.555 $X2=0 $Y2=0
cc_537 N_S_M1018_g N_VGND_c_1340_n 0.00485459f $X=5.55 $Y=0.555 $X2=0 $Y2=0
cc_538 N_S_M1030_g N_VGND_c_1341_n 0.00717665f $X=8.115 $Y=0.655 $X2=0 $Y2=0
cc_539 N_S_M1010_g N_VGND_c_1352_n 0.00512179f $X=4.12 $Y=0.555 $X2=0 $Y2=0
cc_540 N_S_M1018_g N_VGND_c_1352_n 0.00420369f $X=5.55 $Y=0.555 $X2=0 $Y2=0
cc_541 N_S_M1030_g N_VGND_c_1353_n 0.0054895f $X=8.115 $Y=0.655 $X2=0 $Y2=0
cc_542 N_S_M1010_g N_VGND_c_1354_n 0.00915933f $X=4.12 $Y=0.555 $X2=0 $Y2=0
cc_543 N_S_M1018_g N_VGND_c_1354_n 0.00641519f $X=5.55 $Y=0.555 $X2=0 $Y2=0
cc_544 N_S_M1030_g N_VGND_c_1354_n 0.0112878f $X=8.115 $Y=0.655 $X2=0 $Y2=0
cc_545 N_S_M1010_g N_A_839_47#_c_1469_n 0.00346811f $X=4.12 $Y=0.555 $X2=0 $Y2=0
cc_546 N_S_M1018_g N_A_839_47#_c_1471_n 0.00326721f $X=5.55 $Y=0.555 $X2=0 $Y2=0
cc_547 N_A1_c_633_n N_A0_c_753_n 0.00742217f $X=6.93 $Y=1.76 $X2=0 $Y2=0
cc_548 N_A1_c_634_n N_A0_c_753_n 7.23783e-19 $X=6.93 $Y=1.76 $X2=0 $Y2=0
cc_549 N_A1_c_636_n N_A0_c_753_n 0.0243224f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_550 A1 N_A0_c_753_n 0.007435f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_551 N_A1_c_641_n N_A0_c_753_n 0.00766213f $X=6.595 $Y=1.737 $X2=0 $Y2=0
cc_552 N_A1_c_631_n N_A0_c_754_n 0.0109185f $X=4.975 $Y=1.1 $X2=0 $Y2=0
cc_553 N_A1_c_635_n N_A0_c_754_n 0.0136604f $X=4.64 $Y=1.19 $X2=0 $Y2=0
cc_554 N_A1_c_640_n N_A0_c_754_n 2.26938e-19 $X=4.805 $Y=1.19 $X2=0 $Y2=0
cc_555 N_A1_c_631_n N_A0_c_755_n 0.00103272f $X=4.975 $Y=1.1 $X2=0 $Y2=0
cc_556 N_A1_c_636_n N_A0_c_755_n 0.0211558f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_557 N_A1_c_637_n N_A0_c_755_n 0.0021532f $X=4.705 $Y=1.665 $X2=0 $Y2=0
cc_558 N_A1_c_638_n N_A0_c_755_n 0.0142775f $X=4.56 $Y=1.665 $X2=0 $Y2=0
cc_559 N_A1_c_631_n N_A0_c_756_n 0.00920701f $X=4.975 $Y=1.1 $X2=0 $Y2=0
cc_560 N_A1_c_635_n N_A0_c_756_n 0.00101771f $X=4.64 $Y=1.19 $X2=0 $Y2=0
cc_561 N_A1_c_636_n N_A0_c_756_n 0.00349046f $X=6.335 $Y=1.665 $X2=0 $Y2=0
cc_562 N_A1_c_637_n N_A0_c_756_n 0.00276023f $X=4.705 $Y=1.665 $X2=0 $Y2=0
cc_563 N_A1_c_638_n N_A0_c_756_n 0.00408757f $X=4.56 $Y=1.665 $X2=0 $Y2=0
cc_564 N_A1_c_640_n N_A0_c_756_n 0.00736363f $X=4.805 $Y=1.19 $X2=0 $Y2=0
cc_565 N_A1_c_635_n N_A0_c_757_n 0.0119874f $X=4.64 $Y=1.19 $X2=0 $Y2=0
cc_566 N_A1_c_637_n N_A0_c_757_n 4.11066e-19 $X=4.705 $Y=1.665 $X2=0 $Y2=0
cc_567 N_A1_c_638_n N_A0_c_757_n 0.00973739f $X=4.56 $Y=1.665 $X2=0 $Y2=0
cc_568 N_A1_c_640_n N_A0_c_757_n 0.00167437f $X=4.805 $Y=1.19 $X2=0 $Y2=0
cc_569 N_A1_c_633_n N_A0_c_758_n 0.00171942f $X=6.93 $Y=1.76 $X2=0 $Y2=0
cc_570 N_A1_c_634_n N_A0_c_758_n 0.0219699f $X=6.93 $Y=1.76 $X2=0 $Y2=0
cc_571 N_A1_c_641_n N_A0_c_758_n 3.1063e-19 $X=6.595 $Y=1.737 $X2=0 $Y2=0
cc_572 N_A1_c_633_n N_A0_c_759_n 0.0270966f $X=6.93 $Y=1.76 $X2=0 $Y2=0
cc_573 N_A1_c_634_n N_A0_c_759_n 0.00105016f $X=6.93 $Y=1.76 $X2=0 $Y2=0
cc_574 N_A1_c_634_n N_A_1179_311#_M1003_g 0.0450093f $X=6.93 $Y=1.76 $X2=0 $Y2=0
cc_575 N_A1_c_641_n N_A_1179_311#_M1003_g 2.61121e-19 $X=6.595 $Y=1.737 $X2=0
+ $Y2=0
cc_576 N_A1_c_633_n N_A_1179_311#_M1013_g 4.89398e-19 $X=6.93 $Y=1.76 $X2=0
+ $Y2=0
cc_577 N_A1_c_634_n N_A_1179_311#_M1013_g 0.0458655f $X=6.93 $Y=1.76 $X2=0 $Y2=0
cc_578 N_A1_c_634_n N_A_1179_311#_c_856_n 0.00172735f $X=6.93 $Y=1.76 $X2=0
+ $Y2=0
cc_579 N_A1_c_636_n N_A_1179_311#_c_856_n 0.0163422f $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_580 A1 N_A_1179_311#_c_856_n 0.0024718f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_581 N_A1_c_641_n N_A_1179_311#_c_856_n 0.0274506f $X=6.595 $Y=1.737 $X2=0
+ $Y2=0
cc_582 N_A1_c_634_n N_A_1179_311#_c_857_n 0.00837982f $X=6.93 $Y=1.76 $X2=0
+ $Y2=0
cc_583 N_A1_c_636_n N_A_1179_311#_c_857_n 0.00241793f $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_584 A1 N_A_1179_311#_c_857_n 0.0019417f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_585 N_A1_c_641_n N_A_1179_311#_c_857_n 0.00326733f $X=6.595 $Y=1.737 $X2=0
+ $Y2=0
cc_586 N_A1_M1017_g N_A_1179_311#_c_877_n 0.00990584f $X=6.57 $Y=2.595 $X2=0
+ $Y2=0
cc_587 N_A1_M1026_g N_A_1179_311#_c_877_n 0.0123419f $X=7.07 $Y=2.595 $X2=0
+ $Y2=0
cc_588 N_A1_c_634_n N_A_1179_311#_c_877_n 0.00363213f $X=6.93 $Y=1.76 $X2=0
+ $Y2=0
cc_589 N_A1_c_636_n N_A_1179_311#_c_877_n 9.85178e-19 $X=6.335 $Y=1.665 $X2=0
+ $Y2=0
cc_590 A1 N_A_1179_311#_c_877_n 4.07013e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_591 N_A1_c_641_n N_A_1179_311#_c_877_n 0.0444327f $X=6.595 $Y=1.737 $X2=0
+ $Y2=0
cc_592 N_A1_c_633_n N_A_1179_311#_c_858_n 0.0203265f $X=6.93 $Y=1.76 $X2=0 $Y2=0
cc_593 N_A1_c_634_n N_A_1179_311#_c_858_n 0.00272922f $X=6.93 $Y=1.76 $X2=0
+ $Y2=0
cc_594 N_A1_M1026_g N_A_1179_311#_c_880_n 0.00678518f $X=7.07 $Y=2.595 $X2=0
+ $Y2=0
cc_595 N_A1_M1017_g N_VPWR_c_1022_n 0.00358377f $X=6.57 $Y=2.595 $X2=0 $Y2=0
cc_596 N_A1_M1026_g N_VPWR_c_1022_n 0.00357877f $X=7.07 $Y=2.595 $X2=0 $Y2=0
cc_597 N_A1_M1017_g N_VPWR_c_1005_n 0.0056244f $X=6.57 $Y=2.595 $X2=0 $Y2=0
cc_598 N_A1_M1026_g N_VPWR_c_1005_n 0.00582826f $X=7.07 $Y=2.595 $X2=0 $Y2=0
cc_599 N_A1_M1017_g N_A_1243_419#_c_1308_n 0.00821814f $X=6.57 $Y=2.595 $X2=0
+ $Y2=0
cc_600 N_A1_M1026_g N_A_1243_419#_c_1308_n 0.0109638f $X=7.07 $Y=2.595 $X2=0
+ $Y2=0
cc_601 N_A1_M1017_g N_A_1243_419#_c_1311_n 0.00401399f $X=6.57 $Y=2.595 $X2=0
+ $Y2=0
cc_602 N_A1_M1026_g N_A_1243_419#_c_1311_n 4.77867e-19 $X=7.07 $Y=2.595 $X2=0
+ $Y2=0
cc_603 N_A1_M1016_g N_VGND_c_1352_n 0.0035834f $X=4.55 $Y=0.555 $X2=0 $Y2=0
cc_604 N_A1_M1019_g N_VGND_c_1352_n 0.00357877f $X=5.05 $Y=0.555 $X2=0 $Y2=0
cc_605 N_A1_M1016_g N_VGND_c_1354_n 0.00555171f $X=4.55 $Y=0.555 $X2=0 $Y2=0
cc_606 N_A1_M1019_g N_VGND_c_1354_n 0.00580543f $X=5.05 $Y=0.555 $X2=0 $Y2=0
cc_607 N_A1_M1016_g N_A_839_47#_c_1465_n 0.00803937f $X=4.55 $Y=0.555 $X2=0
+ $Y2=0
cc_608 N_A1_M1019_g N_A_839_47#_c_1465_n 0.00955131f $X=5.05 $Y=0.555 $X2=0
+ $Y2=0
cc_609 N_A1_M1016_g N_A_839_47#_c_1469_n 0.00321302f $X=4.55 $Y=0.555 $X2=0
+ $Y2=0
cc_610 N_A1_M1019_g N_A_839_47#_c_1469_n 3.05402e-19 $X=5.05 $Y=0.555 $X2=0
+ $Y2=0
cc_611 N_A0_M1008_g N_A_1179_311#_M1001_g 0.0349635f $X=6.57 $Y=0.555 $X2=0
+ $Y2=0
cc_612 N_A0_c_753_n N_A_1179_311#_M1001_g 0.0122625f $X=6.765 $Y=1.11 $X2=0
+ $Y2=0
cc_613 N_A0_c_758_n N_A_1179_311#_M1001_g 0.00414865f $X=6.93 $Y=1.19 $X2=0
+ $Y2=0
cc_614 N_A0_c_759_n N_A_1179_311#_M1001_g 0.00188847f $X=6.93 $Y=1.11 $X2=0
+ $Y2=0
cc_615 N_A0_M1029_g N_A_1179_311#_M1020_g 0.0249214f $X=7 $Y=0.555 $X2=0 $Y2=0
cc_616 N_A0_c_758_n N_A_1179_311#_M1020_g 0.00583338f $X=6.93 $Y=1.19 $X2=0
+ $Y2=0
cc_617 N_A0_c_753_n N_A_1179_311#_c_856_n 0.0106472f $X=6.765 $Y=1.11 $X2=0
+ $Y2=0
cc_618 N_A0_c_753_n N_A_1179_311#_c_857_n 0.00131941f $X=6.765 $Y=1.11 $X2=0
+ $Y2=0
cc_619 N_A0_M1029_g N_A_1179_311#_c_860_n 4.8735e-19 $X=7 $Y=0.555 $X2=0 $Y2=0
cc_620 N_A0_c_758_n N_A_1179_311#_c_860_n 0.00123483f $X=6.93 $Y=1.19 $X2=0
+ $Y2=0
cc_621 N_A0_c_759_n N_A_1179_311#_c_860_n 0.0089623f $X=6.93 $Y=1.11 $X2=0 $Y2=0
cc_622 N_A0_c_758_n N_A_1179_311#_c_924_n 7.19672e-19 $X=6.93 $Y=1.19 $X2=0
+ $Y2=0
cc_623 N_A0_c_759_n N_A_1179_311#_c_924_n 0.0115636f $X=6.93 $Y=1.11 $X2=0 $Y2=0
cc_624 N_A0_c_758_n N_A_1179_311#_c_862_n 0.00761478f $X=6.93 $Y=1.19 $X2=0
+ $Y2=0
cc_625 N_A0_c_759_n N_A_1179_311#_c_862_n 0.00150854f $X=6.93 $Y=1.11 $X2=0
+ $Y2=0
cc_626 N_A0_M1002_g N_VPWR_c_1021_n 0.00357877f $X=4.64 $Y=2.595 $X2=0 $Y2=0
cc_627 N_A0_M1028_g N_VPWR_c_1021_n 0.00357877f $X=5.07 $Y=2.595 $X2=0 $Y2=0
cc_628 N_A0_M1002_g N_VPWR_c_1005_n 0.00562115f $X=4.64 $Y=2.595 $X2=0 $Y2=0
cc_629 N_A0_M1028_g N_VPWR_c_1005_n 0.00562115f $X=5.07 $Y=2.595 $X2=0 $Y2=0
cc_630 N_A0_M1002_g N_A_843_419#_c_1286_n 0.00941846f $X=4.64 $Y=2.595 $X2=0
+ $Y2=0
cc_631 N_A0_M1028_g N_A_843_419#_c_1286_n 0.00941846f $X=5.07 $Y=2.595 $X2=0
+ $Y2=0
cc_632 N_A0_M1008_g N_VGND_c_1350_n 0.00366111f $X=6.57 $Y=0.555 $X2=0 $Y2=0
cc_633 N_A0_M1029_g N_VGND_c_1350_n 0.00366111f $X=7 $Y=0.555 $X2=0 $Y2=0
cc_634 N_A0_M1008_g N_VGND_c_1354_n 0.00538943f $X=6.57 $Y=0.555 $X2=0 $Y2=0
cc_635 N_A0_M1029_g N_VGND_c_1354_n 0.00563413f $X=7 $Y=0.555 $X2=0 $Y2=0
cc_636 N_A0_M1008_g N_A_1243_47#_c_1488_n 0.00820048f $X=6.57 $Y=0.555 $X2=0
+ $Y2=0
cc_637 N_A0_M1029_g N_A_1243_47#_c_1488_n 0.0119083f $X=7 $Y=0.555 $X2=0 $Y2=0
cc_638 N_A0_c_759_n N_A_1243_47#_c_1488_n 0.00366057f $X=6.93 $Y=1.11 $X2=0
+ $Y2=0
cc_639 N_A_1179_311#_c_879_n N_VPWR_M1023_d 0.00262003f $X=6.185 $Y=2.18 $X2=0
+ $Y2=0
cc_640 N_A_1179_311#_c_912_n N_VPWR_M1013_d 0.00665095f $X=8.255 $Y=2.405 $X2=0
+ $Y2=0
cc_641 N_A_1179_311#_M1003_g N_VPWR_c_1013_n 0.00510249f $X=6.14 $Y=2.595 $X2=0
+ $Y2=0
cc_642 N_A_1179_311#_M1013_g N_VPWR_c_1014_n 0.00708018f $X=7.58 $Y=2.595 $X2=0
+ $Y2=0
cc_643 N_A_1179_311#_c_912_n N_VPWR_c_1014_n 0.0206668f $X=8.255 $Y=2.405 $X2=0
+ $Y2=0
cc_644 N_A_1179_311#_M1003_g N_VPWR_c_1022_n 0.00425023f $X=6.14 $Y=2.595 $X2=0
+ $Y2=0
cc_645 N_A_1179_311#_M1013_g N_VPWR_c_1022_n 0.00564131f $X=7.58 $Y=2.595 $X2=0
+ $Y2=0
cc_646 N_A_1179_311#_c_870_n N_VPWR_c_1023_n 0.0174288f $X=8.34 $Y=2.46 $X2=0
+ $Y2=0
cc_647 N_A_1179_311#_M1000_d N_VPWR_c_1005_n 0.00266928f $X=8.2 $Y=1.835 $X2=0
+ $Y2=0
cc_648 N_A_1179_311#_M1003_g N_VPWR_c_1005_n 0.00634446f $X=6.14 $Y=2.595 $X2=0
+ $Y2=0
cc_649 N_A_1179_311#_M1013_g N_VPWR_c_1005_n 0.00690916f $X=7.58 $Y=2.595 $X2=0
+ $Y2=0
cc_650 N_A_1179_311#_c_912_n N_VPWR_c_1005_n 0.01275f $X=8.255 $Y=2.405 $X2=0
+ $Y2=0
cc_651 N_A_1179_311#_c_880_n N_VPWR_c_1005_n 7.51695e-19 $X=7.45 $Y=2.18 $X2=0
+ $Y2=0
cc_652 N_A_1179_311#_c_870_n N_VPWR_c_1005_n 0.00963639f $X=8.34 $Y=2.46 $X2=0
+ $Y2=0
cc_653 N_A_1179_311#_c_877_n N_A_1243_419#_M1003_s 0.00357657f $X=7.365 $Y=2.18
+ $X2=-0.19 $Y2=-0.245
cc_654 N_A_1179_311#_c_877_n N_A_1243_419#_M1026_s 0.00575034f $X=7.365 $Y=2.18
+ $X2=0 $Y2=0
cc_655 N_A_1179_311#_c_880_n N_A_1243_419#_M1026_s 0.00397016f $X=7.45 $Y=2.18
+ $X2=0 $Y2=0
cc_656 N_A_1179_311#_c_877_n N_A_1243_419#_c_1308_n 0.00281168f $X=7.365 $Y=2.18
+ $X2=0 $Y2=0
cc_657 N_A_1179_311#_M1003_g N_A_1243_419#_c_1311_n 0.00361296f $X=6.14 $Y=2.595
+ $X2=0 $Y2=0
cc_658 N_A_1179_311#_M1013_g N_A_1243_419#_c_1312_n 0.00514296f $X=7.58 $Y=2.595
+ $X2=0 $Y2=0
cc_659 N_A_1179_311#_c_877_n N_A_1243_419#_c_1312_n 0.00577695f $X=7.365 $Y=2.18
+ $X2=0 $Y2=0
cc_660 N_A_1179_311#_c_880_n N_A_1243_419#_c_1312_n 0.00784404f $X=7.45 $Y=2.18
+ $X2=0 $Y2=0
cc_661 N_A_1179_311#_c_859_n N_VGND_M1020_d 0.00305087f $X=8.165 $Y=1.09 $X2=0
+ $Y2=0
cc_662 N_A_1179_311#_M1001_g N_VGND_c_1340_n 0.00485459f $X=6.14 $Y=0.555 $X2=0
+ $Y2=0
cc_663 N_A_1179_311#_M1020_g N_VGND_c_1341_n 0.00976992f $X=7.5 $Y=0.555 $X2=0
+ $Y2=0
cc_664 N_A_1179_311#_c_859_n N_VGND_c_1341_n 0.0233948f $X=8.165 $Y=1.09 $X2=0
+ $Y2=0
cc_665 N_A_1179_311#_c_860_n N_VGND_c_1341_n 0.00259365f $X=7.695 $Y=1.09 $X2=0
+ $Y2=0
cc_666 N_A_1179_311#_M1001_g N_VGND_c_1350_n 0.00421279f $X=6.14 $Y=0.555 $X2=0
+ $Y2=0
cc_667 N_A_1179_311#_M1020_g N_VGND_c_1350_n 0.00548805f $X=7.5 $Y=0.555 $X2=0
+ $Y2=0
cc_668 N_A_1179_311#_c_861_n N_VGND_c_1353_n 0.0210192f $X=8.33 $Y=0.42 $X2=0
+ $Y2=0
cc_669 N_A_1179_311#_M1030_d N_VGND_c_1354_n 0.00231914f $X=8.19 $Y=0.235 $X2=0
+ $Y2=0
cc_670 N_A_1179_311#_M1001_g N_VGND_c_1354_n 0.0062528f $X=6.14 $Y=0.555 $X2=0
+ $Y2=0
cc_671 N_A_1179_311#_M1020_g N_VGND_c_1354_n 0.0106692f $X=7.5 $Y=0.555 $X2=0
+ $Y2=0
cc_672 N_A_1179_311#_c_861_n N_VGND_c_1354_n 0.0125689f $X=8.33 $Y=0.42 $X2=0
+ $Y2=0
cc_673 N_A_1179_311#_M1001_g N_A_1243_47#_c_1488_n 0.0024106f $X=6.14 $Y=0.555
+ $X2=0 $Y2=0
cc_674 N_A_1179_311#_M1020_g N_A_1243_47#_c_1488_n 0.00269452f $X=7.5 $Y=0.555
+ $X2=0 $Y2=0
cc_675 N_A_1179_311#_M1020_g N_A_1243_47#_c_1496_n 0.00596256f $X=7.5 $Y=0.555
+ $X2=0 $Y2=0
cc_676 N_A_1179_311#_c_860_n N_A_1243_47#_c_1496_n 0.00493823f $X=7.695 $Y=1.09
+ $X2=0 $Y2=0
cc_677 N_VPWR_c_1005_n N_X_M1006_d 0.00223559f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_678 N_VPWR_c_1005_n N_X_M1015_d 0.00223559f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_679 N_VPWR_c_1005_n N_X_M1022_d 0.00223559f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_680 N_VPWR_c_1005_n N_X_M1031_d 0.0041489f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_681 N_VPWR_c_1015_n N_X_c_1162_n 0.0189236f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_682 N_VPWR_c_1005_n N_X_c_1162_n 0.0123859f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_683 N_VPWR_M1012_s N_X_c_1153_n 0.00176461f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_684 N_VPWR_c_1008_n N_X_c_1153_n 0.0135055f $X=1.14 $Y=2.32 $X2=0 $Y2=0
cc_685 N_VPWR_c_1017_n N_X_c_1177_n 0.0189236f $X=1.915 $Y=3.33 $X2=0 $Y2=0
cc_686 N_VPWR_c_1005_n N_X_c_1177_n 0.0123859f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_687 N_VPWR_M1021_s N_X_c_1154_n 0.00176461f $X=1.86 $Y=1.835 $X2=0 $Y2=0
cc_688 N_VPWR_c_1009_n N_X_c_1154_n 0.0135055f $X=2 $Y=2.32 $X2=0 $Y2=0
cc_689 N_VPWR_c_1019_n N_X_c_1193_n 0.0189236f $X=2.775 $Y=3.33 $X2=0 $Y2=0
cc_690 N_VPWR_c_1005_n N_X_c_1193_n 0.0123859f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_691 N_VPWR_M1024_s N_X_c_1155_n 0.00176461f $X=2.72 $Y=1.835 $X2=0 $Y2=0
cc_692 N_VPWR_c_1010_n N_X_c_1155_n 0.0135055f $X=2.86 $Y=2.32 $X2=0 $Y2=0
cc_693 N_VPWR_c_1011_n N_X_c_1210_n 0.0153332f $X=3.555 $Y=3.33 $X2=0 $Y2=0
cc_694 N_VPWR_c_1005_n N_X_c_1210_n 0.00945339f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_695 N_VPWR_c_1007_n N_X_c_1217_n 0.00756924f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_696 N_VPWR_c_1007_n X 0.00144727f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_697 N_VPWR_c_1005_n N_A_843_419#_M1007_s 0.00279854f $X=8.4 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_698 N_VPWR_c_1005_n N_A_843_419#_M1028_d 0.00279854f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_699 N_VPWR_c_1021_n N_A_843_419#_c_1286_n 0.0361696f $X=5.69 $Y=3.33 $X2=0
+ $Y2=0
cc_700 N_VPWR_c_1005_n N_A_843_419#_c_1286_n 0.0238254f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_701 N_VPWR_c_1012_n N_A_843_419#_c_1290_n 0.0163663f $X=3.72 $Y=2.885 $X2=0
+ $Y2=0
cc_702 N_VPWR_c_1021_n N_A_843_419#_c_1290_n 0.0196957f $X=5.69 $Y=3.33 $X2=0
+ $Y2=0
cc_703 N_VPWR_c_1005_n N_A_843_419#_c_1290_n 0.0123432f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_704 N_VPWR_c_1021_n N_A_843_419#_c_1291_n 0.0196957f $X=5.69 $Y=3.33 $X2=0
+ $Y2=0
cc_705 N_VPWR_c_1005_n N_A_843_419#_c_1291_n 0.0123432f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_706 N_VPWR_c_1005_n N_A_1243_419#_M1003_s 0.00225167f $X=8.4 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_707 N_VPWR_c_1005_n N_A_1243_419#_M1026_s 0.00288699f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_708 N_VPWR_c_1022_n N_A_1243_419#_c_1308_n 0.0374817f $X=7.745 $Y=3.33 $X2=0
+ $Y2=0
cc_709 N_VPWR_c_1005_n N_A_1243_419#_c_1308_n 0.0239391f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_710 N_VPWR_c_1022_n N_A_1243_419#_c_1311_n 0.0180867f $X=7.745 $Y=3.33 $X2=0
+ $Y2=0
cc_711 N_VPWR_c_1005_n N_A_1243_419#_c_1311_n 0.0122611f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_712 N_VPWR_c_1014_n N_A_1243_419#_c_1312_n 0.0259741f $X=7.91 $Y=2.885 $X2=0
+ $Y2=0
cc_713 N_VPWR_c_1022_n N_A_1243_419#_c_1312_n 0.0200258f $X=7.745 $Y=3.33 $X2=0
+ $Y2=0
cc_714 N_VPWR_c_1005_n N_A_1243_419#_c_1312_n 0.0125293f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_715 N_VPWR_c_1007_n N_VGND_c_1335_n 0.00876255f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_716 N_X_c_1148_n N_VGND_M1005_d 0.00176461f $X=1.405 $Y=1.01 $X2=0 $Y2=0
cc_717 N_X_c_1149_n N_VGND_M1011_d 0.00176461f $X=2.265 $Y=1.01 $X2=0 $Y2=0
cc_718 N_X_c_1150_n N_VGND_M1025_d 0.00250873f $X=3.195 $Y=1.01 $X2=0 $Y2=0
cc_719 N_X_c_1215_n N_VGND_c_1335_n 0.00792678f $X=0.71 $Y=1.01 $X2=0 $Y2=0
cc_720 X N_VGND_c_1335_n 0.00151553f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_721 N_X_c_1148_n N_VGND_c_1336_n 0.0135055f $X=1.405 $Y=1.01 $X2=0 $Y2=0
cc_722 N_X_c_1149_n N_VGND_c_1337_n 0.0135055f $X=2.265 $Y=1.01 $X2=0 $Y2=0
cc_723 N_X_c_1150_n N_VGND_c_1338_n 0.0192006f $X=3.195 $Y=1.01 $X2=0 $Y2=0
cc_724 N_X_c_1150_n N_VGND_c_1339_n 0.00756924f $X=3.195 $Y=1.01 $X2=0 $Y2=0
cc_725 N_X_c_1159_n N_VGND_c_1342_n 0.015091f $X=0.71 $Y=0.38 $X2=0 $Y2=0
cc_726 N_X_c_1173_n N_VGND_c_1344_n 0.015091f $X=1.57 $Y=0.38 $X2=0 $Y2=0
cc_727 N_X_c_1189_n N_VGND_c_1346_n 0.015091f $X=2.43 $Y=0.38 $X2=0 $Y2=0
cc_728 N_X_c_1212_n N_VGND_c_1348_n 0.015091f $X=3.36 $Y=0.38 $X2=0 $Y2=0
cc_729 N_X_M1004_s N_VGND_c_1354_n 0.00225632f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_730 N_X_M1009_s N_VGND_c_1354_n 0.00225632f $X=1.43 $Y=0.235 $X2=0 $Y2=0
cc_731 N_X_M1014_s N_VGND_c_1354_n 0.00225632f $X=2.29 $Y=0.235 $X2=0 $Y2=0
cc_732 N_X_M1027_s N_VGND_c_1354_n 0.00225632f $X=3.22 $Y=0.235 $X2=0 $Y2=0
cc_733 N_X_c_1159_n N_VGND_c_1354_n 0.0121307f $X=0.71 $Y=0.38 $X2=0 $Y2=0
cc_734 N_X_c_1173_n N_VGND_c_1354_n 0.0121307f $X=1.57 $Y=0.38 $X2=0 $Y2=0
cc_735 N_X_c_1189_n N_VGND_c_1354_n 0.0121307f $X=2.43 $Y=0.38 $X2=0 $Y2=0
cc_736 N_X_c_1212_n N_VGND_c_1354_n 0.0121307f $X=3.36 $Y=0.38 $X2=0 $Y2=0
cc_737 N_VGND_c_1354_n N_A_839_47#_M1010_s 0.00223559f $X=8.4 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_738 N_VGND_c_1354_n N_A_839_47#_M1019_d 0.00279854f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_739 N_VGND_c_1352_n N_A_839_47#_c_1465_n 0.0374817f $X=5.68 $Y=0 $X2=0 $Y2=0
cc_740 N_VGND_c_1354_n N_A_839_47#_c_1465_n 0.0239391f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_741 N_VGND_c_1339_n N_A_839_47#_c_1469_n 0.0164929f $X=3.79 $Y=0.38 $X2=0
+ $Y2=0
cc_742 N_VGND_c_1352_n N_A_839_47#_c_1469_n 0.0179506f $X=5.68 $Y=0 $X2=0 $Y2=0
cc_743 N_VGND_c_1354_n N_A_839_47#_c_1469_n 0.0120948f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_744 N_VGND_c_1352_n N_A_839_47#_c_1471_n 0.0194152f $X=5.68 $Y=0 $X2=0 $Y2=0
cc_745 N_VGND_c_1354_n N_A_839_47#_c_1471_n 0.0122756f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_746 N_VGND_c_1354_n N_A_1243_47#_M1001_s 0.00225719f $X=8.4 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_747 N_VGND_c_1354_n N_A_1243_47#_M1029_d 0.00284083f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_748 N_VGND_c_1341_n N_A_1243_47#_c_1488_n 0.0116786f $X=7.83 $Y=0.525 $X2=0
+ $Y2=0
cc_749 N_VGND_c_1350_n N_A_1243_47#_c_1488_n 0.0567053f $X=7.665 $Y=0 $X2=0
+ $Y2=0
cc_750 N_VGND_c_1354_n N_A_1243_47#_c_1488_n 0.0448316f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_751 N_VGND_c_1341_n N_A_1243_47#_c_1496_n 0.0239461f $X=7.83 $Y=0.525 $X2=0
+ $Y2=0
