* File: sky130_fd_sc_lp__nand4b_1.pxi.spice
* Created: Wed Sep  2 10:06:03 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4B_1%A_N N_A_N_M1003_g N_A_N_M1006_g A_N N_A_N_c_56_n
+ N_A_N_c_57_n PM_SKY130_FD_SC_LP__NAND4B_1%A_N
x_PM_SKY130_FD_SC_LP__NAND4B_1%D N_D_M1004_g N_D_M1001_g D N_D_c_82_n N_D_c_83_n
+ PM_SKY130_FD_SC_LP__NAND4B_1%D
x_PM_SKY130_FD_SC_LP__NAND4B_1%C N_C_M1005_g N_C_M1008_g C C C N_C_c_111_n
+ N_C_c_112_n PM_SKY130_FD_SC_LP__NAND4B_1%C
x_PM_SKY130_FD_SC_LP__NAND4B_1%B N_B_M1007_g N_B_M1002_g B B B N_B_c_146_n
+ N_B_c_147_n PM_SKY130_FD_SC_LP__NAND4B_1%B
x_PM_SKY130_FD_SC_LP__NAND4B_1%A_71_131# N_A_71_131#_M1003_s N_A_71_131#_M1006_s
+ N_A_71_131#_M1000_g N_A_71_131#_M1009_g N_A_71_131#_c_185_n
+ N_A_71_131#_c_191_n N_A_71_131#_c_186_n N_A_71_131#_c_187_n
+ N_A_71_131#_c_188_n N_A_71_131#_c_193_n PM_SKY130_FD_SC_LP__NAND4B_1%A_71_131#
x_PM_SKY130_FD_SC_LP__NAND4B_1%VPWR N_VPWR_M1006_d N_VPWR_M1008_d N_VPWR_M1009_d
+ N_VPWR_c_249_n N_VPWR_c_250_n N_VPWR_c_251_n N_VPWR_c_252_n N_VPWR_c_253_n
+ N_VPWR_c_254_n N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_257_n N_VPWR_c_258_n
+ VPWR N_VPWR_c_248_n PM_SKY130_FD_SC_LP__NAND4B_1%VPWR
x_PM_SKY130_FD_SC_LP__NAND4B_1%Y N_Y_M1000_d N_Y_M1001_d N_Y_M1002_d N_Y_c_294_n
+ N_Y_c_295_n N_Y_c_296_n N_Y_c_297_n N_Y_c_309_n N_Y_c_301_n Y Y Y Y Y
+ N_Y_c_291_n PM_SKY130_FD_SC_LP__NAND4B_1%Y
x_PM_SKY130_FD_SC_LP__NAND4B_1%VGND N_VGND_M1003_d N_VGND_c_336_n N_VGND_c_337_n
+ N_VGND_c_338_n VGND N_VGND_c_339_n N_VGND_c_340_n
+ PM_SKY130_FD_SC_LP__NAND4B_1%VGND
cc_1 VNB N_A_N_M1006_g 0.00873217f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.045
cc_2 VNB A_N 0.00491327f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_N_c_56_n 0.0313049f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_4 VNB N_A_N_c_57_n 0.0227123f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.185
cc_5 VNB N_D_M1001_g 0.00808665f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.045
cc_6 VNB D 0.00713688f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_D_c_82_n 0.029896f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_8 VNB N_D_c_83_n 0.0189959f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.185
cc_9 VNB N_C_M1008_g 0.00826622f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.045
cc_10 VNB C 0.00205827f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_C_c_111_n 0.0331915f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_12 VNB N_C_c_112_n 0.0162637f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_13 VNB N_B_M1002_g 0.00824325f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.045
cc_14 VNB B 0.00610876f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_15 VNB N_B_c_146_n 0.0306371f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_16 VNB N_B_c_147_n 0.0172487f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_17 VNB N_A_71_131#_M1000_g 0.0297002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_71_131#_c_185_n 0.0353068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_71_131#_c_186_n 0.00106609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_71_131#_c_187_n 0.028533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_71_131#_c_188_n 0.0209758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_248_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB Y 0.018969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB Y 0.0296645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_291_n 0.029663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_336_n 0.0187121f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.045
cc_27 VNB N_VGND_c_337_n 0.02527f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_28 VNB N_VGND_c_338_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.35
cc_29 VNB N_VGND_c_339_n 0.0628297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_340_n 0.199282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_A_N_M1006_g 0.0291537f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.045
cc_32 VPB N_D_M1001_g 0.0221403f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.045
cc_33 VPB N_C_M1008_g 0.0204684f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.045
cc_34 VPB N_B_M1002_g 0.0204426f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.045
cc_35 VPB N_A_71_131#_M1009_g 0.0217293f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.185
cc_36 VPB N_A_71_131#_c_185_n 0.00301684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_71_131#_c_191_n 0.0288525f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.35
cc_38 VPB N_A_71_131#_c_187_n 0.00662455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_71_131#_c_193_n 0.0415262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_249_n 0.035401f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.35
cc_41 VPB N_VPWR_c_250_n 0.00439683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_251_n 0.0307535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_252_n 0.0258507f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_253_n 0.00795653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_254_n 0.0170386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_255_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_256_n 0.011849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_257_n 0.0157463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_258_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_248_n 0.0792373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB Y 0.0203426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB Y 0.0177964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 N_A_N_M1006_g N_D_M1001_g 0.0203859f $X=0.695 $Y=2.045 $X2=0 $Y2=0
cc_54 A_N D 0.0261418f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_55 N_A_N_c_56_n D 2.86117e-19 $X=0.605 $Y=1.35 $X2=0 $Y2=0
cc_56 A_N N_D_c_82_n 0.00220021f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_57 N_A_N_c_56_n N_D_c_82_n 0.0204447f $X=0.605 $Y=1.35 $X2=0 $Y2=0
cc_58 N_A_N_c_57_n N_D_c_83_n 0.0117676f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_59 N_A_N_M1006_g N_A_71_131#_c_185_n 0.00582323f $X=0.695 $Y=2.045 $X2=0
+ $Y2=0
cc_60 A_N N_A_71_131#_c_185_n 0.0258517f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_61 N_A_N_c_56_n N_A_71_131#_c_185_n 0.00825642f $X=0.605 $Y=1.35 $X2=0 $Y2=0
cc_62 N_A_N_c_57_n N_A_71_131#_c_185_n 0.00504346f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_63 N_A_N_M1006_g N_A_71_131#_c_191_n 0.0158642f $X=0.695 $Y=2.045 $X2=0 $Y2=0
cc_64 A_N N_A_71_131#_c_188_n 0.00581439f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_N_c_56_n N_A_71_131#_c_188_n 0.00536659f $X=0.605 $Y=1.35 $X2=0 $Y2=0
cc_66 N_A_N_c_57_n N_A_71_131#_c_188_n 0.00293284f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_67 A_N N_A_71_131#_c_193_n 0.0268896f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A_N_c_56_n N_A_71_131#_c_193_n 0.00562391f $X=0.605 $Y=1.35 $X2=0 $Y2=0
cc_69 N_A_N_M1006_g N_VPWR_c_249_n 0.0127642f $X=0.695 $Y=2.045 $X2=0 $Y2=0
cc_70 A_N N_VGND_c_336_n 0.0067576f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A_N_c_57_n N_VGND_c_336_n 0.00409434f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_72 N_A_N_c_57_n N_VGND_c_337_n 0.00396943f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_73 N_A_N_c_57_n N_VGND_c_340_n 0.0046122f $X=0.605 $Y=1.185 $X2=0 $Y2=0
cc_74 N_D_M1001_g N_C_M1008_g 0.0304123f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_75 D C 0.0257082f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_76 N_D_c_82_n C 3.67073e-19 $X=1.145 $Y=1.35 $X2=0 $Y2=0
cc_77 N_D_c_83_n C 0.00331368f $X=1.145 $Y=1.185 $X2=0 $Y2=0
cc_78 D N_C_c_111_n 0.0018783f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_79 N_D_c_82_n N_C_c_111_n 0.0421705f $X=1.145 $Y=1.35 $X2=0 $Y2=0
cc_80 N_D_c_83_n N_C_c_112_n 0.0421705f $X=1.145 $Y=1.185 $X2=0 $Y2=0
cc_81 N_D_M1001_g N_A_71_131#_c_191_n 0.0156025f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_82 D N_A_71_131#_c_191_n 0.0211909f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_83 N_D_c_82_n N_A_71_131#_c_191_n 0.00369946f $X=1.145 $Y=1.35 $X2=0 $Y2=0
cc_84 N_D_M1001_g N_VPWR_c_249_n 0.00583221f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_85 N_D_M1001_g N_VPWR_c_254_n 0.00583607f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_86 N_D_M1001_g N_VPWR_c_248_n 0.011804f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_87 D N_VGND_c_336_n 0.00428201f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_D_c_82_n N_VGND_c_336_n 0.00403473f $X=1.145 $Y=1.35 $X2=0 $Y2=0
cc_89 N_D_c_83_n N_VGND_c_336_n 0.00731125f $X=1.145 $Y=1.185 $X2=0 $Y2=0
cc_90 N_D_c_83_n N_VGND_c_339_n 0.00585385f $X=1.145 $Y=1.185 $X2=0 $Y2=0
cc_91 N_D_c_83_n N_VGND_c_340_n 0.0118303f $X=1.145 $Y=1.185 $X2=0 $Y2=0
cc_92 N_C_M1008_g N_B_M1002_g 0.0418775f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_93 C B 0.0923364f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_94 N_C_c_111_n B 0.00199212f $X=1.685 $Y=1.35 $X2=0 $Y2=0
cc_95 N_C_c_112_n B 0.00223426f $X=1.685 $Y=1.185 $X2=0 $Y2=0
cc_96 C N_B_c_146_n 3.47522e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_97 N_C_c_111_n N_B_c_146_n 0.0205559f $X=1.685 $Y=1.35 $X2=0 $Y2=0
cc_98 C N_B_c_147_n 0.00261784f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_99 N_C_c_112_n N_B_c_147_n 0.0329186f $X=1.685 $Y=1.185 $X2=0 $Y2=0
cc_100 N_C_M1008_g N_A_71_131#_c_191_n 0.0111891f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_101 C N_A_71_131#_c_191_n 0.0218531f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_102 N_C_c_111_n N_A_71_131#_c_191_n 0.00240813f $X=1.685 $Y=1.35 $X2=0 $Y2=0
cc_103 N_C_M1008_g N_VPWR_c_250_n 0.00621433f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_104 N_C_M1008_g N_VPWR_c_254_n 0.0054895f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_105 N_C_M1008_g N_VPWR_c_248_n 0.0102691f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_106 N_C_M1008_g N_Y_c_294_n 7.32094e-19 $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_107 N_C_M1008_g N_Y_c_295_n 0.0108383f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_108 N_C_M1008_g N_Y_c_296_n 0.0118389f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_109 N_C_M1008_g N_Y_c_297_n 9.16075e-19 $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_110 C N_VGND_c_339_n 0.010446f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_111 N_C_c_112_n N_VGND_c_339_n 0.00395586f $X=1.685 $Y=1.185 $X2=0 $Y2=0
cc_112 C N_VGND_c_340_n 0.010014f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_113 N_C_c_112_n N_VGND_c_340_n 0.00602252f $X=1.685 $Y=1.185 $X2=0 $Y2=0
cc_114 C A_334_47# 0.00733994f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_115 B N_A_71_131#_M1000_g 0.00858188f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_116 N_B_c_146_n N_A_71_131#_M1000_g 0.020219f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_117 N_B_c_147_n N_A_71_131#_M1000_g 0.029884f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_118 N_B_M1002_g N_A_71_131#_c_191_n 0.0111891f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_119 B N_A_71_131#_c_191_n 0.0297983f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_120 N_B_c_146_n N_A_71_131#_c_191_n 0.00123623f $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_121 N_B_M1002_g N_A_71_131#_c_186_n 0.00112272f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_122 B N_A_71_131#_c_186_n 0.0106994f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_123 N_B_c_146_n N_A_71_131#_c_186_n 5.92853e-19 $X=2.225 $Y=1.35 $X2=0 $Y2=0
cc_124 N_B_M1002_g N_A_71_131#_c_187_n 0.0269117f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B_M1002_g N_VPWR_c_250_n 0.00606107f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B_M1002_g N_VPWR_c_251_n 4.81961e-19 $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B_M1002_g N_VPWR_c_257_n 0.0054895f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_128 N_B_M1002_g N_VPWR_c_248_n 0.0102964f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_129 N_B_M1002_g N_Y_c_295_n 9.07394e-19 $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_130 N_B_M1002_g N_Y_c_296_n 0.0118389f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_131 N_B_M1002_g N_Y_c_297_n 0.0112541f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_132 N_B_M1002_g N_Y_c_301_n 7.32094e-19 $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_133 B Y 0.00756371f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_134 B N_Y_c_291_n 0.0352231f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_135 N_B_c_147_n N_Y_c_291_n 0.0011516f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_136 B N_VGND_c_339_n 0.0133676f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_137 N_B_c_147_n N_VGND_c_339_n 0.00380566f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_138 B N_VGND_c_340_n 0.013609f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_139 N_B_c_147_n N_VGND_c_340_n 0.00607665f $X=2.225 $Y=1.185 $X2=0 $Y2=0
cc_140 B A_334_47# 0.00651476f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_141 B A_442_47# 0.00963833f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_142 N_A_71_131#_c_191_n N_VPWR_M1006_d 0.00298209f $X=2.6 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_71_131#_c_191_n N_VPWR_M1008_d 0.00347969f $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_144 N_A_71_131#_c_191_n N_VPWR_M1009_d 7.94932e-19 $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_145 N_A_71_131#_c_191_n N_VPWR_c_249_n 0.024241f $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_146 N_A_71_131#_M1009_g N_VPWR_c_251_n 0.014154f $X=2.675 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_71_131#_M1009_g N_VPWR_c_257_n 0.00486043f $X=2.675 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_71_131#_M1009_g N_VPWR_c_248_n 0.0082726f $X=2.675 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_71_131#_c_191_n N_Y_M1001_d 0.00176461f $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_150 N_A_71_131#_c_191_n N_Y_M1002_d 0.00176461f $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_151 N_A_71_131#_c_191_n N_Y_c_294_n 0.0153678f $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_152 N_A_71_131#_c_191_n N_Y_c_296_n 0.0398294f $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_153 N_A_71_131#_M1009_g N_Y_c_309_n 0.0140658f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_71_131#_c_191_n N_Y_c_309_n 0.0145239f $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_155 N_A_71_131#_c_187_n N_Y_c_309_n 0.00283209f $X=2.765 $Y=1.51 $X2=0 $Y2=0
cc_156 N_A_71_131#_c_191_n N_Y_c_301_n 0.0153678f $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_157 N_A_71_131#_M1000_g Y 0.00474021f $X=2.675 $Y=0.655 $X2=0 $Y2=0
cc_158 N_A_71_131#_c_186_n Y 0.00793827f $X=2.765 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A_71_131#_c_187_n Y 0.00405119f $X=2.765 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A_71_131#_M1000_g Y 0.00533078f $X=2.675 $Y=0.655 $X2=0 $Y2=0
cc_161 N_A_71_131#_M1009_g Y 0.0065605f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_71_131#_c_191_n Y 0.0147119f $X=2.6 $Y=1.78 $X2=0 $Y2=0
cc_163 N_A_71_131#_c_186_n Y 0.0266309f $X=2.765 $Y=1.51 $X2=0 $Y2=0
cc_164 N_A_71_131#_c_187_n Y 0.00821699f $X=2.765 $Y=1.51 $X2=0 $Y2=0
cc_165 N_A_71_131#_M1000_g N_Y_c_291_n 0.0116838f $X=2.675 $Y=0.655 $X2=0 $Y2=0
cc_166 N_A_71_131#_c_188_n N_VGND_c_337_n 0.00864052f $X=0.48 $Y=0.85 $X2=0
+ $Y2=0
cc_167 N_A_71_131#_M1000_g N_VGND_c_339_n 0.0054895f $X=2.675 $Y=0.655 $X2=0
+ $Y2=0
cc_168 N_A_71_131#_M1000_g N_VGND_c_340_n 0.0113886f $X=2.675 $Y=0.655 $X2=0
+ $Y2=0
cc_169 N_A_71_131#_c_188_n N_VGND_c_340_n 0.0152422f $X=0.48 $Y=0.85 $X2=0 $Y2=0
cc_170 N_VPWR_c_248_n N_Y_M1001_d 0.00293134f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_171 N_VPWR_c_248_n N_Y_M1002_d 0.00380103f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_172 N_VPWR_c_254_n N_Y_c_295_n 0.0165751f $X=1.785 $Y=3.33 $X2=0 $Y2=0
cc_173 N_VPWR_c_248_n N_Y_c_295_n 0.0108194f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_174 N_VPWR_M1008_d N_Y_c_296_n 0.00725795f $X=1.74 $Y=1.835 $X2=0 $Y2=0
cc_175 N_VPWR_c_250_n N_Y_c_296_n 0.0257093f $X=1.95 $Y=2.48 $X2=0 $Y2=0
cc_176 N_VPWR_c_257_n N_Y_c_297_n 0.015688f $X=2.725 $Y=3.33 $X2=0 $Y2=0
cc_177 N_VPWR_c_248_n N_Y_c_297_n 0.00984745f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_178 N_VPWR_M1009_d N_Y_c_309_n 0.00770817f $X=2.75 $Y=1.835 $X2=0 $Y2=0
cc_179 N_VPWR_c_251_n N_Y_c_309_n 0.0190932f $X=2.89 $Y=2.485 $X2=0 $Y2=0
cc_180 N_VPWR_c_251_n Y 0.00313887f $X=2.89 $Y=2.485 $X2=0 $Y2=0
cc_181 N_Y_c_291_n N_VGND_c_339_n 0.0368177f $X=2.89 $Y=0.42 $X2=0 $Y2=0
cc_182 N_Y_M1000_d N_VGND_c_340_n 0.00215158f $X=2.75 $Y=0.235 $X2=0 $Y2=0
cc_183 N_Y_c_291_n N_VGND_c_340_n 0.021122f $X=2.89 $Y=0.42 $X2=0 $Y2=0
cc_184 N_VGND_c_340_n A_262_47# 0.00899413f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_185 N_VGND_c_340_n A_334_47# 0.00923159f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_186 N_VGND_c_340_n A_442_47# 0.0105701f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
