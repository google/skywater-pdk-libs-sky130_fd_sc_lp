* File: sky130_fd_sc_lp__o21ba_1.spice
* Created: Fri Aug 28 11:05:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ba_1.pex.spice"
.subckt sky130_fd_sc_lp__o21ba_1  VNB VPB B1_N A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_84_28#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2772 AS=0.2394 PD=2.03333 PS=2.25 NRD=2.136 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1006 N_A_281_138#_M1006_d N_B1_N_M1006_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1554 AS=0.1386 PD=1.58 PS=1.01667 NRD=30 NRS=78.564 M=1 R=2.8
+ SA=75001 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1002 N_A_494_51#_M1002_d N_A_281_138#_M1002_g N_A_84_28#_M1002_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_494_51#_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1596 AS=0.1176 PD=1.22 PS=1.12 NRD=4.284 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1009 N_A_494_51#_M1009_d N_A1_M1009_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1596 PD=2.21 PS=1.22 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A_84_28#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.319725 AS=0.3339 PD=2.6175 PS=3.05 NRD=5.4569 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.4 A=0.189 P=2.82 MULT=1
MM1000 N_A_281_138#_M1000_d N_B1_N_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1386 AS=0.106575 PD=1.5 PS=0.8725 NRD=21.0987 NRS=46.886 M=1 R=2.8
+ SA=75000.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1001 N_A_84_28#_M1001_d N_A_281_138#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.189 AS=0.3339 PD=1.56 PS=3.05 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 A_584_367# N_A2_M1003_g N_A_84_28#_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.189 PD=1.62 PS=1.56 NRD=19.5424 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_584_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2268 PD=3.05 PS=1.62 NRD=0 NRS=19.5424 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o21ba_1.pxi.spice"
*
.ends
*
*
