* File: sky130_fd_sc_lp__xor2_0.pex.spice
* Created: Wed Sep  2 10:40:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XOR2_0%B 3 7 11 15 17 19 20 26 27 28 29 39 43
c77 15 0 1.31594e-19 $X=1.9 $Y=0.635
c78 11 0 1.56626e-19 $X=1.725 $Y=2.725
r79 43 54 2.90608 $w=2.9e-07 $l=2.1e-07 $layer=LI1_cond $X=1.52 $Y=1.71 $X2=1.73
+ $Y2=1.71
r80 40 54 0.685978 $w=4.18e-07 $l=2.5e-08 $layer=LI1_cond $X=1.73 $Y=1.685
+ $X2=1.73 $Y2=1.71
r81 39 42 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.792 $Y=1.685
+ $X2=1.792 $Y2=1.85
r82 39 41 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.792 $Y=1.685
+ $X2=1.792 $Y2=1.52
r83 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.775
+ $Y=1.685 $X2=1.775 $Y2=1.685
r84 29 40 0.548782 $w=4.18e-07 $l=2e-08 $layer=LI1_cond $X=1.73 $Y=1.665
+ $X2=1.73 $Y2=1.685
r85 28 29 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.73 $Y=1.295
+ $X2=1.73 $Y2=1.665
r86 27 43 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=1.2 $Y=1.71 $X2=1.52
+ $Y2=1.71
r87 26 27 19.0749 $w=2.88e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.71 $X2=1.2
+ $Y2=1.71
r88 25 37 47.1166 $w=5.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.465 $Y=1.69
+ $X2=0.465 $Y2=1.855
r89 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.69 $X2=0.37 $Y2=1.69
r90 22 26 10.5309 $w=2.88e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=1.71
+ $X2=0.72 $Y2=1.71
r91 22 24 3.17836 $w=2.9e-07 $l=1.25e-07 $layer=LI1_cond $X=0.455 $Y=1.71
+ $X2=0.33 $Y2=1.71
r92 20 25 34.9827 $w=5.2e-07 $l=3.4e-07 $layer=POLY_cond $X=0.465 $Y=1.35
+ $X2=0.465 $Y2=1.69
r93 20 35 47.1166 $w=5.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.465 $Y=1.35
+ $X2=0.465 $Y2=1.185
r94 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.35 $X2=0.37 $Y2=1.35
r95 17 24 3.6869 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=0.33 $Y=1.565
+ $X2=0.33 $Y2=1.71
r96 17 19 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=0.33 $Y=1.565
+ $X2=0.33 $Y2=1.35
r97 15 41 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=1.9 $Y=0.635
+ $X2=1.9 $Y2=1.52
r98 11 42 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.725 $Y=2.725
+ $X2=1.725 $Y2=1.85
r99 7 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.65 $Y=0.635
+ $X2=0.65 $Y2=1.185
r100 3 37 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=0.475 $Y=2.725
+ $X2=0.475 $Y2=1.855
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_0%A 3 7 11 15 21 27 29 30 34
c52 30 0 1.31594e-19 $X=1.2 $Y=1.295
c53 11 0 1.56626e-19 $X=1.295 $Y=2.725
r54 30 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.295 $X2=1.17 $Y2=1.295
r55 29 30 26.9779 $w=1.83e-07 $l=4.5e-07 $layer=LI1_cond $X=0.72 $Y=1.302
+ $X2=1.17 $Y2=1.302
r56 26 34 2.37141 $w=3.65e-07 $l=1.5e-08 $layer=POLY_cond $X=1.187 $Y=1.28
+ $X2=1.187 $Y2=1.295
r57 26 27 165.623 $w=1.5e-07 $l=3.23e-07 $layer=POLY_cond $X=1.187 $Y=1.205
+ $X2=1.51 $Y2=1.205
r58 23 26 54.866 $w=1.5e-07 $l=1.07e-07 $layer=POLY_cond $X=1.08 $Y=1.205
+ $X2=1.187 $Y2=1.205
r59 20 34 126.475 $w=3.65e-07 $l=8e-07 $layer=POLY_cond $X=1.187 $Y=2.095
+ $X2=1.187 $Y2=1.295
r60 20 21 55.3787 $w=1.5e-07 $l=1.08e-07 $layer=POLY_cond $X=1.187 $Y=2.17
+ $X2=1.295 $Y2=2.17
r61 17 20 165.111 $w=1.5e-07 $l=3.22e-07 $layer=POLY_cond $X=0.865 $Y=2.17
+ $X2=1.187 $Y2=2.17
r62 13 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.51 $Y=1.13
+ $X2=1.51 $Y2=1.205
r63 13 15 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.51 $Y=1.13
+ $X2=1.51 $Y2=0.635
r64 9 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.295 $Y=2.245
+ $X2=1.295 $Y2=2.17
r65 9 11 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.295 $Y=2.245
+ $X2=1.295 $Y2=2.725
r66 5 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.08 $Y=1.13 $X2=1.08
+ $Y2=1.205
r67 5 7 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.08 $Y=1.13 $X2=1.08
+ $Y2=0.635
r68 1 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.865 $Y=2.245
+ $X2=0.865 $Y2=2.17
r69 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.865 $Y=2.245
+ $X2=0.865 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_0%A_27_481# 1 2 7 8 9 11 14 17 20 22 23 26 28
+ 29 33 34 36 37
r83 36 37 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.29 $Y=2.025 $X2=2.29
+ $Y2=1.625
r84 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.38
+ $Y=1.12 $X2=2.38 $Y2=1.12
r85 31 37 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.34 $Y=1.49
+ $X2=2.34 $Y2=1.625
r86 31 33 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.34 $Y=1.49
+ $X2=2.34 $Y2=1.12
r87 30 33 3.41465 $w=2.68e-07 $l=8e-08 $layer=LI1_cond $X=2.34 $Y=1.04 $X2=2.34
+ $Y2=1.12
r88 28 30 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.205 $Y=0.955
+ $X2=2.34 $Y2=1.04
r89 28 29 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=2.205 $Y=0.955
+ $X2=0.96 $Y2=0.955
r90 24 29 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.845 $Y=0.87
+ $X2=0.96 $Y2=0.955
r91 24 26 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.845 $Y=0.87
+ $X2=0.845 $Y2=0.635
r92 22 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.205 $Y=2.11
+ $X2=2.29 $Y2=2.025
r93 22 23 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=2.205 $Y=2.11
+ $X2=0.425 $Y2=2.11
r94 18 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=2.195
+ $X2=0.425 $Y2=2.11
r95 18 20 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.26 $Y=2.195
+ $X2=0.26 $Y2=2.55
r96 16 34 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.38 $Y=1.105
+ $X2=2.38 $Y2=1.12
r97 12 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=1.105
+ $X2=2.875 $Y2=1.03
r98 12 14 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.875 $Y=1.105
+ $X2=2.875 $Y2=2.155
r99 9 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=0.955
+ $X2=2.875 $Y2=1.03
r100 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.875 $Y=0.955
+ $X2=2.875 $Y2=0.635
r101 8 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.545 $Y=1.03
+ $X2=2.38 $Y2=1.105
r102 7 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.8 $Y=1.03
+ $X2=2.875 $Y2=1.03
r103 7 8 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=2.8 $Y=1.03
+ $X2=2.545 $Y2=1.03
r104 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.405 $X2=0.26 $Y2=2.55
r105 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.725
+ $Y=0.425 $X2=0.865 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_0%VPWR 1 2 9 13 16 17 19 20 21 34 35
r39 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r42 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 21 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 19 28 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 19 20 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.922 $Y2=3.33
r49 18 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 18 20 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.922 $Y2=3.33
r51 16 24 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 16 17 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=1.062 $Y2=3.33
r53 15 28 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.21 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 15 17 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.21 $Y=3.33
+ $X2=1.062 $Y2=3.33
r55 11 20 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.922 $Y=3.245
+ $X2=1.922 $Y2=3.33
r56 11 13 19.2074 $w=2.23e-07 $l=3.75e-07 $layer=LI1_cond $X=1.922 $Y=3.245
+ $X2=1.922 $Y2=2.87
r57 7 17 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.062 $Y=3.245
+ $X2=1.062 $Y2=3.33
r58 7 9 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=1.062 $Y=3.245
+ $X2=1.062 $Y2=2.55
r59 2 13 600 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=1 $X=1.8
+ $Y=2.405 $X2=1.94 $Y2=2.87
r60 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.94
+ $Y=2.405 $X2=1.08 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_0%A_274_481# 1 2 9 11 12 13 17 19
c31 9 0 3.13252e-19 $X=1.51 $Y=2.55
r32 19 21 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.29 $Y=2.45 $X2=2.29
+ $Y2=2.75
r33 15 17 29.2379 $w=2.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.12 $Y=2.665
+ $X2=3.12 $Y2=1.98
r34 14 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=2.75
+ $X2=2.29 $Y2=2.75
r35 13 15 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.985 $Y=2.75
+ $X2=3.12 $Y2=2.665
r36 13 14 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.985 $Y=2.75
+ $X2=2.375 $Y2=2.75
r37 11 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=2.45
+ $X2=2.29 $Y2=2.45
r38 11 12 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.205 $Y=2.45
+ $X2=1.64 $Y2=2.45
r39 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.51 $Y=2.535
+ $X2=1.64 $Y2=2.45
r40 7 9 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.51 $Y=2.535
+ $X2=1.51 $Y2=2.55
r41 2 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.95
+ $Y=1.835 $X2=3.09 $Y2=1.98
r42 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.37
+ $Y=2.405 $X2=1.51 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_0%X 1 2 7 9 11 13 14 15 19 25
r33 19 25 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=2.645 $Y=0.555
+ $X2=2.64 $Y2=0.555
r34 15 19 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=0.555
+ $X2=2.645 $Y2=0.555
r35 15 25 1.58958 $w=2.88e-07 $l=4e-08 $layer=LI1_cond $X=2.6 $Y=0.555 $X2=2.64
+ $Y2=0.555
r36 14 15 17.4853 $w=2.88e-07 $l=4.4e-07 $layer=LI1_cond $X=2.16 $Y=0.555
+ $X2=2.6 $Y2=0.555
r37 11 15 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.73 $Y=0.7 $X2=2.73
+ $Y2=0.555
r38 11 13 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=2.73 $Y=0.7
+ $X2=2.73 $Y2=1.815
r39 7 13 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.68 $Y=1.95
+ $X2=2.68 $Y2=1.815
r40 7 9 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=2.68 $Y=1.95 $X2=2.68
+ $Y2=1.98
r41 2 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=1.835 $X2=2.66 $Y2=1.98
r42 1 15 91 $w=1.7e-07 $l=7.52994e-07 $layer=licon1_NDIFF $count=2 $X=1.975
+ $Y=0.425 $X2=2.65 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__XOR2_0%VGND 1 2 3 10 12 14 18 20 22 24 26 38 42
r38 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r40 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r41 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r42 33 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r43 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r45 27 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=0 $X2=1.295
+ $Y2=0
r46 27 29 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.46 $Y=0 $X2=1.68
+ $Y2=0
r47 26 41 4.20444 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=3.172
+ $Y2=0
r48 26 32 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=0 $X2=2.64
+ $Y2=0
r49 24 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 24 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r51 24 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 20 41 3.08026 $w=2.7e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.12 $Y=0.085
+ $X2=3.172 $Y2=0
r53 20 22 23.4757 $w=2.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.12 $Y=0.085
+ $X2=3.12 $Y2=0.635
r54 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.085
+ $X2=1.295 $Y2=0
r55 16 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.295 $Y=0.085
+ $X2=1.295 $Y2=0.595
r56 15 35 4.16519 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.28
+ $Y2=0
r57 14 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=1.295
+ $Y2=0
r58 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=0.56
+ $Y2=0
r59 10 35 3.27265 $w=2.9e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.28 $Y2=0
r60 10 12 21.8567 $w=2.88e-07 $l=5.5e-07 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.415 $Y2=0.635
r61 3 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.95
+ $Y=0.425 $X2=3.09 $Y2=0.635
r62 2 18 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=1.155
+ $Y=0.425 $X2=1.295 $Y2=0.595
r63 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.425 $X2=0.435 $Y2=0.635
.ends

