* File: sky130_fd_sc_lp__nor3b_m.pex.spice
* Created: Fri Aug 28 10:56:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3B_M%C_N 3 5 6 8 10 11 14 16 17 21
c38 21 0 1.79783e-19 $X=0.27 $Y=1.38
c39 14 0 1.10055e-19 $X=0.635 $Y=0.87
r40 16 17 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r41 16 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.38 $X2=0.27 $Y2=1.38
r42 12 14 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.36 $Y=0.87
+ $X2=0.635 $Y2=0.87
r43 11 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.72
+ $X2=0.27 $Y2=1.38
r44 10 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.215
+ $X2=0.27 $Y2=1.38
r45 6 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.635 $Y=0.795
+ $X2=0.635 $Y2=0.87
r46 6 8 96.4 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=0.635 $Y=0.795 $X2=0.635
+ $Y2=0.495
r47 3 11 72.2097 $w=2.67e-07 $l=4.91935e-07 $layer=POLY_cond $X=0.475 $Y=2.12
+ $X2=0.27 $Y2=1.72
r48 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.475 $Y=2.12 $X2=0.475
+ $Y2=2.405
r49 1 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=0.945
+ $X2=0.36 $Y2=0.87
r50 1 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.36 $Y=0.945
+ $X2=0.36 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_M%A 3 7 11 12 13 14 18 19
c44 7 0 6.71248e-20 $X=1.065 $Y=0.495
c45 3 0 1.9212e-20 $X=1.015 $Y=2.405
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.03
+ $Y=1.27 $X2=1.03 $Y2=1.27
r47 13 14 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.14 $Y=1.295
+ $X2=1.14 $Y2=1.665
r48 13 19 0.738746 $w=3.88e-07 $l=2.5e-08 $layer=LI1_cond $X=1.14 $Y=1.295
+ $X2=1.14 $Y2=1.27
r49 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.03 $Y=1.61
+ $X2=1.03 $Y2=1.27
r50 11 12 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.61
+ $X2=1.03 $Y2=1.775
r51 10 18 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.03 $Y=1.105
+ $X2=1.03 $Y2=1.27
r52 7 10 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.065 $Y=0.495
+ $X2=1.065 $Y2=1.105
r53 3 12 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.015 $Y=2.405
+ $X2=1.015 $Y2=1.775
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_M%B 1 3 6 9 12 14 15 19
c43 14 0 1.9212e-20 $X=1.68 $Y=1.295
c44 12 0 1.87727e-20 $X=1.495 $Y=2.045
r45 19 22 51.4356 $w=3.7e-07 $l=1.95e-07 $layer=POLY_cond $X=1.605 $Y=1.345
+ $X2=1.605 $Y2=1.54
r46 19 21 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.605 $Y=1.345
+ $X2=1.605 $Y2=1.18
r47 14 15 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=1.295
+ $X2=1.66 $Y2=1.665
r48 14 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.625
+ $Y=1.345 $X2=1.625 $Y2=1.345
r49 10 12 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=1.375 $Y=2.045
+ $X2=1.495 $Y2=2.045
r50 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.495 $Y=1.97
+ $X2=1.495 $Y2=2.045
r51 9 22 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.495 $Y=1.97
+ $X2=1.495 $Y2=1.54
r52 6 21 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=1.495 $Y=0.495
+ $X2=1.495 $Y2=1.18
r53 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.375 $Y=2.12
+ $X2=1.375 $Y2=2.045
r54 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.375 $Y=2.12 $X2=1.375
+ $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_M%A_27_439# 1 2 10 11 13 15 18 22 26 28 31 32
+ 35 36 43 45 49 50
c82 45 0 1.55344e-19 $X=0.69 $Y=2.14
c83 43 0 1.79783e-19 $X=0.69 $Y=0.905
c84 26 0 6.71248e-20 $X=0.42 $Y=0.495
r85 50 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=2.945
+ $X2=1.825 $Y2=2.78
r86 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=2.945 $X2=1.825 $Y2=2.945
r87 36 39 7.3171 $w=3.13e-07 $l=2e-07 $layer=LI1_cond $X=0.267 $Y=2.14 $X2=0.267
+ $Y2=2.34
r88 35 49 3.3206 $w=2.93e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=2.927
+ $X2=1.825 $Y2=2.927
r89 34 35 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.74 $Y=2.225
+ $X2=1.74 $Y2=2.78
r90 33 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=2.14
+ $X2=0.69 $Y2=2.14
r91 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.655 $Y=2.14
+ $X2=1.74 $Y2=2.225
r92 32 33 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.655 $Y=2.14
+ $X2=0.775 $Y2=2.14
r93 31 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=2.055
+ $X2=0.69 $Y2=2.14
r94 30 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.99
+ $X2=0.69 $Y2=0.905
r95 30 31 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=0.69 $Y=0.99
+ $X2=0.69 $Y2=2.055
r96 29 36 4.34843 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.425 $Y=2.14
+ $X2=0.267 $Y2=2.14
r97 28 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=2.14
+ $X2=0.69 $Y2=2.14
r98 28 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.605 $Y=2.14
+ $X2=0.425 $Y2=2.14
r99 24 43 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=0.905 $X2=0.69
+ $Y2=0.905
r100 24 26 13.872 $w=2.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.39 $Y=0.82
+ $X2=0.39 $Y2=0.495
r101 20 22 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.925 $Y=0.89
+ $X2=2.105 $Y2=0.89
r102 16 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.895 $Y=2.01
+ $X2=2.105 $Y2=2.01
r103 15 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.105 $Y=1.935
+ $X2=2.105 $Y2=2.01
r104 14 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.105 $Y=0.965
+ $X2=2.105 $Y2=0.89
r105 14 15 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=2.105 $Y=0.965
+ $X2=2.105 $Y2=1.935
r106 11 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=0.815
+ $X2=1.925 $Y2=0.89
r107 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.925 $Y=0.815
+ $X2=1.925 $Y2=0.495
r108 10 53 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.895 $Y=2.405
+ $X2=1.895 $Y2=2.78
r109 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.895 $Y=2.085
+ $X2=1.895 $Y2=2.01
r110 7 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.895 $Y=2.085
+ $X2=1.895 $Y2=2.405
r111 2 39 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.195 $X2=0.26 $Y2=2.34
r112 1 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.295
+ $Y=0.285 $X2=0.42 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_M%VPWR 1 6 8 10 20 21 24
r24 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r26 17 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r27 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.76 $Y2=3.33
r28 15 17 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.2 $Y2=3.33
r29 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.76 $Y2=3.33
r32 10 12 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 8 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r34 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.72
+ $Y2=3.33
r35 8 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245 $X2=0.76
+ $Y2=3.33
r37 4 6 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=2.49
r38 1 6 600 $w=1.7e-07 $l=3.85973e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.195 $X2=0.76 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_M%Y 1 2 3 12 14 15 16 17 38
c34 38 0 1.10055e-19 $X=2.16 $Y=0.925
c35 15 0 1.87727e-20 $X=2.16 $Y=1.295
r36 17 32 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=2.155 $Y=2.035
+ $X2=2.155 $Y2=2.34
r37 16 17 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.155 $Y=1.665
+ $X2=2.155 $Y2=2.035
r38 15 16 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.155 $Y=1.295
+ $X2=2.155 $Y2=1.665
r39 14 38 4.34843 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=0.745
r40 14 15 8.81211 $w=4.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.155 $Y=1.01
+ $X2=2.155 $Y2=1.295
r41 10 38 0.193651 $w=3.15e-07 $l=5e-09 $layer=LI1_cond $X=2.155 $Y=0.745
+ $X2=2.16 $Y2=0.745
r42 10 14 1.01224 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=2.155 $Y=0.745
+ $X2=2.155 $Y2=1.01
r43 10 35 33.8889 $w=3.15e-07 $l=8.75e-07 $layer=LI1_cond $X=2.155 $Y=0.745
+ $X2=1.28 $Y2=0.745
r44 10 12 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=2.155 $Y=0.745
+ $X2=2.155 $Y2=0.43
r45 3 32 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.97
+ $Y=2.195 $X2=2.11 $Y2=2.34
r46 2 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.285 $X2=2.14 $Y2=0.43
r47 1 35 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.285 $X2=1.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_M%VGND 1 2 9 11 15 17 18 19 27 28 31
r33 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r34 28 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r35 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r36 25 31 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.73
+ $Y2=0
r37 25 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2.16
+ $Y2=0
r38 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 19 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r40 19 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r41 17 22 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=0 $X2=0.72
+ $Y2=0
r42 17 18 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.745 $Y=0 $X2=0.84
+ $Y2=0
r43 13 31 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=0.085
+ $X2=1.73 $Y2=0
r44 13 15 17.1645 $w=2.08e-07 $l=3.25e-07 $layer=LI1_cond $X=1.73 $Y=0.085
+ $X2=1.73 $Y2=0.41
r45 12 18 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.84
+ $Y2=0
r46 11 31 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.73
+ $Y2=0
r47 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=0.935
+ $Y2=0
r48 7 18 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=0.085
+ $X2=0.84 $Y2=0
r49 7 9 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=0.84 $Y=0.085
+ $X2=0.84 $Y2=0.43
r50 2 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.285 $X2=1.71 $Y2=0.41
r51 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.71
+ $Y=0.285 $X2=0.85 $Y2=0.43
.ends

