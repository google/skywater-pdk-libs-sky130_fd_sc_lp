* File: sky130_fd_sc_lp__o21ai_2.pxi.spice
* Created: Wed Sep  2 10:16:06 2020
* 
x_PM_SKY130_FD_SC_LP__O21AI_2%A1 N_A1_M1005_g N_A1_M1003_g N_A1_M1007_g
+ N_A1_M1010_g N_A1_c_61_n N_A1_c_69_n N_A1_c_62_n A1 A1 N_A1_c_64_n N_A1_c_65_n
+ PM_SKY130_FD_SC_LP__O21AI_2%A1
x_PM_SKY130_FD_SC_LP__O21AI_2%A2 N_A2_c_136_n N_A2_M1001_g N_A2_M1002_g
+ N_A2_c_138_n N_A2_M1009_g N_A2_M1011_g A2 N_A2_c_140_n N_A2_c_141_n
+ PM_SKY130_FD_SC_LP__O21AI_2%A2
x_PM_SKY130_FD_SC_LP__O21AI_2%B1 N_B1_M1004_g N_B1_M1000_g N_B1_c_191_n
+ N_B1_M1008_g N_B1_M1006_g B1 B1 N_B1_c_194_n PM_SKY130_FD_SC_LP__O21AI_2%B1
x_PM_SKY130_FD_SC_LP__O21AI_2%VPWR N_VPWR_M1003_d N_VPWR_M1007_d N_VPWR_M1006_s
+ N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n N_VPWR_c_238_n
+ VPWR N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_233_n
+ PM_SKY130_FD_SC_LP__O21AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O21AI_2%A_113_367# N_A_113_367#_M1003_s
+ N_A_113_367#_M1011_s N_A_113_367#_c_285_n N_A_113_367#_c_280_n
+ N_A_113_367#_c_281_n N_A_113_367#_c_292_p
+ PM_SKY130_FD_SC_LP__O21AI_2%A_113_367#
x_PM_SKY130_FD_SC_LP__O21AI_2%Y N_Y_M1004_d N_Y_M1002_d N_Y_M1000_d N_Y_c_319_n
+ N_Y_c_295_n N_Y_c_300_n Y Y Y N_Y_c_304_n N_Y_c_306_n Y
+ PM_SKY130_FD_SC_LP__O21AI_2%Y
x_PM_SKY130_FD_SC_LP__O21AI_2%A_30_47# N_A_30_47#_M1005_s N_A_30_47#_M1001_s
+ N_A_30_47#_M1010_s N_A_30_47#_M1008_s N_A_30_47#_c_333_n N_A_30_47#_c_334_n
+ N_A_30_47#_c_340_n N_A_30_47#_c_354_n N_A_30_47#_c_335_n N_A_30_47#_c_346_n
+ N_A_30_47#_c_347_n N_A_30_47#_c_364_n N_A_30_47#_c_336_n N_A_30_47#_c_337_n
+ PM_SKY130_FD_SC_LP__O21AI_2%A_30_47#
x_PM_SKY130_FD_SC_LP__O21AI_2%VGND N_VGND_M1005_d N_VGND_M1009_d N_VGND_c_393_n
+ N_VGND_c_394_n VGND N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n
+ N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n PM_SKY130_FD_SC_LP__O21AI_2%VGND
cc_1 VNB N_A1_M1005_g 0.0307707f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_2 VNB N_A1_M1003_g 0.00184777f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_3 VNB N_A1_M1010_g 0.0267318f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=0.655
cc_4 VNB N_A1_c_61_n 0.00111806f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_5 VNB N_A1_c_62_n 0.00169258f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.605
cc_6 VNB A1 0.00541527f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_7 VNB N_A1_c_64_n 0.0543735f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.46
cc_8 VNB N_A1_c_65_n 0.0234112f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.51
cc_9 VNB N_A2_c_136_n 0.0161793f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.295
cc_10 VNB N_A2_M1002_g 0.00726874f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_11 VNB N_A2_c_138_n 0.0169297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_M1011_g 0.00635208f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.345
cc_13 VNB N_A2_c_140_n 0.00554038f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_14 VNB N_A2_c_141_n 0.0414191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_M1004_g 0.0171179f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_16 VNB N_B1_M1000_g 0.00601414f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_17 VNB N_B1_c_191_n 0.0220461f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.675
cc_18 VNB N_B1_M1006_g 0.00857668f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=0.655
cc_19 VNB B1 0.0179106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_194_n 0.0687608f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_21 VNB N_VPWR_c_233_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_295_n 0.00376151f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.78
cc_23 VNB N_A_30_47#_c_333_n 0.00798915f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.345
cc_24 VNB N_A_30_47#_c_334_n 0.0224525f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=0.655
cc_25 VNB N_A_30_47#_c_335_n 0.00680429f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.78
cc_26 VNB N_A_30_47#_c_336_n 0.00220432f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.46
cc_27 VNB N_A_30_47#_c_337_n 0.0312825f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.345
cc_28 VNB N_VGND_c_393_n 4.20494e-19 $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.675
cc_29 VNB N_VGND_c_394_n 0.00499816f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.345
cc_30 VNB N_VGND_c_395_n 0.0158532f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.78
cc_31 VNB N_VGND_c_396_n 0.0168667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_397_n 0.0382261f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_33 VNB N_VGND_c_398_n 0.191119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_399_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.51
cc_35 VNB N_VGND_c_400_n 0.00634044f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.345
cc_36 VPB N_A1_M1003_g 0.0230824f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_37 VPB N_A1_M1007_g 0.0203232f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=2.465
cc_38 VPB N_A1_c_61_n 0.00819765f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_39 VPB N_A1_c_69_n 0.00827138f $X=-0.19 $Y=1.655 $X2=1.245 $Y2=1.605
cc_40 VPB N_A1_c_62_n 4.83595e-19 $X=-0.19 $Y=1.655 $X2=1.415 $Y2=1.605
cc_41 VPB A1 0.00739377f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.58
cc_42 VPB N_A1_c_65_n 0.0063771f $X=-0.19 $Y=1.655 $X2=1.955 $Y2=1.51
cc_43 VPB N_A2_M1002_g 0.0187161f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_44 VPB N_A2_M1011_g 0.020454f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=1.345
cc_45 VPB N_B1_M1000_g 0.0199365f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_46 VPB N_B1_M1006_g 0.0251154f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=0.655
cc_47 VPB B1 0.00875028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_234_n 0.0108182f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=2.465
cc_49 VPB N_VPWR_c_235_n 0.044414f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_236_n 0.00227295f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.78
cc_51 VPB N_VPWR_c_237_n 0.0116683f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_52 VPB N_VPWR_c_238_n 0.0479442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_239_n 0.0359769f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_54 VPB N_VPWR_c_240_n 0.0149952f $X=-0.19 $Y=1.655 $X2=1.955 $Y2=1.51
cc_55 VPB N_VPWR_c_241_n 0.00519718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_233_n 0.0462495f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_Y_c_295_n 0.00322011f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.78
cc_58 N_A1_M1005_g N_A2_c_136_n 0.0311799f $X=0.49 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_59 N_A1_c_61_n N_A2_M1002_g 9.82602e-19 $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_60 N_A1_c_69_n N_A2_M1002_g 0.0150885f $X=1.245 $Y=1.605 $X2=0 $Y2=0
cc_61 N_A1_c_62_n N_A2_M1002_g 0.00451012f $X=1.415 $Y=1.605 $X2=0 $Y2=0
cc_62 N_A1_c_64_n N_A2_M1002_g 0.029366f $X=0.49 $Y=1.46 $X2=0 $Y2=0
cc_63 N_A1_M1010_g N_A2_c_138_n 0.0262407f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_64 N_A1_M1007_g N_A2_M1011_g 0.036142f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_65 N_A1_c_62_n N_A2_M1011_g 0.011304f $X=1.415 $Y=1.605 $X2=0 $Y2=0
cc_66 A1 N_A2_M1011_g 0.0038453f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_67 N_A1_M1005_g N_A2_c_140_n 0.00622359f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_68 N_A1_c_61_n N_A2_c_140_n 0.0112237f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_69 N_A1_c_69_n N_A2_c_140_n 0.0288546f $X=1.245 $Y=1.605 $X2=0 $Y2=0
cc_70 N_A1_c_62_n N_A2_c_140_n 0.0110987f $X=1.415 $Y=1.605 $X2=0 $Y2=0
cc_71 N_A1_M1005_g N_A2_c_141_n 0.0203806f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_72 N_A1_c_69_n N_A2_c_141_n 0.00527565f $X=1.245 $Y=1.605 $X2=0 $Y2=0
cc_73 N_A1_c_62_n N_A2_c_141_n 0.00785233f $X=1.415 $Y=1.605 $X2=0 $Y2=0
cc_74 A1 N_A2_c_141_n 0.00275462f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_75 N_A1_c_65_n N_A2_c_141_n 0.0105172f $X=1.955 $Y=1.51 $X2=0 $Y2=0
cc_76 N_A1_M1010_g N_B1_M1004_g 0.025183f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_77 N_A1_M1007_g N_B1_M1000_g 0.0317236f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_78 A1 N_B1_M1000_g 0.00512908f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_79 A1 N_B1_c_194_n 0.00475316f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_80 N_A1_c_65_n N_B1_c_194_n 0.0213966f $X=1.955 $Y=1.51 $X2=0 $Y2=0
cc_81 N_A1_c_61_n N_VPWR_M1003_d 0.00242003f $X=0.29 $Y=1.46 $X2=-0.19
+ $Y2=-0.245
cc_82 N_A1_M1003_g N_VPWR_c_235_n 0.0180747f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A1_c_61_n N_VPWR_c_235_n 0.0224433f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_84 N_A1_c_64_n N_VPWR_c_235_n 0.00122589f $X=0.49 $Y=1.46 $X2=0 $Y2=0
cc_85 N_A1_M1007_g N_VPWR_c_236_n 0.0125532f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A1_M1003_g N_VPWR_c_239_n 0.00486043f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A1_M1007_g N_VPWR_c_239_n 0.00544582f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_88 N_A1_M1003_g N_VPWR_c_233_n 0.0082726f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A1_M1007_g N_VPWR_c_233_n 0.00966241f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A1_c_69_n N_A_113_367#_M1003_s 0.00176461f $X=1.245 $Y=1.605 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A1_c_69_n N_A_113_367#_c_280_n 0.0135055f $X=1.245 $Y=1.605 $X2=0 $Y2=0
cc_92 N_A1_c_69_n N_Y_M1002_d 0.00176461f $X=1.245 $Y=1.605 $X2=0 $Y2=0
cc_93 N_A1_M1010_g N_Y_c_295_n 5.81725e-19 $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_94 A1 N_Y_c_295_n 0.0320079f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A1_M1007_g N_Y_c_300_n 8.39609e-19 $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A1_c_69_n N_Y_c_300_n 0.0155633f $X=1.245 $Y=1.605 $X2=0 $Y2=0
cc_97 N_A1_c_62_n Y 0.00848929f $X=1.415 $Y=1.605 $X2=0 $Y2=0
cc_98 A1 Y 0.00833648f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_99 N_A1_M1007_g N_Y_c_304_n 0.0207289f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A1_c_65_n N_Y_c_304_n 8.37766e-19 $X=1.955 $Y=1.51 $X2=0 $Y2=0
cc_101 A1 N_Y_c_306_n 0.0545232f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A1_c_61_n N_A_30_47#_c_333_n 0.0113924f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_103 N_A1_c_64_n N_A_30_47#_c_333_n 0.00555768f $X=0.49 $Y=1.46 $X2=0 $Y2=0
cc_104 N_A1_M1005_g N_A_30_47#_c_340_n 0.0133559f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_105 N_A1_c_61_n N_A_30_47#_c_340_n 0.00254549f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_106 N_A1_M1010_g N_A_30_47#_c_335_n 0.0143523f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_107 N_A1_c_62_n N_A_30_47#_c_335_n 0.0519429f $X=1.415 $Y=1.605 $X2=0 $Y2=0
cc_108 A1 N_A_30_47#_c_335_n 0.0280813f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A1_c_65_n N_A_30_47#_c_335_n 0.00425455f $X=1.955 $Y=1.51 $X2=0 $Y2=0
cc_110 N_A1_M1010_g N_A_30_47#_c_346_n 0.00177471f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_111 N_A1_M1010_g N_A_30_47#_c_347_n 0.00884601f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_112 N_A1_M1010_g N_A_30_47#_c_336_n 5.53867e-19 $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_113 N_A1_c_69_n N_A_30_47#_c_336_n 0.0019245f $X=1.245 $Y=1.605 $X2=0 $Y2=0
cc_114 N_A1_c_62_n N_A_30_47#_c_336_n 0.0100406f $X=1.415 $Y=1.605 $X2=0 $Y2=0
cc_115 N_A1_M1005_g N_VGND_c_393_n 0.0116209f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_116 N_A1_M1010_g N_VGND_c_394_n 0.00733525f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_117 N_A1_M1005_g N_VGND_c_395_n 0.00486043f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_118 N_A1_M1010_g N_VGND_c_397_n 0.00562613f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_119 N_A1_M1005_g N_VGND_c_398_n 0.00549807f $X=0.49 $Y=0.655 $X2=0 $Y2=0
cc_120 N_A1_M1010_g N_VGND_c_398_n 0.0106613f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_121 N_A2_M1002_g N_VPWR_c_235_n 0.00109252f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A2_M1011_g N_VPWR_c_236_n 0.00112044f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A2_M1002_g N_VPWR_c_239_n 0.00357877f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A2_M1011_g N_VPWR_c_239_n 0.00357877f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A2_M1002_g N_VPWR_c_233_n 0.00537654f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A2_M1011_g N_VPWR_c_233_n 0.00580255f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A2_M1002_g N_A_113_367#_c_281_n 0.012237f $X=0.92 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A2_M1011_g N_A_113_367#_c_281_n 0.0139882f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A2_M1011_g N_Y_c_300_n 0.00825361f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A2_M1011_g Y 0.0119028f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A2_M1011_g N_Y_c_306_n 0.00331714f $X=1.35 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A2_c_136_n N_A_30_47#_c_340_n 0.0097033f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_133 N_A2_c_140_n N_A_30_47#_c_340_n 0.0265951f $X=0.94 $Y=1.35 $X2=0 $Y2=0
cc_134 N_A2_c_141_n N_A_30_47#_c_340_n 0.00144439f $X=1.35 $Y=1.35 $X2=0 $Y2=0
cc_135 N_A2_c_138_n N_A_30_47#_c_354_n 0.0107276f $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_136 N_A2_c_138_n N_A_30_47#_c_335_n 0.00721602f $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_137 N_A2_c_138_n N_A_30_47#_c_347_n 6.16399e-19 $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_138 N_A2_c_136_n N_A_30_47#_c_336_n 0.00406336f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_139 N_A2_c_138_n N_A_30_47#_c_336_n 0.00728496f $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_140 N_A2_c_141_n N_A_30_47#_c_336_n 0.00444413f $X=1.35 $Y=1.35 $X2=0 $Y2=0
cc_141 N_A2_c_136_n N_VGND_c_393_n 0.0102417f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_142 N_A2_c_138_n N_VGND_c_393_n 6.49123e-19 $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_143 N_A2_c_138_n N_VGND_c_394_n 0.00683397f $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_144 N_A2_c_136_n N_VGND_c_396_n 0.00486043f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_145 N_A2_c_138_n N_VGND_c_396_n 0.00450273f $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_146 N_A2_c_136_n N_VGND_c_398_n 0.00455156f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_147 N_A2_c_138_n N_VGND_c_398_n 0.0080685f $X=1.35 $Y=1.185 $X2=0 $Y2=0
cc_148 N_B1_M1000_g N_VPWR_c_236_n 0.00207663f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_149 N_B1_M1000_g N_VPWR_c_238_n 7.68283e-19 $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_150 N_B1_M1006_g N_VPWR_c_238_n 0.0162756f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_151 B1 N_VPWR_c_238_n 0.0252511f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_152 N_B1_c_194_n N_VPWR_c_238_n 0.00130751f $X=2.835 $Y=1.35 $X2=0 $Y2=0
cc_153 N_B1_M1000_g N_VPWR_c_240_n 0.00583607f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_154 N_B1_M1006_g N_VPWR_c_240_n 0.00564095f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_155 N_B1_M1000_g N_VPWR_c_233_n 0.0106071f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_156 N_B1_M1006_g N_VPWR_c_233_n 0.00948291f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_157 N_B1_M1004_g N_Y_c_295_n 0.00211518f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_158 N_B1_M1000_g N_Y_c_295_n 0.00383795f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B1_c_191_n N_Y_c_295_n 0.00403031f $X=2.835 $Y=1.185 $X2=0 $Y2=0
cc_160 N_B1_M1006_g N_Y_c_295_n 0.00395223f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_161 B1 N_Y_c_295_n 0.0403036f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B1_c_194_n N_Y_c_295_n 0.0193986f $X=2.835 $Y=1.35 $X2=0 $Y2=0
cc_163 N_B1_M1000_g N_Y_c_304_n 0.021149f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_164 N_B1_M1004_g N_A_30_47#_c_335_n 0.00325239f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_165 N_B1_M1004_g N_A_30_47#_c_346_n 5.89773e-19 $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_166 N_B1_M1004_g N_A_30_47#_c_347_n 0.00854791f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_167 N_B1_c_191_n N_A_30_47#_c_347_n 5.54906e-19 $X=2.835 $Y=1.185 $X2=0 $Y2=0
cc_168 N_B1_M1004_g N_A_30_47#_c_364_n 0.0105205f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_169 N_B1_c_191_n N_A_30_47#_c_364_n 0.0118937f $X=2.835 $Y=1.185 $X2=0 $Y2=0
cc_170 N_B1_M1004_g N_A_30_47#_c_337_n 5.41428e-19 $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_171 N_B1_c_191_n N_A_30_47#_c_337_n 0.00797407f $X=2.835 $Y=1.185 $X2=0 $Y2=0
cc_172 B1 N_A_30_47#_c_337_n 0.0239164f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_173 N_B1_c_194_n N_A_30_47#_c_337_n 0.00711154f $X=2.835 $Y=1.35 $X2=0 $Y2=0
cc_174 N_B1_M1004_g N_VGND_c_397_n 0.00357842f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_175 N_B1_c_191_n N_VGND_c_397_n 0.0035787f $X=2.835 $Y=1.185 $X2=0 $Y2=0
cc_176 N_B1_M1004_g N_VGND_c_398_n 0.00537652f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_177 N_B1_c_191_n N_VGND_c_398_n 0.00629143f $X=2.835 $Y=1.185 $X2=0 $Y2=0
cc_178 N_VPWR_c_233_n N_A_113_367#_M1003_s 0.00376625f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_179 N_VPWR_c_233_n N_A_113_367#_M1011_s 0.00543669f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_239_n N_A_113_367#_c_285_n 0.0135879f $X=2 $Y=3.33 $X2=0 $Y2=0
cc_181 N_VPWR_c_233_n N_A_113_367#_c_285_n 0.00855309f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_239_n N_A_113_367#_c_281_n 0.0581994f $X=2 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_233_n N_A_113_367#_c_281_n 0.0356355f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_233_n N_Y_M1002_d 0.00225186f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_185 N_VPWR_c_233_n N_Y_M1000_d 0.00380103f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_186 N_VPWR_c_240_n N_Y_c_319_n 0.0140491f $X=2.905 $Y=3.33 $X2=0 $Y2=0
cc_187 N_VPWR_c_233_n N_Y_c_319_n 0.0090585f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_188 N_VPWR_M1007_d N_Y_c_304_n 0.00434484f $X=2.01 $Y=1.835 $X2=0 $Y2=0
cc_189 N_VPWR_c_236_n N_Y_c_304_n 0.0180329f $X=2.165 $Y=2.49 $X2=0 $Y2=0
cc_190 N_A_113_367#_c_281_n N_Y_M1002_d 0.00332344f $X=1.475 $Y=2.99 $X2=0.49
+ $Y2=0.655
cc_191 N_A_113_367#_c_281_n N_Y_c_300_n 0.0143397f $X=1.475 $Y=2.99 $X2=0 $Y2=0
cc_192 N_A_113_367#_M1011_s Y 0.00270121f $X=1.425 $Y=1.835 $X2=0.29 $Y2=1.78
cc_193 N_A_113_367#_c_292_p Y 0.0267124f $X=1.64 $Y=2.49 $X2=0.29 $Y2=1.78
cc_194 N_A_113_367#_M1011_s N_Y_c_304_n 0.0013787f $X=1.425 $Y=1.835 $X2=0 $Y2=0
cc_195 N_A_113_367#_M1011_s N_Y_c_306_n 0.00580814f $X=1.425 $Y=1.835 $X2=0.29
+ $Y2=1.46
cc_196 N_Y_c_295_n N_A_30_47#_c_335_n 0.0110235f $X=2.62 $Y=0.76 $X2=0 $Y2=0
cc_197 N_Y_M1004_d N_A_30_47#_c_364_n 0.00332344f $X=2.48 $Y=0.235 $X2=0 $Y2=0
cc_198 N_Y_c_295_n N_A_30_47#_c_364_n 0.0126348f $X=2.62 $Y=0.76 $X2=0 $Y2=0
cc_199 N_Y_M1004_d N_VGND_c_398_n 0.00225186f $X=2.48 $Y=0.235 $X2=0 $Y2=0
cc_200 N_A_30_47#_c_340_n N_VGND_M1005_d 0.00344855f $X=1.04 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_201 N_A_30_47#_c_335_n N_VGND_M1009_d 0.00584231f $X=2.035 $Y=1.09 $X2=0
+ $Y2=0
cc_202 N_A_30_47#_c_340_n N_VGND_c_393_n 0.016709f $X=1.04 $Y=0.93 $X2=0 $Y2=0
cc_203 N_A_30_47#_c_354_n N_VGND_c_394_n 0.0441963f $X=1.135 $Y=0.42 $X2=0 $Y2=0
cc_204 N_A_30_47#_c_335_n N_VGND_c_394_n 0.0239317f $X=2.035 $Y=1.09 $X2=0 $Y2=0
cc_205 N_A_30_47#_c_334_n N_VGND_c_395_n 0.0178111f $X=0.275 $Y=0.42 $X2=0 $Y2=0
cc_206 N_A_30_47#_c_354_n N_VGND_c_396_n 0.0201192f $X=1.135 $Y=0.42 $X2=0 $Y2=0
cc_207 N_A_30_47#_c_346_n N_VGND_c_397_n 0.0183782f $X=2.195 $Y=0.425 $X2=0
+ $Y2=0
cc_208 N_A_30_47#_c_364_n N_VGND_c_397_n 0.0310975f $X=2.905 $Y=0.34 $X2=0 $Y2=0
cc_209 N_A_30_47#_c_337_n N_VGND_c_397_n 0.0198231f $X=3.05 $Y=0.42 $X2=0 $Y2=0
cc_210 N_A_30_47#_M1005_s N_VGND_c_398_n 0.00243868f $X=0.15 $Y=0.235 $X2=0
+ $Y2=0
cc_211 N_A_30_47#_M1001_s N_VGND_c_398_n 0.00252268f $X=0.995 $Y=0.235 $X2=0
+ $Y2=0
cc_212 N_A_30_47#_M1010_s N_VGND_c_398_n 0.00223559f $X=2.05 $Y=0.235 $X2=0
+ $Y2=0
cc_213 N_A_30_47#_M1008_s N_VGND_c_398_n 0.00215158f $X=2.91 $Y=0.235 $X2=0
+ $Y2=0
cc_214 N_A_30_47#_c_334_n N_VGND_c_398_n 0.0100304f $X=0.275 $Y=0.42 $X2=0 $Y2=0
cc_215 N_A_30_47#_c_340_n N_VGND_c_398_n 0.0108383f $X=1.04 $Y=0.93 $X2=0 $Y2=0
cc_216 N_A_30_47#_c_354_n N_VGND_c_398_n 0.0120771f $X=1.135 $Y=0.42 $X2=0 $Y2=0
cc_217 N_A_30_47#_c_346_n N_VGND_c_398_n 0.0121115f $X=2.195 $Y=0.425 $X2=0
+ $Y2=0
cc_218 N_A_30_47#_c_364_n N_VGND_c_398_n 0.0194432f $X=2.905 $Y=0.34 $X2=0 $Y2=0
cc_219 N_A_30_47#_c_337_n N_VGND_c_398_n 0.011956f $X=3.05 $Y=0.42 $X2=0 $Y2=0
