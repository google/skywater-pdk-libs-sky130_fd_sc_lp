# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sleep_sergate_plv_14
  CLASS BLOCK ;
  FOREIGN sky130_fd_sc_lp__sleep_sergate_plv_14 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  PIN SLEEP
    ANTENNAGATEAREA  2.100000 ;
    PORT
      LAYER li1 ;
        RECT 8.255000 0.800000 8.785000 2.830000 ;
    END
  END SLEEP
  PIN VIRTPWR
    ANTENNADIFFAREA  3.710000 ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.120000 3.415000 ;
        RECT 1.055000 1.980000 7.950000 2.240000 ;
        RECT 1.055000 2.840000 8.055000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 1.895000 2.025000 2.065000 2.195000 ;
        RECT 1.895000 2.885000 2.065000 3.055000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.255000 2.025000 2.425000 2.195000 ;
        RECT 2.255000 2.885000 2.425000 3.055000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.450000 2.025000 3.620000 2.195000 ;
        RECT 3.450000 2.885000 3.620000 3.055000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.810000 2.025000 3.980000 2.195000 ;
        RECT 3.810000 2.885000 3.980000 3.055000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.005000 2.025000 5.175000 2.195000 ;
        RECT 5.005000 2.885000 5.175000 3.055000 ;
        RECT 5.365000 2.025000 5.535000 2.195000 ;
        RECT 5.365000 2.885000 5.535000 3.055000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.560000 2.025000 6.730000 2.195000 ;
        RECT 6.560000 2.885000 6.730000 3.055000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 6.920000 2.025000 7.090000 2.195000 ;
        RECT 6.920000 2.885000 7.090000 3.055000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
        RECT 1.845000 1.965000 2.470000 3.085000 ;
        RECT 3.400000 1.965000 4.025000 3.085000 ;
        RECT 4.955000 1.965000 5.580000 3.085000 ;
        RECT 6.510000 1.965000 7.155000 3.085000 ;
    END
  END VIRTPWR
  PIN VPWR
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.055000 2.410000 7.950000 2.670000 ;
      LAYER mcon ;
        RECT 1.115000 2.455000 1.285000 2.625000 ;
        RECT 1.475000 2.455000 1.645000 2.625000 ;
        RECT 2.670000 2.455000 2.840000 2.625000 ;
        RECT 3.030000 2.455000 3.200000 2.625000 ;
        RECT 4.225000 2.455000 4.395000 2.625000 ;
        RECT 4.585000 2.455000 4.755000 2.625000 ;
        RECT 5.780000 2.455000 5.950000 2.625000 ;
        RECT 6.140000 2.455000 6.310000 2.625000 ;
        RECT 7.355000 2.455000 7.525000 2.625000 ;
        RECT 7.715000 2.455000 7.885000 2.625000 ;
      LAYER met1 ;
        RECT 1.055000 2.410000 1.705000 2.670000 ;
        RECT 2.610000 2.410000 3.260000 2.670000 ;
        RECT 4.165000 2.410000 4.815000 2.670000 ;
        RECT 5.720000 2.410000 6.370000 2.670000 ;
        RECT 7.295000 2.410000 7.945000 2.670000 ;
      LAYER met2 ;
        RECT 0.280000 0.000000 8.840000 3.330000 ;
      LAYER via ;
        RECT 1.095000 2.410000 1.355000 2.670000 ;
        RECT 1.415000 2.410000 1.675000 2.670000 ;
        RECT 2.640000 2.410000 2.900000 2.670000 ;
        RECT 2.960000 2.410000 3.220000 2.670000 ;
        RECT 4.195000 2.410000 4.455000 2.670000 ;
        RECT 4.515000 2.410000 4.775000 2.670000 ;
        RECT 5.750000 2.410000 6.010000 2.670000 ;
        RECT 6.070000 2.410000 6.330000 2.670000 ;
        RECT 7.325000 2.410000 7.585000 2.670000 ;
        RECT 7.645000 2.410000 7.905000 2.670000 ;
    END
  END VPWR
END sky130_fd_sc_lp__sleep_sergate_plv_14
