* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfrbp_lp CLK D RESET_B VGND VNB VPB VPWR Q Q_N
X0 a_1712_379# a_662_90# a_1799_379# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_560_90# CLK a_2831_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_3036_367# a_1799_379# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_847_116# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1496_111# a_560_90# a_662_90# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND RESET_B a_2493_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_3222_137# a_1799_379# a_3309_137# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_2451_397# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND a_3222_137# a_3490_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_590_116# a_662_90# a_111_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_590_116# a_662_90# a_692_116# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_484_411# a_560_90# a_590_116# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_1301_67# a_590_116# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 a_2185_397# a_1799_379# a_2102_25# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_2825_48# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1712_379# a_2102_25# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VGND a_560_90# a_1496_111# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_1799_379# a_2185_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_692_116# a_817_90# a_847_116# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_817_90# a_662_90# a_1799_379# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 a_817_90# a_590_116# a_1301_373# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_1301_373# a_590_116# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 a_111_457# a_560_90# a_590_116# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR a_560_90# a_1480_413# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_1480_413# a_560_90# a_662_90# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_1037_457# RESET_B a_590_116# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_3309_137# a_1799_379# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VGND a_1799_379# a_3036_48# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_484_411# a_817_90# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_2831_367# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_2000_51# a_2102_25# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VPWR a_1799_379# a_3036_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 a_3222_137# a_1799_379# a_3309_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 a_817_90# a_590_116# a_1301_67# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X34 a_3036_48# a_1799_379# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X35 a_560_90# CLK a_2825_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_349_116# D a_111_457# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_2102_25# RESET_B a_2451_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 a_2493_51# a_1799_379# a_2102_25# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VPWR a_3222_137# a_3490_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X40 a_3490_53# a_3222_137# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X41 a_111_457# RESET_B a_197_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X42 a_197_457# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X43 a_3490_367# a_3222_137# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X44 a_1799_379# a_560_90# a_817_90# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X45 a_3309_367# a_1799_379# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X46 VGND RESET_B a_349_116# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X47 VPWR D a_27_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X48 VPWR RESET_B a_1037_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X49 a_1799_379# a_560_90# a_2000_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X50 a_27_457# D a_111_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
