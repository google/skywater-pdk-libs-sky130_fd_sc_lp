* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_674_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.079e+12p pd=1.338e+07u as=4.914e+11p ps=3.3e+06u
M1001 a_386_51# D1 a_80_21# VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=2.226e+11p ps=2.21e+06u
M1002 a_458_51# C1 a_386_51# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=0p ps=0u
M1003 a_80_21# D1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=8.442e+11p pd=6.38e+06u as=0p ps=0u
M1004 a_80_21# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_80_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=7.728e+11p ps=6.88e+06u
M1006 a_566_51# B1 a_458_51# VNB nshort w=840000u l=150000u
+  ad=5.502e+11p pd=4.67e+06u as=0p ps=0u
M1007 VPWR a_80_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1008 VGND a_80_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_566_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_674_367# A2 a_80_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_566_51# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_80_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR C1 a_80_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
