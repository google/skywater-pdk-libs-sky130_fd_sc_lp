# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__fahcin_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__fahcin_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.460000 1.345000 0.805000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.759000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.660000 1.180000 5.155000 1.670000 ;
    END
  END B
  PIN CIN
    ANTENNAGATEAREA  0.561000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.245000 1.080000 8.575000 1.410000 ;
    END
  END CIN
  PIN COUT
    ANTENNADIFFAREA  1.564400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 0.295000 6.695000 0.440000 ;
        RECT 6.365000 0.440000 7.555000 0.885000 ;
        RECT 6.525000 0.885000 6.695000 1.960000 ;
        RECT 6.525000 1.960000 6.855000 2.715000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.592200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.825000 0.375000 12.370000 1.075000 ;
        RECT 12.120000 1.075000 12.370000 3.065000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 12.480000 0.085000 ;
        RECT  0.635000  0.085000  0.805000 0.815000 ;
        RECT  5.225000  0.085000  5.555000 0.650000 ;
        RECT  8.245000  0.085000  8.575000 0.900000 ;
        RECT 11.315000  0.085000 11.645000 1.075000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.480000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 12.480000 3.415000 ;
        RECT  0.555000 2.055000  0.885000 3.245000 ;
        RECT  5.145000 2.785000  5.475000 3.245000 ;
        RECT  8.495000 1.940000  8.665000 3.245000 ;
        RECT 11.690000 1.855000 11.940000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 12.480000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.110000 0.265000  0.455000 0.995000 ;
      RECT  0.110000 0.995000  1.155000 1.165000 ;
      RECT  0.110000 1.165000  0.280000 1.960000 ;
      RECT  0.110000 1.960000  0.375000 3.065000 ;
      RECT  0.985000 0.265000  2.570000 0.435000 ;
      RECT  0.985000 0.435000  1.155000 0.995000 ;
      RECT  0.985000 1.165000  1.155000 1.205000 ;
      RECT  0.985000 1.205000  1.360000 1.875000 ;
      RECT  1.065000 1.875000  1.235000 2.895000 ;
      RECT  1.065000 2.895000  3.675000 3.065000 ;
      RECT  1.335000 0.615000  1.585000 0.855000 ;
      RECT  1.335000 0.855000  2.920000 1.025000 ;
      RECT  1.415000 2.055000  1.665000 2.545000 ;
      RECT  1.415000 2.545000  2.665000 2.715000 ;
      RECT  1.565000 1.550000  2.155000 1.780000 ;
      RECT  1.785000 1.205000  2.155000 1.550000 ;
      RECT  1.905000 1.780000  2.155000 2.365000 ;
      RECT  2.320000 0.435000  2.570000 0.675000 ;
      RECT  2.335000 1.025000  2.665000 2.545000 ;
      RECT  2.750000 0.265000  3.700000 0.435000 ;
      RECT  2.750000 0.435000  2.920000 0.855000 ;
      RECT  2.880000 1.875000  3.270000 1.960000 ;
      RECT  2.880000 1.960000  4.025000 2.130000 ;
      RECT  2.880000 2.130000  3.270000 2.715000 ;
      RECT  3.100000 0.615000  3.270000 1.875000 ;
      RECT  3.450000 0.435000  3.700000 1.020000 ;
      RECT  3.450000 1.200000  4.050000 1.370000 ;
      RECT  3.450000 1.370000  3.780000 1.705000 ;
      RECT  3.505000 2.310000  3.675000 2.895000 ;
      RECT  3.855000 2.130000  4.025000 2.895000 ;
      RECT  3.855000 2.895000  4.965000 3.065000 ;
      RECT  3.880000 0.265000  5.045000 0.435000 ;
      RECT  3.880000 0.435000  4.050000 1.200000 ;
      RECT  3.965000 1.550000  4.480000 1.780000 ;
      RECT  4.205000 1.780000  4.480000 2.715000 ;
      RECT  4.230000 0.615000  4.480000 1.550000 ;
      RECT  4.715000 0.435000  5.045000 0.830000 ;
      RECT  4.715000 0.830000  5.635000 1.000000 ;
      RECT  4.715000 1.850000  5.635000 2.020000 ;
      RECT  4.715000 2.020000  5.045000 2.255000 ;
      RECT  4.795000 2.435000  6.345000 2.605000 ;
      RECT  4.795000 2.605000  4.965000 2.895000 ;
      RECT  5.380000 1.000000  5.635000 1.850000 ;
      RECT  5.815000 0.295000  6.185000 0.975000 ;
      RECT  5.815000 0.975000  5.985000 2.255000 ;
      RECT  6.165000 1.455000  6.345000 2.435000 ;
      RECT  6.165000 2.605000  6.345000 2.895000 ;
      RECT  6.165000 2.895000  8.315000 3.065000 ;
      RECT  6.875000 1.065000  7.140000 1.395000 ;
      RECT  6.875000 1.395000  7.075000 1.780000 ;
      RECT  7.265000 1.575000  7.615000 1.745000 ;
      RECT  7.265000 1.745000  7.435000 2.895000 ;
      RECT  7.350000 1.115000  7.615000 1.575000 ;
      RECT  7.615000 1.925000  7.965000 2.715000 ;
      RECT  7.735000 0.295000  8.065000 0.935000 ;
      RECT  7.795000 0.935000  7.965000 1.925000 ;
      RECT  8.145000 1.590000  8.925000 1.760000 ;
      RECT  8.145000 1.760000  8.315000 2.895000 ;
      RECT  8.755000 0.265000  9.775000 0.565000 ;
      RECT  8.755000 0.565000  8.925000 1.590000 ;
      RECT  8.845000 1.940000  9.290000 2.895000 ;
      RECT  8.845000 2.895000 11.510000 3.065000 ;
      RECT  9.120000 0.745000  9.505000 1.335000 ;
      RECT  9.120000 1.335000  9.290000 1.940000 ;
      RECT  9.470000 2.385000 11.160000 2.555000 ;
      RECT  9.470000 2.555000  9.720000 2.715000 ;
      RECT  9.755000 1.135000 10.205000 1.305000 ;
      RECT  9.755000 1.305000  9.925000 2.035000 ;
      RECT  9.755000 2.035000 10.150000 2.205000 ;
      RECT  9.955000 0.265000 11.135000 0.435000 ;
      RECT  9.955000 0.435000 10.205000 1.135000 ;
      RECT 10.105000 1.485000 10.435000 1.815000 ;
      RECT 10.360000 2.735000 10.690000 2.895000 ;
      RECT 10.420000 0.615000 10.785000 1.305000 ;
      RECT 10.615000 1.305000 10.785000 2.205000 ;
      RECT 10.615000 2.205000 11.160000 2.385000 ;
      RECT 10.910000 2.555000 11.160000 2.715000 ;
      RECT 10.965000 0.435000 11.135000 1.255000 ;
      RECT 10.965000 1.255000 11.940000 1.425000 ;
      RECT 11.035000 1.605000 11.365000 1.855000 ;
      RECT 11.035000 1.855000 11.510000 2.025000 ;
      RECT 11.340000 2.025000 11.510000 2.895000 ;
      RECT 11.610000 1.425000 11.940000 1.675000 ;
    LAYER mcon ;
      RECT  1.595000 1.580000  1.765000 1.750000 ;
      RECT  3.995000 1.580000  4.165000 1.750000 ;
      RECT  6.875000 1.580000  7.045000 1.750000 ;
      RECT 10.235000 1.580000 10.405000 1.750000 ;
    LAYER met1 ;
      RECT  1.535000 1.550000  1.825000 1.595000 ;
      RECT  1.535000 1.595000 10.465000 1.735000 ;
      RECT  1.535000 1.735000  1.825000 1.780000 ;
      RECT  3.935000 1.550000  4.225000 1.595000 ;
      RECT  3.935000 1.735000  4.225000 1.780000 ;
      RECT  6.815000 1.550000  7.105000 1.595000 ;
      RECT  6.815000 1.735000  7.105000 1.780000 ;
      RECT 10.175000 1.550000 10.465000 1.595000 ;
      RECT 10.175000 1.735000 10.465000 1.780000 ;
  END
END sky130_fd_sc_lp__fahcin_1
