# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__or4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__or4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.345000 2.315000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.385000 1.920000 2.855000 2.940000 ;
        RECT 2.485000 1.345000 2.855000 1.920000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.025000 1.345000 3.685000 2.940000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.730000 1.535000 5.195000 2.205000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.005000 0.790000 1.175000 ;
        RECT 0.090000 1.175000 0.335000 1.695000 ;
        RECT 0.090000 1.695000 1.715000 1.865000 ;
        RECT 0.610000 0.255000 0.800000 0.655000 ;
        RECT 0.610000 0.655000 1.680000 0.825000 ;
        RECT 0.610000 0.825000 0.790000 1.005000 ;
        RECT 0.610000 1.865000 0.800000 3.075000 ;
        RECT 1.470000 0.485000 1.680000 0.655000 ;
        RECT 1.470000 1.865000 1.715000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.110000  0.085000 0.440000 0.835000 ;
      RECT 0.110000  2.035000 0.440000 3.245000 ;
      RECT 0.505000  1.355000 1.905000 1.525000 ;
      RECT 0.970000  0.085000 1.300000 0.485000 ;
      RECT 0.970000  2.035000 1.300000 3.245000 ;
      RECT 1.735000  0.995000 3.760000 1.005000 ;
      RECT 1.735000  1.005000 4.035000 1.175000 ;
      RECT 1.735000  1.175000 1.905000 1.355000 ;
      RECT 1.850000  0.085000 2.180000 0.825000 ;
      RECT 1.885000  1.920000 2.215000 3.245000 ;
      RECT 2.350000  0.255000 2.560000 0.995000 ;
      RECT 2.730000  0.085000 3.400000 0.825000 ;
      RECT 3.570000  0.255000 3.760000 0.995000 ;
      RECT 3.855000  1.175000 4.035000 1.815000 ;
      RECT 3.855000  1.815000 4.090000 3.075000 ;
      RECT 3.930000  0.085000 4.700000 0.835000 ;
      RECT 4.205000  0.835000 4.700000 1.015000 ;
      RECT 4.215000  1.185000 5.130000 1.355000 ;
      RECT 4.215000  1.355000 4.560000 1.515000 ;
      RECT 4.260000  1.515000 4.560000 2.375000 ;
      RECT 4.260000  2.375000 5.185000 2.545000 ;
      RECT 4.425000  2.715000 4.755000 3.245000 ;
      RECT 4.870000  0.700000 5.130000 1.185000 ;
      RECT 4.925000  2.545000 5.185000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_lp__or4b_4
END LIBRARY
