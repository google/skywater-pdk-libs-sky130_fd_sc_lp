* File: sky130_fd_sc_lp__decap_4.pxi.spice
* Created: Wed Sep  2 09:42:00 2020
* 
x_PM_SKY130_FD_SC_LP__DECAP_4%VGND N_VGND_M1001_s N_VGND_c_23_n N_VGND_M1000_g
+ N_VGND_c_24_n N_VGND_c_25_n N_VGND_c_26_n N_VGND_c_27_n N_VGND_c_28_n VGND
+ N_VGND_c_29_n N_VGND_c_30_n PM_SKY130_FD_SC_LP__DECAP_4%VGND
x_PM_SKY130_FD_SC_LP__DECAP_4%VPWR N_VPWR_M1000_s N_VPWR_c_53_n N_VPWR_c_54_n
+ N_VPWR_c_55_n N_VPWR_c_56_n N_VPWR_c_50_n VPWR N_VPWR_M1001_g N_VPWR_c_59_n
+ N_VPWR_c_52_n PM_SKY130_FD_SC_LP__DECAP_4%VPWR
cc_1 VNB N_VGND_c_23_n 0.0113126f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.935
cc_2 VNB N_VGND_c_24_n 0.012758f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.085
cc_3 VNB N_VGND_c_25_n 0.0607496f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.38
cc_4 VNB N_VGND_c_26_n 0.0118011f $X=-0.19 $Y=-0.245 $X2=1.615 $Y2=0.085
cc_5 VNB N_VGND_c_27_n 0.0371702f $X=-0.19 $Y=-0.245 $X2=1.615 $Y2=0.36
cc_6 VNB N_VGND_c_28_n 0.00314375f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.77
cc_7 VNB N_VGND_c_29_n 0.0280737f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0
cc_8 VNB N_VGND_c_30_n 0.132299f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0
cc_9 VNB N_VPWR_c_50_n 0.0248034f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=1.77
cc_10 VNB N_VPWR_M1001_g 0.123316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_VPWR_c_52_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=0
cc_12 VPB N_VGND_c_23_n 0.0464251f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.935
cc_13 VPB N_VGND_M1000_g 0.0850668f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.595
cc_14 VPB N_VGND_c_28_n 0.0173225f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.77
cc_15 VPB N_VPWR_c_53_n 0.0103989f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.935
cc_16 VPB N_VPWR_c_54_n 0.0425694f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.595
cc_17 VPB N_VPWR_c_55_n 0.0138486f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.38
cc_18 VPB N_VPWR_c_56_n 0.060805f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=1.06
cc_19 VPB N_VPWR_c_50_n 0.00154239f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=1.77
cc_20 VPB N_VPWR_M1001_g 0.00822137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_21 VPB N_VPWR_c_59_n 0.0283919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_52_n 0.047818f $X=-0.19 $Y=1.655 $X2=1.685 $Y2=0
cc_23 N_VGND_M1000_g N_VPWR_c_54_n 0.0546012f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_24 N_VGND_c_28_n N_VPWR_c_54_n 0.0192408f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_25 N_VGND_c_23_n N_VPWR_c_56_n 0.00391118f $X=0.91 $Y=1.935 $X2=0 $Y2=0
cc_26 N_VGND_M1000_g N_VPWR_c_56_n 0.0672708f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_27 N_VGND_c_28_n N_VPWR_c_56_n 0.00754551f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_28 N_VGND_c_23_n N_VPWR_c_50_n 0.00168112f $X=0.91 $Y=1.935 $X2=0 $Y2=0
cc_29 N_VGND_c_27_n N_VPWR_c_50_n 0.0168265f $X=1.615 $Y=0.36 $X2=0 $Y2=0
cc_30 N_VGND_c_28_n N_VPWR_c_50_n 0.00256852f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_31 N_VGND_c_23_n N_VPWR_M1001_g 0.0523192f $X=0.91 $Y=1.935 $X2=0 $Y2=0
cc_32 N_VGND_c_25_n N_VPWR_M1001_g 0.0687615f $X=0.335 $Y=0.38 $X2=0 $Y2=0
cc_33 N_VGND_c_27_n N_VPWR_M1001_g 0.0510153f $X=1.615 $Y=0.36 $X2=0 $Y2=0
cc_34 N_VGND_c_28_n N_VPWR_M1001_g 0.00192223f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_35 N_VGND_c_29_n N_VPWR_M1001_g 0.0370388f $X=1.45 $Y=0 $X2=0 $Y2=0
cc_36 N_VGND_c_30_n N_VPWR_M1001_g 0.0582443f $X=1.68 $Y=0 $X2=0 $Y2=0
cc_37 N_VGND_M1000_g N_VPWR_c_59_n 0.0374291f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_38 N_VGND_M1000_g N_VPWR_c_52_n 0.0588621f $X=0.91 $Y=2.595 $X2=0 $Y2=0
