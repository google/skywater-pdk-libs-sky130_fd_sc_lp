* File: sky130_fd_sc_lp__o221a_4.pxi.spice
* Created: Wed Sep  2 10:18:29 2020
* 
x_PM_SKY130_FD_SC_LP__O221A_4%C1 N_C1_c_119_n N_C1_M1005_g N_C1_M1006_g
+ N_C1_c_121_n N_C1_M1014_g N_C1_M1022_g C1 C1 N_C1_c_124_n
+ PM_SKY130_FD_SC_LP__O221A_4%C1
x_PM_SKY130_FD_SC_LP__O221A_4%B1 N_B1_M1015_g N_B1_M1000_g N_B1_c_163_n
+ N_B1_M1023_g N_B1_M1026_g N_B1_c_165_n N_B1_c_166_n N_B1_c_167_n B1 B1
+ N_B1_c_169_n N_B1_c_170_n N_B1_c_171_n PM_SKY130_FD_SC_LP__O221A_4%B1
x_PM_SKY130_FD_SC_LP__O221A_4%B2 N_B2_M1003_g N_B2_M1009_g N_B2_M1020_g
+ N_B2_M1018_g B2 B2 N_B2_c_253_n PM_SKY130_FD_SC_LP__O221A_4%B2
x_PM_SKY130_FD_SC_LP__O221A_4%A1 N_A1_M1007_g N_A1_M1002_g N_A1_M1011_g
+ N_A1_M1008_g N_A1_c_302_n N_A1_c_303_n A1 N_A1_c_304_n N_A1_c_305_n
+ N_A1_c_306_n N_A1_c_307_n N_A1_c_308_n PM_SKY130_FD_SC_LP__O221A_4%A1
x_PM_SKY130_FD_SC_LP__O221A_4%A2 N_A2_M1016_g N_A2_M1010_g N_A2_M1027_g
+ N_A2_M1017_g A2 N_A2_c_387_n N_A2_c_388_n PM_SKY130_FD_SC_LP__O221A_4%A2
x_PM_SKY130_FD_SC_LP__O221A_4%A_112_65# N_A_112_65#_M1005_d N_A_112_65#_M1006_s
+ N_A_112_65#_M1009_s N_A_112_65#_M1016_s N_A_112_65#_M1004_g
+ N_A_112_65#_M1001_g N_A_112_65#_M1012_g N_A_112_65#_M1013_g
+ N_A_112_65#_M1021_g N_A_112_65#_M1019_g N_A_112_65#_M1024_g
+ N_A_112_65#_M1025_g N_A_112_65#_c_453_n N_A_112_65#_c_442_n
+ N_A_112_65#_c_523_p N_A_112_65#_c_461_n N_A_112_65#_c_472_n
+ N_A_112_65#_c_490_n N_A_112_65#_c_443_n N_A_112_65#_c_444_n
+ N_A_112_65#_c_550_p N_A_112_65#_c_462_n N_A_112_65#_c_464_n
+ N_A_112_65#_c_475_n N_A_112_65#_c_497_n N_A_112_65#_c_445_n
+ PM_SKY130_FD_SC_LP__O221A_4%A_112_65#
x_PM_SKY130_FD_SC_LP__O221A_4%VPWR N_VPWR_M1006_d N_VPWR_M1022_d N_VPWR_M1026_s
+ N_VPWR_M1011_d N_VPWR_M1013_s N_VPWR_M1025_s N_VPWR_c_594_n N_VPWR_c_595_n
+ N_VPWR_c_596_n N_VPWR_c_597_n N_VPWR_c_598_n N_VPWR_c_599_n N_VPWR_c_600_n
+ N_VPWR_c_601_n VPWR N_VPWR_c_602_n N_VPWR_c_603_n N_VPWR_c_604_n
+ N_VPWR_c_605_n N_VPWR_c_606_n N_VPWR_c_607_n N_VPWR_c_608_n N_VPWR_c_609_n
+ N_VPWR_c_610_n N_VPWR_c_593_n PM_SKY130_FD_SC_LP__O221A_4%VPWR
x_PM_SKY130_FD_SC_LP__O221A_4%A_292_367# N_A_292_367#_M1000_d
+ N_A_292_367#_M1018_d N_A_292_367#_c_698_n N_A_292_367#_c_694_n
+ N_A_292_367#_c_706_n N_A_292_367#_c_701_n
+ PM_SKY130_FD_SC_LP__O221A_4%A_292_367#
x_PM_SKY130_FD_SC_LP__O221A_4%A_726_367# N_A_726_367#_M1007_s
+ N_A_726_367#_M1027_d N_A_726_367#_c_714_n N_A_726_367#_c_708_n
+ N_A_726_367#_c_722_n N_A_726_367#_c_709_n
+ PM_SKY130_FD_SC_LP__O221A_4%A_726_367#
x_PM_SKY130_FD_SC_LP__O221A_4%X N_X_M1004_s N_X_M1021_s N_X_M1001_d N_X_M1019_d
+ N_X_c_779_p N_X_c_765_n N_X_c_724_n N_X_c_725_n N_X_c_730_n N_X_c_731_n
+ N_X_c_780_p N_X_c_769_n N_X_c_726_n N_X_c_732_n N_X_c_727_n N_X_c_733_n X X
+ N_X_c_728_n X PM_SKY130_FD_SC_LP__O221A_4%X
x_PM_SKY130_FD_SC_LP__O221A_4%A_29_65# N_A_29_65#_M1005_s N_A_29_65#_M1014_s
+ N_A_29_65#_M1003_s N_A_29_65#_M1023_d N_A_29_65#_c_785_n N_A_29_65#_c_786_n
+ N_A_29_65#_c_787_n N_A_29_65#_c_788_n N_A_29_65#_c_789_n N_A_29_65#_c_790_n
+ PM_SKY130_FD_SC_LP__O221A_4%A_29_65#
x_PM_SKY130_FD_SC_LP__O221A_4%A_284_65# N_A_284_65#_M1015_s N_A_284_65#_M1020_d
+ N_A_284_65#_M1002_d N_A_284_65#_M1017_s N_A_284_65#_c_828_n
+ N_A_284_65#_c_823_n N_A_284_65#_c_824_n N_A_284_65#_c_832_n
+ N_A_284_65#_c_825_n PM_SKY130_FD_SC_LP__O221A_4%A_284_65#
x_PM_SKY130_FD_SC_LP__O221A_4%VGND N_VGND_M1002_s N_VGND_M1010_d N_VGND_M1008_s
+ N_VGND_M1012_d N_VGND_M1024_d N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n
+ N_VGND_c_870_n N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n N_VGND_c_874_n
+ N_VGND_c_875_n N_VGND_c_876_n N_VGND_c_877_n VGND N_VGND_c_878_n
+ N_VGND_c_879_n N_VGND_c_880_n N_VGND_c_881_n N_VGND_c_882_n
+ PM_SKY130_FD_SC_LP__O221A_4%VGND
cc_1 VNB N_C1_c_119_n 0.0201642f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.275
cc_2 VNB N_C1_M1006_g 0.00302368f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_3 VNB N_C1_c_121_n 0.0159488f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.275
cc_4 VNB N_C1_M1022_g 0.00244346f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_5 VNB C1 0.0200912f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_C1_c_124_n 0.0700533f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.44
cc_7 VNB N_B1_M1000_g 0.00272569f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_8 VNB N_B1_c_163_n 0.0189449f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.275
cc_9 VNB N_B1_M1026_g 0.00374192f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=2.465
cc_10 VNB N_B1_c_165_n 0.0111937f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_B1_c_166_n 0.00347631f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.44
cc_12 VNB N_B1_c_167_n 0.0528012f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.44
cc_13 VNB B1 0.00966285f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.44
cc_14 VNB N_B1_c_169_n 0.0283247f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.44
cc_15 VNB N_B1_c_170_n 0.0162867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_171_n 0.00226644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B2_M1003_g 0.0188655f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.745
cc_18 VNB N_B2_M1020_g 0.0192608f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.605
cc_19 VNB B2 0.00265344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B2_c_253_n 0.0297064f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.295
cc_21 VNB N_A1_M1007_g 0.00905845f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.745
cc_22 VNB N_A1_M1011_g 0.00817833f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.745
cc_23 VNB N_A1_c_302_n 0.00316391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_303_n 0.0344468f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.44
cc_25 VNB N_A1_c_304_n 0.0187962f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.295
cc_26 VNB N_A1_c_305_n 0.0309724f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.665
cc_27 VNB N_A1_c_306_n 0.00893373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A1_c_307_n 0.0157574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A1_c_308_n 0.0161904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A2_M1010_g 0.0228946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_M1017_g 0.0218553f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_32 VNB N_A2_c_387_n 0.00310799f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.44
cc_33 VNB N_A2_c_388_n 0.0347114f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.44
cc_34 VNB N_A_112_65#_M1004_g 0.0236724f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_35 VNB N_A_112_65#_M1012_g 0.0219214f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.44
cc_36 VNB N_A_112_65#_M1021_g 0.0219009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_112_65#_M1024_g 0.0264632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_112_65#_c_442_n 0.00114144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_112_65#_c_443_n 7.22757e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_112_65#_c_444_n 0.0036682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_112_65#_c_445_n 0.0733449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_593_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_724_n 0.00304888f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.44
cc_44 VNB N_X_c_725_n 0.00341938f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.44
cc_45 VNB N_X_c_726_n 0.00172363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_X_c_727_n 0.00144499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_X_c_728_n 0.0106328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB X 0.0225555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_29_65#_c_785_n 0.0233564f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_50 VNB N_A_29_65#_c_786_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_29_65#_c_787_n 0.00928796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_29_65#_c_788_n 0.00166139f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.295
cc_53 VNB N_A_29_65#_c_789_n 0.00556476f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.44
cc_54 VNB N_A_29_65#_c_790_n 0.00632187f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.665
cc_55 VNB N_A_284_65#_c_823_n 0.00499622f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.44
cc_56 VNB N_A_284_65#_c_824_n 0.00268692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_284_65#_c_825_n 0.00304778f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.44
cc_58 VNB N_VGND_c_867_n 0.00596559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_868_n 3.20903e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_869_n 0.0163414f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.44
cc_61 VNB N_VGND_c_870_n 0.00397364f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.44
cc_62 VNB N_VGND_c_871_n 3.16049e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_872_n 0.0119606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_873_n 0.0269916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_874_n 0.0761852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_875_n 0.00510557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_876_n 0.0126883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_877_n 0.00436584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_878_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_879_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_880_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_881_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_882_n 0.36665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VPB N_C1_M1006_g 0.0244731f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_75 VPB N_C1_M1022_g 0.0196313f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_76 VPB C1 0.00855959f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_77 VPB N_B1_M1000_g 0.0207397f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_78 VPB N_B1_M1026_g 0.0266837f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_79 VPB N_B2_M1009_g 0.0190473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_B2_M1018_g 0.0182425f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_81 VPB B2 0.00519067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_B2_c_253_n 0.00472401f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.295
cc_83 VPB N_A1_M1007_g 0.0272659f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.745
cc_84 VPB N_A1_M1011_g 0.022018f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.745
cc_85 VPB N_A2_M1016_g 0.0182325f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.745
cc_86 VPB N_A2_M1027_g 0.0190448f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.605
cc_87 VPB N_A2_c_387_n 0.00466831f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.44
cc_88 VPB N_A2_c_388_n 0.00475123f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.44
cc_89 VPB N_A_112_65#_M1001_g 0.0205786f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.44
cc_90 VPB N_A_112_65#_M1013_g 0.0188559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_112_65#_M1019_g 0.0188421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_112_65#_M1025_g 0.0224142f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_112_65#_c_442_n 0.00130642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_112_65#_c_443_n 0.00188545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_112_65#_c_445_n 0.00721304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_594_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.44
cc_97 VPB N_VPWR_c_595_n 0.0469092f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.44
cc_98 VPB N_VPWR_c_596_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_597_n 0.00253106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_598_n 0.00498595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_599_n 3.20903e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_600_n 0.0108182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_601_n 0.0412086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_602_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_603_n 0.0323803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_604_n 0.0345906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_605_n 0.0162141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_606_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_607_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_608_n 0.0125509f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_609_n 0.00631973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_610_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_593_n 0.0450291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_X_c_730_n 0.00304705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_X_c_731_n 0.00202795f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.295
cc_116 VPB N_X_c_732_n 0.010425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_X_c_733_n 0.00144314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB X 0.00506177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 N_C1_M1022_g N_B1_M1000_g 0.0345124f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_120 N_C1_c_121_n B1 0.00338708f $X=0.915 $Y=1.275 $X2=0 $Y2=0
cc_121 N_C1_c_124_n N_B1_c_169_n 0.0215828f $X=0.915 $Y=1.44 $X2=0 $Y2=0
cc_122 N_C1_c_121_n N_B1_c_170_n 0.0176319f $X=0.915 $Y=1.275 $X2=0 $Y2=0
cc_123 N_C1_c_119_n N_A_112_65#_c_453_n 0.00441594f $X=0.485 $Y=1.275 $X2=0
+ $Y2=0
cc_124 N_C1_c_121_n N_A_112_65#_c_453_n 0.0041768f $X=0.915 $Y=1.275 $X2=0 $Y2=0
cc_125 N_C1_c_119_n N_A_112_65#_c_442_n 0.00172473f $X=0.485 $Y=1.275 $X2=0
+ $Y2=0
cc_126 N_C1_M1006_g N_A_112_65#_c_442_n 0.00261835f $X=0.485 $Y=2.465 $X2=0
+ $Y2=0
cc_127 N_C1_c_121_n N_A_112_65#_c_442_n 0.00280302f $X=0.915 $Y=1.275 $X2=0
+ $Y2=0
cc_128 N_C1_M1022_g N_A_112_65#_c_442_n 0.00807208f $X=0.915 $Y=2.465 $X2=0
+ $Y2=0
cc_129 C1 N_A_112_65#_c_442_n 0.0409404f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_130 N_C1_c_124_n N_A_112_65#_c_442_n 0.0202524f $X=0.915 $Y=1.44 $X2=0 $Y2=0
cc_131 N_C1_M1022_g N_A_112_65#_c_461_n 0.0149388f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_132 N_C1_c_119_n N_A_112_65#_c_462_n 0.00635526f $X=0.485 $Y=1.275 $X2=0
+ $Y2=0
cc_133 N_C1_c_121_n N_A_112_65#_c_462_n 0.00301443f $X=0.915 $Y=1.275 $X2=0
+ $Y2=0
cc_134 N_C1_M1022_g N_A_112_65#_c_464_n 0.00157824f $X=0.915 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_C1_M1006_g N_VPWR_c_595_n 0.0193679f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_136 N_C1_M1022_g N_VPWR_c_595_n 7.33921e-19 $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_137 C1 N_VPWR_c_595_n 0.026901f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_138 N_C1_c_124_n N_VPWR_c_595_n 0.0014558f $X=0.915 $Y=1.44 $X2=0 $Y2=0
cc_139 N_C1_M1006_g N_VPWR_c_596_n 6.51893e-19 $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_140 N_C1_M1022_g N_VPWR_c_596_n 0.0128331f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_141 N_C1_M1006_g N_VPWR_c_602_n 0.00486043f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_142 N_C1_M1022_g N_VPWR_c_602_n 0.00564095f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_143 N_C1_M1006_g N_VPWR_c_593_n 0.00824727f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_144 N_C1_M1022_g N_VPWR_c_593_n 0.00948291f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_145 C1 N_A_29_65#_c_785_n 0.0226419f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_146 N_C1_c_124_n N_A_29_65#_c_785_n 0.00190643f $X=0.915 $Y=1.44 $X2=0 $Y2=0
cc_147 N_C1_c_119_n N_A_29_65#_c_786_n 0.0125492f $X=0.485 $Y=1.275 $X2=0 $Y2=0
cc_148 N_C1_c_121_n N_A_29_65#_c_786_n 0.0119687f $X=0.915 $Y=1.275 $X2=0 $Y2=0
cc_149 N_C1_c_119_n N_VGND_c_874_n 0.00302501f $X=0.485 $Y=1.275 $X2=0 $Y2=0
cc_150 N_C1_c_121_n N_VGND_c_874_n 0.00302501f $X=0.915 $Y=1.275 $X2=0 $Y2=0
cc_151 N_C1_c_119_n N_VGND_c_882_n 0.004709f $X=0.485 $Y=1.275 $X2=0 $Y2=0
cc_152 N_C1_c_121_n N_VGND_c_882_n 0.00435646f $X=0.915 $Y=1.275 $X2=0 $Y2=0
cc_153 N_B1_c_165_n N_B2_M1003_g 0.00709446f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_154 N_B1_c_169_n N_B2_M1003_g 0.0214236f $X=1.365 $Y=1.44 $X2=0 $Y2=0
cc_155 N_B1_c_170_n N_B2_M1003_g 0.0266409f $X=1.365 $Y=1.275 $X2=0 $Y2=0
cc_156 N_B1_c_171_n N_B2_M1003_g 0.00733923f $X=1.82 $Y=1.34 $X2=0 $Y2=0
cc_157 N_B1_c_163_n N_B2_M1020_g 0.0292949f $X=2.675 $Y=1.275 $X2=0 $Y2=0
cc_158 N_B1_c_165_n N_B2_M1020_g 0.0104702f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_159 N_B1_c_166_n N_B2_M1020_g 5.85731e-19 $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_160 N_B1_c_171_n N_B2_M1020_g 5.31765e-19 $X=1.82 $Y=1.34 $X2=0 $Y2=0
cc_161 N_B1_M1026_g N_B2_M1018_g 0.0292949f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_162 N_B1_M1000_g B2 2.693e-19 $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_163 N_B1_M1026_g B2 0.0122399f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_164 N_B1_c_165_n B2 0.0537867f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B1_c_166_n B2 0.0140075f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_166 N_B1_c_167_n B2 0.00892545f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_167 N_B1_c_171_n B2 0.0150679f $X=1.82 $Y=1.34 $X2=0 $Y2=0
cc_168 N_B1_M1000_g N_B2_c_253_n 0.0397983f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_169 N_B1_c_165_n N_B2_c_253_n 0.00260948f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B1_c_167_n N_B2_c_253_n 0.0292949f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_171 N_B1_c_171_n N_B2_c_253_n 0.0124852f $X=1.82 $Y=1.34 $X2=0 $Y2=0
cc_172 N_B1_c_166_n N_A1_M1007_g 5.44356e-19 $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_173 N_B1_c_167_n N_A1_M1007_g 0.00384431f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_174 N_B1_c_163_n N_A1_c_302_n 4.14348e-19 $X=2.675 $Y=1.275 $X2=0 $Y2=0
cc_175 N_B1_c_165_n N_A1_c_302_n 0.0124644f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_176 N_B1_c_166_n N_A1_c_302_n 0.016491f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_177 N_B1_c_167_n N_A1_c_302_n 9.31734e-19 $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_178 N_B1_c_163_n N_A1_c_303_n 0.00107883f $X=2.675 $Y=1.275 $X2=0 $Y2=0
cc_179 N_B1_c_165_n N_A1_c_303_n 6.401e-19 $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_180 N_B1_c_166_n N_A1_c_303_n 0.00114031f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_181 N_B1_c_167_n N_A1_c_303_n 0.014794f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_182 N_B1_c_165_n N_A1_c_304_n 5.81256e-19 $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_183 N_B1_c_170_n N_A_112_65#_c_453_n 0.00118912f $X=1.365 $Y=1.275 $X2=0
+ $Y2=0
cc_184 N_B1_M1000_g N_A_112_65#_c_442_n 0.00155491f $X=1.385 $Y=2.465 $X2=0
+ $Y2=0
cc_185 B1 N_A_112_65#_c_442_n 0.03257f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_186 N_B1_c_169_n N_A_112_65#_c_442_n 2.50314e-19 $X=1.365 $Y=1.44 $X2=0 $Y2=0
cc_187 N_B1_M1000_g N_A_112_65#_c_461_n 0.0158967f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_188 B1 N_A_112_65#_c_461_n 0.0329229f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_189 N_B1_c_169_n N_A_112_65#_c_461_n 0.00341407f $X=1.365 $Y=1.44 $X2=0 $Y2=0
cc_190 N_B1_M1026_g N_A_112_65#_c_472_n 0.0167919f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B1_c_166_n N_A_112_65#_c_472_n 0.0115787f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_192 N_B1_c_167_n N_A_112_65#_c_472_n 0.00565263f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_193 N_B1_M1000_g N_A_112_65#_c_475_n 8.92984e-19 $X=1.385 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_B1_M1026_g N_A_112_65#_c_475_n 8.92984e-19 $X=2.675 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_B1_M1000_g N_VPWR_c_596_n 0.0139395f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_196 N_B1_M1026_g N_VPWR_c_597_n 0.0194393f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_197 N_B1_M1000_g N_VPWR_c_603_n 0.00564095f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_198 N_B1_M1026_g N_VPWR_c_603_n 0.00486043f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_199 N_B1_M1000_g N_VPWR_c_593_n 0.00950825f $X=1.385 $Y=2.465 $X2=0 $Y2=0
cc_200 N_B1_M1026_g N_VPWR_c_593_n 0.0082726f $X=2.675 $Y=2.465 $X2=0 $Y2=0
cc_201 N_B1_c_165_n N_A_29_65#_M1003_s 0.00176891f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B1_c_165_n N_A_29_65#_M1023_d 0.00232777f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_203 B1 N_A_29_65#_c_788_n 0.0137135f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_204 N_B1_c_169_n N_A_29_65#_c_788_n 2.59249e-19 $X=1.365 $Y=1.44 $X2=0 $Y2=0
cc_205 N_B1_c_163_n N_A_29_65#_c_789_n 0.00277403f $X=2.675 $Y=1.275 $X2=0 $Y2=0
cc_206 N_B1_c_163_n N_A_29_65#_c_790_n 0.00917604f $X=2.675 $Y=1.275 $X2=0 $Y2=0
cc_207 B1 N_A_29_65#_c_790_n 0.00390375f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_208 N_B1_c_170_n N_A_29_65#_c_790_n 0.0138088f $X=1.365 $Y=1.275 $X2=0 $Y2=0
cc_209 N_B1_c_171_n N_A_284_65#_M1015_s 0.00219477f $X=1.82 $Y=1.34 $X2=-0.19
+ $Y2=-0.245
cc_210 N_B1_c_165_n N_A_284_65#_M1020_d 0.00176891f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_211 B1 N_A_284_65#_c_828_n 0.00738292f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_212 N_B1_c_169_n N_A_284_65#_c_828_n 4.15557e-19 $X=1.365 $Y=1.44 $X2=0 $Y2=0
cc_213 N_B1_c_171_n N_A_284_65#_c_828_n 0.0348267f $X=1.82 $Y=1.34 $X2=0 $Y2=0
cc_214 N_B1_c_163_n N_A_284_65#_c_823_n 2.62132e-19 $X=2.675 $Y=1.275 $X2=0
+ $Y2=0
cc_215 N_B1_c_163_n N_A_284_65#_c_832_n 0.00222917f $X=2.675 $Y=1.275 $X2=0
+ $Y2=0
cc_216 N_B1_c_165_n N_A_284_65#_c_832_n 0.0348267f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B1_c_163_n N_A_284_65#_c_825_n 0.00892373f $X=2.675 $Y=1.275 $X2=0
+ $Y2=0
cc_218 N_B1_c_165_n N_A_284_65#_c_825_n 0.0204095f $X=2.905 $Y=1.16 $X2=0 $Y2=0
cc_219 N_B1_c_167_n N_A_284_65#_c_825_n 0.00126308f $X=2.99 $Y=1.44 $X2=0 $Y2=0
cc_220 N_B1_c_163_n N_VGND_c_867_n 0.00168875f $X=2.675 $Y=1.275 $X2=0 $Y2=0
cc_221 N_B1_c_163_n N_VGND_c_874_n 0.00302501f $X=2.675 $Y=1.275 $X2=0 $Y2=0
cc_222 N_B1_c_170_n N_VGND_c_874_n 0.00302501f $X=1.365 $Y=1.275 $X2=0 $Y2=0
cc_223 N_B1_c_163_n N_VGND_c_882_n 0.00485634f $X=2.675 $Y=1.275 $X2=0 $Y2=0
cc_224 N_B1_c_170_n N_VGND_c_882_n 0.00440224f $X=1.365 $Y=1.275 $X2=0 $Y2=0
cc_225 N_B2_M1009_g N_A_112_65#_c_461_n 0.0129102f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_226 N_B2_M1018_g N_A_112_65#_c_472_n 0.0111034f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_227 B2 N_A_112_65#_c_472_n 0.0362688f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B2_M1009_g N_A_112_65#_c_475_n 0.0110689f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_229 N_B2_M1018_g N_A_112_65#_c_475_n 0.0101708f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_230 B2 N_A_112_65#_c_475_n 0.0150188f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_231 N_B2_c_253_n N_A_112_65#_c_475_n 9.79786e-19 $X=2.245 $Y=1.51 $X2=0 $Y2=0
cc_232 N_B2_M1009_g N_VPWR_c_596_n 0.00105138f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_233 N_B2_M1018_g N_VPWR_c_597_n 0.00115783f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_234 N_B2_M1009_g N_VPWR_c_603_n 0.00357877f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_235 N_B2_M1018_g N_VPWR_c_603_n 0.00357877f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_236 N_B2_M1009_g N_VPWR_c_593_n 0.00537654f $X=1.815 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B2_M1018_g N_VPWR_c_593_n 0.00537654f $X=2.245 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B2_M1009_g N_A_292_367#_c_694_n 0.0114565f $X=1.815 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_B2_M1018_g N_A_292_367#_c_694_n 0.0114565f $X=2.245 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_B2_M1003_g N_A_29_65#_c_790_n 0.0115051f $X=1.815 $Y=0.745 $X2=0 $Y2=0
cc_241 N_B2_M1020_g N_A_29_65#_c_790_n 0.011126f $X=2.245 $Y=0.745 $X2=0 $Y2=0
cc_242 N_B2_M1003_g N_A_284_65#_c_828_n 0.00910195f $X=1.815 $Y=0.745 $X2=0
+ $Y2=0
cc_243 N_B2_M1020_g N_A_284_65#_c_828_n 0.00910195f $X=2.245 $Y=0.745 $X2=0
+ $Y2=0
cc_244 N_B2_M1003_g N_VGND_c_874_n 0.00302501f $X=1.815 $Y=0.745 $X2=0 $Y2=0
cc_245 N_B2_M1020_g N_VGND_c_874_n 0.00302501f $X=2.245 $Y=0.745 $X2=0 $Y2=0
cc_246 N_B2_M1003_g N_VGND_c_882_n 0.0043925f $X=1.815 $Y=0.745 $X2=0 $Y2=0
cc_247 N_B2_M1020_g N_VGND_c_882_n 0.00435646f $X=2.245 $Y=0.745 $X2=0 $Y2=0
cc_248 N_A1_c_302_n N_A2_M1010_g 7.23929e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A1_c_304_n N_A2_M1010_g 0.0387407f $X=3.535 $Y=1.185 $X2=0 $Y2=0
cc_250 N_A1_c_306_n N_A2_M1010_g 5.49816e-19 $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_251 N_A1_c_308_n N_A2_M1010_g 0.0105012f $X=4.465 $Y=1.295 $X2=0 $Y2=0
cc_252 N_A1_M1011_g N_A2_M1027_g 0.0229039f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_253 N_A1_c_305_n N_A2_M1017_g 0.0200703f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_254 N_A1_c_306_n N_A2_M1017_g 0.00800574f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_255 N_A1_c_307_n N_A2_M1017_g 0.0311483f $X=4.935 $Y=1.185 $X2=0 $Y2=0
cc_256 N_A1_c_308_n N_A2_M1017_g 0.00598841f $X=4.465 $Y=1.295 $X2=0 $Y2=0
cc_257 N_A1_M1007_g N_A2_c_387_n 0.00567357f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A1_c_302_n N_A2_c_387_n 0.00726628f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A1_c_303_n N_A2_c_387_n 5.99261e-19 $X=3.535 $Y=1.35 $X2=0 $Y2=0
cc_260 N_A1_c_305_n N_A2_c_387_n 7.35159e-19 $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_261 N_A1_c_306_n N_A2_c_387_n 0.00714502f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_262 N_A1_c_308_n N_A2_c_387_n 0.0312207f $X=4.465 $Y=1.295 $X2=0 $Y2=0
cc_263 N_A1_M1007_g N_A2_c_388_n 0.0421804f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A1_c_302_n N_A2_c_388_n 6.65848e-19 $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A1_c_303_n N_A2_c_388_n 0.00859299f $X=3.535 $Y=1.35 $X2=0 $Y2=0
cc_266 N_A1_c_305_n N_A2_c_388_n 0.0229039f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_267 N_A1_c_306_n N_A2_c_388_n 0.00966833f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_268 N_A1_c_308_n N_A2_c_388_n 0.00388788f $X=4.465 $Y=1.295 $X2=0 $Y2=0
cc_269 N_A1_c_305_n N_A_112_65#_M1004_g 0.0188454f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_270 N_A1_c_306_n N_A_112_65#_M1004_g 0.00205108f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_271 N_A1_c_307_n N_A_112_65#_M1004_g 0.0150513f $X=4.935 $Y=1.185 $X2=0 $Y2=0
cc_272 N_A1_M1007_g N_A_112_65#_c_472_n 0.0176274f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A1_c_302_n N_A_112_65#_c_472_n 0.0095814f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_274 N_A1_c_303_n N_A_112_65#_c_472_n 9.64415e-19 $X=3.535 $Y=1.35 $X2=0 $Y2=0
cc_275 N_A1_M1011_g N_A_112_65#_c_490_n 0.01627f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A1_c_305_n N_A_112_65#_c_490_n 0.00412461f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_277 N_A1_c_306_n N_A_112_65#_c_490_n 0.0190191f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_278 N_A1_M1011_g N_A_112_65#_c_443_n 0.00663693f $X=4.845 $Y=2.465 $X2=0
+ $Y2=0
cc_279 N_A1_M1011_g N_A_112_65#_c_444_n 0.00177586f $X=4.845 $Y=2.465 $X2=0
+ $Y2=0
cc_280 N_A1_c_305_n N_A_112_65#_c_444_n 9.60004e-19 $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_281 N_A1_c_306_n N_A_112_65#_c_444_n 0.0113481f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_282 N_A1_M1007_g N_A_112_65#_c_497_n 8.92984e-19 $X=3.555 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_A1_M1011_g N_A_112_65#_c_497_n 9.54555e-19 $X=4.845 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_A1_M1011_g N_A_112_65#_c_445_n 0.0385082f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_285 N_A1_c_305_n N_A_112_65#_c_445_n 0.00203966f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_286 N_A1_M1007_g N_VPWR_c_597_n 0.0194393f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A1_M1011_g N_VPWR_c_598_n 0.00814344f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_288 N_A1_M1007_g N_VPWR_c_604_n 0.00486043f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_289 N_A1_M1011_g N_VPWR_c_604_n 0.00547432f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_290 N_A1_M1007_g N_VPWR_c_593_n 0.0082726f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A1_M1011_g N_VPWR_c_593_n 0.0102357f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A1_M1011_g N_A_726_367#_c_708_n 0.00198785f $X=4.845 $Y=2.465 $X2=0
+ $Y2=0
cc_293 N_A1_M1011_g N_A_726_367#_c_709_n 0.00755845f $X=4.845 $Y=2.465 $X2=0
+ $Y2=0
cc_294 N_A1_c_306_n N_X_c_725_n 0.00659735f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_295 N_A1_c_302_n N_A_284_65#_c_824_n 0.0223882f $X=3.53 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A1_c_303_n N_A_284_65#_c_824_n 8.54053e-19 $X=3.535 $Y=1.35 $X2=0 $Y2=0
cc_297 N_A1_c_304_n N_A_284_65#_c_824_n 0.012775f $X=3.535 $Y=1.185 $X2=0 $Y2=0
cc_298 N_A1_c_305_n N_A_284_65#_c_824_n 2.68039e-19 $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_299 N_A1_c_307_n N_A_284_65#_c_824_n 0.00290087f $X=4.935 $Y=1.185 $X2=0
+ $Y2=0
cc_300 N_A1_c_308_n N_A_284_65#_c_824_n 0.0751366f $X=4.465 $Y=1.295 $X2=0 $Y2=0
cc_301 N_A1_c_302_n N_VGND_M1002_s 0.00195953f $X=3.53 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_302 N_A1_c_304_n N_VGND_c_867_n 0.0103512f $X=3.535 $Y=1.185 $X2=0 $Y2=0
cc_303 N_A1_c_304_n N_VGND_c_868_n 0.0013251f $X=3.535 $Y=1.185 $X2=0 $Y2=0
cc_304 N_A1_c_307_n N_VGND_c_868_n 0.00137734f $X=4.935 $Y=1.185 $X2=0 $Y2=0
cc_305 N_A1_c_307_n N_VGND_c_869_n 0.00560454f $X=4.935 $Y=1.185 $X2=0 $Y2=0
cc_306 N_A1_c_305_n N_VGND_c_870_n 0.00229172f $X=4.935 $Y=1.35 $X2=0 $Y2=0
cc_307 N_A1_c_307_n N_VGND_c_870_n 0.0015486f $X=4.935 $Y=1.185 $X2=0 $Y2=0
cc_308 N_A1_c_304_n N_VGND_c_876_n 0.00362386f $X=3.535 $Y=1.185 $X2=0 $Y2=0
cc_309 N_A1_c_304_n N_VGND_c_882_n 0.00437379f $X=3.535 $Y=1.185 $X2=0 $Y2=0
cc_310 N_A1_c_307_n N_VGND_c_882_n 0.0100768f $X=4.935 $Y=1.185 $X2=0 $Y2=0
cc_311 N_A2_M1016_g N_A_112_65#_c_472_n 0.0110983f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_312 N_A2_c_387_n N_A_112_65#_c_472_n 0.0110052f $X=4.13 $Y=1.51 $X2=0 $Y2=0
cc_313 N_A2_M1027_g N_A_112_65#_c_490_n 0.0143434f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A2_c_388_n N_A_112_65#_c_490_n 2.1507e-19 $X=4.415 $Y=1.51 $X2=0 $Y2=0
cc_315 N_A2_M1016_g N_A_112_65#_c_497_n 0.0102902f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_316 N_A2_M1027_g N_A_112_65#_c_497_n 0.0112745f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_317 N_A2_c_387_n N_A_112_65#_c_497_n 0.0193049f $X=4.13 $Y=1.51 $X2=0 $Y2=0
cc_318 N_A2_c_388_n N_A_112_65#_c_497_n 6.31337e-19 $X=4.415 $Y=1.51 $X2=0 $Y2=0
cc_319 N_A2_M1016_g N_VPWR_c_597_n 0.00115783f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_320 N_A2_M1016_g N_VPWR_c_604_n 0.00357877f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_321 N_A2_M1027_g N_VPWR_c_604_n 0.00357877f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A2_M1016_g N_VPWR_c_593_n 0.00537654f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_323 N_A2_M1027_g N_VPWR_c_593_n 0.00537654f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_324 N_A2_M1016_g N_A_726_367#_c_708_n 0.0115031f $X=3.985 $Y=2.465 $X2=0
+ $Y2=0
cc_325 N_A2_M1027_g N_A_726_367#_c_708_n 0.0114565f $X=4.415 $Y=2.465 $X2=0
+ $Y2=0
cc_326 N_A2_M1010_g N_A_284_65#_c_824_n 0.0104843f $X=4.055 $Y=0.655 $X2=0 $Y2=0
cc_327 N_A2_M1017_g N_A_284_65#_c_824_n 0.0104843f $X=4.485 $Y=0.655 $X2=0 $Y2=0
cc_328 N_A2_M1010_g N_VGND_c_867_n 0.0013251f $X=4.055 $Y=0.655 $X2=0 $Y2=0
cc_329 N_A2_M1010_g N_VGND_c_868_n 0.00928769f $X=4.055 $Y=0.655 $X2=0 $Y2=0
cc_330 N_A2_M1017_g N_VGND_c_868_n 0.00975952f $X=4.485 $Y=0.655 $X2=0 $Y2=0
cc_331 N_A2_M1017_g N_VGND_c_869_n 0.00362386f $X=4.485 $Y=0.655 $X2=0 $Y2=0
cc_332 N_A2_M1010_g N_VGND_c_876_n 0.00362386f $X=4.055 $Y=0.655 $X2=0 $Y2=0
cc_333 N_A2_M1010_g N_VGND_c_882_n 0.00437379f $X=4.055 $Y=0.655 $X2=0 $Y2=0
cc_334 N_A2_M1017_g N_VGND_c_882_n 0.00437379f $X=4.485 $Y=0.655 $X2=0 $Y2=0
cc_335 N_A_112_65#_c_461_n N_VPWR_M1022_d 0.00501123f $X=1.865 $Y=2.015 $X2=0
+ $Y2=0
cc_336 N_A_112_65#_c_472_n N_VPWR_M1026_s 0.0231566f $X=4.035 $Y=2.015 $X2=0
+ $Y2=0
cc_337 N_A_112_65#_c_490_n N_VPWR_M1011_d 0.00942156f $X=5.2 $Y=2.015 $X2=0
+ $Y2=0
cc_338 N_A_112_65#_c_443_n N_VPWR_M1011_d 0.00118786f $X=5.285 $Y=1.93 $X2=0
+ $Y2=0
cc_339 N_A_112_65#_c_461_n N_VPWR_c_596_n 0.017285f $X=1.865 $Y=2.015 $X2=0
+ $Y2=0
cc_340 N_A_112_65#_c_472_n N_VPWR_c_597_n 0.053689f $X=4.035 $Y=2.015 $X2=0
+ $Y2=0
cc_341 N_A_112_65#_M1001_g N_VPWR_c_598_n 0.00677703f $X=5.42 $Y=2.465 $X2=0
+ $Y2=0
cc_342 N_A_112_65#_c_490_n N_VPWR_c_598_n 0.0260249f $X=5.2 $Y=2.015 $X2=0 $Y2=0
cc_343 N_A_112_65#_M1001_g N_VPWR_c_599_n 7.52465e-19 $X=5.42 $Y=2.465 $X2=0
+ $Y2=0
cc_344 N_A_112_65#_M1013_g N_VPWR_c_599_n 0.0144667f $X=5.85 $Y=2.465 $X2=0
+ $Y2=0
cc_345 N_A_112_65#_M1019_g N_VPWR_c_599_n 0.0143085f $X=6.28 $Y=2.465 $X2=0
+ $Y2=0
cc_346 N_A_112_65#_M1025_g N_VPWR_c_599_n 7.24342e-19 $X=6.71 $Y=2.465 $X2=0
+ $Y2=0
cc_347 N_A_112_65#_M1019_g N_VPWR_c_601_n 7.24342e-19 $X=6.28 $Y=2.465 $X2=0
+ $Y2=0
cc_348 N_A_112_65#_M1025_g N_VPWR_c_601_n 0.0154956f $X=6.71 $Y=2.465 $X2=0
+ $Y2=0
cc_349 N_A_112_65#_c_523_p N_VPWR_c_602_n 0.0131621f $X=0.7 $Y=2.475 $X2=0 $Y2=0
cc_350 N_A_112_65#_M1001_g N_VPWR_c_605_n 0.00585385f $X=5.42 $Y=2.465 $X2=0
+ $Y2=0
cc_351 N_A_112_65#_M1013_g N_VPWR_c_605_n 0.00486043f $X=5.85 $Y=2.465 $X2=0
+ $Y2=0
cc_352 N_A_112_65#_M1019_g N_VPWR_c_606_n 0.00486043f $X=6.28 $Y=2.465 $X2=0
+ $Y2=0
cc_353 N_A_112_65#_M1025_g N_VPWR_c_606_n 0.00486043f $X=6.71 $Y=2.465 $X2=0
+ $Y2=0
cc_354 N_A_112_65#_M1006_s N_VPWR_c_593_n 0.00467071f $X=0.56 $Y=1.835 $X2=0
+ $Y2=0
cc_355 N_A_112_65#_M1009_s N_VPWR_c_593_n 0.00225186f $X=1.89 $Y=1.835 $X2=0
+ $Y2=0
cc_356 N_A_112_65#_M1016_s N_VPWR_c_593_n 0.00225186f $X=4.06 $Y=1.835 $X2=0
+ $Y2=0
cc_357 N_A_112_65#_M1001_g N_VPWR_c_593_n 0.0110861f $X=5.42 $Y=2.465 $X2=0
+ $Y2=0
cc_358 N_A_112_65#_M1013_g N_VPWR_c_593_n 0.00824727f $X=5.85 $Y=2.465 $X2=0
+ $Y2=0
cc_359 N_A_112_65#_M1019_g N_VPWR_c_593_n 0.00824727f $X=6.28 $Y=2.465 $X2=0
+ $Y2=0
cc_360 N_A_112_65#_M1025_g N_VPWR_c_593_n 0.00824727f $X=6.71 $Y=2.465 $X2=0
+ $Y2=0
cc_361 N_A_112_65#_c_523_p N_VPWR_c_593_n 0.00808656f $X=0.7 $Y=2.475 $X2=0
+ $Y2=0
cc_362 N_A_112_65#_c_461_n N_A_292_367#_M1000_d 0.00412021f $X=1.865 $Y=2.015
+ $X2=-0.19 $Y2=-0.245
cc_363 N_A_112_65#_c_472_n N_A_292_367#_M1018_d 0.00353353f $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_364 N_A_112_65#_c_461_n N_A_292_367#_c_698_n 0.0135055f $X=1.865 $Y=2.015
+ $X2=0 $Y2=0
cc_365 N_A_112_65#_M1009_s N_A_292_367#_c_694_n 0.00332344f $X=1.89 $Y=1.835
+ $X2=0 $Y2=0
cc_366 N_A_112_65#_c_475_n N_A_292_367#_c_694_n 0.0159805f $X=2.03 $Y=2.095
+ $X2=0 $Y2=0
cc_367 N_A_112_65#_c_472_n N_A_292_367#_c_701_n 0.0135055f $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_368 N_A_112_65#_c_472_n N_A_726_367#_M1007_s 0.00775942f $X=4.035 $Y=2.015
+ $X2=-0.19 $Y2=-0.245
cc_369 N_A_112_65#_c_490_n N_A_726_367#_M1027_d 0.00448746f $X=5.2 $Y=2.015
+ $X2=0 $Y2=0
cc_370 N_A_112_65#_c_472_n N_A_726_367#_c_714_n 0.0135055f $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_371 N_A_112_65#_M1016_s N_A_726_367#_c_708_n 0.00332344f $X=4.06 $Y=1.835
+ $X2=0 $Y2=0
cc_372 N_A_112_65#_c_497_n N_A_726_367#_c_708_n 0.0159805f $X=4.2 $Y=2.095 $X2=0
+ $Y2=0
cc_373 N_A_112_65#_c_490_n N_A_726_367#_c_709_n 0.0146459f $X=5.2 $Y=2.015 $X2=0
+ $Y2=0
cc_374 N_A_112_65#_M1012_g N_X_c_724_n 0.0136745f $X=5.815 $Y=0.655 $X2=0 $Y2=0
cc_375 N_A_112_65#_M1021_g N_X_c_724_n 0.0138978f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_376 N_A_112_65#_c_550_p N_X_c_724_n 0.0473015f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_377 N_A_112_65#_c_445_n N_X_c_724_n 0.00255374f $X=6.675 $Y=1.49 $X2=0 $Y2=0
cc_378 N_A_112_65#_M1004_g N_X_c_725_n 0.00200648f $X=5.385 $Y=0.655 $X2=0 $Y2=0
cc_379 N_A_112_65#_c_550_p N_X_c_725_n 0.0187574f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_380 N_A_112_65#_c_445_n N_X_c_725_n 0.00265263f $X=6.675 $Y=1.49 $X2=0 $Y2=0
cc_381 N_A_112_65#_M1013_g N_X_c_730_n 0.0130133f $X=5.85 $Y=2.465 $X2=0 $Y2=0
cc_382 N_A_112_65#_M1019_g N_X_c_730_n 0.0131755f $X=6.28 $Y=2.465 $X2=0 $Y2=0
cc_383 N_A_112_65#_c_550_p N_X_c_730_n 0.0473014f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_384 N_A_112_65#_c_445_n N_X_c_730_n 0.00258422f $X=6.675 $Y=1.49 $X2=0 $Y2=0
cc_385 N_A_112_65#_M1001_g N_X_c_731_n 6.55961e-19 $X=5.42 $Y=2.465 $X2=0 $Y2=0
cc_386 N_A_112_65#_c_443_n N_X_c_731_n 0.00947164f $X=5.285 $Y=1.93 $X2=0 $Y2=0
cc_387 N_A_112_65#_c_550_p N_X_c_731_n 0.0154947f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_388 N_A_112_65#_c_445_n N_X_c_731_n 0.00268515f $X=6.675 $Y=1.49 $X2=0 $Y2=0
cc_389 N_A_112_65#_M1024_g N_X_c_726_n 0.0160926f $X=6.675 $Y=0.655 $X2=0 $Y2=0
cc_390 N_A_112_65#_c_550_p N_X_c_726_n 0.00974094f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_391 N_A_112_65#_c_445_n N_X_c_726_n 0.00113866f $X=6.675 $Y=1.49 $X2=0 $Y2=0
cc_392 N_A_112_65#_M1025_g N_X_c_732_n 0.0156161f $X=6.71 $Y=2.465 $X2=0 $Y2=0
cc_393 N_A_112_65#_c_550_p N_X_c_732_n 0.00733859f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_394 N_A_112_65#_c_550_p N_X_c_727_n 0.0154948f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_395 N_A_112_65#_c_445_n N_X_c_727_n 0.00265263f $X=6.675 $Y=1.49 $X2=0 $Y2=0
cc_396 N_A_112_65#_c_550_p N_X_c_733_n 0.0154947f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_397 N_A_112_65#_c_445_n N_X_c_733_n 0.00268515f $X=6.675 $Y=1.49 $X2=0 $Y2=0
cc_398 N_A_112_65#_M1024_g X 0.00414777f $X=6.675 $Y=0.655 $X2=0 $Y2=0
cc_399 N_A_112_65#_c_550_p X 0.0162728f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_400 N_A_112_65#_c_445_n X 0.0160363f $X=6.675 $Y=1.49 $X2=0 $Y2=0
cc_401 N_A_112_65#_M1005_d N_A_29_65#_c_786_n 0.00176461f $X=0.56 $Y=0.325 $X2=0
+ $Y2=0
cc_402 N_A_112_65#_c_453_n N_A_29_65#_c_786_n 0.0159533f $X=0.7 $Y=0.68 $X2=0
+ $Y2=0
cc_403 N_A_112_65#_M1004_g N_VGND_c_870_n 0.00163601f $X=5.385 $Y=0.655 $X2=0
+ $Y2=0
cc_404 N_A_112_65#_c_444_n N_VGND_c_870_n 0.00325583f $X=5.37 $Y=1.485 $X2=0
+ $Y2=0
cc_405 N_A_112_65#_M1004_g N_VGND_c_871_n 6.3872e-19 $X=5.385 $Y=0.655 $X2=0
+ $Y2=0
cc_406 N_A_112_65#_M1012_g N_VGND_c_871_n 0.0108228f $X=5.815 $Y=0.655 $X2=0
+ $Y2=0
cc_407 N_A_112_65#_M1021_g N_VGND_c_871_n 0.0107309f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_408 N_A_112_65#_M1024_g N_VGND_c_871_n 6.22495e-19 $X=6.675 $Y=0.655 $X2=0
+ $Y2=0
cc_409 N_A_112_65#_M1021_g N_VGND_c_873_n 6.25324e-19 $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_410 N_A_112_65#_M1024_g N_VGND_c_873_n 0.0120503f $X=6.675 $Y=0.655 $X2=0
+ $Y2=0
cc_411 N_A_112_65#_M1004_g N_VGND_c_878_n 0.00585385f $X=5.385 $Y=0.655 $X2=0
+ $Y2=0
cc_412 N_A_112_65#_M1012_g N_VGND_c_878_n 0.00486043f $X=5.815 $Y=0.655 $X2=0
+ $Y2=0
cc_413 N_A_112_65#_M1021_g N_VGND_c_879_n 0.00486043f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_414 N_A_112_65#_M1024_g N_VGND_c_879_n 0.00486043f $X=6.675 $Y=0.655 $X2=0
+ $Y2=0
cc_415 N_A_112_65#_M1004_g N_VGND_c_882_n 0.0106551f $X=5.385 $Y=0.655 $X2=0
+ $Y2=0
cc_416 N_A_112_65#_M1012_g N_VGND_c_882_n 0.00824727f $X=5.815 $Y=0.655 $X2=0
+ $Y2=0
cc_417 N_A_112_65#_M1021_g N_VGND_c_882_n 0.00824727f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_418 N_A_112_65#_M1024_g N_VGND_c_882_n 0.00824727f $X=6.675 $Y=0.655 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_593_n N_A_292_367#_M1000_d 0.00307052f $X=6.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_420 N_VPWR_c_593_n N_A_292_367#_M1018_d 0.00376627f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_603_n N_A_292_367#_c_694_n 0.0486406f $X=2.725 $Y=3.33 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_593_n N_A_292_367#_c_694_n 0.0310628f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_603_n N_A_292_367#_c_706_n 0.0132331f $X=2.725 $Y=3.33 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_593_n N_A_292_367#_c_706_n 0.00816431f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_593_n N_A_726_367#_M1007_s 0.00376627f $X=6.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_426 N_VPWR_c_593_n N_A_726_367#_M1027_d 0.00223562f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_604_n N_A_726_367#_c_708_n 0.0519089f $X=4.97 $Y=3.33 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_593_n N_A_726_367#_c_708_n 0.0335966f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_604_n N_A_726_367#_c_722_n 0.0125234f $X=4.97 $Y=3.33 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_593_n N_A_726_367#_c_722_n 0.00738676f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_593_n N_X_M1001_d 0.00536646f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_432 N_VPWR_c_593_n N_X_M1019_d 0.00536646f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_433 N_VPWR_c_605_n N_X_c_765_n 0.0124525f $X=5.9 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_c_593_n N_X_c_765_n 0.00730901f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_435 N_VPWR_M1013_s N_X_c_730_n 0.00180746f $X=5.925 $Y=1.835 $X2=0 $Y2=0
cc_436 N_VPWR_c_599_n N_X_c_730_n 0.0163515f $X=6.065 $Y=2.19 $X2=0 $Y2=0
cc_437 N_VPWR_c_606_n N_X_c_769_n 0.0124525f $X=6.76 $Y=3.33 $X2=0 $Y2=0
cc_438 N_VPWR_c_593_n N_X_c_769_n 0.00730901f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_439 N_VPWR_M1025_s N_X_c_732_n 0.00276041f $X=6.785 $Y=1.835 $X2=0 $Y2=0
cc_440 N_VPWR_c_601_n N_X_c_732_n 0.0229493f $X=6.925 $Y=2.19 $X2=0 $Y2=0
cc_441 N_X_c_724_n N_VGND_M1012_d 0.00180746f $X=6.365 $Y=1.13 $X2=0 $Y2=0
cc_442 N_X_c_726_n N_VGND_M1024_d 6.05921e-19 $X=6.865 $Y=1.13 $X2=0 $Y2=0
cc_443 N_X_c_728_n N_VGND_M1024_d 0.00205561f $X=6.99 $Y=1.215 $X2=0 $Y2=0
cc_444 N_X_c_724_n N_VGND_c_871_n 0.0163515f $X=6.365 $Y=1.13 $X2=0 $Y2=0
cc_445 N_X_c_726_n N_VGND_c_873_n 0.0064684f $X=6.865 $Y=1.13 $X2=0 $Y2=0
cc_446 N_X_c_728_n N_VGND_c_873_n 0.0171078f $X=6.99 $Y=1.215 $X2=0 $Y2=0
cc_447 N_X_c_779_p N_VGND_c_878_n 0.0138717f $X=5.6 $Y=0.42 $X2=0 $Y2=0
cc_448 N_X_c_780_p N_VGND_c_879_n 0.0124525f $X=6.46 $Y=0.42 $X2=0 $Y2=0
cc_449 N_X_M1004_s N_VGND_c_882_n 0.00397496f $X=5.46 $Y=0.235 $X2=0 $Y2=0
cc_450 N_X_M1021_s N_VGND_c_882_n 0.00536646f $X=6.32 $Y=0.235 $X2=0 $Y2=0
cc_451 N_X_c_779_p N_VGND_c_882_n 0.00886411f $X=5.6 $Y=0.42 $X2=0 $Y2=0
cc_452 N_X_c_780_p N_VGND_c_882_n 0.00730901f $X=6.46 $Y=0.42 $X2=0 $Y2=0
cc_453 N_A_29_65#_c_790_n N_A_284_65#_M1015_s 0.00223038f $X=2.725 $Y=0.405
+ $X2=-0.19 $Y2=-0.245
cc_454 N_A_29_65#_c_790_n N_A_284_65#_M1020_d 0.00179729f $X=2.725 $Y=0.405
+ $X2=0 $Y2=0
cc_455 N_A_29_65#_M1003_s N_A_284_65#_c_828_n 0.00336695f $X=1.89 $Y=0.325 $X2=0
+ $Y2=0
cc_456 N_A_29_65#_c_790_n N_A_284_65#_c_828_n 0.0629266f $X=2.725 $Y=0.405 $X2=0
+ $Y2=0
cc_457 N_A_29_65#_M1023_d N_A_284_65#_c_825_n 0.00487561f $X=2.75 $Y=0.325 $X2=0
+ $Y2=0
cc_458 N_A_29_65#_c_789_n N_A_284_65#_c_825_n 0.0199859f $X=2.89 $Y=0.47 $X2=0
+ $Y2=0
cc_459 N_A_29_65#_c_790_n N_A_284_65#_c_825_n 0.00499648f $X=2.725 $Y=0.405
+ $X2=0 $Y2=0
cc_460 N_A_29_65#_c_789_n N_VGND_c_867_n 0.0232212f $X=2.89 $Y=0.47 $X2=0 $Y2=0
cc_461 N_A_29_65#_c_786_n N_VGND_c_874_n 0.0422287f $X=1.035 $Y=0.34 $X2=0 $Y2=0
cc_462 N_A_29_65#_c_787_n N_VGND_c_874_n 0.0186386f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_463 N_A_29_65#_c_788_n N_VGND_c_874_n 0.0165592f $X=1.13 $Y=0.47 $X2=0 $Y2=0
cc_464 N_A_29_65#_c_790_n N_VGND_c_874_n 0.117712f $X=2.725 $Y=0.405 $X2=0 $Y2=0
cc_465 N_A_29_65#_c_786_n N_VGND_c_882_n 0.0238173f $X=1.035 $Y=0.34 $X2=0 $Y2=0
cc_466 N_A_29_65#_c_787_n N_VGND_c_882_n 0.0101082f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_467 N_A_29_65#_c_788_n N_VGND_c_882_n 0.00895533f $X=1.13 $Y=0.47 $X2=0 $Y2=0
cc_468 N_A_29_65#_c_790_n N_VGND_c_882_n 0.0653393f $X=2.725 $Y=0.405 $X2=0
+ $Y2=0
cc_469 N_A_284_65#_c_824_n N_VGND_M1002_s 0.00747177f $X=4.7 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_470 N_A_284_65#_c_824_n N_VGND_M1010_d 0.00336289f $X=4.7 $Y=0.805 $X2=0
+ $Y2=0
cc_471 N_A_284_65#_c_824_n N_VGND_c_867_n 0.0212603f $X=4.7 $Y=0.805 $X2=0 $Y2=0
cc_472 N_A_284_65#_c_824_n N_VGND_c_868_n 0.0165006f $X=4.7 $Y=0.805 $X2=0 $Y2=0
cc_473 N_A_284_65#_c_824_n N_VGND_c_869_n 0.00548336f $X=4.7 $Y=0.805 $X2=0
+ $Y2=0
cc_474 N_A_284_65#_c_823_n N_VGND_c_874_n 0.00172364f $X=3.232 $Y=0.807 $X2=0
+ $Y2=0
cc_475 N_A_284_65#_c_825_n N_VGND_c_874_n 0.00121409f $X=3.135 $Y=0.807 $X2=0
+ $Y2=0
cc_476 N_A_284_65#_c_824_n N_VGND_c_876_n 0.00686768f $X=4.7 $Y=0.805 $X2=0
+ $Y2=0
cc_477 N_A_284_65#_M1002_d N_VGND_c_882_n 0.00356404f $X=3.7 $Y=0.235 $X2=0
+ $Y2=0
cc_478 N_A_284_65#_M1017_s N_VGND_c_882_n 0.00356404f $X=4.56 $Y=0.235 $X2=0
+ $Y2=0
cc_479 N_A_284_65#_c_823_n N_VGND_c_882_n 0.0030156f $X=3.232 $Y=0.807 $X2=0
+ $Y2=0
cc_480 N_A_284_65#_c_824_n N_VGND_c_882_n 0.0266556f $X=4.7 $Y=0.805 $X2=0 $Y2=0
cc_481 N_A_284_65#_c_825_n N_VGND_c_882_n 0.00280399f $X=3.135 $Y=0.807 $X2=0
+ $Y2=0
