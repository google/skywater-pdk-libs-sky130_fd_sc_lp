* NGSPICE file created from sky130_fd_sc_lp__nand2_lp2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand2_lp2 A B VGND VNB VPB VPWR Y
M1000 Y A a_151_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1001 a_151_57# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1002 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=5.7e+11p pd=5.14e+06u as=2.8e+11p ps=2.56e+06u
M1003 Y B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

