* File: sky130_fd_sc_lp__a2111oi_1.pxi.spice
* Created: Fri Aug 28 09:46:33 2020
* 
x_PM_SKY130_FD_SC_LP__A2111OI_1%D1 N_D1_M1002_g N_D1_M1005_g D1 D1 D1 D1
+ N_D1_c_50_n N_D1_c_51_n PM_SKY130_FD_SC_LP__A2111OI_1%D1
x_PM_SKY130_FD_SC_LP__A2111OI_1%C1 N_C1_M1008_g N_C1_M1000_g C1 C1 C1 C1 C1
+ N_C1_c_84_n PM_SKY130_FD_SC_LP__A2111OI_1%C1
x_PM_SKY130_FD_SC_LP__A2111OI_1%B1 N_B1_M1004_g N_B1_c_120_n N_B1_M1009_g B1
+ N_B1_c_122_n PM_SKY130_FD_SC_LP__A2111OI_1%B1
x_PM_SKY130_FD_SC_LP__A2111OI_1%A1 N_A1_M1001_g N_A1_c_152_n N_A1_M1006_g A1 A1
+ N_A1_c_154_n PM_SKY130_FD_SC_LP__A2111OI_1%A1
x_PM_SKY130_FD_SC_LP__A2111OI_1%A2 N_A2_c_183_n N_A2_M1003_g N_A2_M1007_g A2
+ N_A2_c_186_n PM_SKY130_FD_SC_LP__A2111OI_1%A2
x_PM_SKY130_FD_SC_LP__A2111OI_1%Y N_Y_M1002_d N_Y_M1009_d N_Y_M1005_s
+ N_Y_c_207_n N_Y_c_208_n Y Y Y Y Y N_Y_c_241_p N_Y_c_210_n N_Y_c_223_n
+ PM_SKY130_FD_SC_LP__A2111OI_1%Y
x_PM_SKY130_FD_SC_LP__A2111OI_1%A_343_367# N_A_343_367#_M1004_d
+ N_A_343_367#_M1007_d N_A_343_367#_c_270_p N_A_343_367#_c_254_n
+ N_A_343_367#_c_255_n N_A_343_367#_c_256_n
+ PM_SKY130_FD_SC_LP__A2111OI_1%A_343_367#
x_PM_SKY130_FD_SC_LP__A2111OI_1%VPWR N_VPWR_M1001_d N_VPWR_c_277_n
+ N_VPWR_c_278_n N_VPWR_c_279_n VPWR N_VPWR_c_280_n N_VPWR_c_276_n
+ PM_SKY130_FD_SC_LP__A2111OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A2111OI_1%VGND N_VGND_M1002_s N_VGND_M1008_d
+ N_VGND_M1003_d N_VGND_c_311_n N_VGND_c_312_n N_VGND_c_313_n N_VGND_c_314_n
+ N_VGND_c_315_n VGND N_VGND_c_316_n N_VGND_c_317_n
+ PM_SKY130_FD_SC_LP__A2111OI_1%VGND
cc_1 VNB N_D1_M1002_g 0.0293967f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_2 VNB N_D1_c_50_n 0.0043755f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_3 VNB N_D1_c_51_n 0.0272592f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.51
cc_4 VNB N_C1_M1008_g 0.0214429f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_5 VNB N_C1_M1000_g 0.00517185f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.465
cc_6 VNB C1 0.00364013f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_7 VNB N_C1_c_84_n 0.0381186f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_8 VNB N_B1_M1004_g 0.00793252f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_9 VNB N_B1_c_120_n 0.0201258f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.675
cc_10 VNB B1 0.0108019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_c_122_n 0.0335266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_M1001_g 0.00880642f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.655
cc_13 VNB N_A1_c_152_n 0.0171567f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.675
cc_14 VNB A1 0.00792292f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_15 VNB N_A1_c_154_n 0.0302777f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_16 VNB N_A2_c_183_n 0.0219728f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.345
cc_17 VNB N_A2_M1007_g 0.0116674f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.465
cc_18 VNB A2 0.0206727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_186_n 0.0444647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_207_n 0.0254721f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_21 VNB N_Y_c_208_n 0.0085488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Y 0.00309861f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_23 VNB N_Y_c_210_n 0.00263169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_276_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.51
cc_25 VNB N_VGND_c_311_n 0.0117008f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_26 VNB N_VGND_c_312_n 0.0247905f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_27 VNB N_VGND_c_313_n 0.0284864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_314_n 0.0136746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_315_n 0.034093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_316_n 0.026456f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.51
cc_31 VNB N_VGND_c_317_n 0.193373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_D1_M1005_g 0.0230655f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.465
cc_33 VPB N_D1_c_50_n 0.00263031f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.51
cc_34 VPB N_D1_c_51_n 0.00906229f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.51
cc_35 VPB N_C1_M1000_g 0.0192378f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.465
cc_36 VPB C1 0.00292672f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_37 VPB N_B1_M1004_g 0.0221866f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.655
cc_38 VPB N_A1_M1001_g 0.0225851f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.655
cc_39 VPB N_A2_M1007_g 0.0276856f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.465
cc_40 VPB N_Y_c_207_n 0.0559567f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.69
cc_41 VPB N_A_343_367#_c_254_n 0.0139898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_343_367#_c_255_n 0.0080198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_343_367#_c_256_n 0.0437226f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.51
cc_44 VPB N_VPWR_c_277_n 0.005617f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.465
cc_45 VPB N_VPWR_c_278_n 0.0663151f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_46 VPB N_VPWR_c_279_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.69
cc_47 VPB N_VPWR_c_280_n 0.0220565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_276_n 0.0502457f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.51
cc_49 N_D1_M1002_g N_C1_M1008_g 0.0225431f $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_50 N_D1_c_50_n N_C1_M1000_g 0.00387844f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_51 N_D1_c_51_n N_C1_M1000_g 0.0619479f $X=0.71 $Y=1.51 $X2=0 $Y2=0
cc_52 N_D1_M1002_g C1 5.01444e-19 $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_53 N_D1_M1005_g C1 0.00166332f $X=0.71 $Y=2.465 $X2=0 $Y2=0
cc_54 N_D1_c_50_n C1 0.120755f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_55 N_D1_c_51_n C1 0.00419796f $X=0.71 $Y=1.51 $X2=0 $Y2=0
cc_56 N_D1_c_50_n N_C1_c_84_n 0.00117584f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_57 N_D1_c_51_n N_C1_c_84_n 0.0122165f $X=0.71 $Y=1.51 $X2=0 $Y2=0
cc_58 N_D1_c_50_n N_Y_M1005_s 0.0117493f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_59 N_D1_M1002_g N_Y_c_207_n 0.0141289f $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_60 N_D1_M1005_g N_Y_c_207_n 0.0119721f $X=0.71 $Y=2.465 $X2=0 $Y2=0
cc_61 N_D1_c_50_n N_Y_c_207_n 0.118863f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_62 N_D1_M1002_g Y 0.0186917f $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_63 N_D1_c_50_n Y 0.00699286f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_64 N_D1_c_51_n Y 2.38553e-19 $X=0.71 $Y=1.51 $X2=0 $Y2=0
cc_65 N_D1_c_50_n N_Y_c_210_n 0.0182637f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_66 N_D1_c_51_n N_Y_c_210_n 0.00115713f $X=0.71 $Y=1.51 $X2=0 $Y2=0
cc_67 N_D1_c_50_n A_157_367# 0.00922154f $X=0.62 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_68 N_D1_M1005_g N_VPWR_c_278_n 0.00398598f $X=0.71 $Y=2.465 $X2=0 $Y2=0
cc_69 N_D1_c_50_n N_VPWR_c_278_n 0.00743808f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_70 N_D1_M1005_g N_VPWR_c_276_n 0.00698697f $X=0.71 $Y=2.465 $X2=0 $Y2=0
cc_71 N_D1_c_50_n N_VPWR_c_276_n 0.01011f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_72 N_D1_M1002_g N_VGND_c_312_n 0.0106461f $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_73 N_D1_M1002_g N_VGND_c_313_n 0.0058062f $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_74 N_D1_M1002_g N_VGND_c_317_n 0.00927162f $X=0.525 $Y=0.655 $X2=0 $Y2=0
cc_75 N_C1_M1000_g N_B1_M1004_g 0.0650432f $X=1.19 $Y=2.465 $X2=0 $Y2=0
cc_76 C1 N_B1_M1004_g 0.00889712f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_77 N_C1_M1008_g N_B1_c_120_n 0.0123118f $X=1.07 $Y=0.655 $X2=0 $Y2=0
cc_78 N_C1_M1008_g B1 5.28321e-19 $X=1.07 $Y=0.655 $X2=0 $Y2=0
cc_79 C1 B1 0.0246339f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 N_C1_c_84_n B1 0.00194705f $X=1.19 $Y=1.375 $X2=0 $Y2=0
cc_81 N_C1_M1008_g N_B1_c_122_n 4.68129e-19 $X=1.07 $Y=0.655 $X2=0 $Y2=0
cc_82 C1 N_B1_c_122_n 3.09362e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_83 N_C1_c_84_n N_B1_c_122_n 0.0206777f $X=1.19 $Y=1.375 $X2=0 $Y2=0
cc_84 C1 N_Y_c_207_n 0.00810802f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_C1_M1008_g N_Y_c_210_n 0.00388207f $X=1.07 $Y=0.655 $X2=0 $Y2=0
cc_86 N_C1_M1008_g N_Y_c_223_n 0.012357f $X=1.07 $Y=0.655 $X2=0 $Y2=0
cc_87 C1 N_Y_c_223_n 0.0182109f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_C1_c_84_n N_Y_c_223_n 0.00251758f $X=1.19 $Y=1.375 $X2=0 $Y2=0
cc_89 C1 A_157_367# 0.0117726f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_90 C1 N_A_343_367#_c_255_n 0.00350372f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_C1_M1000_g N_VPWR_c_278_n 0.00368922f $X=1.19 $Y=2.465 $X2=0 $Y2=0
cc_92 C1 N_VPWR_c_278_n 0.0119974f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_93 N_C1_M1000_g N_VPWR_c_276_n 0.00567429f $X=1.19 $Y=2.465 $X2=0 $Y2=0
cc_94 C1 N_VPWR_c_276_n 0.010176f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_95 N_C1_M1008_g N_VGND_c_312_n 5.39859e-19 $X=1.07 $Y=0.655 $X2=0 $Y2=0
cc_96 N_C1_M1008_g N_VGND_c_313_n 0.0165784f $X=1.07 $Y=0.655 $X2=0 $Y2=0
cc_97 N_C1_M1008_g N_VGND_c_317_n 0.00530063f $X=1.07 $Y=0.655 $X2=0 $Y2=0
cc_98 N_B1_M1004_g N_A1_M1001_g 0.0385818f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_99 N_B1_c_122_n N_A1_M1001_g 0.0104498f $X=1.85 $Y=1.355 $X2=0 $Y2=0
cc_100 N_B1_c_120_n N_A1_c_152_n 0.0282473f $X=1.85 $Y=1.19 $X2=0 $Y2=0
cc_101 N_B1_c_120_n A1 0.0022272f $X=1.85 $Y=1.19 $X2=0 $Y2=0
cc_102 B1 A1 0.0279408f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B1_c_120_n N_A1_c_154_n 0.0104498f $X=1.85 $Y=1.19 $X2=0 $Y2=0
cc_104 B1 N_A1_c_154_n 3.47656e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B1_c_120_n N_Y_c_223_n 0.015456f $X=1.85 $Y=1.19 $X2=0 $Y2=0
cc_106 B1 N_Y_c_223_n 0.0277509f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_107 N_B1_c_122_n N_Y_c_223_n 0.00132385f $X=1.85 $Y=1.355 $X2=0 $Y2=0
cc_108 N_B1_M1004_g N_A_343_367#_c_255_n 0.00174574f $X=1.64 $Y=2.465 $X2=0
+ $Y2=0
cc_109 B1 N_A_343_367#_c_255_n 0.00725039f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_110 N_B1_c_122_n N_A_343_367#_c_255_n 0.00312269f $X=1.85 $Y=1.355 $X2=0
+ $Y2=0
cc_111 N_B1_M1004_g N_VPWR_c_278_n 0.00585385f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_112 N_B1_M1004_g N_VPWR_c_276_n 0.0114101f $X=1.64 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B1_c_120_n N_VGND_c_313_n 0.0139339f $X=1.85 $Y=1.19 $X2=0 $Y2=0
cc_114 N_B1_c_120_n N_VGND_c_316_n 0.00487821f $X=1.85 $Y=1.19 $X2=0 $Y2=0
cc_115 N_B1_c_120_n N_VGND_c_317_n 0.00496998f $X=1.85 $Y=1.19 $X2=0 $Y2=0
cc_116 N_A1_c_152_n N_A2_c_183_n 0.0459218f $X=2.42 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_117 A1 N_A2_c_183_n 2.81786e-19 $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_118 A1 A2 0.0249238f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_119 N_A1_c_154_n A2 2.02927e-19 $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_120 N_A1_M1001_g N_A2_c_186_n 0.04047f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_121 A1 N_A2_c_186_n 0.00871013f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A1_c_154_n N_A2_c_186_n 0.0459218f $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_123 N_A1_c_152_n Y 0.0320932f $X=2.42 $Y=1.185 $X2=0 $Y2=0
cc_124 A1 Y 0.0490242f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A1_c_154_n Y 0.00530641f $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_126 N_A1_M1001_g N_A_343_367#_c_254_n 0.016527f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_127 A1 N_A_343_367#_c_254_n 0.0369648f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_128 N_A1_c_154_n N_A_343_367#_c_254_n 0.00503928f $X=2.42 $Y=1.35 $X2=0 $Y2=0
cc_129 A1 N_A_343_367#_c_255_n 0.00347299f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A1_M1001_g N_VPWR_c_277_n 0.00926406f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A1_M1001_g N_VPWR_c_278_n 0.00585385f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A1_M1001_g N_VPWR_c_276_n 0.0115207f $X=2.21 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A1_c_152_n N_VGND_c_313_n 0.00125958f $X=2.42 $Y=1.185 $X2=0 $Y2=0
cc_134 N_A1_c_152_n N_VGND_c_316_n 0.00357877f $X=2.42 $Y=1.185 $X2=0 $Y2=0
cc_135 N_A1_c_152_n N_VGND_c_317_n 0.00560459f $X=2.42 $Y=1.185 $X2=0 $Y2=0
cc_136 N_A2_c_183_n Y 0.0151709f $X=2.78 $Y=1.19 $X2=0 $Y2=0
cc_137 N_A2_M1007_g N_A_343_367#_c_254_n 0.0192643f $X=2.78 $Y=2.465 $X2=0 $Y2=0
cc_138 A2 N_A_343_367#_c_254_n 0.0169058f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A2_c_186_n N_A_343_367#_c_254_n 0.00745614f $X=2.99 $Y=1.355 $X2=0
+ $Y2=0
cc_140 N_A2_M1007_g N_VPWR_c_277_n 0.00908039f $X=2.78 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A2_M1007_g N_VPWR_c_280_n 0.00585385f $X=2.78 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A2_M1007_g N_VPWR_c_276_n 0.0121075f $X=2.78 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A2_c_183_n N_VGND_c_315_n 0.00619578f $X=2.78 $Y=1.19 $X2=0 $Y2=0
cc_144 A2 N_VGND_c_315_n 0.0202608f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_145 N_A2_c_186_n N_VGND_c_315_n 0.00596923f $X=2.99 $Y=1.355 $X2=0 $Y2=0
cc_146 N_A2_c_183_n N_VGND_c_316_n 0.0055505f $X=2.78 $Y=1.19 $X2=0 $Y2=0
cc_147 N_A2_c_183_n N_VGND_c_317_n 0.0108209f $X=2.78 $Y=1.19 $X2=0 $Y2=0
cc_148 N_Y_c_207_n N_VPWR_c_278_n 0.0174911f $X=0.28 $Y=1.98 $X2=0 $Y2=0
cc_149 N_Y_M1005_s N_VPWR_c_276_n 0.0100837f $X=0.155 $Y=1.835 $X2=0 $Y2=0
cc_150 N_Y_c_207_n N_VPWR_c_276_n 0.00964167f $X=0.28 $Y=1.98 $X2=0 $Y2=0
cc_151 N_Y_c_208_n N_VGND_M1002_s 0.00289679f $X=0.365 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_152 Y N_VGND_M1002_s 2.87015e-19 $X=0.635 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_153 N_Y_c_223_n N_VGND_M1008_d 0.0165732f $X=1.97 $Y=0.635 $X2=0 $Y2=0
cc_154 N_Y_c_208_n N_VGND_c_312_n 0.0207142f $X=0.365 $Y=1.07 $X2=0 $Y2=0
cc_155 Y N_VGND_c_312_n 0.00326589f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_156 N_Y_c_241_p N_VGND_c_313_n 0.0214254f $X=0.8 $Y=0.42 $X2=0 $Y2=0
cc_157 N_Y_c_223_n N_VGND_c_313_n 0.0435608f $X=1.97 $Y=0.635 $X2=0 $Y2=0
cc_158 Y N_VGND_c_316_n 0.0460537f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_159 N_Y_M1002_d N_VGND_c_317_n 0.00461686f $X=0.6 $Y=0.235 $X2=0 $Y2=0
cc_160 N_Y_M1009_d N_VGND_c_317_n 0.00369641f $X=1.925 $Y=0.235 $X2=0 $Y2=0
cc_161 Y N_VGND_c_317_n 0.0285606f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_162 N_Y_c_241_p N_VGND_c_317_n 0.0127519f $X=0.8 $Y=0.42 $X2=0 $Y2=0
cc_163 N_Y_c_223_n N_VGND_c_317_n 0.0119597f $X=1.97 $Y=0.635 $X2=0 $Y2=0
cc_164 Y A_499_47# 0.00200838f $X=2.555 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_165 A_157_367# N_VPWR_c_276_n 0.00874569f $X=0.785 $Y=1.835 $X2=0.695
+ $Y2=1.51
cc_166 A_253_367# N_VPWR_c_276_n 0.0111504f $X=1.265 $Y=1.835 $X2=3.12 $Y2=3.33
cc_167 N_A_343_367#_c_254_n N_VPWR_M1001_d 0.00362739f $X=2.89 $Y=1.84 $X2=-0.19
+ $Y2=1.655
cc_168 N_A_343_367#_c_254_n N_VPWR_c_277_n 0.0238538f $X=2.89 $Y=1.84 $X2=0
+ $Y2=0
cc_169 N_A_343_367#_c_270_p N_VPWR_c_278_n 0.0222962f $X=1.93 $Y=1.98 $X2=0
+ $Y2=0
cc_170 N_A_343_367#_c_256_n N_VPWR_c_280_n 0.0181659f $X=2.995 $Y=1.98 $X2=0
+ $Y2=0
cc_171 N_A_343_367#_M1004_d N_VPWR_c_276_n 0.00659813f $X=1.715 $Y=1.835 $X2=0
+ $Y2=0
cc_172 N_A_343_367#_M1007_d N_VPWR_c_276_n 0.00336915f $X=2.855 $Y=1.835 $X2=0
+ $Y2=0
cc_173 N_A_343_367#_c_270_p N_VPWR_c_276_n 0.0127519f $X=1.93 $Y=1.98 $X2=0
+ $Y2=0
cc_174 N_A_343_367#_c_256_n N_VPWR_c_276_n 0.0104192f $X=2.995 $Y=1.98 $X2=0
+ $Y2=0
cc_175 N_VGND_c_317_n A_499_47# 0.00168889f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
