* File: sky130_fd_sc_lp__o221a_4.spice
* Created: Fri Aug 28 11:07:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221a_4.pex.spice"
.subckt sky130_fd_sc_lp__o221a_4  VNB VPB C1 B1 B2 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1005 N_A_112_65#_M1005_d N_C1_M1005_g N_A_29_65#_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1014 N_A_112_65#_M1005_d N_C1_M1014_g N_A_29_65#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1015 N_A_29_65#_M1014_s N_B1_M1015_g N_A_284_65#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=5.712 M=1 R=5.6
+ SA=75001.1 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1003 N_A_284_65#_M1015_s N_B2_M1003_g N_A_29_65#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1020 N_A_284_65#_M1020_d N_B2_M1020_g N_A_29_65#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1023 N_A_29_65#_M1023_d N_B1_M1023_g N_A_284_65#_M1020_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_A_284_65#_M1002_d N_A1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_284_65#_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1010_d N_A2_M1017_g N_A_284_65#_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1008 N_A_284_65#_M1017_s N_A1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.856 M=1 R=5.6 SA=75001.5
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1008_s N_A_112_65#_M1004_g N_X_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A_112_65#_M1012_g N_X_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1021 N_VGND_M1012_d N_A_112_65#_M1021_g N_X_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1024_d N_A_112_65#_M1024_g N_X_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_C1_M1006_g N_A_112_65#_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75006.4 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_C1_M1022_g N_A_112_65#_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75006 A=0.189 P=2.82 MULT=1
MM1000 N_A_292_367#_M1000_d N_B1_M1000_g N_VPWR_M1022_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75001.1 SB=75005.5 A=0.189 P=2.82 MULT=1
MM1009 N_A_292_367#_M1000_d N_B2_M1009_g N_A_112_65#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75005.1 A=0.189 P=2.82 MULT=1
MM1018 N_A_292_367#_M1018_d N_B2_M1018_g N_A_112_65#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1026 N_A_292_367#_M1018_d N_B1_M1026_g N_VPWR_M1026_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.4599 PD=1.54 PS=1.99 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75004.2 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1026_s N_A1_M1007_g N_A_726_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.4599 AS=0.1764 PD=1.99 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.3
+ SB=75003.3 A=0.189 P=2.82 MULT=1
MM1016 N_A_726_367#_M1007_s N_A2_M1016_g N_A_112_65#_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1027 N_A_726_367#_M1027_d N_A2_M1027_g N_A_112_65#_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A1_M1011_g N_A_726_367#_M1027_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.26775 AS=0.1764 PD=1.685 PS=1.54 NRD=11.7215 NRS=0 M=1 R=8.4
+ SA=75004.5 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1001 N_X_M1001_d N_A_112_65#_M1001_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.26775 PD=1.54 PS=1.685 NRD=0 NRS=10.9335 M=1 R=8.4 SA=75005.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1013 N_X_M1001_d N_A_112_65#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1019 N_X_M1019_d N_A_112_65#_M1019_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1025 N_X_M1019_d N_A_112_65#_M1025_g N_VPWR_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75006.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=14.1367 P=18.89
*
.include "sky130_fd_sc_lp__o221a_4.pxi.spice"
*
.ends
*
*
