* File: sky130_fd_sc_lp__busdrivernovlpsleep_20.pxi.spice
* Created: Fri Aug 28 10:13:39 2020
* 
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%SLEEP N_SLEEP_M1030_g
+ N_SLEEP_M1026_g N_SLEEP_M1002_g N_SLEEP_M1006_g N_SLEEP_M1013_g
+ N_SLEEP_M1045_g N_SLEEP_M1049_g N_SLEEP_M1015_g N_SLEEP_M1046_g
+ N_SLEEP_c_459_n N_SLEEP_c_450_n N_SLEEP_c_460_n N_SLEEP_c_479_p
+ N_SLEEP_c_461_n N_SLEEP_c_549_p N_SLEEP_c_530_p N_SLEEP_c_531_p SLEEP
+ N_SLEEP_c_462_n N_SLEEP_c_451_n N_SLEEP_c_452_n N_SLEEP_c_453_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%SLEEP
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%TE_B N_TE_B_M1001_g N_TE_B_c_676_n
+ N_TE_B_c_677_n N_TE_B_c_670_n N_TE_B_M1008_g N_TE_B_M1040_g TE_B
+ N_TE_B_c_674_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%TE_B
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_27_47# N_A_27_47#_M1030_s
+ N_A_27_47#_M1026_s N_A_27_47#_M1036_g N_A_27_47#_M1066_g N_A_27_47#_c_729_n
+ N_A_27_47#_c_730_n N_A_27_47#_c_751_n N_A_27_47#_c_731_n N_A_27_47#_c_738_n
+ N_A_27_47#_c_732_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_27_47#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_280_47# N_A_280_47#_M1013_s
+ N_A_280_47#_M1008_s N_A_280_47#_M1001_d N_A_280_47#_M1035_g
+ N_A_280_47#_c_828_n N_A_280_47#_c_829_n N_A_280_47#_c_830_n
+ N_A_280_47#_c_831_n N_A_280_47#_M1011_g N_A_280_47#_M1063_g
+ N_A_280_47#_c_832_n N_A_280_47#_M1042_g N_A_280_47#_c_818_n
+ N_A_280_47#_c_819_n N_A_280_47#_M1037_g N_A_280_47#_c_821_n
+ N_A_280_47#_c_822_n N_A_280_47#_c_823_n N_A_280_47#_M1057_g
+ N_A_280_47#_c_825_n N_A_280_47#_c_983_p N_A_280_47#_c_826_n
+ N_A_280_47#_c_836_n N_A_280_47#_c_859_n N_A_280_47#_c_837_n
+ N_A_280_47#_c_884_n N_A_280_47#_c_838_n N_A_280_47#_c_905_n
+ N_A_280_47#_c_839_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_280_47#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_705_367# N_A_705_367#_M1005_s
+ N_A_705_367#_M1011_s N_A_705_367#_M1016_d N_A_705_367#_M1014_g
+ N_A_705_367#_c_997_n N_A_705_367#_c_998_n N_A_705_367#_c_999_n
+ N_A_705_367#_c_1000_n N_A_705_367#_M1027_g N_A_705_367#_c_1042_n
+ N_A_705_367#_M1004_g N_A_705_367#_c_1001_n N_A_705_367#_c_1002_n
+ N_A_705_367#_c_1045_n N_A_705_367#_M1010_g N_A_705_367#_c_1003_n
+ N_A_705_367#_c_1047_n N_A_705_367#_M1017_g N_A_705_367#_c_1004_n
+ N_A_705_367#_c_1049_n N_A_705_367#_M1019_g N_A_705_367#_c_1005_n
+ N_A_705_367#_c_1051_n N_A_705_367#_M1022_g N_A_705_367#_c_1006_n
+ N_A_705_367#_c_1053_n N_A_705_367#_M1024_g N_A_705_367#_c_1007_n
+ N_A_705_367#_c_1055_n N_A_705_367#_M1028_g N_A_705_367#_c_1008_n
+ N_A_705_367#_c_1057_n N_A_705_367#_M1031_g N_A_705_367#_c_1009_n
+ N_A_705_367#_c_1059_n N_A_705_367#_M1033_g N_A_705_367#_c_1010_n
+ N_A_705_367#_c_1061_n N_A_705_367#_M1034_g N_A_705_367#_c_1011_n
+ N_A_705_367#_c_1063_n N_A_705_367#_M1039_g N_A_705_367#_c_1012_n
+ N_A_705_367#_c_1065_n N_A_705_367#_M1043_g N_A_705_367#_c_1066_n
+ N_A_705_367#_M1051_g N_A_705_367#_c_1067_n N_A_705_367#_M1053_g
+ N_A_705_367#_c_1068_n N_A_705_367#_M1054_g N_A_705_367#_c_1069_n
+ N_A_705_367#_M1060_g N_A_705_367#_c_1070_n N_A_705_367#_M1061_g
+ N_A_705_367#_c_1071_n N_A_705_367#_M1064_g N_A_705_367#_c_1072_n
+ N_A_705_367#_M1070_g N_A_705_367#_c_1073_n N_A_705_367#_M1072_g
+ N_A_705_367#_c_1013_n N_A_705_367#_c_1014_n N_A_705_367#_c_1015_n
+ N_A_705_367#_c_1016_n N_A_705_367#_c_1017_n N_A_705_367#_c_1018_n
+ N_A_705_367#_c_1019_n N_A_705_367#_c_1020_n N_A_705_367#_c_1021_n
+ N_A_705_367#_c_1022_n N_A_705_367#_c_1084_n N_A_705_367#_c_1023_n
+ N_A_705_367#_c_1139_n N_A_705_367#_c_1024_n N_A_705_367#_c_1025_n
+ N_A_705_367#_c_1260_p N_A_705_367#_c_1086_n N_A_705_367#_c_1087_n
+ N_A_705_367#_c_1276_p N_A_705_367#_c_1026_n N_A_705_367#_c_1027_n
+ N_A_705_367#_c_1028_n N_A_705_367#_c_1029_n N_A_705_367#_c_1030_n
+ N_A_705_367#_c_1031_n N_A_705_367#_c_1032_n N_A_705_367#_c_1033_n
+ N_A_705_367#_c_1034_n N_A_705_367#_c_1035_n N_A_705_367#_c_1036_n
+ N_A_705_367#_c_1037_n N_A_705_367#_c_1038_n N_A_705_367#_c_1039_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_705_367#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_407_491# N_A_407_491#_M1063_s
+ N_A_407_491#_M1035_s N_A_407_491#_c_1550_n N_A_407_491#_c_1551_n
+ N_A_407_491#_c_1552_n N_A_407_491#_c_1553_n N_A_407_491#_M1038_g
+ N_A_407_491#_c_1554_n N_A_407_491#_c_1555_n N_A_407_491#_M1050_g
+ N_A_407_491#_c_1556_n N_A_407_491#_M1018_g N_A_407_491#_M1020_g
+ N_A_407_491#_c_1559_n N_A_407_491#_c_1560_n N_A_407_491#_c_1572_n
+ N_A_407_491#_c_1573_n N_A_407_491#_c_1574_n N_A_407_491#_c_1561_n
+ N_A_407_491#_c_1562_n N_A_407_491#_c_1563_n N_A_407_491#_c_1564_n
+ N_A_407_491#_c_1739_p N_A_407_491#_c_1565_n N_A_407_491#_c_1566_n
+ N_A_407_491#_c_1567_n N_A_407_491#_c_1648_p N_A_407_491#_c_1649_p
+ N_A_407_491#_c_1650_p N_A_407_491#_c_1689_p N_A_407_491#_c_1568_n
+ N_A_407_491#_c_1669_p N_A_407_491#_c_1569_n N_A_407_491#_c_1570_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_407_491#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_896_367# N_A_896_367#_M1014_d
+ N_A_896_367#_M1036_s N_A_896_367#_M1057_d N_A_896_367#_c_1764_n
+ N_A_896_367#_c_1774_n N_A_896_367#_M1023_g N_A_896_367#_c_1765_n
+ N_A_896_367#_c_1776_n N_A_896_367#_M1067_g N_A_896_367#_c_1766_n
+ N_A_896_367#_c_1884_p N_A_896_367#_c_1778_n N_A_896_367#_c_1767_n
+ N_A_896_367#_c_1768_n N_A_896_367#_c_1769_n N_A_896_367#_c_1770_n
+ N_A_896_367#_c_1779_n N_A_896_367#_c_1771_n N_A_896_367#_c_1795_n
+ N_A_896_367#_c_1781_n N_A_896_367#_c_1809_n N_A_896_367#_c_1772_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_896_367#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_1486_47# N_A_1486_47#_M1038_d
+ N_A_1486_47#_M1003_d N_A_1486_47#_M1023_d N_A_1486_47#_M1068_g
+ N_A_1486_47#_M1065_g N_A_1486_47#_M1000_g N_A_1486_47#_M1009_g
+ N_A_1486_47#_M1021_g N_A_1486_47#_M1025_g N_A_1486_47#_c_1924_n
+ N_A_1486_47#_M1029_g N_A_1486_47#_c_1925_n N_A_1486_47#_M1032_g
+ N_A_1486_47#_c_1926_n N_A_1486_47#_M1047_g N_A_1486_47#_c_1927_n
+ N_A_1486_47#_M1048_g N_A_1486_47#_c_1928_n N_A_1486_47#_c_1929_n
+ N_A_1486_47#_c_1930_n N_A_1486_47#_M1052_g N_A_1486_47#_c_1931_n
+ N_A_1486_47#_c_1932_n N_A_1486_47#_M1056_g N_A_1486_47#_c_1933_n
+ N_A_1486_47#_c_1934_n N_A_1486_47#_M1058_g N_A_1486_47#_c_1935_n
+ N_A_1486_47#_c_1936_n N_A_1486_47#_M1059_g N_A_1486_47#_c_1937_n
+ N_A_1486_47#_c_1938_n N_A_1486_47#_M1062_g N_A_1486_47#_c_1939_n
+ N_A_1486_47#_c_1940_n N_A_1486_47#_M1073_g N_A_1486_47#_c_1941_n
+ N_A_1486_47#_c_1942_n N_A_1486_47#_c_1943_n N_A_1486_47#_c_1944_n
+ N_A_1486_47#_c_1945_n N_A_1486_47#_c_1946_n N_A_1486_47#_c_1947_n
+ N_A_1486_47#_c_2028_n N_A_1486_47#_c_1948_n N_A_1486_47#_c_1949_n
+ N_A_1486_47#_c_1950_n N_A_1486_47#_c_1951_n N_A_1486_47#_c_1952_n
+ N_A_1486_47#_c_1953_n N_A_1486_47#_c_1954_n N_A_1486_47#_c_1955_n
+ N_A_1486_47#_c_1956_n N_A_1486_47#_c_1957_n N_A_1486_47#_c_1958_n
+ N_A_1486_47#_c_1959_n N_A_1486_47#_c_1960_n N_A_1486_47#_c_1961_n
+ N_A_1486_47#_c_1962_n N_A_1486_47#_c_1963_n N_A_1486_47#_c_1964_n
+ N_A_1486_47#_c_1965_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_1486_47#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A N_A_c_2281_n N_A_M1012_g
+ N_A_M1003_g N_A_c_2282_n N_A_M1044_g N_A_M1071_g N_A_c_2283_n N_A_c_2284_n
+ N_A_c_2285_n N_A_c_2286_n N_A_c_2265_n N_A_c_2266_n N_A_c_2267_n N_A_c_2268_n
+ N_A_M1007_g N_A_c_2289_n N_A_M1016_g N_A_c_2270_n N_A_M1041_g N_A_c_2291_n
+ N_A_M1069_g N_A_c_2272_n N_A_c_2273_n N_A_c_2274_n N_A_c_2275_n N_A_c_2276_n
+ N_A_c_2277_n N_A_c_2278_n N_A_c_2279_n A A
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_2063_47# N_A_2063_47#_M1020_d
+ N_A_2063_47#_M1068_d N_A_2063_47#_M1005_g N_A_2063_47#_c_2481_n
+ N_A_2063_47#_c_2482_n N_A_2063_47#_M1055_g N_A_2063_47#_c_2605_p
+ N_A_2063_47#_c_2483_n N_A_2063_47#_c_2484_n N_A_2063_47#_c_2485_n
+ N_A_2063_47#_c_2486_n N_A_2063_47#_c_2487_n N_A_2063_47#_c_2488_n
+ N_A_2063_47#_c_2489_n N_A_2063_47#_c_2490_n N_A_2063_47#_c_2495_n
+ N_A_2063_47#_c_2496_n N_A_2063_47#_c_2491_n N_A_2063_47#_c_2492_n
+ N_A_2063_47#_c_2493_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_2063_47#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%VPWR N_VPWR_M1026_d N_VPWR_M1049_s
+ N_VPWR_M1027_d N_VPWR_M1012_s N_VPWR_M1018_s N_VPWR_M1015_d N_VPWR_M1046_d
+ N_VPWR_M1004_s N_VPWR_M1010_s N_VPWR_M1019_s N_VPWR_M1024_s N_VPWR_M1031_s
+ N_VPWR_M1034_s N_VPWR_M1043_s N_VPWR_M1053_s N_VPWR_M1060_s N_VPWR_M1064_s
+ N_VPWR_M1072_s N_VPWR_c_2628_n N_VPWR_c_2629_n N_VPWR_c_2630_n N_VPWR_c_2631_n
+ N_VPWR_c_2632_n N_VPWR_c_2633_n N_VPWR_c_2634_n N_VPWR_c_2635_n
+ N_VPWR_c_2636_n N_VPWR_c_2637_n N_VPWR_c_2638_n N_VPWR_c_2639_n
+ N_VPWR_c_2640_n N_VPWR_c_2641_n N_VPWR_c_2642_n N_VPWR_c_2643_n
+ N_VPWR_c_2644_n N_VPWR_c_2645_n N_VPWR_c_2646_n N_VPWR_c_2647_n
+ N_VPWR_c_2648_n N_VPWR_c_2649_n N_VPWR_c_2650_n N_VPWR_c_2651_n
+ N_VPWR_c_2652_n N_VPWR_c_2653_n N_VPWR_c_2654_n N_VPWR_c_2655_n
+ N_VPWR_c_2656_n N_VPWR_c_2657_n N_VPWR_c_2658_n N_VPWR_c_2659_n
+ N_VPWR_c_2660_n N_VPWR_c_2661_n N_VPWR_c_2662_n N_VPWR_c_2663_n
+ N_VPWR_c_2664_n N_VPWR_c_2665_n VPWR N_VPWR_c_2666_n N_VPWR_c_2667_n
+ N_VPWR_c_2668_n N_VPWR_c_2669_n N_VPWR_c_2670_n N_VPWR_c_2671_n
+ N_VPWR_c_2672_n N_VPWR_c_2673_n N_VPWR_c_2627_n N_VPWR_c_2675_n
+ N_VPWR_c_2676_n N_VPWR_c_2677_n N_VPWR_c_2678_n N_VPWR_c_2679_n
+ N_VPWR_c_2680_n N_VPWR_c_2681_n N_VPWR_c_2682_n N_VPWR_c_2683_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%VPWR
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%KAPWR N_KAPWR_M1035_d
+ N_KAPWR_M1042_d N_KAPWR_M1066_d KAPWR N_KAPWR_c_3047_n N_KAPWR_c_3065_n
+ N_KAPWR_c_3048_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%KAPWR
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_1492_367# N_A_1492_367#_M1023_s
+ N_A_1492_367#_M1067_s N_A_1492_367#_M1044_d N_A_1492_367#_c_3248_n
+ N_A_1492_367#_c_3237_n N_A_1492_367#_c_3255_n N_A_1492_367#_c_3238_n
+ N_A_1492_367#_c_3258_n N_A_1492_367#_c_3244_n N_A_1492_367#_c_3260_n
+ N_A_1492_367#_c_3239_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_1492_367#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_2345_367# N_A_2345_367#_M1015_s
+ N_A_2345_367#_M1016_s N_A_2345_367#_M1069_s N_A_2345_367#_c_3306_n
+ N_A_2345_367#_c_3307_n N_A_2345_367#_c_3308_n N_A_2345_367#_c_3327_n
+ N_A_2345_367#_c_3309_n N_A_2345_367#_c_3310_n N_A_2345_367#_c_3311_n
+ N_A_2345_367#_c_3318_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_2345_367#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%Z N_Z_M1000_s N_Z_M1009_s
+ N_Z_M1025_s N_Z_M1032_s N_Z_M1048_s N_Z_M1056_s N_Z_M1059_s N_Z_M1073_s
+ N_Z_M1004_d N_Z_M1017_d N_Z_M1022_d N_Z_M1028_d N_Z_M1033_d N_Z_M1039_d
+ N_Z_M1051_d N_Z_M1054_d N_Z_M1061_d N_Z_M1070_d N_Z_c_3375_n N_Z_c_3564_n
+ N_Z_c_3379_n N_Z_c_3367_n N_Z_c_3393_n Z N_Z_c_3368_n N_Z_c_3369_n
+ N_Z_c_3370_n N_Z_c_3371_n N_Z_c_3372_n N_Z_c_3373_n N_Z_c_3374_n N_Z_c_3454_n
+ N_Z_c_3460_n N_Z_c_3492_n Z PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%Z
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%VGND N_VGND_M1002_d N_VGND_M1045_d
+ N_VGND_M1040_d N_VGND_M1063_d N_VGND_M1038_s N_VGND_M1050_s N_VGND_M1071_s
+ N_VGND_M1065_d N_VGND_M1007_d N_VGND_M1000_d N_VGND_M1021_d N_VGND_M1029_d
+ N_VGND_M1047_d N_VGND_M1052_d N_VGND_M1058_d N_VGND_M1062_d N_VGND_c_3664_n
+ N_VGND_c_3665_n N_VGND_c_3666_n N_VGND_c_3667_n N_VGND_c_3668_n
+ N_VGND_c_3669_n N_VGND_c_3670_n N_VGND_c_3671_n N_VGND_c_3672_n
+ N_VGND_c_3673_n N_VGND_c_3674_n N_VGND_c_3675_n N_VGND_c_3676_n
+ N_VGND_c_3677_n N_VGND_c_3678_n N_VGND_c_3679_n N_VGND_c_3680_n
+ N_VGND_c_3681_n N_VGND_c_3682_n N_VGND_c_3683_n N_VGND_c_3684_n
+ N_VGND_c_3685_n N_VGND_c_3686_n N_VGND_c_3687_n N_VGND_c_3688_n
+ N_VGND_c_3689_n N_VGND_c_3690_n N_VGND_c_3691_n N_VGND_c_3692_n
+ N_VGND_c_3693_n N_VGND_c_3694_n N_VGND_c_3695_n N_VGND_c_3696_n
+ N_VGND_c_3697_n N_VGND_c_3698_n N_VGND_c_3699_n N_VGND_c_3700_n
+ N_VGND_c_3701_n N_VGND_c_3702_n N_VGND_c_3703_n VGND N_VGND_c_3704_n
+ N_VGND_c_3705_n N_VGND_c_3706_n N_VGND_c_3707_n N_VGND_c_3708_n
+ N_VGND_c_3709_n N_VGND_c_3710_n N_VGND_c_3711_n N_VGND_c_3712_n
+ N_VGND_c_3713_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%VGND
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_2519_47# N_A_2519_47#_M1007_s
+ N_A_2519_47#_M1041_s N_A_2519_47#_M1055_d N_A_2519_47#_c_3971_n
+ N_A_2519_47#_c_3956_n N_A_2519_47#_c_3957_n N_A_2519_47#_c_3989_n
+ N_A_2519_47#_c_3990_n N_A_2519_47#_c_3961_n N_A_2519_47#_c_3958_n
+ N_A_2519_47#_c_3959_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_2519_47#
cc_1 VNB N_SLEEP_M1030_g 0.0478893f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_2 VNB N_SLEEP_M1026_g 0.00523536f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.595
cc_3 VNB N_SLEEP_M1002_g 0.0397434f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.445
cc_4 VNB N_SLEEP_M1006_g 0.00475907f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.775
cc_5 VNB N_SLEEP_M1013_g 0.0201503f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=0.655
cc_6 VNB N_SLEEP_M1045_g 0.0195014f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=0.655
cc_7 VNB N_SLEEP_c_450_n 0.0020826f $X=-0.19 $Y=-0.245 $X2=11.95 $Y2=1.445
cc_8 VNB N_SLEEP_c_451_n 0.00863145f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.415
cc_9 VNB N_SLEEP_c_452_n 0.0927393f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.415
cc_10 VNB N_SLEEP_c_453_n 0.049109f $X=-0.19 $Y=-0.245 $X2=12.08 $Y2=1.475
cc_11 VNB N_TE_B_c_670_n 0.00489902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_TE_B_M1008_g 0.0170997f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.445
cc_13 VNB N_TE_B_M1040_g 0.02155f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.775
cc_14 VNB TE_B 0.0069706f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.25
cc_15 VNB N_TE_B_c_674_n 0.0524379f $X=-0.19 $Y=-0.245 $X2=5.785 $Y2=2.095
cc_16 VNB N_A_27_47#_c_729_n 0.0208388f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.775
cc_17 VNB N_A_27_47#_c_730_n 0.00414678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_731_n 0.0498952f $X=-0.19 $Y=-0.245 $X2=5.785 $Y2=2.675
cc_19 VNB N_A_27_47#_c_732_n 0.0550616f $X=-0.19 $Y=-0.245 $X2=11.65 $Y2=1.67
cc_20 VNB N_A_280_47#_M1063_g 0.0371167f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=0.655
cc_21 VNB N_A_280_47#_c_818_n 0.0530071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_280_47#_c_819_n 0.133123f $X=-0.19 $Y=-0.245 $X2=11.65 $Y2=1.67
cc_23 VNB N_A_280_47#_M1037_g 0.0299592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_280_47#_c_821_n 0.0233633f $X=-0.19 $Y=-0.245 $X2=12.08 $Y2=2.465
cc_25 VNB N_A_280_47#_c_822_n 0.0498555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_280_47#_c_823_n 0.0110273f $X=-0.19 $Y=-0.245 $X2=5.71 $Y2=1.93
cc_27 VNB N_A_280_47#_M1057_g 0.00542098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_280_47#_c_825_n 0.0043695f $X=-0.19 $Y=-0.245 $X2=11.95 $Y2=1.445
cc_29 VNB N_A_280_47#_c_826_n 0.00475237f $X=-0.19 $Y=-0.245 $X2=5.645 $Y2=2.035
cc_30 VNB N_A_705_367#_M1014_g 0.035202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_705_367#_c_997_n 0.0565566f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.775
cc_32 VNB N_A_705_367#_c_998_n 0.00675945f $X=-0.19 $Y=-0.245 $X2=1.065
+ $Y2=2.775
cc_33 VNB N_A_705_367#_c_999_n 0.0221419f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.25
cc_34 VNB N_A_705_367#_c_1000_n 0.00957217f $X=-0.19 $Y=-0.245 $X2=1.325
+ $Y2=0.655
cc_35 VNB N_A_705_367#_c_1001_n 0.0103042f $X=-0.19 $Y=-0.245 $X2=5.785
+ $Y2=2.095
cc_36 VNB N_A_705_367#_c_1002_n 0.0052103f $X=-0.19 $Y=-0.245 $X2=5.785
+ $Y2=2.675
cc_37 VNB N_A_705_367#_c_1003_n 0.00532452f $X=-0.19 $Y=-0.245 $X2=11.65
+ $Y2=2.465
cc_38 VNB N_A_705_367#_c_1004_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=12.08
+ $Y2=2.465
cc_39 VNB N_A_705_367#_c_1005_n 0.00536775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_705_367#_c_1006_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=5.355
+ $Y2=2.035
cc_41 VNB N_A_705_367#_c_1007_n 0.00536775f $X=-0.19 $Y=-0.245 $X2=5.5 $Y2=2.035
cc_42 VNB N_A_705_367#_c_1008_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_705_367#_c_1009_n 0.00536775f $X=-0.19 $Y=-0.245 $X2=5.51 $Y2=1.93
cc_44 VNB N_A_705_367#_c_1010_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.415
cc_45 VNB N_A_705_367#_c_1011_n 0.00536775f $X=-0.19 $Y=-0.245 $X2=1.755
+ $Y2=1.415
cc_46 VNB N_A_705_367#_c_1012_n 0.0075543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_705_367#_c_1013_n 0.00430336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_705_367#_c_1014_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_705_367#_c_1015_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_705_367#_c_1016_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_705_367#_c_1017_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_705_367#_c_1018_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_705_367#_c_1019_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_705_367#_c_1020_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_705_367#_c_1021_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_705_367#_c_1022_n 0.00385496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_705_367#_c_1023_n 0.0230132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_705_367#_c_1024_n 0.0044896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_705_367#_c_1025_n 0.00407275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_705_367#_c_1026_n 0.00771272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_705_367#_c_1027_n 8.93368e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_705_367#_c_1028_n 9.9273e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_705_367#_c_1029_n 0.0122055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_705_367#_c_1030_n 0.0010183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_705_367#_c_1031_n 0.00426465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_705_367#_c_1032_n 0.0161415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_705_367#_c_1033_n 0.0024063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_705_367#_c_1034_n 0.00173813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_705_367#_c_1035_n 0.00173813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_705_367#_c_1036_n 0.00173813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_705_367#_c_1037_n 0.216896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_705_367#_c_1038_n 0.0225506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_705_367#_c_1039_n 7.68132e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_407_491#_c_1550_n 0.0197983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_407_491#_c_1551_n 0.0136559f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.25
cc_76 VNB N_A_407_491#_c_1552_n 0.00828505f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.445
cc_77 VNB N_A_407_491#_c_1553_n 0.0210659f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.445
cc_78 VNB N_A_407_491#_c_1554_n 0.0388288f $X=-0.19 $Y=-0.245 $X2=1.065
+ $Y2=2.775
cc_79 VNB N_A_407_491#_c_1555_n 0.0194352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_407_491#_c_1556_n 0.0359803f $X=-0.19 $Y=-0.245 $X2=1.325
+ $Y2=0.655
cc_81 VNB N_A_407_491#_M1018_g 0.0188969f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=1.25
cc_82 VNB N_A_407_491#_M1020_g 0.0335598f $X=-0.19 $Y=-0.245 $X2=5.785 $Y2=2.095
cc_83 VNB N_A_407_491#_c_1559_n 0.0560598f $X=-0.19 $Y=-0.245 $X2=5.785
+ $Y2=2.675
cc_84 VNB N_A_407_491#_c_1560_n 0.00514745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_407_491#_c_1561_n 0.0054889f $X=-0.19 $Y=-0.245 $X2=12.08
+ $Y2=2.465
cc_86 VNB N_A_407_491#_c_1562_n 0.0052449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_407_491#_c_1563_n 0.0188131f $X=-0.19 $Y=-0.245 $X2=5.71 $Y2=1.93
cc_88 VNB N_A_407_491#_c_1564_n 0.0152093f $X=-0.19 $Y=-0.245 $X2=11.95 $Y2=1.47
cc_89 VNB N_A_407_491#_c_1565_n 0.00323848f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=2.035
cc_90 VNB N_A_407_491#_c_1566_n 0.00269144f $X=-0.19 $Y=-0.245 $X2=5.645
+ $Y2=2.035
cc_91 VNB N_A_407_491#_c_1567_n 0.00274797f $X=-0.19 $Y=-0.245 $X2=5.5 $Y2=2.035
cc_92 VNB N_A_407_491#_c_1568_n 0.00918455f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_93 VNB N_A_407_491#_c_1569_n 3.8413e-19 $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.415
cc_94 VNB N_A_407_491#_c_1570_n 0.00368024f $X=-0.19 $Y=-0.245 $X2=0.76
+ $Y2=1.415
cc_95 VNB N_A_896_367#_c_1764_n 0.0110305f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.445
cc_96 VNB N_A_896_367#_c_1765_n 0.0138902f $X=-0.19 $Y=-0.245 $X2=1.065
+ $Y2=2.775
cc_97 VNB N_A_896_367#_c_1766_n 0.0040035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_896_367#_c_1767_n 0.0112146f $X=-0.19 $Y=-0.245 $X2=5.785
+ $Y2=2.675
cc_99 VNB N_A_896_367#_c_1768_n 0.00468969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_896_367#_c_1769_n 0.00743501f $X=-0.19 $Y=-0.245 $X2=12.08
+ $Y2=2.465
cc_101 VNB N_A_896_367#_c_1770_n 0.00299368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_896_367#_c_1771_n 0.00973466f $X=-0.19 $Y=-0.245 $X2=11.95
+ $Y2=1.445
cc_103 VNB N_A_896_367#_c_1772_n 0.0080585f $X=-0.19 $Y=-0.245 $X2=11.865
+ $Y2=2.035
cc_104 VNB N_A_1486_47#_M1065_g 0.0306354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1486_47#_M1000_g 0.023129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1486_47#_M1009_g 0.0180558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1486_47#_M1021_g 0.0180558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1486_47#_M1025_g 0.0180558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1486_47#_c_1924_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=12.08
+ $Y2=2.465
cc_110 VNB N_A_1486_47#_c_1925_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=5.71 $Y2=1.93
cc_111 VNB N_A_1486_47#_c_1926_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1486_47#_c_1927_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=11.95
+ $Y2=1.445
cc_113 VNB N_A_1486_47#_c_1928_n 0.0124835f $X=-0.19 $Y=-0.245 $X2=0.915
+ $Y2=2.035
cc_114 VNB N_A_1486_47#_c_1929_n 0.176985f $X=-0.19 $Y=-0.245 $X2=11.72
+ $Y2=2.035
cc_115 VNB N_A_1486_47#_c_1930_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=5.645
+ $Y2=2.035
cc_116 VNB N_A_1486_47#_c_1931_n 0.0112546f $X=-0.19 $Y=-0.245 $X2=5.5 $Y2=2.035
cc_117 VNB N_A_1486_47#_c_1932_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=11.865
+ $Y2=2.035
cc_118 VNB N_A_1486_47#_c_1933_n 0.0101163f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.95
cc_119 VNB N_A_1486_47#_c_1934_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=5.51 $Y2=1.93
cc_120 VNB N_A_1486_47#_c_1935_n 0.0112546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_1486_47#_c_1936_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.415
cc_122 VNB N_A_1486_47#_c_1937_n 0.0101163f $X=-0.19 $Y=-0.245 $X2=0.76
+ $Y2=1.415
cc_123 VNB N_A_1486_47#_c_1938_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=1.065
+ $Y2=1.415
cc_124 VNB N_A_1486_47#_c_1939_n 0.020322f $X=-0.19 $Y=-0.245 $X2=11.65
+ $Y2=1.475
cc_125 VNB N_A_1486_47#_c_1940_n 0.0200313f $X=-0.19 $Y=-0.245 $X2=11.95
+ $Y2=1.475
cc_126 VNB N_A_1486_47#_c_1941_n 0.024136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_1486_47#_c_1942_n 0.0144693f $X=-0.19 $Y=-0.245 $X2=0.76
+ $Y2=2.035
cc_128 VNB N_A_1486_47#_c_1943_n 0.00578834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_1486_47#_c_1944_n 0.00478657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_1486_47#_c_1945_n 0.00478657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_1486_47#_c_1946_n 0.00478657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_1486_47#_c_1947_n 0.00478657f $X=-0.19 $Y=-0.245 $X2=11.882
+ $Y2=2.035
cc_133 VNB N_A_1486_47#_c_1948_n 0.0115295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_1486_47#_c_1949_n 0.0107928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_1486_47#_c_1950_n 0.00227985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_1486_47#_c_1951_n 0.0080974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_1486_47#_c_1952_n 0.00104784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_1486_47#_c_1953_n 0.0327059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_1486_47#_c_1954_n 0.0019175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_1486_47#_c_1955_n 0.00111797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_1486_47#_c_1956_n 0.0152829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_A_1486_47#_c_1957_n 0.00548335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_1486_47#_c_1958_n 0.00460804f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_1486_47#_c_1959_n 0.015033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_A_1486_47#_c_1960_n 0.0715265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_A_1486_47#_c_1961_n 0.00921911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_1486_47#_c_1962_n 0.00365776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_A_1486_47#_c_1963_n 0.00365776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_A_1486_47#_c_1964_n 0.00273005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_A_1486_47#_c_1965_n 0.00273005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_A_M1003_g 0.0342429f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.595
cc_152 VNB N_A_M1071_g 0.0323419f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.58
cc_153 VNB N_A_c_2265_n 0.0102599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_A_c_2266_n 0.0345499f $X=-0.19 $Y=-0.245 $X2=5.785 $Y2=2.675
cc_155 VNB N_A_c_2267_n 0.00763766f $X=-0.19 $Y=-0.245 $X2=5.785 $Y2=2.675
cc_156 VNB N_A_c_2268_n 0.00210766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_A_M1007_g 0.038982f $X=-0.19 $Y=-0.245 $X2=11.65 $Y2=2.465
cc_158 VNB N_A_c_2270_n 0.0077642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_A_M1041_g 0.0348444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_A_c_2272_n 0.0527294f $X=-0.19 $Y=-0.245 $X2=5.645 $Y2=2.035
cc_161 VNB N_A_c_2273_n 0.0340938f $X=-0.19 $Y=-0.245 $X2=5.5 $Y2=2.035
cc_162 VNB N_A_c_2274_n 0.00379481f $X=-0.19 $Y=-0.245 $X2=5.5 $Y2=2.035
cc_163 VNB N_A_c_2275_n 0.0335918f $X=-0.19 $Y=-0.245 $X2=11.865 $Y2=2.035
cc_164 VNB N_A_c_2276_n 0.0105327f $X=-0.19 $Y=-0.245 $X2=11.865 $Y2=2.035
cc_165 VNB N_A_c_2277_n 0.0941969f $X=-0.19 $Y=-0.245 $X2=11.865 $Y2=2.035
cc_166 VNB N_A_c_2278_n 0.00222282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_A_c_2279_n 0.00326886f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_168 VNB A 0.00448178f $X=-0.19 $Y=-0.245 $X2=5.51 $Y2=1.93
cc_169 VNB N_A_2063_47#_c_2481_n 0.0207339f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.445
cc_170 VNB N_A_2063_47#_c_2482_n 0.018846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_A_2063_47#_c_2483_n 0.00505707f $X=-0.19 $Y=-0.245 $X2=1.755
+ $Y2=1.25
cc_172 VNB N_A_2063_47#_c_2484_n 0.00379473f $X=-0.19 $Y=-0.245 $X2=1.755
+ $Y2=0.655
cc_173 VNB N_A_2063_47#_c_2485_n 0.00137975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_A_2063_47#_c_2486_n 0.00249903f $X=-0.19 $Y=-0.245 $X2=5.785
+ $Y2=2.675
cc_175 VNB N_A_2063_47#_c_2487_n 0.0216394f $X=-0.19 $Y=-0.245 $X2=5.785
+ $Y2=2.675
cc_176 VNB N_A_2063_47#_c_2488_n 0.00385664f $X=-0.19 $Y=-0.245 $X2=11.65
+ $Y2=2.465
cc_177 VNB N_A_2063_47#_c_2489_n 0.00324898f $X=-0.19 $Y=-0.245 $X2=11.65
+ $Y2=2.465
cc_178 VNB N_A_2063_47#_c_2490_n 0.00570023f $X=-0.19 $Y=-0.245 $X2=12.08
+ $Y2=1.67
cc_179 VNB N_A_2063_47#_c_2491_n 0.00127745f $X=-0.19 $Y=-0.245 $X2=11.95
+ $Y2=1.47
cc_180 VNB N_A_2063_47#_c_2492_n 0.0401706f $X=-0.19 $Y=-0.245 $X2=11.95
+ $Y2=1.445
cc_181 VNB N_A_2063_47#_c_2493_n 0.0168593f $X=-0.19 $Y=-0.245 $X2=11.95
+ $Y2=1.445
cc_182 VNB N_VPWR_c_2627_n 0.97968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_Z_c_3367_n 0.0203284f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.415
cc_184 VNB N_Z_c_3368_n 0.00437785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_Z_c_3369_n 0.00437785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_Z_c_3370_n 0.00437785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_Z_c_3371_n 0.00844534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_Z_c_3372_n 0.00549438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_189 VNB N_Z_c_3373_n 0.00549438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_190 VNB N_Z_c_3374_n 0.045274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_191 VNB N_VGND_c_3664_n 0.00928816f $X=-0.19 $Y=-0.245 $X2=5.5 $Y2=2.035
cc_192 VNB N_VGND_c_3665_n 3.22914e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_193 VNB N_VGND_c_3666_n 0.0130914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_194 VNB N_VGND_c_3667_n 0.0108519f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=1.415
cc_195 VNB N_VGND_c_3668_n 0.00277956f $X=-0.19 $Y=-0.245 $X2=1.325 $Y2=1.415
cc_196 VNB N_VGND_c_3669_n 0.0122192f $X=-0.19 $Y=-0.245 $X2=11.65 $Y2=1.475
cc_197 VNB N_VGND_c_3670_n 0.0110989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_198 VNB N_VGND_c_3671_n 0.00546467f $X=-0.19 $Y=-0.245 $X2=0.77 $Y2=2.035
cc_199 VNB N_VGND_c_3672_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_200 VNB N_VGND_c_3673_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.035
cc_201 VNB N_VGND_c_3674_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_202 VNB N_VGND_c_3675_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_203 VNB N_VGND_c_3676_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_204 VNB N_VGND_c_3677_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_205 VNB N_VGND_c_3678_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_206 VNB N_VGND_c_3679_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_207 VNB N_VGND_c_3680_n 0.0290019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_208 VNB N_VGND_c_3681_n 0.0058666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_209 VNB N_VGND_c_3682_n 0.0145469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_210 VNB N_VGND_c_3683_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_211 VNB N_VGND_c_3684_n 0.0151002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_212 VNB N_VGND_c_3685_n 0.00528623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_213 VNB N_VGND_c_3686_n 0.0157231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_214 VNB N_VGND_c_3687_n 0.0179442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_215 VNB N_VGND_c_3688_n 0.0454967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_216 VNB N_VGND_c_3689_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_217 VNB N_VGND_c_3690_n 0.0292503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_218 VNB N_VGND_c_3691_n 0.00563307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_219 VNB N_VGND_c_3692_n 0.0639666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_220 VNB N_VGND_c_3693_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_221 VNB N_VGND_c_3694_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_222 VNB N_VGND_c_3695_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_223 VNB N_VGND_c_3696_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_224 VNB N_VGND_c_3697_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_225 VNB N_VGND_c_3698_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_226 VNB N_VGND_c_3699_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_227 VNB N_VGND_c_3700_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_228 VNB N_VGND_c_3701_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_229 VNB N_VGND_c_3702_n 0.018736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_230 VNB N_VGND_c_3703_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_231 VNB N_VGND_c_3704_n 0.0146622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_232 VNB N_VGND_c_3705_n 0.054046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_233 VNB N_VGND_c_3706_n 0.07403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_234 VNB N_VGND_c_3707_n 1.16202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_235 VNB N_VGND_c_3708_n 0.00885031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_236 VNB N_VGND_c_3709_n 0.0163055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_237 VNB N_VGND_c_3710_n 0.0138218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_238 VNB N_VGND_c_3711_n 0.00510127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_239 VNB N_VGND_c_3712_n 0.00596278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_240 VNB N_VGND_c_3713_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_241 VNB N_A_2519_47#_c_3956_n 0.00471053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_242 VNB N_A_2519_47#_c_3957_n 0.00134066f $X=-0.19 $Y=-0.245 $X2=1.065
+ $Y2=1.58
cc_243 VNB N_A_2519_47#_c_3958_n 0.00737026f $X=-0.19 $Y=-0.245 $X2=1.755
+ $Y2=1.25
cc_244 VNB N_A_2519_47#_c_3959_n 0.014863f $X=-0.19 $Y=-0.245 $X2=5.785
+ $Y2=2.675
cc_245 VPB N_SLEEP_M1026_g 0.0492776f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.595
cc_246 VPB N_SLEEP_M1006_g 0.0519351f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.775
cc_247 VPB N_SLEEP_M1049_g 0.0233442f $X=-0.19 $Y=1.655 $X2=5.785 $Y2=2.675
cc_248 VPB N_SLEEP_M1015_g 0.0191061f $X=-0.19 $Y=1.655 $X2=11.65 $Y2=2.465
cc_249 VPB N_SLEEP_M1046_g 0.0237126f $X=-0.19 $Y=1.655 $X2=12.08 $Y2=2.465
cc_250 VPB N_SLEEP_c_459_n 0.0458767f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=1.93
cc_251 VPB N_SLEEP_c_460_n 0.0148638f $X=-0.19 $Y=1.655 $X2=5.355 $Y2=2.035
cc_252 VPB N_SLEEP_c_461_n 0.017477f $X=-0.19 $Y=1.655 $X2=11.72 $Y2=2.035
cc_253 VPB N_SLEEP_c_462_n 0.0124693f $X=-0.19 $Y=1.655 $X2=5.51 $Y2=1.93
cc_254 VPB N_SLEEP_c_451_n 0.00544351f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=1.415
cc_255 VPB N_SLEEP_c_453_n 0.00872303f $X=-0.19 $Y=1.655 $X2=12.08 $Y2=1.475
cc_256 VPB N_TE_B_M1001_g 0.0436144f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_257 VPB N_TE_B_c_676_n 0.0463758f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.58
cc_258 VPB N_TE_B_c_677_n 0.00695714f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.595
cc_259 VPB N_TE_B_c_670_n 0.00938063f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_27_47#_M1036_g 0.01719f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=1.25
cc_261 VPB N_A_27_47#_M1066_g 0.0216352f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=1.58
cc_262 VPB N_A_27_47#_c_729_n 0.0112908f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.775
cc_263 VPB N_A_27_47#_c_730_n 0.00495812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_27_47#_c_731_n 0.00947783f $X=-0.19 $Y=1.655 $X2=5.785 $Y2=2.675
cc_265 VPB N_A_27_47#_c_738_n 0.00340299f $X=-0.19 $Y=1.655 $X2=5.785 $Y2=2.675
cc_266 VPB N_A_27_47#_c_732_n 0.0470004f $X=-0.19 $Y=1.655 $X2=11.65 $Y2=1.67
cc_267 VPB N_A_280_47#_M1035_g 0.0301355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_280_47#_c_828_n 0.0372888f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.775
cc_269 VPB N_A_280_47#_c_829_n 0.00983351f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=2.775
cc_270 VPB N_A_280_47#_c_830_n 0.0257422f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=1.25
cc_271 VPB N_A_280_47#_c_831_n 0.0198268f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=0.655
cc_272 VPB N_A_280_47#_c_832_n 0.0176315f $X=-0.19 $Y=1.655 $X2=5.785 $Y2=2.095
cc_273 VPB N_A_280_47#_c_819_n 0.0203276f $X=-0.19 $Y=1.655 $X2=11.65 $Y2=1.67
cc_274 VPB N_A_280_47#_M1057_g 0.0396008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_280_47#_c_826_n 0.00218237f $X=-0.19 $Y=1.655 $X2=5.645 $Y2=2.035
cc_276 VPB N_A_280_47#_c_836_n 0.0114219f $X=-0.19 $Y=1.655 $X2=5.5 $Y2=2.035
cc_277 VPB N_A_280_47#_c_837_n 0.0124518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_A_280_47#_c_838_n 2.16534e-19 $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.415
cc_279 VPB N_A_280_47#_c_839_n 8.45823e-19 $X=-0.19 $Y=1.655 $X2=1.065 $Y2=1.415
cc_280 VPB N_A_705_367#_c_1000_n 0.0186906f $X=-0.19 $Y=1.655 $X2=1.325
+ $Y2=0.655
cc_281 VPB N_A_705_367#_M1027_g 0.0340453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_A_705_367#_c_1042_n 0.0189328f $X=-0.19 $Y=1.655 $X2=1.755
+ $Y2=0.655
cc_283 VPB N_A_705_367#_c_1001_n 0.0049292f $X=-0.19 $Y=1.655 $X2=5.785
+ $Y2=2.095
cc_284 VPB N_A_705_367#_c_1002_n 0.00311208f $X=-0.19 $Y=1.655 $X2=5.785
+ $Y2=2.675
cc_285 VPB N_A_705_367#_c_1045_n 0.0155578f $X=-0.19 $Y=1.655 $X2=5.785
+ $Y2=2.675
cc_286 VPB N_A_705_367#_c_1003_n 0.00544413f $X=-0.19 $Y=1.655 $X2=11.65
+ $Y2=2.465
cc_287 VPB N_A_705_367#_c_1047_n 0.0155017f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_A_705_367#_c_1004_n 0.0049292f $X=-0.19 $Y=1.655 $X2=12.08
+ $Y2=2.465
cc_289 VPB N_A_705_367#_c_1049_n 0.0155111f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=1.93
cc_290 VPB N_A_705_367#_c_1005_n 0.00544413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_A_705_367#_c_1051_n 0.0155111f $X=-0.19 $Y=1.655 $X2=11.95
+ $Y2=1.445
cc_292 VPB N_A_705_367#_c_1006_n 0.0049292f $X=-0.19 $Y=1.655 $X2=5.355
+ $Y2=2.035
cc_293 VPB N_A_705_367#_c_1053_n 0.0155111f $X=-0.19 $Y=1.655 $X2=11.72
+ $Y2=2.035
cc_294 VPB N_A_705_367#_c_1007_n 0.00544413f $X=-0.19 $Y=1.655 $X2=5.5 $Y2=2.035
cc_295 VPB N_A_705_367#_c_1055_n 0.0155111f $X=-0.19 $Y=1.655 $X2=11.865
+ $Y2=2.035
cc_296 VPB N_A_705_367#_c_1008_n 0.0049292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_A_705_367#_c_1057_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_A_705_367#_c_1009_n 0.00544413f $X=-0.19 $Y=1.655 $X2=5.51 $Y2=1.93
cc_299 VPB N_A_705_367#_c_1059_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=1.415
cc_300 VPB N_A_705_367#_c_1010_n 0.0049292f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=1.415
cc_301 VPB N_A_705_367#_c_1061_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0.835
+ $Y2=1.415
cc_302 VPB N_A_705_367#_c_1011_n 0.00544413f $X=-0.19 $Y=1.655 $X2=1.755
+ $Y2=1.415
cc_303 VPB N_A_705_367#_c_1063_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_304 VPB N_A_705_367#_c_1012_n 0.0049292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_A_705_367#_c_1065_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_A_705_367#_c_1066_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.035
cc_307 VPB N_A_705_367#_c_1067_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_308 VPB N_A_705_367#_c_1068_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_309 VPB N_A_705_367#_c_1069_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_310 VPB N_A_705_367#_c_1070_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_311 VPB N_A_705_367#_c_1071_n 0.0155152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_312 VPB N_A_705_367#_c_1072_n 0.0157552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_313 VPB N_A_705_367#_c_1073_n 0.0220709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_314 VPB N_A_705_367#_c_1013_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_315 VPB N_A_705_367#_c_1014_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_316 VPB N_A_705_367#_c_1015_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_317 VPB N_A_705_367#_c_1016_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_318 VPB N_A_705_367#_c_1017_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_319 VPB N_A_705_367#_c_1018_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_320 VPB N_A_705_367#_c_1019_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_321 VPB N_A_705_367#_c_1020_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_322 VPB N_A_705_367#_c_1021_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_323 VPB N_A_705_367#_c_1022_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_324 VPB N_A_705_367#_c_1084_n 0.00170855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_325 VPB N_A_705_367#_c_1025_n 0.00470295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_326 VPB N_A_705_367#_c_1086_n 0.0127797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_327 VPB N_A_705_367#_c_1087_n 0.00209965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_328 VPB N_A_705_367#_c_1028_n 0.00189688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_329 VPB N_A_705_367#_c_1029_n 0.0331746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_330 VPB N_A_705_367#_c_1030_n 9.06975e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_331 VPB N_A_705_367#_c_1031_n 0.00144296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_332 VPB N_A_705_367#_c_1032_n 0.0163193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_333 VPB N_A_705_367#_c_1033_n 0.00408636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_334 VPB N_A_705_367#_c_1034_n 0.00187511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_335 VPB N_A_705_367#_c_1035_n 0.00187511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_336 VPB N_A_705_367#_c_1036_n 0.00187511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_337 VPB N_A_705_367#_c_1037_n 0.0534031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_338 VPB N_A_705_367#_c_1038_n 0.00353111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_339 VPB N_A_705_367#_c_1039_n 0.00179737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_340 VPB N_A_407_491#_M1018_g 0.0177917f $X=-0.19 $Y=1.655 $X2=1.755 $Y2=1.25
cc_341 VPB N_A_407_491#_c_1572_n 0.00710636f $X=-0.19 $Y=1.655 $X2=11.65
+ $Y2=2.465
cc_342 VPB N_A_407_491#_c_1573_n 0.00283629f $X=-0.19 $Y=1.655 $X2=12.08
+ $Y2=1.67
cc_343 VPB N_A_407_491#_c_1574_n 0.00308242f $X=-0.19 $Y=1.655 $X2=12.08
+ $Y2=2.465
cc_344 VPB N_A_407_491#_c_1562_n 6.98705e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_345 VPB N_A_896_367#_c_1764_n 0.0174351f $X=-0.19 $Y=1.655 $X2=0.835
+ $Y2=0.445
cc_346 VPB N_A_896_367#_c_1774_n 0.0192172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_347 VPB N_A_896_367#_c_1765_n 0.00700949f $X=-0.19 $Y=1.655 $X2=1.065
+ $Y2=2.775
cc_348 VPB N_A_896_367#_c_1776_n 0.0161951f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=1.25
cc_349 VPB N_A_896_367#_c_1766_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_350 VPB N_A_896_367#_c_1778_n 0.00655073f $X=-0.19 $Y=1.655 $X2=5.785
+ $Y2=2.095
cc_351 VPB N_A_896_367#_c_1779_n 0.0144931f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=1.93
cc_352 VPB N_A_896_367#_c_1771_n 0.00329303f $X=-0.19 $Y=1.655 $X2=11.95
+ $Y2=1.445
cc_353 VPB N_A_896_367#_c_1781_n 0.00133332f $X=-0.19 $Y=1.655 $X2=5.645
+ $Y2=2.035
cc_354 VPB N_A_896_367#_c_1772_n 0.0263723f $X=-0.19 $Y=1.655 $X2=11.865
+ $Y2=2.035
cc_355 VPB N_A_1486_47#_M1068_g 0.0178282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_356 VPB N_A_1486_47#_c_1942_n 0.0137652f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=2.035
cc_357 VPB N_A_1486_47#_c_1948_n 0.00194604f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_358 VPB N_A_c_2281_n 0.0166547f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.25
cc_359 VPB N_A_c_2282_n 0.0169487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_360 VPB N_A_c_2283_n 0.0754222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_361 VPB N_A_c_2284_n 0.110679f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=1.25
cc_362 VPB N_A_c_2285_n 0.00989679f $X=-0.19 $Y=1.655 $X2=1.325 $Y2=0.655
cc_363 VPB N_A_c_2286_n 0.085051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_364 VPB N_A_c_2267_n 0.0141786f $X=-0.19 $Y=1.655 $X2=5.785 $Y2=2.675
cc_365 VPB N_A_c_2268_n 0.00697368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_366 VPB N_A_c_2289_n 0.0219093f $X=-0.19 $Y=1.655 $X2=12.08 $Y2=1.67
cc_367 VPB N_A_c_2270_n 0.00544413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_368 VPB N_A_c_2291_n 0.0199545f $X=-0.19 $Y=1.655 $X2=11.95 $Y2=1.445
cc_369 VPB N_A_c_2272_n 0.0174916f $X=-0.19 $Y=1.655 $X2=5.645 $Y2=2.035
cc_370 VPB N_A_c_2274_n 0.00408568f $X=-0.19 $Y=1.655 $X2=5.5 $Y2=2.035
cc_371 VPB N_A_c_2278_n 0.00505188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_372 VPB N_A_c_2279_n 0.00349565f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_373 VPB N_A_2063_47#_c_2486_n 0.00250237f $X=-0.19 $Y=1.655 $X2=5.785
+ $Y2=2.675
cc_374 VPB N_A_2063_47#_c_2495_n 0.010598f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=1.93
cc_375 VPB N_A_2063_47#_c_2496_n 0.0065842f $X=-0.19 $Y=1.655 $X2=11.882
+ $Y2=1.615
cc_376 VPB N_VPWR_c_2628_n 0.00466824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_377 VPB N_VPWR_c_2629_n 0.00645436f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.415
cc_378 VPB N_VPWR_c_2630_n 0.0150479f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=1.415
cc_379 VPB N_VPWR_c_2631_n 0.002326f $X=-0.19 $Y=1.655 $X2=11.65 $Y2=1.475
cc_380 VPB N_VPWR_c_2632_n 0.021392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_381 VPB N_VPWR_c_2633_n 0.0138734f $X=-0.19 $Y=1.655 $X2=0.77 $Y2=2.035
cc_382 VPB N_VPWR_c_2634_n 0.0184034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_383 VPB N_VPWR_c_2635_n 0.00740105f $X=-0.19 $Y=1.655 $X2=11.882 $Y2=2.035
cc_384 VPB N_VPWR_c_2636_n 0.0110763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_385 VPB N_VPWR_c_2637_n 0.00229788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_386 VPB N_VPWR_c_2638_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_387 VPB N_VPWR_c_2639_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_388 VPB N_VPWR_c_2640_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_389 VPB N_VPWR_c_2641_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_390 VPB N_VPWR_c_2642_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_391 VPB N_VPWR_c_2643_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_392 VPB N_VPWR_c_2644_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_393 VPB N_VPWR_c_2645_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_394 VPB N_VPWR_c_2646_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_395 VPB N_VPWR_c_2647_n 0.0290284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_396 VPB N_VPWR_c_2648_n 0.0267309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_397 VPB N_VPWR_c_2649_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_398 VPB N_VPWR_c_2650_n 0.0131585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_399 VPB N_VPWR_c_2651_n 0.00356964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_400 VPB N_VPWR_c_2652_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_401 VPB N_VPWR_c_2653_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_402 VPB N_VPWR_c_2654_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_403 VPB N_VPWR_c_2655_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_404 VPB N_VPWR_c_2656_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_405 VPB N_VPWR_c_2657_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_406 VPB N_VPWR_c_2658_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_407 VPB N_VPWR_c_2659_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_408 VPB N_VPWR_c_2660_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_409 VPB N_VPWR_c_2661_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_410 VPB N_VPWR_c_2662_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_411 VPB N_VPWR_c_2663_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_412 VPB N_VPWR_c_2664_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_413 VPB N_VPWR_c_2665_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_414 VPB N_VPWR_c_2666_n 0.0178246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_415 VPB N_VPWR_c_2667_n 0.117603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_416 VPB N_VPWR_c_2668_n 0.0477806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_417 VPB N_VPWR_c_2669_n 0.0167833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_418 VPB N_VPWR_c_2670_n 0.0364808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_419 VPB N_VPWR_c_2671_n 0.0382621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_420 VPB N_VPWR_c_2672_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_421 VPB N_VPWR_c_2673_n 0.0199636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_422 VPB N_VPWR_c_2627_n 0.0625959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_423 VPB N_VPWR_c_2675_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_424 VPB N_VPWR_c_2676_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_425 VPB N_VPWR_c_2677_n 0.00376198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_426 VPB N_VPWR_c_2678_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_427 VPB N_VPWR_c_2679_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_428 VPB N_VPWR_c_2680_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_429 VPB N_VPWR_c_2681_n 0.00520459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_430 VPB N_VPWR_c_2682_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_431 VPB N_VPWR_c_2683_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_432 VPB KAPWR 0.0804176f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.445
cc_433 VPB N_KAPWR_c_3047_n 0.00376924f $X=-0.19 $Y=1.655 $X2=1.755 $Y2=1.25
cc_434 VPB N_KAPWR_c_3048_n 0.00278483f $X=-0.19 $Y=1.655 $X2=12.08 $Y2=1.67
cc_435 VPB N_A_1492_367#_c_3237_n 9.03475e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_436 VPB N_A_1492_367#_c_3238_n 0.00334613f $X=-0.19 $Y=1.655 $X2=1.325
+ $Y2=0.655
cc_437 VPB N_A_1492_367#_c_3239_n 0.00625053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_438 VPB N_A_2345_367#_c_3306_n 0.00546202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_439 VPB N_A_2345_367#_c_3307_n 0.00271861f $X=-0.19 $Y=1.655 $X2=1.065
+ $Y2=2.775
cc_440 VPB N_A_2345_367#_c_3308_n 0.00301578f $X=-0.19 $Y=1.655 $X2=1.065
+ $Y2=2.775
cc_441 VPB N_A_2345_367#_c_3309_n 0.00236122f $X=-0.19 $Y=1.655 $X2=1.325
+ $Y2=1.25
cc_442 VPB N_A_2345_367#_c_3310_n 0.00233756f $X=-0.19 $Y=1.655 $X2=1.325
+ $Y2=0.655
cc_443 VPB N_A_2345_367#_c_3311_n 0.00513326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_444 N_SLEEP_c_460_n N_TE_B_M1001_g 0.00373287f $X=5.355 $Y=2.035 $X2=0 $Y2=0
cc_445 N_SLEEP_c_460_n N_TE_B_c_676_n 0.00702438f $X=5.355 $Y=2.035 $X2=0 $Y2=0
cc_446 N_SLEEP_M1006_g N_TE_B_c_677_n 0.0912569f $X=1.065 $Y=2.775 $X2=0 $Y2=0
cc_447 N_SLEEP_c_452_n N_TE_B_c_677_n 0.0324572f $X=1.325 $Y=1.415 $X2=0 $Y2=0
cc_448 N_SLEEP_M1045_g N_TE_B_M1008_g 0.0316992f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_449 N_SLEEP_M1045_g TE_B 0.00347561f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_450 N_SLEEP_M1045_g N_TE_B_c_674_n 0.019512f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_451 N_SLEEP_c_460_n N_A_27_47#_M1036_g 0.00455628f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_452 N_SLEEP_c_459_n N_A_27_47#_M1066_g 0.00820478f $X=5.71 $Y=1.93 $X2=0
+ $Y2=0
cc_453 N_SLEEP_c_460_n N_A_27_47#_M1066_g 0.00871295f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_454 N_SLEEP_c_462_n N_A_27_47#_M1066_g 0.00586016f $X=5.51 $Y=1.93 $X2=0
+ $Y2=0
cc_455 N_SLEEP_M1026_g N_A_27_47#_c_729_n 0.0141342f $X=0.525 $Y=2.595 $X2=0
+ $Y2=0
cc_456 N_SLEEP_M1006_g N_A_27_47#_c_729_n 0.00749461f $X=1.065 $Y=2.775 $X2=0
+ $Y2=0
cc_457 N_SLEEP_c_460_n N_A_27_47#_c_729_n 0.280506f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_458 N_SLEEP_c_479_p N_A_27_47#_c_729_n 0.0229319f $X=0.915 $Y=2.035 $X2=0
+ $Y2=0
cc_459 N_SLEEP_c_451_n N_A_27_47#_c_729_n 0.0271297f $X=0.76 $Y=1.415 $X2=0
+ $Y2=0
cc_460 N_SLEEP_c_452_n N_A_27_47#_c_729_n 0.0104103f $X=1.325 $Y=1.415 $X2=0
+ $Y2=0
cc_461 N_SLEEP_c_451_n N_A_27_47#_c_730_n 5.97957e-19 $X=0.76 $Y=1.415 $X2=0
+ $Y2=0
cc_462 N_SLEEP_c_460_n N_A_27_47#_c_751_n 0.0254252f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_463 N_SLEEP_c_460_n N_A_27_47#_c_738_n 0.0035121f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_464 N_SLEEP_c_462_n N_A_27_47#_c_738_n 0.00180558f $X=5.51 $Y=1.93 $X2=0
+ $Y2=0
cc_465 N_SLEEP_M1030_g N_A_27_47#_c_732_n 0.0296029f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_466 N_SLEEP_M1026_g N_A_27_47#_c_732_n 0.0390841f $X=0.525 $Y=2.595 $X2=0
+ $Y2=0
cc_467 N_SLEEP_M1002_g N_A_27_47#_c_732_n 0.00309257f $X=0.835 $Y=0.445 $X2=0
+ $Y2=0
cc_468 N_SLEEP_M1006_g N_A_27_47#_c_732_n 0.00106881f $X=1.065 $Y=2.775 $X2=0
+ $Y2=0
cc_469 N_SLEEP_c_479_p N_A_27_47#_c_732_n 0.00153655f $X=0.915 $Y=2.035 $X2=0
+ $Y2=0
cc_470 N_SLEEP_c_451_n N_A_27_47#_c_732_n 0.067899f $X=0.76 $Y=1.415 $X2=0 $Y2=0
cc_471 N_SLEEP_c_452_n N_A_27_47#_c_732_n 0.0120573f $X=1.325 $Y=1.415 $X2=0
+ $Y2=0
cc_472 N_SLEEP_c_460_n N_A_280_47#_c_830_n 0.00469684f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_473 N_SLEEP_c_460_n N_A_280_47#_c_831_n 0.00189154f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_474 N_SLEEP_c_460_n N_A_280_47#_c_832_n 0.00402676f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_475 N_SLEEP_c_460_n N_A_280_47#_c_819_n 9.68465e-19 $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_476 N_SLEEP_c_459_n N_A_280_47#_c_822_n 0.0324665f $X=5.71 $Y=1.93 $X2=0
+ $Y2=0
cc_477 N_SLEEP_c_461_n N_A_280_47#_c_822_n 7.05058e-19 $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_478 N_SLEEP_c_462_n N_A_280_47#_c_822_n 0.00305752f $X=5.51 $Y=1.93 $X2=0
+ $Y2=0
cc_479 N_SLEEP_c_460_n N_A_280_47#_c_823_n 0.00385139f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_480 N_SLEEP_c_459_n N_A_280_47#_M1057_g 0.0948103f $X=5.71 $Y=1.93 $X2=0
+ $Y2=0
cc_481 N_SLEEP_c_461_n N_A_280_47#_M1057_g 0.00460927f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_482 N_SLEEP_c_462_n N_A_280_47#_M1057_g 0.00163219f $X=5.51 $Y=1.93 $X2=0
+ $Y2=0
cc_483 N_SLEEP_M1013_g N_A_280_47#_c_826_n 0.00382499f $X=1.325 $Y=0.655 $X2=0
+ $Y2=0
cc_484 N_SLEEP_M1045_g N_A_280_47#_c_826_n 0.00359111f $X=1.755 $Y=0.655 $X2=0
+ $Y2=0
cc_485 N_SLEEP_c_451_n N_A_280_47#_c_826_n 0.0166463f $X=0.76 $Y=1.415 $X2=0
+ $Y2=0
cc_486 N_SLEEP_c_452_n N_A_280_47#_c_826_n 0.0264005f $X=1.325 $Y=1.415 $X2=0
+ $Y2=0
cc_487 N_SLEEP_M1006_g N_A_280_47#_c_836_n 0.003865f $X=1.065 $Y=2.775 $X2=0
+ $Y2=0
cc_488 N_SLEEP_c_460_n N_A_280_47#_c_836_n 0.0295656f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_489 N_SLEEP_c_479_p N_A_280_47#_c_836_n 2.86441e-19 $X=0.915 $Y=2.035 $X2=0
+ $Y2=0
cc_490 N_SLEEP_c_451_n N_A_280_47#_c_836_n 0.00411286f $X=0.76 $Y=1.415 $X2=0
+ $Y2=0
cc_491 N_SLEEP_M1045_g N_A_280_47#_c_859_n 0.0110272f $X=1.755 $Y=0.655 $X2=0
+ $Y2=0
cc_492 N_SLEEP_c_460_n N_A_280_47#_c_837_n 0.015554f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_493 N_SLEEP_c_452_n N_A_280_47#_c_837_n 4.98767e-19 $X=1.325 $Y=1.415 $X2=0
+ $Y2=0
cc_494 N_SLEEP_M1006_g N_A_280_47#_c_839_n 9.88631e-19 $X=1.065 $Y=2.775 $X2=0
+ $Y2=0
cc_495 N_SLEEP_c_460_n N_A_280_47#_c_839_n 0.00195787f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_496 N_SLEEP_c_451_n N_A_280_47#_c_839_n 0.00638111f $X=0.76 $Y=1.415 $X2=0
+ $Y2=0
cc_497 N_SLEEP_c_452_n N_A_280_47#_c_839_n 0.00492897f $X=1.325 $Y=1.415 $X2=0
+ $Y2=0
cc_498 N_SLEEP_c_460_n N_A_705_367#_M1011_s 0.00349198f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_499 N_SLEEP_c_461_n N_A_705_367#_c_1000_n 0.00329157f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_500 N_SLEEP_c_461_n N_A_705_367#_M1027_g 0.00408112f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_501 N_SLEEP_c_460_n N_A_705_367#_c_1084_n 0.0173967f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_502 N_SLEEP_c_462_n N_A_705_367#_c_1023_n 0.011136f $X=5.51 $Y=1.93 $X2=0
+ $Y2=0
cc_503 N_SLEEP_c_459_n N_A_705_367#_c_1025_n 2.45819e-19 $X=5.71 $Y=1.93 $X2=0
+ $Y2=0
cc_504 N_SLEEP_c_461_n N_A_705_367#_c_1025_n 0.00542024f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_505 N_SLEEP_M1015_g N_A_705_367#_c_1029_n 0.00189407f $X=11.65 $Y=2.465 $X2=0
+ $Y2=0
cc_506 N_SLEEP_M1046_g N_A_705_367#_c_1029_n 0.00189569f $X=12.08 $Y=2.465 $X2=0
+ $Y2=0
cc_507 N_SLEEP_c_450_n N_A_705_367#_c_1029_n 0.0179922f $X=11.95 $Y=1.445 $X2=0
+ $Y2=0
cc_508 N_SLEEP_c_461_n N_A_705_367#_c_1029_n 0.398654f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_509 N_SLEEP_c_530_p N_A_705_367#_c_1029_n 0.0229319f $X=11.865 $Y=2.035 $X2=0
+ $Y2=0
cc_510 N_SLEEP_c_531_p N_A_705_367#_c_1029_n 0.0157109f $X=11.865 $Y=2.035 $X2=0
+ $Y2=0
cc_511 N_SLEEP_c_453_n N_A_705_367#_c_1029_n 0.00225159f $X=12.08 $Y=1.475 $X2=0
+ $Y2=0
cc_512 N_SLEEP_c_461_n N_A_705_367#_c_1030_n 0.0253772f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_513 N_SLEEP_c_461_n N_A_705_367#_c_1033_n 0.00338067f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_514 N_SLEEP_c_462_n N_A_705_367#_c_1033_n 0.00389486f $X=5.51 $Y=1.93 $X2=0
+ $Y2=0
cc_515 N_SLEEP_c_461_n N_A_705_367#_c_1039_n 0.00838423f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_516 N_SLEEP_c_461_n N_A_407_491#_M1018_g 0.0044577f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_517 N_SLEEP_c_460_n N_A_407_491#_c_1573_n 0.034048f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_518 N_SLEEP_c_460_n N_A_407_491#_c_1574_n 0.0127257f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_519 N_SLEEP_c_460_n N_A_407_491#_c_1562_n 0.0120229f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_520 N_SLEEP_c_460_n N_A_896_367#_M1036_s 0.00161074f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_521 N_SLEEP_c_461_n N_A_896_367#_c_1764_n 0.00102701f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_522 N_SLEEP_c_461_n N_A_896_367#_c_1774_n 0.00330179f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_523 N_SLEEP_c_461_n N_A_896_367#_c_1776_n 0.00340098f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_524 N_SLEEP_M1049_g N_A_896_367#_c_1778_n 0.0126492f $X=5.785 $Y=2.675 $X2=0
+ $Y2=0
cc_525 N_SLEEP_c_459_n N_A_896_367#_c_1778_n 0.00192973f $X=5.71 $Y=1.93 $X2=0
+ $Y2=0
cc_526 N_SLEEP_c_460_n N_A_896_367#_c_1778_n 0.0148849f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_527 N_SLEEP_c_461_n N_A_896_367#_c_1778_n 0.00978701f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_528 N_SLEEP_c_549_p N_A_896_367#_c_1778_n 0.00129072f $X=5.645 $Y=2.035 $X2=0
+ $Y2=0
cc_529 N_SLEEP_c_462_n N_A_896_367#_c_1778_n 0.0277452f $X=5.51 $Y=1.93 $X2=0
+ $Y2=0
cc_530 N_SLEEP_c_461_n N_A_896_367#_c_1779_n 0.0235519f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_531 N_SLEEP_c_461_n N_A_896_367#_c_1771_n 0.0146753f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_532 N_SLEEP_c_460_n N_A_896_367#_c_1795_n 0.0117722f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_533 N_SLEEP_c_462_n N_A_896_367#_c_1795_n 0.00154713f $X=5.51 $Y=1.93 $X2=0
+ $Y2=0
cc_534 N_SLEEP_M1049_g N_A_896_367#_c_1781_n 0.00215566f $X=5.785 $Y=2.675 $X2=0
+ $Y2=0
cc_535 N_SLEEP_c_459_n N_A_896_367#_c_1781_n 0.00107774f $X=5.71 $Y=1.93 $X2=0
+ $Y2=0
cc_536 N_SLEEP_c_461_n N_A_896_367#_c_1781_n 0.0142665f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_537 N_SLEEP_c_462_n N_A_896_367#_c_1781_n 0.00163075f $X=5.51 $Y=1.93 $X2=0
+ $Y2=0
cc_538 N_SLEEP_c_461_n N_A_896_367#_c_1772_n 0.00121015f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_539 N_SLEEP_c_461_n N_A_1486_47#_M1023_d 0.00199463f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_540 N_SLEEP_c_461_n N_A_1486_47#_M1068_g 0.00439161f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_541 N_SLEEP_c_461_n N_A_1486_47#_c_1948_n 0.0155505f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_542 N_SLEEP_c_450_n N_A_1486_47#_c_1953_n 0.0185924f $X=11.95 $Y=1.445 $X2=0
+ $Y2=0
cc_543 N_SLEEP_c_531_p N_A_1486_47#_c_1953_n 2.05202e-19 $X=11.865 $Y=2.035
+ $X2=0 $Y2=0
cc_544 N_SLEEP_c_453_n N_A_1486_47#_c_1953_n 0.00231107f $X=12.08 $Y=1.475 $X2=0
+ $Y2=0
cc_545 N_SLEEP_c_461_n N_A_1486_47#_c_1958_n 8.46721e-19 $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_546 N_SLEEP_c_461_n N_A_c_2281_n 0.00373978f $X=11.72 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_547 N_SLEEP_c_461_n N_A_c_2282_n 0.00640605f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_548 N_SLEEP_c_461_n N_A_c_2283_n 0.00702949f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_549 N_SLEEP_M1015_g N_A_c_2286_n 0.0373753f $X=11.65 $Y=2.465 $X2=0 $Y2=0
cc_550 N_SLEEP_c_461_n N_A_c_2286_n 0.00572249f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_551 N_SLEEP_c_531_p N_A_c_2286_n 0.00172656f $X=11.865 $Y=2.035 $X2=0 $Y2=0
cc_552 N_SLEEP_c_450_n N_A_c_2266_n 3.06978e-19 $X=11.95 $Y=1.445 $X2=0 $Y2=0
cc_553 N_SLEEP_c_453_n N_A_c_2266_n 0.0150763f $X=12.08 $Y=1.475 $X2=0 $Y2=0
cc_554 N_SLEEP_M1046_g N_A_c_2268_n 0.0150763f $X=12.08 $Y=2.465 $X2=0 $Y2=0
cc_555 N_SLEEP_c_531_p N_A_c_2268_n 0.00101617f $X=11.865 $Y=2.035 $X2=0 $Y2=0
cc_556 N_SLEEP_c_461_n N_A_c_2272_n 0.00140223f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_557 N_SLEEP_c_450_n N_A_c_2273_n 9.71842e-19 $X=11.95 $Y=1.445 $X2=0 $Y2=0
cc_558 N_SLEEP_c_453_n N_A_c_2273_n 0.0248695f $X=12.08 $Y=1.475 $X2=0 $Y2=0
cc_559 N_SLEEP_M1015_g N_A_c_2274_n 0.00221245f $X=11.65 $Y=2.465 $X2=0 $Y2=0
cc_560 N_SLEEP_c_531_p N_A_c_2274_n 3.13669e-19 $X=11.865 $Y=2.035 $X2=0 $Y2=0
cc_561 N_SLEEP_c_453_n N_A_c_2275_n 0.0256294f $X=12.08 $Y=1.475 $X2=0 $Y2=0
cc_562 N_SLEEP_M1015_g N_A_2063_47#_c_2486_n 5.83242e-19 $X=11.65 $Y=2.465 $X2=0
+ $Y2=0
cc_563 N_SLEEP_c_450_n N_A_2063_47#_c_2486_n 0.0128537f $X=11.95 $Y=1.445 $X2=0
+ $Y2=0
cc_564 N_SLEEP_c_531_p N_A_2063_47#_c_2486_n 0.0043544f $X=11.865 $Y=2.035 $X2=0
+ $Y2=0
cc_565 N_SLEEP_c_453_n N_A_2063_47#_c_2486_n 9.95471e-19 $X=12.08 $Y=1.475 $X2=0
+ $Y2=0
cc_566 N_SLEEP_c_450_n N_A_2063_47#_c_2487_n 0.0357796f $X=11.95 $Y=1.445 $X2=0
+ $Y2=0
cc_567 N_SLEEP_c_453_n N_A_2063_47#_c_2487_n 0.00529345f $X=12.08 $Y=1.475 $X2=0
+ $Y2=0
cc_568 N_SLEEP_c_450_n N_A_2063_47#_c_2489_n 0.023939f $X=11.95 $Y=1.445 $X2=0
+ $Y2=0
cc_569 N_SLEEP_c_453_n N_A_2063_47#_c_2489_n 0.00285261f $X=12.08 $Y=1.475 $X2=0
+ $Y2=0
cc_570 N_SLEEP_c_461_n N_A_2063_47#_c_2495_n 0.0190762f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_571 N_SLEEP_M1015_g N_A_2063_47#_c_2496_n 5.77226e-19 $X=11.65 $Y=2.465 $X2=0
+ $Y2=0
cc_572 N_SLEEP_c_461_n N_A_2063_47#_c_2496_n 0.0200864f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_573 N_SLEEP_c_531_p N_A_2063_47#_c_2496_n 0.00363366f $X=11.865 $Y=2.035
+ $X2=0 $Y2=0
cc_574 N_SLEEP_c_479_p N_VPWR_M1026_d 0.00145735f $X=0.915 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_575 N_SLEEP_c_451_n N_VPWR_M1026_d 0.00123652f $X=0.76 $Y=1.415 $X2=-0.19
+ $Y2=-0.245
cc_576 N_SLEEP_c_461_n N_VPWR_M1012_s 0.00450916f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_577 N_SLEEP_c_461_n N_VPWR_M1015_d 0.00427268f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_578 N_SLEEP_M1026_g N_VPWR_c_2628_n 0.0183708f $X=0.525 $Y=2.595 $X2=0 $Y2=0
cc_579 N_SLEEP_M1006_g N_VPWR_c_2628_n 0.00909072f $X=1.065 $Y=2.775 $X2=0 $Y2=0
cc_580 N_SLEEP_c_460_n N_VPWR_c_2628_n 0.0011617f $X=5.355 $Y=2.035 $X2=0 $Y2=0
cc_581 N_SLEEP_c_479_p N_VPWR_c_2628_n 0.00154633f $X=0.915 $Y=2.035 $X2=0 $Y2=0
cc_582 N_SLEEP_c_451_n N_VPWR_c_2628_n 0.0184682f $X=0.76 $Y=1.415 $X2=0 $Y2=0
cc_583 N_SLEEP_M1049_g N_VPWR_c_2629_n 0.0134474f $X=5.785 $Y=2.675 $X2=0 $Y2=0
cc_584 N_SLEEP_c_461_n N_VPWR_c_2630_n 0.00101414f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_585 N_SLEEP_c_461_n N_VPWR_c_2632_n 0.0282924f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_586 N_SLEEP_M1015_g N_VPWR_c_2633_n 0.00215291f $X=11.65 $Y=2.465 $X2=0 $Y2=0
cc_587 N_SLEEP_c_461_n N_VPWR_c_2633_n 0.00960853f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_588 N_SLEEP_c_453_n N_VPWR_c_2633_n 0.00162231f $X=12.08 $Y=1.475 $X2=0 $Y2=0
cc_589 N_SLEEP_M1015_g N_VPWR_c_2634_n 0.00550269f $X=11.65 $Y=2.465 $X2=0 $Y2=0
cc_590 N_SLEEP_M1046_g N_VPWR_c_2634_n 0.00550269f $X=12.08 $Y=2.465 $X2=0 $Y2=0
cc_591 N_SLEEP_M1046_g N_VPWR_c_2635_n 0.00353971f $X=12.08 $Y=2.465 $X2=0 $Y2=0
cc_592 N_SLEEP_M1049_g N_VPWR_c_2648_n 0.00486043f $X=5.785 $Y=2.675 $X2=0 $Y2=0
cc_593 N_SLEEP_M1026_g N_VPWR_c_2666_n 0.00839865f $X=0.525 $Y=2.595 $X2=0 $Y2=0
cc_594 N_SLEEP_M1006_g N_VPWR_c_2667_n 0.00585385f $X=1.065 $Y=2.775 $X2=0 $Y2=0
cc_595 N_SLEEP_M1026_g N_VPWR_c_2627_n 0.00688923f $X=0.525 $Y=2.595 $X2=0 $Y2=0
cc_596 N_SLEEP_M1006_g N_VPWR_c_2627_n 0.00520998f $X=1.065 $Y=2.775 $X2=0 $Y2=0
cc_597 N_SLEEP_M1049_g N_VPWR_c_2627_n 0.00328821f $X=5.785 $Y=2.675 $X2=0 $Y2=0
cc_598 N_SLEEP_M1015_g N_VPWR_c_2627_n 0.00522432f $X=11.65 $Y=2.465 $X2=0 $Y2=0
cc_599 N_SLEEP_M1046_g N_VPWR_c_2627_n 0.00610887f $X=12.08 $Y=2.465 $X2=0 $Y2=0
cc_600 N_SLEEP_c_460_n N_KAPWR_M1035_d 0.00158481f $X=5.355 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_601 N_SLEEP_c_460_n N_KAPWR_M1042_d 6.17359e-19 $X=5.355 $Y=2.035 $X2=0 $Y2=0
cc_602 N_SLEEP_c_460_n N_KAPWR_M1066_d 0.0113862f $X=5.355 $Y=2.035 $X2=0 $Y2=0
cc_603 N_SLEEP_M1026_g KAPWR 0.00915521f $X=0.525 $Y=2.595 $X2=0 $Y2=0
cc_604 N_SLEEP_M1006_g KAPWR 0.00777058f $X=1.065 $Y=2.775 $X2=0 $Y2=0
cc_605 N_SLEEP_M1049_g KAPWR 0.00358348f $X=5.785 $Y=2.675 $X2=0 $Y2=0
cc_606 N_SLEEP_M1015_g KAPWR 0.00306098f $X=11.65 $Y=2.465 $X2=0 $Y2=0
cc_607 N_SLEEP_M1046_g KAPWR 0.00243668f $X=12.08 $Y=2.465 $X2=0 $Y2=0
cc_608 N_SLEEP_c_460_n KAPWR 0.189338f $X=5.355 $Y=2.035 $X2=0 $Y2=0
cc_609 N_SLEEP_c_479_p KAPWR 0.0120637f $X=0.915 $Y=2.035 $X2=0 $Y2=0
cc_610 N_SLEEP_c_461_n KAPWR 0.268169f $X=11.72 $Y=2.035 $X2=0 $Y2=0
cc_611 N_SLEEP_c_549_p KAPWR 0.0123087f $X=5.645 $Y=2.035 $X2=0 $Y2=0
cc_612 N_SLEEP_c_530_p KAPWR 0.0120593f $X=11.865 $Y=2.035 $X2=0 $Y2=0
cc_613 N_SLEEP_c_531_p KAPWR 3.65254e-19 $X=11.865 $Y=2.035 $X2=0 $Y2=0
cc_614 N_SLEEP_c_451_n KAPWR 0.00118658f $X=0.76 $Y=1.415 $X2=0 $Y2=0
cc_615 N_SLEEP_c_460_n N_KAPWR_c_3047_n 0.00348194f $X=5.355 $Y=2.035 $X2=0
+ $Y2=0
cc_616 N_SLEEP_c_460_n N_KAPWR_c_3065_n 0.0205206f $X=5.355 $Y=2.035 $X2=0 $Y2=0
cc_617 N_SLEEP_c_461_n N_A_1492_367#_M1023_s 9.10393e-19 $X=11.72 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_618 N_SLEEP_c_461_n N_A_1492_367#_M1044_d 0.00416605f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_619 N_SLEEP_c_461_n N_A_1492_367#_c_3237_n 0.0186583f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_620 N_SLEEP_c_461_n N_A_1492_367#_c_3238_n 0.0256034f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_621 N_SLEEP_c_461_n N_A_1492_367#_c_3244_n 0.0168032f $X=11.72 $Y=2.035 $X2=0
+ $Y2=0
cc_622 N_SLEEP_c_461_n N_A_1492_367#_c_3239_n 0.00968301f $X=11.72 $Y=2.035
+ $X2=0 $Y2=0
cc_623 N_SLEEP_c_461_n A_2033_373# 0.00482195f $X=11.72 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_624 N_SLEEP_c_530_p N_A_2345_367#_M1015_s 0.00116308f $X=11.865 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_625 N_SLEEP_c_531_p N_A_2345_367#_M1015_s 7.79861e-19 $X=11.865 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_626 N_SLEEP_M1046_g N_A_2345_367#_c_3306_n 0.010696f $X=12.08 $Y=2.465 $X2=0
+ $Y2=0
cc_627 N_SLEEP_c_531_p N_A_2345_367#_c_3306_n 0.00165595f $X=11.865 $Y=2.035
+ $X2=0 $Y2=0
cc_628 N_SLEEP_M1046_g N_A_2345_367#_c_3307_n 0.00356744f $X=12.08 $Y=2.465
+ $X2=0 $Y2=0
cc_629 N_SLEEP_M1046_g N_A_2345_367#_c_3308_n 0.00346098f $X=12.08 $Y=2.465
+ $X2=0 $Y2=0
cc_630 N_SLEEP_M1015_g N_A_2345_367#_c_3318_n 0.00726395f $X=11.65 $Y=2.465
+ $X2=0 $Y2=0
cc_631 N_SLEEP_M1046_g N_A_2345_367#_c_3318_n 0.008392f $X=12.08 $Y=2.465 $X2=0
+ $Y2=0
cc_632 N_SLEEP_c_461_n N_A_2345_367#_c_3318_n 3.93675e-19 $X=11.72 $Y=2.035
+ $X2=0 $Y2=0
cc_633 N_SLEEP_c_530_p N_A_2345_367#_c_3318_n 0.00156246f $X=11.865 $Y=2.035
+ $X2=0 $Y2=0
cc_634 N_SLEEP_c_531_p N_A_2345_367#_c_3318_n 0.0170035f $X=11.865 $Y=2.035
+ $X2=0 $Y2=0
cc_635 N_SLEEP_c_453_n N_A_2345_367#_c_3318_n 3.05781e-19 $X=12.08 $Y=1.475
+ $X2=0 $Y2=0
cc_636 N_SLEEP_M1002_g N_VGND_c_3664_n 0.0103132f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_637 N_SLEEP_M1013_g N_VGND_c_3664_n 0.00228538f $X=1.325 $Y=0.655 $X2=0 $Y2=0
cc_638 N_SLEEP_c_452_n N_VGND_c_3664_n 0.00718274f $X=1.325 $Y=1.415 $X2=0 $Y2=0
cc_639 N_SLEEP_M1013_g N_VGND_c_3665_n 5.83176e-19 $X=1.325 $Y=0.655 $X2=0 $Y2=0
cc_640 N_SLEEP_M1045_g N_VGND_c_3665_n 0.00986287f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_641 N_SLEEP_M1030_g N_VGND_c_3680_n 0.0054895f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_642 N_SLEEP_M1002_g N_VGND_c_3680_n 0.00585385f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_643 N_SLEEP_M1013_g N_VGND_c_3682_n 0.00583607f $X=1.325 $Y=0.655 $X2=0 $Y2=0
cc_644 N_SLEEP_M1045_g N_VGND_c_3682_n 0.00486043f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_645 N_SLEEP_M1030_g N_VGND_c_3707_n 0.0107425f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_646 N_SLEEP_M1002_g N_VGND_c_3707_n 0.0107545f $X=0.835 $Y=0.445 $X2=0 $Y2=0
cc_647 N_SLEEP_M1013_g N_VGND_c_3707_n 0.0106359f $X=1.325 $Y=0.655 $X2=0 $Y2=0
cc_648 N_SLEEP_M1045_g N_VGND_c_3707_n 0.00458264f $X=1.755 $Y=0.655 $X2=0 $Y2=0
cc_649 N_TE_B_c_677_n N_A_27_47#_c_729_n 3.66409e-19 $X=1.5 $Y=1.86 $X2=0 $Y2=0
cc_650 N_TE_B_c_670_n N_A_27_47#_c_729_n 0.0065473f $X=2.155 $Y=1.785 $X2=0
+ $Y2=0
cc_651 TE_B N_A_27_47#_c_729_n 0.0111613f $X=2.15 $Y=1.21 $X2=0 $Y2=0
cc_652 N_TE_B_c_674_n N_A_27_47#_c_729_n 0.00527645f $X=2.615 $Y=1.395 $X2=0
+ $Y2=0
cc_653 N_TE_B_c_674_n N_A_280_47#_c_829_n 0.00610561f $X=2.615 $Y=1.395 $X2=0
+ $Y2=0
cc_654 N_TE_B_c_676_n N_A_280_47#_c_830_n 0.00243495f $X=2.08 $Y=1.86 $X2=0
+ $Y2=0
cc_655 N_TE_B_c_670_n N_A_280_47#_c_819_n 0.00243495f $X=2.155 $Y=1.785 $X2=0
+ $Y2=0
cc_656 TE_B N_A_280_47#_c_819_n 0.00110141f $X=2.15 $Y=1.21 $X2=0 $Y2=0
cc_657 N_TE_B_c_674_n N_A_280_47#_c_819_n 0.024292f $X=2.615 $Y=1.395 $X2=0
+ $Y2=0
cc_658 N_TE_B_c_670_n N_A_280_47#_c_826_n 0.00308784f $X=2.155 $Y=1.785 $X2=0
+ $Y2=0
cc_659 TE_B N_A_280_47#_c_826_n 0.0159345f $X=2.15 $Y=1.21 $X2=0 $Y2=0
cc_660 N_TE_B_c_674_n N_A_280_47#_c_826_n 3.74055e-19 $X=2.615 $Y=1.395 $X2=0
+ $Y2=0
cc_661 N_TE_B_M1001_g N_A_280_47#_c_836_n 0.0281702f $X=1.425 $Y=2.775 $X2=0
+ $Y2=0
cc_662 N_TE_B_c_676_n N_A_280_47#_c_836_n 0.00741343f $X=2.08 $Y=1.86 $X2=0
+ $Y2=0
cc_663 N_TE_B_M1008_g N_A_280_47#_c_859_n 0.00972748f $X=2.185 $Y=0.655 $X2=0
+ $Y2=0
cc_664 N_TE_B_M1040_g N_A_280_47#_c_859_n 0.00187695f $X=2.615 $Y=0.655 $X2=0
+ $Y2=0
cc_665 TE_B N_A_280_47#_c_859_n 0.0251279f $X=2.15 $Y=1.21 $X2=0 $Y2=0
cc_666 N_TE_B_c_674_n N_A_280_47#_c_859_n 0.00211324f $X=2.615 $Y=1.395 $X2=0
+ $Y2=0
cc_667 N_TE_B_c_676_n N_A_280_47#_c_837_n 0.0156717f $X=2.08 $Y=1.86 $X2=0 $Y2=0
cc_668 N_TE_B_c_670_n N_A_280_47#_c_837_n 0.00327152f $X=2.155 $Y=1.785 $X2=0
+ $Y2=0
cc_669 TE_B N_A_280_47#_c_837_n 0.0227594f $X=2.15 $Y=1.21 $X2=0 $Y2=0
cc_670 N_TE_B_c_674_n N_A_280_47#_c_837_n 0.00799004f $X=2.615 $Y=1.395 $X2=0
+ $Y2=0
cc_671 N_TE_B_M1040_g N_A_280_47#_c_884_n 0.00611044f $X=2.615 $Y=0.655 $X2=0
+ $Y2=0
cc_672 N_TE_B_c_670_n N_A_280_47#_c_838_n 9.19395e-19 $X=2.155 $Y=1.785 $X2=0
+ $Y2=0
cc_673 TE_B N_A_280_47#_c_838_n 0.00780662f $X=2.15 $Y=1.21 $X2=0 $Y2=0
cc_674 N_TE_B_c_674_n N_A_280_47#_c_838_n 0.00110519f $X=2.615 $Y=1.395 $X2=0
+ $Y2=0
cc_675 N_TE_B_c_676_n N_A_280_47#_c_839_n 0.00561654f $X=2.08 $Y=1.86 $X2=0
+ $Y2=0
cc_676 N_TE_B_c_677_n N_A_280_47#_c_839_n 0.0046026f $X=1.5 $Y=1.86 $X2=0 $Y2=0
cc_677 N_TE_B_M1001_g N_A_407_491#_c_1572_n 0.00149304f $X=1.425 $Y=2.775 $X2=0
+ $Y2=0
cc_678 N_TE_B_M1001_g N_A_407_491#_c_1574_n 6.97426e-19 $X=1.425 $Y=2.775 $X2=0
+ $Y2=0
cc_679 N_TE_B_c_676_n N_A_407_491#_c_1574_n 0.00556751f $X=2.08 $Y=1.86 $X2=0
+ $Y2=0
cc_680 N_TE_B_M1040_g N_A_407_491#_c_1562_n 0.00465516f $X=2.615 $Y=0.655 $X2=0
+ $Y2=0
cc_681 N_TE_B_c_674_n N_A_407_491#_c_1562_n 3.56531e-19 $X=2.615 $Y=1.395 $X2=0
+ $Y2=0
cc_682 N_TE_B_M1001_g N_VPWR_c_2667_n 0.00549284f $X=1.425 $Y=2.775 $X2=0 $Y2=0
cc_683 N_TE_B_M1001_g N_VPWR_c_2627_n 0.00636695f $X=1.425 $Y=2.775 $X2=0 $Y2=0
cc_684 N_TE_B_M1001_g KAPWR 0.00453421f $X=1.425 $Y=2.775 $X2=0 $Y2=0
cc_685 N_TE_B_M1008_g N_VGND_c_3665_n 0.0099303f $X=2.185 $Y=0.655 $X2=0 $Y2=0
cc_686 N_TE_B_M1040_g N_VGND_c_3665_n 6.06541e-19 $X=2.615 $Y=0.655 $X2=0 $Y2=0
cc_687 N_TE_B_M1040_g N_VGND_c_3666_n 0.00524039f $X=2.615 $Y=0.655 $X2=0 $Y2=0
cc_688 N_TE_B_M1008_g N_VGND_c_3684_n 0.00486043f $X=2.185 $Y=0.655 $X2=0 $Y2=0
cc_689 N_TE_B_M1040_g N_VGND_c_3684_n 0.00571722f $X=2.615 $Y=0.655 $X2=0 $Y2=0
cc_690 N_TE_B_M1008_g N_VGND_c_3707_n 0.00458264f $X=2.185 $Y=0.655 $X2=0 $Y2=0
cc_691 N_TE_B_M1040_g N_VGND_c_3707_n 0.0115803f $X=2.615 $Y=0.655 $X2=0 $Y2=0
cc_692 N_A_27_47#_c_729_n N_A_280_47#_c_830_n 2.19115e-19 $X=4.505 $Y=1.665
+ $X2=0 $Y2=0
cc_693 N_A_27_47#_c_729_n N_A_280_47#_c_831_n 3.66694e-19 $X=4.505 $Y=1.665
+ $X2=0 $Y2=0
cc_694 N_A_27_47#_M1036_g N_A_280_47#_c_832_n 0.0192513f $X=4.405 $Y=2.465 $X2=0
+ $Y2=0
cc_695 N_A_27_47#_c_729_n N_A_280_47#_c_832_n 0.00186897f $X=4.505 $Y=1.665
+ $X2=0 $Y2=0
cc_696 N_A_27_47#_c_731_n N_A_280_47#_c_818_n 0.0375387f $X=4.65 $Y=1.445 $X2=0
+ $Y2=0
cc_697 N_A_27_47#_c_738_n N_A_280_47#_c_818_n 3.24011e-19 $X=4.65 $Y=1.445 $X2=0
+ $Y2=0
cc_698 N_A_27_47#_c_729_n N_A_280_47#_c_819_n 0.0192675f $X=4.505 $Y=1.665 $X2=0
+ $Y2=0
cc_699 N_A_27_47#_c_731_n N_A_280_47#_c_819_n 0.0192513f $X=4.65 $Y=1.445 $X2=0
+ $Y2=0
cc_700 N_A_27_47#_c_738_n N_A_280_47#_c_819_n 0.00138777f $X=4.65 $Y=1.445 $X2=0
+ $Y2=0
cc_701 N_A_27_47#_c_731_n N_A_280_47#_c_821_n 0.0201175f $X=4.65 $Y=1.445 $X2=0
+ $Y2=0
cc_702 N_A_27_47#_c_738_n N_A_280_47#_c_821_n 0.00136891f $X=4.65 $Y=1.445 $X2=0
+ $Y2=0
cc_703 N_A_27_47#_c_729_n N_A_280_47#_c_826_n 0.0194057f $X=4.505 $Y=1.665 $X2=0
+ $Y2=0
cc_704 N_A_27_47#_c_729_n N_A_280_47#_c_859_n 0.0173804f $X=4.505 $Y=1.665 $X2=0
+ $Y2=0
cc_705 N_A_27_47#_c_729_n N_A_280_47#_c_837_n 0.0255369f $X=4.505 $Y=1.665 $X2=0
+ $Y2=0
cc_706 N_A_27_47#_c_729_n N_A_280_47#_c_838_n 0.0218939f $X=4.505 $Y=1.665 $X2=0
+ $Y2=0
cc_707 N_A_27_47#_c_729_n N_A_280_47#_c_905_n 3.62468e-19 $X=4.505 $Y=1.665
+ $X2=0 $Y2=0
cc_708 N_A_27_47#_c_729_n N_A_280_47#_c_839_n 0.00717939f $X=4.505 $Y=1.665
+ $X2=0 $Y2=0
cc_709 N_A_27_47#_c_729_n N_A_705_367#_c_1084_n 0.023097f $X=4.505 $Y=1.665
+ $X2=0 $Y2=0
cc_710 N_A_27_47#_c_751_n N_A_705_367#_c_1084_n 5.23641e-19 $X=4.65 $Y=1.665
+ $X2=0 $Y2=0
cc_711 N_A_27_47#_c_731_n N_A_705_367#_c_1084_n 0.00161001f $X=4.65 $Y=1.445
+ $X2=0 $Y2=0
cc_712 N_A_27_47#_c_738_n N_A_705_367#_c_1084_n 0.0109025f $X=4.65 $Y=1.445
+ $X2=0 $Y2=0
cc_713 N_A_27_47#_c_729_n N_A_705_367#_c_1023_n 0.0191194f $X=4.505 $Y=1.665
+ $X2=0 $Y2=0
cc_714 N_A_27_47#_c_751_n N_A_705_367#_c_1023_n 0.00132654f $X=4.65 $Y=1.665
+ $X2=0 $Y2=0
cc_715 N_A_27_47#_c_731_n N_A_705_367#_c_1023_n 0.00763655f $X=4.65 $Y=1.445
+ $X2=0 $Y2=0
cc_716 N_A_27_47#_c_738_n N_A_705_367#_c_1023_n 0.024374f $X=4.65 $Y=1.445 $X2=0
+ $Y2=0
cc_717 N_A_27_47#_c_729_n N_A_407_491#_c_1573_n 0.00118282f $X=4.505 $Y=1.665
+ $X2=0 $Y2=0
cc_718 N_A_27_47#_c_729_n N_A_407_491#_c_1562_n 0.0169523f $X=4.505 $Y=1.665
+ $X2=0 $Y2=0
cc_719 N_A_27_47#_M1066_g N_A_896_367#_c_1778_n 0.0114517f $X=4.835 $Y=2.465
+ $X2=0 $Y2=0
cc_720 N_A_27_47#_c_738_n N_A_896_367#_c_1778_n 0.00107941f $X=4.65 $Y=1.445
+ $X2=0 $Y2=0
cc_721 N_A_27_47#_c_731_n N_A_896_367#_c_1795_n 4.76986e-19 $X=4.65 $Y=1.445
+ $X2=0 $Y2=0
cc_722 N_A_27_47#_c_738_n N_A_896_367#_c_1795_n 0.0101634f $X=4.65 $Y=1.445
+ $X2=0 $Y2=0
cc_723 N_A_27_47#_c_732_n N_VPWR_c_2628_n 0.0466684f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_724 N_A_27_47#_M1066_g N_VPWR_c_2629_n 0.00452531f $X=4.835 $Y=2.465 $X2=0
+ $Y2=0
cc_725 N_A_27_47#_c_732_n N_VPWR_c_2666_n 0.0210467f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_726 N_A_27_47#_M1036_g N_VPWR_c_2667_n 0.00585385f $X=4.405 $Y=2.465 $X2=0
+ $Y2=0
cc_727 N_A_27_47#_M1066_g N_VPWR_c_2667_n 0.00549506f $X=4.835 $Y=2.465 $X2=0
+ $Y2=0
cc_728 N_A_27_47#_M1026_s N_VPWR_c_2627_n 0.00110569f $X=0.135 $Y=2.095 $X2=0
+ $Y2=0
cc_729 N_A_27_47#_M1036_g N_VPWR_c_2627_n 0.00535018f $X=4.405 $Y=2.465 $X2=0
+ $Y2=0
cc_730 N_A_27_47#_M1066_g N_VPWR_c_2627_n 0.0064266f $X=4.835 $Y=2.465 $X2=0
+ $Y2=0
cc_731 N_A_27_47#_c_732_n N_VPWR_c_2627_n 0.00303861f $X=0.26 $Y=0.42 $X2=0
+ $Y2=0
cc_732 N_A_27_47#_M1036_g KAPWR 0.00347624f $X=4.405 $Y=2.465 $X2=0 $Y2=0
cc_733 N_A_27_47#_M1066_g KAPWR 0.00191564f $X=4.835 $Y=2.465 $X2=0 $Y2=0
cc_734 N_A_27_47#_c_732_n KAPWR 0.0391539f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_735 N_A_27_47#_M1036_g N_KAPWR_c_3065_n 0.00187544f $X=4.405 $Y=2.465 $X2=0
+ $Y2=0
cc_736 N_A_27_47#_c_729_n N_KAPWR_c_3065_n 0.00892118f $X=4.505 $Y=1.665 $X2=0
+ $Y2=0
cc_737 N_A_27_47#_M1066_g N_KAPWR_c_3048_n 0.00376886f $X=4.835 $Y=2.465 $X2=0
+ $Y2=0
cc_738 N_A_27_47#_c_729_n N_VGND_c_3664_n 0.0103868f $X=4.505 $Y=1.665 $X2=0
+ $Y2=0
cc_739 N_A_27_47#_c_732_n N_VGND_c_3664_n 0.0183245f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_740 N_A_27_47#_c_729_n N_VGND_c_3666_n 0.00707505f $X=4.505 $Y=1.665 $X2=0
+ $Y2=0
cc_741 N_A_27_47#_c_732_n N_VGND_c_3680_n 0.0210467f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_742 N_A_27_47#_M1030_s N_VGND_c_3707_n 0.00215158f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_743 N_A_27_47#_c_732_n N_VGND_c_3707_n 0.0125689f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_744 N_A_280_47#_M1037_g N_A_705_367#_M1014_g 0.033599f $X=5.19 $Y=0.445 $X2=0
+ $Y2=0
cc_745 N_A_280_47#_c_822_n N_A_705_367#_c_998_n 0.0472035f $X=6.07 $Y=1.48 $X2=0
+ $Y2=0
cc_746 N_A_280_47#_c_825_n N_A_705_367#_c_998_n 0.033599f $X=5.19 $Y=0.995 $X2=0
+ $Y2=0
cc_747 N_A_280_47#_c_822_n N_A_705_367#_c_999_n 0.0160416f $X=6.07 $Y=1.48 $X2=0
+ $Y2=0
cc_748 N_A_280_47#_M1057_g N_A_705_367#_c_1000_n 0.0442533f $X=6.145 $Y=2.675
+ $X2=0 $Y2=0
cc_749 N_A_280_47#_c_831_n N_A_705_367#_c_1084_n 0.0122139f $X=3.45 $Y=1.715
+ $X2=0 $Y2=0
cc_750 N_A_280_47#_c_832_n N_A_705_367#_c_1084_n 0.00358974f $X=3.975 $Y=1.715
+ $X2=0 $Y2=0
cc_751 N_A_280_47#_c_819_n N_A_705_367#_c_1084_n 0.0335247f $X=4.05 $Y=0.995
+ $X2=0 $Y2=0
cc_752 N_A_280_47#_c_818_n N_A_705_367#_c_1023_n 0.0233579f $X=5.115 $Y=0.995
+ $X2=0 $Y2=0
cc_753 N_A_280_47#_c_819_n N_A_705_367#_c_1023_n 0.00879632f $X=4.05 $Y=0.995
+ $X2=0 $Y2=0
cc_754 N_A_280_47#_c_821_n N_A_705_367#_c_1023_n 0.0100608f $X=5.19 $Y=1.405
+ $X2=0 $Y2=0
cc_755 N_A_280_47#_c_822_n N_A_705_367#_c_1023_n 0.00626021f $X=6.07 $Y=1.48
+ $X2=0 $Y2=0
cc_756 N_A_280_47#_c_825_n N_A_705_367#_c_1023_n 0.00401069f $X=5.19 $Y=0.995
+ $X2=0 $Y2=0
cc_757 N_A_280_47#_c_819_n N_A_705_367#_c_1139_n 0.00790253f $X=4.05 $Y=0.995
+ $X2=0 $Y2=0
cc_758 N_A_280_47#_c_821_n N_A_705_367#_c_1024_n 0.00481054f $X=5.19 $Y=1.405
+ $X2=0 $Y2=0
cc_759 N_A_280_47#_c_822_n N_A_705_367#_c_1024_n 0.0123707f $X=6.07 $Y=1.48
+ $X2=0 $Y2=0
cc_760 N_A_280_47#_c_822_n N_A_705_367#_c_1025_n 0.00317014f $X=6.07 $Y=1.48
+ $X2=0 $Y2=0
cc_761 N_A_280_47#_M1057_g N_A_705_367#_c_1033_n 0.00259081f $X=6.145 $Y=2.675
+ $X2=0 $Y2=0
cc_762 N_A_280_47#_c_822_n N_A_705_367#_c_1039_n 0.00369083f $X=6.07 $Y=1.48
+ $X2=0 $Y2=0
cc_763 N_A_280_47#_M1057_g N_A_705_367#_c_1039_n 0.0104132f $X=6.145 $Y=2.675
+ $X2=0 $Y2=0
cc_764 N_A_280_47#_M1035_g N_A_407_491#_c_1572_n 0.0153997f $X=2.375 $Y=2.775
+ $X2=0 $Y2=0
cc_765 N_A_280_47#_c_829_n N_A_407_491#_c_1572_n 0.00168485f $X=2.45 $Y=2.22
+ $X2=0 $Y2=0
cc_766 N_A_280_47#_c_836_n N_A_407_491#_c_1572_n 0.0578045f $X=1.64 $Y=2.61
+ $X2=0 $Y2=0
cc_767 N_A_280_47#_c_828_n N_A_407_491#_c_1573_n 0.0178196f $X=2.9 $Y=2.22 $X2=0
+ $Y2=0
cc_768 N_A_280_47#_c_829_n N_A_407_491#_c_1573_n 0.00510721f $X=2.45 $Y=2.22
+ $X2=0 $Y2=0
cc_769 N_A_280_47#_c_830_n N_A_407_491#_c_1573_n 0.00334258f $X=2.975 $Y=2.145
+ $X2=0 $Y2=0
cc_770 N_A_280_47#_c_831_n N_A_407_491#_c_1573_n 0.00796025f $X=3.45 $Y=1.715
+ $X2=0 $Y2=0
cc_771 N_A_280_47#_c_819_n N_A_407_491#_c_1573_n 0.0024939f $X=4.05 $Y=0.995
+ $X2=0 $Y2=0
cc_772 N_A_280_47#_c_837_n N_A_407_491#_c_1573_n 0.054714f $X=2.9 $Y=1.845 $X2=0
+ $Y2=0
cc_773 N_A_280_47#_c_829_n N_A_407_491#_c_1574_n 0.00305576f $X=2.45 $Y=2.22
+ $X2=0 $Y2=0
cc_774 N_A_280_47#_c_836_n N_A_407_491#_c_1574_n 0.0135765f $X=1.64 $Y=2.61
+ $X2=0 $Y2=0
cc_775 N_A_280_47#_c_837_n N_A_407_491#_c_1574_n 0.0212076f $X=2.9 $Y=1.845
+ $X2=0 $Y2=0
cc_776 N_A_280_47#_M1063_g N_A_407_491#_c_1561_n 0.0126541f $X=3.565 $Y=0.445
+ $X2=0 $Y2=0
cc_777 N_A_280_47#_c_819_n N_A_407_491#_c_1561_n 0.00393981f $X=4.05 $Y=0.995
+ $X2=0 $Y2=0
cc_778 N_A_280_47#_c_830_n N_A_407_491#_c_1562_n 0.00158825f $X=2.975 $Y=2.145
+ $X2=0 $Y2=0
cc_779 N_A_280_47#_c_831_n N_A_407_491#_c_1562_n 0.00792805f $X=3.45 $Y=1.715
+ $X2=0 $Y2=0
cc_780 N_A_280_47#_M1063_g N_A_407_491#_c_1562_n 0.00587022f $X=3.565 $Y=0.445
+ $X2=0 $Y2=0
cc_781 N_A_280_47#_c_819_n N_A_407_491#_c_1562_n 0.0356455f $X=4.05 $Y=0.995
+ $X2=0 $Y2=0
cc_782 N_A_280_47#_c_837_n N_A_407_491#_c_1562_n 0.0105588f $X=2.9 $Y=1.845
+ $X2=0 $Y2=0
cc_783 N_A_280_47#_c_838_n N_A_407_491#_c_1562_n 0.0286729f $X=3.065 $Y=1.51
+ $X2=0 $Y2=0
cc_784 N_A_280_47#_M1063_g N_A_407_491#_c_1563_n 0.0151958f $X=3.565 $Y=0.445
+ $X2=0 $Y2=0
cc_785 N_A_280_47#_c_819_n N_A_407_491#_c_1563_n 0.0298942f $X=4.05 $Y=0.995
+ $X2=0 $Y2=0
cc_786 N_A_280_47#_M1037_g N_A_407_491#_c_1563_n 0.0130501f $X=5.19 $Y=0.445
+ $X2=0 $Y2=0
cc_787 N_A_280_47#_M1057_g N_A_896_367#_c_1778_n 0.00903174f $X=6.145 $Y=2.675
+ $X2=0 $Y2=0
cc_788 N_A_280_47#_c_822_n N_A_896_367#_c_1770_n 3.18767e-19 $X=6.07 $Y=1.48
+ $X2=0 $Y2=0
cc_789 N_A_280_47#_M1057_g N_A_896_367#_c_1781_n 0.00718137f $X=6.145 $Y=2.675
+ $X2=0 $Y2=0
cc_790 N_A_280_47#_M1057_g N_A_896_367#_c_1809_n 0.00969648f $X=6.145 $Y=2.675
+ $X2=0 $Y2=0
cc_791 N_A_280_47#_c_836_n N_VPWR_c_2628_n 0.0130916f $X=1.64 $Y=2.61 $X2=0
+ $Y2=0
cc_792 N_A_280_47#_M1057_g N_VPWR_c_2629_n 0.00251151f $X=6.145 $Y=2.675 $X2=0
+ $Y2=0
cc_793 N_A_280_47#_M1057_g N_VPWR_c_2648_n 0.00549284f $X=6.145 $Y=2.675 $X2=0
+ $Y2=0
cc_794 N_A_280_47#_M1035_g N_VPWR_c_2667_n 0.0054895f $X=2.375 $Y=2.775 $X2=0
+ $Y2=0
cc_795 N_A_280_47#_c_831_n N_VPWR_c_2667_n 0.00547467f $X=3.45 $Y=1.715 $X2=0
+ $Y2=0
cc_796 N_A_280_47#_c_832_n N_VPWR_c_2667_n 0.00585385f $X=3.975 $Y=1.715 $X2=0
+ $Y2=0
cc_797 N_A_280_47#_c_836_n N_VPWR_c_2667_n 0.0197852f $X=1.64 $Y=2.61 $X2=0
+ $Y2=0
cc_798 N_A_280_47#_M1001_d N_VPWR_c_2627_n 0.00110665f $X=1.5 $Y=2.455 $X2=0
+ $Y2=0
cc_799 N_A_280_47#_M1035_g N_VPWR_c_2627_n 0.00793447f $X=2.375 $Y=2.775 $X2=0
+ $Y2=0
cc_800 N_A_280_47#_c_831_n N_VPWR_c_2627_n 0.00677531f $X=3.45 $Y=1.715 $X2=0
+ $Y2=0
cc_801 N_A_280_47#_c_832_n N_VPWR_c_2627_n 0.00557705f $X=3.975 $Y=1.715 $X2=0
+ $Y2=0
cc_802 N_A_280_47#_M1057_g N_VPWR_c_2627_n 0.00487983f $X=6.145 $Y=2.675 $X2=0
+ $Y2=0
cc_803 N_A_280_47#_c_836_n N_VPWR_c_2627_n 0.00306434f $X=1.64 $Y=2.61 $X2=0
+ $Y2=0
cc_804 N_A_280_47#_c_837_n N_KAPWR_M1035_d 0.0012192f $X=2.9 $Y=1.845 $X2=-0.19
+ $Y2=-0.245
cc_805 N_A_280_47#_M1035_g KAPWR 0.00629849f $X=2.375 $Y=2.775 $X2=0 $Y2=0
cc_806 N_A_280_47#_c_828_n KAPWR 5.68091e-19 $X=2.9 $Y=2.22 $X2=0 $Y2=0
cc_807 N_A_280_47#_c_831_n KAPWR 0.00471376f $X=3.45 $Y=1.715 $X2=0 $Y2=0
cc_808 N_A_280_47#_c_832_n KAPWR 0.00372916f $X=3.975 $Y=1.715 $X2=0 $Y2=0
cc_809 N_A_280_47#_M1057_g KAPWR 0.00357997f $X=6.145 $Y=2.675 $X2=0 $Y2=0
cc_810 N_A_280_47#_c_836_n KAPWR 0.0308293f $X=1.64 $Y=2.61 $X2=0 $Y2=0
cc_811 N_A_280_47#_M1035_g N_KAPWR_c_3047_n 0.0120166f $X=2.375 $Y=2.775 $X2=0
+ $Y2=0
cc_812 N_A_280_47#_c_828_n N_KAPWR_c_3047_n 0.0124708f $X=2.9 $Y=2.22 $X2=0
+ $Y2=0
cc_813 N_A_280_47#_c_831_n N_KAPWR_c_3047_n 0.00760623f $X=3.45 $Y=1.715 $X2=0
+ $Y2=0
cc_814 N_A_280_47#_c_832_n N_KAPWR_c_3065_n 9.93406e-19 $X=3.975 $Y=1.715 $X2=0
+ $Y2=0
cc_815 N_A_280_47#_c_859_n N_VGND_M1045_d 0.00483959f $X=2.305 $Y=0.945 $X2=0
+ $Y2=0
cc_816 N_A_280_47#_c_859_n N_VGND_c_3665_n 0.0167297f $X=2.305 $Y=0.945 $X2=0
+ $Y2=0
cc_817 N_A_280_47#_M1063_g N_VGND_c_3666_n 0.00516038f $X=3.565 $Y=0.445 $X2=0
+ $Y2=0
cc_818 N_A_280_47#_c_819_n N_VGND_c_3666_n 0.00264602f $X=4.05 $Y=0.995 $X2=0
+ $Y2=0
cc_819 N_A_280_47#_c_838_n N_VGND_c_3666_n 0.00462935f $X=3.065 $Y=1.51 $X2=0
+ $Y2=0
cc_820 N_A_280_47#_c_983_p N_VGND_c_3682_n 0.0133395f $X=1.54 $Y=0.42 $X2=0
+ $Y2=0
cc_821 N_A_280_47#_c_884_n N_VGND_c_3684_n 0.0146655f $X=2.4 $Y=0.42 $X2=0 $Y2=0
cc_822 N_A_280_47#_M1063_g N_VGND_c_3686_n 0.00967207f $X=3.565 $Y=0.445 $X2=0
+ $Y2=0
cc_823 N_A_280_47#_M1063_g N_VGND_c_3687_n 0.00420091f $X=3.565 $Y=0.445 $X2=0
+ $Y2=0
cc_824 N_A_280_47#_M1037_g N_VGND_c_3688_n 0.00426565f $X=5.19 $Y=0.445 $X2=0
+ $Y2=0
cc_825 N_A_280_47#_M1013_s N_VGND_c_3707_n 0.00322829f $X=1.4 $Y=0.235 $X2=0
+ $Y2=0
cc_826 N_A_280_47#_M1008_s N_VGND_c_3707_n 0.00253254f $X=2.26 $Y=0.235 $X2=0
+ $Y2=0
cc_827 N_A_280_47#_M1063_g N_VGND_c_3707_n 0.00859912f $X=3.565 $Y=0.445 $X2=0
+ $Y2=0
cc_828 N_A_280_47#_M1037_g N_VGND_c_3707_n 0.00684647f $X=5.19 $Y=0.445 $X2=0
+ $Y2=0
cc_829 N_A_280_47#_c_983_p N_VGND_c_3707_n 0.00828095f $X=1.54 $Y=0.42 $X2=0
+ $Y2=0
cc_830 N_A_280_47#_c_859_n N_VGND_c_3707_n 0.0106723f $X=2.305 $Y=0.945 $X2=0
+ $Y2=0
cc_831 N_A_280_47#_c_884_n N_VGND_c_3707_n 0.00933292f $X=2.4 $Y=0.42 $X2=0
+ $Y2=0
cc_832 N_A_280_47#_M1037_g N_VGND_c_3708_n 0.00528389f $X=5.19 $Y=0.445 $X2=0
+ $Y2=0
cc_833 N_A_705_367#_c_997_n N_A_407_491#_c_1550_n 0.00990093f $X=6.43 $Y=1.12
+ $X2=0 $Y2=0
cc_834 N_A_705_367#_c_1029_n N_A_407_491#_c_1551_n 0.00378739f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_835 N_A_705_367#_c_999_n N_A_407_491#_c_1552_n 0.00990093f $X=6.505 $Y=1.575
+ $X2=0 $Y2=0
cc_836 N_A_705_367#_c_1029_n N_A_407_491#_c_1556_n 7.94408e-19 $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_837 N_A_705_367#_c_1029_n N_A_407_491#_M1018_g 0.00519027f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_838 N_A_705_367#_c_997_n N_A_407_491#_c_1559_n 0.00928501f $X=6.43 $Y=1.12
+ $X2=0 $Y2=0
cc_839 N_A_705_367#_c_1084_n N_A_407_491#_c_1573_n 0.0133627f $X=3.76 $Y=1.96
+ $X2=0 $Y2=0
cc_840 N_A_705_367#_c_1084_n N_A_407_491#_c_1562_n 0.0651163f $X=3.76 $Y=1.96
+ $X2=0 $Y2=0
cc_841 N_A_705_367#_c_1139_n N_A_407_491#_c_1562_n 0.0129498f $X=3.895 $Y=1.07
+ $X2=0 $Y2=0
cc_842 N_A_705_367#_M1014_g N_A_407_491#_c_1563_n 0.00140148f $X=5.55 $Y=0.445
+ $X2=0 $Y2=0
cc_843 N_A_705_367#_c_1023_n N_A_407_491#_c_1563_n 0.112897f $X=5.845 $Y=1.07
+ $X2=0 $Y2=0
cc_844 N_A_705_367#_c_1139_n N_A_407_491#_c_1563_n 0.0175813f $X=3.895 $Y=1.07
+ $X2=0 $Y2=0
cc_845 N_A_705_367#_M1014_g N_A_407_491#_c_1564_n 0.0127946f $X=5.55 $Y=0.445
+ $X2=0 $Y2=0
cc_846 N_A_705_367#_c_997_n N_A_407_491#_c_1564_n 0.00322328f $X=6.43 $Y=1.12
+ $X2=0 $Y2=0
cc_847 N_A_705_367#_c_1023_n N_A_407_491#_c_1564_n 0.00479493f $X=5.845 $Y=1.07
+ $X2=0 $Y2=0
cc_848 N_A_705_367#_c_1029_n N_A_407_491#_c_1566_n 0.0104808f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_849 N_A_705_367#_c_997_n N_A_407_491#_c_1567_n 5.11754e-19 $X=6.43 $Y=1.12
+ $X2=0 $Y2=0
cc_850 N_A_705_367#_c_1029_n N_A_407_491#_c_1569_n 0.00454721f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_851 N_A_705_367#_c_1029_n N_A_896_367#_c_1764_n 0.0114052f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_852 N_A_705_367#_c_1029_n N_A_896_367#_c_1774_n 0.00161676f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_853 N_A_705_367#_c_1029_n N_A_896_367#_c_1765_n 0.00387969f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_854 N_A_705_367#_c_1029_n N_A_896_367#_c_1776_n 0.00159563f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_855 N_A_705_367#_c_1029_n N_A_896_367#_c_1766_n 0.00207758f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_856 N_A_705_367#_c_1025_n N_A_896_367#_c_1778_n 0.00189944f $X=6.015 $Y=1.635
+ $X2=0 $Y2=0
cc_857 N_A_705_367#_c_1039_n N_A_896_367#_c_1778_n 0.00150331f $X=6.335 $Y=1.727
+ $X2=0 $Y2=0
cc_858 N_A_705_367#_M1014_g N_A_896_367#_c_1767_n 0.00482317f $X=5.55 $Y=0.445
+ $X2=0 $Y2=0
cc_859 N_A_705_367#_c_997_n N_A_896_367#_c_1767_n 0.00778057f $X=6.43 $Y=1.12
+ $X2=0 $Y2=0
cc_860 N_A_705_367#_c_1023_n N_A_896_367#_c_1767_n 0.0283388f $X=5.845 $Y=1.07
+ $X2=0 $Y2=0
cc_861 N_A_705_367#_M1014_g N_A_896_367#_c_1768_n 0.0040619f $X=5.55 $Y=0.445
+ $X2=0 $Y2=0
cc_862 N_A_705_367#_c_997_n N_A_896_367#_c_1768_n 0.0130828f $X=6.43 $Y=1.12
+ $X2=0 $Y2=0
cc_863 N_A_705_367#_c_1023_n N_A_896_367#_c_1768_n 0.0134469f $X=5.845 $Y=1.07
+ $X2=0 $Y2=0
cc_864 N_A_705_367#_c_1024_n N_A_896_367#_c_1768_n 0.00301617f $X=5.93 $Y=1.55
+ $X2=0 $Y2=0
cc_865 N_A_705_367#_c_997_n N_A_896_367#_c_1769_n 0.00303517f $X=6.43 $Y=1.12
+ $X2=0 $Y2=0
cc_866 N_A_705_367#_c_999_n N_A_896_367#_c_1769_n 0.0118469f $X=6.505 $Y=1.575
+ $X2=0 $Y2=0
cc_867 N_A_705_367#_c_1000_n N_A_896_367#_c_1769_n 0.00116575f $X=6.575 $Y=1.91
+ $X2=0 $Y2=0
cc_868 N_A_705_367#_c_1029_n N_A_896_367#_c_1769_n 0.00992693f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_869 N_A_705_367#_c_1030_n N_A_896_367#_c_1769_n 0.00673256f $X=6.625 $Y=1.665
+ $X2=0 $Y2=0
cc_870 N_A_705_367#_c_1033_n N_A_896_367#_c_1769_n 0.0254181f $X=6.48 $Y=1.665
+ $X2=0 $Y2=0
cc_871 N_A_705_367#_c_1024_n N_A_896_367#_c_1770_n 0.014358f $X=5.93 $Y=1.55
+ $X2=0 $Y2=0
cc_872 N_A_705_367#_c_1030_n N_A_896_367#_c_1770_n 5.65981e-19 $X=6.625 $Y=1.665
+ $X2=0 $Y2=0
cc_873 N_A_705_367#_c_1039_n N_A_896_367#_c_1770_n 0.0129849f $X=6.335 $Y=1.727
+ $X2=0 $Y2=0
cc_874 N_A_705_367#_c_1000_n N_A_896_367#_c_1779_n 0.00241807f $X=6.575 $Y=1.91
+ $X2=0 $Y2=0
cc_875 N_A_705_367#_M1027_g N_A_896_367#_c_1779_n 0.0098172f $X=6.575 $Y=2.675
+ $X2=0 $Y2=0
cc_876 N_A_705_367#_c_1029_n N_A_896_367#_c_1779_n 0.00126009f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_877 N_A_705_367#_c_1033_n N_A_896_367#_c_1779_n 0.0139257f $X=6.48 $Y=1.665
+ $X2=0 $Y2=0
cc_878 N_A_705_367#_c_999_n N_A_896_367#_c_1771_n 0.00526066f $X=6.505 $Y=1.575
+ $X2=0 $Y2=0
cc_879 N_A_705_367#_c_1000_n N_A_896_367#_c_1771_n 6.94059e-19 $X=6.575 $Y=1.91
+ $X2=0 $Y2=0
cc_880 N_A_705_367#_M1027_g N_A_896_367#_c_1771_n 0.00408777f $X=6.575 $Y=2.675
+ $X2=0 $Y2=0
cc_881 N_A_705_367#_c_1029_n N_A_896_367#_c_1771_n 0.018539f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_882 N_A_705_367#_c_1030_n N_A_896_367#_c_1771_n 4.71905e-19 $X=6.625 $Y=1.665
+ $X2=0 $Y2=0
cc_883 N_A_705_367#_c_1033_n N_A_896_367#_c_1771_n 0.0206727f $X=6.48 $Y=1.665
+ $X2=0 $Y2=0
cc_884 N_A_705_367#_c_1000_n N_A_896_367#_c_1781_n 0.00182326f $X=6.575 $Y=1.91
+ $X2=0 $Y2=0
cc_885 N_A_705_367#_M1027_g N_A_896_367#_c_1781_n 0.0114657f $X=6.575 $Y=2.675
+ $X2=0 $Y2=0
cc_886 N_A_705_367#_c_1033_n N_A_896_367#_c_1781_n 0.0120479f $X=6.48 $Y=1.665
+ $X2=0 $Y2=0
cc_887 N_A_705_367#_c_1039_n N_A_896_367#_c_1781_n 0.00398757f $X=6.335 $Y=1.727
+ $X2=0 $Y2=0
cc_888 N_A_705_367#_M1027_g N_A_896_367#_c_1809_n 0.00666366f $X=6.575 $Y=2.675
+ $X2=0 $Y2=0
cc_889 N_A_705_367#_c_1000_n N_A_896_367#_c_1772_n 0.0216572f $X=6.575 $Y=1.91
+ $X2=0 $Y2=0
cc_890 N_A_705_367#_c_1029_n N_A_896_367#_c_1772_n 0.00210717f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_891 N_A_705_367#_c_1033_n N_A_896_367#_c_1772_n 0.00118121f $X=6.48 $Y=1.665
+ $X2=0 $Y2=0
cc_892 N_A_705_367#_c_1029_n N_A_1486_47#_M1068_g 0.00212115f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_893 N_A_705_367#_c_1012_n N_A_1486_47#_c_1928_n 0.00460862f $X=19.065 $Y=1.65
+ $X2=0 $Y2=0
cc_894 N_A_705_367#_c_1007_n N_A_1486_47#_c_1929_n 0.131316f $X=16.915 $Y=1.65
+ $X2=0 $Y2=0
cc_895 N_A_705_367#_c_1022_n N_A_1486_47#_c_1929_n 0.00460862f $X=18.71 $Y=1.65
+ $X2=0 $Y2=0
cc_896 N_A_705_367#_c_1032_n N_A_1486_47#_c_1929_n 0.00225921f $X=22.285
+ $Y=1.665 $X2=0 $Y2=0
cc_897 N_A_705_367#_c_1037_n N_A_1486_47#_c_1929_n 4.34413e-19 $X=22.265 $Y=1.51
+ $X2=0 $Y2=0
cc_898 N_A_705_367#_c_1034_n N_A_1486_47#_c_1931_n 8.42755e-19 $X=19.345 $Y=1.51
+ $X2=0 $Y2=0
cc_899 N_A_705_367#_c_1035_n N_A_1486_47#_c_1935_n 8.42755e-19 $X=20.205 $Y=1.51
+ $X2=0 $Y2=0
cc_900 N_A_705_367#_c_1036_n N_A_1486_47#_c_1939_n 8.42755e-19 $X=21.065 $Y=1.51
+ $X2=0 $Y2=0
cc_901 N_A_705_367#_c_1029_n N_A_1486_47#_c_1942_n 0.00498952f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_902 N_A_705_367#_c_1032_n N_A_1486_47#_c_1943_n 0.00452657f $X=22.285
+ $Y=1.665 $X2=0 $Y2=0
cc_903 N_A_705_367#_c_1037_n N_A_1486_47#_c_1943_n 0.161537f $X=22.265 $Y=1.51
+ $X2=0 $Y2=0
cc_904 N_A_705_367#_c_1029_n N_A_1486_47#_c_1948_n 0.0165016f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_905 N_A_705_367#_c_1029_n N_A_1486_47#_c_1949_n 0.0388629f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_906 N_A_705_367#_c_1029_n N_A_1486_47#_c_1950_n 0.00619203f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_907 N_A_705_367#_c_1029_n N_A_1486_47#_c_1951_n 0.0527876f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_908 N_A_705_367#_c_1029_n N_A_1486_47#_c_1952_n 0.0239718f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_909 N_A_705_367#_c_1026_n N_A_1486_47#_c_1953_n 0.0198201f $X=14.285 $Y=1.55
+ $X2=0 $Y2=0
cc_910 N_A_705_367#_c_1027_n N_A_1486_47#_c_1953_n 0.00608621f $X=14.222
+ $Y=1.095 $X2=0 $Y2=0
cc_911 N_A_705_367#_c_1029_n N_A_1486_47#_c_1953_n 0.304992f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_912 N_A_705_367#_c_1031_n N_A_1486_47#_c_1953_n 0.00559893f $X=14.68 $Y=1.665
+ $X2=0 $Y2=0
cc_913 N_A_705_367#_c_1029_n N_A_1486_47#_c_1954_n 0.0234815f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_914 N_A_705_367#_c_1003_n N_A_1486_47#_c_1955_n 0.00146859f $X=15.195 $Y=1.65
+ $X2=0 $Y2=0
cc_915 N_A_705_367#_c_1026_n N_A_1486_47#_c_1955_n 0.00209523f $X=14.285 $Y=1.55
+ $X2=0 $Y2=0
cc_916 N_A_705_367#_c_1032_n N_A_1486_47#_c_1955_n 0.372459f $X=22.285 $Y=1.665
+ $X2=0 $Y2=0
cc_917 N_A_705_367#_c_1018_n N_A_1486_47#_c_1956_n 0.00146859f $X=16.99 $Y=1.65
+ $X2=0 $Y2=0
cc_918 N_A_705_367#_c_1029_n N_A_1486_47#_c_1957_n 0.00901644f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_919 N_A_705_367#_c_1029_n N_A_1486_47#_c_1958_n 0.0113327f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_920 N_A_705_367#_c_1013_n N_A_1486_47#_c_1960_n 0.131316f $X=14.84 $Y=1.65
+ $X2=0 $Y2=0
cc_921 N_A_705_367#_c_1026_n N_A_1486_47#_c_1960_n 3.58093e-19 $X=14.285 $Y=1.55
+ $X2=0 $Y2=0
cc_922 N_A_705_367#_c_1027_n N_A_1486_47#_c_1960_n 9.7253e-19 $X=14.222 $Y=1.095
+ $X2=0 $Y2=0
cc_923 N_A_705_367#_c_1031_n N_A_1486_47#_c_1960_n 2.39489e-19 $X=14.68 $Y=1.665
+ $X2=0 $Y2=0
cc_924 N_A_705_367#_c_1032_n N_A_1486_47#_c_1960_n 0.00294233f $X=22.285
+ $Y=1.665 $X2=0 $Y2=0
cc_925 N_A_705_367#_c_1003_n N_A_1486_47#_c_1961_n 0.00142857f $X=15.195 $Y=1.65
+ $X2=0 $Y2=0
cc_926 N_A_705_367#_c_1026_n N_A_1486_47#_c_1961_n 0.00506713f $X=14.285 $Y=1.55
+ $X2=0 $Y2=0
cc_927 N_A_705_367#_c_1032_n N_A_1486_47#_c_1961_n 8.68597e-19 $X=22.285
+ $Y=1.665 $X2=0 $Y2=0
cc_928 N_A_705_367#_c_1005_n N_A_1486_47#_c_1962_n 0.00329165f $X=16.055 $Y=1.65
+ $X2=0 $Y2=0
cc_929 N_A_705_367#_c_1032_n N_A_1486_47#_c_1962_n 0.00149426f $X=22.285
+ $Y=1.665 $X2=0 $Y2=0
cc_930 N_A_705_367#_c_1007_n N_A_1486_47#_c_1963_n 0.00329165f $X=16.915 $Y=1.65
+ $X2=0 $Y2=0
cc_931 N_A_705_367#_c_1032_n N_A_1486_47#_c_1963_n 0.00149426f $X=22.285
+ $Y=1.665 $X2=0 $Y2=0
cc_932 N_A_705_367#_c_1009_n N_A_1486_47#_c_1964_n 0.00329165f $X=17.775 $Y=1.65
+ $X2=0 $Y2=0
cc_933 N_A_705_367#_c_1032_n N_A_1486_47#_c_1964_n 0.00149426f $X=22.285
+ $Y=1.665 $X2=0 $Y2=0
cc_934 N_A_705_367#_c_1011_n N_A_1486_47#_c_1965_n 0.00329165f $X=18.635 $Y=1.65
+ $X2=0 $Y2=0
cc_935 N_A_705_367#_c_1032_n N_A_1486_47#_c_1965_n 0.00149426f $X=22.285
+ $Y=1.665 $X2=0 $Y2=0
cc_936 N_A_705_367#_c_1029_n N_A_c_2281_n 0.00154649f $X=14.5 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_937 N_A_705_367#_c_1029_n N_A_c_2282_n 0.00163123f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_938 N_A_705_367#_c_1029_n N_A_c_2283_n 0.0019639f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_939 N_A_705_367#_c_1029_n N_A_c_2286_n 8.5564e-19 $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_940 N_A_705_367#_c_1029_n N_A_c_2267_n 0.003034f $X=14.5 $Y=1.665 $X2=0 $Y2=0
cc_941 N_A_705_367#_c_1029_n N_A_c_2268_n 0.00191611f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_942 N_A_705_367#_c_1087_n N_A_c_2289_n 0.00157406f $X=13.41 $Y=1.87 $X2=0
+ $Y2=0
cc_943 N_A_705_367#_c_1029_n N_A_c_2289_n 0.00570979f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_944 N_A_705_367#_c_1087_n N_A_c_2270_n 0.00203878f $X=13.41 $Y=1.87 $X2=0
+ $Y2=0
cc_945 N_A_705_367#_c_1029_n N_A_c_2270_n 0.00105254f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_946 N_A_705_367#_c_1026_n N_A_M1041_g 3.64544e-19 $X=14.285 $Y=1.55 $X2=0
+ $Y2=0
cc_947 N_A_705_367#_c_1260_p N_A_c_2291_n 0.0141715f $X=13.245 $Y=1.98 $X2=0
+ $Y2=0
cc_948 N_A_705_367#_c_1086_n N_A_c_2291_n 0.0130694f $X=14.2 $Y=1.87 $X2=0 $Y2=0
cc_949 N_A_705_367#_c_1087_n N_A_c_2291_n 0.00119606f $X=13.41 $Y=1.87 $X2=0
+ $Y2=0
cc_950 N_A_705_367#_c_1028_n N_A_c_2291_n 2.99261e-19 $X=14.37 $Y=1.665 $X2=0
+ $Y2=0
cc_951 N_A_705_367#_c_1029_n N_A_c_2291_n 0.00148605f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_952 N_A_705_367#_c_1029_n N_A_c_2272_n 0.0201994f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_953 N_A_705_367#_c_1029_n N_A_c_2274_n 0.00168794f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_954 N_A_705_367#_c_1029_n N_A_c_2278_n 9.81943e-19 $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_955 N_A_705_367#_c_1028_n N_A_c_2279_n 0.00265957f $X=14.37 $Y=1.665 $X2=0
+ $Y2=0
cc_956 N_A_705_367#_c_1029_n N_A_c_2279_n 0.00214403f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_957 N_A_705_367#_c_1002_n N_A_2063_47#_c_2481_n 0.00726207f $X=14.485 $Y=1.65
+ $X2=0 $Y2=0
cc_958 N_A_705_367#_c_1086_n N_A_2063_47#_c_2481_n 0.00270933f $X=14.2 $Y=1.87
+ $X2=0 $Y2=0
cc_959 N_A_705_367#_c_1026_n N_A_2063_47#_c_2481_n 0.0104899f $X=14.285 $Y=1.55
+ $X2=0 $Y2=0
cc_960 N_A_705_367#_c_1027_n N_A_2063_47#_c_2481_n 0.00340113f $X=14.222
+ $Y=1.095 $X2=0 $Y2=0
cc_961 N_A_705_367#_c_1029_n N_A_2063_47#_c_2481_n 6.29496e-19 $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_962 N_A_705_367#_c_1031_n N_A_2063_47#_c_2481_n 0.00181843f $X=14.68 $Y=1.665
+ $X2=0 $Y2=0
cc_963 N_A_705_367#_c_1276_p N_A_2063_47#_c_2482_n 0.00523642f $X=14.17 $Y=0.815
+ $X2=0 $Y2=0
cc_964 N_A_705_367#_c_1026_n N_A_2063_47#_c_2482_n 0.00237781f $X=14.285 $Y=1.55
+ $X2=0 $Y2=0
cc_965 N_A_705_367#_c_1027_n N_A_2063_47#_c_2482_n 0.00268423f $X=14.222
+ $Y=1.095 $X2=0 $Y2=0
cc_966 N_A_705_367#_c_1029_n N_A_2063_47#_c_2486_n 0.0129669f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_967 N_A_705_367#_c_1029_n N_A_2063_47#_c_2489_n 0.0066187f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_968 N_A_705_367#_c_1086_n N_A_2063_47#_c_2490_n 0.0363169f $X=14.2 $Y=1.87
+ $X2=0 $Y2=0
cc_969 N_A_705_367#_c_1087_n N_A_2063_47#_c_2490_n 0.0167791f $X=13.41 $Y=1.87
+ $X2=0 $Y2=0
cc_970 N_A_705_367#_c_1026_n N_A_2063_47#_c_2490_n 0.0247486f $X=14.285 $Y=1.55
+ $X2=0 $Y2=0
cc_971 N_A_705_367#_c_1029_n N_A_2063_47#_c_2490_n 0.0435512f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_972 N_A_705_367#_c_1029_n N_A_2063_47#_c_2496_n 0.00722937f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_973 N_A_705_367#_c_1002_n N_A_2063_47#_c_2492_n 0.00147739f $X=14.485 $Y=1.65
+ $X2=0 $Y2=0
cc_974 N_A_705_367#_c_1086_n N_A_2063_47#_c_2492_n 0.00656991f $X=14.2 $Y=1.87
+ $X2=0 $Y2=0
cc_975 N_A_705_367#_c_1026_n N_A_2063_47#_c_2492_n 0.0056917f $X=14.285 $Y=1.55
+ $X2=0 $Y2=0
cc_976 N_A_705_367#_c_1029_n N_A_2063_47#_c_2492_n 0.00392599f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_977 N_A_705_367#_c_1026_n N_A_2063_47#_c_2493_n 0.00184046f $X=14.285 $Y=1.55
+ $X2=0 $Y2=0
cc_978 N_A_705_367#_c_1027_n N_A_2063_47#_c_2493_n 4.47617e-19 $X=14.222
+ $Y=1.095 $X2=0 $Y2=0
cc_979 N_A_705_367#_c_1086_n N_VPWR_M1004_s 0.0022499f $X=14.2 $Y=1.87 $X2=0
+ $Y2=0
cc_980 N_A_705_367#_c_1028_n N_VPWR_M1004_s 0.00120577f $X=14.37 $Y=1.665 $X2=0
+ $Y2=0
cc_981 N_A_705_367#_M1027_g N_VPWR_c_2630_n 0.00485222f $X=6.575 $Y=2.675 $X2=0
+ $Y2=0
cc_982 N_A_705_367#_c_1029_n N_VPWR_c_2632_n 0.00990802f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_983 N_A_705_367#_c_1042_n N_VPWR_c_2636_n 0.0142841f $X=14.41 $Y=1.725 $X2=0
+ $Y2=0
cc_984 N_A_705_367#_c_1045_n N_VPWR_c_2636_n 8.40773e-19 $X=14.84 $Y=1.725 $X2=0
+ $Y2=0
cc_985 N_A_705_367#_c_1260_p N_VPWR_c_2636_n 0.00147385f $X=13.245 $Y=1.98 $X2=0
+ $Y2=0
cc_986 N_A_705_367#_c_1086_n N_VPWR_c_2636_n 0.0128494f $X=14.2 $Y=1.87 $X2=0
+ $Y2=0
cc_987 N_A_705_367#_c_1028_n N_VPWR_c_2636_n 0.00807505f $X=14.37 $Y=1.665 $X2=0
+ $Y2=0
cc_988 N_A_705_367#_c_1029_n N_VPWR_c_2636_n 0.00131333f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_989 N_A_705_367#_c_1042_n N_VPWR_c_2637_n 7.78238e-19 $X=14.41 $Y=1.725 $X2=0
+ $Y2=0
cc_990 N_A_705_367#_c_1045_n N_VPWR_c_2637_n 0.0118036f $X=14.84 $Y=1.725 $X2=0
+ $Y2=0
cc_991 N_A_705_367#_c_1047_n N_VPWR_c_2637_n 0.00349139f $X=15.27 $Y=1.725 $X2=0
+ $Y2=0
cc_992 N_A_705_367#_c_1049_n N_VPWR_c_2638_n 0.00344889f $X=15.7 $Y=1.725 $X2=0
+ $Y2=0
cc_993 N_A_705_367#_c_1005_n N_VPWR_c_2638_n 0.0022751f $X=16.055 $Y=1.65 $X2=0
+ $Y2=0
cc_994 N_A_705_367#_c_1051_n N_VPWR_c_2638_n 0.00344889f $X=16.13 $Y=1.725 $X2=0
+ $Y2=0
cc_995 N_A_705_367#_c_1053_n N_VPWR_c_2639_n 0.00344889f $X=16.56 $Y=1.725 $X2=0
+ $Y2=0
cc_996 N_A_705_367#_c_1007_n N_VPWR_c_2639_n 0.0022751f $X=16.915 $Y=1.65 $X2=0
+ $Y2=0
cc_997 N_A_705_367#_c_1055_n N_VPWR_c_2639_n 0.00344889f $X=16.99 $Y=1.725 $X2=0
+ $Y2=0
cc_998 N_A_705_367#_c_1057_n N_VPWR_c_2640_n 0.00344889f $X=17.42 $Y=1.725 $X2=0
+ $Y2=0
cc_999 N_A_705_367#_c_1009_n N_VPWR_c_2640_n 0.0022751f $X=17.775 $Y=1.65 $X2=0
+ $Y2=0
cc_1000 N_A_705_367#_c_1059_n N_VPWR_c_2640_n 0.00344889f $X=17.85 $Y=1.725
+ $X2=0 $Y2=0
cc_1001 N_A_705_367#_c_1059_n N_VPWR_c_2641_n 0.00549284f $X=17.85 $Y=1.725
+ $X2=0 $Y2=0
cc_1002 N_A_705_367#_c_1061_n N_VPWR_c_2641_n 0.00549284f $X=18.28 $Y=1.725
+ $X2=0 $Y2=0
cc_1003 N_A_705_367#_c_1061_n N_VPWR_c_2642_n 0.00344889f $X=18.28 $Y=1.725
+ $X2=0 $Y2=0
cc_1004 N_A_705_367#_c_1011_n N_VPWR_c_2642_n 0.0022751f $X=18.635 $Y=1.65 $X2=0
+ $Y2=0
cc_1005 N_A_705_367#_c_1063_n N_VPWR_c_2642_n 0.00344889f $X=18.71 $Y=1.725
+ $X2=0 $Y2=0
cc_1006 N_A_705_367#_c_1065_n N_VPWR_c_2643_n 0.00344889f $X=19.14 $Y=1.725
+ $X2=0 $Y2=0
cc_1007 N_A_705_367#_c_1066_n N_VPWR_c_2643_n 0.00344889f $X=19.57 $Y=1.725
+ $X2=0 $Y2=0
cc_1008 N_A_705_367#_c_1034_n N_VPWR_c_2643_n 0.00309227f $X=19.345 $Y=1.51
+ $X2=0 $Y2=0
cc_1009 N_A_705_367#_c_1037_n N_VPWR_c_2643_n 6.2031e-19 $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1010 N_A_705_367#_c_1067_n N_VPWR_c_2644_n 0.00344889f $X=20 $Y=1.725 $X2=0
+ $Y2=0
cc_1011 N_A_705_367#_c_1068_n N_VPWR_c_2644_n 0.00344889f $X=20.43 $Y=1.725
+ $X2=0 $Y2=0
cc_1012 N_A_705_367#_c_1035_n N_VPWR_c_2644_n 0.00309227f $X=20.205 $Y=1.51
+ $X2=0 $Y2=0
cc_1013 N_A_705_367#_c_1037_n N_VPWR_c_2644_n 6.2031e-19 $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1014 N_A_705_367#_c_1069_n N_VPWR_c_2645_n 0.00344889f $X=20.86 $Y=1.725
+ $X2=0 $Y2=0
cc_1015 N_A_705_367#_c_1070_n N_VPWR_c_2645_n 0.00344889f $X=21.29 $Y=1.725
+ $X2=0 $Y2=0
cc_1016 N_A_705_367#_c_1036_n N_VPWR_c_2645_n 0.00309227f $X=21.065 $Y=1.51
+ $X2=0 $Y2=0
cc_1017 N_A_705_367#_c_1037_n N_VPWR_c_2645_n 6.2031e-19 $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1018 N_A_705_367#_c_1071_n N_VPWR_c_2646_n 0.00344889f $X=21.72 $Y=1.725
+ $X2=0 $Y2=0
cc_1019 N_A_705_367#_c_1072_n N_VPWR_c_2646_n 0.00344889f $X=22.15 $Y=1.725
+ $X2=0 $Y2=0
cc_1020 N_A_705_367#_c_1037_n N_VPWR_c_2646_n 6.2031e-19 $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1021 N_A_705_367#_c_1038_n N_VPWR_c_2646_n 0.00309227f $X=22.265 $Y=1.51
+ $X2=0 $Y2=0
cc_1022 N_A_705_367#_c_1073_n N_VPWR_c_2647_n 0.00664936f $X=22.58 $Y=1.725
+ $X2=0 $Y2=0
cc_1023 N_A_705_367#_M1027_g N_VPWR_c_2648_n 0.00549284f $X=6.575 $Y=2.675 $X2=0
+ $Y2=0
cc_1024 N_A_705_367#_c_1042_n N_VPWR_c_2650_n 0.00486043f $X=14.41 $Y=1.725
+ $X2=0 $Y2=0
cc_1025 N_A_705_367#_c_1045_n N_VPWR_c_2650_n 0.00486043f $X=14.84 $Y=1.725
+ $X2=0 $Y2=0
cc_1026 N_A_705_367#_c_1047_n N_VPWR_c_2652_n 0.00549284f $X=15.27 $Y=1.725
+ $X2=0 $Y2=0
cc_1027 N_A_705_367#_c_1049_n N_VPWR_c_2652_n 0.00549284f $X=15.7 $Y=1.725 $X2=0
+ $Y2=0
cc_1028 N_A_705_367#_c_1051_n N_VPWR_c_2654_n 0.00549284f $X=16.13 $Y=1.725
+ $X2=0 $Y2=0
cc_1029 N_A_705_367#_c_1053_n N_VPWR_c_2654_n 0.00549284f $X=16.56 $Y=1.725
+ $X2=0 $Y2=0
cc_1030 N_A_705_367#_c_1055_n N_VPWR_c_2656_n 0.00549284f $X=16.99 $Y=1.725
+ $X2=0 $Y2=0
cc_1031 N_A_705_367#_c_1057_n N_VPWR_c_2656_n 0.00549284f $X=17.42 $Y=1.725
+ $X2=0 $Y2=0
cc_1032 N_A_705_367#_c_1063_n N_VPWR_c_2658_n 0.00549284f $X=18.71 $Y=1.725
+ $X2=0 $Y2=0
cc_1033 N_A_705_367#_c_1065_n N_VPWR_c_2658_n 0.00549284f $X=19.14 $Y=1.725
+ $X2=0 $Y2=0
cc_1034 N_A_705_367#_c_1066_n N_VPWR_c_2660_n 0.00549284f $X=19.57 $Y=1.725
+ $X2=0 $Y2=0
cc_1035 N_A_705_367#_c_1067_n N_VPWR_c_2660_n 0.00549284f $X=20 $Y=1.725 $X2=0
+ $Y2=0
cc_1036 N_A_705_367#_c_1068_n N_VPWR_c_2662_n 0.00549284f $X=20.43 $Y=1.725
+ $X2=0 $Y2=0
cc_1037 N_A_705_367#_c_1069_n N_VPWR_c_2662_n 0.00549284f $X=20.86 $Y=1.725
+ $X2=0 $Y2=0
cc_1038 N_A_705_367#_c_1070_n N_VPWR_c_2664_n 0.00549284f $X=21.29 $Y=1.725
+ $X2=0 $Y2=0
cc_1039 N_A_705_367#_c_1071_n N_VPWR_c_2664_n 0.00549284f $X=21.72 $Y=1.725
+ $X2=0 $Y2=0
cc_1040 N_A_705_367#_c_1084_n N_VPWR_c_2667_n 0.0127414f $X=3.76 $Y=1.96 $X2=0
+ $Y2=0
cc_1041 N_A_705_367#_c_1072_n N_VPWR_c_2672_n 0.00549284f $X=22.15 $Y=1.725
+ $X2=0 $Y2=0
cc_1042 N_A_705_367#_c_1073_n N_VPWR_c_2672_n 0.00549284f $X=22.58 $Y=1.725
+ $X2=0 $Y2=0
cc_1043 N_A_705_367#_M1011_s N_VPWR_c_2627_n 0.00215585f $X=3.525 $Y=1.835 $X2=0
+ $Y2=0
cc_1044 N_A_705_367#_M1016_d N_VPWR_c_2627_n 0.00114246f $X=13.105 $Y=1.835
+ $X2=0 $Y2=0
cc_1045 N_A_705_367#_M1027_g N_VPWR_c_2627_n 0.00636983f $X=6.575 $Y=2.675 $X2=0
+ $Y2=0
cc_1046 N_A_705_367#_c_1042_n N_VPWR_c_2627_n 0.00359111f $X=14.41 $Y=1.725
+ $X2=0 $Y2=0
cc_1047 N_A_705_367#_c_1045_n N_VPWR_c_2627_n 0.00359111f $X=14.84 $Y=1.725
+ $X2=0 $Y2=0
cc_1048 N_A_705_367#_c_1047_n N_VPWR_c_2627_n 0.0050448f $X=15.27 $Y=1.725 $X2=0
+ $Y2=0
cc_1049 N_A_705_367#_c_1049_n N_VPWR_c_2627_n 0.0050448f $X=15.7 $Y=1.725 $X2=0
+ $Y2=0
cc_1050 N_A_705_367#_c_1051_n N_VPWR_c_2627_n 0.0050448f $X=16.13 $Y=1.725 $X2=0
+ $Y2=0
cc_1051 N_A_705_367#_c_1053_n N_VPWR_c_2627_n 0.0050448f $X=16.56 $Y=1.725 $X2=0
+ $Y2=0
cc_1052 N_A_705_367#_c_1055_n N_VPWR_c_2627_n 0.0050448f $X=16.99 $Y=1.725 $X2=0
+ $Y2=0
cc_1053 N_A_705_367#_c_1057_n N_VPWR_c_2627_n 0.0050448f $X=17.42 $Y=1.725 $X2=0
+ $Y2=0
cc_1054 N_A_705_367#_c_1059_n N_VPWR_c_2627_n 0.0050448f $X=17.85 $Y=1.725 $X2=0
+ $Y2=0
cc_1055 N_A_705_367#_c_1061_n N_VPWR_c_2627_n 0.0050448f $X=18.28 $Y=1.725 $X2=0
+ $Y2=0
cc_1056 N_A_705_367#_c_1063_n N_VPWR_c_2627_n 0.0050448f $X=18.71 $Y=1.725 $X2=0
+ $Y2=0
cc_1057 N_A_705_367#_c_1065_n N_VPWR_c_2627_n 0.0050448f $X=19.14 $Y=1.725 $X2=0
+ $Y2=0
cc_1058 N_A_705_367#_c_1066_n N_VPWR_c_2627_n 0.0050448f $X=19.57 $Y=1.725 $X2=0
+ $Y2=0
cc_1059 N_A_705_367#_c_1067_n N_VPWR_c_2627_n 0.0050448f $X=20 $Y=1.725 $X2=0
+ $Y2=0
cc_1060 N_A_705_367#_c_1068_n N_VPWR_c_2627_n 0.0050448f $X=20.43 $Y=1.725 $X2=0
+ $Y2=0
cc_1061 N_A_705_367#_c_1069_n N_VPWR_c_2627_n 0.0050448f $X=20.86 $Y=1.725 $X2=0
+ $Y2=0
cc_1062 N_A_705_367#_c_1070_n N_VPWR_c_2627_n 0.0050448f $X=21.29 $Y=1.725 $X2=0
+ $Y2=0
cc_1063 N_A_705_367#_c_1071_n N_VPWR_c_2627_n 0.0050448f $X=21.72 $Y=1.725 $X2=0
+ $Y2=0
cc_1064 N_A_705_367#_c_1072_n N_VPWR_c_2627_n 0.0050448f $X=22.15 $Y=1.725 $X2=0
+ $Y2=0
cc_1065 N_A_705_367#_c_1073_n N_VPWR_c_2627_n 0.0063445f $X=22.58 $Y=1.725 $X2=0
+ $Y2=0
cc_1066 N_A_705_367#_c_1084_n N_VPWR_c_2627_n 0.00206609f $X=3.76 $Y=1.96 $X2=0
+ $Y2=0
cc_1067 N_A_705_367#_M1011_s KAPWR 0.00293013f $X=3.525 $Y=1.835 $X2=0 $Y2=0
cc_1068 N_A_705_367#_M1016_d KAPWR 0.00367316f $X=13.105 $Y=1.835 $X2=0 $Y2=0
cc_1069 N_A_705_367#_M1027_g KAPWR 0.00218356f $X=6.575 $Y=2.675 $X2=0 $Y2=0
cc_1070 N_A_705_367#_c_1042_n KAPWR 0.006024f $X=14.41 $Y=1.725 $X2=0 $Y2=0
cc_1071 N_A_705_367#_c_1045_n KAPWR 0.00227958f $X=14.84 $Y=1.725 $X2=0 $Y2=0
cc_1072 N_A_705_367#_c_1047_n KAPWR 0.00277511f $X=15.27 $Y=1.725 $X2=0 $Y2=0
cc_1073 N_A_705_367#_c_1049_n KAPWR 0.00330943f $X=15.7 $Y=1.725 $X2=0 $Y2=0
cc_1074 N_A_705_367#_c_1051_n KAPWR 0.00330943f $X=16.13 $Y=1.725 $X2=0 $Y2=0
cc_1075 N_A_705_367#_c_1053_n KAPWR 0.00330943f $X=16.56 $Y=1.725 $X2=0 $Y2=0
cc_1076 N_A_705_367#_c_1055_n KAPWR 0.00330943f $X=16.99 $Y=1.725 $X2=0 $Y2=0
cc_1077 N_A_705_367#_c_1057_n KAPWR 0.00330943f $X=17.42 $Y=1.725 $X2=0 $Y2=0
cc_1078 N_A_705_367#_c_1059_n KAPWR 0.00330943f $X=17.85 $Y=1.725 $X2=0 $Y2=0
cc_1079 N_A_705_367#_c_1061_n KAPWR 0.00330943f $X=18.28 $Y=1.725 $X2=0 $Y2=0
cc_1080 N_A_705_367#_c_1063_n KAPWR 0.00330943f $X=18.71 $Y=1.725 $X2=0 $Y2=0
cc_1081 N_A_705_367#_c_1065_n KAPWR 0.00330943f $X=19.14 $Y=1.725 $X2=0 $Y2=0
cc_1082 N_A_705_367#_c_1066_n KAPWR 0.00330943f $X=19.57 $Y=1.725 $X2=0 $Y2=0
cc_1083 N_A_705_367#_c_1067_n KAPWR 0.00330943f $X=20 $Y=1.725 $X2=0 $Y2=0
cc_1084 N_A_705_367#_c_1068_n KAPWR 0.00330943f $X=20.43 $Y=1.725 $X2=0 $Y2=0
cc_1085 N_A_705_367#_c_1069_n KAPWR 0.00330943f $X=20.86 $Y=1.725 $X2=0 $Y2=0
cc_1086 N_A_705_367#_c_1070_n KAPWR 0.00330943f $X=21.29 $Y=1.725 $X2=0 $Y2=0
cc_1087 N_A_705_367#_c_1071_n KAPWR 0.00330943f $X=21.72 $Y=1.725 $X2=0 $Y2=0
cc_1088 N_A_705_367#_c_1072_n KAPWR 0.00330943f $X=22.15 $Y=1.725 $X2=0 $Y2=0
cc_1089 N_A_705_367#_c_1073_n KAPWR 0.00753768f $X=22.58 $Y=1.725 $X2=0 $Y2=0
cc_1090 N_A_705_367#_c_1084_n KAPWR 0.0213093f $X=3.76 $Y=1.96 $X2=0 $Y2=0
cc_1091 N_A_705_367#_c_1260_p KAPWR 0.00833653f $X=13.245 $Y=1.98 $X2=0 $Y2=0
cc_1092 N_A_705_367#_c_1084_n N_KAPWR_c_3047_n 0.0303854f $X=3.76 $Y=1.96 $X2=0
+ $Y2=0
cc_1093 N_A_705_367#_c_1084_n N_KAPWR_c_3065_n 0.0156777f $X=3.76 $Y=1.96 $X2=0
+ $Y2=0
cc_1094 N_A_705_367#_c_1029_n N_A_1492_367#_c_3237_n 0.00892417f $X=14.5
+ $Y=1.665 $X2=0 $Y2=0
cc_1095 N_A_705_367#_c_1029_n N_A_1492_367#_c_3238_n 0.00593911f $X=14.5
+ $Y=1.665 $X2=0 $Y2=0
cc_1096 N_A_705_367#_c_1086_n N_A_2345_367#_M1069_s 0.00308603f $X=14.2 $Y=1.87
+ $X2=0 $Y2=0
cc_1097 N_A_705_367#_c_1029_n N_A_2345_367#_c_3306_n 0.0176781f $X=14.5 $Y=1.665
+ $X2=0 $Y2=0
cc_1098 N_A_705_367#_c_1029_n N_A_2345_367#_c_3307_n 0.00780084f $X=14.5
+ $Y=1.665 $X2=0 $Y2=0
cc_1099 N_A_705_367#_M1016_d N_A_2345_367#_c_3327_n 0.00236976f $X=13.105
+ $Y=1.835 $X2=0 $Y2=0
cc_1100 N_A_705_367#_c_1260_p N_A_2345_367#_c_3327_n 0.01442f $X=13.245 $Y=1.98
+ $X2=0 $Y2=0
cc_1101 N_A_705_367#_c_1086_n N_A_2345_367#_c_3311_n 0.0147623f $X=14.2 $Y=1.87
+ $X2=0 $Y2=0
cc_1102 N_A_705_367#_c_1001_n N_Z_c_3375_n 5.97954e-19 $X=14.765 $Y=1.65 $X2=0
+ $Y2=0
cc_1103 N_A_705_367#_c_1028_n N_Z_c_3375_n 2.27616e-19 $X=14.37 $Y=1.665 $X2=0
+ $Y2=0
cc_1104 N_A_705_367#_c_1029_n N_Z_c_3375_n 5.28259e-19 $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_1105 N_A_705_367#_c_1031_n N_Z_c_3375_n 0.0121334f $X=14.68 $Y=1.665 $X2=0
+ $Y2=0
cc_1106 N_A_705_367#_c_1045_n N_Z_c_3379_n 0.00975003f $X=14.84 $Y=1.725 $X2=0
+ $Y2=0
cc_1107 N_A_705_367#_c_1003_n N_Z_c_3379_n 0.00163567f $X=15.195 $Y=1.65 $X2=0
+ $Y2=0
cc_1108 N_A_705_367#_c_1047_n N_Z_c_3379_n 0.00988676f $X=15.27 $Y=1.725 $X2=0
+ $Y2=0
cc_1109 N_A_705_367#_c_1031_n N_Z_c_3379_n 0.0091072f $X=14.68 $Y=1.665 $X2=0
+ $Y2=0
cc_1110 N_A_705_367#_c_1032_n N_Z_c_3379_n 0.00458049f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1111 N_A_705_367#_c_1045_n N_Z_c_3367_n 0.00107992f $X=14.84 $Y=1.725 $X2=0
+ $Y2=0
cc_1112 N_A_705_367#_c_1047_n N_Z_c_3367_n 0.00602501f $X=15.27 $Y=1.725 $X2=0
+ $Y2=0
cc_1113 N_A_705_367#_c_1004_n N_Z_c_3367_n 0.0088652f $X=15.625 $Y=1.65 $X2=0
+ $Y2=0
cc_1114 N_A_705_367#_c_1049_n N_Z_c_3367_n 0.00573605f $X=15.7 $Y=1.725 $X2=0
+ $Y2=0
cc_1115 N_A_705_367#_c_1051_n N_Z_c_3367_n 6.8716e-19 $X=16.13 $Y=1.725 $X2=0
+ $Y2=0
cc_1116 N_A_705_367#_c_1014_n N_Z_c_3367_n 0.00308303f $X=15.27 $Y=1.65 $X2=0
+ $Y2=0
cc_1117 N_A_705_367#_c_1015_n N_Z_c_3367_n 0.00328496f $X=15.7 $Y=1.65 $X2=0
+ $Y2=0
cc_1118 N_A_705_367#_c_1031_n N_Z_c_3367_n 0.00432657f $X=14.68 $Y=1.665 $X2=0
+ $Y2=0
cc_1119 N_A_705_367#_c_1032_n N_Z_c_3367_n 0.0265363f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1120 N_A_705_367#_c_1045_n N_Z_c_3393_n 8.58142e-19 $X=14.84 $Y=1.725 $X2=0
+ $Y2=0
cc_1121 N_A_705_367#_c_1047_n N_Z_c_3393_n 0.0105614f $X=15.27 $Y=1.725 $X2=0
+ $Y2=0
cc_1122 N_A_705_367#_c_1049_n N_Z_c_3393_n 0.0101966f $X=15.7 $Y=1.725 $X2=0
+ $Y2=0
cc_1123 N_A_705_367#_c_1051_n N_Z_c_3393_n 7.46996e-19 $X=16.13 $Y=1.725 $X2=0
+ $Y2=0
cc_1124 N_A_705_367#_c_1049_n N_Z_c_3368_n 0.0020244f $X=15.7 $Y=1.725 $X2=0
+ $Y2=0
cc_1125 N_A_705_367#_c_1051_n N_Z_c_3368_n 0.0182943f $X=16.13 $Y=1.725 $X2=0
+ $Y2=0
cc_1126 N_A_705_367#_c_1006_n N_Z_c_3368_n 0.0088652f $X=16.485 $Y=1.65 $X2=0
+ $Y2=0
cc_1127 N_A_705_367#_c_1053_n N_Z_c_3368_n 0.0182971f $X=16.56 $Y=1.725 $X2=0
+ $Y2=0
cc_1128 N_A_705_367#_c_1055_n N_Z_c_3368_n 0.00202491f $X=16.99 $Y=1.725 $X2=0
+ $Y2=0
cc_1129 N_A_705_367#_c_1016_n N_Z_c_3368_n 0.00328496f $X=16.13 $Y=1.65 $X2=0
+ $Y2=0
cc_1130 N_A_705_367#_c_1017_n N_Z_c_3368_n 0.00328496f $X=16.56 $Y=1.65 $X2=0
+ $Y2=0
cc_1131 N_A_705_367#_c_1032_n N_Z_c_3368_n 0.0269783f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1132 N_A_705_367#_c_1053_n N_Z_c_3369_n 0.00202491f $X=16.56 $Y=1.725 $X2=0
+ $Y2=0
cc_1133 N_A_705_367#_c_1055_n N_Z_c_3369_n 0.0182971f $X=16.99 $Y=1.725 $X2=0
+ $Y2=0
cc_1134 N_A_705_367#_c_1008_n N_Z_c_3369_n 0.0088652f $X=17.345 $Y=1.65 $X2=0
+ $Y2=0
cc_1135 N_A_705_367#_c_1057_n N_Z_c_3369_n 0.0182971f $X=17.42 $Y=1.725 $X2=0
+ $Y2=0
cc_1136 N_A_705_367#_c_1059_n N_Z_c_3369_n 0.00202491f $X=17.85 $Y=1.725 $X2=0
+ $Y2=0
cc_1137 N_A_705_367#_c_1018_n N_Z_c_3369_n 0.00328496f $X=16.99 $Y=1.65 $X2=0
+ $Y2=0
cc_1138 N_A_705_367#_c_1019_n N_Z_c_3369_n 0.00328496f $X=17.42 $Y=1.65 $X2=0
+ $Y2=0
cc_1139 N_A_705_367#_c_1032_n N_Z_c_3369_n 0.0269783f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1140 N_A_705_367#_c_1057_n N_Z_c_3370_n 0.00202491f $X=17.42 $Y=1.725 $X2=0
+ $Y2=0
cc_1141 N_A_705_367#_c_1059_n N_Z_c_3370_n 0.0182971f $X=17.85 $Y=1.725 $X2=0
+ $Y2=0
cc_1142 N_A_705_367#_c_1010_n N_Z_c_3370_n 0.0088652f $X=18.205 $Y=1.65 $X2=0
+ $Y2=0
cc_1143 N_A_705_367#_c_1061_n N_Z_c_3370_n 0.0182971f $X=18.28 $Y=1.725 $X2=0
+ $Y2=0
cc_1144 N_A_705_367#_c_1063_n N_Z_c_3370_n 0.00202491f $X=18.71 $Y=1.725 $X2=0
+ $Y2=0
cc_1145 N_A_705_367#_c_1020_n N_Z_c_3370_n 0.00328496f $X=17.85 $Y=1.65 $X2=0
+ $Y2=0
cc_1146 N_A_705_367#_c_1021_n N_Z_c_3370_n 0.00328496f $X=18.28 $Y=1.65 $X2=0
+ $Y2=0
cc_1147 N_A_705_367#_c_1032_n N_Z_c_3370_n 0.0269783f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1148 N_A_705_367#_c_1061_n N_Z_c_3371_n 0.00202491f $X=18.28 $Y=1.725 $X2=0
+ $Y2=0
cc_1149 N_A_705_367#_c_1063_n N_Z_c_3371_n 0.0182971f $X=18.71 $Y=1.725 $X2=0
+ $Y2=0
cc_1150 N_A_705_367#_c_1012_n N_Z_c_3371_n 0.0109356f $X=19.065 $Y=1.65 $X2=0
+ $Y2=0
cc_1151 N_A_705_367#_c_1065_n N_Z_c_3371_n 0.0180894f $X=19.14 $Y=1.725 $X2=0
+ $Y2=0
cc_1152 N_A_705_367#_c_1066_n N_Z_c_3371_n 0.00193435f $X=19.57 $Y=1.725 $X2=0
+ $Y2=0
cc_1153 N_A_705_367#_c_1022_n N_Z_c_3371_n 0.00346539f $X=18.71 $Y=1.65 $X2=0
+ $Y2=0
cc_1154 N_A_705_367#_c_1032_n N_Z_c_3371_n 0.0295962f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1155 N_A_705_367#_c_1034_n N_Z_c_3371_n 0.0293342f $X=19.345 $Y=1.51 $X2=0
+ $Y2=0
cc_1156 N_A_705_367#_c_1037_n N_Z_c_3371_n 0.00807773f $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1157 N_A_705_367#_c_1065_n N_Z_c_3372_n 0.00193435f $X=19.14 $Y=1.725 $X2=0
+ $Y2=0
cc_1158 N_A_705_367#_c_1066_n N_Z_c_3372_n 0.0180894f $X=19.57 $Y=1.725 $X2=0
+ $Y2=0
cc_1159 N_A_705_367#_c_1067_n N_Z_c_3372_n 0.0180894f $X=20 $Y=1.725 $X2=0 $Y2=0
cc_1160 N_A_705_367#_c_1068_n N_Z_c_3372_n 0.00193435f $X=20.43 $Y=1.725 $X2=0
+ $Y2=0
cc_1161 N_A_705_367#_c_1032_n N_Z_c_3372_n 0.0270023f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1162 N_A_705_367#_c_1034_n N_Z_c_3372_n 0.0285366f $X=19.345 $Y=1.51 $X2=0
+ $Y2=0
cc_1163 N_A_705_367#_c_1035_n N_Z_c_3372_n 0.0285366f $X=20.205 $Y=1.51 $X2=0
+ $Y2=0
cc_1164 N_A_705_367#_c_1037_n N_Z_c_3372_n 0.0256227f $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1165 N_A_705_367#_c_1067_n N_Z_c_3373_n 0.00193435f $X=20 $Y=1.725 $X2=0
+ $Y2=0
cc_1166 N_A_705_367#_c_1068_n N_Z_c_3373_n 0.0180894f $X=20.43 $Y=1.725 $X2=0
+ $Y2=0
cc_1167 N_A_705_367#_c_1069_n N_Z_c_3373_n 0.0180894f $X=20.86 $Y=1.725 $X2=0
+ $Y2=0
cc_1168 N_A_705_367#_c_1070_n N_Z_c_3373_n 0.00193435f $X=21.29 $Y=1.725 $X2=0
+ $Y2=0
cc_1169 N_A_705_367#_c_1032_n N_Z_c_3373_n 0.0270023f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1170 N_A_705_367#_c_1035_n N_Z_c_3373_n 0.0285366f $X=20.205 $Y=1.51 $X2=0
+ $Y2=0
cc_1171 N_A_705_367#_c_1036_n N_Z_c_3373_n 0.0285366f $X=21.065 $Y=1.51 $X2=0
+ $Y2=0
cc_1172 N_A_705_367#_c_1037_n N_Z_c_3373_n 0.0256227f $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1173 N_A_705_367#_c_1069_n N_Z_c_3374_n 0.00193435f $X=20.86 $Y=1.725 $X2=0
+ $Y2=0
cc_1174 N_A_705_367#_c_1070_n N_Z_c_3374_n 0.0180894f $X=21.29 $Y=1.725 $X2=0
+ $Y2=0
cc_1175 N_A_705_367#_c_1071_n N_Z_c_3374_n 0.0185428f $X=21.72 $Y=1.725 $X2=0
+ $Y2=0
cc_1176 N_A_705_367#_c_1072_n N_Z_c_3374_n 0.00239833f $X=22.15 $Y=1.725 $X2=0
+ $Y2=0
cc_1177 N_A_705_367#_c_1032_n N_Z_c_3374_n 0.0352521f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1178 N_A_705_367#_c_1036_n N_Z_c_3374_n 0.0285366f $X=21.065 $Y=1.51 $X2=0
+ $Y2=0
cc_1179 N_A_705_367#_c_1037_n N_Z_c_3374_n 0.0304401f $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1180 N_A_705_367#_c_1038_n N_Z_c_3374_n 0.0299743f $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1181 N_A_705_367#_c_1071_n N_Z_c_3454_n 0.00136857f $X=21.72 $Y=1.725 $X2=0
+ $Y2=0
cc_1182 N_A_705_367#_c_1072_n N_Z_c_3454_n 0.0128593f $X=22.15 $Y=1.725 $X2=0
+ $Y2=0
cc_1183 N_A_705_367#_c_1073_n N_Z_c_3454_n 0.0239079f $X=22.58 $Y=1.725 $X2=0
+ $Y2=0
cc_1184 N_A_705_367#_c_1032_n N_Z_c_3454_n 0.00101997f $X=22.285 $Y=1.665 $X2=0
+ $Y2=0
cc_1185 N_A_705_367#_c_1037_n N_Z_c_3454_n 6.13936e-19 $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1186 N_A_705_367#_c_1038_n N_Z_c_3454_n 0.0145361f $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1187 N_A_705_367#_c_1042_n N_Z_c_3460_n 0.00770204f $X=14.41 $Y=1.725 $X2=0
+ $Y2=0
cc_1188 N_A_705_367#_c_1045_n N_Z_c_3460_n 0.00357174f $X=14.84 $Y=1.725 $X2=0
+ $Y2=0
cc_1189 N_A_705_367#_c_1003_n N_Z_c_3460_n 4.88914e-19 $X=15.195 $Y=1.65 $X2=0
+ $Y2=0
cc_1190 N_A_705_367#_c_1047_n N_Z_c_3460_n 0.00338438f $X=15.27 $Y=1.725 $X2=0
+ $Y2=0
cc_1191 N_A_705_367#_c_1049_n N_Z_c_3460_n 0.00475577f $X=15.7 $Y=1.725 $X2=0
+ $Y2=0
cc_1192 N_A_705_367#_c_1005_n N_Z_c_3460_n 4.88914e-19 $X=16.055 $Y=1.65 $X2=0
+ $Y2=0
cc_1193 N_A_705_367#_c_1051_n N_Z_c_3460_n 0.00476607f $X=16.13 $Y=1.725 $X2=0
+ $Y2=0
cc_1194 N_A_705_367#_c_1053_n N_Z_c_3460_n 0.00476607f $X=16.56 $Y=1.725 $X2=0
+ $Y2=0
cc_1195 N_A_705_367#_c_1007_n N_Z_c_3460_n 4.88914e-19 $X=16.915 $Y=1.65 $X2=0
+ $Y2=0
cc_1196 N_A_705_367#_c_1055_n N_Z_c_3460_n 0.00476607f $X=16.99 $Y=1.725 $X2=0
+ $Y2=0
cc_1197 N_A_705_367#_c_1057_n N_Z_c_3460_n 0.00476607f $X=17.42 $Y=1.725 $X2=0
+ $Y2=0
cc_1198 N_A_705_367#_c_1009_n N_Z_c_3460_n 4.88914e-19 $X=17.775 $Y=1.65 $X2=0
+ $Y2=0
cc_1199 N_A_705_367#_c_1059_n N_Z_c_3460_n 0.00476607f $X=17.85 $Y=1.725 $X2=0
+ $Y2=0
cc_1200 N_A_705_367#_c_1061_n N_Z_c_3460_n 0.00476607f $X=18.28 $Y=1.725 $X2=0
+ $Y2=0
cc_1201 N_A_705_367#_c_1011_n N_Z_c_3460_n 4.88914e-19 $X=18.635 $Y=1.65 $X2=0
+ $Y2=0
cc_1202 N_A_705_367#_c_1063_n N_Z_c_3460_n 0.00482744f $X=18.71 $Y=1.725 $X2=0
+ $Y2=0
cc_1203 N_A_705_367#_c_1065_n N_Z_c_3460_n 0.00485104f $X=19.14 $Y=1.725 $X2=0
+ $Y2=0
cc_1204 N_A_705_367#_c_1066_n N_Z_c_3460_n 0.00485104f $X=19.57 $Y=1.725 $X2=0
+ $Y2=0
cc_1205 N_A_705_367#_c_1067_n N_Z_c_3460_n 0.00485104f $X=20 $Y=1.725 $X2=0
+ $Y2=0
cc_1206 N_A_705_367#_c_1068_n N_Z_c_3460_n 0.00485104f $X=20.43 $Y=1.725 $X2=0
+ $Y2=0
cc_1207 N_A_705_367#_c_1069_n N_Z_c_3460_n 0.00485104f $X=20.86 $Y=1.725 $X2=0
+ $Y2=0
cc_1208 N_A_705_367#_c_1070_n N_Z_c_3460_n 0.00485104f $X=21.29 $Y=1.725 $X2=0
+ $Y2=0
cc_1209 N_A_705_367#_c_1071_n N_Z_c_3460_n 0.00485104f $X=21.72 $Y=1.725 $X2=0
+ $Y2=0
cc_1210 N_A_705_367#_c_1072_n N_Z_c_3460_n 0.00453899f $X=22.15 $Y=1.725 $X2=0
+ $Y2=0
cc_1211 N_A_705_367#_c_1073_n N_Z_c_3460_n 8.0075e-19 $X=22.58 $Y=1.725 $X2=0
+ $Y2=0
cc_1212 N_A_705_367#_c_1028_n N_Z_c_3460_n 0.00162358f $X=14.37 $Y=1.665 $X2=0
+ $Y2=0
cc_1213 N_A_705_367#_c_1029_n N_Z_c_3460_n 0.791722f $X=14.5 $Y=1.665 $X2=0
+ $Y2=0
cc_1214 N_A_705_367#_c_1031_n N_Z_c_3460_n 0.00203371f $X=14.68 $Y=1.665 $X2=0
+ $Y2=0
cc_1215 N_A_705_367#_c_1034_n N_Z_c_3460_n 8.62013e-19 $X=19.345 $Y=1.51 $X2=0
+ $Y2=0
cc_1216 N_A_705_367#_c_1035_n N_Z_c_3460_n 8.62013e-19 $X=20.205 $Y=1.51 $X2=0
+ $Y2=0
cc_1217 N_A_705_367#_c_1036_n N_Z_c_3460_n 8.62013e-19 $X=21.065 $Y=1.51 $X2=0
+ $Y2=0
cc_1218 N_A_705_367#_c_1038_n N_Z_c_3460_n 0.00404212f $X=22.265 $Y=1.51 $X2=0
+ $Y2=0
cc_1219 N_A_705_367#_c_1047_n N_Z_c_3492_n 4.0679e-19 $X=15.27 $Y=1.725 $X2=0
+ $Y2=0
cc_1220 N_A_705_367#_c_1049_n N_Z_c_3492_n 0.0023483f $X=15.7 $Y=1.725 $X2=0
+ $Y2=0
cc_1221 N_A_705_367#_c_1051_n N_Z_c_3492_n 6.12528e-19 $X=16.13 $Y=1.725 $X2=0
+ $Y2=0
cc_1222 N_A_705_367#_c_1034_n N_VGND_c_3677_n 0.00626246f $X=19.345 $Y=1.51
+ $X2=0 $Y2=0
cc_1223 N_A_705_367#_c_1037_n N_VGND_c_3677_n 3.37033e-19 $X=22.265 $Y=1.51
+ $X2=0 $Y2=0
cc_1224 N_A_705_367#_c_1035_n N_VGND_c_3678_n 0.00626246f $X=20.205 $Y=1.51
+ $X2=0 $Y2=0
cc_1225 N_A_705_367#_c_1037_n N_VGND_c_3678_n 3.37033e-19 $X=22.265 $Y=1.51
+ $X2=0 $Y2=0
cc_1226 N_A_705_367#_c_1036_n N_VGND_c_3679_n 0.00626246f $X=21.065 $Y=1.51
+ $X2=0 $Y2=0
cc_1227 N_A_705_367#_c_1037_n N_VGND_c_3679_n 3.37033e-19 $X=22.265 $Y=1.51
+ $X2=0 $Y2=0
cc_1228 N_A_705_367#_M1014_g N_VGND_c_3688_n 0.00359964f $X=5.55 $Y=0.445 $X2=0
+ $Y2=0
cc_1229 N_A_705_367#_M1005_s N_VGND_c_3707_n 0.00225465f $X=14.03 $Y=0.235 $X2=0
+ $Y2=0
cc_1230 N_A_705_367#_M1014_g N_VGND_c_3707_n 0.00665534f $X=5.55 $Y=0.445 $X2=0
+ $Y2=0
cc_1231 N_A_705_367#_c_1027_n N_A_2519_47#_c_3956_n 0.00794156f $X=14.222
+ $Y=1.095 $X2=0 $Y2=0
cc_1232 N_A_705_367#_M1005_s N_A_2519_47#_c_3961_n 0.00340092f $X=14.03 $Y=0.235
+ $X2=0 $Y2=0
cc_1233 N_A_705_367#_c_1276_p N_A_2519_47#_c_3961_n 0.0158394f $X=14.17 $Y=0.815
+ $X2=0 $Y2=0
cc_1234 N_A_705_367#_c_1001_n N_A_2519_47#_c_3959_n 0.00162515f $X=14.765
+ $Y=1.65 $X2=0 $Y2=0
cc_1235 N_A_705_367#_c_1276_p N_A_2519_47#_c_3959_n 0.0361629f $X=14.17 $Y=0.815
+ $X2=0 $Y2=0
cc_1236 N_A_705_367#_c_1031_n N_A_2519_47#_c_3959_n 0.00580564f $X=14.68
+ $Y=1.665 $X2=0 $Y2=0
cc_1237 N_A_407_491#_c_1564_n N_A_896_367#_M1014_d 0.00653876f $X=6.525 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_1238 N_A_407_491#_c_1560_n N_A_896_367#_c_1764_n 0.0217278f $X=7.355 $Y=1.26
+ $X2=0 $Y2=0
cc_1239 N_A_407_491#_c_1566_n N_A_896_367#_c_1764_n 8.52481e-19 $X=7.395
+ $Y=0.935 $X2=0 $Y2=0
cc_1240 N_A_407_491#_c_1554_n N_A_896_367#_c_1766_n 0.0217278f $X=7.96 $Y=1.26
+ $X2=0 $Y2=0
cc_1241 N_A_407_491#_c_1559_n N_A_896_367#_c_1767_n 0.00583548f $X=6.79 $Y=0.67
+ $X2=0 $Y2=0
cc_1242 N_A_407_491#_c_1563_n N_A_896_367#_c_1767_n 0.0129699f $X=5.285 $Y=0.73
+ $X2=0 $Y2=0
cc_1243 N_A_407_491#_c_1564_n N_A_896_367#_c_1767_n 0.0489967f $X=6.525 $Y=0.35
+ $X2=0 $Y2=0
cc_1244 N_A_407_491#_c_1565_n N_A_896_367#_c_1767_n 0.0169735f $X=6.61 $Y=0.67
+ $X2=0 $Y2=0
cc_1245 N_A_407_491#_c_1550_n N_A_896_367#_c_1768_n 0.00198969f $X=6.865
+ $Y=1.185 $X2=0 $Y2=0
cc_1246 N_A_407_491#_c_1559_n N_A_896_367#_c_1768_n 5.33128e-19 $X=6.79 $Y=0.67
+ $X2=0 $Y2=0
cc_1247 N_A_407_491#_c_1565_n N_A_896_367#_c_1768_n 0.00248455f $X=6.61 $Y=0.67
+ $X2=0 $Y2=0
cc_1248 N_A_407_491#_c_1567_n N_A_896_367#_c_1768_n 0.0143581f $X=6.695 $Y=0.935
+ $X2=0 $Y2=0
cc_1249 N_A_407_491#_c_1551_n N_A_896_367#_c_1769_n 0.0159012f $X=7.28 $Y=1.26
+ $X2=0 $Y2=0
cc_1250 N_A_407_491#_c_1552_n N_A_896_367#_c_1769_n 0.00743002f $X=6.94 $Y=1.26
+ $X2=0 $Y2=0
cc_1251 N_A_407_491#_c_1559_n N_A_896_367#_c_1769_n 0.00113735f $X=6.79 $Y=0.67
+ $X2=0 $Y2=0
cc_1252 N_A_407_491#_c_1566_n N_A_896_367#_c_1769_n 0.0367585f $X=7.395 $Y=0.935
+ $X2=0 $Y2=0
cc_1253 N_A_407_491#_c_1567_n N_A_896_367#_c_1769_n 0.0130548f $X=6.695 $Y=0.935
+ $X2=0 $Y2=0
cc_1254 N_A_407_491#_c_1551_n N_A_896_367#_c_1772_n 0.0217278f $X=7.28 $Y=1.26
+ $X2=0 $Y2=0
cc_1255 N_A_407_491#_c_1566_n N_A_896_367#_c_1772_n 5.85059e-19 $X=7.395
+ $Y=0.935 $X2=0 $Y2=0
cc_1256 N_A_407_491#_c_1566_n N_A_1486_47#_M1038_d 0.00224952f $X=7.395 $Y=0.935
+ $X2=-0.19 $Y2=-0.245
cc_1257 N_A_407_491#_c_1648_p N_A_1486_47#_M1038_d 0.00452263f $X=7.48 $Y=0.85
+ $X2=-0.19 $Y2=-0.245
cc_1258 N_A_407_491#_c_1649_p N_A_1486_47#_M1038_d 0.0130392f $X=8.075 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_1259 N_A_407_491#_c_1650_p N_A_1486_47#_M1038_d 7.79781e-19 $X=7.565 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_1260 N_A_407_491#_c_1568_n N_A_1486_47#_M1003_d 0.0105144f $X=9.985 $Y=0.74
+ $X2=0 $Y2=0
cc_1261 N_A_407_491#_M1020_g N_A_1486_47#_M1065_g 0.0222649f $X=10.24 $Y=0.445
+ $X2=0 $Y2=0
cc_1262 N_A_407_491#_M1018_g N_A_1486_47#_c_1941_n 0.00642768f $X=10.09 $Y=2.285
+ $X2=0 $Y2=0
cc_1263 N_A_407_491#_M1018_g N_A_1486_47#_c_1942_n 0.0809517f $X=10.09 $Y=2.285
+ $X2=0 $Y2=0
cc_1264 N_A_407_491#_c_1553_n N_A_1486_47#_c_2028_n 0.00107255f $X=7.355
+ $Y=1.185 $X2=0 $Y2=0
cc_1265 N_A_407_491#_c_1554_n N_A_1486_47#_c_2028_n 6.26978e-19 $X=7.96 $Y=1.26
+ $X2=0 $Y2=0
cc_1266 N_A_407_491#_c_1566_n N_A_1486_47#_c_2028_n 0.0117969f $X=7.395 $Y=0.935
+ $X2=0 $Y2=0
cc_1267 N_A_407_491#_c_1648_p N_A_1486_47#_c_2028_n 0.0177587f $X=7.48 $Y=0.85
+ $X2=0 $Y2=0
cc_1268 N_A_407_491#_c_1649_p N_A_1486_47#_c_2028_n 0.0122122f $X=8.075 $Y=0.35
+ $X2=0 $Y2=0
cc_1269 N_A_407_491#_c_1554_n N_A_1486_47#_c_1948_n 0.0112967f $X=7.96 $Y=1.26
+ $X2=0 $Y2=0
cc_1270 N_A_407_491#_c_1556_n N_A_1486_47#_c_1949_n 0.0016127f $X=10.09 $Y=1.33
+ $X2=0 $Y2=0
cc_1271 N_A_407_491#_c_1568_n N_A_1486_47#_c_1949_n 0.0915402f $X=9.985 $Y=0.74
+ $X2=0 $Y2=0
cc_1272 N_A_407_491#_c_1569_n N_A_1486_47#_c_1949_n 0.0110821f $X=10.15 $Y=1.16
+ $X2=0 $Y2=0
cc_1273 N_A_407_491#_c_1553_n N_A_1486_47#_c_1950_n 0.00421962f $X=7.355
+ $Y=1.185 $X2=0 $Y2=0
cc_1274 N_A_407_491#_c_1554_n N_A_1486_47#_c_1950_n 0.00727057f $X=7.96 $Y=1.26
+ $X2=0 $Y2=0
cc_1275 N_A_407_491#_c_1555_n N_A_1486_47#_c_1950_n 0.0118963f $X=8.035 $Y=1.185
+ $X2=0 $Y2=0
cc_1276 N_A_407_491#_c_1566_n N_A_1486_47#_c_1950_n 0.00216387f $X=7.395
+ $Y=0.935 $X2=0 $Y2=0
cc_1277 N_A_407_491#_c_1649_p N_A_1486_47#_c_1950_n 0.00299905f $X=8.075 $Y=0.35
+ $X2=0 $Y2=0
cc_1278 N_A_407_491#_c_1669_p N_A_1486_47#_c_1950_n 0.0089265f $X=8.245 $Y=0.74
+ $X2=0 $Y2=0
cc_1279 N_A_407_491#_c_1556_n N_A_1486_47#_c_1951_n 0.00307699f $X=10.09 $Y=1.33
+ $X2=0 $Y2=0
cc_1280 N_A_407_491#_M1018_g N_A_1486_47#_c_1951_n 0.00214297f $X=10.09 $Y=2.285
+ $X2=0 $Y2=0
cc_1281 N_A_407_491#_c_1568_n N_A_1486_47#_c_1951_n 0.00867852f $X=9.985 $Y=0.74
+ $X2=0 $Y2=0
cc_1282 N_A_407_491#_c_1569_n N_A_1486_47#_c_1951_n 0.0265518f $X=10.15 $Y=1.16
+ $X2=0 $Y2=0
cc_1283 N_A_407_491#_c_1556_n N_A_1486_47#_c_1952_n 7.49848e-19 $X=10.09 $Y=1.33
+ $X2=0 $Y2=0
cc_1284 N_A_407_491#_M1018_g N_A_1486_47#_c_1952_n 7.01421e-19 $X=10.09 $Y=2.285
+ $X2=0 $Y2=0
cc_1285 N_A_407_491#_c_1568_n N_A_1486_47#_c_1952_n 0.00141077f $X=9.985 $Y=0.74
+ $X2=0 $Y2=0
cc_1286 N_A_407_491#_c_1569_n N_A_1486_47#_c_1952_n 0.00123014f $X=10.15 $Y=1.16
+ $X2=0 $Y2=0
cc_1287 N_A_407_491#_c_1556_n N_A_1486_47#_c_1954_n 7.14409e-19 $X=10.09 $Y=1.33
+ $X2=0 $Y2=0
cc_1288 N_A_407_491#_M1018_g N_A_1486_47#_c_1954_n 6.64757e-19 $X=10.09 $Y=2.285
+ $X2=0 $Y2=0
cc_1289 N_A_407_491#_c_1569_n N_A_1486_47#_c_1954_n 0.00137314f $X=10.15 $Y=1.16
+ $X2=0 $Y2=0
cc_1290 N_A_407_491#_c_1556_n N_A_1486_47#_c_1957_n 0.00463379f $X=10.09 $Y=1.33
+ $X2=0 $Y2=0
cc_1291 N_A_407_491#_c_1569_n N_A_1486_47#_c_1957_n 0.00773658f $X=10.15 $Y=1.16
+ $X2=0 $Y2=0
cc_1292 N_A_407_491#_c_1556_n N_A_1486_47#_c_1958_n 0.00175188f $X=10.09 $Y=1.33
+ $X2=0 $Y2=0
cc_1293 N_A_407_491#_M1018_g N_A_1486_47#_c_1958_n 0.00464034f $X=10.09 $Y=2.285
+ $X2=0 $Y2=0
cc_1294 N_A_407_491#_c_1569_n N_A_1486_47#_c_1958_n 0.0244555f $X=10.15 $Y=1.16
+ $X2=0 $Y2=0
cc_1295 N_A_407_491#_c_1556_n N_A_1486_47#_c_1959_n 0.0214821f $X=10.09 $Y=1.33
+ $X2=0 $Y2=0
cc_1296 N_A_407_491#_c_1569_n N_A_1486_47#_c_1959_n 4.35733e-19 $X=10.15 $Y=1.16
+ $X2=0 $Y2=0
cc_1297 N_A_407_491#_c_1555_n N_A_M1003_g 0.0174883f $X=8.035 $Y=1.185 $X2=0
+ $Y2=0
cc_1298 N_A_407_491#_c_1689_p N_A_M1003_g 0.00268143f $X=8.16 $Y=0.655 $X2=0
+ $Y2=0
cc_1299 N_A_407_491#_c_1568_n N_A_M1003_g 0.0134897f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1300 N_A_407_491#_c_1556_n N_A_M1071_g 0.00883235f $X=10.09 $Y=1.33 $X2=0
+ $Y2=0
cc_1301 N_A_407_491#_M1020_g N_A_M1071_g 0.00679714f $X=10.24 $Y=0.445 $X2=0
+ $Y2=0
cc_1302 N_A_407_491#_c_1568_n N_A_M1071_g 0.0139865f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1303 N_A_407_491#_c_1569_n N_A_M1071_g 3.38257e-19 $X=10.15 $Y=1.16 $X2=0
+ $Y2=0
cc_1304 N_A_407_491#_c_1570_n N_A_M1071_g 0.0027251f $X=10.15 $Y=0.995 $X2=0
+ $Y2=0
cc_1305 N_A_407_491#_M1018_g N_A_c_2284_n 0.00870829f $X=10.09 $Y=2.285 $X2=0
+ $Y2=0
cc_1306 N_A_407_491#_M1018_g N_A_c_2272_n 0.0328992f $X=10.09 $Y=2.285 $X2=0
+ $Y2=0
cc_1307 N_A_407_491#_M1020_g N_A_2063_47#_c_2484_n 0.00142946f $X=10.24 $Y=0.445
+ $X2=0 $Y2=0
cc_1308 N_A_407_491#_c_1568_n N_A_2063_47#_c_2484_n 0.0130716f $X=9.985 $Y=0.74
+ $X2=0 $Y2=0
cc_1309 N_A_407_491#_M1018_g N_A_2063_47#_c_2495_n 0.00201332f $X=10.09 $Y=2.285
+ $X2=0 $Y2=0
cc_1310 N_A_407_491#_M1018_g N_A_2063_47#_c_2496_n 4.97653e-19 $X=10.09 $Y=2.285
+ $X2=0 $Y2=0
cc_1311 N_A_407_491#_M1018_g N_VPWR_c_2632_n 0.0200637f $X=10.09 $Y=2.285 $X2=0
+ $Y2=0
cc_1312 N_A_407_491#_c_1569_n N_VPWR_c_2632_n 8.02218e-19 $X=10.15 $Y=1.16 $X2=0
+ $Y2=0
cc_1313 N_A_407_491#_c_1572_n N_VPWR_c_2667_n 0.0210467f $X=2.16 $Y=2.61 $X2=0
+ $Y2=0
cc_1314 N_A_407_491#_M1035_s N_VPWR_c_2627_n 0.00110569f $X=2.035 $Y=2.455 $X2=0
+ $Y2=0
cc_1315 N_A_407_491#_c_1572_n N_VPWR_c_2627_n 0.00303861f $X=2.16 $Y=2.61 $X2=0
+ $Y2=0
cc_1316 N_A_407_491#_c_1573_n N_KAPWR_M1035_d 0.00477266f $X=3.335 $Y=2.185
+ $X2=-0.19 $Y2=-0.245
cc_1317 N_A_407_491#_M1018_g KAPWR 0.00321232f $X=10.09 $Y=2.285 $X2=0 $Y2=0
cc_1318 N_A_407_491#_c_1572_n KAPWR 0.02777f $X=2.16 $Y=2.61 $X2=0 $Y2=0
cc_1319 N_A_407_491#_c_1573_n KAPWR 0.00822444f $X=3.335 $Y=2.185 $X2=0 $Y2=0
cc_1320 N_A_407_491#_c_1572_n N_KAPWR_c_3047_n 0.0281622f $X=2.16 $Y=2.61 $X2=0
+ $Y2=0
cc_1321 N_A_407_491#_c_1573_n N_KAPWR_c_3047_n 0.060236f $X=3.335 $Y=2.185 $X2=0
+ $Y2=0
cc_1322 N_A_407_491#_c_1563_n N_VGND_M1063_d 0.0145196f $X=5.285 $Y=0.73 $X2=0
+ $Y2=0
cc_1323 N_A_407_491#_c_1566_n N_VGND_M1038_s 0.00398869f $X=7.395 $Y=0.935 $X2=0
+ $Y2=0
cc_1324 N_A_407_491#_c_1649_p N_VGND_M1050_s 0.00243741f $X=8.075 $Y=0.35 $X2=0
+ $Y2=0
cc_1325 N_A_407_491#_c_1689_p N_VGND_M1050_s 0.00312021f $X=8.16 $Y=0.655 $X2=0
+ $Y2=0
cc_1326 N_A_407_491#_c_1568_n N_VGND_M1050_s 0.0123548f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1327 N_A_407_491#_c_1669_p N_VGND_M1050_s 8.6018e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_1328 N_A_407_491#_c_1568_n N_VGND_M1071_s 0.00640006f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1329 N_A_407_491#_c_1561_n N_VGND_c_3666_n 0.0361421f $X=3.42 $Y=0.815 $X2=0
+ $Y2=0
cc_1330 N_A_407_491#_c_1562_n N_VGND_c_3666_n 0.0108617f $X=3.42 $Y=2.1 $X2=0
+ $Y2=0
cc_1331 N_A_407_491#_c_1553_n N_VGND_c_3667_n 0.0061012f $X=7.355 $Y=1.185 $X2=0
+ $Y2=0
cc_1332 N_A_407_491#_c_1559_n N_VGND_c_3667_n 0.00205946f $X=6.79 $Y=0.67 $X2=0
+ $Y2=0
cc_1333 N_A_407_491#_c_1564_n N_VGND_c_3667_n 0.0104094f $X=6.525 $Y=0.35 $X2=0
+ $Y2=0
cc_1334 N_A_407_491#_c_1565_n N_VGND_c_3667_n 0.012722f $X=6.61 $Y=0.67 $X2=0
+ $Y2=0
cc_1335 N_A_407_491#_c_1566_n N_VGND_c_3667_n 0.0197903f $X=7.395 $Y=0.935 $X2=0
+ $Y2=0
cc_1336 N_A_407_491#_c_1555_n N_VGND_c_3668_n 0.00327414f $X=8.035 $Y=1.185
+ $X2=0 $Y2=0
cc_1337 N_A_407_491#_c_1649_p N_VGND_c_3668_n 0.0145956f $X=8.075 $Y=0.35 $X2=0
+ $Y2=0
cc_1338 N_A_407_491#_c_1689_p N_VGND_c_3668_n 0.00227704f $X=8.16 $Y=0.655 $X2=0
+ $Y2=0
cc_1339 N_A_407_491#_c_1568_n N_VGND_c_3668_n 0.0212616f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1340 N_A_407_491#_M1020_g N_VGND_c_3669_n 0.00486043f $X=10.24 $Y=0.445 $X2=0
+ $Y2=0
cc_1341 N_A_407_491#_M1020_g N_VGND_c_3670_n 5.71707e-19 $X=10.24 $Y=0.445 $X2=0
+ $Y2=0
cc_1342 N_A_407_491#_c_1563_n N_VGND_c_3686_n 0.103441f $X=5.285 $Y=0.73 $X2=0
+ $Y2=0
cc_1343 N_A_407_491#_c_1561_n N_VGND_c_3687_n 0.0177128f $X=3.42 $Y=0.815 $X2=0
+ $Y2=0
cc_1344 N_A_407_491#_c_1563_n N_VGND_c_3687_n 0.00247188f $X=5.285 $Y=0.73 $X2=0
+ $Y2=0
cc_1345 N_A_407_491#_c_1559_n N_VGND_c_3688_n 0.0071072f $X=6.79 $Y=0.67 $X2=0
+ $Y2=0
cc_1346 N_A_407_491#_c_1563_n N_VGND_c_3688_n 0.00262235f $X=5.285 $Y=0.73 $X2=0
+ $Y2=0
cc_1347 N_A_407_491#_c_1564_n N_VGND_c_3688_n 0.0735058f $X=6.525 $Y=0.35 $X2=0
+ $Y2=0
cc_1348 N_A_407_491#_c_1739_p N_VGND_c_3688_n 0.0087245f $X=5.455 $Y=0.35 $X2=0
+ $Y2=0
cc_1349 N_A_407_491#_c_1553_n N_VGND_c_3690_n 0.00532738f $X=7.355 $Y=1.185
+ $X2=0 $Y2=0
cc_1350 N_A_407_491#_c_1555_n N_VGND_c_3690_n 0.00359916f $X=8.035 $Y=1.185
+ $X2=0 $Y2=0
cc_1351 N_A_407_491#_c_1649_p N_VGND_c_3690_n 0.0378378f $X=8.075 $Y=0.35 $X2=0
+ $Y2=0
cc_1352 N_A_407_491#_c_1650_p N_VGND_c_3690_n 0.0093013f $X=7.565 $Y=0.35 $X2=0
+ $Y2=0
cc_1353 N_A_407_491#_c_1568_n N_VGND_c_3690_n 0.00282537f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1354 N_A_407_491#_M1063_s N_VGND_c_3707_n 0.00215817f $X=3.225 $Y=0.235 $X2=0
+ $Y2=0
cc_1355 N_A_407_491#_c_1553_n N_VGND_c_3707_n 0.00813154f $X=7.355 $Y=1.185
+ $X2=0 $Y2=0
cc_1356 N_A_407_491#_c_1555_n N_VGND_c_3707_n 0.00665845f $X=8.035 $Y=1.185
+ $X2=0 $Y2=0
cc_1357 N_A_407_491#_M1020_g N_VGND_c_3707_n 0.0083335f $X=10.24 $Y=0.445 $X2=0
+ $Y2=0
cc_1358 N_A_407_491#_c_1559_n N_VGND_c_3707_n 0.00730016f $X=6.79 $Y=0.67 $X2=0
+ $Y2=0
cc_1359 N_A_407_491#_c_1561_n N_VGND_c_3707_n 0.0120687f $X=3.42 $Y=0.815 $X2=0
+ $Y2=0
cc_1360 N_A_407_491#_c_1563_n N_VGND_c_3707_n 0.0145779f $X=5.285 $Y=0.73 $X2=0
+ $Y2=0
cc_1361 N_A_407_491#_c_1564_n N_VGND_c_3707_n 0.045872f $X=6.525 $Y=0.35 $X2=0
+ $Y2=0
cc_1362 N_A_407_491#_c_1739_p N_VGND_c_3707_n 0.00654039f $X=5.455 $Y=0.35 $X2=0
+ $Y2=0
cc_1363 N_A_407_491#_c_1566_n N_VGND_c_3707_n 0.0148749f $X=7.395 $Y=0.935 $X2=0
+ $Y2=0
cc_1364 N_A_407_491#_c_1649_p N_VGND_c_3707_n 0.0249084f $X=8.075 $Y=0.35 $X2=0
+ $Y2=0
cc_1365 N_A_407_491#_c_1650_p N_VGND_c_3707_n 0.00641662f $X=7.565 $Y=0.35 $X2=0
+ $Y2=0
cc_1366 N_A_407_491#_c_1568_n N_VGND_c_3707_n 0.0274073f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1367 N_A_407_491#_c_1568_n N_VGND_c_3709_n 0.0100997f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1368 N_A_407_491#_c_1556_n N_VGND_c_3710_n 5.58057e-19 $X=10.09 $Y=1.33 $X2=0
+ $Y2=0
cc_1369 N_A_407_491#_M1020_g N_VGND_c_3710_n 0.00814187f $X=10.24 $Y=0.445 $X2=0
+ $Y2=0
cc_1370 N_A_407_491#_c_1568_n N_VGND_c_3710_n 0.0484577f $X=9.985 $Y=0.74 $X2=0
+ $Y2=0
cc_1371 N_A_407_491#_c_1569_n N_VGND_c_3710_n 9.36914e-19 $X=10.15 $Y=1.16 $X2=0
+ $Y2=0
cc_1372 N_A_407_491#_c_1739_p A_1053_47# 9.53517e-19 $X=5.455 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_1373 N_A_896_367#_c_1774_n N_A_1486_47#_c_1948_n 0.00335423f $X=7.8 $Y=1.725
+ $X2=0 $Y2=0
cc_1374 N_A_896_367#_c_1765_n N_A_1486_47#_c_1948_n 0.0139951f $X=8.155 $Y=1.65
+ $X2=0 $Y2=0
cc_1375 N_A_896_367#_c_1776_n N_A_1486_47#_c_1948_n 0.00335423f $X=8.23 $Y=1.725
+ $X2=0 $Y2=0
cc_1376 N_A_896_367#_c_1765_n N_A_1486_47#_c_1949_n 0.00603375f $X=8.155 $Y=1.65
+ $X2=0 $Y2=0
cc_1377 N_A_896_367#_c_1766_n N_A_1486_47#_c_1950_n 0.00108865f $X=7.8 $Y=1.65
+ $X2=0 $Y2=0
cc_1378 N_A_896_367#_c_1769_n N_A_1486_47#_c_1950_n 7.94705e-19 $X=6.97 $Y=1.285
+ $X2=0 $Y2=0
cc_1379 N_A_896_367#_c_1776_n N_A_c_2281_n 0.0129622f $X=8.23 $Y=1.725 $X2=-0.19
+ $Y2=-0.245
cc_1380 N_A_896_367#_c_1765_n N_A_c_2272_n 0.0129622f $X=8.155 $Y=1.65 $X2=0
+ $Y2=0
cc_1381 N_A_896_367#_c_1778_n N_VPWR_M1049_s 0.00441857f $X=6.195 $Y=2.41 $X2=0
+ $Y2=0
cc_1382 N_A_896_367#_c_1778_n N_VPWR_c_2629_n 0.0193944f $X=6.195 $Y=2.41 $X2=0
+ $Y2=0
cc_1383 N_A_896_367#_c_1809_n N_VPWR_c_2629_n 0.00922356f $X=6.36 $Y=2.41 $X2=0
+ $Y2=0
cc_1384 N_A_896_367#_c_1779_n N_VPWR_c_2630_n 0.0171884f $X=6.97 $Y=2.17 $X2=0
+ $Y2=0
cc_1385 N_A_896_367#_c_1781_n N_VPWR_c_2630_n 0.0256862f $X=6.36 $Y=2.17 $X2=0
+ $Y2=0
cc_1386 N_A_896_367#_c_1809_n N_VPWR_c_2648_n 0.0177952f $X=6.36 $Y=2.41 $X2=0
+ $Y2=0
cc_1387 N_A_896_367#_c_1884_p N_VPWR_c_2667_n 0.0134452f $X=4.62 $Y=2.565 $X2=0
+ $Y2=0
cc_1388 N_A_896_367#_c_1774_n N_VPWR_c_2668_n 0.0035993f $X=7.8 $Y=1.725 $X2=0
+ $Y2=0
cc_1389 N_A_896_367#_c_1776_n N_VPWR_c_2668_n 0.0035993f $X=8.23 $Y=1.725 $X2=0
+ $Y2=0
cc_1390 N_A_896_367#_M1036_s N_VPWR_c_2627_n 0.00124018f $X=4.48 $Y=1.835 $X2=0
+ $Y2=0
cc_1391 N_A_896_367#_M1057_d N_VPWR_c_2627_n 0.00113524f $X=6.22 $Y=2.255 $X2=0
+ $Y2=0
cc_1392 N_A_896_367#_c_1774_n N_VPWR_c_2627_n 0.00605454f $X=7.8 $Y=1.725 $X2=0
+ $Y2=0
cc_1393 N_A_896_367#_c_1776_n N_VPWR_c_2627_n 0.00478018f $X=8.23 $Y=1.725 $X2=0
+ $Y2=0
cc_1394 N_A_896_367#_c_1884_p N_VPWR_c_2627_n 0.00215193f $X=4.62 $Y=2.565 $X2=0
+ $Y2=0
cc_1395 N_A_896_367#_c_1809_n N_VPWR_c_2627_n 0.00302007f $X=6.36 $Y=2.41 $X2=0
+ $Y2=0
cc_1396 N_A_896_367#_c_1778_n N_KAPWR_M1066_d 0.00560077f $X=6.195 $Y=2.41 $X2=0
+ $Y2=0
cc_1397 N_A_896_367#_M1036_s KAPWR 5.22398e-19 $X=4.48 $Y=1.835 $X2=0 $Y2=0
cc_1398 N_A_896_367#_c_1774_n KAPWR 0.00303402f $X=7.8 $Y=1.725 $X2=0 $Y2=0
cc_1399 N_A_896_367#_c_1776_n KAPWR 0.00303402f $X=8.23 $Y=1.725 $X2=0 $Y2=0
cc_1400 N_A_896_367#_c_1884_p KAPWR 0.0208779f $X=4.62 $Y=2.565 $X2=0 $Y2=0
cc_1401 N_A_896_367#_c_1778_n KAPWR 0.0269087f $X=6.195 $Y=2.41 $X2=0 $Y2=0
cc_1402 N_A_896_367#_c_1779_n KAPWR 0.0125073f $X=6.97 $Y=2.17 $X2=0 $Y2=0
cc_1403 N_A_896_367#_c_1809_n KAPWR 0.0301183f $X=6.36 $Y=2.41 $X2=0 $Y2=0
cc_1404 N_A_896_367#_c_1795_n N_KAPWR_c_3065_n 0.0117665f $X=4.62 $Y=2.225 $X2=0
+ $Y2=0
cc_1405 N_A_896_367#_c_1884_p N_KAPWR_c_3048_n 0.0166469f $X=4.62 $Y=2.565 $X2=0
+ $Y2=0
cc_1406 N_A_896_367#_c_1778_n N_KAPWR_c_3048_n 0.0184133f $X=6.195 $Y=2.41 $X2=0
+ $Y2=0
cc_1407 N_A_896_367#_c_1778_n A_1172_451# 0.00286996f $X=6.195 $Y=2.41 $X2=-0.19
+ $Y2=-0.245
cc_1408 N_A_896_367#_c_1774_n N_A_1492_367#_c_3248_n 6.00691e-19 $X=7.8 $Y=1.725
+ $X2=0 $Y2=0
cc_1409 N_A_896_367#_c_1764_n N_A_1492_367#_c_3237_n 0.00937288f $X=7.725
+ $Y=1.65 $X2=0 $Y2=0
cc_1410 N_A_896_367#_c_1774_n N_A_1492_367#_c_3237_n 0.013915f $X=7.8 $Y=1.725
+ $X2=0 $Y2=0
cc_1411 N_A_896_367#_c_1776_n N_A_1492_367#_c_3237_n 8.63529e-19 $X=8.23
+ $Y=1.725 $X2=0 $Y2=0
cc_1412 N_A_896_367#_c_1779_n N_A_1492_367#_c_3237_n 0.0098661f $X=6.97 $Y=2.17
+ $X2=0 $Y2=0
cc_1413 N_A_896_367#_c_1771_n N_A_1492_367#_c_3237_n 0.0132278f $X=7.135 $Y=1.74
+ $X2=0 $Y2=0
cc_1414 N_A_896_367#_c_1772_n N_A_1492_367#_c_3237_n 7.98572e-19 $X=7.135
+ $Y=1.65 $X2=0 $Y2=0
cc_1415 N_A_896_367#_c_1774_n N_A_1492_367#_c_3255_n 0.00807446f $X=7.8 $Y=1.725
+ $X2=0 $Y2=0
cc_1416 N_A_896_367#_c_1776_n N_A_1492_367#_c_3255_n 0.00802789f $X=8.23
+ $Y=1.725 $X2=0 $Y2=0
cc_1417 N_A_896_367#_c_1776_n N_A_1492_367#_c_3238_n 0.0060471f $X=8.23 $Y=1.725
+ $X2=0 $Y2=0
cc_1418 N_A_896_367#_c_1774_n N_A_1492_367#_c_3258_n 6.16883e-19 $X=7.8 $Y=1.725
+ $X2=0 $Y2=0
cc_1419 N_A_896_367#_c_1776_n N_A_1492_367#_c_3258_n 0.00578295f $X=8.23
+ $Y=1.725 $X2=0 $Y2=0
cc_1420 N_A_896_367#_c_1776_n N_A_1492_367#_c_3260_n 0.00182707f $X=8.23
+ $Y=1.725 $X2=0 $Y2=0
cc_1421 N_A_896_367#_M1014_d N_VGND_c_3707_n 0.00266576f $X=5.625 $Y=0.235 $X2=0
+ $Y2=0
cc_1422 N_A_1486_47#_c_1948_n N_A_M1003_g 0.0021851f $X=8.015 $Y=1.98 $X2=0
+ $Y2=0
cc_1423 N_A_1486_47#_c_1949_n N_A_M1003_g 0.0136333f $X=9.455 $Y=1.08 $X2=0
+ $Y2=0
cc_1424 N_A_1486_47#_c_1950_n N_A_M1003_g 2.90194e-19 $X=8.11 $Y=1.11 $X2=0
+ $Y2=0
cc_1425 N_A_1486_47#_c_1952_n N_A_M1003_g 0.00103507f $X=9.745 $Y=1.295 $X2=0
+ $Y2=0
cc_1426 N_A_1486_47#_c_1957_n N_A_M1003_g 0.00167293f $X=9.6 $Y=1.295 $X2=0
+ $Y2=0
cc_1427 N_A_1486_47#_c_1949_n N_A_M1071_g 0.0121466f $X=9.455 $Y=1.08 $X2=0
+ $Y2=0
cc_1428 N_A_1486_47#_c_1952_n N_A_M1071_g 0.00440528f $X=9.745 $Y=1.295 $X2=0
+ $Y2=0
cc_1429 N_A_1486_47#_c_1957_n N_A_M1071_g 0.00866095f $X=9.6 $Y=1.295 $X2=0
+ $Y2=0
cc_1430 N_A_1486_47#_M1068_g N_A_c_2284_n 0.00871667f $X=10.45 $Y=2.285 $X2=0
+ $Y2=0
cc_1431 N_A_1486_47#_M1065_g N_A_c_2265_n 0.0067428f $X=10.67 $Y=0.445 $X2=0
+ $Y2=0
cc_1432 N_A_1486_47#_c_1953_n N_A_c_2266_n 0.00288109f $X=14.92 $Y=1.295 $X2=0
+ $Y2=0
cc_1433 N_A_1486_47#_c_1953_n N_A_M1007_g 0.00205883f $X=14.92 $Y=1.295 $X2=0
+ $Y2=0
cc_1434 N_A_1486_47#_c_1953_n N_A_M1041_g 0.00194256f $X=14.92 $Y=1.295 $X2=0
+ $Y2=0
cc_1435 N_A_1486_47#_c_1948_n N_A_c_2272_n 0.00599912f $X=8.015 $Y=1.98 $X2=0
+ $Y2=0
cc_1436 N_A_1486_47#_c_1949_n N_A_c_2272_n 0.0156542f $X=9.455 $Y=1.08 $X2=0
+ $Y2=0
cc_1437 N_A_1486_47#_c_1957_n N_A_c_2272_n 0.0156388f $X=9.6 $Y=1.295 $X2=0
+ $Y2=0
cc_1438 N_A_1486_47#_c_1953_n N_A_c_2273_n 0.00304573f $X=14.92 $Y=1.295 $X2=0
+ $Y2=0
cc_1439 N_A_1486_47#_c_1958_n N_A_c_2273_n 6.13516e-19 $X=10.57 $Y=1.295 $X2=0
+ $Y2=0
cc_1440 N_A_1486_47#_c_1959_n N_A_c_2273_n 0.0326668f $X=10.69 $Y=1.16 $X2=0
+ $Y2=0
cc_1441 N_A_1486_47#_M1068_g N_A_c_2274_n 0.0138261f $X=10.45 $Y=2.285 $X2=0
+ $Y2=0
cc_1442 N_A_1486_47#_c_1942_n N_A_c_2274_n 0.0077399f $X=10.615 $Y=1.69 $X2=0
+ $Y2=0
cc_1443 N_A_1486_47#_M1065_g N_A_c_2275_n 0.00325661f $X=10.67 $Y=0.445 $X2=0
+ $Y2=0
cc_1444 N_A_1486_47#_M1065_g A 6.20888e-19 $X=10.67 $Y=0.445 $X2=0 $Y2=0
cc_1445 N_A_1486_47#_c_1953_n A 0.00199402f $X=14.92 $Y=1.295 $X2=0 $Y2=0
cc_1446 N_A_1486_47#_c_1953_n N_A_2063_47#_c_2481_n 0.00665425f $X=14.92
+ $Y=1.295 $X2=0 $Y2=0
cc_1447 N_A_1486_47#_c_1955_n N_A_2063_47#_c_2482_n 2.65929e-19 $X=15.035
+ $Y=1.295 $X2=0 $Y2=0
cc_1448 N_A_1486_47#_c_1960_n N_A_2063_47#_c_2482_n 0.00926198f $X=15.625 $Y=1.2
+ $X2=0 $Y2=0
cc_1449 N_A_1486_47#_c_1961_n N_A_2063_47#_c_2482_n 8.65471e-19 $X=15.065 $Y=1.2
+ $X2=0 $Y2=0
cc_1450 N_A_1486_47#_M1065_g N_A_2063_47#_c_2483_n 0.011988f $X=10.67 $Y=0.445
+ $X2=0 $Y2=0
cc_1451 N_A_1486_47#_c_1953_n N_A_2063_47#_c_2483_n 0.0062871f $X=14.92 $Y=1.295
+ $X2=0 $Y2=0
cc_1452 N_A_1486_47#_c_1954_n N_A_2063_47#_c_2483_n 7.67525e-19 $X=10.715
+ $Y=1.295 $X2=0 $Y2=0
cc_1453 N_A_1486_47#_c_1958_n N_A_2063_47#_c_2483_n 0.0173982f $X=10.57 $Y=1.295
+ $X2=0 $Y2=0
cc_1454 N_A_1486_47#_c_1959_n N_A_2063_47#_c_2483_n 0.00484373f $X=10.69 $Y=1.16
+ $X2=0 $Y2=0
cc_1455 N_A_1486_47#_c_1951_n N_A_2063_47#_c_2484_n 0.00263275f $X=10.425
+ $Y=1.295 $X2=0 $Y2=0
cc_1456 N_A_1486_47#_c_1954_n N_A_2063_47#_c_2484_n 0.00302244f $X=10.715
+ $Y=1.295 $X2=0 $Y2=0
cc_1457 N_A_1486_47#_c_1958_n N_A_2063_47#_c_2484_n 0.00525667f $X=10.57
+ $Y=1.295 $X2=0 $Y2=0
cc_1458 N_A_1486_47#_c_1959_n N_A_2063_47#_c_2484_n 6.67758e-19 $X=10.69 $Y=1.16
+ $X2=0 $Y2=0
cc_1459 N_A_1486_47#_M1065_g N_A_2063_47#_c_2485_n 0.00275516f $X=10.67 $Y=0.445
+ $X2=0 $Y2=0
cc_1460 N_A_1486_47#_M1068_g N_A_2063_47#_c_2486_n 0.002305f $X=10.45 $Y=2.285
+ $X2=0 $Y2=0
cc_1461 N_A_1486_47#_c_1953_n N_A_2063_47#_c_2486_n 0.0190398f $X=14.92 $Y=1.295
+ $X2=0 $Y2=0
cc_1462 N_A_1486_47#_c_1954_n N_A_2063_47#_c_2486_n 5.43417e-19 $X=10.715
+ $Y=1.295 $X2=0 $Y2=0
cc_1463 N_A_1486_47#_c_1958_n N_A_2063_47#_c_2486_n 0.0380996f $X=10.57 $Y=1.295
+ $X2=0 $Y2=0
cc_1464 N_A_1486_47#_c_1959_n N_A_2063_47#_c_2486_n 0.00347397f $X=10.69 $Y=1.16
+ $X2=0 $Y2=0
cc_1465 N_A_1486_47#_c_1953_n N_A_2063_47#_c_2487_n 0.0413075f $X=14.92 $Y=1.295
+ $X2=0 $Y2=0
cc_1466 N_A_1486_47#_c_1953_n N_A_2063_47#_c_2488_n 0.00870395f $X=14.92
+ $Y=1.295 $X2=0 $Y2=0
cc_1467 N_A_1486_47#_c_1953_n N_A_2063_47#_c_2489_n 0.00680367f $X=14.92
+ $Y=1.295 $X2=0 $Y2=0
cc_1468 N_A_1486_47#_c_1953_n N_A_2063_47#_c_2490_n 0.0527918f $X=14.92 $Y=1.295
+ $X2=0 $Y2=0
cc_1469 N_A_1486_47#_M1068_g N_A_2063_47#_c_2495_n 0.0136494f $X=10.45 $Y=2.285
+ $X2=0 $Y2=0
cc_1470 N_A_1486_47#_M1068_g N_A_2063_47#_c_2496_n 0.00309056f $X=10.45 $Y=2.285
+ $X2=0 $Y2=0
cc_1471 N_A_1486_47#_c_1942_n N_A_2063_47#_c_2496_n 0.00714038f $X=10.615
+ $Y=1.69 $X2=0 $Y2=0
cc_1472 N_A_1486_47#_c_1958_n N_A_2063_47#_c_2496_n 0.0175369f $X=10.57 $Y=1.295
+ $X2=0 $Y2=0
cc_1473 N_A_1486_47#_M1065_g N_A_2063_47#_c_2491_n 0.00105159f $X=10.67 $Y=0.445
+ $X2=0 $Y2=0
cc_1474 N_A_1486_47#_c_1958_n N_A_2063_47#_c_2491_n 0.0113191f $X=10.57 $Y=1.295
+ $X2=0 $Y2=0
cc_1475 N_A_1486_47#_c_1959_n N_A_2063_47#_c_2491_n 9.70073e-19 $X=10.69 $Y=1.16
+ $X2=0 $Y2=0
cc_1476 N_A_1486_47#_c_1953_n N_A_2063_47#_c_2492_n 0.00929668f $X=14.92
+ $Y=1.295 $X2=0 $Y2=0
cc_1477 N_A_1486_47#_M1068_g N_VPWR_c_2632_n 0.00344549f $X=10.45 $Y=2.285 $X2=0
+ $Y2=0
cc_1478 N_A_1486_47#_c_1957_n N_VPWR_c_2632_n 0.00101432f $X=9.6 $Y=1.295 $X2=0
+ $Y2=0
cc_1479 N_A_1486_47#_M1023_d N_VPWR_c_2627_n 0.00114355f $X=7.875 $Y=1.835 $X2=0
+ $Y2=0
cc_1480 N_A_1486_47#_M1023_d KAPWR 0.0012473f $X=7.875 $Y=1.835 $X2=0 $Y2=0
cc_1481 N_A_1486_47#_M1068_g KAPWR 0.00440817f $X=10.45 $Y=2.285 $X2=0 $Y2=0
cc_1482 N_A_1486_47#_c_1948_n KAPWR 0.00906391f $X=8.015 $Y=1.98 $X2=0 $Y2=0
cc_1483 N_A_1486_47#_c_1948_n N_A_1492_367#_c_3237_n 0.0360913f $X=8.015 $Y=1.98
+ $X2=0 $Y2=0
cc_1484 N_A_1486_47#_M1023_d N_A_1492_367#_c_3255_n 0.00242215f $X=7.875
+ $Y=1.835 $X2=0 $Y2=0
cc_1485 N_A_1486_47#_c_1948_n N_A_1492_367#_c_3255_n 0.0117275f $X=8.015 $Y=1.98
+ $X2=0 $Y2=0
cc_1486 N_A_1486_47#_c_1948_n N_A_1492_367#_c_3238_n 0.0218145f $X=8.015 $Y=1.98
+ $X2=0 $Y2=0
cc_1487 N_A_1486_47#_c_1949_n N_A_1492_367#_c_3238_n 0.00419213f $X=9.455
+ $Y=1.08 $X2=0 $Y2=0
cc_1488 N_A_1486_47#_c_1948_n N_A_1492_367#_c_3258_n 0.00854184f $X=8.015
+ $Y=1.98 $X2=0 $Y2=0
cc_1489 N_A_1486_47#_c_1960_n N_Z_c_3379_n 0.00147174f $X=15.625 $Y=1.2 $X2=0
+ $Y2=0
cc_1490 N_A_1486_47#_c_1961_n N_Z_c_3379_n 0.00349691f $X=15.065 $Y=1.2 $X2=0
+ $Y2=0
cc_1491 N_A_1486_47#_M1000_g N_Z_c_3367_n 0.0126545f $X=15.7 $Y=0.555 $X2=0
+ $Y2=0
cc_1492 N_A_1486_47#_M1009_g N_Z_c_3367_n 6.57936e-19 $X=16.13 $Y=0.555 $X2=0
+ $Y2=0
cc_1493 N_A_1486_47#_c_1929_n N_Z_c_3367_n 0.00440309f $X=18.785 $Y=1.06 $X2=0
+ $Y2=0
cc_1494 N_A_1486_47#_c_1956_n N_Z_c_3367_n 0.0353753f $X=18.505 $Y=1.295 $X2=0
+ $Y2=0
cc_1495 N_A_1486_47#_c_1960_n N_Z_c_3367_n 0.0230572f $X=15.625 $Y=1.2 $X2=0
+ $Y2=0
cc_1496 N_A_1486_47#_c_1961_n N_Z_c_3367_n 0.0256972f $X=15.065 $Y=1.2 $X2=0
+ $Y2=0
cc_1497 N_A_1486_47#_c_1962_n N_Z_c_3367_n 0.0256972f $X=15.925 $Y=1.2 $X2=0
+ $Y2=0
cc_1498 N_A_1486_47#_M1000_g N_Z_c_3368_n 6.57936e-19 $X=15.7 $Y=0.555 $X2=0
+ $Y2=0
cc_1499 N_A_1486_47#_M1009_g N_Z_c_3368_n 0.0113519f $X=16.13 $Y=0.555 $X2=0
+ $Y2=0
cc_1500 N_A_1486_47#_M1021_g N_Z_c_3368_n 0.0113519f $X=16.56 $Y=0.555 $X2=0
+ $Y2=0
cc_1501 N_A_1486_47#_M1025_g N_Z_c_3368_n 6.57936e-19 $X=16.99 $Y=0.555 $X2=0
+ $Y2=0
cc_1502 N_A_1486_47#_c_1929_n N_Z_c_3368_n 0.022527f $X=18.785 $Y=1.06 $X2=0
+ $Y2=0
cc_1503 N_A_1486_47#_c_1956_n N_Z_c_3368_n 0.0353753f $X=18.505 $Y=1.295 $X2=0
+ $Y2=0
cc_1504 N_A_1486_47#_c_1962_n N_Z_c_3368_n 0.0256972f $X=15.925 $Y=1.2 $X2=0
+ $Y2=0
cc_1505 N_A_1486_47#_c_1963_n N_Z_c_3368_n 0.0256972f $X=16.765 $Y=1.2 $X2=0
+ $Y2=0
cc_1506 N_A_1486_47#_M1021_g N_Z_c_3369_n 6.57936e-19 $X=16.56 $Y=0.555 $X2=0
+ $Y2=0
cc_1507 N_A_1486_47#_M1025_g N_Z_c_3369_n 0.0113519f $X=16.99 $Y=0.555 $X2=0
+ $Y2=0
cc_1508 N_A_1486_47#_c_1924_n N_Z_c_3369_n 0.00987762f $X=17.42 $Y=0.985 $X2=0
+ $Y2=0
cc_1509 N_A_1486_47#_c_1925_n N_Z_c_3369_n 5.10745e-19 $X=17.85 $Y=0.985 $X2=0
+ $Y2=0
cc_1510 N_A_1486_47#_c_1929_n N_Z_c_3369_n 0.024478f $X=18.785 $Y=1.06 $X2=0
+ $Y2=0
cc_1511 N_A_1486_47#_c_1956_n N_Z_c_3369_n 0.0353753f $X=18.505 $Y=1.295 $X2=0
+ $Y2=0
cc_1512 N_A_1486_47#_c_1963_n N_Z_c_3369_n 0.0256972f $X=16.765 $Y=1.2 $X2=0
+ $Y2=0
cc_1513 N_A_1486_47#_c_1964_n N_Z_c_3369_n 0.0256972f $X=17.645 $Y=1.2 $X2=0
+ $Y2=0
cc_1514 N_A_1486_47#_c_1924_n N_Z_c_3370_n 5.10745e-19 $X=17.42 $Y=0.985 $X2=0
+ $Y2=0
cc_1515 N_A_1486_47#_c_1925_n N_Z_c_3370_n 0.00987762f $X=17.85 $Y=0.985 $X2=0
+ $Y2=0
cc_1516 N_A_1486_47#_c_1926_n N_Z_c_3370_n 0.00987762f $X=18.28 $Y=0.985 $X2=0
+ $Y2=0
cc_1517 N_A_1486_47#_c_1927_n N_Z_c_3370_n 5.10745e-19 $X=18.71 $Y=0.985 $X2=0
+ $Y2=0
cc_1518 N_A_1486_47#_c_1929_n N_Z_c_3370_n 0.0265644f $X=18.785 $Y=1.06 $X2=0
+ $Y2=0
cc_1519 N_A_1486_47#_c_1956_n N_Z_c_3370_n 0.0353753f $X=18.505 $Y=1.295 $X2=0
+ $Y2=0
cc_1520 N_A_1486_47#_c_1964_n N_Z_c_3370_n 0.0256972f $X=17.645 $Y=1.2 $X2=0
+ $Y2=0
cc_1521 N_A_1486_47#_c_1965_n N_Z_c_3370_n 0.0256972f $X=18.505 $Y=1.2 $X2=0
+ $Y2=0
cc_1522 N_A_1486_47#_c_1926_n N_Z_c_3371_n 5.10745e-19 $X=18.28 $Y=0.985 $X2=0
+ $Y2=0
cc_1523 N_A_1486_47#_c_1927_n N_Z_c_3371_n 0.00987762f $X=18.71 $Y=0.985 $X2=0
+ $Y2=0
cc_1524 N_A_1486_47#_c_1928_n N_Z_c_3371_n 0.0109356f $X=19.065 $Y=1.06 $X2=0
+ $Y2=0
cc_1525 N_A_1486_47#_c_1929_n N_Z_c_3371_n 0.00850001f $X=18.785 $Y=1.06 $X2=0
+ $Y2=0
cc_1526 N_A_1486_47#_c_1930_n N_Z_c_3371_n 0.00987762f $X=19.14 $Y=0.985 $X2=0
+ $Y2=0
cc_1527 N_A_1486_47#_c_1932_n N_Z_c_3371_n 5.10745e-19 $X=19.57 $Y=0.985 $X2=0
+ $Y2=0
cc_1528 N_A_1486_47#_c_1943_n N_Z_c_3371_n 0.00446221f $X=19.14 $Y=1.06 $X2=0
+ $Y2=0
cc_1529 N_A_1486_47#_c_1956_n N_Z_c_3371_n 0.00871004f $X=18.505 $Y=1.295 $X2=0
+ $Y2=0
cc_1530 N_A_1486_47#_c_1965_n N_Z_c_3371_n 0.0256915f $X=18.505 $Y=1.2 $X2=0
+ $Y2=0
cc_1531 N_A_1486_47#_c_1930_n N_Z_c_3372_n 5.10745e-19 $X=19.14 $Y=0.985 $X2=0
+ $Y2=0
cc_1532 N_A_1486_47#_c_1932_n N_Z_c_3372_n 0.00987762f $X=19.57 $Y=0.985 $X2=0
+ $Y2=0
cc_1533 N_A_1486_47#_c_1933_n N_Z_c_3372_n 0.0088652f $X=19.925 $Y=1.06 $X2=0
+ $Y2=0
cc_1534 N_A_1486_47#_c_1934_n N_Z_c_3372_n 0.00987762f $X=20 $Y=0.985 $X2=0
+ $Y2=0
cc_1535 N_A_1486_47#_c_1936_n N_Z_c_3372_n 5.10745e-19 $X=20.43 $Y=0.985 $X2=0
+ $Y2=0
cc_1536 N_A_1486_47#_c_1944_n N_Z_c_3372_n 0.00428178f $X=19.57 $Y=1.06 $X2=0
+ $Y2=0
cc_1537 N_A_1486_47#_c_1945_n N_Z_c_3372_n 0.00428178f $X=20 $Y=1.06 $X2=0 $Y2=0
cc_1538 N_A_1486_47#_c_1934_n N_Z_c_3373_n 5.09252e-19 $X=20 $Y=0.985 $X2=0
+ $Y2=0
cc_1539 N_A_1486_47#_c_1936_n N_Z_c_3373_n 0.00983119f $X=20.43 $Y=0.985 $X2=0
+ $Y2=0
cc_1540 N_A_1486_47#_c_1937_n N_Z_c_3373_n 0.0088652f $X=20.785 $Y=1.06 $X2=0
+ $Y2=0
cc_1541 N_A_1486_47#_c_1938_n N_Z_c_3373_n 0.00983119f $X=20.86 $Y=0.985 $X2=0
+ $Y2=0
cc_1542 N_A_1486_47#_c_1940_n N_Z_c_3373_n 5.09252e-19 $X=21.29 $Y=0.985 $X2=0
+ $Y2=0
cc_1543 N_A_1486_47#_c_1946_n N_Z_c_3373_n 0.00428178f $X=20.43 $Y=1.06 $X2=0
+ $Y2=0
cc_1544 N_A_1486_47#_c_1947_n N_Z_c_3373_n 0.00428178f $X=20.86 $Y=1.06 $X2=0
+ $Y2=0
cc_1545 N_A_1486_47#_c_1938_n N_Z_c_3374_n 5.10745e-19 $X=20.86 $Y=0.985 $X2=0
+ $Y2=0
cc_1546 N_A_1486_47#_c_1939_n N_Z_c_3374_n 0.00731f $X=21.215 $Y=1.06 $X2=0
+ $Y2=0
cc_1547 N_A_1486_47#_c_1940_n N_Z_c_3374_n 0.010768f $X=21.29 $Y=0.985 $X2=0
+ $Y2=0
cc_1548 N_A_1486_47#_c_1949_n N_VGND_M1050_s 0.00637658f $X=9.455 $Y=1.08 $X2=0
+ $Y2=0
cc_1549 N_A_1486_47#_c_1949_n N_VGND_M1071_s 0.00243229f $X=9.455 $Y=1.08 $X2=0
+ $Y2=0
cc_1550 N_A_1486_47#_M1065_g N_VGND_c_3669_n 0.00354752f $X=10.67 $Y=0.445 $X2=0
+ $Y2=0
cc_1551 N_A_1486_47#_M1065_g N_VGND_c_3670_n 0.00757954f $X=10.67 $Y=0.445 $X2=0
+ $Y2=0
cc_1552 N_A_1486_47#_M1000_g N_VGND_c_3672_n 0.00271808f $X=15.7 $Y=0.555 $X2=0
+ $Y2=0
cc_1553 N_A_1486_47#_M1009_g N_VGND_c_3672_n 0.00271808f $X=16.13 $Y=0.555 $X2=0
+ $Y2=0
cc_1554 N_A_1486_47#_c_1929_n N_VGND_c_3672_n 7.91474e-19 $X=18.785 $Y=1.06
+ $X2=0 $Y2=0
cc_1555 N_A_1486_47#_c_1956_n N_VGND_c_3672_n 0.00100776f $X=18.505 $Y=1.295
+ $X2=0 $Y2=0
cc_1556 N_A_1486_47#_c_1962_n N_VGND_c_3672_n 0.0130159f $X=15.925 $Y=1.2 $X2=0
+ $Y2=0
cc_1557 N_A_1486_47#_M1021_g N_VGND_c_3673_n 0.00271808f $X=16.56 $Y=0.555 $X2=0
+ $Y2=0
cc_1558 N_A_1486_47#_M1025_g N_VGND_c_3673_n 0.00271808f $X=16.99 $Y=0.555 $X2=0
+ $Y2=0
cc_1559 N_A_1486_47#_c_1929_n N_VGND_c_3673_n 7.91474e-19 $X=18.785 $Y=1.06
+ $X2=0 $Y2=0
cc_1560 N_A_1486_47#_c_1956_n N_VGND_c_3673_n 0.00100776f $X=18.505 $Y=1.295
+ $X2=0 $Y2=0
cc_1561 N_A_1486_47#_c_1963_n N_VGND_c_3673_n 0.0130159f $X=16.765 $Y=1.2 $X2=0
+ $Y2=0
cc_1562 N_A_1486_47#_c_1924_n N_VGND_c_3674_n 0.00271808f $X=17.42 $Y=0.985
+ $X2=0 $Y2=0
cc_1563 N_A_1486_47#_c_1925_n N_VGND_c_3674_n 0.00271808f $X=17.85 $Y=0.985
+ $X2=0 $Y2=0
cc_1564 N_A_1486_47#_c_1929_n N_VGND_c_3674_n 0.00254294f $X=18.785 $Y=1.06
+ $X2=0 $Y2=0
cc_1565 N_A_1486_47#_c_1956_n N_VGND_c_3674_n 0.00100776f $X=18.505 $Y=1.295
+ $X2=0 $Y2=0
cc_1566 N_A_1486_47#_c_1964_n N_VGND_c_3674_n 0.0130158f $X=17.645 $Y=1.2 $X2=0
+ $Y2=0
cc_1567 N_A_1486_47#_c_1925_n N_VGND_c_3675_n 0.0054895f $X=17.85 $Y=0.985 $X2=0
+ $Y2=0
cc_1568 N_A_1486_47#_c_1926_n N_VGND_c_3675_n 0.0054895f $X=18.28 $Y=0.985 $X2=0
+ $Y2=0
cc_1569 N_A_1486_47#_c_1926_n N_VGND_c_3676_n 0.00271808f $X=18.28 $Y=0.985
+ $X2=0 $Y2=0
cc_1570 N_A_1486_47#_c_1927_n N_VGND_c_3676_n 0.00271808f $X=18.71 $Y=0.985
+ $X2=0 $Y2=0
cc_1571 N_A_1486_47#_c_1929_n N_VGND_c_3676_n 0.00254294f $X=18.785 $Y=1.06
+ $X2=0 $Y2=0
cc_1572 N_A_1486_47#_c_1956_n N_VGND_c_3676_n 0.00100776f $X=18.505 $Y=1.295
+ $X2=0 $Y2=0
cc_1573 N_A_1486_47#_c_1965_n N_VGND_c_3676_n 0.0130158f $X=18.505 $Y=1.2 $X2=0
+ $Y2=0
cc_1574 N_A_1486_47#_c_1930_n N_VGND_c_3677_n 0.00271808f $X=19.14 $Y=0.985
+ $X2=0 $Y2=0
cc_1575 N_A_1486_47#_c_1931_n N_VGND_c_3677_n 0.0026233f $X=19.495 $Y=1.06 $X2=0
+ $Y2=0
cc_1576 N_A_1486_47#_c_1932_n N_VGND_c_3677_n 0.00271808f $X=19.57 $Y=0.985
+ $X2=0 $Y2=0
cc_1577 N_A_1486_47#_c_1934_n N_VGND_c_3678_n 0.00271808f $X=20 $Y=0.985 $X2=0
+ $Y2=0
cc_1578 N_A_1486_47#_c_1935_n N_VGND_c_3678_n 0.0026233f $X=20.355 $Y=1.06 $X2=0
+ $Y2=0
cc_1579 N_A_1486_47#_c_1936_n N_VGND_c_3678_n 0.00271808f $X=20.43 $Y=0.985
+ $X2=0 $Y2=0
cc_1580 N_A_1486_47#_c_1938_n N_VGND_c_3679_n 0.00271808f $X=20.86 $Y=0.985
+ $X2=0 $Y2=0
cc_1581 N_A_1486_47#_c_1939_n N_VGND_c_3679_n 0.0026233f $X=21.215 $Y=1.06 $X2=0
+ $Y2=0
cc_1582 N_A_1486_47#_c_1940_n N_VGND_c_3679_n 0.00271808f $X=21.29 $Y=0.985
+ $X2=0 $Y2=0
cc_1583 N_A_1486_47#_M1000_g N_VGND_c_3692_n 0.0054895f $X=15.7 $Y=0.555 $X2=0
+ $Y2=0
cc_1584 N_A_1486_47#_M1009_g N_VGND_c_3694_n 0.0054895f $X=16.13 $Y=0.555 $X2=0
+ $Y2=0
cc_1585 N_A_1486_47#_M1021_g N_VGND_c_3694_n 0.0054895f $X=16.56 $Y=0.555 $X2=0
+ $Y2=0
cc_1586 N_A_1486_47#_M1025_g N_VGND_c_3696_n 0.0054895f $X=16.99 $Y=0.555 $X2=0
+ $Y2=0
cc_1587 N_A_1486_47#_c_1924_n N_VGND_c_3696_n 0.0054895f $X=17.42 $Y=0.985 $X2=0
+ $Y2=0
cc_1588 N_A_1486_47#_c_1927_n N_VGND_c_3698_n 0.0054895f $X=18.71 $Y=0.985 $X2=0
+ $Y2=0
cc_1589 N_A_1486_47#_c_1930_n N_VGND_c_3698_n 0.0054895f $X=19.14 $Y=0.985 $X2=0
+ $Y2=0
cc_1590 N_A_1486_47#_c_1932_n N_VGND_c_3700_n 0.0054895f $X=19.57 $Y=0.985 $X2=0
+ $Y2=0
cc_1591 N_A_1486_47#_c_1934_n N_VGND_c_3700_n 0.0054895f $X=20 $Y=0.985 $X2=0
+ $Y2=0
cc_1592 N_A_1486_47#_c_1936_n N_VGND_c_3702_n 0.00549117f $X=20.43 $Y=0.985
+ $X2=0 $Y2=0
cc_1593 N_A_1486_47#_c_1938_n N_VGND_c_3702_n 0.00549117f $X=20.86 $Y=0.985
+ $X2=0 $Y2=0
cc_1594 N_A_1486_47#_c_1940_n N_VGND_c_3706_n 0.0054895f $X=21.29 $Y=0.985 $X2=0
+ $Y2=0
cc_1595 N_A_1486_47#_M1038_d N_VGND_c_3707_n 0.00432472f $X=7.43 $Y=0.235 $X2=0
+ $Y2=0
cc_1596 N_A_1486_47#_M1003_d N_VGND_c_3707_n 0.00557193f $X=8.87 $Y=0.235 $X2=0
+ $Y2=0
cc_1597 N_A_1486_47#_M1065_g N_VGND_c_3707_n 0.00423947f $X=10.67 $Y=0.445 $X2=0
+ $Y2=0
cc_1598 N_A_1486_47#_M1000_g N_VGND_c_3707_n 0.0110927f $X=15.7 $Y=0.555 $X2=0
+ $Y2=0
cc_1599 N_A_1486_47#_M1009_g N_VGND_c_3707_n 0.00979301f $X=16.13 $Y=0.555 $X2=0
+ $Y2=0
cc_1600 N_A_1486_47#_M1021_g N_VGND_c_3707_n 0.00979301f $X=16.56 $Y=0.555 $X2=0
+ $Y2=0
cc_1601 N_A_1486_47#_M1025_g N_VGND_c_3707_n 0.00979301f $X=16.99 $Y=0.555 $X2=0
+ $Y2=0
cc_1602 N_A_1486_47#_c_1924_n N_VGND_c_3707_n 0.00979301f $X=17.42 $Y=0.985
+ $X2=0 $Y2=0
cc_1603 N_A_1486_47#_c_1925_n N_VGND_c_3707_n 0.00979301f $X=17.85 $Y=0.985
+ $X2=0 $Y2=0
cc_1604 N_A_1486_47#_c_1926_n N_VGND_c_3707_n 0.00979301f $X=18.28 $Y=0.985
+ $X2=0 $Y2=0
cc_1605 N_A_1486_47#_c_1927_n N_VGND_c_3707_n 0.00979301f $X=18.71 $Y=0.985
+ $X2=0 $Y2=0
cc_1606 N_A_1486_47#_c_1930_n N_VGND_c_3707_n 0.00979301f $X=19.14 $Y=0.985
+ $X2=0 $Y2=0
cc_1607 N_A_1486_47#_c_1932_n N_VGND_c_3707_n 0.00979301f $X=19.57 $Y=0.985
+ $X2=0 $Y2=0
cc_1608 N_A_1486_47#_c_1934_n N_VGND_c_3707_n 0.00979301f $X=20 $Y=0.985 $X2=0
+ $Y2=0
cc_1609 N_A_1486_47#_c_1936_n N_VGND_c_3707_n 0.00979311f $X=20.43 $Y=0.985
+ $X2=0 $Y2=0
cc_1610 N_A_1486_47#_c_1938_n N_VGND_c_3707_n 0.00979311f $X=20.86 $Y=0.985
+ $X2=0 $Y2=0
cc_1611 N_A_1486_47#_c_1940_n N_VGND_c_3707_n 0.0110927f $X=21.29 $Y=0.985 $X2=0
+ $Y2=0
cc_1612 N_A_1486_47#_M1065_g N_VGND_c_3710_n 5.95653e-19 $X=10.67 $Y=0.445 $X2=0
+ $Y2=0
cc_1613 N_A_1486_47#_c_1953_n N_A_2519_47#_c_3956_n 0.0256561f $X=14.92 $Y=1.295
+ $X2=0 $Y2=0
cc_1614 N_A_1486_47#_c_1953_n N_A_2519_47#_c_3957_n 0.00553971f $X=14.92
+ $Y=1.295 $X2=0 $Y2=0
cc_1615 N_A_1486_47#_c_1953_n N_A_2519_47#_c_3959_n 0.00821049f $X=14.92
+ $Y=1.295 $X2=0 $Y2=0
cc_1616 N_A_1486_47#_c_1960_n N_A_2519_47#_c_3959_n 6.57308e-19 $X=15.625 $Y=1.2
+ $X2=0 $Y2=0
cc_1617 N_A_1486_47#_c_1961_n N_A_2519_47#_c_3959_n 0.0044621f $X=15.065 $Y=1.2
+ $X2=0 $Y2=0
cc_1618 N_A_c_2265_n N_A_2063_47#_c_2483_n 0.00307498f $X=11.235 $Y=0.86 $X2=0
+ $Y2=0
cc_1619 N_A_c_2275_n N_A_2063_47#_c_2483_n 0.00112333f $X=11.647 $Y=0.687 $X2=0
+ $Y2=0
cc_1620 A N_A_2063_47#_c_2483_n 0.00803147f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1621 N_A_c_2265_n N_A_2063_47#_c_2485_n 0.00679754f $X=11.235 $Y=0.86 $X2=0
+ $Y2=0
cc_1622 N_A_c_2273_n N_A_2063_47#_c_2485_n 9.11108e-19 $X=11.15 $Y=1.575 $X2=0
+ $Y2=0
cc_1623 N_A_c_2286_n N_A_2063_47#_c_2486_n 0.00406364f $X=11.14 $Y=3.075 $X2=0
+ $Y2=0
cc_1624 N_A_c_2273_n N_A_2063_47#_c_2486_n 0.0123378f $X=11.15 $Y=1.575 $X2=0
+ $Y2=0
cc_1625 N_A_c_2274_n N_A_2063_47#_c_2486_n 0.003897f $X=11.15 $Y=1.725 $X2=0
+ $Y2=0
cc_1626 N_A_c_2266_n N_A_2063_47#_c_2487_n 0.0110461f $X=12.44 $Y=1.575 $X2=0
+ $Y2=0
cc_1627 N_A_M1007_g N_A_2063_47#_c_2487_n 3.11937e-19 $X=12.935 $Y=0.655 $X2=0
+ $Y2=0
cc_1628 N_A_c_2273_n N_A_2063_47#_c_2487_n 0.010719f $X=11.15 $Y=1.575 $X2=0
+ $Y2=0
cc_1629 N_A_c_2276_n N_A_2063_47#_c_2487_n 0.0152262f $X=11.4 $Y=0.687 $X2=0
+ $Y2=0
cc_1630 A N_A_2063_47#_c_2487_n 0.0667321f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1631 N_A_c_2266_n N_A_2063_47#_c_2488_n 0.00570167f $X=12.44 $Y=1.575 $X2=0
+ $Y2=0
cc_1632 N_A_M1007_g N_A_2063_47#_c_2488_n 8.84125e-19 $X=12.935 $Y=0.655 $X2=0
+ $Y2=0
cc_1633 N_A_c_2266_n N_A_2063_47#_c_2489_n 0.00371922f $X=12.44 $Y=1.575 $X2=0
+ $Y2=0
cc_1634 N_A_c_2268_n N_A_2063_47#_c_2489_n 0.00209488f $X=12.515 $Y=1.65 $X2=0
+ $Y2=0
cc_1635 N_A_c_2266_n N_A_2063_47#_c_2490_n 0.00727954f $X=12.44 $Y=1.575 $X2=0
+ $Y2=0
cc_1636 N_A_c_2267_n N_A_2063_47#_c_2490_n 0.00922189f $X=12.86 $Y=1.65 $X2=0
+ $Y2=0
cc_1637 N_A_c_2268_n N_A_2063_47#_c_2490_n 0.0012938f $X=12.515 $Y=1.65 $X2=0
+ $Y2=0
cc_1638 N_A_M1007_g N_A_2063_47#_c_2490_n 0.0139339f $X=12.935 $Y=0.655 $X2=0
+ $Y2=0
cc_1639 N_A_c_2270_n N_A_2063_47#_c_2490_n 0.00714878f $X=13.385 $Y=1.65 $X2=0
+ $Y2=0
cc_1640 N_A_M1041_g N_A_2063_47#_c_2490_n 0.0125543f $X=13.46 $Y=0.655 $X2=0
+ $Y2=0
cc_1641 N_A_c_2278_n N_A_2063_47#_c_2490_n 0.00532433f $X=12.982 $Y=1.65 $X2=0
+ $Y2=0
cc_1642 N_A_c_2279_n N_A_2063_47#_c_2490_n 0.00187458f $X=13.46 $Y=1.65 $X2=0
+ $Y2=0
cc_1643 N_A_c_2284_n N_A_2063_47#_c_2495_n 0.00541204f $X=11.065 $Y=3.15 $X2=0
+ $Y2=0
cc_1644 N_A_c_2286_n N_A_2063_47#_c_2495_n 0.0106945f $X=11.14 $Y=3.075 $X2=0
+ $Y2=0
cc_1645 N_A_c_2286_n N_A_2063_47#_c_2496_n 0.00846917f $X=11.14 $Y=3.075 $X2=0
+ $Y2=0
cc_1646 N_A_c_2273_n N_A_2063_47#_c_2491_n 0.00192837f $X=11.15 $Y=1.575 $X2=0
+ $Y2=0
cc_1647 N_A_M1041_g N_A_2063_47#_c_2492_n 0.0277978f $X=13.46 $Y=0.655 $X2=0
+ $Y2=0
cc_1648 N_A_M1041_g N_A_2063_47#_c_2493_n 0.0228319f $X=13.46 $Y=0.655 $X2=0
+ $Y2=0
cc_1649 N_A_c_2281_n N_VPWR_c_2631_n 0.00351376f $X=8.66 $Y=1.715 $X2=0 $Y2=0
cc_1650 N_A_c_2282_n N_VPWR_c_2631_n 0.00822433f $X=9.09 $Y=1.715 $X2=0 $Y2=0
cc_1651 N_A_c_2283_n N_VPWR_c_2631_n 7.62468e-19 $X=9.58 $Y=3.075 $X2=0 $Y2=0
cc_1652 N_A_c_2282_n N_VPWR_c_2632_n 4.19165e-19 $X=9.09 $Y=1.715 $X2=0 $Y2=0
cc_1653 N_A_c_2283_n N_VPWR_c_2632_n 0.0224336f $X=9.58 $Y=3.075 $X2=0 $Y2=0
cc_1654 N_A_c_2284_n N_VPWR_c_2632_n 0.0233904f $X=11.065 $Y=3.15 $X2=0 $Y2=0
cc_1655 N_A_c_2286_n N_VPWR_c_2633_n 0.016741f $X=11.14 $Y=3.075 $X2=0 $Y2=0
cc_1656 N_A_c_2289_n N_VPWR_c_2635_n 0.00225841f $X=13.03 $Y=1.725 $X2=0 $Y2=0
cc_1657 N_A_c_2291_n N_VPWR_c_2636_n 0.00363222f $X=13.46 $Y=1.725 $X2=0 $Y2=0
cc_1658 N_A_c_2281_n N_VPWR_c_2668_n 0.0054778f $X=8.66 $Y=1.715 $X2=0 $Y2=0
cc_1659 N_A_c_2282_n N_VPWR_c_2669_n 0.00486043f $X=9.09 $Y=1.715 $X2=0 $Y2=0
cc_1660 N_A_c_2285_n N_VPWR_c_2669_n 0.00796123f $X=9.655 $Y=3.15 $X2=0 $Y2=0
cc_1661 N_A_c_2284_n N_VPWR_c_2670_n 0.0387249f $X=11.065 $Y=3.15 $X2=0 $Y2=0
cc_1662 N_A_c_2289_n N_VPWR_c_2671_n 0.00357842f $X=13.03 $Y=1.725 $X2=0 $Y2=0
cc_1663 N_A_c_2291_n N_VPWR_c_2671_n 0.00357877f $X=13.46 $Y=1.725 $X2=0 $Y2=0
cc_1664 N_A_c_2281_n N_VPWR_c_2627_n 0.00490302f $X=8.66 $Y=1.715 $X2=0 $Y2=0
cc_1665 N_A_c_2282_n N_VPWR_c_2627_n 0.00361338f $X=9.09 $Y=1.715 $X2=0 $Y2=0
cc_1666 N_A_c_2284_n N_VPWR_c_2627_n 0.025376f $X=11.065 $Y=3.15 $X2=0 $Y2=0
cc_1667 N_A_c_2285_n N_VPWR_c_2627_n 0.00457585f $X=9.655 $Y=3.15 $X2=0 $Y2=0
cc_1668 N_A_c_2289_n N_VPWR_c_2627_n 0.00605388f $X=13.03 $Y=1.725 $X2=0 $Y2=0
cc_1669 N_A_c_2291_n N_VPWR_c_2627_n 0.00605389f $X=13.46 $Y=1.725 $X2=0 $Y2=0
cc_1670 N_A_c_2281_n KAPWR 0.00191104f $X=8.66 $Y=1.715 $X2=0 $Y2=0
cc_1671 N_A_c_2282_n KAPWR 0.00192048f $X=9.09 $Y=1.715 $X2=0 $Y2=0
cc_1672 N_A_c_2283_n KAPWR 0.00891568f $X=9.58 $Y=3.075 $X2=0 $Y2=0
cc_1673 N_A_c_2284_n KAPWR 0.00910781f $X=11.065 $Y=3.15 $X2=0 $Y2=0
cc_1674 N_A_c_2286_n KAPWR 0.0102074f $X=11.14 $Y=3.075 $X2=0 $Y2=0
cc_1675 N_A_c_2289_n KAPWR 0.00610801f $X=13.03 $Y=1.725 $X2=0 $Y2=0
cc_1676 N_A_c_2291_n KAPWR 0.00696289f $X=13.46 $Y=1.725 $X2=0 $Y2=0
cc_1677 N_A_c_2281_n N_A_1492_367#_c_3238_n 0.0113008f $X=8.66 $Y=1.715 $X2=0
+ $Y2=0
cc_1678 N_A_c_2282_n N_A_1492_367#_c_3238_n 0.00294186f $X=9.09 $Y=1.715 $X2=0
+ $Y2=0
cc_1679 N_A_c_2281_n N_A_1492_367#_c_3258_n 0.00729651f $X=8.66 $Y=1.715 $X2=0
+ $Y2=0
cc_1680 N_A_c_2282_n N_A_1492_367#_c_3258_n 5.33199e-19 $X=9.09 $Y=1.715 $X2=0
+ $Y2=0
cc_1681 N_A_c_2281_n N_A_1492_367#_c_3244_n 0.00817057f $X=8.66 $Y=1.715 $X2=0
+ $Y2=0
cc_1682 N_A_c_2282_n N_A_1492_367#_c_3244_n 0.00932616f $X=9.09 $Y=1.715 $X2=0
+ $Y2=0
cc_1683 N_A_c_2272_n N_A_1492_367#_c_3244_n 0.00187703f $X=9.405 $Y=1.562 $X2=0
+ $Y2=0
cc_1684 N_A_c_2281_n N_A_1492_367#_c_3260_n 4.0679e-19 $X=8.66 $Y=1.715 $X2=0
+ $Y2=0
cc_1685 N_A_c_2282_n N_A_1492_367#_c_3239_n 5.74483e-19 $X=9.09 $Y=1.715 $X2=0
+ $Y2=0
cc_1686 N_A_c_2283_n N_A_1492_367#_c_3239_n 0.00693331f $X=9.58 $Y=3.075 $X2=0
+ $Y2=0
cc_1687 N_A_c_2272_n N_A_1492_367#_c_3239_n 0.00367995f $X=9.405 $Y=1.562 $X2=0
+ $Y2=0
cc_1688 N_A_c_2268_n N_A_2345_367#_c_3306_n 0.00529777f $X=12.515 $Y=1.65 $X2=0
+ $Y2=0
cc_1689 N_A_c_2267_n N_A_2345_367#_c_3307_n 0.00409996f $X=12.86 $Y=1.65 $X2=0
+ $Y2=0
cc_1690 N_A_c_2289_n N_A_2345_367#_c_3307_n 0.00375656f $X=13.03 $Y=1.725 $X2=0
+ $Y2=0
cc_1691 N_A_c_2289_n N_A_2345_367#_c_3308_n 0.00731319f $X=13.03 $Y=1.725 $X2=0
+ $Y2=0
cc_1692 N_A_c_2291_n N_A_2345_367#_c_3308_n 4.94364e-19 $X=13.46 $Y=1.725 $X2=0
+ $Y2=0
cc_1693 N_A_c_2289_n N_A_2345_367#_c_3327_n 0.0110776f $X=13.03 $Y=1.725 $X2=0
+ $Y2=0
cc_1694 N_A_c_2291_n N_A_2345_367#_c_3327_n 0.0121982f $X=13.46 $Y=1.725 $X2=0
+ $Y2=0
cc_1695 N_A_c_2289_n N_A_2345_367#_c_3309_n 8.83566e-19 $X=13.03 $Y=1.725 $X2=0
+ $Y2=0
cc_1696 N_A_c_2291_n N_A_2345_367#_c_3311_n 0.00351247f $X=13.46 $Y=1.725 $X2=0
+ $Y2=0
cc_1697 N_A_M1003_g N_VGND_c_3668_n 0.0118244f $X=8.795 $Y=0.655 $X2=0 $Y2=0
cc_1698 N_A_M1071_g N_VGND_c_3668_n 0.00118042f $X=9.405 $Y=0.655 $X2=0 $Y2=0
cc_1699 A N_VGND_c_3670_n 0.00117226f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1700 N_A_M1007_g N_VGND_c_3671_n 0.00396327f $X=12.935 $Y=0.655 $X2=0 $Y2=0
cc_1701 N_A_M1041_g N_VGND_c_3671_n 0.00416483f $X=13.46 $Y=0.655 $X2=0 $Y2=0
cc_1702 N_A_M1041_g N_VGND_c_3692_n 0.00585385f $X=13.46 $Y=0.655 $X2=0 $Y2=0
cc_1703 N_A_M1007_g N_VGND_c_3705_n 0.00548839f $X=12.935 $Y=0.655 $X2=0 $Y2=0
cc_1704 N_A_c_2275_n N_VGND_c_3705_n 0.0240071f $X=11.647 $Y=0.687 $X2=0 $Y2=0
cc_1705 A N_VGND_c_3705_n 0.0281312f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1706 N_A_M1003_g N_VGND_c_3707_n 0.00353651f $X=8.795 $Y=0.655 $X2=0 $Y2=0
cc_1707 N_A_M1071_g N_VGND_c_3707_n 0.00464467f $X=9.405 $Y=0.655 $X2=0 $Y2=0
cc_1708 N_A_c_2265_n N_VGND_c_3707_n 0.00644231f $X=11.235 $Y=0.86 $X2=0 $Y2=0
cc_1709 N_A_M1007_g N_VGND_c_3707_n 0.0113729f $X=12.935 $Y=0.655 $X2=0 $Y2=0
cc_1710 N_A_M1041_g N_VGND_c_3707_n 0.0111968f $X=13.46 $Y=0.655 $X2=0 $Y2=0
cc_1711 N_A_c_2275_n N_VGND_c_3707_n 0.0343746f $X=11.647 $Y=0.687 $X2=0 $Y2=0
cc_1712 A N_VGND_c_3707_n 0.0324641f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1713 N_A_M1003_g N_VGND_c_3709_n 0.00241817f $X=8.795 $Y=0.655 $X2=0 $Y2=0
cc_1714 N_A_M1071_g N_VGND_c_3709_n 0.00355956f $X=9.405 $Y=0.655 $X2=0 $Y2=0
cc_1715 N_A_M1003_g N_VGND_c_3710_n 0.00118809f $X=8.795 $Y=0.655 $X2=0 $Y2=0
cc_1716 N_A_M1071_g N_VGND_c_3710_n 0.0105319f $X=9.405 $Y=0.655 $X2=0 $Y2=0
cc_1717 N_A_M1007_g N_A_2519_47#_c_3971_n 0.00963624f $X=12.935 $Y=0.655 $X2=0
+ $Y2=0
cc_1718 N_A_M1041_g N_A_2519_47#_c_3971_n 7.89445e-19 $X=13.46 $Y=0.655 $X2=0
+ $Y2=0
cc_1719 N_A_c_2277_n N_A_2519_47#_c_3971_n 0.00664308f $X=12.365 $Y=0.687 $X2=0
+ $Y2=0
cc_1720 A N_A_2519_47#_c_3971_n 0.0158119f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1721 N_A_M1007_g N_A_2519_47#_c_3956_n 0.0116375f $X=12.935 $Y=0.655 $X2=0
+ $Y2=0
cc_1722 N_A_M1041_g N_A_2519_47#_c_3956_n 0.0157982f $X=13.46 $Y=0.655 $X2=0
+ $Y2=0
cc_1723 N_A_c_2278_n N_A_2519_47#_c_3956_n 7.12423e-19 $X=12.982 $Y=1.65 $X2=0
+ $Y2=0
cc_1724 N_A_c_2267_n N_A_2519_47#_c_3957_n 3.75089e-19 $X=12.86 $Y=1.65 $X2=0
+ $Y2=0
cc_1725 N_A_M1007_g N_A_2519_47#_c_3957_n 0.00236445f $X=12.935 $Y=0.655 $X2=0
+ $Y2=0
cc_1726 N_A_c_2277_n N_A_2519_47#_c_3957_n 0.00198898f $X=12.365 $Y=0.687 $X2=0
+ $Y2=0
cc_1727 N_A_M1007_g N_A_2519_47#_c_3958_n 0.00205246f $X=12.935 $Y=0.655 $X2=0
+ $Y2=0
cc_1728 N_A_c_2277_n N_A_2519_47#_c_3958_n 2.78591e-19 $X=12.365 $Y=0.687 $X2=0
+ $Y2=0
cc_1729 A N_A_2519_47#_c_3958_n 0.00193934f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1730 N_A_2063_47#_c_2495_n N_VPWR_c_2632_n 0.0213669f $X=10.665 $Y=2.01 $X2=0
+ $Y2=0
cc_1731 N_A_2063_47#_c_2496_n N_VPWR_c_2632_n 0.0048356f $X=11.055 $Y=1.93 $X2=0
+ $Y2=0
cc_1732 N_A_2063_47#_c_2495_n N_VPWR_c_2633_n 0.0163084f $X=10.665 $Y=2.01 $X2=0
+ $Y2=0
cc_1733 N_A_2063_47#_c_2495_n N_VPWR_c_2670_n 0.00703609f $X=10.665 $Y=2.01
+ $X2=0 $Y2=0
cc_1734 N_A_2063_47#_c_2495_n N_VPWR_c_2627_n 8.9012e-19 $X=10.665 $Y=2.01 $X2=0
+ $Y2=0
cc_1735 N_A_2063_47#_c_2495_n KAPWR 0.0188316f $X=10.665 $Y=2.01 $X2=0 $Y2=0
cc_1736 N_A_2063_47#_c_2490_n N_A_2345_367#_c_3307_n 0.00445005f $X=13.91
+ $Y=1.44 $X2=0 $Y2=0
cc_1737 N_A_2063_47#_c_2483_n N_VGND_M1065_d 0.00218537f $X=10.97 $Y=0.73 $X2=0
+ $Y2=0
cc_1738 N_A_2063_47#_c_2605_p N_VGND_c_3669_n 0.0115363f $X=10.455 $Y=0.47 $X2=0
+ $Y2=0
cc_1739 N_A_2063_47#_c_2483_n N_VGND_c_3669_n 0.00240763f $X=10.97 $Y=0.73 $X2=0
+ $Y2=0
cc_1740 N_A_2063_47#_c_2483_n N_VGND_c_3670_n 0.0202356f $X=10.97 $Y=0.73 $X2=0
+ $Y2=0
cc_1741 N_A_2063_47#_c_2482_n N_VGND_c_3692_n 0.00359964f $X=14.385 $Y=1.185
+ $X2=0 $Y2=0
cc_1742 N_A_2063_47#_c_2493_n N_VGND_c_3692_n 0.0035993f $X=13.91 $Y=1.185 $X2=0
+ $Y2=0
cc_1743 N_A_2063_47#_c_2483_n N_VGND_c_3705_n 0.001776f $X=10.97 $Y=0.73 $X2=0
+ $Y2=0
cc_1744 N_A_2063_47#_M1020_d N_VGND_c_3707_n 0.00401354f $X=10.315 $Y=0.235
+ $X2=0 $Y2=0
cc_1745 N_A_2063_47#_c_2482_n N_VGND_c_3707_n 0.00665257f $X=14.385 $Y=1.185
+ $X2=0 $Y2=0
cc_1746 N_A_2063_47#_c_2605_p N_VGND_c_3707_n 0.0072329f $X=10.455 $Y=0.47 $X2=0
+ $Y2=0
cc_1747 N_A_2063_47#_c_2483_n N_VGND_c_3707_n 0.0084857f $X=10.97 $Y=0.73 $X2=0
+ $Y2=0
cc_1748 N_A_2063_47#_c_2493_n N_VGND_c_3707_n 0.00552708f $X=13.91 $Y=1.185
+ $X2=0 $Y2=0
cc_1749 N_A_2063_47#_c_2490_n N_A_2519_47#_c_3956_n 0.063271f $X=13.91 $Y=1.44
+ $X2=0 $Y2=0
cc_1750 N_A_2063_47#_c_2492_n N_A_2519_47#_c_3956_n 0.00366108f $X=13.91 $Y=1.26
+ $X2=0 $Y2=0
cc_1751 N_A_2063_47#_c_2493_n N_A_2519_47#_c_3956_n 0.00234543f $X=13.91
+ $Y=1.185 $X2=0 $Y2=0
cc_1752 N_A_2063_47#_c_2487_n N_A_2519_47#_c_3957_n 0.00988015f $X=12.285
+ $Y=1.042 $X2=0 $Y2=0
cc_1753 N_A_2063_47#_c_2490_n N_A_2519_47#_c_3957_n 0.0139193f $X=13.91 $Y=1.44
+ $X2=0 $Y2=0
cc_1754 N_A_2063_47#_c_2493_n N_A_2519_47#_c_3989_n 6.00691e-19 $X=13.91
+ $Y=1.185 $X2=0 $Y2=0
cc_1755 N_A_2063_47#_c_2482_n N_A_2519_47#_c_3990_n 6.41262e-19 $X=14.385
+ $Y=1.185 $X2=0 $Y2=0
cc_1756 N_A_2063_47#_c_2493_n N_A_2519_47#_c_3990_n 0.00785343f $X=13.91
+ $Y=1.185 $X2=0 $Y2=0
cc_1757 N_A_2063_47#_c_2482_n N_A_2519_47#_c_3961_n 0.0105245f $X=14.385
+ $Y=1.185 $X2=0 $Y2=0
cc_1758 N_A_2063_47#_c_2493_n N_A_2519_47#_c_3961_n 0.0105769f $X=13.91 $Y=1.185
+ $X2=0 $Y2=0
cc_1759 N_A_2063_47#_c_2482_n N_A_2519_47#_c_3959_n 0.00511944f $X=14.385
+ $Y=1.185 $X2=0 $Y2=0
cc_1760 N_VPWR_c_2627_n A_228_491# 0.00170373f $X=23.28 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1761 N_VPWR_c_2627_n N_KAPWR_M1035_d 0.00414155f $X=23.28 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1762 N_VPWR_c_2627_n N_KAPWR_M1042_d 0.00127595f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1763 N_VPWR_c_2627_n N_KAPWR_M1066_d 0.00112543f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1764 N_VPWR_M1026_d KAPWR 6.59763e-19 $X=0.65 $Y=2.095 $X2=0 $Y2=0
cc_1765 N_VPWR_M1027_d KAPWR 7.37933e-19 $X=6.65 $Y=2.255 $X2=0 $Y2=0
cc_1766 N_VPWR_M1012_s KAPWR 5.21092e-19 $X=8.735 $Y=1.835 $X2=0 $Y2=0
cc_1767 N_VPWR_M1015_d KAPWR 8.34407e-19 $X=11.31 $Y=1.835 $X2=0 $Y2=0
cc_1768 N_VPWR_M1046_d KAPWR 0.00247367f $X=12.155 $Y=1.835 $X2=0 $Y2=0
cc_1769 N_VPWR_M1010_s KAPWR 7.83613e-19 $X=14.915 $Y=1.835 $X2=0 $Y2=0
cc_1770 N_VPWR_M1019_s KAPWR 0.00204076f $X=15.775 $Y=1.835 $X2=0 $Y2=0
cc_1771 N_VPWR_M1024_s KAPWR 0.00204076f $X=16.635 $Y=1.835 $X2=0 $Y2=0
cc_1772 N_VPWR_M1031_s KAPWR 0.00204076f $X=17.495 $Y=1.835 $X2=0 $Y2=0
cc_1773 N_VPWR_M1034_s KAPWR 0.00204076f $X=18.355 $Y=1.835 $X2=0 $Y2=0
cc_1774 N_VPWR_M1043_s KAPWR 0.00204076f $X=19.215 $Y=1.835 $X2=0 $Y2=0
cc_1775 N_VPWR_M1053_s KAPWR 0.00204076f $X=20.075 $Y=1.835 $X2=0 $Y2=0
cc_1776 N_VPWR_M1060_s KAPWR 0.00204076f $X=20.935 $Y=1.835 $X2=0 $Y2=0
cc_1777 N_VPWR_M1064_s KAPWR 0.00204076f $X=21.795 $Y=1.835 $X2=0 $Y2=0
cc_1778 N_VPWR_M1072_s KAPWR 0.00244555f $X=22.655 $Y=1.835 $X2=0 $Y2=0
cc_1779 N_VPWR_c_2628_n KAPWR 0.0309633f $X=0.79 $Y=2.43 $X2=0 $Y2=0
cc_1780 N_VPWR_c_2629_n KAPWR 0.0269172f $X=5.57 $Y=2.83 $X2=0 $Y2=0
cc_1781 N_VPWR_c_2630_n KAPWR 0.0249891f $X=6.79 $Y=2.6 $X2=0 $Y2=0
cc_1782 N_VPWR_c_2631_n KAPWR 0.0199096f $X=8.875 $Y=2.835 $X2=0 $Y2=0
cc_1783 N_VPWR_c_2632_n KAPWR 0.0353158f $X=9.875 $Y=2.01 $X2=0 $Y2=0
cc_1784 N_VPWR_c_2633_n KAPWR 0.0290786f $X=11.435 $Y=2.485 $X2=0 $Y2=0
cc_1785 N_VPWR_c_2634_n KAPWR 0.00197582f $X=12.2 $Y=3.33 $X2=0 $Y2=0
cc_1786 N_VPWR_c_2635_n KAPWR 0.0152854f $X=12.295 $Y=2.9 $X2=0 $Y2=0
cc_1787 N_VPWR_c_2636_n KAPWR 0.0374775f $X=14.195 $Y=2.27 $X2=0 $Y2=0
cc_1788 N_VPWR_c_2637_n KAPWR 0.022083f $X=15.055 $Y=2.475 $X2=0 $Y2=0
cc_1789 N_VPWR_c_2638_n KAPWR 0.0172617f $X=15.915 $Y=2.455 $X2=0 $Y2=0
cc_1790 N_VPWR_c_2639_n KAPWR 0.0172617f $X=16.775 $Y=2.455 $X2=0 $Y2=0
cc_1791 N_VPWR_c_2640_n KAPWR 0.0172617f $X=17.635 $Y=2.455 $X2=0 $Y2=0
cc_1792 N_VPWR_c_2641_n KAPWR 0.00206353f $X=18.41 $Y=3.33 $X2=0 $Y2=0
cc_1793 N_VPWR_c_2642_n KAPWR 0.0172617f $X=18.495 $Y=2.455 $X2=0 $Y2=0
cc_1794 N_VPWR_c_2643_n KAPWR 0.0172617f $X=19.355 $Y=2.455 $X2=0 $Y2=0
cc_1795 N_VPWR_c_2644_n KAPWR 0.0172617f $X=20.215 $Y=2.455 $X2=0 $Y2=0
cc_1796 N_VPWR_c_2645_n KAPWR 0.0172617f $X=21.075 $Y=2.455 $X2=0 $Y2=0
cc_1797 N_VPWR_c_2646_n KAPWR 0.0172617f $X=21.935 $Y=2.455 $X2=0 $Y2=0
cc_1798 N_VPWR_c_2647_n KAPWR 0.0350235f $X=22.795 $Y=2.455 $X2=0 $Y2=0
cc_1799 N_VPWR_c_2648_n KAPWR 0.00352976f $X=6.705 $Y=3.33 $X2=0 $Y2=0
cc_1800 N_VPWR_c_2650_n KAPWR 0.00194996f $X=14.89 $Y=3.33 $X2=0 $Y2=0
cc_1801 N_VPWR_c_2652_n KAPWR 0.00206353f $X=15.83 $Y=3.33 $X2=0 $Y2=0
cc_1802 N_VPWR_c_2654_n KAPWR 0.00206353f $X=16.69 $Y=3.33 $X2=0 $Y2=0
cc_1803 N_VPWR_c_2656_n KAPWR 0.00206353f $X=17.55 $Y=3.33 $X2=0 $Y2=0
cc_1804 N_VPWR_c_2658_n KAPWR 0.00206353f $X=19.27 $Y=3.33 $X2=0 $Y2=0
cc_1805 N_VPWR_c_2660_n KAPWR 0.00206353f $X=20.13 $Y=3.33 $X2=0 $Y2=0
cc_1806 N_VPWR_c_2662_n KAPWR 0.00206353f $X=20.99 $Y=3.33 $X2=0 $Y2=0
cc_1807 N_VPWR_c_2664_n KAPWR 0.00206353f $X=21.85 $Y=3.33 $X2=0 $Y2=0
cc_1808 N_VPWR_c_2666_n KAPWR 0.00136244f $X=0.625 $Y=3.33 $X2=0 $Y2=0
cc_1809 N_VPWR_c_2667_n KAPWR 0.0114317f $X=5.405 $Y=3.33 $X2=0 $Y2=0
cc_1810 N_VPWR_c_2668_n KAPWR 0.0045498f $X=8.78 $Y=3.33 $X2=0 $Y2=0
cc_1811 N_VPWR_c_2669_n KAPWR 0.00227968f $X=9.71 $Y=3.33 $X2=0 $Y2=0
cc_1812 N_VPWR_c_2670_n KAPWR 0.00579737f $X=11.27 $Y=3.33 $X2=0 $Y2=0
cc_1813 N_VPWR_c_2671_n KAPWR 0.00280393f $X=14.025 $Y=3.33 $X2=0 $Y2=0
cc_1814 N_VPWR_c_2672_n KAPWR 0.00206353f $X=22.71 $Y=3.33 $X2=0 $Y2=0
cc_1815 N_VPWR_c_2673_n KAPWR 0.00262962f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1816 N_VPWR_c_2627_n KAPWR 2.4233f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1817 N_VPWR_c_2667_n N_KAPWR_c_3047_n 0.0604494f $X=5.405 $Y=3.33 $X2=0 $Y2=0
cc_1818 N_VPWR_c_2627_n N_KAPWR_c_3047_n 0.008401f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1819 N_VPWR_c_2667_n N_KAPWR_c_3065_n 0.0122542f $X=5.405 $Y=3.33 $X2=0 $Y2=0
cc_1820 N_VPWR_c_2627_n N_KAPWR_c_3065_n 0.00238443f $X=23.28 $Y=3.33 $X2=0
+ $Y2=0
cc_1821 N_VPWR_c_2629_n N_KAPWR_c_3048_n 0.0235402f $X=5.57 $Y=2.83 $X2=0 $Y2=0
cc_1822 N_VPWR_c_2667_n N_KAPWR_c_3048_n 0.014625f $X=5.405 $Y=3.33 $X2=0 $Y2=0
cc_1823 N_VPWR_c_2627_n N_KAPWR_c_3048_n 0.00294717f $X=23.28 $Y=3.33 $X2=0
+ $Y2=0
cc_1824 N_VPWR_c_2627_n A_1172_451# 0.00128403f $X=23.28 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1825 N_VPWR_c_2627_n N_A_1492_367#_M1023_s 0.00126783f $X=23.28 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_1826 N_VPWR_c_2627_n N_A_1492_367#_M1067_s 0.00113524f $X=23.28 $Y=3.33 $X2=0
+ $Y2=0
cc_1827 N_VPWR_c_2627_n N_A_1492_367#_M1044_d 0.00116866f $X=23.28 $Y=3.33 $X2=0
+ $Y2=0
cc_1828 N_VPWR_c_2630_n N_A_1492_367#_c_3248_n 0.00534048f $X=6.79 $Y=2.6 $X2=0
+ $Y2=0
cc_1829 N_VPWR_c_2668_n N_A_1492_367#_c_3248_n 0.0145445f $X=8.78 $Y=3.33 $X2=0
+ $Y2=0
cc_1830 N_VPWR_c_2627_n N_A_1492_367#_c_3248_n 0.00231855f $X=23.28 $Y=3.33
+ $X2=0 $Y2=0
cc_1831 N_VPWR_c_2630_n N_A_1492_367#_c_3237_n 0.0122501f $X=6.79 $Y=2.6 $X2=0
+ $Y2=0
cc_1832 N_VPWR_c_2668_n N_A_1492_367#_c_3255_n 0.0280869f $X=8.78 $Y=3.33 $X2=0
+ $Y2=0
cc_1833 N_VPWR_c_2627_n N_A_1492_367#_c_3255_n 0.00406229f $X=23.28 $Y=3.33
+ $X2=0 $Y2=0
cc_1834 N_VPWR_c_2631_n N_A_1492_367#_c_3258_n 0.0188707f $X=8.875 $Y=2.835
+ $X2=0 $Y2=0
cc_1835 N_VPWR_c_2668_n N_A_1492_367#_c_3258_n 0.0179231f $X=8.78 $Y=3.33 $X2=0
+ $Y2=0
cc_1836 N_VPWR_c_2627_n N_A_1492_367#_c_3258_n 0.00303682f $X=23.28 $Y=3.33
+ $X2=0 $Y2=0
cc_1837 N_VPWR_M1012_s N_A_1492_367#_c_3244_n 0.00308831f $X=8.735 $Y=1.835
+ $X2=0 $Y2=0
cc_1838 N_VPWR_c_2631_n N_A_1492_367#_c_3244_n 0.013575f $X=8.875 $Y=2.835 $X2=0
+ $Y2=0
cc_1839 N_VPWR_c_2631_n N_A_1492_367#_c_3239_n 0.0181395f $X=8.875 $Y=2.835
+ $X2=0 $Y2=0
cc_1840 N_VPWR_c_2632_n N_A_1492_367#_c_3239_n 0.0452137f $X=9.875 $Y=2.01 $X2=0
+ $Y2=0
cc_1841 N_VPWR_c_2669_n N_A_1492_367#_c_3239_n 0.0167395f $X=9.71 $Y=3.33 $X2=0
+ $Y2=0
cc_1842 N_VPWR_c_2627_n N_A_1492_367#_c_3239_n 0.00244519f $X=23.28 $Y=3.33
+ $X2=0 $Y2=0
cc_1843 N_VPWR_c_2627_n N_A_2345_367#_M1015_s 0.00114229f $X=23.28 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_1844 N_VPWR_c_2627_n N_A_2345_367#_M1016_s 0.00110569f $X=23.28 $Y=3.33 $X2=0
+ $Y2=0
cc_1845 N_VPWR_c_2627_n N_A_2345_367#_M1069_s 0.0011057f $X=23.28 $Y=3.33 $X2=0
+ $Y2=0
cc_1846 N_VPWR_M1046_d N_A_2345_367#_c_3306_n 0.00665866f $X=12.155 $Y=1.835
+ $X2=0 $Y2=0
cc_1847 N_VPWR_c_2635_n N_A_2345_367#_c_3306_n 0.0110201f $X=12.295 $Y=2.9 $X2=0
+ $Y2=0
cc_1848 N_VPWR_c_2635_n N_A_2345_367#_c_3308_n 0.00253838f $X=12.295 $Y=2.9
+ $X2=0 $Y2=0
cc_1849 N_VPWR_c_2671_n N_A_2345_367#_c_3327_n 0.0344117f $X=14.025 $Y=3.33
+ $X2=0 $Y2=0
cc_1850 N_VPWR_c_2627_n N_A_2345_367#_c_3327_n 0.00493963f $X=23.28 $Y=3.33
+ $X2=0 $Y2=0
cc_1851 N_VPWR_c_2635_n N_A_2345_367#_c_3309_n 0.0215602f $X=12.295 $Y=2.9 $X2=0
+ $Y2=0
cc_1852 N_VPWR_c_2671_n N_A_2345_367#_c_3309_n 0.0211865f $X=14.025 $Y=3.33
+ $X2=0 $Y2=0
cc_1853 N_VPWR_c_2627_n N_A_2345_367#_c_3309_n 0.00305633f $X=23.28 $Y=3.33
+ $X2=0 $Y2=0
cc_1854 N_VPWR_c_2636_n N_A_2345_367#_c_3310_n 0.0222939f $X=14.195 $Y=2.27
+ $X2=0 $Y2=0
cc_1855 N_VPWR_c_2671_n N_A_2345_367#_c_3310_n 0.0175634f $X=14.025 $Y=3.33
+ $X2=0 $Y2=0
cc_1856 N_VPWR_c_2627_n N_A_2345_367#_c_3310_n 0.0023387f $X=23.28 $Y=3.33 $X2=0
+ $Y2=0
cc_1857 N_VPWR_c_2636_n N_A_2345_367#_c_3311_n 0.0442579f $X=14.195 $Y=2.27
+ $X2=0 $Y2=0
cc_1858 N_VPWR_c_2633_n N_A_2345_367#_c_3318_n 0.023916f $X=11.435 $Y=2.485
+ $X2=0 $Y2=0
cc_1859 N_VPWR_c_2634_n N_A_2345_367#_c_3318_n 0.0151334f $X=12.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1860 N_VPWR_c_2635_n N_A_2345_367#_c_3318_n 0.0139819f $X=12.295 $Y=2.9 $X2=0
+ $Y2=0
cc_1861 N_VPWR_c_2627_n N_A_2345_367#_c_3318_n 0.00309906f $X=23.28 $Y=3.33
+ $X2=0 $Y2=0
cc_1862 N_VPWR_c_2627_n N_Z_M1004_d 0.00157848f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1863 N_VPWR_c_2627_n N_Z_M1017_d 0.00113524f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1864 N_VPWR_c_2627_n N_Z_M1022_d 0.00113524f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1865 N_VPWR_c_2627_n N_Z_M1028_d 0.00113524f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1866 N_VPWR_c_2627_n N_Z_M1033_d 0.00113524f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1867 N_VPWR_c_2627_n N_Z_M1039_d 0.00113524f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1868 N_VPWR_c_2627_n N_Z_M1051_d 0.00113524f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1869 N_VPWR_c_2627_n N_Z_M1054_d 0.00113524f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1870 N_VPWR_c_2627_n N_Z_M1061_d 0.00113524f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1871 N_VPWR_c_2627_n N_Z_M1070_d 0.00113524f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1872 N_VPWR_c_2636_n N_Z_c_3564_n 0.0366036f $X=14.195 $Y=2.27 $X2=0 $Y2=0
cc_1873 N_VPWR_c_2637_n N_Z_c_3564_n 0.0294041f $X=15.055 $Y=2.475 $X2=0 $Y2=0
cc_1874 N_VPWR_c_2650_n N_Z_c_3564_n 0.0110337f $X=14.89 $Y=3.33 $X2=0 $Y2=0
cc_1875 N_VPWR_c_2627_n N_Z_c_3564_n 0.00158132f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1876 N_VPWR_M1010_s N_Z_c_3379_n 0.00278715f $X=14.915 $Y=1.835 $X2=0 $Y2=0
cc_1877 N_VPWR_c_2637_n N_Z_c_3379_n 0.0135053f $X=15.055 $Y=2.475 $X2=0 $Y2=0
cc_1878 N_VPWR_c_2637_n N_Z_c_3393_n 0.0302022f $X=15.055 $Y=2.475 $X2=0 $Y2=0
cc_1879 N_VPWR_c_2638_n N_Z_c_3393_n 0.030864f $X=15.915 $Y=2.455 $X2=0 $Y2=0
cc_1880 N_VPWR_c_2652_n N_Z_c_3393_n 0.0177952f $X=15.83 $Y=3.33 $X2=0 $Y2=0
cc_1881 N_VPWR_c_2627_n N_Z_c_3393_n 0.00302007f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1882 N_VPWR_c_2638_n N_Z_c_3368_n 0.030864f $X=15.915 $Y=2.455 $X2=0 $Y2=0
cc_1883 N_VPWR_c_2639_n N_Z_c_3368_n 0.030864f $X=16.775 $Y=2.455 $X2=0 $Y2=0
cc_1884 N_VPWR_c_2654_n N_Z_c_3368_n 0.0177952f $X=16.69 $Y=3.33 $X2=0 $Y2=0
cc_1885 N_VPWR_c_2627_n N_Z_c_3368_n 0.00302007f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1886 N_VPWR_c_2639_n N_Z_c_3369_n 0.030864f $X=16.775 $Y=2.455 $X2=0 $Y2=0
cc_1887 N_VPWR_c_2640_n N_Z_c_3369_n 0.030864f $X=17.635 $Y=2.455 $X2=0 $Y2=0
cc_1888 N_VPWR_c_2656_n N_Z_c_3369_n 0.0177952f $X=17.55 $Y=3.33 $X2=0 $Y2=0
cc_1889 N_VPWR_c_2627_n N_Z_c_3369_n 0.00302007f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1890 N_VPWR_c_2640_n N_Z_c_3370_n 0.030864f $X=17.635 $Y=2.455 $X2=0 $Y2=0
cc_1891 N_VPWR_c_2641_n N_Z_c_3370_n 0.0177952f $X=18.41 $Y=3.33 $X2=0 $Y2=0
cc_1892 N_VPWR_c_2642_n N_Z_c_3370_n 0.030864f $X=18.495 $Y=2.455 $X2=0 $Y2=0
cc_1893 N_VPWR_c_2627_n N_Z_c_3370_n 0.00302007f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1894 N_VPWR_c_2642_n N_Z_c_3371_n 0.030864f $X=18.495 $Y=2.455 $X2=0 $Y2=0
cc_1895 N_VPWR_c_2643_n N_Z_c_3371_n 0.030864f $X=19.355 $Y=2.455 $X2=0 $Y2=0
cc_1896 N_VPWR_c_2658_n N_Z_c_3371_n 0.0177952f $X=19.27 $Y=3.33 $X2=0 $Y2=0
cc_1897 N_VPWR_c_2627_n N_Z_c_3371_n 0.00302007f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1898 N_VPWR_c_2643_n N_Z_c_3372_n 0.030864f $X=19.355 $Y=2.455 $X2=0 $Y2=0
cc_1899 N_VPWR_c_2644_n N_Z_c_3372_n 0.030864f $X=20.215 $Y=2.455 $X2=0 $Y2=0
cc_1900 N_VPWR_c_2660_n N_Z_c_3372_n 0.0177952f $X=20.13 $Y=3.33 $X2=0 $Y2=0
cc_1901 N_VPWR_c_2627_n N_Z_c_3372_n 0.00302007f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1902 N_VPWR_c_2644_n N_Z_c_3373_n 0.030864f $X=20.215 $Y=2.455 $X2=0 $Y2=0
cc_1903 N_VPWR_c_2645_n N_Z_c_3373_n 0.030864f $X=21.075 $Y=2.455 $X2=0 $Y2=0
cc_1904 N_VPWR_c_2662_n N_Z_c_3373_n 0.0177952f $X=20.99 $Y=3.33 $X2=0 $Y2=0
cc_1905 N_VPWR_c_2627_n N_Z_c_3373_n 0.00302007f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1906 N_VPWR_c_2645_n N_Z_c_3374_n 0.030864f $X=21.075 $Y=2.455 $X2=0 $Y2=0
cc_1907 N_VPWR_c_2646_n N_Z_c_3374_n 0.030864f $X=21.935 $Y=2.455 $X2=0 $Y2=0
cc_1908 N_VPWR_c_2664_n N_Z_c_3374_n 0.0177952f $X=21.85 $Y=3.33 $X2=0 $Y2=0
cc_1909 N_VPWR_c_2627_n N_Z_c_3374_n 0.00302007f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1910 N_VPWR_c_2646_n N_Z_c_3454_n 0.030864f $X=21.935 $Y=2.455 $X2=0 $Y2=0
cc_1911 N_VPWR_c_2647_n N_Z_c_3454_n 0.030919f $X=22.795 $Y=2.455 $X2=0 $Y2=0
cc_1912 N_VPWR_c_2672_n N_Z_c_3454_n 0.0177952f $X=22.71 $Y=3.33 $X2=0 $Y2=0
cc_1913 N_VPWR_c_2627_n N_Z_c_3454_n 0.00302007f $X=23.28 $Y=3.33 $X2=0 $Y2=0
cc_1914 N_VPWR_M1010_s N_Z_c_3460_n 0.00408427f $X=14.915 $Y=1.835 $X2=0 $Y2=0
cc_1915 N_VPWR_M1019_s N_Z_c_3460_n 0.00446486f $X=15.775 $Y=1.835 $X2=0 $Y2=0
cc_1916 N_VPWR_M1024_s N_Z_c_3460_n 0.00446486f $X=16.635 $Y=1.835 $X2=0 $Y2=0
cc_1917 N_VPWR_M1031_s N_Z_c_3460_n 0.00446486f $X=17.495 $Y=1.835 $X2=0 $Y2=0
cc_1918 N_VPWR_M1034_s N_Z_c_3460_n 0.00446486f $X=18.355 $Y=1.835 $X2=0 $Y2=0
cc_1919 N_VPWR_M1043_s N_Z_c_3460_n 0.00428354f $X=19.215 $Y=1.835 $X2=0 $Y2=0
cc_1920 N_VPWR_M1053_s N_Z_c_3460_n 0.00428354f $X=20.075 $Y=1.835 $X2=0 $Y2=0
cc_1921 N_VPWR_M1060_s N_Z_c_3460_n 0.00428354f $X=20.935 $Y=1.835 $X2=0 $Y2=0
cc_1922 N_VPWR_M1064_s N_Z_c_3460_n 0.00411203f $X=21.795 $Y=1.835 $X2=0 $Y2=0
cc_1923 N_VPWR_c_2636_n N_Z_c_3460_n 4.67603e-19 $X=14.195 $Y=2.27 $X2=0 $Y2=0
cc_1924 N_VPWR_c_2637_n N_Z_c_3460_n 0.00306514f $X=15.055 $Y=2.475 $X2=0 $Y2=0
cc_1925 N_VPWR_c_2638_n N_Z_c_3460_n 0.00667189f $X=15.915 $Y=2.455 $X2=0 $Y2=0
cc_1926 N_VPWR_c_2639_n N_Z_c_3460_n 0.00667189f $X=16.775 $Y=2.455 $X2=0 $Y2=0
cc_1927 N_VPWR_c_2640_n N_Z_c_3460_n 0.00667189f $X=17.635 $Y=2.455 $X2=0 $Y2=0
cc_1928 N_VPWR_c_2642_n N_Z_c_3460_n 0.00667189f $X=18.495 $Y=2.455 $X2=0 $Y2=0
cc_1929 N_VPWR_c_2643_n N_Z_c_3460_n 0.00329183f $X=19.355 $Y=2.455 $X2=0 $Y2=0
cc_1930 N_VPWR_c_2644_n N_Z_c_3460_n 0.00329183f $X=20.215 $Y=2.455 $X2=0 $Y2=0
cc_1931 N_VPWR_c_2645_n N_Z_c_3460_n 0.00329183f $X=21.075 $Y=2.455 $X2=0 $Y2=0
cc_1932 N_VPWR_c_2646_n N_Z_c_3460_n 0.00329183f $X=21.935 $Y=2.455 $X2=0 $Y2=0
cc_1933 A_228_491# KAPWR 0.00407501f $X=1.14 $Y=2.455 $X2=15.775 $Y2=1.835
cc_1934 KAPWR A_1172_451# 0.00255125f $X=0.07 $Y=2.675 $X2=-0.19 $Y2=1.655
cc_1935 KAPWR N_A_1492_367#_M1023_s 7.90696e-19 $X=0.07 $Y=2.675 $X2=-0.19
+ $Y2=1.655
cc_1936 KAPWR N_A_1492_367#_M1044_d 5.21092e-19 $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1937 KAPWR N_A_1492_367#_c_3248_n 0.004468f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1938 KAPWR N_A_1492_367#_c_3237_n 0.0225426f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1939 KAPWR N_A_1492_367#_c_3255_n 0.0159925f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1940 KAPWR N_A_1492_367#_c_3258_n 0.0288558f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1941 KAPWR N_A_1492_367#_c_3244_n 0.0107217f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1942 KAPWR N_A_1492_367#_c_3239_n 0.0226892f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1943 KAPWR A_2033_373# 0.00304573f $X=0.07 $Y=2.675 $X2=-0.19 $Y2=1.655
cc_1944 KAPWR N_A_2345_367#_M1069_s 0.00218578f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1945 KAPWR N_A_2345_367#_c_3306_n 0.0237469f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1946 KAPWR N_A_2345_367#_c_3308_n 0.0247828f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1947 KAPWR N_A_2345_367#_c_3327_n 0.0239751f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1948 KAPWR N_A_2345_367#_c_3309_n 0.0109089f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1949 KAPWR N_A_2345_367#_c_3310_n 0.00867691f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1950 KAPWR N_A_2345_367#_c_3311_n 0.0190984f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1951 KAPWR N_A_2345_367#_c_3318_n 0.025488f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1952 KAPWR N_Z_M1004_d 0.0017802f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1953 KAPWR N_Z_c_3564_n 0.0168728f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1954 KAPWR N_Z_c_3379_n 0.00371135f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1955 KAPWR N_Z_c_3393_n 0.0271478f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1956 KAPWR N_Z_c_3368_n 0.0271478f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1957 KAPWR N_Z_c_3369_n 0.0271478f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1958 KAPWR N_Z_c_3370_n 0.0271478f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1959 KAPWR N_Z_c_3371_n 0.0271478f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1960 KAPWR N_Z_c_3372_n 0.0271478f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1961 KAPWR N_Z_c_3373_n 0.0271478f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1962 KAPWR N_Z_c_3374_n 0.0271478f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1963 KAPWR N_Z_c_3454_n 0.0276761f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1964 KAPWR N_Z_c_3460_n 0.371306f $X=0.07 $Y=2.675 $X2=0 $Y2=0
cc_1965 N_Z_c_3370_n N_VGND_c_3675_n 0.0189236f $X=18.065 $Y=0.36 $X2=0 $Y2=0
cc_1966 N_Z_c_3367_n N_VGND_c_3692_n 0.0210192f $X=15.485 $Y=0.36 $X2=0 $Y2=0
cc_1967 N_Z_c_3368_n N_VGND_c_3694_n 0.0189236f $X=16.345 $Y=0.36 $X2=0 $Y2=0
cc_1968 N_Z_c_3369_n N_VGND_c_3696_n 0.0189236f $X=17.205 $Y=0.36 $X2=0 $Y2=0
cc_1969 N_Z_c_3371_n N_VGND_c_3698_n 0.0189236f $X=18.925 $Y=0.36 $X2=0 $Y2=0
cc_1970 N_Z_c_3372_n N_VGND_c_3700_n 0.0189236f $X=19.785 $Y=0.36 $X2=0 $Y2=0
cc_1971 N_Z_c_3373_n N_VGND_c_3702_n 0.0183421f $X=20.645 $Y=0.36 $X2=0 $Y2=0
cc_1972 N_Z_c_3374_n N_VGND_c_3706_n 0.0210192f $X=21.505 $Y=0.36 $X2=0 $Y2=0
cc_1973 N_Z_M1000_s N_VGND_c_3707_n 0.00231914f $X=15.34 $Y=0.235 $X2=0 $Y2=0
cc_1974 N_Z_M1009_s N_VGND_c_3707_n 0.00223559f $X=16.205 $Y=0.235 $X2=0 $Y2=0
cc_1975 N_Z_M1025_s N_VGND_c_3707_n 0.00223559f $X=17.065 $Y=0.235 $X2=0 $Y2=0
cc_1976 N_Z_M1032_s N_VGND_c_3707_n 0.00223559f $X=17.925 $Y=0.235 $X2=0 $Y2=0
cc_1977 N_Z_M1048_s N_VGND_c_3707_n 0.00223559f $X=18.785 $Y=0.235 $X2=0 $Y2=0
cc_1978 N_Z_M1056_s N_VGND_c_3707_n 0.00223559f $X=19.645 $Y=0.235 $X2=0 $Y2=0
cc_1979 N_Z_M1059_s N_VGND_c_3707_n 0.00223667f $X=20.505 $Y=0.235 $X2=0 $Y2=0
cc_1980 N_Z_M1073_s N_VGND_c_3707_n 0.00231914f $X=21.365 $Y=0.235 $X2=0 $Y2=0
cc_1981 N_Z_c_3367_n N_VGND_c_3707_n 0.0125689f $X=15.485 $Y=0.36 $X2=0 $Y2=0
cc_1982 N_Z_c_3368_n N_VGND_c_3707_n 0.0123859f $X=16.345 $Y=0.36 $X2=0 $Y2=0
cc_1983 N_Z_c_3369_n N_VGND_c_3707_n 0.0123859f $X=17.205 $Y=0.36 $X2=0 $Y2=0
cc_1984 N_Z_c_3370_n N_VGND_c_3707_n 0.0123859f $X=18.065 $Y=0.36 $X2=0 $Y2=0
cc_1985 N_Z_c_3371_n N_VGND_c_3707_n 0.0123859f $X=18.925 $Y=0.36 $X2=0 $Y2=0
cc_1986 N_Z_c_3372_n N_VGND_c_3707_n 0.0123859f $X=19.785 $Y=0.36 $X2=0 $Y2=0
cc_1987 N_Z_c_3373_n N_VGND_c_3707_n 0.0123555f $X=20.645 $Y=0.36 $X2=0 $Y2=0
cc_1988 N_Z_c_3374_n N_VGND_c_3707_n 0.0125689f $X=21.505 $Y=0.36 $X2=0 $Y2=0
cc_1989 N_Z_c_3367_n N_A_2519_47#_c_3959_n 0.0290655f $X=15.485 $Y=0.36 $X2=0
+ $Y2=0
cc_1990 A_110_47# N_VGND_c_3707_n 0.00899413f $X=0.55 $Y=0.235 $X2=23.28 $Y2=0
cc_1991 N_VGND_c_3707_n A_1053_47# 0.00176519f $X=23.28 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1992 N_VGND_c_3707_n N_A_2519_47#_M1007_s 0.00217209f $X=23.28 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1993 N_VGND_c_3707_n N_A_2519_47#_M1041_s 0.00416069f $X=23.28 $Y=0 $X2=0
+ $Y2=0
cc_1994 N_VGND_c_3707_n N_A_2519_47#_M1055_d 0.00253158f $X=23.28 $Y=0 $X2=0
+ $Y2=0
cc_1995 N_VGND_M1007_d N_A_2519_47#_c_3956_n 0.00289819f $X=13.01 $Y=0.235 $X2=0
+ $Y2=0
cc_1996 N_VGND_c_3671_n N_A_2519_47#_c_3956_n 0.0203217f $X=13.205 $Y=0.59 $X2=0
+ $Y2=0
cc_1997 N_VGND_c_3692_n N_A_2519_47#_c_3989_n 0.0193086f $X=15.83 $Y=0 $X2=0
+ $Y2=0
cc_1998 N_VGND_c_3707_n N_A_2519_47#_c_3989_n 0.0125808f $X=23.28 $Y=0 $X2=0
+ $Y2=0
cc_1999 N_VGND_c_3692_n N_A_2519_47#_c_3961_n 0.0327749f $X=15.83 $Y=0 $X2=0
+ $Y2=0
cc_2000 N_VGND_c_3707_n N_A_2519_47#_c_3961_n 0.022395f $X=23.28 $Y=0 $X2=0
+ $Y2=0
cc_2001 N_VGND_c_3705_n N_A_2519_47#_c_3958_n 0.0154057f $X=13.055 $Y=0 $X2=0
+ $Y2=0
cc_2002 N_VGND_c_3707_n N_A_2519_47#_c_3958_n 0.0119195f $X=23.28 $Y=0 $X2=0
+ $Y2=0
cc_2003 N_VGND_c_3692_n N_A_2519_47#_c_3959_n 0.0165434f $X=15.83 $Y=0 $X2=0
+ $Y2=0
cc_2004 N_VGND_c_3707_n N_A_2519_47#_c_3959_n 0.00967329f $X=23.28 $Y=0 $X2=0
+ $Y2=0
