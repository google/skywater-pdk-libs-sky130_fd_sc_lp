* File: sky130_fd_sc_lp__dlclkp_lp.pex.spice
* Created: Wed Sep  2 09:46:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%A_80_21# 1 2 9 13 17 21 25 27 30 32 33 36
+ 37 40 42 48 51 55 57
c150 57 0 2.16197e-19 $X=4.815 $Y=2.48
c151 37 0 1.88043e-19 $X=2.545 $Y=1.615
r152 59 60 17.0922 $w=2.82e-07 $l=1e-07 $layer=POLY_cond $X=0.475 $Y=1.23
+ $X2=0.575 $Y2=1.23
r153 54 57 12.7703 $w=3.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.405 $Y=2.5
+ $X2=4.815 $Y2=2.5
r154 54 55 6.04704 $w=3.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=2.5
+ $X2=4.32 $Y2=2.5
r155 48 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.645 $Y=1.285
+ $X2=1.645 $Y2=1.12
r156 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.645
+ $Y=1.285 $X2=1.645 $Y2=1.285
r157 42 54 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.405 $Y=2.315
+ $X2=4.405 $Y2=2.5
r158 41 51 2.99516 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=4.405 $Y=1.145
+ $X2=4.325 $Y2=1.02
r159 41 42 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.405 $Y=1.145
+ $X2=4.405 $Y2=2.315
r160 40 55 163.754 $w=1.68e-07 $l=2.51e-06 $layer=LI1_cond $X=1.81 $Y=2.6
+ $X2=4.32 $Y2=2.6
r161 37 68 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.545 $Y=1.615
+ $X2=2.545 $Y2=1.78
r162 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.545
+ $Y=1.615 $X2=2.545 $Y2=1.615
r163 34 47 15.7266 $w=2.56e-07 $l=3.3e-07 $layer=LI1_cond $X=1.645 $Y=1.615
+ $X2=1.645 $Y2=1.285
r164 34 36 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=1.81 $Y=1.615
+ $X2=2.545 $Y2=1.615
r165 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.725 $Y=2.515
+ $X2=1.81 $Y2=2.6
r166 32 34 9.24244 $w=2.56e-07 $l=2.0106e-07 $layer=LI1_cond $X=1.725 $Y=1.78
+ $X2=1.645 $Y2=1.615
r167 32 33 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.725 $Y=1.78
+ $X2=1.725 $Y2=2.515
r168 30 60 5.98227 $w=2.82e-07 $l=3.5e-08 $layer=POLY_cond $X=0.61 $Y=1.23
+ $X2=0.575 $Y2=1.23
r169 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.23 $X2=0.61 $Y2=1.23
r170 27 47 2.62109 $w=2.56e-07 $l=5.5e-08 $layer=LI1_cond $X=1.645 $Y=1.23
+ $X2=1.645 $Y2=1.285
r171 27 29 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=1.48 $Y=1.23
+ $X2=0.61 $Y2=1.23
r172 25 68 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.505 $Y=2.595
+ $X2=2.505 $Y2=1.78
r173 21 64 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.735 $Y=0.445
+ $X2=1.735 $Y2=1.12
r174 15 30 38.4574 $w=2.82e-07 $l=2.96226e-07 $layer=POLY_cond $X=0.835 $Y=1.065
+ $X2=0.61 $Y2=1.23
r175 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.835 $Y=1.065
+ $X2=0.835 $Y2=0.445
r176 11 60 5.69241 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.395
+ $X2=0.575 $Y2=1.23
r177 11 13 298.144 $w=2.5e-07 $l=1.2e-06 $layer=POLY_cond $X=0.575 $Y=1.395
+ $X2=0.575 $Y2=2.595
r178 7 59 17.5183 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.065
+ $X2=0.475 $Y2=1.23
r179 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.475 $Y=1.065
+ $X2=0.475 $Y2=0.445
r180 2 57 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=4.67
+ $Y=2.095 $X2=4.815 $Y2=2.48
r181 1 51 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.18
+ $Y=0.925 $X2=4.325 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%GATE 3 7 9 12 14 17 18 19
c48 12 0 1.88697e-19 $X=1.345 $Y=0.805
r49 17 20 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.77
+ $X2=1.105 $Y2=1.935
r50 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.77
+ $X2=1.105 $Y2=1.605
r51 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=1.77 $X2=1.105 $Y2=1.77
r52 14 18 8.44936 $w=5.43e-07 $l=3.85e-07 $layer=LI1_cond $X=0.72 $Y=1.877
+ $X2=1.105 $Y2=1.877
r53 10 12 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.195 $Y=0.805
+ $X2=1.345 $Y2=0.805
r54 7 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.345 $Y=0.73
+ $X2=1.345 $Y2=0.805
r55 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.345 $Y=0.73 $X2=1.345
+ $Y2=0.445
r56 5 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.195 $Y=0.88
+ $X2=1.195 $Y2=0.805
r57 5 19 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=1.195 $Y=0.88
+ $X2=1.195 $Y2=1.605
r58 3 20 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.145 $Y=2.595
+ $X2=1.145 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%A_27_47# 1 2 9 11 12 13 14 15 17 20 26 28
+ 30 31 32
c89 32 0 1.88043e-19 $X=2.255 $Y=0.8
r90 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.255
+ $Y=0.93 $X2=2.255 $Y2=0.93
r91 32 35 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.255 $Y=0.8
+ $X2=2.255 $Y2=0.93
r92 30 31 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.285 $Y=2.495
+ $X2=0.285 $Y2=2.33
r93 27 28 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=0.8
+ $X2=0.26 $Y2=0.8
r94 26 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=0.8
+ $X2=2.255 $Y2=0.8
r95 26 27 108.626 $w=1.68e-07 $l=1.665e-06 $layer=LI1_cond $X=2.09 $Y=0.8
+ $X2=0.425 $Y2=0.8
r96 22 28 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.18 $Y=0.885
+ $X2=0.26 $Y2=0.8
r97 22 31 94.2727 $w=1.68e-07 $l=1.445e-06 $layer=LI1_cond $X=0.18 $Y=0.885
+ $X2=0.18 $Y2=2.33
r98 18 28 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.715
+ $X2=0.26 $Y2=0.8
r99 18 20 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.26 $Y=0.715
+ $X2=0.26 $Y2=0.47
r100 15 36 38.924 $w=3.61e-07 $l=1.90526e-07 $layer=POLY_cond $X=2.165 $Y=0.765
+ $X2=2.22 $Y2=0.93
r101 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.165 $Y=0.765
+ $X2=2.165 $Y2=0.445
r102 13 36 38.924 $w=3.61e-07 $l=2.18746e-07 $layer=POLY_cond $X=2.095 $Y=1.095
+ $X2=2.22 $Y2=0.93
r103 13 14 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=2.095 $Y=1.095
+ $X2=2.095 $Y2=1.69
r104 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.02 $Y=1.765
+ $X2=2.095 $Y2=1.69
r105 11 12 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=2.02 $Y=1.765
+ $X2=1.76 $Y2=1.765
r106 7 12 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=1.635 $Y=1.84
+ $X2=1.76 $Y2=1.765
r107 7 9 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.635 $Y=1.84
+ $X2=1.635 $Y2=2.595
r108 2 30 300 $w=1.7e-07 $l=4.66905e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.095 $X2=0.31 $Y2=2.495
r109 1 20 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%A_584_21# 1 2 9 13 15 17 20 22 25 27 28 31
+ 32 33 36 37 39 43 48 54 56
c160 37 0 3.57943e-19 $X=6.11 $Y=1.71
c161 36 0 1.04487e-19 $X=6.11 $Y=1.71
c162 31 0 1.54238e-19 $X=4.755 $Y=1.965
c163 15 0 2.81132e-20 $X=5.835 $Y=1.42
r164 55 56 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.895 $Y=1.41
+ $X2=4.055 $Y2=1.41
r165 53 54 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=4.03 $Y=0.47
+ $X2=4.195 $Y2=0.47
r166 50 53 3.79463 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=3.895 $Y=0.47
+ $X2=4.03 $Y2=0.47
r167 46 48 6.77778 $w=1.78e-07 $l=1.1e-07 $layer=LI1_cond $X=3.945 $Y=2.245
+ $X2=4.055 $Y2=2.245
r168 43 60 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.55
+ $X2=3.085 $Y2=1.715
r169 43 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.55
+ $X2=3.085 $Y2=1.385
r170 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.085
+ $Y=1.55 $X2=3.085 $Y2=1.55
r171 39 42 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.085 $Y=1.41
+ $X2=3.085 $Y2=1.55
r172 37 63 4.1913 $w=3.45e-07 $l=3e-08 $layer=POLY_cond $X=6.11 $Y=1.647
+ $X2=6.14 $Y2=1.647
r173 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.11
+ $Y=1.71 $X2=6.11 $Y2=1.71
r174 34 36 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.11 $Y=1.965
+ $X2=6.11 $Y2=1.71
r175 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.945 $Y=2.05
+ $X2=6.11 $Y2=1.965
r176 32 33 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=5.945 $Y=2.05
+ $X2=4.84 $Y2=2.05
r177 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.755 $Y=1.965
+ $X2=4.84 $Y2=2.05
r178 30 31 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.755 $Y=0.675
+ $X2=4.755 $Y2=1.965
r179 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.67 $Y=0.59
+ $X2=4.755 $Y2=0.675
r180 28 54 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.67 $Y=0.59
+ $X2=4.195 $Y2=0.59
r181 27 48 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.055 $Y=2.155
+ $X2=4.055 $Y2=2.245
r182 26 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=1.495
+ $X2=4.055 $Y2=1.41
r183 26 27 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.055 $Y=1.495
+ $X2=4.055 $Y2=2.155
r184 25 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=1.325
+ $X2=3.895 $Y2=1.41
r185 24 50 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.895 $Y=0.675
+ $X2=3.895 $Y2=0.47
r186 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.895 $Y=0.675
+ $X2=3.895 $Y2=1.325
r187 23 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=1.41
+ $X2=3.085 $Y2=1.41
r188 22 55 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.81 $Y=1.41
+ $X2=3.895 $Y2=1.41
r189 22 23 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.81 $Y=1.41
+ $X2=3.25 $Y2=1.41
r190 18 63 10.3696 $w=2.5e-07 $l=2.28e-07 $layer=POLY_cond $X=6.14 $Y=1.875
+ $X2=6.14 $Y2=1.647
r191 18 20 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=6.14 $Y=1.875
+ $X2=6.14 $Y2=2.595
r192 15 37 38.4203 $w=3.45e-07 $l=3.71551e-07 $layer=POLY_cond $X=5.835 $Y=1.42
+ $X2=6.11 $Y2=1.647
r193 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.835 $Y=1.42
+ $X2=5.835 $Y2=1.135
r194 13 60 218.639 $w=2.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.075 $Y=2.595
+ $X2=3.075 $Y2=1.715
r195 9 59 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.995 $Y=0.445 $X2=2.995
+ $Y2=1.385
r196 2 46 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=2.095 $X2=3.945 $Y2=2.245
r197 1 53 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.89
+ $Y=0.235 $X2=4.03 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%A_352_419# 1 2 9 15 19 21 25 30 31 33 37
+ 41 42 46 49
r106 42 50 32.0725 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.632 $Y=1.77
+ $X2=3.632 $Y2=1.935
r107 42 49 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.632 $Y=1.77
+ $X2=3.632 $Y2=1.605
r108 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.625
+ $Y=1.77 $X2=3.625 $Y2=1.77
r109 38 41 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=3.515 $Y=1.805
+ $X2=3.625 $Y2=1.805
r110 36 38 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.515 $Y=1.935
+ $X2=3.515 $Y2=1.805
r111 36 37 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.515 $Y=1.935
+ $X2=3.515 $Y2=2.075
r112 34 46 19.0514 $w=2.53e-07 $l=1e-07 $layer=POLY_cond $X=3.465 $Y=0.98
+ $X2=3.565 $Y2=0.98
r113 34 44 7.62055 $w=2.53e-07 $l=4e-08 $layer=POLY_cond $X=3.465 $Y=0.98
+ $X2=3.425 $Y2=0.98
r114 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.465
+ $Y=0.98 $X2=3.465 $Y2=0.98
r115 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.77 $Y=0.98
+ $X2=3.465 $Y2=0.98
r116 30 31 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.685 $Y=0.815
+ $X2=2.77 $Y2=0.98
r117 29 30 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.685 $Y=0.535
+ $X2=2.685 $Y2=0.815
r118 25 37 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.43 $Y=2.205
+ $X2=3.515 $Y2=2.075
r119 25 27 52.7464 $w=2.58e-07 $l=1.19e-06 $layer=LI1_cond $X=3.43 $Y=2.205
+ $X2=2.24 $Y2=2.205
r120 21 29 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.6 $Y=0.4
+ $X2=2.685 $Y2=0.535
r121 21 23 27.744 $w=2.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.6 $Y=0.4 $X2=1.95
+ $Y2=0.4
r122 17 46 47.6285 $w=2.53e-07 $l=3.22102e-07 $layer=POLY_cond $X=3.815 $Y=0.815
+ $X2=3.565 $Y2=0.98
r123 17 19 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.815 $Y=0.815
+ $X2=3.815 $Y2=0.445
r124 15 50 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.68 $Y=2.595
+ $X2=3.68 $Y2=1.935
r125 11 46 14.9957 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.565 $Y=1.145
+ $X2=3.565 $Y2=0.98
r126 11 49 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.565 $Y=1.145
+ $X2=3.565 $Y2=1.605
r127 7 44 14.9957 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=0.815
+ $X2=3.425 $Y2=0.98
r128 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.425 $Y=0.815
+ $X2=3.425 $Y2=0.445
r129 2 27 600 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=1 $X=1.76
+ $Y=2.095 $X2=2.24 $Y2=2.245
r130 1 23 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.81
+ $Y=0.235 $X2=1.95 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%CLK 1 3 4 5 6 8 11 13 15 18 20 27
c52 18 0 2.16197e-19 $X=5.61 $Y=2.595
c53 11 0 3.29628e-19 $X=5.08 $Y=2.595
r54 25 27 39.576 $w=4.08e-07 $l=3.35e-07 $layer=POLY_cond $X=5.11 $Y=1.707
+ $X2=5.445 $Y2=1.707
r55 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.11
+ $Y=1.62 $X2=5.11 $Y2=1.62
r56 23 25 3.54412 $w=4.08e-07 $l=3e-08 $layer=POLY_cond $X=5.08 $Y=1.707
+ $X2=5.11 $Y2=1.707
r57 22 23 7.67892 $w=4.08e-07 $l=6.5e-08 $layer=POLY_cond $X=5.015 $Y=1.707
+ $X2=5.08 $Y2=1.707
r58 20 26 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.52 $Y=1.62
+ $X2=5.11 $Y2=1.62
r59 16 27 19.4926 $w=4.08e-07 $l=3.25198e-07 $layer=POLY_cond $X=5.61 $Y=1.96
+ $X2=5.445 $Y2=1.707
r60 16 18 157.768 $w=2.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.61 $Y=1.96
+ $X2=5.61 $Y2=2.595
r61 13 27 26.3468 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=5.445 $Y=1.455
+ $X2=5.445 $Y2=1.707
r62 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.445 $Y=1.455
+ $X2=5.445 $Y2=1.135
r63 9 23 14.2339 $w=2.5e-07 $l=2.53e-07 $layer=POLY_cond $X=5.08 $Y=1.96
+ $X2=5.08 $Y2=1.707
r64 9 11 157.768 $w=2.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.08 $Y=1.96
+ $X2=5.08 $Y2=2.595
r65 6 22 26.3468 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=5.015 $Y=1.455
+ $X2=5.015 $Y2=1.707
r66 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.015 $Y=1.455
+ $X2=5.015 $Y2=1.135
r67 4 22 29.1132 $w=4.08e-07 $l=2.11197e-07 $layer=POLY_cond $X=4.94 $Y=1.53
+ $X2=5.015 $Y2=1.707
r68 4 5 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=4.94 $Y=1.53
+ $X2=4.615 $Y2=1.53
r69 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.54 $Y=1.455
+ $X2=4.615 $Y2=1.53
r70 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.54 $Y=1.455 $X2=4.54
+ $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%A_1147_419# 1 2 9 13 17 23 26 29 31 33 34
+ 36 38 39 46 47
c70 38 0 3.7271e-19 $X=5.875 $Y=2.48
c71 31 0 2.81132e-20 $X=6.485 $Y=0.99
c72 26 0 1.04487e-19 $X=6.65 $Y=1.575
c73 23 0 1.60623e-19 $X=6.705 $Y=0.98
r74 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.65
+ $Y=1.07 $X2=6.65 $Y2=1.07
r75 39 42 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=6.05 $Y=0.99
+ $X2=6.05 $Y2=1.135
r76 36 47 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.57 $Y=2.315
+ $X2=6.57 $Y2=1.575
r77 34 47 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=6.622 $Y=1.438
+ $X2=6.622 $Y2=1.575
r78 33 45 2.80348 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=6.622 $Y=1.075
+ $X2=6.622 $Y2=0.99
r79 33 34 15.2122 $w=2.73e-07 $l=3.63e-07 $layer=LI1_cond $X=6.622 $Y=1.075
+ $X2=6.622 $Y2=1.438
r80 32 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.215 $Y=0.99
+ $X2=6.05 $Y2=0.99
r81 31 45 4.51856 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=6.485 $Y=0.99
+ $X2=6.622 $Y2=0.99
r82 31 32 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.485 $Y=0.99
+ $X2=6.215 $Y2=0.99
r83 30 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.04 $Y=2.4
+ $X2=5.875 $Y2=2.4
r84 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.485 $Y=2.4
+ $X2=6.57 $Y2=2.315
r85 29 30 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.485 $Y=2.4
+ $X2=6.04 $Y2=2.4
r86 25 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.65 $Y=1.41
+ $X2=6.65 $Y2=1.07
r87 25 26 31.2043 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.65 $Y=1.41
+ $X2=6.65 $Y2=1.575
r88 22 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.65 $Y=1.055
+ $X2=6.65 $Y2=1.07
r89 22 23 28.2021 $w=1.5e-07 $l=5.5e-08 $layer=POLY_cond $X=6.65 $Y=0.98
+ $X2=6.705 $Y2=0.98
r90 19 22 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=6.345 $Y=0.98
+ $X2=6.65 $Y2=0.98
r91 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.705 $Y=0.905
+ $X2=6.705 $Y2=0.98
r92 15 17 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=6.705 $Y=0.905
+ $X2=6.705 $Y2=0.445
r93 13 26 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=6.67 $Y=2.595
+ $X2=6.67 $Y2=1.575
r94 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.345 $Y=0.905
+ $X2=6.345 $Y2=0.98
r95 7 9 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=6.345 $Y=0.905
+ $X2=6.345 $Y2=0.445
r96 2 38 300 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=2 $X=5.735
+ $Y=2.095 $X2=5.875 $Y2=2.48
r97 1 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.91
+ $Y=0.925 $X2=6.05 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%VPWR 1 2 3 4 17 21 25 29 32 33 35 36 37 52
+ 58 59 62 65
r82 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r83 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r84 59 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r85 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r86 56 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.57 $Y=3.33
+ $X2=6.405 $Y2=3.33
r87 56 58 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.57 $Y=3.33
+ $X2=6.96 $Y2=3.33
r88 55 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r89 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r90 52 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.24 $Y=3.33
+ $X2=6.405 $Y2=3.33
r91 52 54 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.24 $Y=3.33 $X2=6
+ $Y2=3.33
r92 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r93 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r94 47 50 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r96 42 45 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r97 42 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 41 44 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r99 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r100 39 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.84 $Y2=3.33
r101 39 41 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.2 $Y2=3.33
r102 37 51 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r103 37 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r104 37 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 35 50 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.18 $Y=3.33
+ $X2=5.345 $Y2=3.33
r107 34 54 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.51 $Y=3.33 $X2=6
+ $Y2=3.33
r108 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=3.33
+ $X2=5.345 $Y2=3.33
r109 32 44 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.18 $Y=3.33 $X2=3.12
+ $Y2=3.33
r110 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=3.33
+ $X2=3.345 $Y2=3.33
r111 31 47 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.51 $Y=3.33 $X2=3.6
+ $Y2=3.33
r112 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.51 $Y=3.33
+ $X2=3.345 $Y2=3.33
r113 27 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=3.245
+ $X2=6.405 $Y2=3.33
r114 27 29 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=6.405 $Y=3.245
+ $X2=6.405 $Y2=2.89
r115 23 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=3.245
+ $X2=5.345 $Y2=3.33
r116 23 25 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=5.345 $Y=3.245
+ $X2=5.345 $Y2=2.48
r117 19 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=3.245
+ $X2=3.345 $Y2=3.33
r118 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.345 $Y=3.245
+ $X2=3.345 $Y2=2.95
r119 15 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=3.245
+ $X2=0.84 $Y2=3.33
r120 15 17 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.84 $Y=3.245
+ $X2=0.84 $Y2=2.495
r121 4 29 600 $w=1.7e-07 $l=8.62163e-07 $layer=licon1_PDIFF $count=1 $X=6.265
+ $Y=2.095 $X2=6.405 $Y2=2.89
r122 3 25 300 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=2 $X=5.205
+ $Y=2.095 $X2=5.345 $Y2=2.48
r123 2 21 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=2.095 $X2=3.345 $Y2=2.95
r124 1 17 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=0.7
+ $Y=2.095 $X2=0.84 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%GCLK 1 2 10 13 14 15 30 32
r22 20 32 0.739303 $w=2.63e-07 $l=1.7e-08 $layer=LI1_cond $X=6.977 $Y=2.052
+ $X2=6.977 $Y2=2.035
r23 14 15 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=6.977 $Y=2.405
+ $X2=6.977 $Y2=2.775
r24 14 23 7.17559 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=6.977 $Y=2.405
+ $X2=6.977 $Y2=2.24
r25 13 32 1.47861 $w=2.63e-07 $l=3.4e-08 $layer=LI1_cond $X=6.977 $Y=2.001
+ $X2=6.977 $Y2=2.035
r26 13 30 4.99921 $w=2.63e-07 $l=8.1e-08 $layer=LI1_cond $X=6.977 $Y=2.001
+ $X2=6.977 $Y2=1.92
r27 13 23 6.69722 $w=2.63e-07 $l=1.54e-07 $layer=LI1_cond $X=6.977 $Y=2.086
+ $X2=6.977 $Y2=2.24
r28 13 20 1.47861 $w=2.63e-07 $l=3.4e-08 $layer=LI1_cond $X=6.977 $Y=2.086
+ $X2=6.977 $Y2=2.052
r29 12 30 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=7.025 $Y=0.675
+ $X2=7.025 $Y2=1.92
r30 10 12 9.79758 $w=3.53e-07 $l=2.05e-07 $layer=LI1_cond $X=6.932 $Y=0.47
+ $X2=6.932 $Y2=0.675
r31 2 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.795
+ $Y=2.095 $X2=6.935 $Y2=2.24
r32 1 10 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=6.78
+ $Y=0.235 $X2=6.92 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLCLKP_LP%VGND 1 2 3 4 15 17 21 25 27 31 33 34 35 37
+ 51 52 55 58 61
c87 17 0 1.88697e-19 $X=3.045 $Y=0
r88 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r89 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r90 56 59 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r91 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 52 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6
+ $Y2=0
r93 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r94 49 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.13
+ $Y2=0
r95 49 51 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.96
+ $Y2=0
r96 48 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r97 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r98 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r99 42 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.21
+ $Y2=0
r100 42 44 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.6
+ $Y2=0
r101 40 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r102 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r103 37 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.05
+ $Y2=0
r104 37 39 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0
+ $X2=0.72 $Y2=0
r105 35 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r106 35 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r107 35 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r108 33 47 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.065 $Y=0 $X2=5.04
+ $Y2=0
r109 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=0 $X2=5.23
+ $Y2=0
r110 29 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0
r111 29 31 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0.445
r112 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.23
+ $Y2=0
r113 27 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.965 $Y=0 $X2=6.13
+ $Y2=0
r114 27 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.965 $Y=0
+ $X2=5.395 $Y2=0
r115 23 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.23 $Y=0.085
+ $X2=5.23 $Y2=0
r116 23 25 35.0971 $w=3.28e-07 $l=1.005e-06 $layer=LI1_cond $X=5.23 $Y=0.085
+ $X2=5.23 $Y2=1.09
r117 19 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r118 19 21 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.425
r119 18 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=0 $X2=1.05
+ $Y2=0
r120 17 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.21
+ $Y2=0
r121 17 18 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=3.045 $Y=0
+ $X2=1.215 $Y2=0
r122 13 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.05 $Y=0.085
+ $X2=1.05 $Y2=0
r123 13 15 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.05 $Y=0.085
+ $X2=1.05 $Y2=0.415
r124 4 31 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.985
+ $Y=0.235 $X2=6.13 $Y2=0.445
r125 3 25 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.09
+ $Y=0.925 $X2=5.23 $Y2=1.09
r126 2 21 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.235 $X2=3.21 $Y2=0.425
r127 1 15 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.05 $Y2=0.415
.ends

