* File: sky130_fd_sc_lp__o2bb2a_m.pxi.spice
* Created: Fri Aug 28 11:12:17 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2A_M%A_85_187# N_A_85_187#_M1003_s N_A_85_187#_M1000_d
+ N_A_85_187#_M1001_g N_A_85_187#_M1006_g N_A_85_187#_c_82_n N_A_85_187#_c_83_n
+ N_A_85_187#_c_84_n N_A_85_187#_c_85_n N_A_85_187#_c_86_n N_A_85_187#_c_91_n
+ N_A_85_187#_c_87_n N_A_85_187#_c_92_n N_A_85_187#_c_88_n N_A_85_187#_c_94_n
+ PM_SKY130_FD_SC_LP__O2BB2A_M%A_85_187#
x_PM_SKY130_FD_SC_LP__O2BB2A_M%A1_N N_A1_N_M1011_g N_A1_N_M1007_g N_A1_N_c_156_n
+ N_A1_N_c_157_n A1_N A1_N N_A1_N_c_158_n N_A1_N_c_159_n
+ PM_SKY130_FD_SC_LP__O2BB2A_M%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2A_M%A2_N N_A2_N_M1008_g N_A2_N_M1002_g N_A2_N_c_200_n
+ N_A2_N_c_201_n A2_N A2_N A2_N N_A2_N_c_203_n PM_SKY130_FD_SC_LP__O2BB2A_M%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2A_M%A_209_535# N_A_209_535#_M1008_d
+ N_A_209_535#_M1011_d N_A_209_535#_c_244_n N_A_209_535#_M1000_g
+ N_A_209_535#_M1003_g N_A_209_535#_c_247_n N_A_209_535#_c_248_n
+ N_A_209_535#_c_249_n N_A_209_535#_c_263_n N_A_209_535#_c_242_n
+ N_A_209_535#_c_243_n N_A_209_535#_c_250_n
+ PM_SKY130_FD_SC_LP__O2BB2A_M%A_209_535#
x_PM_SKY130_FD_SC_LP__O2BB2A_M%B2 N_B2_M1009_g N_B2_M1004_g N_B2_c_316_n
+ N_B2_c_317_n B2 B2 B2 N_B2_c_314_n PM_SKY130_FD_SC_LP__O2BB2A_M%B2
x_PM_SKY130_FD_SC_LP__O2BB2A_M%B1 N_B1_c_355_n N_B1_M1010_g N_B1_M1005_g
+ N_B1_c_357_n B1 B1 B1 N_B1_c_359_n PM_SKY130_FD_SC_LP__O2BB2A_M%B1
x_PM_SKY130_FD_SC_LP__O2BB2A_M%X N_X_M1006_s N_X_M1001_s N_X_c_386_n X X X X X X
+ N_X_c_385_n PM_SKY130_FD_SC_LP__O2BB2A_M%X
x_PM_SKY130_FD_SC_LP__O2BB2A_M%VPWR N_VPWR_M1001_d N_VPWR_M1002_d N_VPWR_M1010_d
+ N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n
+ N_VPWR_c_409_n N_VPWR_c_410_n VPWR N_VPWR_c_411_n N_VPWR_c_412_n
+ N_VPWR_c_403_n N_VPWR_c_414_n PM_SKY130_FD_SC_LP__O2BB2A_M%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2A_M%VGND N_VGND_M1006_d N_VGND_M1004_d N_VGND_c_458_n
+ N_VGND_c_459_n N_VGND_c_460_n N_VGND_c_461_n VGND N_VGND_c_462_n
+ N_VGND_c_463_n N_VGND_c_464_n PM_SKY130_FD_SC_LP__O2BB2A_M%VGND
x_PM_SKY130_FD_SC_LP__O2BB2A_M%A_487_167# N_A_487_167#_M1003_d
+ N_A_487_167#_M1005_d N_A_487_167#_c_501_n N_A_487_167#_c_498_n
+ N_A_487_167#_c_499_n PM_SKY130_FD_SC_LP__O2BB2A_M%A_487_167#
cc_1 VNB N_A_85_187#_M1001_g 0.00268362f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.885
cc_2 VNB N_A_85_187#_M1006_g 0.0294748f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.445
cc_3 VNB N_A_85_187#_c_82_n 0.0253766f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.44
cc_4 VNB N_A_85_187#_c_83_n 0.0173144f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.605
cc_5 VNB N_A_85_187#_c_84_n 0.0011811f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.1
cc_6 VNB N_A_85_187#_c_85_n 0.0186596f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.1
cc_7 VNB N_A_85_187#_c_86_n 0.0246327f $X=-0.19 $Y=-0.245 $X2=2.04 $Y2=1.66
cc_8 VNB N_A_85_187#_c_87_n 0.00769594f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=1.11
cc_9 VNB N_A_85_187#_c_88_n 0.00161779f $X=-0.19 $Y=-0.245 $X2=2.207 $Y2=1.66
cc_10 VNB N_A1_N_M1007_g 0.0589478f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.605
cc_11 VNB N_A2_N_M1008_g 0.0202563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_N_M1002_g 0.0113859f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.605
cc_13 VNB N_A2_N_c_200_n 0.0254027f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.935
cc_14 VNB N_A2_N_c_201_n 0.0174745f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.445
cc_15 VNB A2_N 0.0116135f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.445
cc_16 VNB N_A2_N_c_203_n 0.0176203f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.1
cc_17 VNB N_A_209_535#_M1003_g 0.0398019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_209_535#_c_242_n 0.0106337f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=1.11
cc_19 VNB N_A_209_535#_c_243_n 0.0434107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B2_M1004_g 0.0236355f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.605
cc_21 VNB B2 0.00131438f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.445
cc_22 VNB N_B2_c_314_n 0.0146571f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.1
cc_23 VNB N_B1_M1005_g 0.0433033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB B1 0.00947924f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.1
cc_25 VNB X 0.0465526f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.445
cc_26 VNB N_X_c_385_n 0.0196285f $X=-0.19 $Y=-0.245 $X2=2.505 $Y2=2.835
cc_27 VNB N_VPWR_c_403_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_458_n 0.00494119f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.935
cc_29 VNB N_VGND_c_459_n 0.0320711f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.1
cc_30 VNB N_VGND_c_460_n 0.0526927f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.605
cc_31 VNB N_VGND_c_461_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.575
cc_32 VNB N_VGND_c_462_n 0.0228276f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.745
cc_33 VNB N_VGND_c_463_n 0.247045f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=2.67
cc_34 VNB N_VGND_c_464_n 0.026361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_487_167#_c_498_n 0.0159138f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.935
cc_36 VNB N_A_487_167#_c_499_n 0.00557763f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.445
cc_37 VPB N_A_85_187#_M1001_g 0.0694802f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.885
cc_38 VPB N_A_85_187#_c_86_n 0.0158665f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=1.66
cc_39 VPB N_A_85_187#_c_91_n 0.0028571f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.66
cc_40 VPB N_A_85_187#_c_92_n 0.0138268f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=2.67
cc_41 VPB N_A_85_187#_c_88_n 0.00182796f $X=-0.19 $Y=1.655 $X2=2.207 $Y2=1.66
cc_42 VPB N_A_85_187#_c_94_n 0.00604385f $X=-0.19 $Y=1.655 $X2=2.505 $Y2=2.835
cc_43 VPB N_A1_N_M1011_g 0.0194631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A1_N_M1007_g 0.00939624f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.605
cc_45 VPB N_A1_N_c_156_n 0.0209194f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.935
cc_46 VPB N_A1_N_c_157_n 0.0159361f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.445
cc_47 VPB N_A1_N_c_158_n 0.0152753f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.605
cc_48 VPB N_A1_N_c_159_n 0.00691937f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.575
cc_49 VPB N_A2_N_M1002_g 0.0674346f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.605
cc_50 VPB N_A_209_535#_c_244_n 0.103714f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.605
cc_51 VPB N_A_209_535#_M1000_g 0.0223459f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.885
cc_52 VPB N_A_209_535#_M1003_g 0.0114521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_209_535#_c_247_n 0.0061914f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.935
cc_54 VPB N_A_209_535#_c_248_n 0.00874553f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.44
cc_55 VPB N_A_209_535#_c_249_n 5.86919e-19 $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.605
cc_56 VPB N_A_209_535#_c_250_n 0.00814623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_B2_M1009_g 0.0340578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_B2_c_316_n 0.0209311f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.935
cc_59 VPB N_B2_c_317_n 0.0158337f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.445
cc_60 VPB B2 0.012376f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.445
cc_61 VPB N_B2_c_314_n 6.18422e-19 $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.1
cc_62 VPB N_B1_c_355_n 0.021073f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=0.835
cc_63 VPB N_B1_M1005_g 0.00267497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_B1_c_357_n 0.0813784f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.935
cc_65 VPB B1 0.0363852f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.1
cc_66 VPB N_B1_c_359_n 0.018372f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.1
cc_67 VPB N_X_c_386_n 0.0145804f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.885
cc_68 VPB X 0.0482713f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.445
cc_69 VPB N_VPWR_c_404_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.445
cc_70 VPB N_VPWR_c_405_n 0.00564356f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.935
cc_71 VPB N_VPWR_c_406_n 0.0125984f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.1
cc_72 VPB N_VPWR_c_407_n 0.0206563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_408_n 0.00631563f $X=-0.19 $Y=1.655 $X2=2.04 $Y2=1.66
cc_74 VPB N_VPWR_c_409_n 0.0307644f $X=-0.19 $Y=1.655 $X2=2.145 $Y2=1.575
cc_75 VPB N_VPWR_c_410_n 0.00510247f $X=-0.19 $Y=1.655 $X2=2.145 $Y2=1.11
cc_76 VPB N_VPWR_c_411_n 0.0173969f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.745
cc_77 VPB N_VPWR_c_412_n 0.0142356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_403_n 0.0519618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_414_n 0.00436274f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 N_A_85_187#_M1001_g N_A1_N_M1011_g 0.0142543f $X=0.5 $Y=2.885 $X2=0 $Y2=0
cc_81 N_A_85_187#_M1001_g N_A1_N_M1007_g 0.00733167f $X=0.5 $Y=2.885 $X2=0 $Y2=0
cc_82 N_A_85_187#_M1006_g N_A1_N_M1007_g 0.0217355f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A_85_187#_c_84_n N_A1_N_M1007_g 0.00240837f $X=0.59 $Y=1.1 $X2=0 $Y2=0
cc_84 N_A_85_187#_c_85_n N_A1_N_M1007_g 0.0412566f $X=0.59 $Y=1.1 $X2=0 $Y2=0
cc_85 N_A_85_187#_c_86_n N_A1_N_M1007_g 0.0149569f $X=2.04 $Y=1.66 $X2=0 $Y2=0
cc_86 N_A_85_187#_M1001_g N_A1_N_c_158_n 0.0399204f $X=0.5 $Y=2.885 $X2=0 $Y2=0
cc_87 N_A_85_187#_c_86_n N_A1_N_c_158_n 0.00512433f $X=2.04 $Y=1.66 $X2=0 $Y2=0
cc_88 N_A_85_187#_M1001_g N_A1_N_c_159_n 0.00518856f $X=0.5 $Y=2.885 $X2=0 $Y2=0
cc_89 N_A_85_187#_c_83_n N_A1_N_c_159_n 6.67744e-19 $X=0.59 $Y=1.605 $X2=0 $Y2=0
cc_90 N_A_85_187#_c_86_n N_A1_N_c_159_n 0.0329913f $X=2.04 $Y=1.66 $X2=0 $Y2=0
cc_91 N_A_85_187#_c_91_n N_A1_N_c_159_n 0.00345972f $X=0.675 $Y=1.66 $X2=0 $Y2=0
cc_92 N_A_85_187#_c_86_n N_A2_N_M1002_g 0.0142937f $X=2.04 $Y=1.66 $X2=0 $Y2=0
cc_93 N_A_85_187#_c_87_n N_A2_N_M1002_g 0.00265175f $X=2.145 $Y=1.11 $X2=0 $Y2=0
cc_94 N_A_85_187#_c_86_n N_A2_N_c_201_n 0.00505609f $X=2.04 $Y=1.66 $X2=0 $Y2=0
cc_95 N_A_85_187#_c_84_n A2_N 0.017234f $X=0.59 $Y=1.1 $X2=0 $Y2=0
cc_96 N_A_85_187#_c_86_n A2_N 0.0391406f $X=2.04 $Y=1.66 $X2=0 $Y2=0
cc_97 N_A_85_187#_c_87_n A2_N 0.0182034f $X=2.145 $Y=1.11 $X2=0 $Y2=0
cc_98 N_A_85_187#_c_87_n N_A2_N_c_203_n 0.00533743f $X=2.145 $Y=1.11 $X2=0 $Y2=0
cc_99 N_A_85_187#_c_86_n N_A_209_535#_c_244_n 0.010019f $X=2.04 $Y=1.66 $X2=0
+ $Y2=0
cc_100 N_A_85_187#_c_92_n N_A_209_535#_c_244_n 0.0287746f $X=2.29 $Y=2.67 $X2=0
+ $Y2=0
cc_101 N_A_85_187#_c_88_n N_A_209_535#_c_244_n 0.00854459f $X=2.207 $Y=1.66
+ $X2=0 $Y2=0
cc_102 N_A_85_187#_c_94_n N_A_209_535#_c_244_n 0.00166951f $X=2.505 $Y=2.835
+ $X2=0 $Y2=0
cc_103 N_A_85_187#_c_92_n N_A_209_535#_M1000_g 0.00573231f $X=2.29 $Y=2.67 $X2=0
+ $Y2=0
cc_104 N_A_85_187#_c_94_n N_A_209_535#_M1000_g 0.0113967f $X=2.505 $Y=2.835
+ $X2=0 $Y2=0
cc_105 N_A_85_187#_c_87_n N_A_209_535#_M1003_g 0.00830652f $X=2.145 $Y=1.11
+ $X2=0 $Y2=0
cc_106 N_A_85_187#_c_92_n N_A_209_535#_M1003_g 0.00297932f $X=2.29 $Y=2.67 $X2=0
+ $Y2=0
cc_107 N_A_85_187#_c_88_n N_A_209_535#_M1003_g 0.0113118f $X=2.207 $Y=1.66 $X2=0
+ $Y2=0
cc_108 N_A_85_187#_c_86_n N_A_209_535#_c_248_n 0.00621544f $X=2.04 $Y=1.66 $X2=0
+ $Y2=0
cc_109 N_A_85_187#_c_92_n N_A_209_535#_c_248_n 0.0123662f $X=2.29 $Y=2.67 $X2=0
+ $Y2=0
cc_110 N_A_85_187#_c_86_n N_A_209_535#_c_249_n 0.00528397f $X=2.04 $Y=1.66 $X2=0
+ $Y2=0
cc_111 N_A_85_187#_c_86_n N_A_209_535#_c_263_n 0.0245291f $X=2.04 $Y=1.66 $X2=0
+ $Y2=0
cc_112 N_A_85_187#_c_92_n N_A_209_535#_c_263_n 0.0231566f $X=2.29 $Y=2.67 $X2=0
+ $Y2=0
cc_113 N_A_85_187#_c_87_n N_A_209_535#_c_242_n 0.0100893f $X=2.145 $Y=1.11 $X2=0
+ $Y2=0
cc_114 N_A_85_187#_c_87_n N_A_209_535#_c_243_n 0.00147028f $X=2.145 $Y=1.11
+ $X2=0 $Y2=0
cc_115 N_A_85_187#_c_92_n N_B2_M1009_g 0.00330074f $X=2.29 $Y=2.67 $X2=0 $Y2=0
cc_116 N_A_85_187#_c_92_n N_B2_c_316_n 0.00151353f $X=2.29 $Y=2.67 $X2=0 $Y2=0
cc_117 N_A_85_187#_c_92_n B2 0.0568091f $X=2.29 $Y=2.67 $X2=0 $Y2=0
cc_118 N_A_85_187#_c_88_n B2 0.0135033f $X=2.207 $Y=1.66 $X2=0 $Y2=0
cc_119 N_A_85_187#_c_94_n B2 0.00444698f $X=2.505 $Y=2.835 $X2=0 $Y2=0
cc_120 N_A_85_187#_M1001_g N_X_c_386_n 8.03018e-19 $X=0.5 $Y=2.885 $X2=0 $Y2=0
cc_121 N_A_85_187#_M1006_g X 0.00849345f $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_85_187#_c_84_n X 0.0437496f $X=0.59 $Y=1.1 $X2=0 $Y2=0
cc_123 N_A_85_187#_c_85_n X 0.0447458f $X=0.59 $Y=1.1 $X2=0 $Y2=0
cc_124 N_A_85_187#_c_91_n X 0.0129659f $X=0.675 $Y=1.66 $X2=0 $Y2=0
cc_125 N_A_85_187#_M1006_g N_X_c_385_n 5.84046e-19 $X=0.61 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_85_187#_c_85_n N_X_c_385_n 0.00298608f $X=0.59 $Y=1.1 $X2=0 $Y2=0
cc_127 N_A_85_187#_M1001_g N_VPWR_c_404_n 0.00998194f $X=0.5 $Y=2.885 $X2=0
+ $Y2=0
cc_128 N_A_85_187#_c_94_n N_VPWR_c_409_n 0.0160652f $X=2.505 $Y=2.835 $X2=0
+ $Y2=0
cc_129 N_A_85_187#_M1001_g N_VPWR_c_411_n 0.00564095f $X=0.5 $Y=2.885 $X2=0
+ $Y2=0
cc_130 N_A_85_187#_M1000_d N_VPWR_c_403_n 0.00253815f $X=2.365 $Y=2.675 $X2=0
+ $Y2=0
cc_131 N_A_85_187#_M1001_g N_VPWR_c_403_n 0.0106196f $X=0.5 $Y=2.885 $X2=0 $Y2=0
cc_132 N_A_85_187#_c_94_n N_VPWR_c_403_n 0.0140646f $X=2.505 $Y=2.835 $X2=0
+ $Y2=0
cc_133 N_A_85_187#_M1006_g N_VGND_c_458_n 0.00288714f $X=0.61 $Y=0.445 $X2=0
+ $Y2=0
cc_134 N_A_85_187#_c_85_n N_VGND_c_458_n 8.82489e-19 $X=0.59 $Y=1.1 $X2=0 $Y2=0
cc_135 N_A_85_187#_M1006_g N_VGND_c_463_n 0.0118413f $X=0.61 $Y=0.445 $X2=0
+ $Y2=0
cc_136 N_A_85_187#_M1006_g N_VGND_c_464_n 0.00585385f $X=0.61 $Y=0.445 $X2=0
+ $Y2=0
cc_137 N_A_85_187#_c_87_n N_A_487_167#_c_499_n 0.00992277f $X=2.145 $Y=1.11
+ $X2=0 $Y2=0
cc_138 N_A1_N_M1007_g N_A2_N_M1008_g 0.0369491f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A1_N_M1011_g N_A2_N_M1002_g 0.016497f $X=0.97 $Y=2.885 $X2=0 $Y2=0
cc_140 N_A1_N_c_159_n N_A2_N_M1002_g 0.00200973f $X=0.95 $Y=2.01 $X2=0 $Y2=0
cc_141 N_A1_N_c_156_n N_A2_N_c_200_n 0.0369491f $X=0.95 $Y=2.35 $X2=0 $Y2=0
cc_142 N_A1_N_c_157_n N_A2_N_c_201_n 0.0369491f $X=0.95 $Y=2.515 $X2=0 $Y2=0
cc_143 N_A1_N_M1007_g A2_N 0.0147716f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A1_N_c_158_n N_A2_N_c_203_n 0.0369491f $X=0.95 $Y=2.01 $X2=0 $Y2=0
cc_145 N_A1_N_M1011_g N_A_209_535#_c_247_n 9.36826e-19 $X=0.97 $Y=2.885 $X2=0
+ $Y2=0
cc_146 N_A1_N_c_157_n N_A_209_535#_c_247_n 3.57326e-19 $X=0.95 $Y=2.515 $X2=0
+ $Y2=0
cc_147 N_A1_N_c_159_n N_A_209_535#_c_247_n 0.00315367f $X=0.95 $Y=2.01 $X2=0
+ $Y2=0
cc_148 N_A1_N_c_156_n N_A_209_535#_c_249_n 5.70835e-19 $X=0.95 $Y=2.35 $X2=0
+ $Y2=0
cc_149 N_A1_N_c_159_n N_A_209_535#_c_249_n 0.0109094f $X=0.95 $Y=2.01 $X2=0
+ $Y2=0
cc_150 N_A1_N_c_159_n N_A_209_535#_c_263_n 0.00949516f $X=0.95 $Y=2.01 $X2=0
+ $Y2=0
cc_151 N_A1_N_c_157_n N_A_209_535#_c_250_n 9.74091e-19 $X=0.95 $Y=2.515 $X2=0
+ $Y2=0
cc_152 N_A1_N_c_159_n N_A_209_535#_c_250_n 0.00261692f $X=0.95 $Y=2.01 $X2=0
+ $Y2=0
cc_153 N_A1_N_c_159_n X 0.0303615f $X=0.95 $Y=2.01 $X2=0 $Y2=0
cc_154 N_A1_N_M1011_g N_VPWR_c_404_n 0.00729534f $X=0.97 $Y=2.885 $X2=0 $Y2=0
cc_155 N_A1_N_c_157_n N_VPWR_c_404_n 0.00242751f $X=0.95 $Y=2.515 $X2=0 $Y2=0
cc_156 N_A1_N_c_159_n N_VPWR_c_404_n 0.0102988f $X=0.95 $Y=2.01 $X2=0 $Y2=0
cc_157 N_A1_N_M1011_g N_VPWR_c_407_n 0.00564095f $X=0.97 $Y=2.885 $X2=0 $Y2=0
cc_158 N_A1_N_M1011_g N_VPWR_c_403_n 0.00528686f $X=0.97 $Y=2.885 $X2=0 $Y2=0
cc_159 N_A1_N_c_157_n N_VPWR_c_403_n 9.08567e-19 $X=0.95 $Y=2.515 $X2=0 $Y2=0
cc_160 N_A1_N_c_159_n N_VPWR_c_403_n 0.00712958f $X=0.95 $Y=2.01 $X2=0 $Y2=0
cc_161 N_A1_N_M1007_g N_VGND_c_458_n 0.00288714f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A1_N_M1007_g N_VGND_c_460_n 0.00585385f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A1_N_M1007_g N_VGND_c_463_n 0.0105559f $X=1.04 $Y=0.445 $X2=0 $Y2=0
cc_164 A2_N N_A_209_535#_M1008_d 0.00411513f $X=1.115 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A2_N_M1002_g N_A_209_535#_c_244_n 0.0421555f $X=1.4 $Y=2.885 $X2=0
+ $Y2=0
cc_166 A2_N N_A_209_535#_M1003_g 0.00534072f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_167 N_A2_N_c_203_n N_A_209_535#_M1003_g 0.00745607f $X=1.49 $Y=0.955 $X2=0
+ $Y2=0
cc_168 N_A2_N_M1002_g N_A_209_535#_c_247_n 0.00879027f $X=1.4 $Y=2.885 $X2=0
+ $Y2=0
cc_169 N_A2_N_M1002_g N_A_209_535#_c_249_n 0.00811287f $X=1.4 $Y=2.885 $X2=0
+ $Y2=0
cc_170 N_A2_N_M1002_g N_A_209_535#_c_263_n 0.00132734f $X=1.4 $Y=2.885 $X2=0
+ $Y2=0
cc_171 N_A2_N_M1008_g N_A_209_535#_c_242_n 0.00509951f $X=1.4 $Y=0.445 $X2=0
+ $Y2=0
cc_172 A2_N N_A_209_535#_c_242_n 0.011276f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_173 N_A2_N_M1008_g N_A_209_535#_c_243_n 0.00323102f $X=1.4 $Y=0.445 $X2=0
+ $Y2=0
cc_174 A2_N N_A_209_535#_c_243_n 3.10683e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A2_N_M1002_g N_A_209_535#_c_250_n 0.012588f $X=1.4 $Y=2.885 $X2=0 $Y2=0
cc_176 A2_N N_X_c_385_n 6.61694e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_177 N_A2_N_M1002_g N_VPWR_c_404_n 0.00137831f $X=1.4 $Y=2.885 $X2=0 $Y2=0
cc_178 N_A2_N_M1002_g N_VPWR_c_405_n 0.00767552f $X=1.4 $Y=2.885 $X2=0 $Y2=0
cc_179 N_A2_N_M1002_g N_VPWR_c_407_n 0.00373071f $X=1.4 $Y=2.885 $X2=0 $Y2=0
cc_180 N_A2_N_M1002_g N_VPWR_c_403_n 0.0068865f $X=1.4 $Y=2.885 $X2=0 $Y2=0
cc_181 N_A2_N_M1008_g N_VGND_c_460_n 0.00398598f $X=1.4 $Y=0.445 $X2=0 $Y2=0
cc_182 A2_N N_VGND_c_460_n 0.0130493f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_183 N_A2_N_M1008_g N_VGND_c_463_n 0.00689053f $X=1.4 $Y=0.445 $X2=0 $Y2=0
cc_184 A2_N N_VGND_c_463_n 0.0176255f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_185 A2_N A_223_47# 0.00139886f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_186 N_A_209_535#_M1003_g N_B2_M1004_g 0.0200367f $X=2.36 $Y=1.045 $X2=0 $Y2=0
cc_187 N_A_209_535#_c_244_n N_B2_c_316_n 0.0351867f $X=2.29 $Y=2.515 $X2=0 $Y2=0
cc_188 N_A_209_535#_M1000_g N_B2_c_317_n 0.0198761f $X=2.29 $Y=2.885 $X2=0 $Y2=0
cc_189 N_A_209_535#_c_244_n B2 0.0017851f $X=2.29 $Y=2.515 $X2=0 $Y2=0
cc_190 N_A_209_535#_M1003_g B2 0.00266489f $X=2.36 $Y=1.045 $X2=0 $Y2=0
cc_191 N_A_209_535#_M1003_g N_B2_c_314_n 0.0153105f $X=2.36 $Y=1.045 $X2=0 $Y2=0
cc_192 N_A_209_535#_c_244_n N_VPWR_c_405_n 0.00812717f $X=2.29 $Y=2.515 $X2=0
+ $Y2=0
cc_193 N_A_209_535#_M1000_g N_VPWR_c_405_n 0.00805545f $X=2.29 $Y=2.885 $X2=0
+ $Y2=0
cc_194 N_A_209_535#_c_248_n N_VPWR_c_405_n 0.0139881f $X=1.695 $Y=2.35 $X2=0
+ $Y2=0
cc_195 N_A_209_535#_c_250_n N_VPWR_c_407_n 0.016805f $X=1.43 $Y=2.835 $X2=0
+ $Y2=0
cc_196 N_A_209_535#_M1000_g N_VPWR_c_409_n 0.00373071f $X=2.29 $Y=2.885 $X2=0
+ $Y2=0
cc_197 N_A_209_535#_M1011_d N_VPWR_c_403_n 0.00252989f $X=1.045 $Y=2.675 $X2=0
+ $Y2=0
cc_198 N_A_209_535#_c_244_n N_VPWR_c_403_n 0.00468299f $X=2.29 $Y=2.515 $X2=0
+ $Y2=0
cc_199 N_A_209_535#_M1000_g N_VPWR_c_403_n 0.0068865f $X=2.29 $Y=2.885 $X2=0
+ $Y2=0
cc_200 N_A_209_535#_c_250_n N_VPWR_c_403_n 0.01516f $X=1.43 $Y=2.835 $X2=0 $Y2=0
cc_201 N_A_209_535#_M1003_g N_VGND_c_459_n 0.00391431f $X=2.36 $Y=1.045 $X2=0
+ $Y2=0
cc_202 N_A_209_535#_c_242_n N_VGND_c_459_n 0.0134416f $X=2.34 $Y=0.44 $X2=0
+ $Y2=0
cc_203 N_A_209_535#_c_243_n N_VGND_c_459_n 0.00688791f $X=2.34 $Y=0.44 $X2=0
+ $Y2=0
cc_204 N_A_209_535#_c_242_n N_VGND_c_460_n 0.034353f $X=2.34 $Y=0.44 $X2=0 $Y2=0
cc_205 N_A_209_535#_c_243_n N_VGND_c_460_n 0.00861782f $X=2.34 $Y=0.44 $X2=0
+ $Y2=0
cc_206 N_A_209_535#_M1008_d N_VGND_c_463_n 0.0113943f $X=1.475 $Y=0.235 $X2=0
+ $Y2=0
cc_207 N_A_209_535#_c_242_n N_VGND_c_463_n 0.0221088f $X=2.34 $Y=0.44 $X2=0
+ $Y2=0
cc_208 N_A_209_535#_c_243_n N_VGND_c_463_n 0.0110351f $X=2.34 $Y=0.44 $X2=0
+ $Y2=0
cc_209 N_A_209_535#_c_243_n N_A_487_167#_c_501_n 8.10213e-19 $X=2.34 $Y=0.44
+ $X2=0 $Y2=0
cc_210 N_A_209_535#_M1003_g N_A_487_167#_c_499_n 0.00132343f $X=2.36 $Y=1.045
+ $X2=0 $Y2=0
cc_211 N_B2_M1004_g N_B1_M1005_g 0.018572f $X=2.79 $Y=1.045 $X2=0 $Y2=0
cc_212 B2 N_B1_M1005_g 0.00211534f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_213 N_B2_c_314_n N_B1_M1005_g 0.0138545f $X=2.81 $Y=1.665 $X2=0 $Y2=0
cc_214 N_B2_M1009_g N_B1_c_357_n 0.0579745f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_215 N_B2_c_317_n N_B1_c_357_n 0.0138545f $X=2.81 $Y=2.17 $X2=0 $Y2=0
cc_216 B2 N_B1_c_357_n 0.0029842f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_217 N_B2_M1009_g B1 3.67947e-19 $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_218 B2 B1 0.0475003f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_219 N_B2_c_314_n B1 0.00181479f $X=2.81 $Y=1.665 $X2=0 $Y2=0
cc_220 N_B2_c_316_n N_B1_c_359_n 0.0138545f $X=2.81 $Y=2.005 $X2=0 $Y2=0
cc_221 N_B2_M1009_g N_VPWR_c_406_n 0.00204602f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_222 N_B2_M1009_g N_VPWR_c_409_n 0.00585385f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_223 N_B2_M1009_g N_VPWR_c_403_n 0.00639038f $X=2.72 $Y=2.885 $X2=0 $Y2=0
cc_224 B2 N_VPWR_c_403_n 0.0133021f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B2_M1004_g N_VGND_c_459_n 0.00661257f $X=2.79 $Y=1.045 $X2=0 $Y2=0
cc_226 N_B2_M1004_g N_VGND_c_460_n 0.00308772f $X=2.79 $Y=1.045 $X2=0 $Y2=0
cc_227 N_B2_M1004_g N_VGND_c_463_n 0.00404023f $X=2.79 $Y=1.045 $X2=0 $Y2=0
cc_228 N_B2_M1004_g N_A_487_167#_c_498_n 0.0140204f $X=2.79 $Y=1.045 $X2=0 $Y2=0
cc_229 B2 N_A_487_167#_c_498_n 0.021428f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_230 N_B2_c_314_n N_A_487_167#_c_498_n 0.00411751f $X=2.81 $Y=1.665 $X2=0
+ $Y2=0
cc_231 B2 N_A_487_167#_c_499_n 0.0104508f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_232 N_B2_c_314_n N_A_487_167#_c_499_n 0.00102667f $X=2.81 $Y=1.665 $X2=0
+ $Y2=0
cc_233 N_B1_c_355_n N_VPWR_c_406_n 0.011235f $X=3.08 $Y=2.56 $X2=0 $Y2=0
cc_234 N_B1_c_357_n N_VPWR_c_406_n 0.00822039f $X=3.35 $Y=2.41 $X2=0 $Y2=0
cc_235 B1 N_VPWR_c_406_n 0.00898021f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_236 N_B1_c_355_n N_VPWR_c_409_n 0.00486043f $X=3.08 $Y=2.56 $X2=0 $Y2=0
cc_237 N_B1_c_357_n N_VPWR_c_412_n 0.00107984f $X=3.35 $Y=2.41 $X2=0 $Y2=0
cc_238 N_B1_c_355_n N_VPWR_c_403_n 0.00818711f $X=3.08 $Y=2.56 $X2=0 $Y2=0
cc_239 N_B1_c_357_n N_VPWR_c_403_n 0.00149216f $X=3.35 $Y=2.41 $X2=0 $Y2=0
cc_240 B1 N_VPWR_c_403_n 0.009764f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_241 N_B1_M1005_g N_VGND_c_459_n 0.0126541f $X=3.26 $Y=1.045 $X2=0 $Y2=0
cc_242 N_B1_M1005_g N_VGND_c_462_n 0.00308772f $X=3.26 $Y=1.045 $X2=0 $Y2=0
cc_243 N_B1_M1005_g N_VGND_c_463_n 0.00404023f $X=3.26 $Y=1.045 $X2=0 $Y2=0
cc_244 N_B1_M1005_g N_A_487_167#_c_498_n 0.017675f $X=3.26 $Y=1.045 $X2=0 $Y2=0
cc_245 B1 N_A_487_167#_c_498_n 0.0256306f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_246 N_B1_c_359_n N_A_487_167#_c_498_n 9.84594e-19 $X=3.35 $Y=1.865 $X2=0
+ $Y2=0
cc_247 N_X_c_386_n N_VPWR_c_411_n 0.00980051f $X=0.285 $Y=2.82 $X2=0 $Y2=0
cc_248 N_X_M1001_s N_VPWR_c_403_n 0.0034811f $X=0.16 $Y=2.675 $X2=0 $Y2=0
cc_249 N_X_c_386_n N_VPWR_c_403_n 0.00857705f $X=0.285 $Y=2.82 $X2=0 $Y2=0
cc_250 N_X_M1006_s N_VGND_c_463_n 0.0034811f $X=0.27 $Y=0.235 $X2=0 $Y2=0
cc_251 N_X_c_385_n N_VGND_c_463_n 0.0125588f $X=0.395 $Y=0.51 $X2=0 $Y2=0
cc_252 N_X_c_385_n N_VGND_c_464_n 0.0145747f $X=0.395 $Y=0.51 $X2=0 $Y2=0
cc_253 N_VPWR_c_403_n A_559_535# 0.00395178f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_254 N_VGND_c_463_n A_223_47# 0.00197491f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_255 N_VGND_M1004_d N_A_487_167#_c_498_n 0.00224299f $X=2.865 $Y=0.835 $X2=0
+ $Y2=0
cc_256 N_VGND_c_459_n N_A_487_167#_c_498_n 0.0165599f $X=3.025 $Y=0.96 $X2=0
+ $Y2=0
