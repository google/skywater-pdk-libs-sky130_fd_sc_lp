* File: sky130_fd_sc_lp__nand4b_m.spice
* Created: Fri Aug 28 10:52:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4b_m.pex.spice"
.subckt sky130_fd_sc_lp__nand4b_m  VNB VPB A_N D C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* D	D
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_N_M1003_g N_A_35_392#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.12285 AS=0.1113 PD=1.005 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1008 A_271_52# N_D_M1008_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.12285 PD=0.63 PS=1.005 NRD=14.28 NRS=87.132 M=1 R=2.8 SA=75000.9
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1009 A_343_52# N_C_M1009_g A_271_52# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75001.3 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1001 A_451_52# N_B_M1001_g A_343_52# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=39.996 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_A_35_392#_M1007_g A_451_52# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_N_M1005_g N_A_35_392#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1302 AS=0.1113 PD=1.04 PS=1.37 NRD=159.471 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_D_M1004_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1302 PD=0.7 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_C_M1000_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_B_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_35_392#_M1002_g N_Y_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__nand4b_m.pxi.spice"
*
.ends
*
*
