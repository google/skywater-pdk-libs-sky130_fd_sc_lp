# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__or4bb_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 1.210000 1.355000 1.755000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 1.345000 1.890000 1.755000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.365000 1.750000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.875000 0.955000 6.155000 1.750000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.465000 0.895000 5.225000 1.145000 ;
        RECT 3.790000 1.745000 5.225000 1.915000 ;
        RECT 3.790000 1.915000 3.980000 3.075000 ;
        RECT 4.650000 1.915000 4.840000 3.075000 ;
        RECT 4.890000 1.145000 5.225000 1.745000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.355000  0.730000 0.705000 1.040000 ;
      RECT 0.355000  1.920000 0.705000 1.925000 ;
      RECT 0.355000  1.925000 2.350000 2.095000 ;
      RECT 0.355000  2.095000 0.685000 2.210000 ;
      RECT 0.535000  1.040000 0.705000 1.920000 ;
      RECT 0.875000  0.085000 1.195000 1.040000 ;
      RECT 0.895000  2.265000 1.225000 3.245000 ;
      RECT 1.365000  0.255000 1.695000 0.995000 ;
      RECT 1.365000  0.995000 2.700000 1.040000 ;
      RECT 1.525000  1.040000 2.700000 1.165000 ;
      RECT 1.865000  0.085000 2.195000 0.815000 ;
      RECT 2.100000  1.345000 2.350000 1.925000 ;
      RECT 2.365000  0.255000 2.700000 0.995000 ;
      RECT 2.530000  1.165000 2.700000 1.755000 ;
      RECT 2.530000  1.755000 3.540000 1.925000 ;
      RECT 2.765000  1.925000 3.095000 3.075000 ;
      RECT 2.870000  0.555000 5.865000 0.715000 ;
      RECT 2.870000  0.715000 5.705000 0.725000 ;
      RECT 2.870000  0.725000 3.130000 1.545000 ;
      RECT 2.880000  0.085000 3.210000 0.385000 ;
      RECT 3.290000  2.095000 3.620000 3.245000 ;
      RECT 3.300000  1.325000 4.720000 1.575000 ;
      RECT 3.300000  1.575000 3.540000 1.755000 ;
      RECT 3.955000  0.085000 4.285000 0.385000 ;
      RECT 4.150000  2.085000 4.480000 3.245000 ;
      RECT 4.990000  0.085000 5.320000 0.385000 ;
      RECT 5.010000  2.085000 5.340000 3.245000 ;
      RECT 5.510000  0.725000 5.705000 1.920000 ;
      RECT 5.510000  1.920000 5.865000 2.210000 ;
      RECT 5.535000  0.310000 5.865000 0.555000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__or4bb_4
