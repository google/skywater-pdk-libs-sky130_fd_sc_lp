* File: sky130_fd_sc_lp__o2bb2a_2.spice
* Created: Fri Aug 28 11:11:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2a_2.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2a_2  VNB VPB B1 B2 A2_N A1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1_N	A1_N
* A2_N	A2_N
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_B1_M1004_g N_A_67_47#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_A_67_47#_M1003_d N_B2_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_222_367#_M1009_d N_A_300_21#_M1009_g N_A_67_47#_M1003_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 A_585_47# N_A2_N_M1011_g N_A_300_21#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A1_N_M1012_g A_585_47# VNB NSHORT L=0.15 W=0.42 AD=0.098
+ AS=0.0441 PD=0.85 PS=0.63 NRD=24.276 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_222_367#_M1002_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.196 PD=1.12 PS=1.7 NRD=0 NRS=4.992 M=1 R=5.6 SA=75000.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1006 N_X_M1002_d N_A_222_367#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 A_150_367# N_B1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.7 A=0.096 P=1.58 MULT=1
MM1010 N_A_222_367#_M1010_d N_B2_M1010_g A_150_367# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=16.9223 NRS=15.3857 M=1 R=4.26667
+ SA=75000.6 SB=75003.4 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A_300_21#_M1007_g N_A_222_367#_M1010_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2656 AS=0.1248 PD=1.47 PS=1.03 NRD=61.5625 NRS=16.9223 M=1
+ R=4.26667 SA=75001.1 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_300_21#_M1000_d N_A2_N_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2656 PD=0.92 PS=1.47 NRD=0 NRS=107.72 M=1 R=4.26667
+ SA=75002.1 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A1_N_M1008_g N_A_300_21#_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.197625 AS=0.0896 PD=1.29347 PS=0.92 NRD=240.084 NRS=0 M=1
+ R=4.26667 SA=75002.5 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1008_d N_A_222_367#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.389075 AS=0.1764 PD=2.54653 PS=1.54 NRD=2.0685 NRS=0 M=1 R=8.4 SA=75001.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A_222_367#_M1013_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
c_89 VPB 0 1.02291e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o2bb2a_2.pxi.spice"
*
.ends
*
*
