* File: sky130_fd_sc_lp__buf_m.pxi.spice
* Created: Fri Aug 28 10:10:50 2020
* 
x_PM_SKY130_FD_SC_LP__BUF_M%A_47_178# N_A_47_178#_M1002_d N_A_47_178#_M1001_d
+ N_A_47_178#_c_34_n N_A_47_178#_c_35_n N_A_47_178#_M1000_g N_A_47_178#_M1003_g
+ N_A_47_178#_c_36_n N_A_47_178#_c_41_n N_A_47_178#_c_42_n N_A_47_178#_c_43_n
+ N_A_47_178#_c_37_n N_A_47_178#_c_38_n N_A_47_178#_c_45_n
+ PM_SKY130_FD_SC_LP__BUF_M%A_47_178#
x_PM_SKY130_FD_SC_LP__BUF_M%A N_A_M1002_g N_A_c_95_n N_A_M1001_g N_A_c_92_n
+ N_A_c_97_n A A A N_A_c_94_n PM_SKY130_FD_SC_LP__BUF_M%A
x_PM_SKY130_FD_SC_LP__BUF_M%X N_X_M1000_s N_X_M1003_s X X X X X X N_X_c_137_n
+ PM_SKY130_FD_SC_LP__BUF_M%X
x_PM_SKY130_FD_SC_LP__BUF_M%VPWR N_VPWR_M1003_d N_VPWR_c_154_n N_VPWR_c_155_n
+ N_VPWR_c_156_n VPWR N_VPWR_c_157_n N_VPWR_c_153_n
+ PM_SKY130_FD_SC_LP__BUF_M%VPWR
x_PM_SKY130_FD_SC_LP__BUF_M%VGND N_VGND_M1000_d N_VGND_c_172_n N_VGND_c_173_n
+ N_VGND_c_174_n VGND N_VGND_c_175_n N_VGND_c_176_n
+ PM_SKY130_FD_SC_LP__BUF_M%VGND
cc_1 VNB N_A_47_178#_c_34_n 0.0399887f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.85
cc_2 VNB N_A_47_178#_c_35_n 0.0219614f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.89
cc_3 VNB N_A_47_178#_c_36_n 0.0267354f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.965
cc_4 VNB N_A_47_178#_c_37_n 0.0231648f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.93
cc_5 VNB N_A_47_178#_c_38_n 0.0026978f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.495
cc_6 VNB N_A_M1002_g 0.0422695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_c_92_n 0.00313241f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.89
cc_8 VNB A 0.00618114f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.86
cc_9 VNB N_A_c_94_n 0.072241f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=2.1
cc_10 VNB N_X_c_137_n 0.032181f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.015
cc_11 VNB N_VPWR_c_153_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_172_n 0.00798166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_173_n 0.0194501f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.89
cc_14 VNB N_VGND_c_174_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.56
cc_15 VNB N_VGND_c_175_n 0.0209787f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.965
cc_16 VNB N_VGND_c_176_n 0.123334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VPB N_A_47_178#_c_34_n 0.0139922f $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.85
cc_18 VPB N_A_47_178#_M1003_g 0.0418156f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.86
cc_19 VPB N_A_47_178#_c_41_n 0.00297844f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.015
cc_20 VPB N_A_47_178#_c_42_n 0.0707366f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.015
cc_21 VPB N_A_47_178#_c_43_n 0.00813905f $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.795
cc_22 VPB N_A_47_178#_c_37_n 0.00299073f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.93
cc_23 VPB N_A_47_178#_c_45_n 5.14497e-19 $X=-0.19 $Y=1.655 $X2=1.12 $Y2=2.015
cc_24 VPB N_A_c_95_n 0.0197663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 VPB N_A_c_92_n 0.0580438f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.89
cc_26 VPB N_A_c_97_n 0.0341167f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.18
cc_27 VPB A 0.00288691f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.86
cc_28 VPB N_X_c_137_n 0.0417274f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.015
cc_29 VPB N_VPWR_c_154_n 0.00567558f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_155_n 0.0191968f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.89
cc_31 VPB N_VPWR_c_156_n 0.0040126f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.56
cc_32 VPB N_VPWR_c_157_n 0.0211061f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.965
cc_33 VPB N_VPWR_c_153_n 0.0583098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 N_A_47_178#_c_34_n N_A_M1002_g 0.00506654f $X=0.31 $Y=1.85 $X2=0 $Y2=0
cc_35 N_A_47_178#_c_35_n N_A_M1002_g 0.0195183f $X=0.475 $Y=0.89 $X2=0 $Y2=0
cc_36 N_A_47_178#_c_37_n N_A_M1002_g 0.0157142f $X=1.14 $Y=1.93 $X2=0 $Y2=0
cc_37 N_A_47_178#_c_38_n N_A_M1002_g 4.64676e-19 $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_38 N_A_47_178#_c_43_n N_A_c_95_n 0.00316026f $X=1.12 $Y=2.795 $X2=0 $Y2=0
cc_39 N_A_47_178#_M1003_g N_A_c_92_n 0.00182353f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_40 N_A_47_178#_c_42_n N_A_c_92_n 0.018171f $X=0.71 $Y=2.015 $X2=0 $Y2=0
cc_41 N_A_47_178#_c_43_n N_A_c_92_n 0.0156198f $X=1.12 $Y=2.795 $X2=0 $Y2=0
cc_42 N_A_47_178#_c_37_n N_A_c_92_n 0.0176236f $X=1.14 $Y=1.93 $X2=0 $Y2=0
cc_43 N_A_47_178#_c_45_n N_A_c_92_n 0.0108117f $X=1.12 $Y=2.015 $X2=0 $Y2=0
cc_44 N_A_47_178#_M1003_g N_A_c_97_n 0.0209615f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_45 N_A_47_178#_c_41_n N_A_c_97_n 0.00516243f $X=1.015 $Y=2.015 $X2=0 $Y2=0
cc_46 N_A_47_178#_c_42_n N_A_c_97_n 0.00326016f $X=0.71 $Y=2.015 $X2=0 $Y2=0
cc_47 N_A_47_178#_c_43_n N_A_c_97_n 0.0182483f $X=1.12 $Y=2.795 $X2=0 $Y2=0
cc_48 N_A_47_178#_c_34_n A 0.00542815f $X=0.31 $Y=1.85 $X2=0 $Y2=0
cc_49 N_A_47_178#_c_35_n A 0.00175393f $X=0.475 $Y=0.89 $X2=0 $Y2=0
cc_50 N_A_47_178#_c_41_n A 0.0183938f $X=1.015 $Y=2.015 $X2=0 $Y2=0
cc_51 N_A_47_178#_c_42_n A 0.00183591f $X=0.71 $Y=2.015 $X2=0 $Y2=0
cc_52 N_A_47_178#_c_37_n A 0.0632293f $X=1.14 $Y=1.93 $X2=0 $Y2=0
cc_53 N_A_47_178#_c_34_n N_A_c_94_n 0.0171342f $X=0.31 $Y=1.85 $X2=0 $Y2=0
cc_54 N_A_47_178#_c_41_n N_A_c_94_n 0.00509287f $X=1.015 $Y=2.015 $X2=0 $Y2=0
cc_55 N_A_47_178#_c_42_n N_A_c_94_n 0.0131494f $X=0.71 $Y=2.015 $X2=0 $Y2=0
cc_56 N_A_47_178#_c_37_n N_A_c_94_n 0.0276054f $X=1.14 $Y=1.93 $X2=0 $Y2=0
cc_57 N_A_47_178#_c_38_n N_A_c_94_n 7.24074e-19 $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_58 N_A_47_178#_c_45_n N_A_c_94_n 0.00151481f $X=1.12 $Y=2.015 $X2=0 $Y2=0
cc_59 N_A_47_178#_c_34_n N_X_c_137_n 0.0315464f $X=0.31 $Y=1.85 $X2=0 $Y2=0
cc_60 N_A_47_178#_c_35_n N_X_c_137_n 0.00401643f $X=0.475 $Y=0.89 $X2=0 $Y2=0
cc_61 N_A_47_178#_M1003_g N_X_c_137_n 0.0135978f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_62 N_A_47_178#_c_36_n N_X_c_137_n 0.00875433f $X=0.475 $Y=0.965 $X2=0 $Y2=0
cc_63 N_A_47_178#_c_41_n N_X_c_137_n 0.0124012f $X=1.015 $Y=2.015 $X2=0 $Y2=0
cc_64 N_A_47_178#_c_42_n N_X_c_137_n 0.0203517f $X=0.71 $Y=2.015 $X2=0 $Y2=0
cc_65 N_A_47_178#_c_43_n N_X_c_137_n 0.0156484f $X=1.12 $Y=2.795 $X2=0 $Y2=0
cc_66 N_A_47_178#_M1003_g N_VPWR_c_154_n 0.00284446f $X=0.475 $Y=2.86 $X2=0
+ $Y2=0
cc_67 N_A_47_178#_c_41_n N_VPWR_c_154_n 0.0049357f $X=1.015 $Y=2.015 $X2=0 $Y2=0
cc_68 N_A_47_178#_c_42_n N_VPWR_c_154_n 0.00354513f $X=0.71 $Y=2.015 $X2=0 $Y2=0
cc_69 N_A_47_178#_M1003_g N_VPWR_c_155_n 0.00560159f $X=0.475 $Y=2.86 $X2=0
+ $Y2=0
cc_70 N_A_47_178#_c_43_n N_VPWR_c_157_n 0.00795263f $X=1.12 $Y=2.795 $X2=0 $Y2=0
cc_71 N_A_47_178#_M1003_g N_VPWR_c_153_n 0.0113779f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_72 N_A_47_178#_c_43_n N_VPWR_c_153_n 0.0075889f $X=1.12 $Y=2.795 $X2=0 $Y2=0
cc_73 N_A_47_178#_c_35_n N_VGND_c_172_n 0.00319474f $X=0.475 $Y=0.89 $X2=0 $Y2=0
cc_74 N_A_47_178#_c_38_n N_VGND_c_172_n 0.00123197f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_75 N_A_47_178#_c_35_n N_VGND_c_173_n 0.00478016f $X=0.475 $Y=0.89 $X2=0 $Y2=0
cc_76 N_A_47_178#_c_38_n N_VGND_c_175_n 0.00999378f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_77 N_A_47_178#_c_35_n N_VGND_c_176_n 0.00956748f $X=0.475 $Y=0.89 $X2=0 $Y2=0
cc_78 N_A_47_178#_c_38_n N_VGND_c_176_n 0.00774102f $X=1.12 $Y=0.495 $X2=0 $Y2=0
cc_79 N_A_M1002_g N_X_c_137_n 3.44994e-19 $X=0.905 $Y=0.56 $X2=0 $Y2=0
cc_80 A N_X_c_137_n 0.0469976f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_81 N_A_c_94_n N_X_c_137_n 0.00134568f $X=1.19 $Y=1.445 $X2=0 $Y2=0
cc_82 N_A_c_95_n N_VPWR_c_154_n 0.00284446f $X=0.905 $Y=2.54 $X2=0 $Y2=0
cc_83 N_A_c_95_n N_VPWR_c_157_n 0.00560159f $X=0.905 $Y=2.54 $X2=0 $Y2=0
cc_84 N_A_c_95_n N_VPWR_c_153_n 0.0114239f $X=0.905 $Y=2.54 $X2=0 $Y2=0
cc_85 N_A_c_97_n N_VPWR_c_153_n 0.00183521f $X=1.19 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A_M1002_g N_VGND_c_172_n 0.00286691f $X=0.905 $Y=0.56 $X2=0 $Y2=0
cc_87 A N_VGND_c_172_n 0.012617f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A_c_94_n N_VGND_c_172_n 7.97056e-19 $X=1.19 $Y=1.445 $X2=0 $Y2=0
cc_89 N_A_M1002_g N_VGND_c_175_n 0.00478016f $X=0.905 $Y=0.56 $X2=0 $Y2=0
cc_90 N_A_M1002_g N_VGND_c_176_n 0.00827221f $X=0.905 $Y=0.56 $X2=0 $Y2=0
cc_91 A N_VGND_c_176_n 0.00340668f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_92 N_X_c_137_n N_VPWR_c_155_n 0.00795263f $X=0.26 $Y=0.625 $X2=0 $Y2=0
cc_93 N_X_c_137_n N_VPWR_c_153_n 0.0075889f $X=0.26 $Y=0.625 $X2=0 $Y2=0
cc_94 N_X_c_137_n N_VGND_c_173_n 0.00590349f $X=0.26 $Y=0.625 $X2=0 $Y2=0
cc_95 N_X_c_137_n N_VGND_c_176_n 0.00715453f $X=0.26 $Y=0.625 $X2=0 $Y2=0
