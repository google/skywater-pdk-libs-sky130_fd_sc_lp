* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfxtp_lp CLK D VGND VNB VPB VPWR Q
X0 a_629_125# a_263_409# a_747_79# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_270_57# a_27_57# a_263_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR a_1429_383# a_1583_285# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_1626_75# a_1583_285# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_1429_383# a_1784_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_747_79# a_1355_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_27_57# a_263_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_902_125# a_1005_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_1583_285# a_2054_92# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_112_57# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_27_57# CLK a_112_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND a_27_57# a_270_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_2054_92# a_1583_285# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR D a_629_125# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VPWR a_747_79# a_1005_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_27_57# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_1429_383# a_263_409# a_1535_383# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_1005_99# a_263_409# a_1429_383# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1429_383# a_27_57# a_1626_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_747_79# a_263_409# a_902_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1355_125# a_747_79# a_1005_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1535_383# a_1583_285# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_1005_99# a_27_57# a_1429_383# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X23 VGND D a_543_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_629_125# a_27_57# a_747_79# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_962_371# a_1005_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X26 a_747_79# a_27_57# a_962_371# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 a_1784_75# a_1429_383# a_1583_285# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_543_125# D a_629_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR a_1583_285# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
