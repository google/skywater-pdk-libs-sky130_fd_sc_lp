* NGSPICE file created from sky130_fd_sc_lp__dfbbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dfbbn_2 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
M1000 VGND a_1746_137# a_1698_163# VNB nshort w=420000u l=150000u
+  ad=2.4516e+12p pd=2.023e+07u as=1.008e+11p ps=1.32e+06u
M1001 VGND RESET_B a_1191_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1002 VGND a_113_57# a_223_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1003 a_1018_60# a_1191_21# a_789_78# VNB nshort w=640000u l=150000u
+  ad=3.648e+11p pd=3.7e+06u as=3.69e+11p ps=2.81e+06u
M1004 a_1746_137# a_1542_428# a_1911_119# VNB nshort w=640000u l=150000u
+  ad=3.5555e+11p pd=2.67e+06u as=3.776e+11p ps=3.74e+06u
M1005 a_1447_379# a_789_78# VPWR VPB phighvt w=840000u l=150000u
+  ad=3.15875e+11p pd=2.82e+06u as=4.10265e+12p ps=2.971e+07u
M1006 VPWR a_1746_137# a_2618_131# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1007 Q a_2618_131# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1008 Q_N a_1746_137# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1009 VPWR a_1191_21# a_2048_428# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1010 a_789_78# a_549_449# a_1018_60# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_1746_137# Q_N VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1012 a_463_449# D VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1013 a_549_449# a_223_119# a_463_449# VNB nshort w=420000u l=150000u
+  ad=2.2125e+11p pd=1.94e+06u as=0p ps=0u
M1014 a_1746_137# SET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1015 a_1698_163# a_223_119# a_1542_428# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.643e+11p ps=2.47e+06u
M1016 a_1644_506# a_113_57# a_1542_428# VPB phighvt w=420000u l=150000u
+  ad=2.919e+11p pd=2.23e+06u as=2.6985e+11p ps=2.4e+06u
M1017 a_1018_60# SET_B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_2618_131# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1019 a_1542_428# a_113_57# a_1447_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.304e+11p ps=2e+06u
M1020 a_1542_428# a_223_119# a_1447_379# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_1746_137# a_1644_506# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_2048_428# a_1542_428# a_1746_137# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_549_449# a_113_57# a_463_449# VPB phighvt w=420000u l=150000u
+  ad=2.73e+11p pd=2.14e+06u as=1.176e+11p ps=1.4e+06u
M1024 a_789_78# SET_B VPWR VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1025 a_113_57# CLK_N VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1026 VPWR RESET_B a_1191_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1027 VPWR a_2618_131# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND a_1746_137# Q_N VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Q_N a_1746_137# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_709_449# a_223_119# a_549_449# VPB phighvt w=420000u l=150000u
+  ad=1.68e+11p pd=1.64e+06u as=0p ps=0u
M1031 a_1911_119# SET_B VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND a_1746_137# a_2618_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1033 VGND a_2618_131# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_113_57# CLK_N VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1035 VPWR a_113_57# a_223_119# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1036 VPWR a_1191_21# a_1119_379# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=3.024e+11p ps=2.4e+06u
M1037 VGND a_789_78# a_705_104# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
M1038 a_1911_119# a_1191_21# a_1746_137# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR a_789_78# a_709_449# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1119_379# a_549_449# a_789_78# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_705_104# a_113_57# a_549_449# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_463_449# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1447_119# a_789_78# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

