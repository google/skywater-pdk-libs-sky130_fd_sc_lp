* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
X0 Y a_27_535# a_312_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_27_535# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_27_535# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_672_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_312_367# C a_229_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_672_367# B a_229_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR A a_672_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 Y a_27_535# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_229_367# B a_672_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VGND a_27_535# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_312_367# a_27_535# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_229_367# C a_312_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
