* File: sky130_fd_sc_lp__or4bb_1.pxi.spice
* Created: Fri Aug 28 11:26:23 2020
* 
x_PM_SKY130_FD_SC_LP__OR4BB_1%C_N N_C_N_M1011_g N_C_N_M1008_g N_C_N_c_91_n
+ N_C_N_c_92_n N_C_N_c_93_n C_N C_N N_C_N_c_95_n PM_SKY130_FD_SC_LP__OR4BB_1%C_N
x_PM_SKY130_FD_SC_LP__OR4BB_1%D_N N_D_N_M1003_g N_D_N_M1009_g N_D_N_c_131_n D_N
+ D_N N_D_N_c_135_n N_D_N_c_132_n PM_SKY130_FD_SC_LP__OR4BB_1%D_N
x_PM_SKY130_FD_SC_LP__OR4BB_1%A_196_535# N_A_196_535#_M1009_d
+ N_A_196_535#_M1003_d N_A_196_535#_c_170_n N_A_196_535#_c_171_n
+ N_A_196_535#_M1010_g N_A_196_535#_M1000_g N_A_196_535#_c_173_n
+ N_A_196_535#_c_180_n N_A_196_535#_c_181_n N_A_196_535#_c_174_n
+ N_A_196_535#_c_175_n N_A_196_535#_c_176_n N_A_196_535#_c_177_n
+ PM_SKY130_FD_SC_LP__OR4BB_1%A_196_535#
x_PM_SKY130_FD_SC_LP__OR4BB_1%A_27_535# N_A_27_535#_M1008_s N_A_27_535#_M1011_s
+ N_A_27_535#_M1004_g N_A_27_535#_M1002_g N_A_27_535#_c_240_n
+ N_A_27_535#_c_241_n N_A_27_535#_c_242_n N_A_27_535#_c_250_n
+ N_A_27_535#_c_243_n N_A_27_535#_c_244_n N_A_27_535#_c_245_n
+ N_A_27_535#_c_246_n N_A_27_535#_c_247_n N_A_27_535#_c_248_n
+ PM_SKY130_FD_SC_LP__OR4BB_1%A_27_535#
x_PM_SKY130_FD_SC_LP__OR4BB_1%B N_B_M1013_g N_B_M1005_g B N_B_c_322_n
+ N_B_c_323_n N_B_c_324_n PM_SKY130_FD_SC_LP__OR4BB_1%B
x_PM_SKY130_FD_SC_LP__OR4BB_1%A N_A_M1007_g N_A_M1006_g A A A N_A_c_360_n
+ PM_SKY130_FD_SC_LP__OR4BB_1%A
x_PM_SKY130_FD_SC_LP__OR4BB_1%A_332_391# N_A_332_391#_M1010_d
+ N_A_332_391#_M1013_d N_A_332_391#_M1000_s N_A_332_391#_M1001_g
+ N_A_332_391#_M1012_g N_A_332_391#_c_408_n N_A_332_391#_c_395_n
+ N_A_332_391#_c_396_n N_A_332_391#_c_397_n N_A_332_391#_c_398_n
+ N_A_332_391#_c_399_n N_A_332_391#_c_400_n N_A_332_391#_c_401_n
+ N_A_332_391#_c_406_n N_A_332_391#_c_402_n N_A_332_391#_c_445_n
+ N_A_332_391#_c_403_n PM_SKY130_FD_SC_LP__OR4BB_1%A_332_391#
x_PM_SKY130_FD_SC_LP__OR4BB_1%VPWR N_VPWR_M1011_d N_VPWR_M1006_d N_VPWR_c_486_n
+ N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n VPWR N_VPWR_c_490_n
+ N_VPWR_c_491_n N_VPWR_c_485_n N_VPWR_c_493_n PM_SKY130_FD_SC_LP__OR4BB_1%VPWR
x_PM_SKY130_FD_SC_LP__OR4BB_1%X N_X_M1012_d N_X_M1001_d N_X_c_533_n N_X_c_534_n
+ X X X X N_X_c_532_n PM_SKY130_FD_SC_LP__OR4BB_1%X
x_PM_SKY130_FD_SC_LP__OR4BB_1%VGND N_VGND_M1008_d N_VGND_M1010_s N_VGND_M1004_d
+ N_VGND_M1007_d N_VGND_c_549_n N_VGND_c_550_n N_VGND_c_551_n N_VGND_c_552_n
+ VGND N_VGND_c_553_n N_VGND_c_554_n N_VGND_c_555_n N_VGND_c_556_n
+ N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n N_VGND_c_560_n N_VGND_c_561_n
+ PM_SKY130_FD_SC_LP__OR4BB_1%VGND
cc_1 VNB N_C_N_M1011_g 0.0131635f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_2 VNB N_C_N_c_91_n 0.0196719f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.765
cc_3 VNB N_C_N_c_92_n 0.023176f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.27
cc_4 VNB N_C_N_c_93_n 0.0163664f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.435
cc_5 VNB C_N 0.00646837f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_C_N_c_95_n 0.0162376f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.93
cc_7 VNB N_D_N_M1009_g 0.0528049f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.445
cc_8 VNB N_D_N_c_131_n 0.0112696f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_9 VNB N_D_N_c_132_n 0.00345589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_196_535#_c_170_n 0.0101575f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.93
cc_11 VNB N_A_196_535#_c_171_n 0.0270966f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.27
cc_12 VNB N_A_196_535#_M1000_g 0.013836f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.93
cc_13 VNB N_A_196_535#_c_173_n 0.0322753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_196_535#_c_174_n 0.00825998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_196_535#_c_175_n 0.0147655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_196_535#_c_176_n 0.0300758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_196_535#_c_177_n 0.0193466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_535#_c_240_n 0.0167621f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.93
cc_19 VNB N_A_27_535#_c_241_n 0.00853853f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.93
cc_20 VNB N_A_27_535#_c_242_n 0.0482576f $X=-0.19 $Y=-0.245 $X2=0.677 $Y2=0.925
cc_21 VNB N_A_27_535#_c_243_n 0.0143057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_535#_c_244_n 0.0061878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_535#_c_245_n 0.00159834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_535#_c_246_n 0.0156314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_535#_c_247_n 0.015089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_535#_c_248_n 0.0279881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_M1005_g 0.024834f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.445
cc_28 VNB N_B_c_322_n 0.0285838f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.435
cc_29 VNB N_B_c_323_n 0.00579758f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_30 VNB N_B_c_324_n 0.0167732f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_31 VNB N_A_M1007_g 0.0579281f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_32 VNB N_A_332_391#_M1001_g 0.00775413f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_33 VNB N_A_332_391#_c_395_n 0.00743608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_332_391#_c_396_n 0.00253571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_332_391#_c_397_n 8.99882e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_332_391#_c_398_n 0.0044919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_332_391#_c_399_n 0.012703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_332_391#_c_400_n 0.00990589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_332_391#_c_401_n 0.037602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_332_391#_c_402_n 0.00732342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_332_391#_c_403_n 0.0211127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_485_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_532_n 0.062609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_549_n 0.00232471f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.93
cc_45 VNB N_VGND_c_550_n 0.00583457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_551_n 4.06069e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_552_n 0.00494777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_553_n 0.0165364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_554_n 0.0139386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_555_n 0.0188323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_556_n 0.0152818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_557_n 0.231072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_558_n 0.0233782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_559_n 0.00484254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_560_n 0.00436942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_561_n 0.00455727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VPB N_C_N_M1011_g 0.0717697f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_58 VPB N_D_N_M1003_g 0.027991f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_59 VPB D_N 0.0209375f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_D_N_c_135_n 0.0289141f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=0.93
cc_61 VPB N_D_N_c_132_n 0.020996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_196_535#_c_170_n 0.0608954f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=0.93
cc_63 VPB N_A_196_535#_M1000_g 0.0276945f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=0.93
cc_64 VPB N_A_196_535#_c_180_n 0.0140673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_196_535#_c_181_n 0.0550212f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_27_535#_M1002_g 0.0186472f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_27_535#_c_250_n 0.0626308f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=0.93
cc_68 VPB N_A_27_535#_c_244_n 0.00640089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_27_535#_c_245_n 8.85151e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_27_535#_c_246_n 0.0120818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_27_535#_c_247_n 0.0165792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_B_M1005_g 0.0220141f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.445
cc_73 VPB N_A_M1007_g 0.0384508f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_74 VPB A 0.0214971f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=1.435
cc_75 VPB N_A_c_360_n 0.0535722f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=1.295
cc_76 VPB N_A_332_391#_M1001_g 0.0267564f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_77 VPB N_A_332_391#_c_397_n 0.00264377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_332_391#_c_406_n 0.00397565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_486_n 0.00522139f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=0.765
cc_80 VPB N_VPWR_c_487_n 0.0166236f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_81 VPB N_VPWR_c_488_n 0.0649395f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=0.93
cc_82 VPB N_VPWR_c_489_n 0.00574453f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=0.925
cc_83 VPB N_VPWR_c_490_n 0.0172362f $X=-0.19 $Y=1.655 $X2=0.677 $Y2=0.93
cc_84 VPB N_VPWR_c_491_n 0.0194887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_485_n 0.0685913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_493_n 0.00497572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_X_c_533_n 0.045918f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=0.765
cc_88 VPB N_X_c_534_n 0.00946635f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_89 VPB N_X_c_532_n 0.00889774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 N_C_N_M1011_g N_D_N_M1003_g 0.0202202f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_91 N_C_N_c_91_n N_D_N_M1009_g 0.012194f $X=0.53 $Y=0.765 $X2=0 $Y2=0
cc_92 C_N N_D_N_M1009_g 0.017128f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_93 N_C_N_c_95_n N_D_N_M1009_g 0.0432012f $X=0.53 $Y=0.93 $X2=0 $Y2=0
cc_94 N_C_N_M1011_g N_D_N_c_131_n 0.00559852f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_95 N_C_N_M1011_g D_N 0.0042882f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_96 N_C_N_M1011_g N_D_N_c_135_n 0.0162096f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_97 N_C_N_M1011_g N_D_N_c_132_n 0.0148381f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_98 C_N N_A_196_535#_c_173_n 5.83707e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_99 C_N N_A_196_535#_c_174_n 8.01585e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_100 C_N N_A_196_535#_c_175_n 0.0276536f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_101 C_N N_A_196_535#_c_176_n 0.00137768f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_102 N_C_N_M1011_g N_A_27_535#_c_242_n 0.00640807f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_103 N_C_N_c_91_n N_A_27_535#_c_242_n 0.00486785f $X=0.53 $Y=0.765 $X2=0 $Y2=0
cc_104 C_N N_A_27_535#_c_242_n 0.0520159f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_105 N_C_N_c_95_n N_A_27_535#_c_242_n 0.0162962f $X=0.53 $Y=0.93 $X2=0 $Y2=0
cc_106 N_C_N_M1011_g N_A_27_535#_c_250_n 0.0286313f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_107 N_C_N_c_91_n N_A_27_535#_c_243_n 0.00374726f $X=0.53 $Y=0.765 $X2=0 $Y2=0
cc_108 C_N N_A_27_535#_c_243_n 0.0034134f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_109 N_C_N_c_95_n N_A_27_535#_c_243_n 0.00276121f $X=0.53 $Y=0.93 $X2=0 $Y2=0
cc_110 N_C_N_c_93_n N_A_27_535#_c_244_n 0.0011869f $X=0.53 $Y=1.435 $X2=0 $Y2=0
cc_111 N_C_N_M1011_g N_A_27_535#_c_247_n 0.0186784f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_112 N_C_N_c_93_n N_A_27_535#_c_247_n 0.00139286f $X=0.53 $Y=1.435 $X2=0 $Y2=0
cc_113 C_N N_A_27_535#_c_247_n 0.0375945f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_114 N_C_N_M1011_g N_VPWR_c_486_n 0.00316145f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_115 N_C_N_M1011_g N_VPWR_c_490_n 0.00585385f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_116 N_C_N_M1011_g N_VPWR_c_485_n 0.0117692f $X=0.475 $Y=2.885 $X2=0 $Y2=0
cc_117 N_C_N_c_91_n N_VGND_c_549_n 0.00288325f $X=0.53 $Y=0.765 $X2=0 $Y2=0
cc_118 C_N N_VGND_c_549_n 0.0187241f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_119 N_C_N_c_91_n N_VGND_c_557_n 0.00706509f $X=0.53 $Y=0.765 $X2=0 $Y2=0
cc_120 C_N N_VGND_c_557_n 0.00706402f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_121 N_C_N_c_91_n N_VGND_c_558_n 0.0054833f $X=0.53 $Y=0.765 $X2=0 $Y2=0
cc_122 N_C_N_c_95_n N_VGND_c_558_n 3.19661e-19 $X=0.53 $Y=0.93 $X2=0 $Y2=0
cc_123 N_D_N_M1003_g N_A_196_535#_c_170_n 0.0173173f $X=0.905 $Y=2.885 $X2=0
+ $Y2=0
cc_124 N_D_N_c_131_n N_A_196_535#_c_170_n 0.0337542f $X=0.995 $Y=1.585 $X2=0
+ $Y2=0
cc_125 D_N N_A_196_535#_c_170_n 0.0105255f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_126 N_D_N_c_135_n N_A_196_535#_c_170_n 0.0181384f $X=0.955 $Y=2.22 $X2=0
+ $Y2=0
cc_127 N_D_N_M1009_g N_A_196_535#_c_173_n 0.00682193f $X=0.98 $Y=0.445 $X2=0
+ $Y2=0
cc_128 D_N N_A_196_535#_c_180_n 0.0264529f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_129 N_D_N_c_135_n N_A_196_535#_c_180_n 5.56561e-19 $X=0.955 $Y=2.22 $X2=0
+ $Y2=0
cc_130 N_D_N_M1009_g N_A_196_535#_c_174_n 0.00498506f $X=0.98 $Y=0.445 $X2=0
+ $Y2=0
cc_131 N_D_N_M1009_g N_A_196_535#_c_175_n 0.0035222f $X=0.98 $Y=0.445 $X2=0
+ $Y2=0
cc_132 N_D_N_M1009_g N_A_196_535#_c_176_n 0.0111144f $X=0.98 $Y=0.445 $X2=0
+ $Y2=0
cc_133 D_N N_A_27_535#_c_250_n 0.0442145f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_134 N_D_N_c_131_n N_A_27_535#_c_247_n 6.65464e-19 $X=0.995 $Y=1.585 $X2=0
+ $Y2=0
cc_135 D_N N_A_27_535#_c_247_n 0.0475354f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_136 N_D_N_c_135_n N_A_27_535#_c_247_n 0.00106549f $X=0.955 $Y=2.22 $X2=0
+ $Y2=0
cc_137 N_D_N_c_132_n N_A_27_535#_c_247_n 0.0161244f $X=0.955 $Y=2.055 $X2=0
+ $Y2=0
cc_138 D_N N_A_332_391#_c_406_n 0.0172342f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_139 N_D_N_M1003_g N_VPWR_c_486_n 0.00316145f $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_140 D_N N_VPWR_c_486_n 0.0182727f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_141 N_D_N_M1003_g N_VPWR_c_488_n 0.00585385f $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_142 N_D_N_M1003_g N_VPWR_c_485_n 0.00756726f $X=0.905 $Y=2.885 $X2=0 $Y2=0
cc_143 D_N N_VPWR_c_485_n 0.00736445f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_144 N_D_N_M1009_g N_VGND_c_549_n 0.00743965f $X=0.98 $Y=0.445 $X2=0 $Y2=0
cc_145 N_D_N_M1009_g N_VGND_c_550_n 0.00214139f $X=0.98 $Y=0.445 $X2=0 $Y2=0
cc_146 N_D_N_M1009_g N_VGND_c_553_n 0.00525069f $X=0.98 $Y=0.445 $X2=0 $Y2=0
cc_147 N_D_N_M1009_g N_VGND_c_557_n 0.0103725f $X=0.98 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A_196_535#_c_177_n N_A_27_535#_c_240_n 0.011568f $X=1.767 $Y=0.765
+ $X2=0 $Y2=0
cc_149 N_A_196_535#_c_176_n N_A_27_535#_c_241_n 0.00754808f $X=1.695 $Y=0.93
+ $X2=0 $Y2=0
cc_150 N_A_196_535#_M1000_g N_A_27_535#_c_245_n 5.27994e-19 $X=2 $Y=2.165 $X2=0
+ $Y2=0
cc_151 N_A_196_535#_M1000_g N_A_27_535#_c_246_n 0.0394498f $X=2 $Y=2.165 $X2=0
+ $Y2=0
cc_152 N_A_196_535#_c_170_n N_A_27_535#_c_247_n 0.0176554f $X=1.415 $Y=2.755
+ $X2=0 $Y2=0
cc_153 N_A_196_535#_M1000_g N_A_27_535#_c_247_n 0.0144547f $X=2 $Y=2.165 $X2=0
+ $Y2=0
cc_154 N_A_196_535#_c_173_n N_A_27_535#_c_247_n 0.00176192f $X=2 $Y=1.36 $X2=0
+ $Y2=0
cc_155 N_A_196_535#_c_175_n N_A_27_535#_c_247_n 0.0368005f $X=1.695 $Y=0.93
+ $X2=0 $Y2=0
cc_156 N_A_196_535#_c_173_n N_A_27_535#_c_248_n 0.0394498f $X=2 $Y=1.36 $X2=0
+ $Y2=0
cc_157 N_A_196_535#_c_175_n N_A_27_535#_c_248_n 4.7474e-19 $X=1.695 $Y=0.93
+ $X2=0 $Y2=0
cc_158 N_A_196_535#_c_176_n N_A_27_535#_c_248_n 0.0145116f $X=1.695 $Y=0.93
+ $X2=0 $Y2=0
cc_159 N_A_196_535#_c_170_n A 0.0051146f $X=1.415 $Y=2.755 $X2=0 $Y2=0
cc_160 N_A_196_535#_M1000_g A 0.00636405f $X=2 $Y=2.165 $X2=0 $Y2=0
cc_161 N_A_196_535#_c_180_n A 0.0171195f $X=1.62 $Y=2.92 $X2=0 $Y2=0
cc_162 N_A_196_535#_c_181_n A 0.00177763f $X=1.62 $Y=2.92 $X2=0 $Y2=0
cc_163 N_A_196_535#_M1000_g N_A_332_391#_c_408_n 0.0115755f $X=2 $Y=2.165 $X2=0
+ $Y2=0
cc_164 N_A_196_535#_c_174_n N_A_332_391#_c_395_n 0.00438417f $X=1.195 $Y=0.445
+ $X2=0 $Y2=0
cc_165 N_A_196_535#_c_175_n N_A_332_391#_c_395_n 0.0328735f $X=1.695 $Y=0.93
+ $X2=0 $Y2=0
cc_166 N_A_196_535#_c_177_n N_A_332_391#_c_395_n 0.00552971f $X=1.767 $Y=0.765
+ $X2=0 $Y2=0
cc_167 N_A_196_535#_c_171_n N_A_332_391#_c_396_n 8.90226e-19 $X=1.767 $Y=1.285
+ $X2=0 $Y2=0
cc_168 N_A_196_535#_c_173_n N_A_332_391#_c_396_n 0.00416684f $X=2 $Y=1.36 $X2=0
+ $Y2=0
cc_169 N_A_196_535#_c_175_n N_A_332_391#_c_396_n 0.013937f $X=1.695 $Y=0.93
+ $X2=0 $Y2=0
cc_170 N_A_196_535#_c_170_n N_A_332_391#_c_406_n 0.00475494f $X=1.415 $Y=2.755
+ $X2=0 $Y2=0
cc_171 N_A_196_535#_c_180_n N_A_332_391#_c_406_n 0.00755477f $X=1.62 $Y=2.92
+ $X2=0 $Y2=0
cc_172 N_A_196_535#_c_181_n N_A_332_391#_c_406_n 9.96055e-19 $X=1.62 $Y=2.92
+ $X2=0 $Y2=0
cc_173 N_A_196_535#_c_180_n N_VPWR_c_488_n 0.0434973f $X=1.62 $Y=2.92 $X2=0
+ $Y2=0
cc_174 N_A_196_535#_c_181_n N_VPWR_c_488_n 0.00783734f $X=1.62 $Y=2.92 $X2=0
+ $Y2=0
cc_175 N_A_196_535#_M1003_d N_VPWR_c_485_n 0.00222647f $X=0.98 $Y=2.675 $X2=0
+ $Y2=0
cc_176 N_A_196_535#_M1000_g N_VPWR_c_485_n 0.00348423f $X=2 $Y=2.165 $X2=0 $Y2=0
cc_177 N_A_196_535#_c_180_n N_VPWR_c_485_n 0.0278542f $X=1.62 $Y=2.92 $X2=0
+ $Y2=0
cc_178 N_A_196_535#_c_181_n N_VPWR_c_485_n 0.0149333f $X=1.62 $Y=2.92 $X2=0
+ $Y2=0
cc_179 N_A_196_535#_c_174_n N_VGND_c_550_n 0.0245336f $X=1.195 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_196_535#_c_175_n N_VGND_c_550_n 0.0211376f $X=1.695 $Y=0.93 $X2=0
+ $Y2=0
cc_181 N_A_196_535#_c_176_n N_VGND_c_550_n 0.00809343f $X=1.695 $Y=0.93 $X2=0
+ $Y2=0
cc_182 N_A_196_535#_c_177_n N_VGND_c_550_n 0.00796437f $X=1.767 $Y=0.765 $X2=0
+ $Y2=0
cc_183 N_A_196_535#_c_177_n N_VGND_c_551_n 5.76268e-19 $X=1.767 $Y=0.765 $X2=0
+ $Y2=0
cc_184 N_A_196_535#_c_174_n N_VGND_c_553_n 0.0153188f $X=1.195 $Y=0.445 $X2=0
+ $Y2=0
cc_185 N_A_196_535#_c_176_n N_VGND_c_553_n 3.91476e-19 $X=1.695 $Y=0.93 $X2=0
+ $Y2=0
cc_186 N_A_196_535#_c_177_n N_VGND_c_554_n 0.00564095f $X=1.767 $Y=0.765 $X2=0
+ $Y2=0
cc_187 N_A_196_535#_M1009_d N_VGND_c_557_n 0.00337718f $X=1.055 $Y=0.235 $X2=0
+ $Y2=0
cc_188 N_A_196_535#_c_174_n N_VGND_c_557_n 0.0102015f $X=1.195 $Y=0.445 $X2=0
+ $Y2=0
cc_189 N_A_196_535#_c_175_n N_VGND_c_557_n 0.00798375f $X=1.695 $Y=0.93 $X2=0
+ $Y2=0
cc_190 N_A_196_535#_c_176_n N_VGND_c_557_n 5.61188e-19 $X=1.695 $Y=0.93 $X2=0
+ $Y2=0
cc_191 N_A_196_535#_c_177_n N_VGND_c_557_n 0.00961799f $X=1.767 $Y=0.765 $X2=0
+ $Y2=0
cc_192 N_A_27_535#_M1002_g N_B_M1005_g 0.0215932f $X=2.36 $Y=2.165 $X2=0 $Y2=0
cc_193 N_A_27_535#_c_245_n N_B_M1005_g 3.06707e-19 $X=2.45 $Y=1.63 $X2=0 $Y2=0
cc_194 N_A_27_535#_c_246_n N_B_M1005_g 0.0211763f $X=2.45 $Y=1.63 $X2=0 $Y2=0
cc_195 N_A_27_535#_c_248_n N_B_M1005_g 0.0108359f $X=2.45 $Y=1.465 $X2=0 $Y2=0
cc_196 N_A_27_535#_c_241_n N_B_c_322_n 0.0199701f $X=2.345 $Y=0.915 $X2=0 $Y2=0
cc_197 N_A_27_535#_c_241_n N_B_c_323_n 0.0019369f $X=2.345 $Y=0.915 $X2=0 $Y2=0
cc_198 N_A_27_535#_c_240_n N_B_c_324_n 0.0104785f $X=2.345 $Y=0.765 $X2=0 $Y2=0
cc_199 N_A_27_535#_M1002_g A 0.0131317f $X=2.36 $Y=2.165 $X2=0 $Y2=0
cc_200 N_A_27_535#_M1002_g N_A_332_391#_c_408_n 0.0105109f $X=2.36 $Y=2.165
+ $X2=0 $Y2=0
cc_201 N_A_27_535#_c_246_n N_A_332_391#_c_408_n 0.00391065f $X=2.45 $Y=1.63
+ $X2=0 $Y2=0
cc_202 N_A_27_535#_c_247_n N_A_332_391#_c_408_n 0.0444538f $X=2.285 $Y=1.665
+ $X2=0 $Y2=0
cc_203 N_A_27_535#_c_240_n N_A_332_391#_c_395_n 0.00293004f $X=2.345 $Y=0.765
+ $X2=0 $Y2=0
cc_204 N_A_27_535#_c_241_n N_A_332_391#_c_395_n 0.00289423f $X=2.345 $Y=0.915
+ $X2=0 $Y2=0
cc_205 N_A_27_535#_c_248_n N_A_332_391#_c_395_n 0.00537973f $X=2.45 $Y=1.465
+ $X2=0 $Y2=0
cc_206 N_A_27_535#_c_247_n N_A_332_391#_c_396_n 0.0144987f $X=2.285 $Y=1.665
+ $X2=0 $Y2=0
cc_207 N_A_27_535#_M1002_g N_A_332_391#_c_397_n 0.00278486f $X=2.36 $Y=2.165
+ $X2=0 $Y2=0
cc_208 N_A_27_535#_c_245_n N_A_332_391#_c_397_n 0.0194098f $X=2.45 $Y=1.63 $X2=0
+ $Y2=0
cc_209 N_A_27_535#_c_246_n N_A_332_391#_c_397_n 9.87041e-19 $X=2.45 $Y=1.63
+ $X2=0 $Y2=0
cc_210 N_A_27_535#_c_246_n N_A_332_391#_c_399_n 0.00159052f $X=2.45 $Y=1.63
+ $X2=0 $Y2=0
cc_211 N_A_27_535#_c_248_n N_A_332_391#_c_399_n 0.00228905f $X=2.45 $Y=1.465
+ $X2=0 $Y2=0
cc_212 N_A_27_535#_c_247_n N_A_332_391#_c_406_n 0.0203904f $X=2.285 $Y=1.665
+ $X2=0 $Y2=0
cc_213 N_A_27_535#_c_241_n N_A_332_391#_c_402_n 7.45437e-19 $X=2.345 $Y=0.915
+ $X2=0 $Y2=0
cc_214 N_A_27_535#_c_245_n N_A_332_391#_c_402_n 0.0237947f $X=2.45 $Y=1.63 $X2=0
+ $Y2=0
cc_215 N_A_27_535#_c_246_n N_A_332_391#_c_402_n 0.00438376f $X=2.45 $Y=1.63
+ $X2=0 $Y2=0
cc_216 N_A_27_535#_c_247_n N_A_332_391#_c_402_n 0.00138747f $X=2.285 $Y=1.665
+ $X2=0 $Y2=0
cc_217 N_A_27_535#_c_248_n N_A_332_391#_c_402_n 0.0149758f $X=2.45 $Y=1.465
+ $X2=0 $Y2=0
cc_218 N_A_27_535#_c_250_n N_VPWR_c_490_n 0.0170509f $X=0.26 $Y=2.885 $X2=0
+ $Y2=0
cc_219 N_A_27_535#_M1011_s N_VPWR_c_485_n 0.00255119f $X=0.135 $Y=2.675 $X2=0
+ $Y2=0
cc_220 N_A_27_535#_c_250_n N_VPWR_c_485_n 0.0116369f $X=0.26 $Y=2.885 $X2=0
+ $Y2=0
cc_221 N_A_27_535#_c_240_n N_VGND_c_550_n 5.73654e-19 $X=2.345 $Y=0.765 $X2=0
+ $Y2=0
cc_222 N_A_27_535#_c_240_n N_VGND_c_551_n 0.0070681f $X=2.345 $Y=0.765 $X2=0
+ $Y2=0
cc_223 N_A_27_535#_c_240_n N_VGND_c_554_n 0.00564095f $X=2.345 $Y=0.765 $X2=0
+ $Y2=0
cc_224 N_A_27_535#_c_241_n N_VGND_c_554_n 4.04329e-19 $X=2.345 $Y=0.915 $X2=0
+ $Y2=0
cc_225 N_A_27_535#_M1008_s N_VGND_c_557_n 0.00233781f $X=0.19 $Y=0.235 $X2=0
+ $Y2=0
cc_226 N_A_27_535#_c_240_n N_VGND_c_557_n 0.00961799f $X=2.345 $Y=0.765 $X2=0
+ $Y2=0
cc_227 N_A_27_535#_c_241_n N_VGND_c_557_n 5.53504e-19 $X=2.345 $Y=0.915 $X2=0
+ $Y2=0
cc_228 N_A_27_535#_c_243_n N_VGND_c_557_n 0.015474f $X=0.335 $Y=0.445 $X2=0
+ $Y2=0
cc_229 N_A_27_535#_c_243_n N_VGND_c_558_n 0.0222161f $X=0.335 $Y=0.445 $X2=0
+ $Y2=0
cc_230 N_B_c_322_n N_A_M1007_g 0.107025f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_231 N_B_c_323_n N_A_M1007_g 2.89286e-19 $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_232 N_B_c_324_n N_A_M1007_g 0.0123927f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_233 N_B_M1005_g A 0.0123009f $X=2.9 $Y=2.165 $X2=0 $Y2=0
cc_234 N_B_M1005_g N_A_c_360_n 0.00552254f $X=2.9 $Y=2.165 $X2=0 $Y2=0
cc_235 N_B_M1005_g N_A_332_391#_c_408_n 0.00838516f $X=2.9 $Y=2.165 $X2=0 $Y2=0
cc_236 N_B_c_323_n N_A_332_391#_c_395_n 0.0167736f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_237 N_B_M1005_g N_A_332_391#_c_397_n 0.0127601f $X=2.9 $Y=2.165 $X2=0 $Y2=0
cc_238 N_B_c_322_n N_A_332_391#_c_398_n 0.00444071f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_239 N_B_c_323_n N_A_332_391#_c_398_n 0.0181463f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_240 N_B_c_324_n N_A_332_391#_c_398_n 0.00208975f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_241 N_B_M1005_g N_A_332_391#_c_399_n 0.0139364f $X=2.9 $Y=2.165 $X2=0 $Y2=0
cc_242 N_B_c_322_n N_A_332_391#_c_402_n 0.00469133f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_243 N_B_c_323_n N_A_332_391#_c_402_n 0.0374792f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_244 N_B_c_322_n N_A_332_391#_c_445_n 8.93904e-19 $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_245 N_B_c_323_n N_A_332_391#_c_445_n 0.00169789f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_246 N_B_c_322_n N_VGND_c_551_n 0.00242887f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_247 N_B_c_323_n N_VGND_c_551_n 0.0196346f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_248 N_B_c_324_n N_VGND_c_551_n 0.00822034f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_249 N_B_c_322_n N_VGND_c_555_n 7.13906e-19 $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_250 N_B_c_324_n N_VGND_c_555_n 0.00564095f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_251 N_B_c_322_n N_VGND_c_557_n 9.35314e-19 $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_252 N_B_c_323_n N_VGND_c_557_n 0.00664607f $X=2.81 $Y=0.93 $X2=0 $Y2=0
cc_253 N_B_c_324_n N_VGND_c_557_n 0.00514335f $X=2.81 $Y=0.765 $X2=0 $Y2=0
cc_254 N_A_M1007_g N_A_332_391#_M1001_g 0.0273585f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_255 N_A_M1007_g N_A_332_391#_c_408_n 5.82194e-19 $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_256 A N_A_332_391#_c_408_n 0.0543926f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_257 N_A_M1007_g N_A_332_391#_c_397_n 0.00242271f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_258 N_A_M1007_g N_A_332_391#_c_398_n 0.0147844f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A_M1007_g N_A_332_391#_c_399_n 0.0143858f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_260 N_A_M1007_g N_A_332_391#_c_400_n 0.00407557f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_261 N_A_M1007_g N_A_332_391#_c_401_n 0.0213482f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_262 N_A_M1007_g N_A_332_391#_c_445_n 0.00764371f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_263 N_A_M1007_g N_A_332_391#_c_403_n 0.0157428f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_264 N_A_M1007_g N_VPWR_c_487_n 0.0124021f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_265 A N_VPWR_c_487_n 0.0543891f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_266 A N_VPWR_c_488_n 0.0531622f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_267 N_A_c_360_n N_VPWR_c_488_n 0.0124786f $X=3.26 $Y=2.91 $X2=0 $Y2=0
cc_268 A N_VPWR_c_485_n 0.0423988f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_269 N_A_c_360_n N_VPWR_c_485_n 0.0153244f $X=3.26 $Y=2.91 $X2=0 $Y2=0
cc_270 A A_415_391# 0.00106797f $X=3.035 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_271 A A_487_391# 0.00303654f $X=3.035 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_272 A A_595_391# 0.00433668f $X=3.035 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_273 N_A_M1007_g N_VGND_c_551_n 0.00114336f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_274 N_A_M1007_g N_VGND_c_552_n 0.00916805f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_275 N_A_M1007_g N_VGND_c_555_n 0.00377881f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_276 N_A_M1007_g N_VGND_c_557_n 0.00619706f $X=3.26 $Y=0.445 $X2=0 $Y2=0
cc_277 N_A_332_391#_M1001_g N_VPWR_c_487_n 0.00598076f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_278 N_A_332_391#_c_397_n N_VPWR_c_487_n 0.00556715f $X=2.88 $Y=1.965 $X2=0
+ $Y2=0
cc_279 N_A_332_391#_c_400_n N_VPWR_c_487_n 0.0176131f $X=3.71 $Y=1.36 $X2=0
+ $Y2=0
cc_280 N_A_332_391#_c_401_n N_VPWR_c_487_n 0.00280627f $X=3.71 $Y=1.36 $X2=0
+ $Y2=0
cc_281 N_A_332_391#_M1001_g N_VPWR_c_491_n 0.00585385f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_282 N_A_332_391#_M1001_g N_VPWR_c_485_n 0.012875f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_A_332_391#_c_408_n A_415_391# 0.00204597f $X=2.795 $Y=2.05 $X2=-0.19
+ $Y2=-0.245
cc_284 N_A_332_391#_c_408_n A_487_391# 0.00709855f $X=2.795 $Y=2.05 $X2=-0.19
+ $Y2=-0.245
cc_285 N_A_332_391#_M1001_g N_X_c_534_n 0.00341053f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_286 N_A_332_391#_c_401_n N_X_c_534_n 0.00102138f $X=3.71 $Y=1.36 $X2=0 $Y2=0
cc_287 N_A_332_391#_M1001_g N_X_c_532_n 0.0112229f $X=3.785 $Y=2.465 $X2=0 $Y2=0
cc_288 N_A_332_391#_c_398_n N_X_c_532_n 0.00378093f $X=3.24 $Y=1.195 $X2=0 $Y2=0
cc_289 N_A_332_391#_c_400_n N_X_c_532_n 0.0271104f $X=3.71 $Y=1.36 $X2=0 $Y2=0
cc_290 N_A_332_391#_c_403_n N_X_c_532_n 0.0147307f $X=3.732 $Y=1.195 $X2=0 $Y2=0
cc_291 N_A_332_391#_c_402_n N_VGND_c_551_n 7.33655e-19 $X=2.795 $Y=1.36 $X2=0
+ $Y2=0
cc_292 N_A_332_391#_c_398_n N_VGND_c_552_n 0.031021f $X=3.24 $Y=1.195 $X2=0
+ $Y2=0
cc_293 N_A_332_391#_c_400_n N_VGND_c_552_n 0.0221599f $X=3.71 $Y=1.36 $X2=0
+ $Y2=0
cc_294 N_A_332_391#_c_401_n N_VGND_c_552_n 0.00530449f $X=3.71 $Y=1.36 $X2=0
+ $Y2=0
cc_295 N_A_332_391#_c_445_n N_VGND_c_552_n 0.0256962f $X=3.24 $Y=0.445 $X2=0
+ $Y2=0
cc_296 N_A_332_391#_c_403_n N_VGND_c_552_n 0.0152762f $X=3.732 $Y=1.195 $X2=0
+ $Y2=0
cc_297 N_A_332_391#_c_395_n N_VGND_c_554_n 0.0119705f $X=2.145 $Y=0.445 $X2=0
+ $Y2=0
cc_298 N_A_332_391#_c_445_n N_VGND_c_555_n 0.0196454f $X=3.24 $Y=0.445 $X2=0
+ $Y2=0
cc_299 N_A_332_391#_c_403_n N_VGND_c_556_n 0.00486043f $X=3.732 $Y=1.195 $X2=0
+ $Y2=0
cc_300 N_A_332_391#_M1010_d N_VGND_c_557_n 0.00343705f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_301 N_A_332_391#_M1013_d N_VGND_c_557_n 0.00246149f $X=2.905 $Y=0.235 $X2=0
+ $Y2=0
cc_302 N_A_332_391#_c_395_n N_VGND_c_557_n 0.00875646f $X=2.145 $Y=0.445 $X2=0
+ $Y2=0
cc_303 N_A_332_391#_c_445_n N_VGND_c_557_n 0.0138301f $X=3.24 $Y=0.445 $X2=0
+ $Y2=0
cc_304 N_A_332_391#_c_403_n N_VGND_c_557_n 0.00917987f $X=3.732 $Y=1.195 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_485_n N_X_M1001_d 0.00336915f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_306 N_VPWR_c_491_n N_X_c_533_n 0.023184f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_307 N_VPWR_c_485_n N_X_c_533_n 0.0131407f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_487_n N_X_c_534_n 0.00131283f $X=3.57 $Y=1.98 $X2=0 $Y2=0
cc_309 N_X_c_532_n N_VGND_c_556_n 0.018528f $X=4.06 $Y=0.42 $X2=0 $Y2=0
cc_310 N_X_M1012_d N_VGND_c_557_n 0.00371702f $X=3.92 $Y=0.235 $X2=0 $Y2=0
cc_311 N_X_c_532_n N_VGND_c_557_n 0.0104192f $X=4.06 $Y=0.42 $X2=0 $Y2=0
