* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
X0 VGND a_1891_47# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 Q a_1891_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR RESET_B a_595_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_1449_133# a_1475_426# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Q a_1891_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_829_119# a_731_405# a_905_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR RESET_B a_1475_426# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 Q a_1891_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND a_1891_47# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_1891_47# a_1255_449# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_27_90# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 Q a_1891_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VPWR a_1891_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 a_731_405# a_216_462# a_1255_449# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 a_1891_47# a_1255_449# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_595_535# a_27_90# a_689_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 VPWR a_595_535# a_731_405# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 a_27_90# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_595_535# a_216_462# a_829_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VPWR D a_340_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VGND a_27_90# a_216_462# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VGND RESET_B a_531_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_340_535# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_340_535# a_27_90# a_595_535# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_1891_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_1475_426# a_1255_449# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_905_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_731_405# a_27_90# a_1255_449# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X28 a_1255_449# a_27_90# a_1449_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_1697_133# a_1255_449# a_1475_426# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_689_535# a_731_405# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_340_535# a_216_462# a_595_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VPWR a_27_90# a_216_462# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X33 a_531_119# D a_340_535# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VGND a_595_535# a_731_405# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 VGND RESET_B a_1697_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_1255_449# a_216_462# a_1380_488# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 a_1380_488# a_1475_426# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
