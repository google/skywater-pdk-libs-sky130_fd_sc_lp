* File: sky130_fd_sc_lp__o41a_1.pxi.spice
* Created: Wed Sep  2 10:27:26 2020
* 
x_PM_SKY130_FD_SC_LP__O41A_1%A_155_23# N_A_155_23#_M1002_s N_A_155_23#_M1010_d
+ N_A_155_23#_c_68_n N_A_155_23#_M1001_g N_A_155_23#_M1008_g N_A_155_23#_c_70_n
+ N_A_155_23#_c_71_n N_A_155_23#_c_77_p N_A_155_23#_c_101_p N_A_155_23#_c_78_p
+ N_A_155_23#_c_79_p N_A_155_23#_c_72_n N_A_155_23#_c_73_n
+ PM_SKY130_FD_SC_LP__O41A_1%A_155_23#
x_PM_SKY130_FD_SC_LP__O41A_1%B1 N_B1_M1010_g N_B1_M1002_g B1 N_B1_c_122_n
+ N_B1_c_123_n PM_SKY130_FD_SC_LP__O41A_1%B1
x_PM_SKY130_FD_SC_LP__O41A_1%A4 N_A4_M1000_g N_A4_M1005_g A4 A4 A4 A4
+ N_A4_c_157_n N_A4_c_158_n PM_SKY130_FD_SC_LP__O41A_1%A4
x_PM_SKY130_FD_SC_LP__O41A_1%A3 N_A3_M1006_g N_A3_M1004_g A3 A3 A3 A3
+ N_A3_c_195_n N_A3_c_196_n PM_SKY130_FD_SC_LP__O41A_1%A3
x_PM_SKY130_FD_SC_LP__O41A_1%A2 N_A2_M1007_g N_A2_M1009_g A2 A2 A2 A2
+ N_A2_c_234_n N_A2_c_235_n A2 PM_SKY130_FD_SC_LP__O41A_1%A2
x_PM_SKY130_FD_SC_LP__O41A_1%A1 N_A1_M1011_g N_A1_M1003_g A1 N_A1_c_271_n
+ N_A1_c_272_n PM_SKY130_FD_SC_LP__O41A_1%A1
x_PM_SKY130_FD_SC_LP__O41A_1%X N_X_M1001_s N_X_M1008_s X X X X X X X N_X_c_296_n
+ PM_SKY130_FD_SC_LP__O41A_1%X
x_PM_SKY130_FD_SC_LP__O41A_1%VPWR N_VPWR_M1008_d N_VPWR_M1003_d N_VPWR_c_311_n
+ N_VPWR_c_312_n N_VPWR_c_313_n VPWR N_VPWR_c_314_n N_VPWR_c_315_n
+ N_VPWR_c_316_n N_VPWR_c_310_n PM_SKY130_FD_SC_LP__O41A_1%VPWR
x_PM_SKY130_FD_SC_LP__O41A_1%VGND N_VGND_M1001_d N_VGND_M1005_d N_VGND_M1007_d
+ N_VGND_c_362_n N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n
+ VGND N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n N_VGND_c_370_n
+ N_VGND_c_371_n N_VGND_c_372_n PM_SKY130_FD_SC_LP__O41A_1%VGND
x_PM_SKY130_FD_SC_LP__O41A_1%A_375_49# N_A_375_49#_M1002_d N_A_375_49#_M1004_d
+ N_A_375_49#_M1011_d N_A_375_49#_c_448_n N_A_375_49#_c_414_n
+ N_A_375_49#_c_415_n N_A_375_49#_c_427_n N_A_375_49#_c_416_n
+ N_A_375_49#_c_417_n N_A_375_49#_c_418_n PM_SKY130_FD_SC_LP__O41A_1%A_375_49#
cc_1 VNB N_A_155_23#_c_68_n 0.022531f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.195
cc_2 VNB N_A_155_23#_M1008_g 0.00841824f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.465
cc_3 VNB N_A_155_23#_c_70_n 0.00257556f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.925
cc_4 VNB N_A_155_23#_c_71_n 0.00797466f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.42
cc_5 VNB N_A_155_23#_c_72_n 0.0299615f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.26
cc_6 VNB N_A_155_23#_c_73_n 0.037382f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.36
cc_7 VNB N_B1_M1002_g 0.0291049f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.195
cc_8 VNB N_B1_c_122_n 0.003958f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.925
cc_9 VNB N_B1_c_123_n 0.0273426f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.995
cc_10 VNB N_A4_M1005_g 0.0257532f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.195
cc_11 VNB N_A4_c_157_n 0.0239216f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.42
cc_12 VNB N_A4_c_158_n 0.0029157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A3_M1004_g 0.0257474f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.195
cc_14 VNB N_A3_c_195_n 0.0242844f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.42
cc_15 VNB N_A3_c_196_n 0.00463619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_M1007_g 0.025264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_234_n 0.0240294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_235_n 0.00360173f $X=-0.19 $Y=-0.245 $X2=1.655 $Y2=2.012
cc_19 VNB N_A1_M1011_g 0.0296502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_M1003_g 0.00154344f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.195
cc_21 VNB N_A1_c_271_n 0.0533793f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.525
cc_22 VNB N_A1_c_272_n 0.0122349f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.925
cc_23 VNB X 0.0272814f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=0.665
cc_24 VNB X 0.0165371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_296_n 0.0297953f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.995
cc_26 VNB N_VPWR_c_310_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_362_n 0.00867586f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.465
cc_28 VNB N_VGND_c_363_n 0.00599613f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.995
cc_29 VNB N_VGND_c_364_n 0.0059479f $X=-0.19 $Y=-0.245 $X2=1.655 $Y2=2.012
cc_30 VNB N_VGND_c_365_n 0.0303463f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=2.91
cc_31 VNB N_VGND_c_366_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=2.91
cc_32 VNB N_VGND_c_367_n 0.023753f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.36
cc_33 VNB N_VGND_c_368_n 0.0182639f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.36
cc_34 VNB N_VGND_c_369_n 0.0193877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_370_n 0.239941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_371_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_372_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_375_49#_c_414_n 0.00603542f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.525
cc_39 VNB N_A_375_49#_c_415_n 0.00854014f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.925
cc_40 VNB N_A_375_49#_c_416_n 0.013185f $X=-0.19 $Y=-0.245 $X2=1.655 $Y2=2.012
cc_41 VNB N_A_375_49#_c_417_n 0.0289544f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=2.91
cc_42 VNB N_A_375_49#_c_418_n 0.0090164f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.26
cc_43 VPB N_A_155_23#_M1008_g 0.02565f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.465
cc_44 VPB N_A_155_23#_c_70_n 0.0038112f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=1.925
cc_45 VPB N_B1_M1010_g 0.021521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_B1_c_122_n 0.00268066f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=1.925
cc_47 VPB N_B1_c_123_n 0.00698171f $X=-0.19 $Y=1.655 $X2=1.565 $Y2=0.995
cc_48 VPB N_A4_M1000_g 0.0206415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A4_c_157_n 0.00819544f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.42
cc_50 VPB N_A4_c_158_n 0.00267032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A3_M1006_g 0.0196024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A3_c_195_n 0.00635236f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=0.42
cc_53 VPB N_A3_c_196_n 0.00238465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A2_M1009_g 0.0197678f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.195
cc_55 VPB A2 0.0013524f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=0.665
cc_56 VPB N_A2_c_234_n 0.00638194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A1_M1003_g 0.0266609f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.195
cc_58 VPB N_A1_c_272_n 0.0097044f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=1.925
cc_59 VPB X 0.0870315f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_311_n 0.00557321f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=0.665
cc_61 VPB N_VPWR_c_312_n 0.0129531f $X=-0.19 $Y=1.655 $X2=1.035 $Y2=2.465
cc_62 VPB N_VPWR_c_313_n 0.0503368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_314_n 0.0309953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_315_n 0.0644349f $X=-0.19 $Y=1.655 $X2=1.82 $Y2=2.91
cc_65 VPB N_VPWR_c_316_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0.85 $Y2=1.36
cc_66 VPB N_VPWR_c_310_n 0.0491418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 N_A_155_23#_M1008_g N_B1_M1010_g 0.0201967f $X=1.035 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A_155_23#_c_77_p N_B1_M1010_g 0.0133518f $X=1.655 $Y=2.012 $X2=0 $Y2=0
cc_69 N_A_155_23#_c_78_p N_B1_M1010_g 7.47598e-19 $X=1.78 $Y=2.1 $X2=0 $Y2=0
cc_70 N_A_155_23#_c_79_p N_B1_M1010_g 0.0123107f $X=1.82 $Y=2.91 $X2=0 $Y2=0
cc_71 N_A_155_23#_c_72_n N_B1_M1002_g 0.00668794f $X=1.34 $Y=1.26 $X2=0 $Y2=0
cc_72 N_A_155_23#_c_73_n N_B1_M1002_g 0.00184162f $X=1.035 $Y=1.36 $X2=0 $Y2=0
cc_73 N_A_155_23#_c_70_n N_B1_c_122_n 0.0167536f $X=1.34 $Y=1.925 $X2=0 $Y2=0
cc_74 N_A_155_23#_c_77_p N_B1_c_122_n 0.00418166f $X=1.655 $Y=2.012 $X2=0 $Y2=0
cc_75 N_A_155_23#_c_78_p N_B1_c_122_n 0.0188216f $X=1.78 $Y=2.1 $X2=0 $Y2=0
cc_76 N_A_155_23#_c_72_n N_B1_c_122_n 0.0244296f $X=1.34 $Y=1.26 $X2=0 $Y2=0
cc_77 N_A_155_23#_c_70_n N_B1_c_123_n 0.00424553f $X=1.34 $Y=1.925 $X2=0 $Y2=0
cc_78 N_A_155_23#_c_78_p N_B1_c_123_n 0.00110665f $X=1.78 $Y=2.1 $X2=0 $Y2=0
cc_79 N_A_155_23#_c_72_n N_B1_c_123_n 0.00583278f $X=1.34 $Y=1.26 $X2=0 $Y2=0
cc_80 N_A_155_23#_c_73_n N_B1_c_123_n 0.0201967f $X=1.035 $Y=1.36 $X2=0 $Y2=0
cc_81 N_A_155_23#_c_78_p N_A4_M1000_g 7.389e-19 $X=1.78 $Y=2.1 $X2=0 $Y2=0
cc_82 N_A_155_23#_c_79_p N_A4_M1000_g 0.00541955f $X=1.82 $Y=2.91 $X2=0 $Y2=0
cc_83 N_A_155_23#_c_70_n N_A4_c_158_n 0.0037169f $X=1.34 $Y=1.925 $X2=0 $Y2=0
cc_84 N_A_155_23#_c_68_n X 0.0106555f $X=0.85 $Y=1.195 $X2=0 $Y2=0
cc_85 N_A_155_23#_c_72_n X 0.0232925f $X=1.34 $Y=1.26 $X2=0 $Y2=0
cc_86 N_A_155_23#_M1008_g X 0.0124789f $X=1.035 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A_155_23#_c_70_n X 0.00302057f $X=1.34 $Y=1.925 $X2=0 $Y2=0
cc_88 N_A_155_23#_c_72_n X 0.0159211f $X=1.34 $Y=1.26 $X2=0 $Y2=0
cc_89 N_A_155_23#_c_73_n X 0.00355657f $X=1.035 $Y=1.36 $X2=0 $Y2=0
cc_90 N_A_155_23#_c_70_n N_VPWR_M1008_d 0.00270126f $X=1.34 $Y=1.925 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A_155_23#_c_77_p N_VPWR_M1008_d 0.00229969f $X=1.655 $Y=2.012 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_155_23#_c_101_p N_VPWR_M1008_d 0.00476405f $X=1.425 $Y=2.012 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_155_23#_M1008_g N_VPWR_c_311_n 0.00816956f $X=1.035 $Y=2.465 $X2=0
+ $Y2=0
cc_94 N_A_155_23#_c_77_p N_VPWR_c_311_n 0.00387621f $X=1.655 $Y=2.012 $X2=0
+ $Y2=0
cc_95 N_A_155_23#_c_101_p N_VPWR_c_311_n 0.0152373f $X=1.425 $Y=2.012 $X2=0
+ $Y2=0
cc_96 N_A_155_23#_M1008_g N_VPWR_c_314_n 0.00585385f $X=1.035 $Y=2.465 $X2=0
+ $Y2=0
cc_97 N_A_155_23#_c_79_p N_VPWR_c_315_n 0.0153681f $X=1.82 $Y=2.91 $X2=0 $Y2=0
cc_98 N_A_155_23#_M1010_d N_VPWR_c_310_n 0.00925041f $X=1.68 $Y=1.835 $X2=0
+ $Y2=0
cc_99 N_A_155_23#_M1008_g N_VPWR_c_310_n 0.0123757f $X=1.035 $Y=2.465 $X2=0
+ $Y2=0
cc_100 N_A_155_23#_c_79_p N_VPWR_c_310_n 0.00945867f $X=1.82 $Y=2.91 $X2=0 $Y2=0
cc_101 N_A_155_23#_c_72_n N_VGND_M1001_d 0.00243438f $X=1.34 $Y=1.26 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_155_23#_c_68_n N_VGND_c_362_n 0.0125878f $X=0.85 $Y=1.195 $X2=0 $Y2=0
cc_103 N_A_155_23#_c_71_n N_VGND_c_362_n 0.0427038f $X=1.585 $Y=0.42 $X2=0 $Y2=0
cc_104 N_A_155_23#_c_72_n N_VGND_c_362_n 0.0229447f $X=1.34 $Y=1.26 $X2=0 $Y2=0
cc_105 N_A_155_23#_c_73_n N_VGND_c_362_n 7.95552e-19 $X=1.035 $Y=1.36 $X2=0
+ $Y2=0
cc_106 N_A_155_23#_c_71_n N_VGND_c_365_n 0.0188755f $X=1.585 $Y=0.42 $X2=0 $Y2=0
cc_107 N_A_155_23#_c_68_n N_VGND_c_367_n 0.00477554f $X=0.85 $Y=1.195 $X2=0
+ $Y2=0
cc_108 N_A_155_23#_M1002_s N_VGND_c_370_n 0.00264482f $X=1.46 $Y=0.245 $X2=0
+ $Y2=0
cc_109 N_A_155_23#_c_68_n N_VGND_c_370_n 0.00955784f $X=0.85 $Y=1.195 $X2=0
+ $Y2=0
cc_110 N_A_155_23#_c_71_n N_VGND_c_370_n 0.0111968f $X=1.585 $Y=0.42 $X2=0 $Y2=0
cc_111 N_A_155_23#_c_72_n N_A_375_49#_c_415_n 0.00786427f $X=1.34 $Y=1.26 $X2=0
+ $Y2=0
cc_112 N_B1_M1010_g N_A4_M1000_g 0.026581f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B1_M1002_g N_A4_M1005_g 0.0232458f $X=1.8 $Y=0.665 $X2=0 $Y2=0
cc_114 N_B1_c_122_n N_A4_c_157_n 0.00133066f $X=1.71 $Y=1.51 $X2=0 $Y2=0
cc_115 N_B1_c_123_n N_A4_c_157_n 0.0214174f $X=1.8 $Y=1.51 $X2=0 $Y2=0
cc_116 N_B1_M1010_g N_A4_c_158_n 0.00104466f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B1_c_122_n N_A4_c_158_n 0.0329562f $X=1.71 $Y=1.51 $X2=0 $Y2=0
cc_118 N_B1_c_123_n N_A4_c_158_n 9.68304e-19 $X=1.8 $Y=1.51 $X2=0 $Y2=0
cc_119 N_B1_M1010_g N_VPWR_c_311_n 0.00816956f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B1_M1010_g N_VPWR_c_315_n 0.0054895f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_121 N_B1_M1010_g N_VPWR_c_310_n 0.0105206f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_122 N_B1_M1002_g N_VGND_c_362_n 0.00308748f $X=1.8 $Y=0.665 $X2=0 $Y2=0
cc_123 N_B1_M1002_g N_VGND_c_365_n 0.00575161f $X=1.8 $Y=0.665 $X2=0 $Y2=0
cc_124 N_B1_M1002_g N_VGND_c_370_n 0.0121037f $X=1.8 $Y=0.665 $X2=0 $Y2=0
cc_125 N_B1_M1002_g N_A_375_49#_c_415_n 8.60087e-19 $X=1.8 $Y=0.665 $X2=0 $Y2=0
cc_126 N_B1_c_122_n N_A_375_49#_c_415_n 0.00216446f $X=1.71 $Y=1.51 $X2=0 $Y2=0
cc_127 N_A4_M1000_g N_A3_M1006_g 0.0338957f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A4_c_158_n N_A3_M1006_g 0.00314103f $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A4_M1005_g N_A3_M1004_g 0.0289901f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_130 N_A4_c_157_n N_A3_c_195_n 0.0204266f $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A4_c_158_n N_A3_c_195_n 2.89053e-19 $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A4_M1000_g N_A3_c_196_n 0.00435948f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A4_c_157_n N_A3_c_196_n 0.00226005f $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A4_c_158_n N_A3_c_196_n 0.13214f $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A4_M1000_g N_VPWR_c_315_n 0.00376756f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A4_c_158_n N_VPWR_c_315_n 0.00958105f $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_137 N_A4_M1000_g N_VPWR_c_310_n 0.00626345f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A4_c_158_n N_VPWR_c_310_n 0.0088053f $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_139 N_A4_c_158_n A_447_367# 0.011031f $X=2.25 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_140 N_A4_M1005_g N_VGND_c_363_n 0.00674143f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_141 N_A4_M1005_g N_VGND_c_365_n 0.00575161f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_142 N_A4_M1005_g N_VGND_c_370_n 0.0110467f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_143 N_A4_M1005_g N_A_375_49#_c_414_n 0.0145773f $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_144 N_A4_c_157_n N_A_375_49#_c_414_n 0.0032799f $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_145 N_A4_c_158_n N_A_375_49#_c_414_n 0.0141056f $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_146 N_A4_c_157_n N_A_375_49#_c_415_n 5.08317e-19 $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_147 N_A4_c_158_n N_A_375_49#_c_415_n 0.00663832f $X=2.25 $Y=1.51 $X2=0 $Y2=0
cc_148 N_A4_M1005_g N_A_375_49#_c_427_n 8.88496e-19 $X=2.23 $Y=0.665 $X2=0 $Y2=0
cc_149 N_A3_M1004_g N_A2_M1007_g 0.0250312f $X=2.81 $Y=0.665 $X2=0 $Y2=0
cc_150 N_A3_M1006_g N_A2_M1009_g 0.060168f $X=2.79 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A3_c_196_n N_A2_M1009_g 0.0101506f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_152 N_A3_M1006_g A2 0.00126863f $X=2.79 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A3_c_196_n A2 0.0652951f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_154 N_A3_c_195_n N_A2_c_234_n 0.020645f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_155 N_A3_c_196_n N_A2_c_234_n 0.00143766f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_156 N_A3_c_195_n N_A2_c_235_n 8.68844e-19 $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A3_c_196_n N_A2_c_235_n 0.0168235f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A3_M1006_g N_VPWR_c_315_n 0.00376756f $X=2.79 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A3_c_196_n N_VPWR_c_315_n 0.0168469f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A3_M1006_g N_VPWR_c_310_n 0.00602234f $X=2.79 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A3_c_196_n N_VPWR_c_310_n 0.0158226f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_162 N_A3_c_196_n A_447_367# 0.0138622f $X=2.79 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_163 N_A3_c_196_n A_573_367# 0.0133859f $X=2.79 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_164 N_A3_M1004_g N_VGND_c_363_n 0.00660861f $X=2.81 $Y=0.665 $X2=0 $Y2=0
cc_165 N_A3_M1004_g N_VGND_c_368_n 0.00539298f $X=2.81 $Y=0.665 $X2=0 $Y2=0
cc_166 N_A3_M1004_g N_VGND_c_370_n 0.0102217f $X=2.81 $Y=0.665 $X2=0 $Y2=0
cc_167 N_A3_M1004_g N_A_375_49#_c_414_n 0.0118338f $X=2.81 $Y=0.665 $X2=0 $Y2=0
cc_168 N_A3_c_195_n N_A_375_49#_c_414_n 7.73559e-19 $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A3_c_196_n N_A_375_49#_c_414_n 0.0283294f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A3_M1004_g N_A_375_49#_c_427_n 0.0113147f $X=2.81 $Y=0.665 $X2=0 $Y2=0
cc_171 N_A3_M1004_g N_A_375_49#_c_418_n 0.00179232f $X=2.81 $Y=0.665 $X2=0 $Y2=0
cc_172 N_A3_c_195_n N_A_375_49#_c_418_n 5.46117e-19 $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A3_c_196_n N_A_375_49#_c_418_n 0.00826793f $X=2.79 $Y=1.51 $X2=0 $Y2=0
cc_174 N_A2_M1007_g N_A1_M1011_g 0.0253971f $X=3.24 $Y=0.665 $X2=0 $Y2=0
cc_175 N_A2_M1009_g N_A1_M1003_g 0.0408443f $X=3.24 $Y=2.465 $X2=0 $Y2=0
cc_176 A2 N_A1_M1003_g 0.00626479f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_177 N_A2_c_234_n N_A1_c_271_n 0.0214632f $X=3.33 $Y=1.51 $X2=0 $Y2=0
cc_178 N_A2_c_235_n N_A1_c_271_n 0.00626479f $X=3.33 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A2_c_234_n N_A1_c_272_n 3.88071e-19 $X=3.33 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A2_c_235_n N_A1_c_272_n 0.0272941f $X=3.33 $Y=1.51 $X2=0 $Y2=0
cc_181 N_A2_M1009_g N_VPWR_c_315_n 0.00531141f $X=3.24 $Y=2.465 $X2=0 $Y2=0
cc_182 A2 N_VPWR_c_315_n 0.0159684f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_183 N_A2_M1009_g N_VPWR_c_310_n 0.00991678f $X=3.24 $Y=2.465 $X2=0 $Y2=0
cc_184 A2 N_VPWR_c_310_n 0.01525f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_185 A2 A_663_367# 0.0128018f $X=3.515 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_186 N_A2_M1007_g N_VGND_c_364_n 0.00640369f $X=3.24 $Y=0.665 $X2=0 $Y2=0
cc_187 N_A2_M1007_g N_VGND_c_368_n 0.00539298f $X=3.24 $Y=0.665 $X2=0 $Y2=0
cc_188 N_A2_M1007_g N_VGND_c_370_n 0.0101176f $X=3.24 $Y=0.665 $X2=0 $Y2=0
cc_189 N_A2_M1007_g N_A_375_49#_c_427_n 0.0110943f $X=3.24 $Y=0.665 $X2=0 $Y2=0
cc_190 N_A2_M1007_g N_A_375_49#_c_416_n 0.0120535f $X=3.24 $Y=0.665 $X2=0 $Y2=0
cc_191 N_A2_c_234_n N_A_375_49#_c_416_n 0.00419993f $X=3.33 $Y=1.51 $X2=0 $Y2=0
cc_192 N_A2_c_235_n N_A_375_49#_c_416_n 0.030172f $X=3.33 $Y=1.51 $X2=0 $Y2=0
cc_193 N_A2_M1007_g N_A_375_49#_c_418_n 0.00185816f $X=3.24 $Y=0.665 $X2=0 $Y2=0
cc_194 N_A2_c_235_n N_A_375_49#_c_418_n 0.00138319f $X=3.33 $Y=1.51 $X2=0 $Y2=0
cc_195 N_A1_M1003_g N_VPWR_c_313_n 0.00663507f $X=3.78 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A1_c_271_n N_VPWR_c_313_n 0.00159592f $X=4.03 $Y=1.46 $X2=0 $Y2=0
cc_197 N_A1_c_272_n N_VPWR_c_313_n 0.0237552f $X=4.03 $Y=1.46 $X2=0 $Y2=0
cc_198 N_A1_M1003_g N_VPWR_c_315_n 0.00585385f $X=3.78 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A1_M1003_g N_VPWR_c_310_n 0.0119068f $X=3.78 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A1_M1011_g N_VGND_c_364_n 0.00321818f $X=3.78 $Y=0.665 $X2=0 $Y2=0
cc_201 N_A1_M1011_g N_VGND_c_369_n 0.00575161f $X=3.78 $Y=0.665 $X2=0 $Y2=0
cc_202 N_A1_M1011_g N_VGND_c_370_n 0.0118051f $X=3.78 $Y=0.665 $X2=0 $Y2=0
cc_203 N_A1_M1011_g N_A_375_49#_c_427_n 3.91265e-19 $X=3.78 $Y=0.665 $X2=0 $Y2=0
cc_204 N_A1_M1011_g N_A_375_49#_c_416_n 0.0198947f $X=3.78 $Y=0.665 $X2=0 $Y2=0
cc_205 N_A1_c_271_n N_A_375_49#_c_416_n 0.00789219f $X=4.03 $Y=1.46 $X2=0 $Y2=0
cc_206 N_A1_c_272_n N_A_375_49#_c_416_n 0.0222271f $X=4.03 $Y=1.46 $X2=0 $Y2=0
cc_207 X N_VPWR_c_314_n 0.0586673f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_208 N_X_M1008_s N_VPWR_c_310_n 0.00618284f $X=0.355 $Y=1.835 $X2=0 $Y2=0
cc_209 X N_VPWR_c_310_n 0.0326573f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_210 N_X_c_296_n N_VGND_c_367_n 0.0449262f $X=0.295 $Y=0.4 $X2=0 $Y2=0
cc_211 N_X_M1001_s N_VGND_c_370_n 0.00642262f $X=0.17 $Y=0.245 $X2=0 $Y2=0
cc_212 N_X_c_296_n N_VGND_c_370_n 0.0249948f $X=0.295 $Y=0.4 $X2=0 $Y2=0
cc_213 N_VPWR_c_310_n A_447_367# 0.00998614f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_214 N_VPWR_c_310_n A_573_367# 0.00978224f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_215 N_VPWR_c_310_n A_663_367# 0.00365493f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_216 N_VGND_c_370_n N_A_375_49#_M1002_d 0.00258346f $X=4.08 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_217 N_VGND_c_370_n N_A_375_49#_M1004_d 0.00223559f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_370_n N_A_375_49#_M1011_d 0.00229694f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_365_n N_A_375_49#_c_448_n 0.015291f $X=2.35 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_370_n N_A_375_49#_c_448_n 0.0104192f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_M1005_d N_A_375_49#_c_414_n 0.00366523f $X=2.305 $Y=0.245 $X2=0
+ $Y2=0
cc_222 N_VGND_c_363_n N_A_375_49#_c_414_n 0.0257093f $X=2.515 $Y=0.37 $X2=0
+ $Y2=0
cc_223 N_VGND_c_368_n N_A_375_49#_c_427_n 0.0189236f $X=3.36 $Y=0 $X2=0 $Y2=0
cc_224 N_VGND_c_370_n N_A_375_49#_c_427_n 0.0123859f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_M1007_d N_A_375_49#_c_416_n 0.00306511f $X=3.315 $Y=0.245 $X2=0
+ $Y2=0
cc_226 N_VGND_c_364_n N_A_375_49#_c_416_n 0.022455f $X=3.525 $Y=0.37 $X2=0 $Y2=0
cc_227 N_VGND_c_369_n N_A_375_49#_c_417_n 0.0192303f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_370_n N_A_375_49#_c_417_n 0.0115856f $X=4.08 $Y=0 $X2=0 $Y2=0
