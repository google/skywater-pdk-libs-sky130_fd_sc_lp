* File: sky130_fd_sc_lp__a32o_1.pxi.spice
* Created: Wed Sep  2 09:27:34 2020
* 
x_PM_SKY130_FD_SC_LP__A32O_1%A_80_21# N_A_80_21#_M1004_d N_A_80_21#_M1003_d
+ N_A_80_21#_c_55_n N_A_80_21#_M1006_g N_A_80_21#_M1005_g N_A_80_21#_c_57_n
+ N_A_80_21#_c_58_n N_A_80_21#_c_68_p N_A_80_21#_c_130_p N_A_80_21#_c_63_n
+ N_A_80_21#_c_112_p N_A_80_21#_c_90_p N_A_80_21#_c_59_n N_A_80_21#_c_86_p
+ N_A_80_21#_c_60_n PM_SKY130_FD_SC_LP__A32O_1%A_80_21#
x_PM_SKY130_FD_SC_LP__A32O_1%A3 N_A3_M1008_g N_A3_M1002_g A3 N_A3_c_147_n
+ N_A3_c_148_n PM_SKY130_FD_SC_LP__A32O_1%A3
x_PM_SKY130_FD_SC_LP__A32O_1%A2 N_A2_M1000_g N_A2_M1007_g A2 N_A2_c_184_n
+ N_A2_c_185_n PM_SKY130_FD_SC_LP__A32O_1%A2
x_PM_SKY130_FD_SC_LP__A32O_1%A1 N_A1_c_215_n N_A1_M1004_g N_A1_M1009_g A1
+ N_A1_c_217_n N_A1_c_218_n PM_SKY130_FD_SC_LP__A32O_1%A1
x_PM_SKY130_FD_SC_LP__A32O_1%B1 N_B1_M1003_g N_B1_M1001_g B1 B1 N_B1_c_251_n
+ N_B1_c_252_n PM_SKY130_FD_SC_LP__A32O_1%B1
x_PM_SKY130_FD_SC_LP__A32O_1%B2 N_B2_M1010_g N_B2_M1011_g B2 B2 N_B2_c_284_n
+ PM_SKY130_FD_SC_LP__A32O_1%B2
x_PM_SKY130_FD_SC_LP__A32O_1%X N_X_M1006_s N_X_M1005_s X X X X X X X N_X_c_306_n
+ X PM_SKY130_FD_SC_LP__A32O_1%X
x_PM_SKY130_FD_SC_LP__A32O_1%VPWR N_VPWR_M1005_d N_VPWR_M1000_d N_VPWR_c_323_n
+ N_VPWR_c_324_n N_VPWR_c_325_n VPWR N_VPWR_c_326_n N_VPWR_c_322_n
+ N_VPWR_c_328_n N_VPWR_c_329_n PM_SKY130_FD_SC_LP__A32O_1%VPWR
x_PM_SKY130_FD_SC_LP__A32O_1%A_249_367# N_A_249_367#_M1008_d
+ N_A_249_367#_M1009_d N_A_249_367#_M1011_d N_A_249_367#_c_374_n
+ N_A_249_367#_c_379_n N_A_249_367#_c_375_n N_A_249_367#_c_393_n
+ N_A_249_367#_c_376_n N_A_249_367#_c_370_n N_A_249_367#_c_371_n
+ PM_SKY130_FD_SC_LP__A32O_1%A_249_367#
x_PM_SKY130_FD_SC_LP__A32O_1%VGND N_VGND_M1006_d N_VGND_M1010_d N_VGND_c_399_n
+ N_VGND_c_400_n VGND N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n
+ N_VGND_c_404_n PM_SKY130_FD_SC_LP__A32O_1%VGND
cc_1 VNB N_A_80_21#_c_55_n 0.0207782f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_A_80_21#_M1005_g 0.00766764f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_3 VNB N_A_80_21#_c_57_n 0.00217516f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.33
cc_4 VNB N_A_80_21#_c_58_n 0.00133699f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.705
cc_5 VNB N_A_80_21#_c_59_n 0.00330423f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.35
cc_6 VNB N_A_80_21#_c_60_n 0.0362598f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.35
cc_7 VNB N_A3_M1008_g 0.0073033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A3 0.00470223f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_9 VNB N_A3_c_147_n 0.0308884f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_10 VNB N_A3_c_148_n 0.0194953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_M1000_g 0.00904011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A2 0.00194146f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_13 VNB N_A2_c_184_n 0.0343133f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.465
cc_14 VNB N_A2_c_185_n 0.0174923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_215_n 0.0202546f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=0.235
cc_16 VNB N_A1_M1009_g 0.00853686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_217_n 0.00287441f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.025
cc_18 VNB N_A1_c_218_n 0.0352347f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.33
cc_19 VNB N_B1_M1003_g 0.00773905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B1 0.0166705f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_21 VNB N_B1_c_251_n 0.0276346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_252_n 0.0184743f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.33
cc_23 VNB N_B2_M1010_g 0.0227402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B2_M1011_g 0.00658167f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_25 VNB B2 0.0222133f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_26 VNB N_B2_c_284_n 0.049615f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.515
cc_27 VNB N_X_c_306_n 0.0607521f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=1.98
cc_28 VNB N_VPWR_c_322_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.515
cc_29 VNB N_VGND_c_399_n 0.0114821f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_30 VNB N_VGND_c_400_n 0.033989f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_31 VNB N_VGND_c_401_n 0.0161285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_402_n 0.0607664f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=0.94
cc_33 VNB N_VGND_c_403_n 0.0120967f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.35
cc_34 VNB N_VGND_c_404_n 0.209623f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.35
cc_35 VPB N_A_80_21#_M1005_g 0.0234587f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_36 VPB N_A_80_21#_c_58_n 4.84152e-19 $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.705
cc_37 VPB N_A_80_21#_c_63_n 0.0305729f $X=-0.19 $Y=1.655 $X2=2.92 $Y2=1.79
cc_38 VPB N_A3_M1008_g 0.0198121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A2_M1000_g 0.0219492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A1_M1009_g 0.0219691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_B1_M1003_g 0.0194596f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_B2_M1011_g 0.0260984f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_43 VPB B2 0.00919227f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_44 VPB X 0.0594156f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_45 VPB N_X_c_306_n 0.010228f $X=-0.19 $Y=1.655 $X2=3.085 $Y2=1.98
cc_46 VPB N_VPWR_c_323_n 0.00220706f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.465
cc_47 VPB N_VPWR_c_324_n 0.0156025f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.33
cc_48 VPB N_VPWR_c_325_n 0.00217586f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.94
cc_49 VPB N_VPWR_c_326_n 0.0363632f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.35
cc_50 VPB N_VPWR_c_322_n 0.0477842f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.515
cc_51 VPB N_VPWR_c_328_n 0.0249317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_329_n 0.0115892f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.35
cc_53 VPB N_A_249_367#_c_370_n 0.00746637f $X=-0.19 $Y=1.655 $X2=3.085 $Y2=1.875
cc_54 VPB N_A_249_367#_c_371_n 0.0374083f $X=-0.19 $Y=1.655 $X2=3.085 $Y2=1.98
cc_55 N_A_80_21#_M1005_g N_A3_M1008_g 0.0338848f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_56 N_A_80_21#_c_58_n N_A3_M1008_g 0.00365555f $X=0.8 $Y=1.705 $X2=0 $Y2=0
cc_57 N_A_80_21#_c_63_n N_A3_M1008_g 0.014675f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_58 N_A_80_21#_c_57_n A3 0.026015f $X=0.7 $Y=1.33 $X2=0 $Y2=0
cc_59 N_A_80_21#_c_68_p A3 0.0182007f $X=2.24 $Y=0.94 $X2=0 $Y2=0
cc_60 N_A_80_21#_c_63_n A3 0.0207668f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_60_n A3 2.81528e-19 $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_62 N_A_80_21#_M1005_g N_A3_c_147_n 5.06359e-19 $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_63 N_A_80_21#_c_57_n N_A3_c_147_n 0.00221465f $X=0.7 $Y=1.33 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_68_p N_A3_c_147_n 0.0036803f $X=2.24 $Y=0.94 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_63_n N_A3_c_147_n 0.00376271f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_60_n N_A3_c_147_n 0.0198604f $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_67 N_A_80_21#_c_55_n N_A3_c_148_n 0.0104545f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_57_n N_A3_c_148_n 0.00399897f $X=0.7 $Y=1.33 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_68_p N_A3_c_148_n 0.0132032f $X=2.24 $Y=0.94 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_60_n N_A3_c_148_n 2.42073e-19 $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_63_n N_A2_M1000_g 0.0118971f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_68_p A2 0.0213035f $X=2.24 $Y=0.94 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_63_n A2 0.0254327f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_68_p N_A2_c_184_n 0.00472955f $X=2.24 $Y=0.94 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_63_n N_A2_c_184_n 0.00133774f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_68_p N_A2_c_185_n 0.0124958f $X=2.24 $Y=0.94 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_86_p N_A2_c_185_n 0.00291174f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_68_p N_A1_c_215_n 0.00951859f $X=2.24 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_79 N_A_80_21#_c_86_p N_A1_c_215_n 0.0169475f $X=2.755 $Y=0.38 $X2=-0.19
+ $Y2=-0.245
cc_80 N_A_80_21#_c_63_n N_A1_M1009_g 0.0158158f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_90_p N_A1_M1009_g 7.68849e-19 $X=3.085 $Y=1.98 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_68_p N_A1_c_217_n 0.010592f $X=2.24 $Y=0.94 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_63_n N_A1_c_217_n 0.0210056f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_86_p N_A1_c_217_n 0.00757357f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_63_n N_A1_c_218_n 0.00593102f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_86_p N_A1_c_218_n 0.00896929f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_63_n N_B1_M1003_g 0.0139055f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_90_p N_B1_M1003_g 0.0126461f $X=3.085 $Y=1.98 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_63_n B1 0.0516284f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_86_p B1 0.0279833f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_63_n N_B1_c_251_n 0.00451068f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_86_p N_B1_c_251_n 0.00450532f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_86_p N_B1_c_252_n 0.0159643f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_86_p N_B2_M1010_g 0.00208412f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_63_n N_B2_M1011_g 0.00331168f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_63_n B2 0.00398213f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_59_n X 0.0011453f $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_60_n X 0.0048644f $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_55_n N_X_c_306_n 0.0134624f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_100 N_A_80_21#_M1005_g N_X_c_306_n 0.00636511f $X=0.665 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_57_n N_X_c_306_n 0.0361093f $X=0.7 $Y=1.33 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_58_n N_X_c_306_n 0.00783259f $X=0.8 $Y=1.705 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_112_p N_X_c_306_n 0.00659728f $X=0.885 $Y=1.79 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_63_n N_VPWR_M1005_d 0.00184604f $X=2.92 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_105 N_A_80_21#_c_112_p N_VPWR_M1005_d 0.00111404f $X=0.885 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_106 N_A_80_21#_c_63_n N_VPWR_M1000_d 0.00672213f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_107 N_A_80_21#_M1005_g N_VPWR_c_323_n 0.0157388f $X=0.665 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_A_80_21#_c_63_n N_VPWR_c_323_n 0.00991684f $X=2.92 $Y=1.79 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_112_p N_VPWR_c_323_n 0.00755868f $X=0.885 $Y=1.79 $X2=0
+ $Y2=0
cc_110 N_A_80_21#_M1003_d N_VPWR_c_322_n 0.00257355f $X=2.935 $Y=1.835 $X2=0
+ $Y2=0
cc_111 N_A_80_21#_M1005_g N_VPWR_c_322_n 0.00962569f $X=0.665 $Y=2.465 $X2=0
+ $Y2=0
cc_112 N_A_80_21#_M1005_g N_VPWR_c_328_n 0.00505556f $X=0.665 $Y=2.465 $X2=0
+ $Y2=0
cc_113 N_A_80_21#_c_63_n N_A_249_367#_M1008_d 0.00176461f $X=2.92 $Y=1.79
+ $X2=-0.19 $Y2=-0.245
cc_114 N_A_80_21#_c_63_n N_A_249_367#_M1009_d 0.00176461f $X=2.92 $Y=1.79 $X2=0
+ $Y2=0
cc_115 N_A_80_21#_c_63_n N_A_249_367#_c_374_n 0.0153678f $X=2.92 $Y=1.79 $X2=0
+ $Y2=0
cc_116 N_A_80_21#_c_63_n N_A_249_367#_c_375_n 0.0748484f $X=2.92 $Y=1.79 $X2=0
+ $Y2=0
cc_117 N_A_80_21#_M1003_d N_A_249_367#_c_376_n 0.00412427f $X=2.935 $Y=1.835
+ $X2=0 $Y2=0
cc_118 N_A_80_21#_c_90_p N_A_249_367#_c_376_n 0.0166396f $X=3.085 $Y=1.98 $X2=0
+ $Y2=0
cc_119 N_A_80_21#_c_57_n N_VGND_M1006_d 6.80172e-19 $X=0.7 $Y=1.33 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_80_21#_c_68_p N_VGND_M1006_d 0.00793859f $X=2.24 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_121 N_A_80_21#_c_130_p N_VGND_M1006_d 0.00432374f $X=0.885 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_80_21#_c_86_p N_VGND_c_400_n 0.0272671f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_55_n N_VGND_c_401_n 0.00565872f $X=0.475 $Y=1.185 $X2=0
+ $Y2=0
cc_124 N_A_80_21#_c_86_p N_VGND_c_402_n 0.043533f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_55_n N_VGND_c_403_n 0.0122534f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_68_p N_VGND_c_403_n 0.0198543f $X=2.24 $Y=0.94 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_130_p N_VGND_c_403_n 0.0248045f $X=0.885 $Y=0.94 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_60_n N_VGND_c_403_n 7.44406e-19 $X=0.665 $Y=1.35 $X2=0 $Y2=0
cc_129 N_A_80_21#_M1004_d N_VGND_c_404_n 0.00514095f $X=2.265 $Y=0.235 $X2=0
+ $Y2=0
cc_130 N_A_80_21#_c_55_n N_VGND_c_404_n 0.00950365f $X=0.475 $Y=1.185 $X2=0
+ $Y2=0
cc_131 N_A_80_21#_c_68_p N_VGND_c_404_n 0.0338082f $X=2.24 $Y=0.94 $X2=0 $Y2=0
cc_132 N_A_80_21#_c_130_p N_VGND_c_404_n 0.00216895f $X=0.885 $Y=0.94 $X2=0
+ $Y2=0
cc_133 N_A_80_21#_c_86_p N_VGND_c_404_n 0.0259931f $X=2.755 $Y=0.38 $X2=0 $Y2=0
cc_134 N_A_80_21#_c_68_p A_263_47# 0.0103214f $X=2.24 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A_80_21#_c_68_p A_356_47# 0.0117901f $X=2.24 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A3_M1008_g N_A2_M1000_g 0.0259984f $X=1.17 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A3_c_147_n N_A2_M1000_g 0.010661f $X=1.15 $Y=1.36 $X2=0 $Y2=0
cc_138 A3 A2 0.0253991f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A3_c_147_n A2 3.84419e-19 $X=1.15 $Y=1.36 $X2=0 $Y2=0
cc_140 A3 N_A2_c_184_n 0.00184765f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A3_c_148_n N_A2_c_184_n 0.010661f $X=1.145 $Y=1.195 $X2=0 $Y2=0
cc_142 N_A3_c_148_n N_A2_c_185_n 0.0455886f $X=1.145 $Y=1.195 $X2=0 $Y2=0
cc_143 N_A3_M1008_g N_VPWR_c_323_n 0.00684568f $X=1.17 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A3_M1008_g N_VPWR_c_324_n 0.00549284f $X=1.17 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A3_M1008_g N_VPWR_c_325_n 5.07426e-19 $X=1.17 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A3_M1008_g N_VPWR_c_322_n 0.0101093f $X=1.17 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A3_M1008_g N_A_249_367#_c_374_n 0.00268536f $X=1.17 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A3_M1008_g N_A_249_367#_c_379_n 0.00893581f $X=1.17 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A3_c_148_n N_VGND_c_402_n 0.00468308f $X=1.145 $Y=1.195 $X2=0 $Y2=0
cc_150 N_A3_c_148_n N_VGND_c_403_n 0.0189103f $X=1.145 $Y=1.195 $X2=0 $Y2=0
cc_151 N_A3_c_148_n N_VGND_c_404_n 0.00460479f $X=1.145 $Y=1.195 $X2=0 $Y2=0
cc_152 N_A2_c_184_n N_A1_c_215_n 0.0176441f $X=1.695 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A2_c_185_n N_A1_c_215_n 0.04193f $X=1.7 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_154 N_A2_M1000_g N_A1_M1009_g 0.015324f $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_155 A2 N_A1_c_217_n 0.0229817f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A2_c_184_n N_A1_c_217_n 0.0019281f $X=1.695 $Y=1.35 $X2=0 $Y2=0
cc_157 N_A2_M1000_g N_A1_c_218_n 2.35166e-19 $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_158 A2 N_A1_c_218_n 4.08683e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A2_M1000_g N_VPWR_c_324_n 0.00486043f $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A2_M1000_g N_VPWR_c_325_n 0.013855f $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A2_M1000_g N_VPWR_c_322_n 0.0082726f $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A2_M1000_g N_A_249_367#_c_375_n 0.0136831f $X=1.6 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A2_c_185_n N_VGND_c_402_n 0.00585385f $X=1.7 $Y=1.185 $X2=0 $Y2=0
cc_164 N_A2_c_185_n N_VGND_c_403_n 0.0032075f $X=1.7 $Y=1.185 $X2=0 $Y2=0
cc_165 N_A2_c_185_n N_VGND_c_404_n 0.00685103f $X=1.7 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A1_c_218_n N_B1_M1003_g 0.0306637f $X=2.43 $Y=1.36 $X2=0 $Y2=0
cc_167 N_A1_c_217_n B1 0.0246001f $X=2.28 $Y=1.36 $X2=0 $Y2=0
cc_168 N_A1_c_218_n B1 0.00265856f $X=2.43 $Y=1.36 $X2=0 $Y2=0
cc_169 N_A1_c_215_n N_B1_c_251_n 3.34595e-19 $X=2.19 $Y=1.195 $X2=0 $Y2=0
cc_170 N_A1_c_217_n N_B1_c_251_n 2.42841e-19 $X=2.28 $Y=1.36 $X2=0 $Y2=0
cc_171 N_A1_c_218_n N_B1_c_251_n 0.0200136f $X=2.43 $Y=1.36 $X2=0 $Y2=0
cc_172 N_A1_c_215_n N_B1_c_252_n 0.00690602f $X=2.19 $Y=1.195 $X2=0 $Y2=0
cc_173 N_A1_M1009_g N_VPWR_c_325_n 0.014802f $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A1_M1009_g N_VPWR_c_326_n 0.00486043f $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A1_M1009_g N_VPWR_c_322_n 0.0082726f $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A1_M1009_g N_A_249_367#_c_375_n 0.0136831f $X=2.43 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A1_c_215_n N_VGND_c_402_n 0.0054895f $X=2.19 $Y=1.195 $X2=0 $Y2=0
cc_178 N_A1_c_215_n N_VGND_c_404_n 0.00711786f $X=2.19 $Y=1.195 $X2=0 $Y2=0
cc_179 B1 N_B2_M1010_g 0.00317278f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_180 N_B1_c_252_n N_B2_M1010_g 0.0425966f $X=2.88 $Y=1.185 $X2=0 $Y2=0
cc_181 B1 B2 0.0257059f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_182 N_B1_c_251_n B2 2.05521e-19 $X=2.88 $Y=1.35 $X2=0 $Y2=0
cc_183 N_B1_M1003_g N_B2_c_284_n 0.0364699f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_184 N_B1_c_251_n N_B2_c_284_n 0.0425966f $X=2.88 $Y=1.35 $X2=0 $Y2=0
cc_185 N_B1_M1003_g N_VPWR_c_325_n 0.00115783f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_186 N_B1_M1003_g N_VPWR_c_326_n 0.00357877f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_187 N_B1_M1003_g N_VPWR_c_322_n 0.00550473f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_188 N_B1_M1003_g N_A_249_367#_c_376_n 0.0119874f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_189 N_B1_c_252_n N_VGND_c_400_n 0.00340288f $X=2.88 $Y=1.185 $X2=0 $Y2=0
cc_190 N_B1_c_252_n N_VGND_c_402_n 0.0054895f $X=2.88 $Y=1.185 $X2=0 $Y2=0
cc_191 N_B1_c_252_n N_VGND_c_404_n 0.0105069f $X=2.88 $Y=1.185 $X2=0 $Y2=0
cc_192 N_B2_M1011_g N_VPWR_c_326_n 0.00357877f $X=3.33 $Y=2.465 $X2=0 $Y2=0
cc_193 N_B2_M1011_g N_VPWR_c_322_n 0.00644349f $X=3.33 $Y=2.465 $X2=0 $Y2=0
cc_194 N_B2_M1011_g N_A_249_367#_c_376_n 0.0124156f $X=3.33 $Y=2.465 $X2=0 $Y2=0
cc_195 B2 N_A_249_367#_c_371_n 0.0232478f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_196 N_B2_c_284_n N_A_249_367#_c_371_n 0.00132803f $X=3.555 $Y=1.375 $X2=0
+ $Y2=0
cc_197 N_B2_M1010_g N_VGND_c_400_n 0.0231855f $X=3.33 $Y=0.655 $X2=0 $Y2=0
cc_198 B2 N_VGND_c_400_n 0.0229723f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_199 N_B2_c_284_n N_VGND_c_400_n 0.0021552f $X=3.555 $Y=1.375 $X2=0 $Y2=0
cc_200 N_B2_M1010_g N_VGND_c_402_n 0.00486043f $X=3.33 $Y=0.655 $X2=0 $Y2=0
cc_201 N_B2_M1010_g N_VGND_c_404_n 0.00818711f $X=3.33 $Y=0.655 $X2=0 $Y2=0
cc_202 N_X_M1005_s N_VPWR_c_322_n 0.00371702f $X=0.325 $Y=1.835 $X2=0 $Y2=0
cc_203 X N_VPWR_c_322_n 0.0174172f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_204 X N_VPWR_c_328_n 0.0314316f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_205 N_X_c_306_n N_VGND_c_401_n 0.0174563f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_206 N_X_M1006_s N_VGND_c_404_n 0.0040649f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_207 N_X_c_306_n N_VGND_c_404_n 0.00963639f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_208 N_VPWR_c_322_n N_A_249_367#_M1008_d 0.00380321f $X=3.6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_209 N_VPWR_c_322_n N_A_249_367#_M1009_d 0.00376626f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_322_n N_A_249_367#_M1011_d 0.00215159f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_324_n N_A_249_367#_c_379_n 0.0147495f $X=1.65 $Y=3.33 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_322_n N_A_249_367#_c_379_n 0.00979951f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_213 N_VPWR_M1000_d N_A_249_367#_c_375_n 0.0146615f $X=1.675 $Y=1.835 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_325_n N_A_249_367#_c_375_n 0.0496211f $X=2.215 $Y=2.5 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_326_n N_A_249_367#_c_393_n 0.0128782f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_322_n N_A_249_367#_c_393_n 0.00777554f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_326_n N_A_249_367#_c_376_n 0.0372417f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_218 N_VPWR_c_322_n N_A_249_367#_c_376_n 0.023676f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_219 N_VPWR_c_326_n N_A_249_367#_c_370_n 0.0189827f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_220 N_VPWR_c_322_n N_A_249_367#_c_370_n 0.0112745f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VGND_c_404_n A_263_47# 0.00469308f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_222 N_VGND_c_404_n A_356_47# 0.00499105f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_223 N_VGND_c_404_n A_609_47# 0.00899413f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
