* File: sky130_fd_sc_lp__o32ai_lp.spice
* Created: Fri Aug 28 11:18:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32ai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o32ai_lp  VNB VPB B1 B2 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_Y_M1009_d N_B1_M1009_g N_A_27_179#_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1533 PD=0.7 PS=1.57 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.3
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1003 N_A_27_179#_M1003_d N_B2_M1003_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.11125 AS=0.0588 PD=0.99 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A3_M1005_g N_A_27_179#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1281 AS=0.11125 PD=1.03 PS=0.99 NRD=71.424 NRS=22.848 M=1 R=2.8 SA=75001
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_A_27_179#_M1006_d N_A2_M1006_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1281 PD=0.7 PS=1.03 NRD=0 NRS=22.848 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A1_M1007_g N_A_27_179#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1533 AS=0.0588 PD=1.57 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1008 A_134_419# N_B1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g A_134_419# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1002 A_338_419# N_A3_M1002_g N_Y_M1000_d VPB PHIGHVT L=0.25 W=1 AD=0.1875
+ AS=0.14 PD=1.375 PS=1.28 NRD=26.0828 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1004 A_463_419# N_A2_M1004_g A_338_419# VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.1875 PD=1.32 PS=1.375 NRD=20.6653 NRS=26.0828 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_463_419# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=20.6653 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o32ai_lp.pxi.spice"
*
.ends
*
*
