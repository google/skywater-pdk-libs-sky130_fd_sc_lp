* File: sky130_fd_sc_lp__clkbuf_4.pex.spice
* Created: Wed Sep  2 09:38:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUF_4%A 3 6 8 11 13
r32 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.94
+ $X2=0.51 $Y2=1.105
r33 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.94
+ $X2=0.51 $Y2=0.775
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=0.94 $X2=0.51 $Y2=0.94
r35 8 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=0.94 $X2=0.51
+ $Y2=0.94
r36 6 14 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.105
r37 3 13 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_4%A_27_47# 1 2 9 13 17 21 25 29 33 37 40 43
+ 51 54 60 62 63 74
r96 73 74 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=2.245 $Y=1.37
+ $X2=2.25 $Y2=1.37
r97 70 71 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.815 $Y=1.37
+ $X2=1.82 $Y2=1.37
r98 69 70 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=1.39 $Y=1.37
+ $X2=1.815 $Y2=1.37
r99 68 69 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.385 $Y=1.37
+ $X2=1.39 $Y2=1.37
r100 64 66 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.955 $Y=1.37
+ $X2=0.96 $Y2=1.37
r101 57 60 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.44 $X2=0.26
+ $Y2=0.44
r102 55 73 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=1.92 $Y=1.37
+ $X2=2.245 $Y2=1.37
r103 55 71 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.92 $Y=1.37 $X2=1.82
+ $Y2=1.37
r104 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.37 $X2=1.92 $Y2=1.37
r105 52 68 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.24 $Y=1.37
+ $X2=1.385 $Y2=1.37
r106 52 66 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=1.24 $Y=1.37
+ $X2=0.96 $Y2=1.37
r107 51 63 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=1.37
+ $X2=1.075 $Y2=1.37
r108 51 54 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.24 $Y=1.37
+ $X2=1.92 $Y2=1.37
r109 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.24
+ $Y=1.37 $X2=1.24 $Y2=1.37
r110 48 62 1.05597 $w=2.6e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=1.405
+ $X2=0.24 $Y2=1.405
r111 48 63 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.395 $Y=1.405
+ $X2=1.075 $Y2=1.405
r112 43 45 31.7851 $w=3.08e-07 $l=8.55e-07 $layer=LI1_cond $X=0.24 $Y=2.04
+ $X2=0.24 $Y2=2.895
r113 41 62 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=0.24 $Y=1.535
+ $X2=0.24 $Y2=1.405
r114 41 43 18.7737 $w=3.08e-07 $l=5.05e-07 $layer=LI1_cond $X=0.24 $Y=1.535
+ $X2=0.24 $Y2=2.04
r115 40 62 5.51899 $w=2.4e-07 $l=1.61245e-07 $layer=LI1_cond $X=0.17 $Y=1.275
+ $X2=0.24 $Y2=1.405
r116 39 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.605
+ $X2=0.17 $Y2=0.44
r117 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=0.605
+ $X2=0.17 $Y2=1.275
r118 35 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.205
+ $X2=2.25 $Y2=1.37
r119 35 37 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=2.25 $Y=1.205
+ $X2=2.25 $Y2=0.445
r120 31 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.245 $Y=1.535
+ $X2=2.245 $Y2=1.37
r121 31 33 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.245 $Y=1.535
+ $X2=2.245 $Y2=2.465
r122 27 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=1.205
+ $X2=1.82 $Y2=1.37
r123 27 29 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.82 $Y=1.205
+ $X2=1.82 $Y2=0.445
r124 23 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.535
+ $X2=1.815 $Y2=1.37
r125 23 25 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=1.815 $Y=1.535
+ $X2=1.815 $Y2=2.465
r126 19 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.205
+ $X2=1.39 $Y2=1.37
r127 19 21 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.39 $Y=1.205
+ $X2=1.39 $Y2=0.445
r128 15 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.535
+ $X2=1.385 $Y2=1.37
r129 15 17 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=1.385 $Y=1.535
+ $X2=1.385 $Y2=2.465
r130 11 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.205
+ $X2=0.96 $Y2=1.37
r131 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.96 $Y=1.205
+ $X2=0.96 $Y2=0.445
r132 7 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.535
+ $X2=0.955 $Y2=1.37
r133 7 9 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=0.955 $Y=1.535
+ $X2=0.955 $Y2=2.465
r134 2 45 400 $w=1.7e-07 $l=1.12076e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.895
r135 2 43 400 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.04
r136 1 60 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_4%VPWR 1 2 3 12 18 22 24 29 30 31 33 42 47 51
r40 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 42 50 4.13232 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.607 $Y2=3.33
r45 42 44 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 41 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 38 47 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 38 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 36 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 33 47 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 33 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 31 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 31 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 29 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 29 30 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.475 $Y=3.33
+ $X2=1.602 $Y2=3.33
r58 28 44 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 28 30 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.73 $Y=3.33
+ $X2=1.602 $Y2=3.33
r60 24 27 28.3056 $w=2.83e-07 $l=7e-07 $layer=LI1_cond $X=2.477 $Y=2.23
+ $X2=2.477 $Y2=2.93
r61 22 50 3.26635 $w=2.85e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.477 $Y=3.245
+ $X2=2.607 $Y2=3.33
r62 22 27 12.7375 $w=2.83e-07 $l=3.15e-07 $layer=LI1_cond $X=2.477 $Y=3.245
+ $X2=2.477 $Y2=2.93
r63 18 21 31.6357 $w=2.53e-07 $l=7e-07 $layer=LI1_cond $X=1.602 $Y=2.23
+ $X2=1.602 $Y2=2.93
r64 16 30 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.602 $Y=3.245
+ $X2=1.602 $Y2=3.33
r65 16 21 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=1.602 $Y=3.245
+ $X2=1.602 $Y2=2.93
r66 12 15 31.7851 $w=3.08e-07 $l=8.55e-07 $layer=LI1_cond $X=0.72 $Y=2.04
+ $X2=0.72 $Y2=2.895
r67 10 47 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r68 10 15 13.0115 $w=3.08e-07 $l=3.5e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.895
r69 3 27 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.835 $X2=2.46 $Y2=2.93
r70 3 24 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.835 $X2=2.46 $Y2=2.23
r71 2 21 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.93
r72 2 18 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.23
r73 1 15 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.895
r74 1 12 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 38 39
+ 50
r61 45 50 1.40715 $w=5.08e-07 $l=6e-08 $layer=LI1_cond $X=2.51 $Y=1.725 $X2=2.51
+ $Y2=1.665
r62 44 51 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=2.51 $Y=0.9
+ $X2=2.035 $Y2=0.9
r63 39 45 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=1.81
+ $X2=2.51 $Y2=1.81
r64 39 50 0.304883 $w=5.08e-07 $l=1.3e-08 $layer=LI1_cond $X=2.51 $Y=1.652
+ $X2=2.51 $Y2=1.665
r65 38 39 8.37255 $w=5.08e-07 $l=3.57e-07 $layer=LI1_cond $X=2.51 $Y=1.295
+ $X2=2.51 $Y2=1.652
r66 38 44 6.33218 $w=5.08e-07 $l=2.7e-07 $layer=LI1_cond $X=2.51 $Y=1.295
+ $X2=2.51 $Y2=1.025
r67 37 44 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=0.9 $X2=2.51
+ $Y2=0.9
r68 33 35 37.8976 $w=2.58e-07 $l=8.55e-07 $layer=LI1_cond $X=2.035 $Y=2.04
+ $X2=2.035 $Y2=2.895
r69 31 45 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.035 $Y=1.81
+ $X2=2.51 $Y2=1.81
r70 31 33 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=2.035 $Y=1.895
+ $X2=2.035 $Y2=2.04
r71 27 51 0.475901 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=0.775
+ $X2=2.035 $Y2=0.9
r72 27 29 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=2.035 $Y=0.775
+ $X2=2.035 $Y2=0.44
r73 25 31 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.905 $Y=1.81
+ $X2=2.035 $Y2=1.81
r74 25 26 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.905 $Y=1.81
+ $X2=1.305 $Y2=1.81
r75 23 51 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.905 $Y=0.9
+ $X2=2.035 $Y2=0.9
r76 23 24 27.6586 $w=2.48e-07 $l=6e-07 $layer=LI1_cond $X=1.905 $Y=0.9 $X2=1.305
+ $Y2=0.9
r77 19 21 37.8976 $w=2.58e-07 $l=8.55e-07 $layer=LI1_cond $X=1.175 $Y=2.04
+ $X2=1.175 $Y2=2.895
r78 17 26 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.175 $Y=1.895
+ $X2=1.305 $Y2=1.81
r79 17 19 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.175 $Y=1.895
+ $X2=1.175 $Y2=2.04
r80 13 24 6.8199 $w=2.5e-07 $l=1.82071e-07 $layer=LI1_cond $X=1.175 $Y=0.775
+ $X2=1.305 $Y2=0.9
r81 13 15 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.175 $Y=0.775
+ $X2=1.175 $Y2=0.44
r82 4 35 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.835 $X2=2.03 $Y2=2.895
r83 4 33 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=1.835 $X2=2.03 $Y2=2.04
r84 3 21 400 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.895
r85 3 19 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.04
r86 2 29 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.035 $Y2=0.44
r87 1 15 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.175 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_4%VGND 1 2 3 12 16 18 20 23 24 25 27 36 41 45
r44 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r45 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r47 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 36 44 4.09394 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.607
+ $Y2=0
r49 36 38 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.335 $Y=0 $X2=2.16
+ $Y2=0
r50 35 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 32 41 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.692
+ $Y2=0
r53 32 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.2
+ $Y2=0
r54 30 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r55 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r56 27 41 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.692
+ $Y2=0
r57 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.24
+ $Y2=0
r58 25 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r59 25 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r60 23 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.2
+ $Y2=0
r61 23 24 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.602
+ $Y2=0
r62 22 38 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.73 $Y=0 $X2=2.16
+ $Y2=0
r63 22 24 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.73 $Y=0 $X2=1.602
+ $Y2=0
r64 18 44 3.26612 $w=2.8e-07 $l=1.69245e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.607 $Y2=0
r65 18 20 14.6113 $w=2.78e-07 $l=3.55e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0.44
r66 14 24 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.602 $Y2=0
r67 14 16 16.0438 $w=2.53e-07 $l=3.55e-07 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.602 $Y2=0.44
r68 10 41 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0
r69 10 12 14.877 $w=2.73e-07 $l=3.55e-07 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0.44
r70 3 20 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.465 $Y2=0.44
r71 2 16 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.235 $X2=1.605 $Y2=0.44
r72 1 12 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.44
.ends

