* File: sky130_fd_sc_lp__o21ai_1.spice
* Created: Wed Sep  2 10:15:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ai_1.pex.spice"
.subckt sky130_fd_sc_lp__o21ai_1  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A1_M1003_g N_A_29_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1596 AS=0.2226 PD=1.22 PS=2.21 NRD=4.284 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1000 N_A_29_47#_M1000_d N_A2_M1000_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1596 PD=1.12 PS=1.22 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_B1_M1005_g N_A_29_47#_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 A_112_367# N_A1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A2_M1001_g A_112_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2835
+ AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2835 PD=3.05 PS=1.71 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.2895 P=8.33
*
.include "sky130_fd_sc_lp__o21ai_1.pxi.spice"
*
.ends
*
*
