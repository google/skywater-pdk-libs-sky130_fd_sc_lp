* File: sky130_fd_sc_lp__and2_lp.pex.spice
* Created: Wed Sep  2 09:30:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2_LP%B 3 7 11 18 19 21 23 25 34
r37 23 25 8.56892 $w=6.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.815
+ $X2=1.2 $Y2=1.815
r38 23 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.72
+ $Y=1.645 $X2=0.72 $Y2=1.645
r39 21 23 8.56892 $w=6.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.815
+ $X2=0.72 $Y2=1.815
r40 18 34 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.72 $Y=2 $X2=0.72
+ $Y2=1.645
r41 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.72 $Y=2.075
+ $X2=0.99 $Y2=2.075
r42 15 18 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.63 $Y=2.075 $X2=0.72
+ $Y2=2.075
r43 14 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.48
+ $X2=0.72 $Y2=1.645
r44 9 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.99 $Y=2.15 $X2=0.99
+ $Y2=2.075
r45 9 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.99 $Y=2.15 $X2=0.99
+ $Y2=2.55
r46 7 14 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.81 $Y=1.08 $X2=0.81
+ $Y2=1.48
r47 1 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.63 $Y=2.15 $X2=0.63
+ $Y2=2.075
r48 1 3 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.63 $Y=2.15 $X2=0.63
+ $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP%A 1 3 5 6 8 9 12 13 15 19 21 22 23 27
c59 23 0 1.5113e-19 $X=1.68 $Y=0.555
c60 5 0 1.00686e-19 $X=1.42 $Y=2.08
r61 27 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=0.515
+ $X2=1.68 $Y2=0.68
r62 23 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=0.515 $X2=1.68 $Y2=0.515
r63 22 23 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.515
+ $X2=1.68 $Y2=0.515
r64 18 19 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.42 $Y=1.475
+ $X2=1.71 $Y2=1.475
r65 16 18 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.2 $Y=1.475
+ $X2=1.42 $Y2=1.475
r66 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.78 $Y=2.23
+ $X2=1.78 $Y2=2.55
r67 12 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.71 $Y=1.4 $X2=1.71
+ $Y2=1.475
r68 12 30 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=1.71 $Y=1.4 $X2=1.71
+ $Y2=0.68
r69 10 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.495 $Y=2.155
+ $X2=1.42 $Y2=2.155
r70 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.705 $Y=2.155
+ $X2=1.78 $Y2=2.23
r71 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.705 $Y=2.155
+ $X2=1.495 $Y2=2.155
r72 6 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.42 $Y=2.23 $X2=1.42
+ $Y2=2.155
r73 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.42 $Y=2.23 $X2=1.42
+ $Y2=2.55
r74 5 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.42 $Y=2.08 $X2=1.42
+ $Y2=2.155
r75 4 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.42 $Y=1.55 $X2=1.42
+ $Y2=1.475
r76 4 5 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.42 $Y=1.55 $X2=1.42
+ $Y2=2.08
r77 1 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.2 $Y=1.4 $X2=1.2
+ $Y2=1.475
r78 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.2 $Y=1.4 $X2=1.2
+ $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP%A_213_468# 1 2 9 13 17 21 24 25 32 38 40 45
c77 40 0 1.00686e-19 $X=2.19 $Y=1.235
c78 13 0 1.5113e-19 $X=2.395 $Y=0.67
r79 44 45 15.7369 $w=5.36e-07 $l=1.75e-07 $layer=POLY_cond $X=2.395 $Y=1.405
+ $X2=2.57 $Y2=1.405
r80 43 44 16.6362 $w=5.36e-07 $l=1.85e-07 $layer=POLY_cond $X=2.21 $Y=1.405
+ $X2=2.395 $Y2=1.405
r81 41 43 1.79851 $w=5.36e-07 $l=2e-08 $layer=POLY_cond $X=2.19 $Y=1.405
+ $X2=2.21 $Y2=1.405
r82 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.19
+ $Y=1.235 $X2=2.19 $Y2=1.235
r83 37 38 7.19996 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=1.08
+ $X2=1.655 $Y2=1.08
r84 35 37 4.03026 $w=4.58e-07 $l=1.55e-07 $layer=LI1_cond $X=1.415 $Y=1.08
+ $X2=1.57 $Y2=1.08
r85 30 32 9.49062 $w=4.58e-07 $l=3.65e-07 $layer=LI1_cond $X=1.205 $Y=2.55
+ $X2=1.57 $Y2=2.55
r86 25 40 4.85386 $w=1.7e-07 $l=1.81659e-07 $layer=LI1_cond $X=2.025 $Y=1.225
+ $X2=2.19 $Y2=1.19
r87 25 38 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.025 $Y=1.225
+ $X2=1.655 $Y2=1.225
r88 24 32 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.57 $Y=2.32 $X2=1.57
+ $Y2=2.55
r89 23 37 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.57 $Y=1.31 $X2=1.57
+ $Y2=1.08
r90 23 24 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.57 $Y=1.31
+ $X2=1.57 $Y2=2.32
r91 19 45 19.334 $w=5.36e-07 $l=4.29244e-07 $layer=POLY_cond $X=2.785 $Y=1.07
+ $X2=2.57 $Y2=1.405
r92 19 21 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.785 $Y=1.07
+ $X2=2.785 $Y2=0.67
r93 15 45 33.1734 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.57 $Y=1.74
+ $X2=2.57 $Y2=1.405
r94 15 17 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.57 $Y=1.74 $X2=2.57
+ $Y2=2.55
r95 11 44 33.1734 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.395 $Y=1.07
+ $X2=2.395 $Y2=1.405
r96 11 13 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.395 $Y=1.07
+ $X2=2.395 $Y2=0.67
r97 7 43 33.1734 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.21 $Y=1.74
+ $X2=2.21 $Y2=1.405
r98 7 9 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.21 $Y=1.74 $X2=2.21
+ $Y2=2.55
r99 2 30 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=2.34 $X2=1.205 $Y2=2.55
r100 1 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.275
+ $Y=0.87 $X2=1.415 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP%VPWR 1 2 7 9 13 16 17 18 31 32
r36 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 28 31 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r40 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 23 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 22 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r43 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 20 35 4.50438 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=0.58 $Y=3.33 $X2=0.29
+ $Y2=3.33
r45 20 22 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 18 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 18 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 18 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 16 25 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=3.33 $X2=1.68
+ $Y2=3.33
r51 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=1.995 $Y2=3.33
r52 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=3.245
+ $X2=1.995 $Y2=3.33
r53 11 13 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.995 $Y=3.245
+ $X2=1.995 $Y2=2.55
r54 7 35 3.26179 $w=3.3e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.415 $Y=3.245
+ $X2=0.29 $Y2=3.33
r55 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.415 $Y=3.245
+ $X2=0.415 $Y2=2.55
r56 2 13 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=2.34 $X2=1.995 $Y2=2.55
r57 1 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.27
+ $Y=2.34 $X2=0.415 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP%X 1 2 7 8 9 10 11 12 13
c14 7 0 6.97414e-20 $X=3.12 $Y=0.555
r15 13 57 3.79039 $w=7.08e-07 $l=2.25e-07 $layer=LI1_cond $X=2.88 $Y=2.775
+ $X2=2.88 $Y2=2.55
r16 12 57 2.4427 $w=7.08e-07 $l=1.45e-07 $layer=LI1_cond $X=2.88 $Y=2.405
+ $X2=2.88 $Y2=2.55
r17 11 12 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=2.035
+ $X2=2.88 $Y2=2.405
r18 10 11 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=2.035
r19 9 10 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=1.295
+ $X2=2.88 $Y2=1.665
r20 8 9 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=0.925 $X2=2.88
+ $Y2=1.295
r21 8 40 4.29577 $w=7.08e-07 $l=2.55e-07 $layer=LI1_cond $X=2.88 $Y=0.925
+ $X2=2.88 $Y2=0.67
r22 7 40 1.93731 $w=7.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.88 $Y=0.555
+ $X2=2.88 $Y2=0.67
r23 2 57 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=2.34 $X2=2.785 $Y2=2.55
r24 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.86
+ $Y=0.46 $X2=3 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LP__AND2_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r36 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r37 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r38 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r39 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.18
+ $Y2=0
r41 27 29 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=3.12
+ $Y2=0
r42 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.595
+ $Y2=0
r43 23 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.76 $Y=0 $X2=1.68
+ $Y2=0
r44 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=2.18
+ $Y2=0
r45 22 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=1.68
+ $Y2=0
r46 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.595
+ $Y2=0
r49 17 19 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.24
+ $Y2=0
r50 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r51 15 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r52 15 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0
r54 11 13 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0.67
r55 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0.085
+ $X2=0.595 $Y2=0
r56 7 9 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=0.595 $Y=0.085
+ $X2=0.595 $Y2=1.08
r57 2 13 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.035
+ $Y=0.46 $X2=2.18 $Y2=0.67
r58 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.45
+ $Y=0.87 $X2=0.595 $Y2=1.08
.ends

