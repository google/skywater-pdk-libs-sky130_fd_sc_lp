* File: sky130_fd_sc_lp__bufinv_8.pxi.spice
* Created: Fri Aug 28 10:11:30 2020
* 
x_PM_SKY130_FD_SC_LP__BUFINV_8%A_82_23# N_A_82_23#_M1002_d N_A_82_23#_M1008_d
+ N_A_82_23#_M1001_s N_A_82_23#_M1010_s N_A_82_23#_M1004_g N_A_82_23#_M1000_g
+ N_A_82_23#_M1005_g N_A_82_23#_M1003_g N_A_82_23#_M1007_g N_A_82_23#_M1006_g
+ N_A_82_23#_M1013_g N_A_82_23#_M1009_g N_A_82_23#_M1014_g N_A_82_23#_M1011_g
+ N_A_82_23#_M1016_g N_A_82_23#_M1017_g N_A_82_23#_M1022_g N_A_82_23#_M1019_g
+ N_A_82_23#_M1023_g N_A_82_23#_M1020_g N_A_82_23#_c_169_p N_A_82_23#_c_119_n
+ N_A_82_23#_c_120_n N_A_82_23#_c_121_n N_A_82_23#_c_122_n N_A_82_23#_c_137_n
+ N_A_82_23#_c_123_n N_A_82_23#_c_138_n N_A_82_23#_c_181_p N_A_82_23#_c_259_p
+ N_A_82_23#_c_124_n N_A_82_23#_c_125_n N_A_82_23#_c_139_n N_A_82_23#_c_126_n
+ PM_SKY130_FD_SC_LP__BUFINV_8%A_82_23#
x_PM_SKY130_FD_SC_LP__BUFINV_8%A_876_23# N_A_876_23#_M1018_d N_A_876_23#_M1012_d
+ N_A_876_23#_M1002_g N_A_876_23#_M1001_g N_A_876_23#_M1008_g
+ N_A_876_23#_M1010_g N_A_876_23#_M1015_g N_A_876_23#_M1021_g
+ N_A_876_23#_c_275_n N_A_876_23#_c_276_n N_A_876_23#_c_277_n
+ N_A_876_23#_c_278_n N_A_876_23#_c_344_p N_A_876_23#_c_308_p
+ N_A_876_23#_c_325_p N_A_876_23#_c_279_n N_A_876_23#_c_286_n
+ N_A_876_23#_c_287_n N_A_876_23#_c_280_n N_A_876_23#_c_281_n
+ PM_SKY130_FD_SC_LP__BUFINV_8%A_876_23#
x_PM_SKY130_FD_SC_LP__BUFINV_8%A N_A_M1018_g N_A_M1012_g A A N_A_c_364_n
+ N_A_c_365_n PM_SKY130_FD_SC_LP__BUFINV_8%A
x_PM_SKY130_FD_SC_LP__BUFINV_8%VPWR N_VPWR_M1000_s N_VPWR_M1003_s N_VPWR_M1009_s
+ N_VPWR_M1017_s N_VPWR_M1020_s N_VPWR_M1001_d N_VPWR_M1021_d N_VPWR_c_392_n
+ N_VPWR_c_393_n N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n
+ N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n
+ N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n
+ VPWR N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_391_n N_VPWR_c_411_n
+ N_VPWR_c_412_n N_VPWR_c_413_n PM_SKY130_FD_SC_LP__BUFINV_8%VPWR
x_PM_SKY130_FD_SC_LP__BUFINV_8%Y N_Y_M1004_s N_Y_M1007_s N_Y_M1014_s N_Y_M1022_s
+ N_Y_M1000_d N_Y_M1006_d N_Y_M1011_d N_Y_M1019_d N_Y_c_574_p N_Y_c_492_n
+ N_Y_c_552_n N_Y_c_493_n N_Y_c_499_n N_Y_c_575_p N_Y_c_556_n N_Y_c_494_n
+ N_Y_c_500_n N_Y_c_576_p N_Y_c_560_n N_Y_c_495_n N_Y_c_501_n N_Y_c_573_p
+ N_Y_c_564_n N_Y_c_496_n N_Y_c_502_n N_Y_c_497_n N_Y_c_503_n Y Y
+ PM_SKY130_FD_SC_LP__BUFINV_8%Y
x_PM_SKY130_FD_SC_LP__BUFINV_8%VGND N_VGND_M1004_d N_VGND_M1005_d N_VGND_M1013_d
+ N_VGND_M1016_d N_VGND_M1023_d N_VGND_M1002_s N_VGND_M1015_s N_VGND_c_585_n
+ N_VGND_c_586_n N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n
+ N_VGND_c_591_n N_VGND_c_592_n N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n
+ N_VGND_c_596_n N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n N_VGND_c_600_n
+ VGND N_VGND_c_601_n N_VGND_c_602_n N_VGND_c_603_n N_VGND_c_604_n
+ N_VGND_c_605_n N_VGND_c_606_n PM_SKY130_FD_SC_LP__BUFINV_8%VGND
cc_1 VNB N_A_82_23#_M1004_g 0.0288076f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.665
cc_2 VNB N_A_82_23#_M1005_g 0.0215624f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.665
cc_3 VNB N_A_82_23#_M1007_g 0.0215892f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.665
cc_4 VNB N_A_82_23#_M1013_g 0.021612f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=0.665
cc_5 VNB N_A_82_23#_M1014_g 0.021612f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=0.665
cc_6 VNB N_A_82_23#_M1016_g 0.021612f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=0.665
cc_7 VNB N_A_82_23#_M1022_g 0.021612f $X=-0.19 $Y=-0.245 $X2=3.065 $Y2=0.665
cc_8 VNB N_A_82_23#_M1023_g 0.0277989f $X=-0.19 $Y=-0.245 $X2=3.495 $Y2=0.665
cc_9 VNB N_A_82_23#_c_119_n 0.0382211f $X=-0.19 $Y=-0.245 $X2=3.87 $Y2=1.49
cc_10 VNB N_A_82_23#_c_120_n 0.00839373f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=0.48
cc_11 VNB N_A_82_23#_c_121_n 0.00285707f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=1.395
cc_12 VNB N_A_82_23#_c_122_n 0.00128445f $X=-0.19 $Y=-0.245 $X2=4.125 $Y2=1.755
cc_13 VNB N_A_82_23#_c_123_n 0.00577664f $X=-0.19 $Y=-0.245 $X2=5.005 $Y2=1.14
cc_14 VNB N_A_82_23#_c_124_n 0.00402709f $X=-0.19 $Y=-0.245 $X2=4.182 $Y2=1.14
cc_15 VNB N_A_82_23#_c_125_n 0.00135588f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=1.49
cc_16 VNB N_A_82_23#_c_126_n 0.136968f $X=-0.19 $Y=-0.245 $X2=3.57 $Y2=1.49
cc_17 VNB N_A_876_23#_M1002_g 0.0266395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_876_23#_M1008_g 0.0213871f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.655
cc_19 VNB N_A_876_23#_M1015_g 0.0215864f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.655
cc_20 VNB N_A_876_23#_c_275_n 0.00126482f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.665
cc_21 VNB N_A_876_23#_c_276_n 0.00228919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_876_23#_c_277_n 4.22924e-19 $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.465
cc_23 VNB N_A_876_23#_c_278_n 0.00753526f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.465
cc_24 VNB N_A_876_23#_c_279_n 0.0235964f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.655
cc_25 VNB N_A_876_23#_c_280_n 0.00119098f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=0.665
cc_26 VNB N_A_876_23#_c_281_n 0.0504698f $X=-0.19 $Y=-0.245 $X2=3.065 $Y2=0.665
cc_27 VNB N_A_M1012_g 0.00722944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB A 0.0204051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_c_364_n 0.0376492f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.325
cc_30 VNB N_A_c_365_n 0.0232711f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.665
cc_31 VNB N_VPWR_c_391_n 0.263193f $X=-0.19 $Y=-0.245 $X2=4.207 $Y2=2.05
cc_32 VNB N_Y_c_492_n 0.0288682f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=1.325
cc_33 VNB N_Y_c_493_n 0.00243905f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=2.465
cc_34 VNB N_Y_c_494_n 0.00240399f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.655
cc_35 VNB N_Y_c_495_n 0.00625533f $X=-0.19 $Y=-0.245 $X2=3.065 $Y2=0.665
cc_36 VNB N_Y_c_496_n 0.00210048f $X=-0.19 $Y=-0.245 $X2=4.03 $Y2=1.49
cc_37 VNB N_Y_c_497_n 0.00210048f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.49
cc_38 VNB N_VGND_c_585_n 0.0112246f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.665
cc_39 VNB N_VGND_c_586_n 0.033976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_587_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_588_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_589_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_590_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=0.665
cc_44 VNB N_VGND_c_591_n 0.0114389f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.465
cc_45 VNB N_VGND_c_592_n 0.0166301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_593_n 5.00113e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_594_n 6.09197e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_595_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=0.665
cc_49 VNB N_VGND_c_596_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_597_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=2.465
cc_51 VNB N_VGND_c_598_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=2.465
cc_52 VNB N_VGND_c_599_n 0.0166024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_600_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=3.065 $Y2=1.325
cc_54 VNB N_VGND_c_601_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=3.495 $Y2=2.465
cc_55 VNB N_VGND_c_602_n 0.01589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_603_n 0.315897f $X=-0.19 $Y=-0.245 $X2=3.87 $Y2=1.49
cc_57 VNB N_VGND_c_604_n 0.00538573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_605_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=4.125 $Y2=1.585
cc_59 VNB N_VGND_c_606_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=4.207 $Y2=2.05
cc_60 VPB N_A_82_23#_M1000_g 0.0236063f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_61 VPB N_A_82_23#_M1003_g 0.0190127f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=2.465
cc_62 VPB N_A_82_23#_M1006_g 0.0190396f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=2.465
cc_63 VPB N_A_82_23#_M1009_g 0.0190623f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.465
cc_64 VPB N_A_82_23#_M1011_g 0.0190623f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=2.465
cc_65 VPB N_A_82_23#_M1017_g 0.0190623f $X=-0.19 $Y=1.655 $X2=2.635 $Y2=2.465
cc_66 VPB N_A_82_23#_M1019_g 0.0190623f $X=-0.19 $Y=1.655 $X2=3.065 $Y2=2.465
cc_67 VPB N_A_82_23#_M1020_g 0.0242057f $X=-0.19 $Y=1.655 $X2=3.495 $Y2=2.465
cc_68 VPB N_A_82_23#_c_119_n 0.0159998f $X=-0.19 $Y=1.655 $X2=3.87 $Y2=1.49
cc_69 VPB N_A_82_23#_c_122_n 0.00218608f $X=-0.19 $Y=1.655 $X2=4.125 $Y2=1.755
cc_70 VPB N_A_82_23#_c_137_n 0.0117115f $X=-0.19 $Y=1.655 $X2=4.24 $Y2=2.05
cc_71 VPB N_A_82_23#_c_138_n 0.00471999f $X=-0.19 $Y=1.655 $X2=4.97 $Y2=1.84
cc_72 VPB N_A_82_23#_c_139_n 0.00444587f $X=-0.19 $Y=1.655 $X2=4.207 $Y2=1.84
cc_73 VPB N_A_82_23#_c_126_n 0.0168787f $X=-0.19 $Y=1.655 $X2=3.57 $Y2=1.49
cc_74 VPB N_A_876_23#_M1001_g 0.0233678f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.325
cc_75 VPB N_A_876_23#_M1010_g 0.0190365f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.325
cc_76 VPB N_A_876_23#_M1021_g 0.0188007f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.325
cc_77 VPB N_A_876_23#_c_277_n 0.00121394f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.465
cc_78 VPB N_A_876_23#_c_286_n 0.00755006f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=2.465
cc_79 VPB N_A_876_23#_c_287_n 0.0346949f $X=-0.19 $Y=1.655 $X2=2.635 $Y2=1.325
cc_80 VPB N_A_876_23#_c_281_n 0.00467327f $X=-0.19 $Y=1.655 $X2=3.065 $Y2=0.665
cc_81 VPB N_A_M1012_g 0.0251806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB A 0.01001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_392_n 0.0111987f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=0.665
cc_84 VPB N_VPWR_c_393_n 0.0431542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_394_n 0.00400996f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.665
cc_86 VPB N_VPWR_c_395_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_396_n 0.00400996f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.465
cc_88 VPB N_VPWR_c_397_n 0.0166954f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=0.665
cc_89 VPB N_VPWR_c_398_n 0.0153363f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=2.465
cc_90 VPB N_VPWR_c_399_n 0.0184035f $X=-0.19 $Y=1.655 $X2=2.635 $Y2=0.665
cc_91 VPB N_VPWR_c_400_n 0.00402346f $X=-0.19 $Y=1.655 $X2=2.635 $Y2=2.465
cc_92 VPB N_VPWR_c_401_n 4.05231e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_402_n 0.0166954f $X=-0.19 $Y=1.655 $X2=3.065 $Y2=2.465
cc_94 VPB N_VPWR_c_403_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_404_n 0.0166954f $X=-0.19 $Y=1.655 $X2=3.495 $Y2=0.665
cc_96 VPB N_VPWR_c_405_n 0.00497514f $X=-0.19 $Y=1.655 $X2=3.495 $Y2=0.665
cc_97 VPB N_VPWR_c_406_n 0.0166954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_407_n 0.00497514f $X=-0.19 $Y=1.655 $X2=3.495 $Y2=1.655
cc_99 VPB N_VPWR_c_408_n 0.0148515f $X=-0.19 $Y=1.655 $X2=4.182 $Y2=0.48
cc_100 VPB N_VPWR_c_409_n 0.0161053f $X=-0.19 $Y=1.655 $X2=4.207 $Y2=1.925
cc_101 VPB N_VPWR_c_391_n 0.0534491f $X=-0.19 $Y=1.655 $X2=4.207 $Y2=2.05
cc_102 VPB N_VPWR_c_411_n 0.00555219f $X=-0.19 $Y=1.655 $X2=4.335 $Y2=1.14
cc_103 VPB N_VPWR_c_412_n 0.00487897f $X=-0.19 $Y=1.655 $X2=5.082 $Y2=1.925
cc_104 VPB N_VPWR_c_413_n 0.00436868f $X=-0.19 $Y=1.655 $X2=5.082 $Y2=2.84
cc_105 VPB N_Y_c_492_n 0.0141773f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=1.325
cc_106 VPB N_Y_c_499_n 0.00243905f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=1.325
cc_107 VPB N_Y_c_500_n 0.00240399f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=2.465
cc_108 VPB N_Y_c_501_n 0.005492f $X=-0.19 $Y=1.655 $X2=3.065 $Y2=1.655
cc_109 VPB N_Y_c_502_n 0.00210048f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.49
cc_110 VPB N_Y_c_503_n 0.00210048f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=1.49
cc_111 N_A_82_23#_c_121_n N_A_876_23#_M1002_g 0.00502654f $X=4.12 $Y=1.395 $X2=0
+ $Y2=0
cc_112 N_A_82_23#_c_123_n N_A_876_23#_M1002_g 0.0157901f $X=5.005 $Y=1.14 $X2=0
+ $Y2=0
cc_113 N_A_82_23#_c_138_n N_A_876_23#_M1001_g 0.0150208f $X=4.97 $Y=1.84 $X2=0
+ $Y2=0
cc_114 N_A_82_23#_c_123_n N_A_876_23#_M1008_g 0.0138902f $X=5.005 $Y=1.14 $X2=0
+ $Y2=0
cc_115 N_A_82_23#_c_138_n N_A_876_23#_M1010_g 0.013934f $X=4.97 $Y=1.84 $X2=0
+ $Y2=0
cc_116 N_A_82_23#_c_123_n N_A_876_23#_M1015_g 0.00133885f $X=5.005 $Y=1.14 $X2=0
+ $Y2=0
cc_117 N_A_82_23#_c_138_n N_A_876_23#_M1021_g 7.75488e-19 $X=4.97 $Y=1.84 $X2=0
+ $Y2=0
cc_118 N_A_82_23#_c_123_n N_A_876_23#_c_275_n 0.0593531f $X=5.005 $Y=1.14 $X2=0
+ $Y2=0
cc_119 N_A_82_23#_c_138_n N_A_876_23#_c_275_n 0.0596739f $X=4.97 $Y=1.84 $X2=0
+ $Y2=0
cc_120 N_A_82_23#_c_125_n N_A_876_23#_c_275_n 0.016761f $X=4.12 $Y=1.49 $X2=0
+ $Y2=0
cc_121 N_A_82_23#_c_123_n N_A_876_23#_c_276_n 0.011281f $X=5.005 $Y=1.14 $X2=0
+ $Y2=0
cc_122 N_A_82_23#_c_138_n N_A_876_23#_c_277_n 0.008696f $X=4.97 $Y=1.84 $X2=0
+ $Y2=0
cc_123 N_A_82_23#_c_119_n N_A_876_23#_c_281_n 0.011358f $X=3.87 $Y=1.49 $X2=0
+ $Y2=0
cc_124 N_A_82_23#_c_122_n N_A_876_23#_c_281_n 0.00498787f $X=4.125 $Y=1.755
+ $X2=0 $Y2=0
cc_125 N_A_82_23#_c_123_n N_A_876_23#_c_281_n 0.00497162f $X=5.005 $Y=1.14 $X2=0
+ $Y2=0
cc_126 N_A_82_23#_c_138_n N_A_876_23#_c_281_n 0.00497162f $X=4.97 $Y=1.84 $X2=0
+ $Y2=0
cc_127 N_A_82_23#_c_125_n N_A_876_23#_c_281_n 7.83897e-19 $X=4.12 $Y=1.49 $X2=0
+ $Y2=0
cc_128 N_A_82_23#_c_138_n N_VPWR_M1001_d 0.00176461f $X=4.97 $Y=1.84 $X2=0 $Y2=0
cc_129 N_A_82_23#_M1000_g N_VPWR_c_393_n 0.00343774f $X=0.485 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_A_82_23#_M1003_g N_VPWR_c_394_n 0.0016342f $X=0.915 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_A_82_23#_M1006_g N_VPWR_c_394_n 0.0016342f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_A_82_23#_M1009_g N_VPWR_c_395_n 0.0016342f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_133 N_A_82_23#_M1011_g N_VPWR_c_395_n 0.0016342f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_82_23#_M1017_g N_VPWR_c_396_n 0.0016342f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_135 N_A_82_23#_M1019_g N_VPWR_c_396_n 0.0016342f $X=3.065 $Y=2.465 $X2=0
+ $Y2=0
cc_136 N_A_82_23#_M1019_g N_VPWR_c_397_n 0.00585385f $X=3.065 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A_82_23#_M1020_g N_VPWR_c_397_n 0.00585385f $X=3.495 $Y=2.465 $X2=0
+ $Y2=0
cc_138 N_A_82_23#_M1020_g N_VPWR_c_398_n 0.00512358f $X=3.495 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_82_23#_c_169_p N_VPWR_c_398_n 0.0153099f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_140 N_A_82_23#_c_119_n N_VPWR_c_398_n 0.00677564f $X=3.87 $Y=1.49 $X2=0 $Y2=0
cc_141 N_A_82_23#_c_137_n N_VPWR_c_398_n 0.0932477f $X=4.24 $Y=2.05 $X2=0 $Y2=0
cc_142 N_A_82_23#_c_139_n N_VPWR_c_398_n 0.00745028f $X=4.207 $Y=1.84 $X2=0
+ $Y2=0
cc_143 N_A_82_23#_c_137_n N_VPWR_c_399_n 0.0192838f $X=4.24 $Y=2.05 $X2=0 $Y2=0
cc_144 N_A_82_23#_c_138_n N_VPWR_c_400_n 0.0135055f $X=4.97 $Y=1.84 $X2=0 $Y2=0
cc_145 N_A_82_23#_M1000_g N_VPWR_c_402_n 0.00585385f $X=0.485 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_82_23#_M1003_g N_VPWR_c_402_n 0.00585385f $X=0.915 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_82_23#_M1006_g N_VPWR_c_404_n 0.00585385f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_82_23#_M1009_g N_VPWR_c_404_n 0.00585385f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_82_23#_M1011_g N_VPWR_c_406_n 0.00585385f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_82_23#_M1017_g N_VPWR_c_406_n 0.00585385f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_82_23#_c_181_p N_VPWR_c_408_n 0.0121496f $X=5.1 $Y=2.05 $X2=0 $Y2=0
cc_152 N_A_82_23#_M1001_s N_VPWR_c_391_n 0.00237481f $X=4.115 $Y=1.835 $X2=0
+ $Y2=0
cc_153 N_A_82_23#_M1010_s N_VPWR_c_391_n 0.00424013f $X=4.96 $Y=1.835 $X2=0
+ $Y2=0
cc_154 N_A_82_23#_M1000_g N_VPWR_c_391_n 0.0115721f $X=0.485 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_82_23#_M1003_g N_VPWR_c_391_n 0.0106302f $X=0.915 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_82_23#_M1006_g N_VPWR_c_391_n 0.0106302f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_82_23#_M1009_g N_VPWR_c_391_n 0.0106302f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A_82_23#_M1011_g N_VPWR_c_391_n 0.0106302f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A_82_23#_M1017_g N_VPWR_c_391_n 0.0106302f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_82_23#_M1019_g N_VPWR_c_391_n 0.0106302f $X=3.065 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_82_23#_M1020_g N_VPWR_c_391_n 0.0121372f $X=3.495 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_82_23#_c_137_n N_VPWR_c_391_n 0.0128214f $X=4.24 $Y=2.05 $X2=0 $Y2=0
cc_163 N_A_82_23#_c_181_p N_VPWR_c_391_n 0.00858612f $X=5.1 $Y=2.05 $X2=0 $Y2=0
cc_164 N_A_82_23#_M1004_g N_Y_c_492_n 0.0177921f $X=0.485 $Y=0.665 $X2=0 $Y2=0
cc_165 N_A_82_23#_M1000_g N_Y_c_492_n 0.0191524f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A_82_23#_M1005_g N_Y_c_492_n 0.00327942f $X=0.915 $Y=0.665 $X2=0 $Y2=0
cc_167 N_A_82_23#_M1003_g N_Y_c_492_n 0.00327942f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A_82_23#_c_169_p N_Y_c_492_n 0.0159839f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_169 N_A_82_23#_c_126_n N_Y_c_492_n 0.0343684f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_170 N_A_82_23#_M1005_g N_Y_c_493_n 0.0164752f $X=0.915 $Y=0.665 $X2=0 $Y2=0
cc_171 N_A_82_23#_M1007_g N_Y_c_493_n 0.0150449f $X=1.345 $Y=0.665 $X2=0 $Y2=0
cc_172 N_A_82_23#_c_169_p N_Y_c_493_n 0.0314731f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_173 N_A_82_23#_c_126_n N_Y_c_493_n 0.00243542f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_174 N_A_82_23#_M1003_g N_Y_c_499_n 0.0158126f $X=0.915 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A_82_23#_M1006_g N_Y_c_499_n 0.0141989f $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_82_23#_c_169_p N_Y_c_499_n 0.0314731f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_177 N_A_82_23#_c_126_n N_Y_c_499_n 0.00243542f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_178 N_A_82_23#_M1013_g N_Y_c_494_n 0.0150738f $X=1.775 $Y=0.665 $X2=0 $Y2=0
cc_179 N_A_82_23#_M1014_g N_Y_c_494_n 0.0150738f $X=2.205 $Y=0.665 $X2=0 $Y2=0
cc_180 N_A_82_23#_c_169_p N_Y_c_494_n 0.0420697f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_181 N_A_82_23#_c_126_n N_Y_c_494_n 0.00243542f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_182 N_A_82_23#_M1009_g N_Y_c_500_n 0.0141989f $X=1.775 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_82_23#_M1011_g N_Y_c_500_n 0.0141989f $X=2.205 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_82_23#_c_169_p N_Y_c_500_n 0.0420697f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_185 N_A_82_23#_c_126_n N_Y_c_500_n 0.00243542f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_186 N_A_82_23#_M1016_g N_Y_c_495_n 0.0150272f $X=2.635 $Y=0.665 $X2=0 $Y2=0
cc_187 N_A_82_23#_M1022_g N_Y_c_495_n 0.0147309f $X=3.065 $Y=0.665 $X2=0 $Y2=0
cc_188 N_A_82_23#_M1023_g N_Y_c_495_n 0.00254815f $X=3.495 $Y=0.665 $X2=0 $Y2=0
cc_189 N_A_82_23#_c_169_p N_Y_c_495_n 0.0632027f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_190 N_A_82_23#_c_124_n N_Y_c_495_n 0.00550621f $X=4.182 $Y=1.14 $X2=0 $Y2=0
cc_191 N_A_82_23#_c_126_n N_Y_c_495_n 0.00497162f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_192 N_A_82_23#_M1017_g N_Y_c_501_n 0.0141523f $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A_82_23#_M1019_g N_Y_c_501_n 0.0139969f $X=3.065 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A_82_23#_M1020_g N_Y_c_501_n 0.00147576f $X=3.495 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A_82_23#_c_169_p N_Y_c_501_n 0.0632027f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_196 N_A_82_23#_c_139_n N_Y_c_501_n 0.0030341f $X=4.207 $Y=1.84 $X2=0 $Y2=0
cc_197 N_A_82_23#_c_126_n N_Y_c_501_n 0.00497162f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_198 N_A_82_23#_c_169_p N_Y_c_496_n 0.021133f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_199 N_A_82_23#_c_126_n N_Y_c_496_n 0.00253619f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_200 N_A_82_23#_c_169_p N_Y_c_502_n 0.021133f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_201 N_A_82_23#_c_126_n N_Y_c_502_n 0.00253619f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_202 N_A_82_23#_c_169_p N_Y_c_497_n 0.021133f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_203 N_A_82_23#_c_126_n N_Y_c_497_n 0.00253619f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_204 N_A_82_23#_c_169_p N_Y_c_503_n 0.021133f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_205 N_A_82_23#_c_126_n N_Y_c_503_n 0.00253619f $X=3.57 $Y=1.49 $X2=0 $Y2=0
cc_206 N_A_82_23#_c_123_n N_VGND_M1002_s 0.00176461f $X=5.005 $Y=1.14 $X2=0
+ $Y2=0
cc_207 N_A_82_23#_M1004_g N_VGND_c_586_n 0.00430204f $X=0.485 $Y=0.665 $X2=0
+ $Y2=0
cc_208 N_A_82_23#_M1005_g N_VGND_c_587_n 0.00159325f $X=0.915 $Y=0.665 $X2=0
+ $Y2=0
cc_209 N_A_82_23#_M1007_g N_VGND_c_587_n 0.00159325f $X=1.345 $Y=0.665 $X2=0
+ $Y2=0
cc_210 N_A_82_23#_M1013_g N_VGND_c_588_n 0.00159325f $X=1.775 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_82_23#_M1014_g N_VGND_c_588_n 0.00159325f $X=2.205 $Y=0.665 $X2=0
+ $Y2=0
cc_212 N_A_82_23#_M1016_g N_VGND_c_589_n 0.00159325f $X=2.635 $Y=0.665 $X2=0
+ $Y2=0
cc_213 N_A_82_23#_M1022_g N_VGND_c_589_n 0.00159325f $X=3.065 $Y=0.665 $X2=0
+ $Y2=0
cc_214 N_A_82_23#_M1022_g N_VGND_c_590_n 0.00575161f $X=3.065 $Y=0.665 $X2=0
+ $Y2=0
cc_215 N_A_82_23#_M1023_g N_VGND_c_590_n 0.00575161f $X=3.495 $Y=0.665 $X2=0
+ $Y2=0
cc_216 N_A_82_23#_M1023_g N_VGND_c_591_n 0.00469772f $X=3.495 $Y=0.665 $X2=0
+ $Y2=0
cc_217 N_A_82_23#_c_169_p N_VGND_c_591_n 0.012215f $X=4.03 $Y=1.49 $X2=0 $Y2=0
cc_218 N_A_82_23#_c_119_n N_VGND_c_591_n 0.00621934f $X=3.87 $Y=1.49 $X2=0 $Y2=0
cc_219 N_A_82_23#_c_120_n N_VGND_c_591_n 0.0653608f $X=4.23 $Y=0.48 $X2=0 $Y2=0
cc_220 N_A_82_23#_c_124_n N_VGND_c_591_n 0.0013115f $X=4.182 $Y=1.14 $X2=0 $Y2=0
cc_221 N_A_82_23#_c_120_n N_VGND_c_592_n 0.0210232f $X=4.23 $Y=0.48 $X2=0 $Y2=0
cc_222 N_A_82_23#_c_123_n N_VGND_c_593_n 0.0170777f $X=5.005 $Y=1.14 $X2=0 $Y2=0
cc_223 N_A_82_23#_M1004_g N_VGND_c_595_n 0.00575161f $X=0.485 $Y=0.665 $X2=0
+ $Y2=0
cc_224 N_A_82_23#_M1005_g N_VGND_c_595_n 0.00575161f $X=0.915 $Y=0.665 $X2=0
+ $Y2=0
cc_225 N_A_82_23#_M1007_g N_VGND_c_597_n 0.00575161f $X=1.345 $Y=0.665 $X2=0
+ $Y2=0
cc_226 N_A_82_23#_M1013_g N_VGND_c_597_n 0.00575161f $X=1.775 $Y=0.665 $X2=0
+ $Y2=0
cc_227 N_A_82_23#_M1014_g N_VGND_c_599_n 0.00575161f $X=2.205 $Y=0.665 $X2=0
+ $Y2=0
cc_228 N_A_82_23#_M1016_g N_VGND_c_599_n 0.00575161f $X=2.635 $Y=0.665 $X2=0
+ $Y2=0
cc_229 N_A_82_23#_c_259_p N_VGND_c_601_n 0.0124525f $X=5.1 $Y=0.48 $X2=0 $Y2=0
cc_230 N_A_82_23#_M1002_d N_VGND_c_603_n 0.00381169f $X=4.105 $Y=0.245 $X2=0
+ $Y2=0
cc_231 N_A_82_23#_M1008_d N_VGND_c_603_n 0.00545212f $X=4.96 $Y=0.245 $X2=0
+ $Y2=0
cc_232 N_A_82_23#_M1004_g N_VGND_c_603_n 0.0115696f $X=0.485 $Y=0.665 $X2=0
+ $Y2=0
cc_233 N_A_82_23#_M1005_g N_VGND_c_603_n 0.0105815f $X=0.915 $Y=0.665 $X2=0
+ $Y2=0
cc_234 N_A_82_23#_M1007_g N_VGND_c_603_n 0.0105815f $X=1.345 $Y=0.665 $X2=0
+ $Y2=0
cc_235 N_A_82_23#_M1013_g N_VGND_c_603_n 0.0105815f $X=1.775 $Y=0.665 $X2=0
+ $Y2=0
cc_236 N_A_82_23#_M1014_g N_VGND_c_603_n 0.0105815f $X=2.205 $Y=0.665 $X2=0
+ $Y2=0
cc_237 N_A_82_23#_M1016_g N_VGND_c_603_n 0.0105815f $X=2.635 $Y=0.665 $X2=0
+ $Y2=0
cc_238 N_A_82_23#_M1022_g N_VGND_c_603_n 0.0105815f $X=3.065 $Y=0.665 $X2=0
+ $Y2=0
cc_239 N_A_82_23#_M1023_g N_VGND_c_603_n 0.0119274f $X=3.495 $Y=0.665 $X2=0
+ $Y2=0
cc_240 N_A_82_23#_c_120_n N_VGND_c_603_n 0.0117799f $X=4.23 $Y=0.48 $X2=0 $Y2=0
cc_241 N_A_82_23#_c_259_p N_VGND_c_603_n 0.00730901f $X=5.1 $Y=0.48 $X2=0 $Y2=0
cc_242 N_A_876_23#_M1021_g N_A_M1012_g 0.0281514f $X=5.315 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A_876_23#_c_277_n N_A_M1012_g 0.00513935f $X=5.47 $Y=1.97 $X2=0 $Y2=0
cc_244 N_A_876_23#_c_308_p N_A_M1012_g 0.0146839f $X=5.865 $Y=2.055 $X2=0 $Y2=0
cc_245 N_A_876_23#_M1015_g A 5.14553e-19 $X=5.315 $Y=0.665 $X2=0 $Y2=0
cc_246 N_A_876_23#_c_276_n A 0.0127034f $X=5.47 $Y=1.395 $X2=0 $Y2=0
cc_247 N_A_876_23#_c_277_n A 0.014769f $X=5.47 $Y=1.97 $X2=0 $Y2=0
cc_248 N_A_876_23#_c_278_n A 0.0314086f $X=5.865 $Y=0.955 $X2=0 $Y2=0
cc_249 N_A_876_23#_c_308_p A 0.00721495f $X=5.865 $Y=2.055 $X2=0 $Y2=0
cc_250 N_A_876_23#_c_286_n A 0.0231742f $X=5.995 $Y=2.14 $X2=0 $Y2=0
cc_251 N_A_876_23#_c_280_n A 0.0146216f $X=5.47 $Y=1.49 $X2=0 $Y2=0
cc_252 N_A_876_23#_c_278_n N_A_c_364_n 0.00103212f $X=5.865 $Y=0.955 $X2=0 $Y2=0
cc_253 N_A_876_23#_c_286_n N_A_c_364_n 5.78882e-19 $X=5.995 $Y=2.14 $X2=0 $Y2=0
cc_254 N_A_876_23#_c_280_n N_A_c_364_n 0.0015461f $X=5.47 $Y=1.49 $X2=0 $Y2=0
cc_255 N_A_876_23#_c_281_n N_A_c_364_n 0.0281514f $X=5.315 $Y=1.49 $X2=0 $Y2=0
cc_256 N_A_876_23#_M1015_g N_A_c_365_n 0.0281514f $X=5.315 $Y=0.665 $X2=0 $Y2=0
cc_257 N_A_876_23#_c_276_n N_A_c_365_n 0.00507626f $X=5.47 $Y=1.395 $X2=0 $Y2=0
cc_258 N_A_876_23#_c_278_n N_A_c_365_n 0.0146839f $X=5.865 $Y=0.955 $X2=0 $Y2=0
cc_259 N_A_876_23#_c_277_n N_VPWR_M1021_d 0.00150539f $X=5.47 $Y=1.97 $X2=0
+ $Y2=0
cc_260 N_A_876_23#_c_308_p N_VPWR_M1021_d 0.00278079f $X=5.865 $Y=2.055 $X2=0
+ $Y2=0
cc_261 N_A_876_23#_c_325_p N_VPWR_M1021_d 0.00118409f $X=5.555 $Y=2.055 $X2=0
+ $Y2=0
cc_262 N_A_876_23#_M1001_g N_VPWR_c_398_n 0.00353963f $X=4.455 $Y=2.465 $X2=0
+ $Y2=0
cc_263 N_A_876_23#_M1001_g N_VPWR_c_399_n 0.00585385f $X=4.455 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A_876_23#_M1001_g N_VPWR_c_400_n 0.00170737f $X=4.455 $Y=2.465 $X2=0
+ $Y2=0
cc_265 N_A_876_23#_M1010_g N_VPWR_c_400_n 0.00158314f $X=4.885 $Y=2.465 $X2=0
+ $Y2=0
cc_266 N_A_876_23#_M1010_g N_VPWR_c_401_n 7.70828e-19 $X=4.885 $Y=2.465 $X2=0
+ $Y2=0
cc_267 N_A_876_23#_M1021_g N_VPWR_c_401_n 0.0142077f $X=5.315 $Y=2.465 $X2=0
+ $Y2=0
cc_268 N_A_876_23#_c_308_p N_VPWR_c_401_n 0.0064684f $X=5.865 $Y=2.055 $X2=0
+ $Y2=0
cc_269 N_A_876_23#_c_325_p N_VPWR_c_401_n 0.010031f $X=5.555 $Y=2.055 $X2=0
+ $Y2=0
cc_270 N_A_876_23#_M1010_g N_VPWR_c_408_n 0.00585385f $X=4.885 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_876_23#_M1021_g N_VPWR_c_408_n 0.00486043f $X=5.315 $Y=2.465 $X2=0
+ $Y2=0
cc_272 N_A_876_23#_c_287_n N_VPWR_c_409_n 0.0157867f $X=5.96 $Y=2.815 $X2=0
+ $Y2=0
cc_273 N_A_876_23#_M1012_d N_VPWR_c_391_n 0.00376532f $X=5.82 $Y=1.835 $X2=0
+ $Y2=0
cc_274 N_A_876_23#_M1001_g N_VPWR_c_391_n 0.0120435f $X=4.455 $Y=2.465 $X2=0
+ $Y2=0
cc_275 N_A_876_23#_M1010_g N_VPWR_c_391_n 0.0106302f $X=4.885 $Y=2.465 $X2=0
+ $Y2=0
cc_276 N_A_876_23#_M1021_g N_VPWR_c_391_n 0.00835506f $X=5.315 $Y=2.465 $X2=0
+ $Y2=0
cc_277 N_A_876_23#_c_287_n N_VPWR_c_391_n 0.00993371f $X=5.96 $Y=2.815 $X2=0
+ $Y2=0
cc_278 N_A_876_23#_c_276_n N_VGND_M1015_s 4.94306e-19 $X=5.47 $Y=1.395 $X2=0
+ $Y2=0
cc_279 N_A_876_23#_c_278_n N_VGND_M1015_s 0.00278079f $X=5.865 $Y=0.955 $X2=0
+ $Y2=0
cc_280 N_A_876_23#_c_344_p N_VGND_M1015_s 0.00119515f $X=5.555 $Y=0.955 $X2=0
+ $Y2=0
cc_281 N_A_876_23#_M1002_g N_VGND_c_591_n 0.00252213f $X=4.455 $Y=0.665 $X2=0
+ $Y2=0
cc_282 N_A_876_23#_M1002_g N_VGND_c_592_n 0.00477554f $X=4.455 $Y=0.665 $X2=0
+ $Y2=0
cc_283 N_A_876_23#_M1002_g N_VGND_c_593_n 0.0111654f $X=4.455 $Y=0.665 $X2=0
+ $Y2=0
cc_284 N_A_876_23#_M1008_g N_VGND_c_593_n 0.010557f $X=4.885 $Y=0.665 $X2=0
+ $Y2=0
cc_285 N_A_876_23#_M1015_g N_VGND_c_593_n 6.31723e-19 $X=5.315 $Y=0.665 $X2=0
+ $Y2=0
cc_286 N_A_876_23#_M1008_g N_VGND_c_594_n 5.79385e-19 $X=4.885 $Y=0.665 $X2=0
+ $Y2=0
cc_287 N_A_876_23#_M1015_g N_VGND_c_594_n 0.0104338f $X=5.315 $Y=0.665 $X2=0
+ $Y2=0
cc_288 N_A_876_23#_c_278_n N_VGND_c_594_n 0.0064684f $X=5.865 $Y=0.955 $X2=0
+ $Y2=0
cc_289 N_A_876_23#_c_344_p N_VGND_c_594_n 0.0101184f $X=5.555 $Y=0.955 $X2=0
+ $Y2=0
cc_290 N_A_876_23#_M1008_g N_VGND_c_601_n 0.00477554f $X=4.885 $Y=0.665 $X2=0
+ $Y2=0
cc_291 N_A_876_23#_M1015_g N_VGND_c_601_n 0.00477554f $X=5.315 $Y=0.665 $X2=0
+ $Y2=0
cc_292 N_A_876_23#_c_279_n N_VGND_c_602_n 0.0192173f $X=5.98 $Y=0.48 $X2=0 $Y2=0
cc_293 N_A_876_23#_M1018_d N_VGND_c_603_n 0.00389211f $X=5.82 $Y=0.245 $X2=0
+ $Y2=0
cc_294 N_A_876_23#_M1002_g N_VGND_c_603_n 0.00960399f $X=4.455 $Y=0.665 $X2=0
+ $Y2=0
cc_295 N_A_876_23#_M1008_g N_VGND_c_603_n 0.0083043f $X=4.885 $Y=0.665 $X2=0
+ $Y2=0
cc_296 N_A_876_23#_M1015_g N_VGND_c_603_n 0.0083043f $X=5.315 $Y=0.665 $X2=0
+ $Y2=0
cc_297 N_A_876_23#_c_279_n N_VGND_c_603_n 0.010808f $X=5.98 $Y=0.48 $X2=0 $Y2=0
cc_298 N_A_M1012_g N_VPWR_c_401_n 0.0158322f $X=5.745 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A_M1012_g N_VPWR_c_409_n 0.00486043f $X=5.745 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A_M1012_g N_VPWR_c_391_n 0.00937921f $X=5.745 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A_c_365_n N_VGND_c_594_n 0.0113834f $X=5.835 $Y=1.21 $X2=0 $Y2=0
cc_302 N_A_c_365_n N_VGND_c_602_n 0.00477554f $X=5.835 $Y=1.21 $X2=0 $Y2=0
cc_303 N_A_c_365_n N_VGND_c_603_n 0.0092553f $X=5.835 $Y=1.21 $X2=0 $Y2=0
cc_304 N_VPWR_c_391_n N_Y_M1000_d 0.00302344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_305 N_VPWR_c_391_n N_Y_M1006_d 0.00302344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_306 N_VPWR_c_391_n N_Y_M1011_d 0.00302344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_307 N_VPWR_c_391_n N_Y_M1019_d 0.00302344f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_M1000_s N_Y_c_492_n 0.00272521f $X=0.145 $Y=1.835 $X2=0 $Y2=0
cc_309 N_VPWR_c_393_n N_Y_c_492_n 0.0224079f $X=0.27 $Y=2.26 $X2=0 $Y2=0
cc_310 N_VPWR_c_402_n N_Y_c_552_n 0.0132609f $X=1 $Y=3.33 $X2=0 $Y2=0
cc_311 N_VPWR_c_391_n N_Y_c_552_n 0.00993371f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_312 N_VPWR_M1003_s N_Y_c_499_n 0.00176461f $X=0.99 $Y=1.835 $X2=0 $Y2=0
cc_313 N_VPWR_c_394_n N_Y_c_499_n 0.0135055f $X=1.13 $Y=2.26 $X2=0 $Y2=0
cc_314 N_VPWR_c_404_n N_Y_c_556_n 0.0132609f $X=1.86 $Y=3.33 $X2=0 $Y2=0
cc_315 N_VPWR_c_391_n N_Y_c_556_n 0.00993371f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_316 N_VPWR_M1009_s N_Y_c_500_n 0.00176461f $X=1.85 $Y=1.835 $X2=0 $Y2=0
cc_317 N_VPWR_c_395_n N_Y_c_500_n 0.0135055f $X=1.99 $Y=2.26 $X2=0 $Y2=0
cc_318 N_VPWR_c_406_n N_Y_c_560_n 0.0132609f $X=2.72 $Y=3.33 $X2=0 $Y2=0
cc_319 N_VPWR_c_391_n N_Y_c_560_n 0.00993371f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_M1017_s N_Y_c_501_n 0.00176461f $X=2.71 $Y=1.835 $X2=0 $Y2=0
cc_321 N_VPWR_c_396_n N_Y_c_501_n 0.0135055f $X=2.85 $Y=2.26 $X2=0 $Y2=0
cc_322 N_VPWR_c_397_n N_Y_c_564_n 0.0132609f $X=3.58 $Y=3.33 $X2=0 $Y2=0
cc_323 N_VPWR_c_391_n N_Y_c_564_n 0.00993371f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_324 N_Y_c_493_n N_VGND_M1005_d 0.00176461f $X=1.43 $Y=1.14 $X2=0 $Y2=0
cc_325 N_Y_c_494_n N_VGND_M1013_d 0.00176461f $X=2.29 $Y=1.14 $X2=0 $Y2=0
cc_326 N_Y_c_495_n N_VGND_M1016_d 0.00176461f $X=3.15 $Y=1.14 $X2=0 $Y2=0
cc_327 N_Y_c_492_n N_VGND_c_586_n 0.0249306f $X=0.7 $Y=1.925 $X2=0 $Y2=0
cc_328 N_Y_c_493_n N_VGND_c_587_n 0.0135055f $X=1.43 $Y=1.14 $X2=0 $Y2=0
cc_329 N_Y_c_494_n N_VGND_c_588_n 0.0135055f $X=2.29 $Y=1.14 $X2=0 $Y2=0
cc_330 N_Y_c_495_n N_VGND_c_589_n 0.0135055f $X=3.15 $Y=1.14 $X2=0 $Y2=0
cc_331 N_Y_c_573_p N_VGND_c_590_n 0.0149362f $X=3.28 $Y=0.48 $X2=0 $Y2=0
cc_332 N_Y_c_574_p N_VGND_c_595_n 0.0149362f $X=0.7 $Y=0.48 $X2=0 $Y2=0
cc_333 N_Y_c_575_p N_VGND_c_597_n 0.0149362f $X=1.56 $Y=0.48 $X2=0 $Y2=0
cc_334 N_Y_c_576_p N_VGND_c_599_n 0.0149362f $X=2.42 $Y=0.48 $X2=0 $Y2=0
cc_335 N_Y_M1004_s N_VGND_c_603_n 0.003017f $X=0.56 $Y=0.245 $X2=0 $Y2=0
cc_336 N_Y_M1007_s N_VGND_c_603_n 0.003017f $X=1.42 $Y=0.245 $X2=0 $Y2=0
cc_337 N_Y_M1014_s N_VGND_c_603_n 0.003017f $X=2.28 $Y=0.245 $X2=0 $Y2=0
cc_338 N_Y_M1022_s N_VGND_c_603_n 0.003017f $X=3.14 $Y=0.245 $X2=0 $Y2=0
cc_339 N_Y_c_574_p N_VGND_c_603_n 0.0100304f $X=0.7 $Y=0.48 $X2=0 $Y2=0
cc_340 N_Y_c_575_p N_VGND_c_603_n 0.0100304f $X=1.56 $Y=0.48 $X2=0 $Y2=0
cc_341 N_Y_c_576_p N_VGND_c_603_n 0.0100304f $X=2.42 $Y=0.48 $X2=0 $Y2=0
cc_342 N_Y_c_573_p N_VGND_c_603_n 0.0100304f $X=3.28 $Y=0.48 $X2=0 $Y2=0
