* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__maj3_m A B C VGND VNB VPB VPWR X
X0 a_34_57# C a_121_425# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_285_425# B a_34_57# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_34_57# B a_449_425# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_449_425# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_121_425# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_285_57# B a_34_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_34_57# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_34_57# C a_121_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR A a_285_425# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_34_57# B a_449_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_121_57# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND A a_285_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_449_57# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VGND a_34_57# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
