* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or2_lp A B VGND VNB VPB VPWR X
X0 a_484_114# a_196_114# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR A a_154_468# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND A a_118_114# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_435_490# a_196_114# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_118_114# A a_196_114# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_282_114# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_154_468# B a_196_114# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_196_114# B a_282_114# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_196_114# a_484_114# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_196_114# a_435_490# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
