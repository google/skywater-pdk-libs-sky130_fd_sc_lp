* File: sky130_fd_sc_lp__o311ai_m.pex.spice
* Created: Wed Sep  2 10:24:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311AI_M%A1 5 8 10 11 12 13 14 19 21
c36 21 0 1.9934e-19 $X=0.442 $Y=0.94
c37 12 0 6.45684e-20 $X=0.24 $Y=0.925
c38 11 0 2.20127e-20 $X=0.472 $Y=1.61
r39 19 21 47.6426 $w=4.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.442 $Y=1.105
+ $X2=0.442 $Y2=0.94
r40 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.37
+ $Y=1.105 $X2=0.37 $Y2=1.105
r41 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.305 $Y=1.295
+ $X2=0.305 $Y2=1.665
r42 13 20 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=0.305 $Y=1.295
+ $X2=0.305 $Y2=1.105
r43 12 20 6.91466 $w=2.98e-07 $l=1.8e-07 $layer=LI1_cond $X=0.305 $Y=0.925
+ $X2=0.305 $Y2=1.105
r44 10 11 45.8863 $w=4.75e-07 $l=1.5e-07 $layer=POLY_cond $X=0.472 $Y=1.46
+ $X2=0.472 $Y2=1.61
r45 8 11 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.665 $Y=2.225
+ $X2=0.665 $Y2=1.61
r46 5 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.605 $Y=0.62
+ $X2=0.605 $Y2=0.94
r47 1 19 8.43012 $w=4.75e-07 $l=7.2e-08 $layer=POLY_cond $X=0.442 $Y=1.177
+ $X2=0.442 $Y2=1.105
r48 1 10 33.1351 $w=4.75e-07 $l=2.83e-07 $layer=POLY_cond $X=0.442 $Y=1.177
+ $X2=0.442 $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_M%A2 4 7 10 11 12
c42 12 0 1.72357e-19 $X=0.72 $Y=2.775
c43 10 0 1.11965e-19 $X=1.03 $Y=1.515
c44 7 0 1.9934e-19 $X=1.035 $Y=0.62
r45 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=2.94 $X2=0.77 $Y2=2.94
r46 12 16 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=2.775
+ $X2=0.77 $Y2=2.94
r47 11 15 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.95 $Y=2.94 $X2=0.77
+ $Y2=2.94
r48 9 10 69.5192 $w=1.6e-07 $l=1.5e-07 $layer=POLY_cond $X=1.03 $Y=1.365
+ $X2=1.03 $Y2=1.515
r49 7 9 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=1.035 $Y=0.62
+ $X2=1.035 $Y2=1.365
r50 4 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.025 $Y=2.225
+ $X2=1.025 $Y2=1.515
r51 2 11 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.025 $Y=2.775
+ $X2=0.95 $Y2=2.94
r52 2 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.025 $Y=2.775
+ $X2=1.025 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_M%A3 4 9 11 12 14 15 16 22
c45 22 0 1.72357e-19 $X=1.505 $Y=2.94
c46 12 0 1.62223e-19 $X=1.405 $Y=1.905
r47 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.505
+ $Y=2.94 $X2=1.505 $Y2=2.94
r48 19 22 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.385 $Y=2.94
+ $X2=1.505 $Y2=2.94
r49 16 23 6.02022 $w=3.33e-07 $l=1.75e-07 $layer=LI1_cond $X=1.68 $Y=2.857
+ $X2=1.505 $Y2=2.857
r50 15 23 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=2.857
+ $X2=1.505 $Y2=2.857
r51 13 14 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.445 $Y=1.11
+ $X2=1.445 $Y2=1.26
r52 11 12 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.405 $Y=1.755
+ $X2=1.405 $Y2=1.905
r53 11 14 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.425 $Y=1.755
+ $X2=1.425 $Y2=1.26
r54 9 13 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.465 $Y=0.62
+ $X2=1.465 $Y2=1.11
r55 4 12 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.385 $Y=2.225
+ $X2=1.385 $Y2=1.905
r56 2 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=2.775
+ $X2=1.385 $Y2=2.94
r57 2 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.385 $Y=2.775
+ $X2=1.385 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_M%B1 3 7 9 10 11 16
c43 7 0 9.31808e-20 $X=1.895 $Y=0.62
r44 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.665
+ $X2=1.905 $Y2=1.83
r45 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.665
+ $X2=1.905 $Y2=1.5
r46 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.905
+ $Y=1.665 $X2=1.905 $Y2=1.665
r47 11 17 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=1.905 $Y2=1.665
r48 10 17 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.905 $Y2=1.665
r49 9 10 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.665 $X2=1.68
+ $Y2=1.665
r50 7 18 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=1.895 $Y=0.62
+ $X2=1.895 $Y2=1.5
r51 3 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.815 $Y=2.225
+ $X2=1.815 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_M%C1 3 6 9 10 12 13 14 15 20 21 22
r39 21 22 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.625 $Y=1.12
+ $X2=2.625 $Y2=1.055
r40 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.61
+ $Y=1.12 $X2=2.61 $Y2=1.12
r41 14 15 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.625 $Y=1.295
+ $X2=2.625 $Y2=1.665
r42 14 21 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=2.625 $Y=1.295
+ $X2=2.625 $Y2=1.12
r43 13 22 8.04083 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=2.625 $Y=0.925
+ $X2=2.625 $Y2=1.055
r44 11 20 35.3689 $w=4.45e-07 $l=2.83e-07 $layer=POLY_cond $X=2.552 $Y=1.403
+ $X2=2.552 $Y2=1.12
r45 11 12 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=2.552 $Y=1.403
+ $X2=2.552 $Y2=1.625
r46 10 20 1.87468 $w=4.45e-07 $l=1.5e-08 $layer=POLY_cond $X=2.552 $Y=1.105
+ $X2=2.552 $Y2=1.12
r47 9 10 44.9281 $w=4.45e-07 $l=1.5e-07 $layer=POLY_cond $X=2.477 $Y=0.955
+ $X2=2.477 $Y2=1.105
r48 6 12 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.405 $Y=2.225 $X2=2.405
+ $Y2=1.625
r49 3 9 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.255 $Y=0.62
+ $X2=2.255 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_M%VPWR 1 2 7 9 13 15 17 27 28 34
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.11 $Y2=3.33
r44 25 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r49 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 18 31 3.5042 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r51 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=2.11 $Y2=3.33
r53 17 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 15 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 15 21 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.11 $Y2=3.33
r57 11 13 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.11 $Y2=2.365
r58 7 31 3.33969 $w=1.9e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.212 $Y2=3.33
r59 7 9 55.7464 $w=1.88e-07 $l=9.55e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.33 $Y2=2.29
r60 2 13 600 $w=1.7e-07 $l=4.46654e-07 $layer=licon1_PDIFF $count=1 $X=1.89
+ $Y=2.015 $X2=2.11 $Y2=2.365
r61 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=2.015 $X2=0.34 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_M%Y 1 2 3 14 15 17 18 20 22 23 24 29 30 31 32
c77 15 0 1.62223e-19 $X=1.705 $Y=2.015
r78 31 32 12.5394 $w=3.38e-07 $l=2.85e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.32
r79 30 31 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=2.035
r80 29 30 12.5394 $w=3.38e-07 $l=2.85e-07 $layer=LI1_cond $X=0.72 $Y=1.38
+ $X2=0.72 $Y2=1.665
r81 24 27 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=2.62 $Y=2.015
+ $X2=2.62 $Y2=2.16
r82 23 29 47.8763 $w=3.38e-07 $l=1.37e-06 $layer=LI1_cond $X=2.175 $Y=1.295
+ $X2=0.805 $Y2=1.295
r83 22 32 24.8274 $w=3.38e-07 $l=6.9e-07 $layer=LI1_cond $X=1.495 $Y=2.405
+ $X2=0.805 $Y2=2.405
r84 18 20 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=2.345 $Y=0.555
+ $X2=2.47 $Y2=0.555
r85 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.26 $Y=1.21
+ $X2=2.175 $Y2=1.295
r86 16 18 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.26 $Y=0.66
+ $X2=2.345 $Y2=0.555
r87 16 17 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.26 $Y=0.66
+ $X2=2.26 $Y2=1.21
r88 14 24 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.515 $Y=2.015
+ $X2=2.62 $Y2=2.015
r89 14 15 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.515 $Y=2.015
+ $X2=1.705 $Y2=2.015
r90 11 22 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.6 $Y=2.32
+ $X2=1.495 $Y2=2.405
r91 11 13 8.45022 $w=2.08e-07 $l=1.6e-07 $layer=LI1_cond $X=1.6 $Y=2.32 $X2=1.6
+ $Y2=2.16
r92 10 15 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.6 $Y=2.1
+ $X2=1.705 $Y2=2.015
r93 10 13 3.16883 $w=2.08e-07 $l=6e-08 $layer=LI1_cond $X=1.6 $Y=2.1 $X2=1.6
+ $Y2=2.16
r94 3 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=2.015 $X2=2.62 $Y2=2.16
r95 2 13 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=2.015 $X2=1.6 $Y2=2.16
r96 1 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.33
+ $Y=0.41 $X2=2.47 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_M%VGND 1 2 7 9 13 15 17 27 28 34
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 25 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r41 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r42 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r43 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.25
+ $Y2=0
r44 22 24 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.68
+ $Y2=0
r45 21 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r46 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r47 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 18 31 4.53571 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.277
+ $Y2=0
r49 18 20 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.72
+ $Y2=0
r50 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=0 $X2=1.25
+ $Y2=0
r51 17 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.085 $Y=0 $X2=0.72
+ $Y2=0
r52 15 25 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r53 15 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r54 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=0.085
+ $X2=1.25 $Y2=0
r55 11 13 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.25 $Y=0.085
+ $X2=1.25 $Y2=0.555
r56 7 31 3.23047 $w=3.3e-07 $l=1.49579e-07 $layer=LI1_cond $X=0.39 $Y=0.085
+ $X2=0.277 $Y2=0
r57 7 9 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.39 $Y=0.085 $X2=0.39
+ $Y2=0.555
r58 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.11
+ $Y=0.41 $X2=1.25 $Y2=0.555
r59 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.265
+ $Y=0.41 $X2=0.39 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_M%A_136_82# 1 2 9 11 12 15
c20 15 0 2.49048e-19 $X=1.68 $Y=0.685
c21 12 0 2.20127e-20 $X=0.905 $Y=0.925
c22 11 0 4.73962e-20 $X=1.595 $Y=0.925
c23 9 0 5.58598e-19 $X=0.82 $Y=0.685
r24 13 15 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.69 $Y=0.84
+ $X2=1.69 $Y2=0.685
r25 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.595 $Y=0.925
+ $X2=1.69 $Y2=0.84
r26 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.595 $Y=0.925
+ $X2=0.905 $Y2=0.925
r27 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.82 $Y=0.84
+ $X2=0.905 $Y2=0.925
r28 7 9 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.82 $Y=0.84 $X2=0.82
+ $Y2=0.685
r29 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.41 $X2=1.68 $Y2=0.685
r30 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.68
+ $Y=0.41 $X2=0.82 $Y2=0.685
.ends

