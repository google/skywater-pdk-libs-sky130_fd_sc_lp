* File: sky130_fd_sc_lp__nand4b_2.pex.spice
* Created: Wed Sep  2 10:06:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4B_2%A_N 2 5 7 8 11 13 16 17
c36 17 0 1.00394e-19 $X=0.27 $Y=1.12
r37 16 18 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.327 $Y=1.12
+ $X2=0.327 $Y2=0.955
r38 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r39 13 17 0.608175 $w=5.88e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=1.33 $X2=0.27
+ $Y2=1.33
r40 9 11 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.8 $Y=1.625 $X2=0.8
+ $Y2=2.045
r41 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.725 $Y=1.55
+ $X2=0.8 $Y2=1.625
r42 7 8 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.725 $Y=1.55 $X2=0.55
+ $Y2=1.55
r43 5 18 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.475 $Y=0.465
+ $X2=0.475 $Y2=0.955
r44 2 8 36.6125 $w=1.5e-07 $l=2.57787e-07 $layer=POLY_cond $X=0.327 $Y=1.475
+ $X2=0.55 $Y2=1.55
r45 1 16 7.12377 $w=4.45e-07 $l=5.7e-08 $layer=POLY_cond $X=0.327 $Y=1.177
+ $X2=0.327 $Y2=1.12
r46 1 2 37.2436 $w=4.45e-07 $l=2.98e-07 $layer=POLY_cond $X=0.327 $Y=1.177
+ $X2=0.327 $Y2=1.475
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%A_27_51# 1 2 9 13 17 21 25 27 28 30 32 35
+ 41 43 47
c82 47 0 1.00394e-19 $X=1.855 $Y=1.51
c83 35 0 1.37013e-19 $X=1.59 $Y=1.51
r84 39 41 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=0.585 $Y=2.06
+ $X2=0.695 $Y2=2.06
r85 36 47 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.59 $Y=1.51
+ $X2=1.855 $Y2=1.51
r86 36 44 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.51
+ $X2=1.425 $Y2=1.51
r87 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.59
+ $Y=1.51 $X2=1.59 $Y2=1.51
r88 33 43 0.47666 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=0.785 $Y=1.53 $X2=0.695
+ $Y2=1.53
r89 33 35 40.3355 $w=2.28e-07 $l=8.05e-07 $layer=LI1_cond $X=0.785 $Y=1.53
+ $X2=1.59 $Y2=1.53
r90 32 41 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=1.895
+ $X2=0.695 $Y2=2.06
r91 31 43 6.30264 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=0.695 $Y=1.645
+ $X2=0.695 $Y2=1.53
r92 31 32 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.695 $Y=1.645
+ $X2=0.695 $Y2=1.895
r93 30 43 6.30264 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=0.695 $Y=1.415
+ $X2=0.695 $Y2=1.53
r94 29 30 33.8889 $w=1.78e-07 $l=5.5e-07 $layer=LI1_cond $X=0.695 $Y=0.865
+ $X2=0.695 $Y2=1.415
r95 27 29 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.605 $Y=0.78
+ $X2=0.695 $Y2=0.865
r96 27 28 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.605 $Y=0.78
+ $X2=0.345 $Y2=0.78
r97 23 28 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.25 $Y=0.695
+ $X2=0.345 $Y2=0.78
r98 23 25 13.4258 $w=1.88e-07 $l=2.3e-07 $layer=LI1_cond $X=0.25 $Y=0.695
+ $X2=0.25 $Y2=0.465
r99 19 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.675
+ $X2=1.855 $Y2=1.51
r100 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.855 $Y=1.675
+ $X2=1.855 $Y2=2.465
r101 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=1.51
r102 15 17 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=0.745
r103 11 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.675
+ $X2=1.425 $Y2=1.51
r104 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.425 $Y=1.675
+ $X2=1.425 $Y2=2.465
r105 7 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=1.51
r106 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.425 $Y=1.345 $X2=1.425
+ $Y2=0.745
r107 2 39 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.46
+ $Y=1.835 $X2=0.585 $Y2=2.06
r108 1 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.255 $X2=0.26 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%B 3 7 11 15 17 18 25
c53 25 0 1.37013e-19 $X=2.795 $Y=1.51
c54 15 0 7.17626e-20 $X=2.855 $Y=0.745
r55 25 26 9.23962 $w=3.13e-07 $l=6e-08 $layer=POLY_cond $X=2.795 $Y=1.51
+ $X2=2.855 $Y2=1.51
r56 23 25 52.3578 $w=3.13e-07 $l=3.4e-07 $layer=POLY_cond $X=2.455 $Y=1.51
+ $X2=2.795 $Y2=1.51
r57 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.455
+ $Y=1.51 $X2=2.455 $Y2=1.51
r58 21 23 15.3994 $w=3.13e-07 $l=1e-07 $layer=POLY_cond $X=2.355 $Y=1.51
+ $X2=2.455 $Y2=1.51
r59 18 24 6.36424 $w=3.33e-07 $l=1.85e-07 $layer=LI1_cond $X=2.64 $Y=1.582
+ $X2=2.455 $Y2=1.582
r60 17 24 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=2.16 $Y=1.582
+ $X2=2.455 $Y2=1.582
r61 13 26 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.345
+ $X2=2.855 $Y2=1.51
r62 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.855 $Y=1.345
+ $X2=2.855 $Y2=0.745
r63 9 25 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.675
+ $X2=2.795 $Y2=1.51
r64 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.795 $Y=1.675
+ $X2=2.795 $Y2=2.465
r65 5 21 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.675
+ $X2=2.355 $Y2=1.51
r66 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.355 $Y=1.675
+ $X2=2.355 $Y2=2.465
r67 1 21 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.345
+ $X2=2.355 $Y2=1.51
r68 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.355 $Y=1.345 $X2=2.355
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%C 3 7 11 15 17 18 19 28
c53 28 0 1.48228e-19 $X=4.335 $Y=1.51
c54 19 0 5.33186e-20 $X=4.56 $Y=1.665
r55 26 28 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.245 $Y=1.51
+ $X2=4.335 $Y2=1.51
r56 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.245
+ $Y=1.51 $X2=4.245 $Y2=1.51
r57 23 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.905 $Y=1.51
+ $X2=4.245 $Y2=1.51
r58 19 27 11.1698 $w=3.23e-07 $l=3.15e-07 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=4.245 $Y2=1.587
r59 18 27 5.85086 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=1.587
+ $X2=4.245 $Y2=1.587
r60 17 18 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.587
+ $X2=4.08 $Y2=1.587
r61 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.335 $Y=1.675
+ $X2=4.335 $Y2=1.51
r62 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.335 $Y=1.675
+ $X2=4.335 $Y2=2.465
r63 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.335 $Y=1.345
+ $X2=4.335 $Y2=1.51
r64 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.335 $Y=1.345
+ $X2=4.335 $Y2=0.765
r65 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.905 $Y=1.675
+ $X2=3.905 $Y2=1.51
r66 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.905 $Y=1.675
+ $X2=3.905 $Y2=2.465
r67 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.905 $Y=1.345
+ $X2=3.905 $Y2=1.51
r68 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.905 $Y=1.345
+ $X2=3.905 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%D 3 7 11 15 17 18 27
c39 18 0 1.48228e-19 $X=5.52 $Y=1.665
c40 11 0 5.33186e-20 $X=5.195 $Y=2.465
r41 26 27 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.195 $Y=1.51
+ $X2=5.205 $Y2=1.51
r42 24 26 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=5.1 $Y=1.51
+ $X2=5.195 $Y2=1.51
r43 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.1
+ $Y=1.51 $X2=5.1 $Y2=1.51
r44 21 24 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=4.765 $Y=1.51
+ $X2=5.1 $Y2=1.51
r45 18 25 14.8931 $w=3.23e-07 $l=4.2e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.1 $Y2=1.587
r46 17 25 2.12759 $w=3.23e-07 $l=6e-08 $layer=LI1_cond $X=5.04 $Y=1.587 $X2=5.1
+ $Y2=1.587
r47 13 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.205 $Y=1.345
+ $X2=5.205 $Y2=1.51
r48 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.205 $Y=1.345
+ $X2=5.205 $Y2=0.765
r49 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.195 $Y=1.675
+ $X2=5.195 $Y2=1.51
r50 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.195 $Y=1.675
+ $X2=5.195 $Y2=2.465
r51 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.765 $Y=1.675
+ $X2=4.765 $Y2=1.51
r52 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.765 $Y=1.675
+ $X2=4.765 $Y2=2.465
r53 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.765 $Y=1.345
+ $X2=4.765 $Y2=1.51
r54 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.765 $Y=1.345
+ $X2=4.765 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%VPWR 1 2 3 4 5 18 24 28 30 32 36 38 43 48
+ 53 58 64 67 70 78 82
r73 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r74 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r76 70 74 11.5356 $w=1.008e-06 $l=9.55e-07 $layer=LI1_cond $X=3.35 $Y=2.375
+ $X2=3.35 $Y2=3.33
r77 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r79 62 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r80 62 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r82 59 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.715 $Y=3.33
+ $X2=4.55 $Y2=3.33
r83 59 61 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.715 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 58 81 4.59886 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=5.245 $Y=3.33
+ $X2=5.502 $Y2=3.33
r85 58 61 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.245 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 57 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 57 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r88 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r89 54 74 11.793 $w=1.7e-07 $l=5.05e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.35 $Y2=3.33
r90 54 56 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.385 $Y=3.33
+ $X2=4.55 $Y2=3.33
r92 53 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.385 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 52 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r95 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=3.33
+ $X2=2.105 $Y2=3.33
r96 49 51 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.27 $Y=3.33 $X2=2.64
+ $Y2=3.33
r97 48 74 11.793 $w=1.7e-07 $l=5.05e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=3.35 $Y2=3.33
r98 48 51 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r100 47 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r101 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 44 64 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.145 $Y2=3.33
r103 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=2.105 $Y2=3.33
r105 43 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 41 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 38 64 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.145 $Y2=3.33
r109 38 40 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.72 $Y2=3.33
r110 36 75 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r111 36 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 32 35 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=5.41 $Y=2.005
+ $X2=5.41 $Y2=2.95
r113 30 81 3.16731 $w=3.3e-07 $l=1.27609e-07 $layer=LI1_cond $X=5.41 $Y=3.245
+ $X2=5.502 $Y2=3.33
r114 30 35 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.41 $Y=3.245
+ $X2=5.41 $Y2=2.95
r115 26 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=3.33
r116 26 28 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=2.39
r117 22 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=3.245
+ $X2=2.105 $Y2=3.33
r118 22 24 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.105 $Y=3.245
+ $X2=2.105 $Y2=2.385
r119 18 21 14.8604 $w=3.78e-07 $l=4.9e-07 $layer=LI1_cond $X=1.145 $Y=1.98
+ $X2=1.145 $Y2=2.47
r120 16 64 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=3.33
r121 16 21 23.5038 $w=3.78e-07 $l=7.75e-07 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=2.47
r122 5 35 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.27
+ $Y=1.835 $X2=5.41 $Y2=2.95
r123 5 32 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=5.27
+ $Y=1.835 $X2=5.41 $Y2=2.005
r124 4 28 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=4.41
+ $Y=1.835 $X2=4.55 $Y2=2.39
r125 3 70 200 $w=1.7e-07 $l=1.05603e-06 $layer=licon1_PDIFF $count=3 $X=2.87
+ $Y=1.835 $X2=3.69 $Y2=2.375
r126 3 70 200 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=3 $X=2.87
+ $Y=1.835 $X2=3.01 $Y2=2.375
r127 2 24 300 $w=1.7e-07 $l=6.31467e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.835 $X2=2.105 $Y2=2.385
r128 1 21 300 $w=1.7e-07 $l=7.84825e-07 $layer=licon1_PDIFF $count=2 $X=0.875
+ $Y=1.835 $X2=1.21 $Y2=2.47
r129 1 18 600 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=0.875
+ $Y=1.835 $X2=1.04 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%Y 1 2 3 4 5 18 20 22 24 26 27 29 30 32 34
+ 40 41 42 43 52 55 62 67
r79 43 55 5.28167 $w=1.85e-07 $l=9.5e-08 $layer=LI1_cond $X=4.12 $Y=2.02
+ $X2=4.025 $Y2=2.02
r80 43 67 13.7558 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.12 $Y=2.12
+ $X2=4.12 $Y2=2.455
r81 43 55 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=4.01 $Y=2.02
+ $X2=4.025 $Y2=2.02
r82 42 43 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=3.6 $Y=2.02 $X2=4.01
+ $Y2=2.02
r83 42 56 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=3.6 $Y=2.02 $X2=3.215
+ $Y2=2.02
r84 41 52 7.31317 $w=2e-07 $l=1.55e-07 $layer=LI1_cond $X=3.06 $Y=2.02 $X2=2.905
+ $Y2=2.02
r85 41 56 7.31317 $w=2e-07 $l=1.55e-07 $layer=LI1_cond $X=3.06 $Y=2.02 $X2=3.215
+ $Y2=2.02
r86 40 53 6.27338 $w=1.85e-07 $l=1.18e-07 $layer=LI1_cond $X=2.557 $Y=2.02
+ $X2=2.675 $Y2=2.02
r87 40 62 12.1936 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=2.557 $Y=2.12
+ $X2=2.557 $Y2=2.455
r88 40 52 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=2.7 $Y=2.02
+ $X2=2.905 $Y2=2.02
r89 40 53 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=2.7 $Y=2.02
+ $X2=2.675 $Y2=2.02
r90 32 39 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=2.09 $X2=4.98
+ $Y2=2.005
r91 32 34 47.866 $w=1.88e-07 $l=8.2e-07 $layer=LI1_cond $X=4.98 $Y=2.09 $X2=4.98
+ $Y2=2.91
r92 31 43 5.28167 $w=1.85e-07 $l=1.02225e-07 $layer=LI1_cond $X=4.215 $Y=2.005
+ $X2=4.12 $Y2=2.02
r93 30 39 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.885 $Y=2.005
+ $X2=4.98 $Y2=2.005
r94 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.885 $Y=2.005
+ $X2=4.215 $Y2=2.005
r95 29 41 0.176625 $w=3.1e-07 $l=1e-07 $layer=LI1_cond $X=3.06 $Y=1.92 $X2=3.06
+ $Y2=2.02
r96 28 29 25.0935 $w=3.08e-07 $l=6.75e-07 $layer=LI1_cond $X=3.06 $Y=1.245
+ $X2=3.06 $Y2=1.92
r97 26 28 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.905 $Y=1.16
+ $X2=3.06 $Y2=1.245
r98 26 27 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=2.905 $Y=1.16
+ $X2=1.805 $Y2=1.16
r99 25 37 4.42198 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.77 $Y=2.005
+ $X2=1.637 $Y2=2.005
r100 24 40 6.27338 $w=1.85e-07 $l=1.24274e-07 $layer=LI1_cond $X=2.44 $Y=2.005
+ $X2=2.557 $Y2=2.02
r101 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.44 $Y=2.005
+ $X2=1.77 $Y2=2.005
r102 20 37 2.82608 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.637 $Y=2.09
+ $X2=1.637 $Y2=2.005
r103 20 22 35.6605 $w=2.63e-07 $l=8.2e-07 $layer=LI1_cond $X=1.637 $Y=2.09
+ $X2=1.637 $Y2=2.91
r104 16 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.64 $Y=1.075
+ $X2=1.805 $Y2=1.16
r105 16 18 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=1.64 $Y=1.075
+ $X2=1.64 $Y2=0.68
r106 5 39 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=4.84
+ $Y=1.835 $X2=4.98 $Y2=2.085
r107 5 34 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.84
+ $Y=1.835 $X2=4.98 $Y2=2.91
r108 4 43 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=3.98
+ $Y=1.835 $X2=4.12 $Y2=2.035
r109 4 67 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=3.98
+ $Y=1.835 $X2=4.12 $Y2=2.455
r110 3 40 600 $w=1.7e-07 $l=2.33238e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.835 $X2=2.58 $Y2=2.005
r111 3 62 300 $w=1.7e-07 $l=6.90941e-07 $layer=licon1_PDIFF $count=2 $X=2.43
+ $Y=1.835 $X2=2.58 $Y2=2.455
r112 2 37 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=2.085
r113 2 22 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=2.91
r114 1 18 91 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.325 $X2=1.64 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%VGND 1 2 9 13 15 17 22 32 33 36 39
r57 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r58 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r59 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r60 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r61 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=4.99
+ $Y2=0
r62 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.155 $Y=0 $X2=5.52
+ $Y2=0
r63 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r64 28 29 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r65 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r66 25 28 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r67 25 26 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r68 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r69 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r70 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=0 $X2=4.99
+ $Y2=0
r71 22 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.825 $Y=0 $X2=4.56
+ $Y2=0
r72 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r73 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r74 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r75 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r76 15 29 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.56
+ $Y2=0
r77 15 26 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.2
+ $Y2=0
r78 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0
r79 11 13 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0.47
r80 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r81 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0.42
r82 2 13 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=4.84
+ $Y=0.345 $X2=4.99 $Y2=0.47
r83 1 9 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.255 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%A_217_65# 1 2 3 12 14 15 19 21 23 24
c41 14 0 7.17626e-20 $X=1.975 $Y=0.34
r42 23 24 5.31268 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=3.07 $Y=0.775
+ $X2=2.975 $Y2=0.775
r43 21 24 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.305 $Y=0.815
+ $X2=2.975 $Y2=0.815
r44 17 21 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.14 $Y=0.725
+ $X2=2.305 $Y2=0.815
r45 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.14 $Y=0.725
+ $X2=2.14 $Y2=0.45
r46 16 19 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.45
r47 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=2.14 $Y2=0.425
r48 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=1.305 $Y2=0.34
r49 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.175 $Y=0.425
+ $X2=1.305 $Y2=0.34
r50 10 12 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=1.175 $Y=0.425
+ $X2=1.175 $Y2=0.47
r51 3 23 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.325 $X2=3.07 $Y2=0.81
r52 2 19 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.325 $X2=2.14 $Y2=0.45
r53 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.325 $X2=1.21 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%A_486_65# 1 2 7 11 13
r28 13 16 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=0.34
+ $X2=2.64 $Y2=0.47
r29 9 11 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.12 $Y=0.425
+ $X2=4.12 $Y2=0.47
r30 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=0.34
+ $X2=2.64 $Y2=0.34
r31 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.955 $Y=0.34
+ $X2=4.12 $Y2=0.425
r32 7 8 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=3.955 $Y=0.34
+ $X2=2.805 $Y2=0.34
r33 2 11 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.98
+ $Y=0.345 $X2=4.12 $Y2=0.47
r34 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.325 $X2=2.64 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_2%A_697_69# 1 2 3 12 14 15 18 20 24 26
r43 22 24 24.4894 $w=2.78e-07 $l=5.95e-07 $layer=LI1_cond $X=5.465 $Y=1.085
+ $X2=5.465 $Y2=0.49
r44 21 26 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.655 $Y=1.17 $X2=4.555
+ $Y2=1.17
r45 20 22 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=5.325 $Y=1.17
+ $X2=5.465 $Y2=1.085
r46 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.325 $Y=1.17
+ $X2=4.655 $Y2=1.17
r47 16 26 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=1.085
+ $X2=4.555 $Y2=1.17
r48 16 18 32.9955 $w=1.98e-07 $l=5.95e-07 $layer=LI1_cond $X=4.555 $Y=1.085
+ $X2=4.555 $Y2=0.49
r49 14 26 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.455 $Y=1.17 $X2=4.555
+ $Y2=1.17
r50 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.455 $Y=1.17
+ $X2=3.775 $Y2=1.17
r51 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.61 $Y=1.085
+ $X2=3.775 $Y2=1.17
r52 10 12 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.61 $Y=1.085
+ $X2=3.61 $Y2=0.68
r53 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.28
+ $Y=0.345 $X2=5.42 $Y2=0.49
r54 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.41
+ $Y=0.345 $X2=4.55 $Y2=0.49
r55 1 12 91 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=2 $X=3.485
+ $Y=0.345 $X2=3.61 $Y2=0.68
.ends

