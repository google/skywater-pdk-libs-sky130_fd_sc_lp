* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4b_m A B C D_N VGND VNB VPB VPWR Y
X0 Y a_33_68# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR A a_312_496# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_312_496# B a_384_496# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_384_496# C a_456_496# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_33_68# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_33_68# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_456_496# a_33_68# Y VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
