* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
X0 VGND a_609_485# a_795_423# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_574_47# a_200_481# a_609_485# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_609_485# a_310_485# a_754_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_27_481# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VGND GATE_N a_200_481# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_795_423# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_754_47# a_795_423# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_795_423# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR a_609_485# a_795_423# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR GATE_N a_200_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_310_485# a_200_481# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_27_481# a_537_485# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 VGND a_27_481# a_574_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 Q a_795_423# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 Q a_795_423# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VGND a_795_423# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_310_485# a_200_481# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_27_481# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 Q a_795_423# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_717_485# a_795_423# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 Q a_795_423# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VPWR a_795_423# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_609_485# a_200_481# a_717_485# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_537_485# a_310_485# a_609_485# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
