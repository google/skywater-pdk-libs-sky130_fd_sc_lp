* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor2_2 A B VGND VNB VPB VPWR X
X0 a_814_65# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 X B a_814_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND B a_149_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND A a_149_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_149_65# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND a_149_65# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR A a_149_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_149_65# B a_149_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR B a_532_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND A a_814_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_532_367# a_149_65# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_814_65# B X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 X a_149_65# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_149_367# B a_149_65# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_532_367# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_532_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_149_65# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 X a_149_65# a_532_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR A a_532_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_149_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
