* NGSPICE file created from sky130_fd_sc_lp__nor3_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor3_lp A B C VGND VNB VPB VPWR Y
M1000 a_173_57# C Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.373e+11p ps=2.81e+06u
M1001 a_297_409# C Y VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=2.85e+11p ps=2.57e+06u
M1002 VGND C a_173_57# VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=0p ps=0u
M1003 Y B a_331_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 VPWR A a_395_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=3.2e+11p ps=2.64e+06u
M1005 a_395_409# B a_297_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_331_57# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_489_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1008 a_489_57# A Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

