# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.940000 1.140000 2.270000 1.765000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.785000 0.375000 8.050000 3.075000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.425000 2.490000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.095000  0.085000 0.425000 0.670000 ;
      RECT 0.095000  2.660000 0.425000 3.245000 ;
      RECT 0.595000  0.330000 1.040000 3.050000 ;
      RECT 1.210000  0.640000 1.585000 1.935000 ;
      RECT 1.210000  1.935000 2.270000 2.105000 ;
      RECT 1.210000  2.105000 1.420000 2.865000 ;
      RECT 1.590000  2.285000 1.920000 3.245000 ;
      RECT 1.755000  0.085000 2.035000 0.970000 ;
      RECT 2.090000  2.105000 2.270000 2.760000 ;
      RECT 2.090000  2.760000 3.690000 2.940000 ;
      RECT 2.225000  0.640000 2.620000 0.970000 ;
      RECT 2.440000  0.970000 2.620000 1.220000 ;
      RECT 2.440000  1.220000 2.630000 2.590000 ;
      RECT 2.790000  0.640000 3.060000 0.865000 ;
      RECT 2.790000  0.865000 3.340000 1.035000 ;
      RECT 2.800000  1.385000 2.970000 2.760000 ;
      RECT 3.140000  1.035000 3.340000 1.055000 ;
      RECT 3.140000  1.055000 4.425000 1.225000 ;
      RECT 3.140000  1.225000 3.350000 2.590000 ;
      RECT 3.520000  0.085000 4.425000 0.885000 ;
      RECT 3.520000  2.285000 5.165000 2.455000 ;
      RECT 3.520000  2.455000 3.690000 2.760000 ;
      RECT 3.605000  1.405000 3.935000 1.915000 ;
      RECT 3.605000  1.915000 4.815000 2.115000 ;
      RECT 3.975000  2.625000 4.305000 3.245000 ;
      RECT 4.175000  1.225000 4.425000 1.675000 ;
      RECT 4.595000  0.585000 4.805000 1.915000 ;
      RECT 4.975000  1.295000 5.305000 1.475000 ;
      RECT 4.985000  1.475000 5.305000 1.555000 ;
      RECT 4.985000  1.555000 5.165000 2.285000 ;
      RECT 5.145000  0.645000 5.655000 1.125000 ;
      RECT 5.335000  1.875000 5.655000 2.755000 ;
      RECT 5.485000  1.125000 6.825000 1.295000 ;
      RECT 5.485000  1.295000 5.655000 1.875000 ;
      RECT 6.000000  0.085000 6.520000 0.945000 ;
      RECT 6.025000  1.465000 6.355000 1.635000 ;
      RECT 6.025000  1.635000 7.435000 1.645000 ;
      RECT 6.025000  1.645000 7.165000 1.805000 ;
      RECT 6.150000  1.975000 6.530000 3.245000 ;
      RECT 6.565000  1.295000 6.825000 1.455000 ;
      RECT 6.690000  0.415000 7.165000 0.945000 ;
      RECT 6.750000  1.805000 7.165000 2.755000 ;
      RECT 6.995000  0.945000 7.165000 1.425000 ;
      RECT 6.995000  1.425000 7.435000 1.635000 ;
      RECT 7.335000  0.085000 7.615000 1.255000 ;
      RECT 7.335000  1.815000 7.615000 3.245000 ;
      RECT 8.220000  0.085000 8.455000 1.255000 ;
      RECT 8.220000  1.815000 8.455000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_lp__dfxtp_2
END LIBRARY
