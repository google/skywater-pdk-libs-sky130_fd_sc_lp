* File: sky130_fd_sc_lp__and4_lp.spice
* Created: Wed Sep  2 09:33:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4_lp.pex.spice"
.subckt sky130_fd_sc_lp__and4_lp  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1000 A_230_55# N_D_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1659 PD=0.66 PS=1.63 NRD=18.564 NRS=31.428 M=1 R=2.8 SA=75000.3
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1014 A_308_55# N_C_M1014_g A_230_55# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=44.28 NRS=18.564 M=1 R=2.8 SA=75000.7 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1001 A_422_55# N_B_M1001_g A_308_55# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=44.28 M=1 R=2.8 SA=75001.3 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_186_485#_M1002_d N_A_M1002_g A_422_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_720_55# N_A_186_485#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_X_M1010_d N_A_186_485#_M1010_g A_720_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_114_485# N_D_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.1197 PD=0.63 PS=1.41 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.8
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_186_485#_M1004_d N_D_M1004_g A_114_485# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1011 A_272_485# N_C_M1011_g N_A_186_485#_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1015 N_VPWR_M1015_d N_C_M1015_g A_272_485# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.4 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1007 A_430_485# N_B_M1007_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.8 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_186_485#_M1003_d N_B_M1003_g A_430_485# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.1
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1013 A_588_485# N_A_M1013_g N_A_186_485#_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g A_588_485# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.9 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1008 A_746_485# N_A_186_485#_M1008_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75003.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_186_485#_M1009_g A_746_485# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75003.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__and4_lp.pxi.spice"
*
.ends
*
*
