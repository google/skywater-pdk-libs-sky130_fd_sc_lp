* File: sky130_fd_sc_lp__dfsbp_2.spice
* Created: Fri Aug 28 10:22:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfsbp_2.pex.spice"
.subckt sky130_fd_sc_lp__dfsbp_2  VNB VPB CLK D SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1002 N_A_129_179#_M1002_d N_CLK_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1512 PD=1.37 PS=1.56 NRD=0 NRS=1.428 M=1 R=2.8
+ SA=75000.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_A_129_179#_M1036_g N_A_191_21#_M1036_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1491 AS=0.1197 PD=1.13 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1032 N_A_507_125#_M1032_d N_D_M1032_g N_VGND_M1036_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1491 PD=0.7 PS=1.13 NRD=0 NRS=99.996 M=1 R=2.8 SA=75001.1
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1033 N_A_593_125#_M1033_d N_A_129_179#_M1033_g N_A_507_125#_M1032_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 A_679_125# N_A_191_21#_M1021_g N_A_593_125#_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_721_99#_M1025_g A_679_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1512 AS=0.0441 PD=1.56 PS=0.63 NRD=1.428 NRS=14.28 M=1 R=2.8 SA=75002.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1023 A_996_169# N_A_593_125#_M1023_g N_A_721_99#_M1023_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_SET_B_M1022_g A_996_169# VNB NSHORT L=0.15 W=0.42
+ AD=0.0855057 AS=0.0441 PD=0.80434 PS=0.63 NRD=28.56 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_1173_125#_M1003_d N_A_593_125#_M1003_g N_VGND_M1022_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.130294 PD=1.81 PS=1.22566 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 N_A_1360_451#_M1020_d N_A_129_179#_M1020_g N_A_1280_159#_M1020_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0855057 AS=0.1113 PD=0.80434 PS=1.37 NRD=12.852
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1026 N_A_1173_125#_M1026_d N_A_191_21#_M1026_g N_A_1360_451#_M1020_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.3179 AS=0.130294 PD=2.7 PS=1.22566 NRD=82.812
+ NRS=9.372 M=1 R=4.26667 SA=75000.5 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1011 A_1677_91# N_A_1533_258#_M1011_g N_A_1280_159#_M1011_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_SET_B_M1014_g A_1677_91# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_1360_451#_M1007_g N_A_1533_258#_M1007_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=28.56 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1015 N_Q_N_M1015_d N_A_1360_451#_M1015_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1030 N_Q_N_M1015_d N_A_1360_451#_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=6.78 M=1 R=5.6 SA=75000.9
+ SB=75000.5 A=0.126 P=1.98 MULT=1
MM1018 N_A_2227_367#_M1018_d N_A_1360_451#_M1018_g N_VGND_M1030_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0896 PD=1.37 PS=0.81 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_Q_M1012_d N_A_2227_367#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1027 N_Q_M1012_d N_A_2227_367#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_129_179#_M1000_d N_CLK_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_A_129_179#_M1006_g N_A_191_21#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.165072 AS=0.1696 PD=1.55774 PS=1.81 NRD=36.9178 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1008 N_A_507_125#_M1008_d N_D_M1008_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.108328 PD=0.7 PS=1.02226 NRD=0 NRS=56.2829 M=1 R=2.8 SA=75000.7
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1037 N_A_593_125#_M1037_d N_A_191_21#_M1037_g N_A_507_125#_M1008_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=16.4101 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75004 A=0.063 P=1.14 MULT=1
MM1028 A_701_535# N_A_129_179#_M1028_g N_A_593_125#_M1037_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=23.443 NRS=2.3443 M=1 R=2.8
+ SA=75001.6 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1031 N_VPWR_M1031_d N_A_721_99#_M1031_g A_701_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.16485 AS=0.0441 PD=1.205 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.9
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1019 N_A_721_99#_M1019_d N_A_593_125#_M1019_g N_VPWR_M1031_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.20265 AS=0.16485 PD=1.385 PS=1.205 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002.8 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_SET_B_M1017_g N_A_721_99#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0896 AS=0.20265 PD=0.81 PS=1.385 NRD=44.5417 NRS=0 M=1 R=2.8
+ SA=75004 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 A_1288_451# N_A_593_125#_M1010_g N_VPWR_M1017_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.0882 AS=0.1792 PD=1.05 PS=1.62 NRD=11.7215 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1009 N_A_1360_451#_M1009_d N_A_129_179#_M1009_g A_1288_451# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1862 AS=0.0882 PD=1.64 PS=1.05 NRD=2.3443 NRS=11.7215 M=1 R=5.6
+ SA=75002.7 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1029 A_1468_451# N_A_191_21#_M1029_g N_A_1360_451#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.06825 AS=0.0931 PD=0.745 PS=0.82 NRD=50.4123 NRS=46.886 M=1 R=2.8
+ SA=75001.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A_1533_258#_M1013_g A_1468_451# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.06825 PD=0.7 PS=0.745 NRD=0 NRS=50.4123 M=1 R=2.8
+ SA=75001.6 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_1360_451#_M1005_d N_SET_B_M1005_g N_VPWR_M1013_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_A_1360_451#_M1024_g N_A_1533_258#_M1024_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=46.886 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1024_d N_A_1360_451#_M1004_g N_Q_N_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.4 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1035 N_VPWR_M1035_d N_A_1360_451#_M1035_g N_Q_N_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.268115 AS=0.1764 PD=2.16853 PS=1.54 NRD=4.9447 NRS=0 M=1 R=8.4
+ SA=75000.8 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1034 N_A_2227_367#_M1034_d N_A_1360_451#_M1034_g N_VPWR_M1035_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.136185 PD=1.81 PS=1.10147 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A_2227_367#_M1001_g N_Q_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_A_2227_367#_M1016_g N_Q_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX38_noxref VNB VPB NWDIODE A=24.8791 P=30.41
*
.include "sky130_fd_sc_lp__dfsbp_2.pxi.spice"
*
.ends
*
*
