* File: sky130_fd_sc_lp__or4_1.pex.spice
* Created: Wed Sep  2 10:31:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4_1%D 3 7 9 10 11 16
r33 16 19 82.4947 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=0.36 $Y=1.005
+ $X2=0.36 $Y2=1.51
r34 16 18 46.8261 $w=5.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.36 $Y=1.005
+ $X2=0.36 $Y2=0.84
r35 10 11 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.247 $Y=1.295
+ $X2=0.247 $Y2=1.665
r36 9 10 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.247 $Y=0.925
+ $X2=0.247 $Y2=1.295
r37 9 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r38 7 19 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=0.54 $Y=2.61 $X2=0.54
+ $Y2=1.51
r39 3 18 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.51 $Y=0.445
+ $X2=0.51 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_1%C 3 7 11 12 13 14 18 19
c40 19 0 1.04888e-19 $X=0.99 $Y=1.07
r41 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.99
+ $Y=1.07 $X2=0.99 $Y2=1.07
r42 13 14 7.76402 $w=5.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.87 $Y=1.295
+ $X2=0.87 $Y2=1.665
r43 13 19 4.72136 $w=5.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.87 $Y=1.295
+ $X2=0.87 $Y2=1.07
r44 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.99 $Y=1.41
+ $X2=0.99 $Y2=1.07
r45 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.41
+ $X2=0.99 $Y2=1.575
r46 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=0.905
+ $X2=0.99 $Y2=1.07
r47 7 10 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.94 $Y=0.445
+ $X2=0.94 $Y2=0.905
r48 3 12 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=0.9 $Y=2.61 $X2=0.9
+ $Y2=1.575
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_1%B 3 6 9 11 12 16 17
c45 9 0 1.04888e-19 $X=1.71 $Y=0.445
r46 16 18 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.575 $Y=1.17
+ $X2=1.575 $Y2=1.005
r47 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.56
+ $Y=1.17 $X2=1.56 $Y2=1.17
r48 11 12 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.585 $Y=1.295
+ $X2=1.585 $Y2=1.665
r49 11 17 3.79093 $w=3.78e-07 $l=1.25e-07 $layer=LI1_cond $X=1.585 $Y=1.295
+ $X2=1.585 $Y2=1.17
r50 9 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.71 $Y=0.445
+ $X2=1.71 $Y2=1.005
r51 5 16 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=1.575 $Y=1.215
+ $X2=1.575 $Y2=1.17
r52 5 6 33.1044 $w=4.2e-07 $l=2.5e-07 $layer=POLY_cond $X=1.575 $Y=1.215
+ $X2=1.575 $Y2=1.465
r53 1 6 69.0671 $w=3.28e-07 $l=6.07413e-07 $layer=POLY_cond $X=1.26 $Y=1.935
+ $X2=1.575 $Y2=1.465
r54 1 3 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.26 $Y=1.935
+ $X2=1.26 $Y2=2.61
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_1%A 1 3 4 5 7 10 12 15 16
c55 15 0 1.09618e-19 $X=2.16 $Y=1.51
r56 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.51
+ $X2=2.16 $Y2=1.675
r57 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.51 $X2=2.16 $Y2=1.51
r58 12 16 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=1.51
r59 8 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.345
+ $X2=2.16 $Y2=1.51
r60 8 10 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.16 $Y=1.345 $X2=2.16
+ $Y2=0.445
r61 7 17 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.07 $Y=2.145 $X2=2.07
+ $Y2=1.675
r62 4 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.995 $Y=2.22
+ $X2=2.07 $Y2=2.145
r63 4 5 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.995 $Y=2.22 $X2=1.695
+ $Y2=2.22
r64 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.62 $Y=2.295
+ $X2=1.695 $Y2=2.22
r65 1 3 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.62 $Y=2.295 $X2=1.62
+ $Y2=2.61
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_1%A_40_480# 1 2 3 10 12 15 19 22 25 27 28 31 34
+ 35 36 37 42 44 45 46 50
c105 45 0 1.09618e-19 $X=2.165 $Y=2.095
r106 45 46 7.84131 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=2.165 $Y=2.095
+ $X2=2.335 $Y2=2.095
r107 43 50 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.73 $Y=1.35
+ $X2=2.885 $Y2=1.35
r108 43 47 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.73 $Y=1.35 $X2=2.65
+ $Y2=1.35
r109 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.73
+ $Y=1.35 $X2=2.73 $Y2=1.35
r110 40 42 26.7367 $w=2.48e-07 $l=5.8e-07 $layer=LI1_cond $X=2.69 $Y=1.93
+ $X2=2.69 $Y2=1.35
r111 39 42 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2.69 $Y=1.245
+ $X2=2.69 $Y2=1.35
r112 37 40 6.85268 $w=2.2e-07 $l=1.71391e-07 $layer=LI1_cond $X=2.565 $Y=2.04
+ $X2=2.69 $Y2=1.93
r113 37 46 12.0483 $w=2.18e-07 $l=2.3e-07 $layer=LI1_cond $X=2.565 $Y=2.04
+ $X2=2.335 $Y2=2.04
r114 35 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.565 $Y=1.16
+ $X2=2.69 $Y2=1.245
r115 35 36 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.565 $Y=1.16
+ $X2=2.115 $Y2=1.16
r116 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.03 $Y=1.075
+ $X2=2.115 $Y2=1.16
r117 33 44 4.02809 $w=2.27e-07 $l=1.1025e-07 $layer=LI1_cond $X=2.03 $Y=0.815
+ $X2=1.972 $Y2=0.73
r118 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.03 $Y=0.815
+ $X2=2.03 $Y2=1.075
r119 29 44 4.02809 $w=2.27e-07 $l=8.5e-08 $layer=LI1_cond $X=1.972 $Y=0.645
+ $X2=1.972 $Y2=0.73
r120 29 31 8.08732 $w=2.83e-07 $l=2e-07 $layer=LI1_cond $X=1.972 $Y=0.645
+ $X2=1.972 $Y2=0.445
r121 27 44 2.40986 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1.83 $Y=0.73
+ $X2=1.972 $Y2=0.73
r122 27 28 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.83 $Y=0.73
+ $X2=0.82 $Y2=0.73
r123 23 28 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.71 $Y=0.645
+ $X2=0.82 $Y2=0.73
r124 23 25 10.4768 $w=2.18e-07 $l=2e-07 $layer=LI1_cond $X=0.71 $Y=0.645
+ $X2=0.71 $Y2=0.445
r125 22 45 74.2439 $w=2.58e-07 $l=1.675e-06 $layer=LI1_cond $X=0.49 $Y=2.13
+ $X2=2.165 $Y2=2.13
r126 17 22 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=0.325 $Y=2.26
+ $X2=0.49 $Y2=2.13
r127 17 19 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.325 $Y=2.26
+ $X2=0.325 $Y2=2.61
r128 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.515
+ $X2=2.885 $Y2=1.35
r129 13 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.885 $Y=1.515
+ $X2=2.885 $Y2=2.465
r130 10 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.185
+ $X2=2.65 $Y2=1.35
r131 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.65 $Y=1.185
+ $X2=2.65 $Y2=0.655
r132 3 19 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=2.4 $X2=0.325 $Y2=2.61
r133 2 31 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=1.785
+ $Y=0.235 $X2=1.945 $Y2=0.445
r134 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.235 $X2=0.725 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_1%VPWR 1 4 6 11 13 14
r28 22 25 0.364179 $w=1.005e-06 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=2.867
+ $X2=2.67 $Y2=2.867
r29 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 20 22 4.49154 $w=1.005e-06 $l=3.7e-07 $layer=LI1_cond $X=2.27 $Y=2.867
+ $X2=2.64 $Y2=2.867
r31 17 20 7.16219 $w=1.005e-06 $l=5.9e-07 $layer=LI1_cond $X=1.68 $Y=2.867
+ $X2=2.27 $Y2=2.867
r32 14 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r34 11 25 12.8781 $w=1.005e-06 $l=5.39225e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.67 $Y2=2.867
r35 11 13 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 8 9 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33 $X2=0.24
+ $Y2=3.33
r37 6 17 10.9965 $w=1.005e-06 $l=4.67973e-07 $layer=LI1_cond $X=1.67 $Y=3.33
+ $X2=1.68 $Y2=2.867
r38 6 8 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.67 $Y=3.33 $X2=0.24
+ $Y2=3.33
r39 4 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 4 9 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 4 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 1 25 600 $w=1.7e-07 $l=1.21937e-06 $layer=licon1_PDIFF $count=1 $X=1.695
+ $Y=2.4 $X2=2.67 $Y2=2.95
r43 1 25 600 $w=1.7e-07 $l=1.01661e-06 $layer=licon1_PDIFF $count=1 $X=1.695
+ $Y=2.4 $X2=2.67 $Y2=2.485
r44 1 20 300 $w=1.7e-07 $l=6.71844e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=2.4 $X2=2.27 $Y2=2.61
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_1%X 1 2 7 8 9 10 11 12 13 24 41
r17 24 46 0.853661 $w=2.68e-07 $l=2e-08 $layer=LI1_cond $X=3.14 $Y=0.925
+ $X2=3.14 $Y2=0.905
r18 13 38 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.14 $Y=2.775
+ $X2=3.14 $Y2=2.91
r19 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=2.405
+ $X2=3.14 $Y2=2.775
r20 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.14 $Y=1.98
+ $X2=3.14 $Y2=2.405
r21 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.14 $Y=1.665
+ $X2=3.14 $Y2=1.98
r22 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=1.295
+ $X2=3.14 $Y2=1.665
r23 8 46 4.074 $w=5.73e-07 $l=3.3e-08 $layer=LI1_cond $X=2.987 $Y=0.872
+ $X2=2.987 $Y2=0.905
r24 8 9 14.4269 $w=2.68e-07 $l=3.38e-07 $layer=LI1_cond $X=3.14 $Y=0.957
+ $X2=3.14 $Y2=1.295
r25 8 24 1.36586 $w=2.68e-07 $l=3.2e-08 $layer=LI1_cond $X=3.14 $Y=0.957
+ $X2=3.14 $Y2=0.925
r26 7 8 6.59403 $w=5.73e-07 $l=3.17e-07 $layer=LI1_cond $X=2.987 $Y=0.555
+ $X2=2.987 $Y2=0.872
r27 7 41 3.64024 $w=5.73e-07 $l=1.75e-07 $layer=LI1_cond $X=2.987 $Y=0.555
+ $X2=2.987 $Y2=0.38
r28 2 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.91
r29 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=1.98
r30 1 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.725
+ $Y=0.235 $X2=2.865 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_1%VGND 1 2 3 10 12 16 21 22 23 35 36 44 47
r48 46 47 9.89636 $w=5.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=0.195
+ $X2=1.66 $Y2=0.195
r49 42 46 6.30077 $w=5.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=0.195
+ $X2=1.495 $Y2=0.195
r50 42 44 10.8575 $w=5.58e-07 $l=2.1e-07 $layer=LI1_cond $X=1.2 $Y=0.195
+ $X2=0.99 $Y2=0.195
r51 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r54 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r55 32 47 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.66
+ $Y2=0
r56 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r57 29 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r58 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r59 28 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.99
+ $Y2=0
r60 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 26 39 4.42822 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r62 26 28 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r63 23 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r64 23 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r65 21 32 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.16
+ $Y2=0
r66 21 22 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.407
+ $Y2=0
r67 20 35 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.12
+ $Y2=0
r68 20 22 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.407
+ $Y2=0
r69 16 18 16.9339 $w=2.43e-07 $l=3.6e-07 $layer=LI1_cond $X=2.407 $Y=0.38
+ $X2=2.407 $Y2=0.74
r70 14 22 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.407 $Y=0.085
+ $X2=2.407 $Y2=0
r71 14 16 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=2.407 $Y=0.085
+ $X2=2.407 $Y2=0.38
r72 10 39 3.08945 $w=3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.215 $Y2=0
r73 10 12 13.8293 $w=2.98e-07 $l=3.6e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.445
r74 3 18 182 $w=1.7e-07 $l=5.96678e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.235 $X2=2.435 $Y2=0.74
r75 3 16 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.235 $X2=2.435 $Y2=0.38
r76 2 46 91 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.235 $X2=1.495 $Y2=0.38
r77 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.235 $X2=0.295 $Y2=0.445
.ends

