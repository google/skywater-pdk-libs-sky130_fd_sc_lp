* File: sky130_fd_sc_lp__dfxtp_lp.pex.spice
* Created: Wed Sep  2 09:45:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%CLK 3 7 11 15 17 18 19 23
c44 23 0 2.79125e-19 $X=0.62 $Y=1.34
r45 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.62
+ $Y=1.34 $X2=0.62 $Y2=1.34
r46 19 24 9.85642 $w=3.78e-07 $l=3.25e-07 $layer=LI1_cond $X=0.645 $Y=1.665
+ $X2=0.645 $Y2=1.34
r47 18 24 1.36474 $w=3.78e-07 $l=4.5e-08 $layer=LI1_cond $X=0.645 $Y=1.295
+ $X2=0.645 $Y2=1.34
r48 16 23 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=0.597 $Y=1.658
+ $X2=0.597 $Y2=1.34
r49 16 17 33.9275 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.597 $Y=1.658
+ $X2=0.597 $Y2=1.845
r50 15 23 2.22462 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=0.597 $Y=1.325
+ $X2=0.597 $Y2=1.34
r51 7 17 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.66 $Y=2.545 $X2=0.66
+ $Y2=1.845
r52 1 15 24.6308 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=0.665 $Y=1.175
+ $X2=0.665 $Y2=1.325
r53 1 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.845 $Y=1.175
+ $X2=0.845 $Y2=0.495
r54 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.485 $Y=1.175
+ $X2=0.485 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%D 3 4 6 8 10 12 14 15 18 19
c43 15 0 1.11272e-19 $X=2.64 $Y=1.295
r44 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.55
+ $Y=1.335 $X2=2.55 $Y2=1.335
r45 18 21 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.55 $Y=1.245 $X2=2.55
+ $Y2=1.335
r46 18 19 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.245
+ $X2=2.55 $Y2=1.17
r47 15 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=1.335 $X2=2.55
+ $Y2=1.335
r48 14 22 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.16 $Y=1.335
+ $X2=2.55 $Y2=1.335
r49 10 13 21.6156 $w=2.33e-07 $l=8.44097e-08 $layer=POLY_cond $X=3.07 $Y=1.17
+ $X2=3.05 $Y2=1.245
r50 10 12 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.07 $Y=1.17
+ $X2=3.07 $Y2=0.835
r51 6 13 38.8528 $w=2.5e-07 $l=2e-07 $layer=POLY_cond $X=3.05 $Y=1.445 $X2=3.05
+ $Y2=1.245
r52 6 8 188.825 $w=2.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.05 $Y=1.445 $X2=3.05
+ $Y2=2.205
r53 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.245
+ $X2=2.55 $Y2=1.245
r54 4 13 13.0941 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.925 $Y=1.245
+ $X2=3.05 $Y2=1.245
r55 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.925 $Y=1.245
+ $X2=2.715 $Y2=1.245
r56 3 19 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.64 $Y=0.835
+ $X2=2.64 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%A_263_409# 1 2 7 9 12 14 17 19 21 24 25 26
+ 29 32 35 37 39 44 45 47 48 50 51 52 54 55 56 58 59 61 64 69 73 78
c192 69 0 2.18075e-19 $X=7.5 $Y=1.3
c193 44 0 1.78866e-19 $X=4.62 $Y=1.32
c194 39 0 6.06529e-20 $X=3.55 $Y=1.38
c195 26 0 8.68493e-20 $X=7.55 $Y=1.785
c196 24 0 1.11272e-19 $X=3.87 $Y=1.365
r197 77 78 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.435 $Y=1.32
+ $X2=4.36 $Y2=1.32
r198 73 83 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.51 $Y=1.38
+ $X2=7.51 $Y2=1.545
r199 73 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.51 $Y=1.38
+ $X2=7.51 $Y2=1.215
r200 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.51
+ $Y=1.38 $X2=7.51 $Y2=1.38
r201 69 72 2.97405 $w=3.08e-07 $l=8e-08 $layer=LI1_cond $X=7.5 $Y=1.3 $X2=7.5
+ $Y2=1.38
r202 61 63 10.6751 $w=3.38e-07 $l=2.3e-07 $layer=LI1_cond $X=1.845 $Y=0.495
+ $X2=1.845 $Y2=0.725
r203 58 59 9.86413 $w=5.53e-07 $l=1.65e-07 $layer=LI1_cond $X=1.567 $Y=2.19
+ $X2=1.567 $Y2=2.025
r204 55 69 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.345 $Y=1.3
+ $X2=7.5 $Y2=1.3
r205 55 56 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.345 $Y=1.3
+ $X2=6.68 $Y2=1.3
r206 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.595 $Y=1.215
+ $X2=6.68 $Y2=1.3
r207 53 54 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.595 $Y=1.035
+ $X2=6.595 $Y2=1.215
r208 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.51 $Y=0.95
+ $X2=6.595 $Y2=1.035
r209 51 52 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.51 $Y=0.95
+ $X2=6.14 $Y2=0.95
r210 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.055 $Y=0.865
+ $X2=6.14 $Y2=0.95
r211 49 50 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.055 $Y=0.625
+ $X2=6.055 $Y2=0.865
r212 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.97 $Y=0.54
+ $X2=6.055 $Y2=0.625
r213 47 48 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=5.97 $Y=0.54
+ $X2=4.715 $Y2=0.54
r214 45 77 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=4.62 $Y=1.32
+ $X2=4.435 $Y2=1.32
r215 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.62
+ $Y=1.32 $X2=4.62 $Y2=1.32
r216 42 48 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.62 $Y=0.625
+ $X2=4.715 $Y2=0.54
r217 42 44 40.5694 $w=1.88e-07 $l=6.95e-07 $layer=LI1_cond $X=4.62 $Y=0.625
+ $X2=4.62 $Y2=1.32
r218 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.38 $X2=3.55 $Y2=1.38
r219 37 67 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.02 $Y=1.38
+ $X2=3.02 $Y2=1.765
r220 37 39 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.105 $Y=1.38
+ $X2=3.55 $Y2=1.38
r221 36 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=1.765
+ $X2=1.76 $Y2=1.765
r222 35 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=1.765
+ $X2=3.02 $Y2=1.765
r223 35 36 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=2.935 $Y=1.765
+ $X2=1.845 $Y2=1.765
r224 33 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=1.85
+ $X2=1.76 $Y2=1.765
r225 33 59 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.76 $Y=1.85
+ $X2=1.76 $Y2=2.025
r226 32 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=1.68
+ $X2=1.76 $Y2=1.765
r227 32 63 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.76 $Y=1.68
+ $X2=1.76 $Y2=0.725
r228 27 58 2.41371 $w=5.53e-07 $l=1.12e-07 $layer=LI1_cond $X=1.567 $Y=2.302
+ $X2=1.567 $Y2=2.19
r229 27 29 12.8875 $w=5.53e-07 $l=5.98e-07 $layer=LI1_cond $X=1.567 $Y=2.302
+ $X2=1.567 $Y2=2.9
r230 26 83 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.6 $Y=1.785
+ $X2=7.6 $Y2=1.545
r231 24 40 51.2926 $w=3.6e-07 $l=3.2e-07 $layer=POLY_cond $X=3.87 $Y=1.365
+ $X2=3.55 $Y2=1.365
r232 24 25 20.0758 $w=2.55e-07 $l=1.8e-07 $layer=POLY_cond $X=3.87 $Y=1.365
+ $X2=3.87 $Y2=1.185
r233 19 26 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=7.55 $Y=1.91
+ $X2=7.55 $Y2=1.785
r234 19 21 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.55 $Y=1.91
+ $X2=7.55 $Y2=2.415
r235 17 82 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=7.5 $Y=0.835
+ $X2=7.5 $Y2=1.215
r236 12 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.435 $Y=1.155
+ $X2=4.435 $Y2=1.32
r237 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.435 $Y=1.155
+ $X2=4.435 $Y2=0.835
r238 11 25 20.0758 $w=2.55e-07 $l=1.83712e-07 $layer=POLY_cond $X=4.02 $Y=1.26
+ $X2=3.87 $Y2=1.185
r239 11 78 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.02 $Y=1.26
+ $X2=4.36 $Y2=1.26
r240 7 25 5.58633 $w=2.5e-07 $l=5.74108e-07 $layer=POLY_cond $X=3.995 $Y=1.7
+ $X2=3.87 $Y2=1.185
r241 7 9 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.995 $Y=1.7
+ $X2=3.995 $Y2=2.205
r242 2 58 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=2.045 $X2=1.455 $Y2=2.19
r243 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.315
+ $Y=2.045 $X2=1.455 $Y2=2.9
r244 1 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.71
+ $Y=0.285 $X2=1.85 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%A_1005_99# 1 2 7 9 12 16 17 19 20 23 27 29
+ 32 34 36
c105 29 0 1.20974e-20 $X=7.835 $Y=0.95
c106 17 0 1.07714e-19 $X=5.34 $Y=1.32
r107 40 42 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.1 $Y=1.32
+ $X2=5.26 $Y2=1.32
r108 36 38 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=7.28 $Y=0.82
+ $X2=7.28 $Y2=0.95
r109 31 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.92 $Y=1.035
+ $X2=7.92 $Y2=1.725
r110 30 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.445 $Y=0.95
+ $X2=7.28 $Y2=0.95
r111 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.835 $Y=0.95
+ $X2=7.92 $Y2=1.035
r112 29 30 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.835 $Y=0.95
+ $X2=7.445 $Y2=0.95
r113 28 34 8.61065 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=6.84 $Y=1.81
+ $X2=6.675 $Y2=1.79
r114 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.835 $Y=1.81
+ $X2=7.92 $Y2=1.725
r115 27 28 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=7.835 $Y=1.81
+ $X2=6.84 $Y2=1.81
r116 23 25 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=6.675 $Y=2.31
+ $X2=6.675 $Y2=2.77
r117 21 34 0.89609 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=6.675 $Y=1.895
+ $X2=6.675 $Y2=1.79
r118 21 23 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=6.675 $Y=1.895
+ $X2=6.675 $Y2=2.31
r119 19 34 8.61065 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=6.51 $Y=1.81
+ $X2=6.675 $Y2=1.79
r120 19 20 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=6.51 $Y=1.81
+ $X2=5.44 $Y2=1.81
r121 17 42 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.34 $Y=1.32 $X2=5.26
+ $Y2=1.32
r122 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.34
+ $Y=1.32 $X2=5.34 $Y2=1.32
r123 14 20 6.85817 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=5.342 $Y=1.725
+ $X2=5.44 $Y2=1.81
r124 14 16 23.035 $w=1.93e-07 $l=4.05e-07 $layer=LI1_cond $X=5.342 $Y=1.725
+ $X2=5.342 $Y2=1.32
r125 10 42 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.26 $Y=1.485
+ $X2=5.26 $Y2=1.32
r126 10 12 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=5.26 $Y=1.485
+ $X2=5.26 $Y2=2.205
r127 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.1 $Y=1.155
+ $X2=5.1 $Y2=1.32
r128 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.1 $Y=1.155 $X2=5.1
+ $Y2=0.835
r129 2 34 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=6.455
+ $Y=1.705 $X2=6.675 $Y2=1.85
r130 2 25 600 $w=1.7e-07 $l=1.16984e-06 $layer=licon1_PDIFF $count=1 $X=6.455
+ $Y=1.705 $X2=6.675 $Y2=2.77
r131 2 23 600 $w=1.7e-07 $l=7.06488e-07 $layer=licon1_PDIFF $count=1 $X=6.455
+ $Y=1.705 $X2=6.675 $Y2=2.31
r132 1 36 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=7.135
+ $Y=0.625 $X2=7.28 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%A_747_79# 1 2 9 13 15 19 21 26 29 33 36 37
+ 38 40 41 43 47 52
c124 19 0 1.20974e-20 $X=7.06 $Y=0.835
c125 15 0 9.2555e-20 $X=6.985 $Y=1.29
r126 51 52 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.7 $Y=1.38
+ $X2=6.775 $Y2=1.38
r127 50 51 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=6.33 $Y=1.38
+ $X2=6.7 $Y2=1.38
r128 44 50 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.165 $Y=1.38
+ $X2=6.33 $Y2=1.38
r129 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.165
+ $Y=1.38 $X2=6.165 $Y2=1.38
r130 41 43 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.79 $Y=1.38
+ $X2=6.165 $Y2=1.38
r131 40 41 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.705 $Y=1.215
+ $X2=5.79 $Y2=1.38
r132 39 40 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.705 $Y=0.975
+ $X2=5.705 $Y2=1.215
r133 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.62 $Y=0.89
+ $X2=5.705 $Y2=0.975
r134 37 38 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.62 $Y=0.89
+ $X2=5.065 $Y2=0.89
r135 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.98 $Y=0.975
+ $X2=5.065 $Y2=0.89
r136 35 36 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.98 $Y=0.975
+ $X2=4.98 $Y2=1.685
r137 34 47 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.505 $Y=1.77
+ $X2=4.34 $Y2=1.77
r138 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.895 $Y=1.77
+ $X2=4.98 $Y2=1.685
r139 33 34 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.895 $Y=1.77
+ $X2=4.505 $Y2=1.77
r140 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.34 $Y=2.28
+ $X2=4.34 $Y2=2.71
r141 27 47 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=1.855
+ $X2=4.34 $Y2=1.77
r142 27 29 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.34 $Y=1.855
+ $X2=4.34 $Y2=2.28
r143 26 47 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.26 $Y=1.685
+ $X2=4.34 $Y2=1.77
r144 25 26 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=4.26 $Y=0.685
+ $X2=4.26 $Y2=1.685
r145 21 25 7.59919 $w=3.1e-07 $l=1.92873e-07 $layer=LI1_cond $X=4.175 $Y=0.53
+ $X2=4.26 $Y2=0.685
r146 21 23 11.1527 $w=3.08e-07 $l=3e-07 $layer=LI1_cond $X=4.175 $Y=0.53
+ $X2=3.875 $Y2=0.53
r147 17 19 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=7.06 $Y=1.215
+ $X2=7.06 $Y2=0.835
r148 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.985 $Y=1.29
+ $X2=7.06 $Y2=1.215
r149 15 52 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.985 $Y=1.29
+ $X2=6.775 $Y2=1.29
r150 11 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.7 $Y=1.215
+ $X2=6.7 $Y2=1.38
r151 11 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=6.7 $Y=1.215
+ $X2=6.7 $Y2=0.835
r152 7 50 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.33 $Y=1.545
+ $X2=6.33 $Y2=1.38
r153 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.33 $Y=1.545
+ $X2=6.33 $Y2=2.205
r154 2 47 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=1.705 $X2=4.34 $Y2=1.85
r155 2 31 600 $w=1.7e-07 $l=1.10956e-06 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=1.705 $X2=4.34 $Y2=2.71
r156 2 29 600 $w=1.7e-07 $l=6.7611e-07 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=1.705 $X2=4.34 $Y2=2.28
r157 1 23 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3.735
+ $Y=0.395 $X2=3.875 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%A_27_57# 1 2 9 11 13 14 16 17 18 20 22 23
+ 24 25 26 29 31 35 37 41 43 45 46 52 53 54 57 63 65 69 71 72 74 75
c175 74 0 1.99528e-19 $X=1.33 $Y=0.99
c176 35 0 2.73522e-19 $X=4.685 $Y=2.355
c177 29 0 6.06529e-20 $X=3.66 $Y=0.605
c178 17 0 1.67093e-19 $X=1.995 $Y=0.855
r179 74 75 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.33
+ $Y=0.99 $X2=1.33 $Y2=0.99
r180 71 72 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.332 $Y=2.19
+ $X2=0.332 $Y2=2.025
r181 66 69 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=0.91
+ $X2=0.27 $Y2=0.91
r182 65 74 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=0.91
+ $X2=1.33 $Y2=0.91
r183 65 66 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.165 $Y=0.91
+ $X2=0.435 $Y2=0.91
r184 61 71 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=0.332 $Y=2.252
+ $X2=0.332 $Y2=2.19
r185 61 63 17.0343 $w=4.53e-07 $l=6.48e-07 $layer=LI1_cond $X=0.332 $Y=2.252
+ $X2=0.332 $Y2=2.9
r186 59 69 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.19 $Y=0.995
+ $X2=0.27 $Y2=0.91
r187 59 72 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.19 $Y=0.995
+ $X2=0.19 $Y2=2.025
r188 55 69 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=0.825
+ $X2=0.27 $Y2=0.91
r189 55 57 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.27 $Y=0.825
+ $X2=0.27 $Y2=0.495
r190 50 75 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.33 $Y=0.93 $X2=1.33
+ $Y2=0.99
r191 50 51 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.33 $Y=0.855
+ $X2=1.635 $Y2=0.855
r192 47 50 28.2021 $w=1.5e-07 $l=5.5e-08 $layer=POLY_cond $X=1.275 $Y=0.855
+ $X2=1.33 $Y2=0.855
r193 46 75 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.33 $Y=1.33
+ $X2=1.33 $Y2=0.99
r194 43 45 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=8.055 $Y=0.255
+ $X2=8.055 $Y2=0.585
r195 39 41 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.02 $Y=3.075
+ $X2=7.02 $Y2=2.415
r196 38 54 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.81 $Y=3.15
+ $X2=4.685 $Y2=3.15
r197 37 39 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=6.895 $Y=3.15
+ $X2=7.02 $Y2=3.075
r198 37 38 1069.12 $w=1.5e-07 $l=2.085e-06 $layer=POLY_cond $X=6.895 $Y=3.15
+ $X2=4.81 $Y2=3.15
r199 33 54 1.63566 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.685 $Y=3.075
+ $X2=4.685 $Y2=3.15
r200 33 35 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=4.685 $Y=3.075
+ $X2=4.685 $Y2=2.355
r201 32 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.735 $Y=0.18
+ $X2=3.66 $Y2=0.18
r202 31 43 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.98 $Y=0.18
+ $X2=8.055 $Y2=0.255
r203 31 32 2176.69 $w=1.5e-07 $l=4.245e-06 $layer=POLY_cond $X=7.98 $Y=0.18
+ $X2=3.735 $Y2=0.18
r204 27 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.66 $Y=0.255
+ $X2=3.66 $Y2=0.18
r205 27 29 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.66 $Y=0.255
+ $X2=3.66 $Y2=0.605
r206 25 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.585 $Y=0.18
+ $X2=3.66 $Y2=0.18
r207 25 26 705.053 $w=1.5e-07 $l=1.375e-06 $layer=POLY_cond $X=3.585 $Y=0.18
+ $X2=2.21 $Y2=0.18
r208 23 54 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.56 $Y=3.15
+ $X2=4.685 $Y2=3.15
r209 23 24 1238.33 $w=1.5e-07 $l=2.415e-06 $layer=POLY_cond $X=4.56 $Y=3.15
+ $X2=2.145 $Y2=3.15
r210 22 52 20.4101 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.135 $Y=0.78
+ $X2=2.102 $Y2=0.855
r211 21 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.135 $Y=0.255
+ $X2=2.21 $Y2=0.18
r212 21 22 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.135 $Y=0.255
+ $X2=2.135 $Y2=0.78
r213 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.07 $Y=3.075
+ $X2=2.145 $Y2=3.15
r214 19 52 20.4101 $w=1.5e-07 $l=8.95824e-08 $layer=POLY_cond $X=2.07 $Y=0.93
+ $X2=2.102 $Y2=0.855
r215 19 20 1099.88 $w=1.5e-07 $l=2.145e-06 $layer=POLY_cond $X=2.07 $Y=0.93
+ $X2=2.07 $Y2=3.075
r216 18 51 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.71 $Y=0.855
+ $X2=1.635 $Y2=0.855
r217 17 52 5.30422 $w=1.5e-07 $l=1.07e-07 $layer=POLY_cond $X=1.995 $Y=0.855
+ $X2=2.102 $Y2=0.855
r218 17 18 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.995 $Y=0.855
+ $X2=1.71 $Y2=0.855
r219 14 51 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.635 $Y=0.78
+ $X2=1.635 $Y2=0.855
r220 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.635 $Y=0.78
+ $X2=1.635 $Y2=0.495
r221 11 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.275 $Y=0.78
+ $X2=1.275 $Y2=0.855
r222 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.275 $Y=0.78
+ $X2=1.275 $Y2=0.495
r223 7 46 64.9888 $w=2.67e-07 $l=4.24264e-07 $layer=POLY_cond $X=1.19 $Y=1.69
+ $X2=1.33 $Y2=1.33
r224 7 9 212.428 $w=2.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.19 $Y=1.69
+ $X2=1.19 $Y2=2.545
r225 2 71 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.25
+ $Y=2.045 $X2=0.395 $Y2=2.19
r226 2 63 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.25
+ $Y=2.045 $X2=0.395 $Y2=2.9
r227 1 57 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.27 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%A_1583_285# 1 2 9 13 17 19 21 25 27 33 34
+ 36 37 38 40 45 46 50 56
c111 33 0 7.9537e-20 $X=8.68 $Y=1.59
c112 27 0 1.2552e-19 $X=8.49 $Y=1.59
r113 58 59 8.23016 $w=2.52e-07 $l=1.7e-07 $layer=LI1_cond $X=9.555 $Y=1.67
+ $X2=9.555 $Y2=1.84
r114 54 56 6.54089 $w=3.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.42 $Y=0.54
+ $X2=9.63 $Y2=0.54
r115 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.25
+ $Y=1.25 $X2=10.25 $Y2=1.25
r116 48 50 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.25 $Y=1.585
+ $X2=10.25 $Y2=1.25
r117 47 58 3.04159 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.72 $Y=1.67
+ $X2=9.555 $Y2=1.67
r118 46 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.085 $Y=1.67
+ $X2=10.25 $Y2=1.585
r119 46 47 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=10.085 $Y=1.67
+ $X2=9.72 $Y2=1.67
r120 45 58 5.41258 $w=2.52e-07 $l=1.16619e-07 $layer=LI1_cond $X=9.63 $Y=1.585
+ $X2=9.555 $Y2=1.67
r121 44 56 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=9.63 $Y=0.725
+ $X2=9.63 $Y2=0.54
r122 44 45 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=9.63 $Y=0.725
+ $X2=9.63 $Y2=1.585
r123 40 42 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=9.555 $Y=2.06
+ $X2=9.555 $Y2=2.77
r124 38 59 3.85419 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.555 $Y=1.925
+ $X2=9.555 $Y2=1.84
r125 38 40 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=9.555 $Y=1.925
+ $X2=9.555 $Y2=2.06
r126 36 59 3.04159 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.39 $Y=1.84
+ $X2=9.555 $Y2=1.84
r127 36 37 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=9.39 $Y=1.84
+ $X2=8.845 $Y2=1.84
r128 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.68
+ $Y=1.59 $X2=8.68 $Y2=1.59
r129 31 37 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=8.69 $Y=1.755
+ $X2=8.845 $Y2=1.84
r130 31 33 6.13397 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=8.69 $Y=1.755
+ $X2=8.69 $Y2=1.59
r131 28 30 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=8.04 $Y=1.59
+ $X2=8.415 $Y2=1.59
r132 27 34 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=8.49 $Y=1.59
+ $X2=8.68 $Y2=1.59
r133 27 30 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.49 $Y=1.59
+ $X2=8.415 $Y2=1.59
r134 23 51 31.7333 $w=2.68e-07 $l=2.68093e-07 $layer=POLY_cond $X=10.555
+ $Y=1.085 $X2=10.357 $Y2=1.25
r135 23 25 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=10.555 $Y=1.085
+ $X2=10.555 $Y2=0.67
r136 19 51 59.2023 $w=5.37e-07 $l=5.69838e-07 $layer=POLY_cond $X=10.495
+ $Y=1.755 $X2=10.357 $Y2=1.25
r137 19 21 180.129 $w=2.5e-07 $l=7.25e-07 $layer=POLY_cond $X=10.495 $Y=1.755
+ $X2=10.495 $Y2=2.48
r138 15 51 31.7333 $w=2.68e-07 $l=2.32282e-07 $layer=POLY_cond $X=10.195
+ $Y=1.085 $X2=10.357 $Y2=1.25
r139 15 17 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=10.195 $Y=1.085
+ $X2=10.195 $Y2=0.67
r140 11 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.415 $Y=1.425
+ $X2=8.415 $Y2=1.59
r141 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.415 $Y=1.425
+ $X2=8.415 $Y2=0.585
r142 7 28 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.04 $Y=1.755
+ $X2=8.04 $Y2=1.59
r143 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.04 $Y=1.755
+ $X2=8.04 $Y2=2.415
r144 2 42 400 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=9.335
+ $Y=1.915 $X2=9.555 $Y2=2.77
r145 2 40 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=9.335
+ $Y=1.915 $X2=9.555 $Y2=2.06
r146 1 54 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.28
+ $Y=0.375 $X2=9.42 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%A_1429_383# 1 2 7 9 12 14 16 21 24 27 29 34
+ 36 37 42 43 45 46
c94 36 0 8.68493e-20 $X=8.27 $Y=2.075
c95 21 0 7.9537e-20 $X=9.22 $Y=1.055
r96 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.22
+ $Y=1.07 $X2=9.22 $Y2=1.07
r97 38 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=1.08
+ $X2=8.27 $Y2=1.08
r98 37 45 4.60557 $w=1.7e-07 $l=1.76068e-07 $layer=LI1_cond $X=9.055 $Y=1.08
+ $X2=9.21 $Y2=1.035
r99 37 38 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=9.055 $Y=1.08
+ $X2=8.355 $Y2=1.08
r100 35 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.27 $Y=1.165
+ $X2=8.27 $Y2=1.08
r101 35 36 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=8.27 $Y=1.165
+ $X2=8.27 $Y2=2.075
r102 34 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.27 $Y=0.995
+ $X2=8.27 $Y2=1.08
r103 33 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.27 $Y=0.685
+ $X2=8.27 $Y2=0.995
r104 29 33 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.185 $Y=0.52
+ $X2=8.27 $Y2=0.685
r105 29 31 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=8.185 $Y=0.52
+ $X2=7.84 $Y2=0.52
r106 28 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=2.16
+ $X2=7.285 $Y2=2.16
r107 27 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.185 $Y=2.16
+ $X2=8.27 $Y2=2.075
r108 27 28 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=8.185 $Y=2.16
+ $X2=7.45 $Y2=2.16
r109 23 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.22 $Y=1.41
+ $X2=9.22 $Y2=1.07
r110 23 24 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.22 $Y=1.41
+ $X2=9.22 $Y2=1.575
r111 21 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.22 $Y=1.055
+ $X2=9.22 $Y2=1.07
r112 19 21 7.69149 $w=1.5e-07 $l=1.5e-08 $layer=POLY_cond $X=9.205 $Y=0.98
+ $X2=9.22 $Y2=0.98
r113 17 19 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=8.845 $Y=0.98
+ $X2=9.205 $Y2=0.98
r114 14 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.205 $Y=0.905
+ $X2=9.205 $Y2=0.98
r115 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.205 $Y=0.905
+ $X2=9.205 $Y2=0.585
r116 12 24 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=9.21 $Y=2.415
+ $X2=9.21 $Y2=1.575
r117 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.845 $Y=0.905
+ $X2=8.845 $Y2=0.98
r118 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.845 $Y=0.905
+ $X2=8.845 $Y2=0.585
r119 2 42 300 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_PDIFF $count=2 $X=7.145
+ $Y=1.915 $X2=7.285 $Y2=2.24
r120 1 31 182 $w=1.7e-07 $l=3.13129e-07 $layer=licon1_NDIFF $count=1 $X=7.575
+ $Y=0.625 $X2=7.84 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%VPWR 1 2 3 4 5 18 24 28 32 36 41 42 44 45
+ 47 48 49 55 62 84 85 88 91
c92 28 0 1.07714e-19 $X=5.525 $Y=2.4
r93 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r94 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r95 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r96 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r97 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r98 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.88 $Y=3.33 $X2=9.84
+ $Y2=3.33
r99 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r100 76 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r101 75 76 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r102 73 76 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6 $Y=3.33 $X2=8.4
+ $Y2=3.33
r103 72 75 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=8.4
+ $Y2=3.33
r104 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r105 70 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.69 $Y=3.33
+ $X2=5.525 $Y2=3.33
r106 70 72 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.69 $Y=3.33 $X2=6
+ $Y2=3.33
r107 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 66 69 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 66 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 65 68 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r111 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 63 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=3.33
+ $X2=2.705 $Y2=3.33
r113 63 65 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.87 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 62 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.36 $Y=3.33
+ $X2=5.525 $Y2=3.33
r115 62 68 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.36 $Y=3.33
+ $X2=5.04 $Y2=3.33
r116 61 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r120 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r121 55 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=3.33
+ $X2=2.705 $Y2=3.33
r122 55 60 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.54 $Y=3.33
+ $X2=2.16 $Y2=3.33
r123 53 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 49 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r126 49 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r127 49 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 47 81 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=10.065 $Y=3.33
+ $X2=9.84 $Y2=3.33
r129 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.065 $Y=3.33
+ $X2=10.23 $Y2=3.33
r130 46 84 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=10.395 $Y=3.33
+ $X2=10.8 $Y2=3.33
r131 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.395 $Y=3.33
+ $X2=10.23 $Y2=3.33
r132 44 75 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.4 $Y2=3.33
r133 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.7 $Y2=3.33
r134 43 78 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=8.865 $Y=3.33
+ $X2=8.88 $Y2=3.33
r135 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.865 $Y=3.33
+ $X2=8.7 $Y2=3.33
r136 41 52 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.76 $Y=3.33 $X2=0.72
+ $Y2=3.33
r137 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=3.33
+ $X2=0.925 $Y2=3.33
r138 40 57 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=1.2 $Y2=3.33
r139 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.925 $Y2=3.33
r140 36 39 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=10.23 $Y=2.125
+ $X2=10.23 $Y2=2.835
r141 34 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.23 $Y=3.245
+ $X2=10.23 $Y2=3.33
r142 34 39 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.23 $Y=3.245
+ $X2=10.23 $Y2=2.835
r143 30 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.7 $Y=3.245 $X2=8.7
+ $Y2=3.33
r144 30 32 34.0495 $w=3.28e-07 $l=9.75e-07 $layer=LI1_cond $X=8.7 $Y=3.245
+ $X2=8.7 $Y2=2.27
r145 26 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.525 $Y=3.245
+ $X2=5.525 $Y2=3.33
r146 26 28 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=5.525 $Y=3.245
+ $X2=5.525 $Y2=2.4
r147 22 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=3.245
+ $X2=2.705 $Y2=3.33
r148 22 24 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=2.705 $Y=3.245
+ $X2=2.705 $Y2=2.195
r149 18 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.925 $Y=2.19
+ $X2=0.925 $Y2=2.9
r150 16 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=3.33
r151 16 21 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.925 $Y=3.245
+ $X2=0.925 $Y2=2.9
r152 5 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.085
+ $Y=1.98 $X2=10.23 $Y2=2.835
r153 5 36 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.085
+ $Y=1.98 $X2=10.23 $Y2=2.125
r154 4 32 300 $w=1.7e-07 $l=6.90036e-07 $layer=licon1_PDIFF $count=2 $X=8.165
+ $Y=1.915 $X2=8.7 $Y2=2.27
r155 3 28 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=1.705 $X2=5.525 $Y2=2.4
r156 2 24 300 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_PDIFF $count=2 $X=2.56
+ $Y=1.705 $X2=2.705 $Y2=2.195
r157 1 21 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.785
+ $Y=2.045 $X2=0.925 $Y2=2.9
r158 1 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.785
+ $Y=2.045 $X2=0.925 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%A_629_125# 1 2 9 13 14 15 18 20
c42 15 0 9.46556e-20 $X=3.825 $Y=1.81
c43 14 0 1.17622e-19 $X=3.53 $Y=0.95
r44 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.91 $Y=1.035
+ $X2=3.91 $Y2=1.725
r45 16 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=1.81
+ $X2=3.45 $Y2=1.81
r46 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.825 $Y=1.81
+ $X2=3.91 $Y2=1.725
r47 15 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.825 $Y=1.81
+ $X2=3.615 $Y2=1.81
r48 13 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.825 $Y=0.95
+ $X2=3.91 $Y2=1.035
r49 13 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.825 $Y=0.95
+ $X2=3.53 $Y2=0.95
r50 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.365 $Y=0.865
+ $X2=3.53 $Y2=0.95
r51 7 9 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.365 $Y=0.865
+ $X2=3.365 $Y2=0.705
r52 2 20 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=3.175
+ $Y=1.705 $X2=3.45 $Y2=1.89
r53 1 9 182 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.625 $X2=3.365 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%Q 1 2 9 13 14 15 16 34
r18 22 34 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=10.765 $Y=1.61
+ $X2=10.765 $Y2=1.665
r19 16 36 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=10.765 $Y=1.68
+ $X2=10.765 $Y2=1.78
r20 16 34 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=10.765 $Y=1.68
+ $X2=10.765 $Y2=1.665
r21 16 22 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=10.765 $Y=1.595
+ $X2=10.765 $Y2=1.61
r22 15 16 10.1686 $w=3.38e-07 $l=3e-07 $layer=LI1_cond $X=10.765 $Y=1.295
+ $X2=10.765 $Y2=1.595
r23 14 15 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.765 $Y=0.925
+ $X2=10.765 $Y2=1.295
r24 14 27 8.64332 $w=3.38e-07 $l=2.55e-07 $layer=LI1_cond $X=10.765 $Y=0.925
+ $X2=10.765 $Y2=0.67
r25 13 27 3.89797 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=10.765 $Y=0.555
+ $X2=10.765 $Y2=0.67
r26 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=10.76 $Y=2.125
+ $X2=10.76 $Y2=2.835
r27 9 36 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=10.76 $Y=2.125
+ $X2=10.76 $Y2=1.78
r28 2 11 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.98 $X2=10.76 $Y2=2.835
r29 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.98 $X2=10.76 $Y2=2.125
r30 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.63
+ $Y=0.46 $X2=10.77 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_LP%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 43 44 45 47 56 77 78 81 84
c121 37 0 1.67093e-19 $X=2.26 $Y=0
r122 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r123 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r124 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r125 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r126 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r127 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r128 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r129 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r130 69 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r131 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r132 66 69 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r133 66 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r134 65 68 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r135 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r136 63 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.57 $Y=0 $X2=6.445
+ $Y2=0
r137 63 65 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=6.57 $Y=0 $X2=6.96
+ $Y2=0
r138 62 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r139 61 62 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6 $Y=0 $X2=6
+ $Y2=0
r140 58 61 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=6
+ $Y2=0
r141 58 59 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r142 56 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.32 $Y=0 $X2=6.445
+ $Y2=0
r143 56 61 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.32 $Y=0 $X2=6
+ $Y2=0
r144 55 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r145 55 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r146 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r147 52 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.06
+ $Y2=0
r148 52 54 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=2.16
+ $Y2=0
r149 50 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r150 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r151 47 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.06
+ $Y2=0
r152 47 49 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.72 $Y2=0
r153 45 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r154 45 59 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=2.64 $Y2=0
r155 43 74 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=9.895 $Y=0 $X2=9.84
+ $Y2=0
r156 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.895 $Y=0
+ $X2=10.02 $Y2=0
r157 42 77 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=10.145 $Y=0
+ $X2=10.8 $Y2=0
r158 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.145 $Y=0
+ $X2=10.02 $Y2=0
r159 40 68 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.545 $Y=0 $X2=8.4
+ $Y2=0
r160 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.545 $Y=0 $X2=8.67
+ $Y2=0
r161 39 71 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.88
+ $Y2=0
r162 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.67
+ $Y2=0
r163 37 54 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.16
+ $Y2=0
r164 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.425
+ $Y2=0
r165 36 58 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.64
+ $Y2=0
r166 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.425
+ $Y2=0
r167 32 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.02 $Y=0.085
+ $X2=10.02 $Y2=0
r168 32 34 26.9672 $w=2.48e-07 $l=5.85e-07 $layer=LI1_cond $X=10.02 $Y=0.085
+ $X2=10.02 $Y2=0.67
r169 28 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.67 $Y=0.085
+ $X2=8.67 $Y2=0
r170 28 30 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=8.67 $Y=0.085
+ $X2=8.67 $Y2=0.585
r171 24 84 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.445 $Y=0.085
+ $X2=6.445 $Y2=0
r172 24 26 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=6.445 $Y=0.085
+ $X2=6.445 $Y2=0.52
r173 20 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0
r174 20 22 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0.795
r175 16 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=0.085
+ $X2=1.06 $Y2=0
r176 16 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.06 $Y=0.085
+ $X2=1.06 $Y2=0.455
r177 5 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=9.835
+ $Y=0.46 $X2=9.98 $Y2=0.67
r178 4 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.49
+ $Y=0.375 $X2=8.63 $Y2=0.585
r179 3 26 182 $w=1.7e-07 $l=1.28143e-06 $layer=licon1_NDIFF $count=1 $X=5.175
+ $Y=0.625 $X2=6.405 $Y2=0.52
r180 2 22 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=2.285
+ $Y=0.625 $X2=2.425 $Y2=0.795
r181 1 18 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=0.92
+ $Y=0.285 $X2=1.06 $Y2=0.455
.ends

