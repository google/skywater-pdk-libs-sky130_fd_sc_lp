* File: sky130_fd_sc_lp__o21ai_m.pxi.spice
* Created: Fri Aug 28 11:05:20 2020
* 
x_PM_SKY130_FD_SC_LP__O21AI_M%A1 N_A1_c_44_n N_A1_M1004_g N_A1_M1005_g
+ N_A1_c_47_n A1 A1 A1 N_A1_c_48_n N_A1_c_49_n PM_SKY130_FD_SC_LP__O21AI_M%A1
x_PM_SKY130_FD_SC_LP__O21AI_M%A2 N_A2_M1003_g N_A2_M1000_g N_A2_c_76_n A2 A2
+ N_A2_c_78_n PM_SKY130_FD_SC_LP__O21AI_M%A2
x_PM_SKY130_FD_SC_LP__O21AI_M%B1 N_B1_M1002_g N_B1_M1001_g N_B1_c_109_n
+ N_B1_c_110_n B1 B1 N_B1_c_111_n N_B1_c_112_n PM_SKY130_FD_SC_LP__O21AI_M%B1
x_PM_SKY130_FD_SC_LP__O21AI_M%VPWR N_VPWR_M1005_s N_VPWR_M1001_d N_VPWR_c_144_n
+ N_VPWR_c_145_n N_VPWR_c_146_n N_VPWR_c_147_n VPWR N_VPWR_c_148_n
+ N_VPWR_c_143_n PM_SKY130_FD_SC_LP__O21AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O21AI_M%Y N_Y_M1002_d N_Y_M1003_d N_Y_c_169_n N_Y_c_170_n
+ N_Y_c_172_n Y Y PM_SKY130_FD_SC_LP__O21AI_M%Y
x_PM_SKY130_FD_SC_LP__O21AI_M%A_27_51# N_A_27_51#_M1004_s N_A_27_51#_M1000_d
+ N_A_27_51#_c_199_n N_A_27_51#_c_200_n N_A_27_51#_c_201_n N_A_27_51#_c_209_n
+ PM_SKY130_FD_SC_LP__O21AI_M%A_27_51#
x_PM_SKY130_FD_SC_LP__O21AI_M%VGND N_VGND_M1004_d N_VGND_c_222_n VGND
+ N_VGND_c_223_n N_VGND_c_224_n N_VGND_c_225_n N_VGND_c_226_n
+ PM_SKY130_FD_SC_LP__O21AI_M%VGND
cc_1 VNB N_A1_c_44_n 0.0285971f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.413
cc_2 VNB N_A1_M1004_g 0.0317798f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.465
cc_3 VNB N_A1_M1005_g 0.00184732f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.38
cc_4 VNB N_A1_c_47_n 0.0326676f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.625
cc_5 VNB N_A1_c_48_n 0.0326498f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_6 VNB N_A1_c_49_n 0.00111806f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_7 VNB N_A2_M1000_g 0.0606645f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.625
cc_8 VNB N_B1_M1002_g 0.0370784f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.955
cc_9 VNB N_B1_c_109_n 0.0236573f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.625
cc_10 VNB N_B1_c_110_n 0.00489944f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_B1_c_111_n 0.0169359f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.12
cc_12 VNB N_B1_c_112_n 0.00905268f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.12
cc_13 VNB N_VPWR_c_143_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_Y_c_169_n 0.048869f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.38
cc_15 VNB N_Y_c_170_n 0.0104829f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_A_27_51#_c_199_n 4.08405e-19 $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.38
cc_17 VNB N_A_27_51#_c_200_n 0.0216577f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.625
cc_18 VNB N_A_27_51#_c_201_n 0.00846785f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_VGND_c_222_n 0.00100404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_223_n 0.0157759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_224_n 0.0301611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_225_n 0.13937f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.12
cc_23 VNB N_VGND_c_226_n 0.00460801f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=0.955
cc_24 VPB N_A1_M1005_g 0.0457475f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.38
cc_25 VPB N_A1_c_49_n 0.0212435f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_26 VPB N_A2_M1003_g 0.0136488f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.465
cc_27 VPB N_A2_M1000_g 0.0138207f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.625
cc_28 VPB N_A2_c_76_n 0.013027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB A2 0.0136243f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_30 VPB N_A2_c_78_n 0.0433373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_B1_M1001_g 0.03964f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.625
cc_32 VPB N_B1_c_110_n 0.0115915f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_33 VPB N_B1_c_112_n 0.00287993f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.12
cc_34 VPB N_VPWR_c_144_n 0.0115529f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.625
cc_35 VPB N_VPWR_c_145_n 0.0422583f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.38
cc_36 VPB N_VPWR_c_146_n 0.0133915f $X=-0.19 $Y=1.655 $X2=0.337 $Y2=1.625
cc_37 VPB N_VPWR_c_147_n 0.0308268f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_38 VPB N_VPWR_c_148_n 0.0283973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_143_n 0.064695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_Y_c_169_n 0.013436f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.38
cc_41 VPB N_Y_c_172_n 0.0212399f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_42 VPB Y 0.0141723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 N_A1_M1004_g N_A2_M1000_g 0.0660085f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_44 N_A1_c_49_n N_A2_M1000_g 0.00325925f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_45 N_A1_M1005_g N_A2_c_76_n 0.0479292f $X=0.475 $Y=2.38 $X2=0 $Y2=0
cc_46 N_A1_c_49_n N_A2_c_76_n 2.77616e-19 $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_47 N_A1_M1005_g A2 2.13366e-19 $X=0.475 $Y=2.38 $X2=0 $Y2=0
cc_48 N_A1_c_49_n N_B1_c_112_n 0.0188023f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_49 N_A1_M1005_g N_VPWR_c_145_n 0.00905675f $X=0.475 $Y=2.38 $X2=0 $Y2=0
cc_50 N_A1_c_49_n N_VPWR_c_145_n 0.0203964f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_51 N_A1_M1005_g N_VPWR_c_148_n 0.00298903f $X=0.475 $Y=2.38 $X2=0 $Y2=0
cc_52 N_A1_M1005_g N_VPWR_c_143_n 0.00368577f $X=0.475 $Y=2.38 $X2=0 $Y2=0
cc_53 N_A1_M1005_g Y 0.00869853f $X=0.475 $Y=2.38 $X2=0 $Y2=0
cc_54 N_A1_c_49_n Y 0.0152592f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_55 N_A1_M1004_g N_A_27_51#_c_199_n 3.52891e-19 $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_56 N_A1_M1004_g N_A_27_51#_c_200_n 0.0159169f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_57 N_A1_c_48_n N_A_27_51#_c_200_n 0.00155403f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_58 N_A1_c_49_n N_A_27_51#_c_200_n 0.00809969f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_59 N_A1_c_48_n N_A_27_51#_c_201_n 0.00552095f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_60 N_A1_c_49_n N_A_27_51#_c_201_n 0.0158108f $X=0.29 $Y=1.12 $X2=0 $Y2=0
cc_61 N_A1_M1004_g N_VGND_c_222_n 0.011607f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_62 N_A1_M1004_g N_VGND_c_223_n 0.00345529f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_63 N_A1_M1004_g N_VGND_c_225_n 0.00505351f $X=0.475 $Y=0.465 $X2=0 $Y2=0
cc_64 N_A2_M1000_g N_B1_M1002_g 0.0280157f $X=0.905 $Y=0.465 $X2=0 $Y2=0
cc_65 N_A2_M1003_g N_B1_M1001_g 0.0134345f $X=0.835 $Y=2.38 $X2=0 $Y2=0
cc_66 N_A2_M1000_g N_B1_M1001_g 0.0124055f $X=0.905 $Y=0.465 $X2=0 $Y2=0
cc_67 A2 N_B1_M1001_g 3.14667e-19 $X=1.115 $Y=2.69 $X2=0 $Y2=0
cc_68 N_A2_M1000_g N_B1_c_111_n 0.0331774f $X=0.905 $Y=0.465 $X2=0 $Y2=0
cc_69 N_A2_M1000_g N_B1_c_112_n 0.00804396f $X=0.905 $Y=0.465 $X2=0 $Y2=0
cc_70 N_A2_M1003_g N_VPWR_c_145_n 0.00270784f $X=0.835 $Y=2.38 $X2=0 $Y2=0
cc_71 A2 N_VPWR_c_145_n 0.0232674f $X=1.115 $Y=2.69 $X2=0 $Y2=0
cc_72 N_A2_c_78_n N_VPWR_c_145_n 0.00274674f $X=0.925 $Y=2.915 $X2=0 $Y2=0
cc_73 A2 N_VPWR_c_147_n 0.0234427f $X=1.115 $Y=2.69 $X2=0 $Y2=0
cc_74 N_A2_c_78_n N_VPWR_c_147_n 0.00357657f $X=0.925 $Y=2.915 $X2=0 $Y2=0
cc_75 A2 N_VPWR_c_148_n 0.0287548f $X=1.115 $Y=2.69 $X2=0 $Y2=0
cc_76 N_A2_c_78_n N_VPWR_c_148_n 0.00811075f $X=0.925 $Y=2.915 $X2=0 $Y2=0
cc_77 A2 N_VPWR_c_143_n 0.0234443f $X=1.115 $Y=2.69 $X2=0 $Y2=0
cc_78 N_A2_c_78_n N_VPWR_c_143_n 0.0112003f $X=0.925 $Y=2.915 $X2=0 $Y2=0
cc_79 N_A2_M1003_g Y 0.0119051f $X=0.835 $Y=2.38 $X2=0 $Y2=0
cc_80 N_A2_c_76_n Y 0.0168446f $X=0.87 $Y=2.06 $X2=0 $Y2=0
cc_81 A2 Y 0.0388131f $X=1.115 $Y=2.69 $X2=0 $Y2=0
cc_82 N_A2_c_78_n Y 8.54323e-19 $X=0.925 $Y=2.915 $X2=0 $Y2=0
cc_83 N_A2_M1000_g N_A_27_51#_c_200_n 0.0159066f $X=0.905 $Y=0.465 $X2=0 $Y2=0
cc_84 N_A2_M1000_g N_A_27_51#_c_209_n 2.03427e-19 $X=0.905 $Y=0.465 $X2=0 $Y2=0
cc_85 N_A2_M1000_g N_VGND_c_222_n 0.00851777f $X=0.905 $Y=0.465 $X2=0 $Y2=0
cc_86 N_A2_M1000_g N_VGND_c_224_n 0.00345529f $X=0.905 $Y=0.465 $X2=0 $Y2=0
cc_87 N_A2_M1000_g N_VGND_c_225_n 0.00421603f $X=0.905 $Y=0.465 $X2=0 $Y2=0
cc_88 N_B1_M1001_g N_VPWR_c_147_n 0.00475733f $X=1.375 $Y=2.38 $X2=0 $Y2=0
cc_89 N_B1_M1001_g N_VPWR_c_148_n 0.00359559f $X=1.375 $Y=2.38 $X2=0 $Y2=0
cc_90 N_B1_M1001_g N_VPWR_c_143_n 0.00438782f $X=1.375 $Y=2.38 $X2=0 $Y2=0
cc_91 N_B1_M1002_g N_Y_c_169_n 0.0109037f $X=1.335 $Y=0.465 $X2=0 $Y2=0
cc_92 N_B1_M1001_g N_Y_c_169_n 0.00593338f $X=1.375 $Y=2.38 $X2=0 $Y2=0
cc_93 N_B1_c_111_n N_Y_c_169_n 0.0163648f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_94 N_B1_c_112_n N_Y_c_169_n 0.048424f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_95 N_B1_M1002_g N_Y_c_170_n 0.00187228f $X=1.335 $Y=0.465 $X2=0 $Y2=0
cc_96 N_B1_c_111_n N_Y_c_170_n 0.0026968f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_97 N_B1_c_112_n N_Y_c_170_n 0.00133188f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_98 N_B1_M1001_g N_Y_c_172_n 0.0166825f $X=1.375 $Y=2.38 $X2=0 $Y2=0
cc_99 N_B1_c_110_n N_Y_c_172_n 0.00342508f $X=1.385 $Y=1.75 $X2=0 $Y2=0
cc_100 N_B1_M1001_g Y 0.0042387f $X=1.375 $Y=2.38 $X2=0 $Y2=0
cc_101 N_B1_c_110_n Y 5.93163e-19 $X=1.385 $Y=1.75 $X2=0 $Y2=0
cc_102 N_B1_c_112_n Y 0.0280456f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_103 N_B1_M1002_g N_A_27_51#_c_200_n 0.00227506f $X=1.335 $Y=0.465 $X2=0 $Y2=0
cc_104 N_B1_c_112_n N_A_27_51#_c_200_n 0.00814522f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_105 N_B1_M1002_g N_VGND_c_222_n 0.00148754f $X=1.335 $Y=0.465 $X2=0 $Y2=0
cc_106 N_B1_M1002_g N_VGND_c_224_n 0.00558812f $X=1.335 $Y=0.465 $X2=0 $Y2=0
cc_107 N_B1_M1002_g N_VGND_c_225_n 0.0115469f $X=1.335 $Y=0.465 $X2=0 $Y2=0
cc_108 N_VPWR_c_147_n N_Y_c_172_n 0.0159014f $X=1.59 $Y=2.445 $X2=0 $Y2=0
cc_109 N_VPWR_c_145_n Y 0.0097157f $X=0.26 $Y=2.445 $X2=0 $Y2=0
cc_110 A_110_434# Y 0.0043102f $X=0.55 $Y=2.17 $X2=1.115 $Y2=1.95
cc_111 N_Y_c_169_n N_A_27_51#_c_200_n 0.00756459f $X=1.735 $Y=1.93 $X2=0 $Y2=0
cc_112 N_Y_c_169_n N_A_27_51#_c_209_n 0.00109941f $X=1.735 $Y=1.93 $X2=0 $Y2=0
cc_113 N_Y_c_170_n N_VGND_c_224_n 0.0120436f $X=1.735 $Y=0.53 $X2=0 $Y2=0
cc_114 N_Y_c_170_n N_VGND_c_225_n 0.0139713f $X=1.735 $Y=0.53 $X2=0 $Y2=0
cc_115 N_A_27_51#_c_200_n N_VGND_c_222_n 0.0193682f $X=1.035 $Y=0.77 $X2=0 $Y2=0
cc_116 N_A_27_51#_c_199_n N_VGND_c_223_n 0.00750141f $X=0.26 $Y=0.53 $X2=0 $Y2=0
cc_117 N_A_27_51#_c_200_n N_VGND_c_223_n 0.00271048f $X=1.035 $Y=0.77 $X2=0
+ $Y2=0
cc_118 N_A_27_51#_c_200_n N_VGND_c_224_n 0.00271048f $X=1.035 $Y=0.77 $X2=0
+ $Y2=0
cc_119 N_A_27_51#_c_209_n N_VGND_c_224_n 0.00711705f $X=1.12 $Y=0.53 $X2=0 $Y2=0
cc_120 N_A_27_51#_c_199_n N_VGND_c_225_n 0.00679726f $X=0.26 $Y=0.53 $X2=0 $Y2=0
cc_121 N_A_27_51#_c_200_n N_VGND_c_225_n 0.0100561f $X=1.035 $Y=0.77 $X2=0 $Y2=0
cc_122 N_A_27_51#_c_209_n N_VGND_c_225_n 0.00679726f $X=1.12 $Y=0.53 $X2=0 $Y2=0
