* File: sky130_fd_sc_lp__maj3_4.spice
* Created: Fri Aug 28 10:43:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__maj3_4.pex.spice"
.subckt sky130_fd_sc_lp__maj3_4  VNB VPB C A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C	C
* VPB	VPB
* VNB	VNB
MM1002 A_154_47# N_C_M1002_g N_A_65_367#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.2394 PD=1.08 PS=2.25 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.3 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g A_154_47# VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1008 PD=1.12 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75000.6 SB=75003.9
+ A=0.126 P=1.98 MULT=1
MM1010 A_318_47# N_A_M1010_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.1176 PD=1.08 PS=1.12 NRD=9.276 NRS=0 M=1 R=5.6 SA=75001 SB=75003.5
+ A=0.126 P=1.98 MULT=1
MM1011 N_A_65_367#_M1011_d N_B_M1011_g A_318_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1008 PD=1.12 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75001.4
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1017 A_482_47# N_B_M1017_g N_A_65_367#_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.1176 PD=1.08 PS=1.12 NRD=9.276 NRS=0 M=1 R=5.6 SA=75001.8
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1016_d N_C_M1016_g A_482_47# VNB NSHORT L=0.15 W=0.84 AD=0.2121
+ AS=0.1008 PD=1.345 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75002.2 SB=75002.3
+ A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1016_d N_A_65_367#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2121 AS=0.1176 PD=1.345 PS=1.12 NRD=32.136 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_65_367#_M1004_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1323 AS=0.1176 PD=1.155 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1004_d N_A_65_367#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1323 AS=0.1344 PD=1.155 PS=1.16 NRD=4.992 NRS=0 M=1 R=5.6 SA=75003.8
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A_65_367#_M1012_g N_X_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.273 AS=0.1344 PD=2.33 PS=1.16 NRD=5.712 NRS=5.712 M=1 R=5.6 SA=75004.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1014 A_154_367# N_C_M1014_g N_A_65_367#_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.3717 PD=1.5 PS=3.11 NRD=10.1455 NRS=1.5563 M=1 R=8.4 SA=75000.2
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_154_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.1764
+ AS=0.1512 PD=1.54 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75000.6 SB=75003.9
+ A=0.189 P=2.82 MULT=1
MM1008 A_318_367# N_A_M1008_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1512
+ AS=0.1764 PD=1.5 PS=1.54 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75001 SB=75003.4
+ A=0.189 P=2.82 MULT=1
MM1018 N_A_65_367#_M1018_d N_B_M1018_g A_318_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1512 PD=1.54 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75001.4
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1009 A_482_367# N_B_M1009_g N_A_65_367#_M1018_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.1764 PD=1.5 PS=1.54 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1019_d N_C_M1019_g A_482_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2646
+ AS=0.1512 PD=1.68 PS=1.5 NRD=9.3772 NRS=10.1455 M=1 R=8.4 SA=75002.2
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1019_d N_A_65_367#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.1764 PD=1.68 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A_65_367#_M1007_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2772 AS=0.1764 PD=1.7 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1007_d N_A_65_367#_M1013_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2772 AS=0.1764 PD=1.7 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4 SA=75003.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1015 N_VPWR_M1015_d N_A_65_367#_M1015_g N_X_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.5559 P=15.05
*
.include "sky130_fd_sc_lp__maj3_4.pxi.spice"
*
.ends
*
*
