# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__lsbufiso0p_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__lsbufiso0p_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  6.660000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.678000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 1.530000 1.245000 2.135000 ;
        RECT 1.075000 2.135000 1.245000 2.775000 ;
        RECT 1.075000 2.775000 1.645000 3.075000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.978000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.835000 4.505000 3.420000 4.910000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.714400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.285000 3.590000 4.565000 4.320000 ;
        RECT 4.285000 4.320000 6.145000 4.490000 ;
        RECT 5.815000 3.585000 6.145000 4.320000 ;
        RECT 5.815000 4.490000 6.145000 6.405000 ;
    END
  END X
  PIN DESTPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 6.575000 6.720000 6.745000 ;
        RECT 3.570000 5.420000 3.740000 6.575000 ;
        RECT 5.040000 5.420000 5.355000 6.575000 ;
      LAYER mcon ;
        RECT 0.155000 6.575000 0.325000 6.745000 ;
        RECT 0.635000 6.575000 0.805000 6.745000 ;
        RECT 1.115000 6.575000 1.285000 6.745000 ;
        RECT 1.595000 6.575000 1.765000 6.745000 ;
        RECT 2.075000 6.575000 2.245000 6.745000 ;
        RECT 2.555000 6.575000 2.725000 6.745000 ;
        RECT 3.035000 6.575000 3.205000 6.745000 ;
        RECT 3.515000 6.575000 3.685000 6.745000 ;
        RECT 3.995000 6.575000 4.165000 6.745000 ;
        RECT 4.475000 6.575000 4.645000 6.745000 ;
        RECT 4.955000 6.575000 5.125000 6.745000 ;
        RECT 5.435000 6.575000 5.605000 6.745000 ;
        RECT 5.915000 6.575000 6.085000 6.745000 ;
        RECT 6.395000 6.575000 6.565000 6.745000 ;
      LAYER met1 ;
        RECT 0.000000 6.415000 6.720000 6.905000 ;
    END
  END DESTPWR
  PIN DESTVPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.090000 5.220000 0.390000 6.395000 ;
        RECT 6.330000 5.220000 6.630000 6.395000 ;
    END
  END DESTVPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 2.145000 3.415000 ;
        RECT 0.090000 1.890000 0.390000 3.245000 ;
        RECT 0.090000 3.415000 0.390000 4.770000 ;
        RECT 0.575000 2.305000 0.905000 3.245000 ;
        RECT 2.700000 3.245000 6.720000 3.415000 ;
        RECT 2.700000 3.415000 3.030000 4.240000 ;
        RECT 2.710000 2.430000 3.040000 3.245000 ;
        RECT 5.025000 3.415000 5.355000 3.880000 ;
        RECT 6.330000 1.890000 6.630000 3.245000 ;
        RECT 6.330000 3.415000 6.630000 4.770000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.075000 6.720000 3.565000 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.265000 0.390000 1.440000 ;
        RECT 6.330000 0.265000 6.630000 1.440000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.720000 0.085000 ;
        RECT 0.575000  0.085000 0.905000 1.175000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.575000 3.585000 0.855000 4.650000 ;
      RECT 0.575000 4.650000 1.690000 4.820000 ;
      RECT 0.575000 4.820000 0.830000 5.435000 ;
      RECT 0.575000 5.435000 0.925000 6.405000 ;
      RECT 1.000000 4.990000 1.330000 5.265000 ;
      RECT 1.160000 5.265000 1.330000 5.355000 ;
      RECT 1.160000 5.355000 2.325000 5.465000 ;
      RECT 1.160000 5.465000 2.485000 5.525000 ;
      RECT 1.365000 0.265000 1.715000 1.360000 ;
      RECT 1.365000 3.585000 2.485000 3.755000 ;
      RECT 1.365000 3.755000 1.645000 4.480000 ;
      RECT 1.365000 5.695000 1.695000 6.235000 ;
      RECT 1.365000 6.235000 3.390000 6.405000 ;
      RECT 1.415000 1.360000 1.715000 2.435000 ;
      RECT 1.415000 2.435000 2.145000 2.605000 ;
      RECT 1.520000 4.820000 1.690000 5.010000 ;
      RECT 1.520000 5.010000 1.930000 5.185000 ;
      RECT 1.815000 2.605000 2.145000 3.075000 ;
      RECT 2.155000 4.070000 2.485000 4.400000 ;
      RECT 2.155000 4.400000 2.325000 5.355000 ;
      RECT 2.155000 5.525000 2.485000 6.055000 ;
      RECT 2.315000 2.330000 2.530000 3.090000 ;
      RECT 2.315000 3.090000 2.485000 3.585000 ;
      RECT 2.495000 4.935000 2.665000 5.080000 ;
      RECT 2.495000 5.080000 4.160000 5.250000 ;
      RECT 2.495000 5.250000 2.745000 5.295000 ;
      RECT 3.060000 5.465000 3.390000 6.235000 ;
      RECT 3.490000 3.585000 4.080000 3.915000 ;
      RECT 3.490000 3.915000 3.820000 4.240000 ;
      RECT 3.590000 4.240000 3.815000 4.740000 ;
      RECT 3.590000 4.740000 4.530000 4.910000 ;
      RECT 3.990000 5.250000 4.160000 6.235000 ;
      RECT 3.990000 6.235000 4.870000 6.405000 ;
      RECT 4.330000 4.910000 4.530000 6.055000 ;
      RECT 4.700000 4.660000 5.580000 4.990000 ;
      RECT 4.700000 4.990000 4.870000 6.235000 ;
  END
END sky130_fd_sc_lp__lsbufiso0p_lp
