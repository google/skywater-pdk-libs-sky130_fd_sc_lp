* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_m A0 A1 S VGND VNB VPB VPWR X
X0 X a_123_269# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_441_125# a_483_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR S a_329_501# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 X a_123_269# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND S a_483_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_261_125# A1 a_123_269# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_487_501# a_483_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_123_269# A1 a_487_501# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_329_501# A0 a_123_269# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VGND S a_261_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_123_269# A0 a_441_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR S a_483_99# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
