* File: sky130_fd_sc_lp__sdfsbp_2.pex.spice
* Created: Fri Aug 28 11:29:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%SCE 2 5 9 13 17 21 25 29 30 32 33 34 35 47
+ 60
c93 30 0 2.4535e-19 $X=2.255 $Y=1.33
r94 45 47 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.72 $Y=2.01
+ $X2=0.905 $Y2=2.01
r95 42 45 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=0.475 $Y=2.01
+ $X2=0.72 $Y2=2.01
r96 35 60 13.5564 $w=2.43e-07 $l=2.65e-07 $layer=LI1_cond $X=0.72 $Y=2.367
+ $X2=0.985 $Y2=2.367
r97 34 35 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.72 $Y=2.01
+ $X2=0.72 $Y2=2.245
r98 34 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=2.01 $X2=0.72 $Y2=2.01
r99 33 34 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=2.01
r100 32 33 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.295
+ $X2=0.72 $Y2=1.665
r101 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.255
+ $Y=1.33 $X2=2.255 $Y2=1.33
r102 27 29 42.1794 $w=2.48e-07 $l=9.15e-07 $layer=LI1_cond $X=2.215 $Y=2.245
+ $X2=2.215 $Y2=1.33
r103 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.09 $Y=2.33
+ $X2=2.215 $Y2=2.245
r104 25 60 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.09 $Y=2.33
+ $X2=0.985 $Y2=2.33
r105 24 30 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.165
+ $X2=2.255 $Y2=1.33
r106 19 21 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=0.475 $Y=1.53
+ $X2=0.725 $Y2=1.53
r107 17 24 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.28 $Y=0.445
+ $X2=2.28 $Y2=1.165
r108 11 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=2.175
+ $X2=0.905 $Y2=2.01
r109 11 13 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.905 $Y=2.175
+ $X2=0.905 $Y2=2.655
r110 7 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.725 $Y=1.455
+ $X2=0.725 $Y2=1.53
r111 7 9 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.725 $Y=1.455
+ $X2=0.725 $Y2=0.445
r112 3 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=2.175
+ $X2=0.475 $Y2=2.01
r113 3 5 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.475 $Y=2.175
+ $X2=0.475 $Y2=2.655
r114 2 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.845
+ $X2=0.475 $Y2=2.01
r115 1 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.605
+ $X2=0.475 $Y2=1.53
r116 1 2 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.475 $Y=1.605
+ $X2=0.475 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%D 3 7 8 11 14 15 16 17 26 28
c54 8 0 2.5644e-19 $X=1.515 $Y=1.945
r55 26 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=0.93
+ $X2=1.715 $Y2=0.765
r56 16 17 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.657 $Y=1.295
+ $X2=1.657 $Y2=1.665
r57 15 16 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.657 $Y=0.925
+ $X2=1.657 $Y2=1.295
r58 15 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.715
+ $Y=0.93 $X2=1.715 $Y2=0.93
r59 14 15 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.657 $Y=0.555
+ $X2=1.657 $Y2=0.925
r60 13 17 6.06549 $w=2.83e-07 $l=1.5e-07 $layer=LI1_cond $X=1.657 $Y=1.815
+ $X2=1.657 $Y2=1.665
r61 11 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.98
+ $X2=1.355 $Y2=2.145
r62 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.355
+ $Y=1.98 $X2=1.355 $Y2=1.98
r63 8 13 6.83516 $w=2.6e-07 $l=1.9653e-07 $layer=LI1_cond $X=1.515 $Y=1.945
+ $X2=1.657 $Y2=1.815
r64 8 10 7.09196 $w=2.58e-07 $l=1.6e-07 $layer=LI1_cond $X=1.515 $Y=1.945
+ $X2=1.355 $Y2=1.945
r65 7 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.625 $Y=0.445
+ $X2=1.625 $Y2=0.765
r66 3 24 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.265 $Y=2.655
+ $X2=1.265 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%A_27_467# 1 2 9 11 12 15 19 22 24 29 34 35
c65 12 0 1.94743e-19 $X=1.34 $Y=1.41
r66 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.175
+ $Y=0.98 $X2=1.175 $Y2=0.98
r67 31 32 5.31754 $w=5.63e-07 $l=8.5e-08 $layer=LI1_cond $X=0.377 $Y=0.9
+ $X2=0.377 $Y2=0.985
r68 29 31 9.73798 $w=5.63e-07 $l=4.6e-07 $layer=LI1_cond $X=0.377 $Y=0.44
+ $X2=0.377 $Y2=0.9
r69 25 31 7.93092 $w=1.7e-07 $l=2.83e-07 $layer=LI1_cond $X=0.66 $Y=0.9
+ $X2=0.377 $Y2=0.9
r70 24 34 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=0.9 $X2=1.2
+ $Y2=0.9
r71 24 25 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.055 $Y=0.9
+ $X2=0.66 $Y2=0.9
r72 22 32 66.2655 $w=2.58e-07 $l=1.495e-06 $layer=LI1_cond $X=0.225 $Y=2.48
+ $X2=0.225 $Y2=0.985
r73 19 35 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.175 $Y=1.335
+ $X2=1.175 $Y2=0.98
r74 18 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=0.815
+ $X2=1.175 $Y2=0.98
r75 13 15 599.936 $w=1.5e-07 $l=1.17e-06 $layer=POLY_cond $X=1.805 $Y=1.485
+ $X2=1.805 $Y2=2.655
r76 12 19 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.34 $Y=1.41
+ $X2=1.175 $Y2=1.335
r77 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.73 $Y=1.41
+ $X2=1.805 $Y2=1.485
r78 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.73 $Y=1.41
+ $X2=1.34 $Y2=1.41
r79 9 18 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.265 $Y=0.445
+ $X2=1.265 $Y2=0.815
r80 2 22 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.335 $X2=0.26 $Y2=2.48
r81 1 29 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.385
+ $Y=0.235 $X2=0.51 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%SCD 1 3 4 5 8 11 12 14 15 16 17 21
r56 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.795
+ $Y=1.745 $X2=2.795 $Y2=1.745
r57 17 22 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=2.7 $Y=2.035 $X2=2.7
+ $Y2=1.745
r58 16 22 2.4262 $w=3.78e-07 $l=8e-08 $layer=LI1_cond $X=2.7 $Y=1.665 $X2=2.7
+ $Y2=1.745
r59 15 21 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.795 $Y=2.075
+ $X2=2.795 $Y2=1.745
r60 14 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.58
+ $X2=2.795 $Y2=1.745
r61 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.705 $Y=0.925
+ $X2=2.705 $Y2=1.58
r62 11 12 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=2.672 $Y=0.775
+ $X2=2.672 $Y2=0.925
r63 8 11 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.64 $Y=0.445 $X2=2.64
+ $Y2=0.775
r64 4 15 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.63 $Y=2.15
+ $X2=2.795 $Y2=2.075
r65 4 5 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.63 $Y=2.15 $X2=2.39
+ $Y2=2.15
r66 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.315 $Y=2.225
+ $X2=2.39 $Y2=2.15
r67 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.315 $Y=2.225
+ $X2=2.315 $Y2=2.655
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%CLK 1 3 6 8 15
c43 15 0 1.0849e-19 $X=3.28 $Y=0.93
c44 8 0 1.99828e-19 $X=3.12 $Y=0.925
r45 13 15 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=3.16 $Y=0.93
+ $X2=3.28 $Y2=0.93
r46 10 13 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.07 $Y=0.93 $X2=3.16
+ $Y2=0.93
r47 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.16
+ $Y=0.93 $X2=3.16 $Y2=0.93
r48 4 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.28 $Y=1.095
+ $X2=3.28 $Y2=0.93
r49 4 6 799.915 $w=1.5e-07 $l=1.56e-06 $layer=POLY_cond $X=3.28 $Y=1.095
+ $X2=3.28 $Y2=2.655
r50 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=0.765
+ $X2=3.07 $Y2=0.93
r51 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.07 $Y=0.765 $X2=3.07
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%A_920_73# 1 2 7 11 15 19 21 25 29 31 32 33
+ 37 38 44 45 50 59
c157 50 0 1.86354e-19 $X=8.13 $Y=1.635
c158 45 0 4.28533e-20 $X=5.21 $Y=1.65
c159 38 0 1.49559e-20 $X=9.05 $Y=1.535
c160 32 0 1.43576e-19 $X=6.43 $Y=1.635
c161 19 0 6.29478e-20 $X=9.045 $Y=0.915
r162 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.13 $Y=1.635
+ $X2=8.13 $Y2=1.94
r163 49 59 17.7787 $w=2.44e-07 $l=9e-08 $layer=POLY_cond $X=6.26 $Y=1.68
+ $X2=6.17 $Y2=1.68
r164 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.26
+ $Y=1.68 $X2=6.26 $Y2=1.68
r165 45 56 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=5.21 $Y=1.65
+ $X2=5.21 $Y2=1.77
r166 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.21
+ $Y=1.65 $X2=5.21 $Y2=1.65
r167 42 44 8.26701 $w=6.78e-07 $l=4.7e-07 $layer=LI1_cond $X=4.74 $Y=1.825
+ $X2=5.21 $Y2=1.825
r168 38 63 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.05 $Y=1.535
+ $X2=9.05 $Y2=1.625
r169 38 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.05 $Y=1.535
+ $X2=9.05 $Y2=1.37
r170 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.05
+ $Y=1.535 $X2=9.05 $Y2=1.535
r171 35 37 14.1839 $w=2.58e-07 $l=3.2e-07 $layer=LI1_cond $X=9.015 $Y=1.855
+ $X2=9.015 $Y2=1.535
r172 34 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.215 $Y=1.94
+ $X2=8.13 $Y2=1.94
r173 33 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=8.885 $Y=1.94
+ $X2=9.015 $Y2=1.855
r174 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.885 $Y=1.94
+ $X2=8.215 $Y2=1.94
r175 32 48 8.78963 $w=3.27e-07 $l=1.91181e-07 $layer=LI1_cond $X=6.43 $Y=1.635
+ $X2=6.26 $Y2=1.68
r176 31 50 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.045 $Y=1.635
+ $X2=8.13 $Y2=1.635
r177 31 32 99.5101 $w=1.78e-07 $l=1.615e-06 $layer=LI1_cond $X=8.045 $Y=1.635
+ $X2=6.43 $Y2=1.635
r178 27 42 4.97917 $w=3.3e-07 $l=3.4e-07 $layer=LI1_cond $X=4.74 $Y=1.485
+ $X2=4.74 $Y2=1.825
r179 27 29 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=4.74 $Y=1.485
+ $X2=4.74 $Y2=0.565
r180 23 25 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=9.445 $Y=1.7
+ $X2=9.445 $Y2=2.67
r181 22 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.215 $Y=1.625
+ $X2=9.05 $Y2=1.625
r182 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.37 $Y=1.625
+ $X2=9.445 $Y2=1.7
r183 21 22 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=9.37 $Y=1.625
+ $X2=9.215 $Y2=1.625
r184 19 62 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.045 $Y=0.915
+ $X2=9.045 $Y2=1.37
r185 13 59 14.1583 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.17 $Y=1.515
+ $X2=6.17 $Y2=1.68
r186 13 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.17 $Y=1.515
+ $X2=6.17 $Y2=0.805
r187 9 59 59.2623 $w=2.44e-07 $l=3.73497e-07 $layer=POLY_cond $X=5.87 $Y=1.845
+ $X2=6.17 $Y2=1.68
r188 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.87 $Y=1.845
+ $X2=5.87 $Y2=2.525
r189 8 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.375 $Y=1.77
+ $X2=5.21 $Y2=1.77
r190 7 9 21.9219 $w=2.44e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.795 $Y=1.77
+ $X2=5.87 $Y2=1.845
r191 7 8 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=5.795 $Y=1.77
+ $X2=5.375 $Y2=1.77
r192 2 42 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.945 $X2=4.74 $Y2=2.07
r193 1 29 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=4.6
+ $Y=0.365 $X2=4.74 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%A_1291_93# 1 2 7 9 10 12 14 17 21 25 30 32
+ 34 36 39 42 43 44 45 46 50
c151 34 0 1.78649e-19 $X=9.315 $Y=2.29
c152 14 0 1.96969e-19 $X=6.74 $Y=1.825
c153 10 0 2.48299e-19 $X=6.66 $Y=2.205
r154 50 52 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.83 $Y=0.95
+ $X2=8.83 $Y2=1.115
r155 46 48 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.13 $Y=2.29
+ $X2=8.13 $Y2=2.385
r156 44 45 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.79 $Y=0.837
+ $X2=7.96 $Y2=0.837
r157 41 43 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.465 $Y=2.495
+ $X2=7.63 $Y2=2.495
r158 41 42 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.465 $Y=2.495
+ $X2=7.3 $Y2=2.495
r159 38 39 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=9.4 $Y=1.2
+ $X2=9.4 $Y2=2.205
r160 37 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.915 $Y=1.115
+ $X2=8.83 $Y2=1.115
r161 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.315 $Y=1.115
+ $X2=9.4 $Y2=1.2
r162 36 37 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.315 $Y=1.115
+ $X2=8.915 $Y2=1.115
r163 35 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.215 $Y=2.29
+ $X2=8.13 $Y2=2.29
r164 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.315 $Y=2.29
+ $X2=9.4 $Y2=2.205
r165 34 35 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=9.315 $Y=2.29
+ $X2=8.215 $Y2=2.29
r166 32 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=0.95
+ $X2=8.83 $Y2=0.95
r167 32 45 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.745 $Y=0.95
+ $X2=7.96 $Y2=0.95
r168 30 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.045 $Y=2.385
+ $X2=8.13 $Y2=2.385
r169 30 43 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.045 $Y=2.385
+ $X2=7.63 $Y2=2.385
r170 28 44 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.36 $Y=0.805
+ $X2=7.79 $Y2=0.805
r171 25 42 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.965 $Y=2.385
+ $X2=7.3 $Y2=2.385
r172 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.8
+ $Y=1.99 $X2=6.8 $Y2=1.99
r173 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.8 $Y=2.3
+ $X2=6.965 $Y2=2.385
r174 19 21 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.8 $Y=2.3 $X2=6.8
+ $Y2=1.99
r175 15 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.53 $Y=1.2
+ $X2=6.74 $Y2=1.2
r176 14 22 38.7725 $w=3.49e-07 $l=1.81659e-07 $layer=POLY_cond $X=6.74 $Y=1.825
+ $X2=6.775 $Y2=1.99
r177 13 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.74 $Y=1.275
+ $X2=6.74 $Y2=1.2
r178 13 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.74 $Y=1.275
+ $X2=6.74 $Y2=1.825
r179 10 22 45.6779 $w=3.49e-07 $l=2.66364e-07 $layer=POLY_cond $X=6.66 $Y=2.205
+ $X2=6.775 $Y2=1.99
r180 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.66 $Y=2.205
+ $X2=6.66 $Y2=2.525
r181 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.53 $Y=1.125
+ $X2=6.53 $Y2=1.2
r182 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.53 $Y=1.125
+ $X2=6.53 $Y2=0.805
r183 2 41 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.325
+ $Y=2.315 $X2=7.465 $Y2=2.525
r184 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=7.235
+ $Y=0.595 $X2=7.36 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%A_1163_119# 1 2 9 11 13 16 18 20 23 29 33
+ 37 38 40 41 42 45 46 47
c129 47 0 1.69947e-19 $X=7.505 $Y=1.257
c130 41 0 2.70218e-20 $X=6.037 $Y=2.02
c131 40 0 4.4433e-20 $X=5.972 $Y=1.242
c132 33 0 1.49559e-20 $X=8.385 $Y=1.29
r133 45 48 15.7745 $w=2.75e-07 $l=9e-08 $layer=POLY_cond $X=7.34 $Y=1.29
+ $X2=7.25 $Y2=1.29
r134 44 47 8.99284 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=1.257
+ $X2=7.505 $Y2=1.257
r135 44 46 8.30985 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=1.257
+ $X2=7.175 $Y2=1.257
r136 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.34
+ $Y=1.29 $X2=7.34 $Y2=1.29
r137 41 42 8.67671 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=6.037 $Y=2.02
+ $X2=6.037 $Y2=2.19
r138 38 53 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=8.48 $Y=1.51
+ $X2=8.6 $Y2=1.51
r139 38 51 10.7111 $w=3.15e-07 $l=7e-08 $layer=POLY_cond $X=8.48 $Y=1.51
+ $X2=8.41 $Y2=1.51
r140 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.48
+ $Y=1.51 $X2=8.48 $Y2=1.51
r141 35 37 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=8.48 $Y=1.375
+ $X2=8.48 $Y2=1.51
r142 33 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.385 $Y=1.29
+ $X2=8.48 $Y2=1.375
r143 33 47 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=8.385 $Y=1.29
+ $X2=7.505 $Y2=1.29
r144 32 40 1.79954 $w=2.05e-07 $l=1.48e-07 $layer=LI1_cond $X=6.12 $Y=1.242
+ $X2=5.972 $Y2=1.242
r145 32 46 57.0776 $w=2.03e-07 $l=1.055e-06 $layer=LI1_cond $X=6.12 $Y=1.242
+ $X2=7.175 $Y2=1.242
r146 29 42 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.1 $Y=2.525
+ $X2=6.1 $Y2=2.19
r147 25 40 4.64645 $w=2.32e-07 $l=1.30365e-07 $layer=LI1_cond $X=5.91 $Y=1.345
+ $X2=5.972 $Y2=1.242
r148 25 41 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=5.91 $Y=1.345
+ $X2=5.91 $Y2=2.02
r149 21 40 4.64645 $w=2.32e-07 $l=1.02e-07 $layer=LI1_cond $X=5.972 $Y=1.14
+ $X2=5.972 $Y2=1.242
r150 21 23 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=5.972 $Y=1.14
+ $X2=5.972 $Y2=0.805
r151 18 53 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.6 $Y=1.345
+ $X2=8.6 $Y2=1.51
r152 18 20 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.6 $Y=1.345
+ $X2=8.6 $Y2=0.915
r153 14 51 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.41 $Y=1.675
+ $X2=8.41 $Y2=1.51
r154 14 16 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=8.41 $Y=1.675
+ $X2=8.41 $Y2=2.315
r155 11 45 41.1891 $w=2.75e-07 $l=3.06594e-07 $layer=POLY_cond $X=7.575 $Y=1.125
+ $X2=7.34 $Y2=1.29
r156 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.575 $Y=1.125
+ $X2=7.575 $Y2=0.805
r157 7 48 16.9318 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.25 $Y=1.455
+ $X2=7.25 $Y2=1.29
r158 7 9 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=7.25 $Y=1.455
+ $X2=7.25 $Y2=2.525
r159 2 29 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.945
+ $Y=2.315 $X2=6.085 $Y2=2.525
r160 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.815
+ $Y=0.595 $X2=5.955 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%SET_B 3 7 9 11 14 16 17 18 19 23 24 25 26
+ 31 34 35 40 41
c129 35 0 2.54e-20 $X=10.8 $Y=1.795
c130 34 0 1.1803e-19 $X=10.8 $Y=1.795
c131 26 0 2.91077e-19 $X=7.585 $Y=2.035
c132 19 0 1.40653e-19 $X=10.47 $Y=2.225
r133 39 41 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=7.7 $Y=1.99
+ $X2=7.935 $Y2=1.99
r134 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.7
+ $Y=1.99 $X2=7.7 $Y2=1.99
r135 36 39 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=7.68 $Y=1.99 $X2=7.7
+ $Y2=1.99
r136 35 50 14.0096 $w=1.88e-07 $l=2.4e-07 $layer=LI1_cond $X=10.8 $Y=1.795
+ $X2=10.8 $Y2=2.035
r137 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.8
+ $Y=1.795 $X2=10.8 $Y2=1.795
r138 31 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r139 29 40 12.7504 $w=2.33e-07 $l=2.6e-07 $layer=LI1_cond $X=7.44 $Y=2.012
+ $X2=7.7 $Y2=2.012
r140 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=2.035
+ $X2=7.44 $Y2=2.035
r141 26 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=2.035
+ $X2=7.44 $Y2=2.035
r142 25 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r143 25 26 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=7.585 $Y2=2.035
r144 24 34 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=10.8 $Y=2.15
+ $X2=10.8 $Y2=1.795
r145 23 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.8 $Y=1.63
+ $X2=10.8 $Y2=1.795
r146 20 23 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=10.71 $Y=1.275
+ $X2=10.71 $Y2=1.63
r147 18 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=10.635 $Y=2.225
+ $X2=10.8 $Y2=2.15
r148 18 19 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.635 $Y=2.225
+ $X2=10.47 $Y2=2.225
r149 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.635 $Y=1.2
+ $X2=10.71 $Y2=1.275
r150 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=10.635 $Y=1.2
+ $X2=10.365 $Y2=1.2
r151 12 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.395 $Y=2.3
+ $X2=10.47 $Y2=2.225
r152 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.395 $Y=2.3
+ $X2=10.395 $Y2=2.67
r153 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.29 $Y=1.125
+ $X2=10.365 $Y2=1.2
r154 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.29 $Y=1.125
+ $X2=10.29 $Y2=0.805
r155 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.935 $Y=1.825
+ $X2=7.935 $Y2=1.99
r156 5 7 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=7.935 $Y=1.825
+ $X2=7.935 $Y2=0.805
r157 1 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.68 $Y=2.155
+ $X2=7.68 $Y2=1.99
r158 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.68 $Y=2.155
+ $X2=7.68 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%A_629_47# 1 2 10 14 15 16 17 18 21 23 27 29
+ 33 37 39 40 41 47 50 52 55
c131 55 0 1.99828e-19 $X=4.24 $Y=1.06
c132 52 0 4.28533e-20 $X=3.745 $Y=1.23
c133 21 0 4.4433e-20 $X=5.74 $Y=0.805
r134 55 58 81.9121 $w=5.25e-07 $l=5.05e-07 $layer=POLY_cond $X=4.337 $Y=1.06
+ $X2=4.337 $Y2=1.565
r135 55 57 47.2626 $w=5.25e-07 $l=1.65e-07 $layer=POLY_cond $X=4.337 $Y=1.06
+ $X2=4.337 $Y2=0.895
r136 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.24
+ $Y=1.06 $X2=4.24 $Y2=1.06
r137 52 54 9.6624 $w=6.25e-07 $l=4.95e-07 $layer=LI1_cond $X=3.745 $Y=1.23
+ $X2=4.24 $Y2=1.23
r138 51 52 4.88 $w=6.25e-07 $l=2.5e-07 $layer=LI1_cond $X=3.495 $Y=1.23
+ $X2=3.745 $Y2=1.23
r139 50 52 3.4964 $w=3.9e-07 $l=3.35e-07 $layer=LI1_cond $X=3.745 $Y=0.895
+ $X2=3.745 $Y2=1.23
r140 49 50 8.56945 $w=3.88e-07 $l=2.9e-07 $layer=LI1_cond $X=3.745 $Y=0.605
+ $X2=3.745 $Y2=0.895
r141 45 51 7.86514 $w=1.9e-07 $l=3.35e-07 $layer=LI1_cond $X=3.495 $Y=1.565
+ $X2=3.495 $Y2=1.23
r142 45 47 52.244 $w=1.88e-07 $l=8.95e-07 $layer=LI1_cond $X=3.495 $Y=1.565
+ $X2=3.495 $Y2=2.46
r143 41 49 6.87824 $w=3.3e-07 $l=2.64953e-07 $layer=LI1_cond $X=3.55 $Y=0.44
+ $X2=3.745 $Y2=0.605
r144 41 43 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.55 $Y=0.44
+ $X2=3.285 $Y2=0.44
r145 35 37 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=9.57 $Y=0.255
+ $X2=9.57 $Y2=0.805
r146 31 33 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=8.92 $Y=3.075
+ $X2=8.92 $Y2=2.46
r147 30 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.375 $Y=3.15
+ $X2=6.3 $Y2=3.15
r148 29 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.845 $Y=3.15
+ $X2=8.92 $Y2=3.075
r149 29 30 1266.53 $w=1.5e-07 $l=2.47e-06 $layer=POLY_cond $X=8.845 $Y=3.15
+ $X2=6.375 $Y2=3.15
r150 25 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.3 $Y=3.075
+ $X2=6.3 $Y2=3.15
r151 25 27 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.3 $Y=3.075
+ $X2=6.3 $Y2=2.525
r152 24 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.815 $Y=0.18
+ $X2=5.74 $Y2=0.18
r153 23 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.495 $Y=0.18
+ $X2=9.57 $Y2=0.255
r154 23 24 1886.98 $w=1.5e-07 $l=3.68e-06 $layer=POLY_cond $X=9.495 $Y=0.18
+ $X2=5.815 $Y2=0.18
r155 19 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.74 $Y=0.255
+ $X2=5.74 $Y2=0.18
r156 19 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.74 $Y=0.255
+ $X2=5.74 $Y2=0.805
r157 17 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.225 $Y=3.15
+ $X2=6.3 $Y2=3.15
r158 17 18 833.245 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=6.225 $Y=3.15
+ $X2=4.6 $Y2=3.15
r159 15 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.665 $Y=0.18
+ $X2=5.74 $Y2=0.18
r160 15 16 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=5.665 $Y=0.18
+ $X2=4.6 $Y2=0.18
r161 14 58 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.525 $Y=2.265
+ $X2=4.525 $Y2=1.565
r162 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.525 $Y=3.075
+ $X2=4.6 $Y2=3.15
r163 12 14 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.525 $Y=3.075
+ $X2=4.525 $Y2=2.265
r164 10 57 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.525 $Y=0.575
+ $X2=4.525 $Y2=0.895
r165 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.525 $Y=0.255
+ $X2=4.6 $Y2=0.18
r166 7 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.525 $Y=0.255
+ $X2=4.525 $Y2=0.575
r167 2 47 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.355
+ $Y=2.335 $X2=3.495 $Y2=2.46
r168 1 43 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.235 $X2=3.285 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%A_1946_369# 1 2 9 13 17 20 21 24 26 28 33
+ 34 36
c92 17 0 1.11454e-19 $X=10.18 $Y=1.68
c93 9 0 1.78649e-19 $X=9.805 $Y=2.67
r94 32 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=11.84 $Y=1.255
+ $X2=11.84 $Y2=1.815
r95 28 33 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.755 $Y=1.98
+ $X2=11.84 $Y2=1.815
r96 28 30 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=11.755 $Y=1.98
+ $X2=11.5 $Y2=1.98
r97 27 34 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.38 $Y=1.17
+ $X2=11.25 $Y2=1.17
r98 26 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.755 $Y=1.17
+ $X2=11.84 $Y2=1.255
r99 26 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.755 $Y=1.17
+ $X2=11.38 $Y2=1.17
r100 22 34 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=11.25 $Y=1.085
+ $X2=11.25 $Y2=1.17
r101 22 24 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=11.25 $Y=1.085
+ $X2=11.25 $Y2=0.875
r102 20 34 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.12 $Y=1.17
+ $X2=11.25 $Y2=1.17
r103 20 21 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=11.12 $Y=1.17
+ $X2=10.345 $Y2=1.17
r104 18 36 36.5152 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=10.18 $Y=1.755
+ $X2=9.93 $Y2=1.755
r105 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.18
+ $Y=1.68 $X2=10.18 $Y2=1.68
r106 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.18 $Y=1.255
+ $X2=10.345 $Y2=1.17
r107 15 17 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=10.18 $Y=1.255
+ $X2=10.18 $Y2=1.68
r108 11 36 21.2229 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.93 $Y=1.515
+ $X2=9.93 $Y2=1.755
r109 11 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=9.93 $Y=1.515
+ $X2=9.93 $Y2=0.805
r110 7 36 18.2576 $w=3.3e-07 $l=2.95973e-07 $layer=POLY_cond $X=9.805 $Y=1.995
+ $X2=9.93 $Y2=1.755
r111 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=9.805 $Y=1.995
+ $X2=9.805 $Y2=2.67
r112 2 30 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=11.375
+ $Y=1.835 $X2=11.5 $Y2=1.98
r113 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=11.16
+ $Y=0.665 $X2=11.285 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%A_1799_408# 1 2 3 12 16 18 22 26 30 34 36
+ 37 40 44 51 53 57 62 64 65 68 69 70 74 75 77 80 85
c175 85 0 2.54e-20 $X=11.79 $Y=1.51
c176 75 0 1.1803e-19 $X=11.235 $Y=1.535
c177 74 0 1.29912e-19 $X=11.15 $Y=2.505
c178 62 0 2.91996e-20 $X=9.75 $Y=2.155
c179 57 0 1.63067e-19 $X=9.665 $Y=0.725
r180 84 85 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.715 $Y=1.51
+ $X2=11.79 $Y2=1.51
r181 83 84 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=11.5 $Y=1.51
+ $X2=11.715 $Y2=1.51
r182 78 83 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.41 $Y=1.51
+ $X2=11.5 $Y2=1.51
r183 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.41
+ $Y=1.51 $X2=11.41 $Y2=1.51
r184 75 77 9.16716 $w=2.18e-07 $l=1.75e-07 $layer=LI1_cond $X=11.235 $Y=1.535
+ $X2=11.41 $Y2=1.535
r185 73 75 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=11.15 $Y=1.645
+ $X2=11.235 $Y2=1.535
r186 73 74 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=11.15 $Y=1.645
+ $X2=11.15 $Y2=2.505
r187 70 72 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=10.535 $Y=2.67
+ $X2=10.61 $Y2=2.67
r188 69 74 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.065 $Y=2.67
+ $X2=11.15 $Y2=2.505
r189 69 72 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=11.065 $Y=2.67
+ $X2=10.61 $Y2=2.67
r190 68 70 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.45 $Y=2.505
+ $X2=10.535 $Y2=2.67
r191 67 68 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.45 $Y=2.335
+ $X2=10.45 $Y2=2.505
r192 66 80 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.835 $Y=2.245
+ $X2=9.75 $Y2=2.245
r193 65 67 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=10.365 $Y=2.245
+ $X2=10.45 $Y2=2.335
r194 65 66 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=10.365 $Y=2.245
+ $X2=9.835 $Y2=2.245
r195 63 80 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.75 $Y=2.335 $X2=9.75
+ $Y2=2.245
r196 63 64 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.75 $Y=2.335
+ $X2=9.75 $Y2=2.555
r197 62 80 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.75 $Y=2.155 $X2=9.75
+ $Y2=2.245
r198 61 62 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=9.75 $Y=0.86
+ $X2=9.75 $Y2=2.155
r199 57 61 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=9.665 $Y=0.725
+ $X2=9.75 $Y2=0.86
r200 57 59 15.5793 $w=2.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.665 $Y=0.725
+ $X2=9.3 $Y2=0.725
r201 53 64 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.665 $Y=2.72
+ $X2=9.75 $Y2=2.555
r202 53 55 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=9.665 $Y=2.72
+ $X2=9.135 $Y2=2.72
r203 50 51 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=13.045 $Y=1.42
+ $X2=13.195 $Y2=1.42
r204 48 49 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=12.52 $Y=1.42
+ $X2=12.67 $Y2=1.42
r205 47 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.24 $Y=1.42
+ $X2=12.52 $Y2=1.42
r206 46 47 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=12.09 $Y=1.42
+ $X2=12.24 $Y2=1.42
r207 42 51 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.195 $Y=1.495
+ $X2=13.195 $Y2=1.42
r208 42 44 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.195 $Y=1.495
+ $X2=13.195 $Y2=2.155
r209 38 50 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.045 $Y=1.345
+ $X2=13.045 $Y2=1.42
r210 38 40 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=13.045 $Y=1.345
+ $X2=13.045 $Y2=0.455
r211 37 49 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.745 $Y=1.42
+ $X2=12.67 $Y2=1.42
r212 36 50 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.97 $Y=1.42
+ $X2=13.045 $Y2=1.42
r213 36 37 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=12.97 $Y=1.42
+ $X2=12.745 $Y2=1.42
r214 32 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.67 $Y=1.495
+ $X2=12.67 $Y2=1.42
r215 32 34 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=12.67 $Y=1.495
+ $X2=12.67 $Y2=2.465
r216 28 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.52 $Y=1.345
+ $X2=12.52 $Y2=1.42
r217 28 30 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=12.52 $Y=1.345
+ $X2=12.52 $Y2=0.665
r218 24 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.24 $Y=1.495
+ $X2=12.24 $Y2=1.42
r219 24 26 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=12.24 $Y=1.495
+ $X2=12.24 $Y2=2.465
r220 20 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.09 $Y=1.345
+ $X2=12.09 $Y2=1.42
r221 20 22 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=12.09 $Y=1.345
+ $X2=12.09 $Y2=0.665
r222 18 46 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.015 $Y=1.42
+ $X2=12.09 $Y2=1.42
r223 18 85 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=12.015 $Y=1.42
+ $X2=11.79 $Y2=1.42
r224 14 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.715 $Y=1.675
+ $X2=11.715 $Y2=1.51
r225 14 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=11.715 $Y=1.675
+ $X2=11.715 $Y2=2.045
r226 10 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.5 $Y=1.345
+ $X2=11.5 $Y2=1.51
r227 10 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=11.5 $Y=1.345 $X2=11.5
+ $Y2=0.875
r228 3 72 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=10.47
+ $Y=2.46 $X2=10.61 $Y2=2.67
r229 2 55 600 $w=1.7e-07 $l=7.46726e-07 $layer=licon1_PDIFF $count=1 $X=8.995
+ $Y=2.04 $X2=9.135 $Y2=2.72
r230 1 59 182 $w=1.7e-07 $l=2.47386e-07 $layer=licon1_NDIFF $count=1 $X=9.12
+ $Y=0.595 $X2=9.3 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%A_2624_49# 1 2 9 13 17 21 24 27 31 37 39 44
r58 43 44 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=14.405 $Y=1.44
+ $X2=14.835 $Y2=1.44
r59 35 37 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=13.26 $Y=0.455
+ $X2=13.37 $Y2=0.455
r60 32 43 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=14.27 $Y=1.44
+ $X2=14.405 $Y2=1.44
r61 32 40 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=14.27 $Y=1.44
+ $X2=14.035 $Y2=1.44
r62 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=14.27
+ $Y=1.44 $X2=14.27 $Y2=1.44
r63 29 39 0.499868 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=13.575 $Y=1.44
+ $X2=13.42 $Y2=1.44
r64 29 31 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=13.575 $Y=1.44
+ $X2=14.27 $Y2=1.44
r65 25 39 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=13.42 $Y=1.605
+ $X2=13.42 $Y2=1.44
r66 25 27 13.9408 $w=3.08e-07 $l=3.75e-07 $layer=LI1_cond $X=13.42 $Y=1.605
+ $X2=13.42 $Y2=1.98
r67 24 39 6.26932 $w=2.6e-07 $l=1.88348e-07 $layer=LI1_cond $X=13.37 $Y=1.275
+ $X2=13.42 $Y2=1.44
r68 23 37 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=13.37 $Y=0.62
+ $X2=13.37 $Y2=0.455
r69 23 24 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=13.37 $Y=0.62
+ $X2=13.37 $Y2=1.275
r70 19 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.835 $Y=1.605
+ $X2=14.835 $Y2=1.44
r71 19 21 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=14.835 $Y=1.605
+ $X2=14.835 $Y2=2.465
r72 15 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.835 $Y=1.275
+ $X2=14.835 $Y2=1.44
r73 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=14.835 $Y=1.275
+ $X2=14.835 $Y2=0.655
r74 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.405 $Y=1.605
+ $X2=14.405 $Y2=1.44
r75 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=14.405 $Y=1.605
+ $X2=14.405 $Y2=2.465
r76 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.035 $Y=1.275
+ $X2=14.035 $Y2=1.44
r77 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=14.035 $Y=1.275
+ $X2=14.035 $Y2=0.655
r78 2 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=13.27
+ $Y=1.835 $X2=13.41 $Y2=1.98
r79 1 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.12
+ $Y=0.245 $X2=13.26 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 57 63 67 69 74 75 77 78 80 81 83 84 86 87 88 90 95 110 136 140 146 149 156 159
+ 163
r168 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r169 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r170 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r171 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r172 149 152 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.61 $Y=3.07
+ $X2=2.61 $Y2=3.33
r173 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r174 144 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r175 144 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r176 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r177 141 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.355 $Y=3.33
+ $X2=14.19 $Y2=3.33
r178 141 143 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=14.355 $Y=3.33
+ $X2=14.64 $Y2=3.33
r179 140 162 4.14267 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=14.945 $Y=3.33
+ $X2=15.152 $Y2=3.33
r180 140 143 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=14.945 $Y=3.33
+ $X2=14.64 $Y2=3.33
r181 139 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r182 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r183 136 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.025 $Y=3.33
+ $X2=14.19 $Y2=3.33
r184 136 138 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=14.025 $Y=3.33
+ $X2=13.68 $Y2=3.33
r185 135 139 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r186 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r187 132 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r188 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r189 129 132 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.76 $Y2=3.33
r190 128 131 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=10.32 $Y=3.33
+ $X2=11.76 $Y2=3.33
r191 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r192 126 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r193 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r194 123 126 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.84 $Y2=3.33
r195 122 125 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.84 $Y2=3.33
r196 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r197 120 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r198 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r199 117 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.12 $Y=3.33
+ $X2=6.955 $Y2=3.33
r200 117 119 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.12 $Y=3.33
+ $X2=7.92 $Y2=3.33
r201 116 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r202 115 116 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r203 113 116 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r204 112 115 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r205 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r206 110 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.79 $Y=3.33
+ $X2=6.955 $Y2=3.33
r207 110 115 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.79 $Y=3.33
+ $X2=6.48 $Y2=3.33
r208 109 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r209 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r210 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r211 106 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r212 105 108 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r213 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r214 103 152 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.61 $Y2=3.33
r215 103 105 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=3.12 $Y2=3.33
r216 102 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r217 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r218 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r219 99 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r220 98 101 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r221 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r222 96 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r223 96 98 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r224 95 152 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.61 $Y2=3.33
r225 95 101 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.16 $Y2=3.33
r226 93 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r227 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r228 90 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r229 90 92 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r230 88 120 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=7.92 $Y2=3.33
r231 88 157 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=6.96 $Y2=3.33
r232 86 134 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=12.755 $Y=3.33
+ $X2=12.72 $Y2=3.33
r233 86 87 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.755 $Y=3.33
+ $X2=12.925 $Y2=3.33
r234 85 138 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=13.095 $Y=3.33
+ $X2=13.68 $Y2=3.33
r235 85 87 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=13.095 $Y=3.33
+ $X2=12.925 $Y2=3.33
r236 83 131 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=11.86 $Y=3.33
+ $X2=11.76 $Y2=3.33
r237 83 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.86 $Y=3.33
+ $X2=11.99 $Y2=3.33
r238 82 134 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=12.12 $Y=3.33
+ $X2=12.72 $Y2=3.33
r239 82 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.12 $Y=3.33
+ $X2=11.99 $Y2=3.33
r240 80 125 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.005 $Y=3.33
+ $X2=9.84 $Y2=3.33
r241 80 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=10.005 $Y=3.33
+ $X2=10.1 $Y2=3.33
r242 79 128 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=10.32 $Y2=3.33
r243 79 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=10.1 $Y2=3.33
r244 77 119 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=7.95 $Y=3.33
+ $X2=7.92 $Y2=3.33
r245 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.95 $Y=3.33
+ $X2=8.115 $Y2=3.33
r246 76 122 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.28 $Y=3.33
+ $X2=8.4 $Y2=3.33
r247 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=3.33
+ $X2=8.115 $Y2=3.33
r248 74 108 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.1 $Y=3.33 $X2=4.08
+ $Y2=3.33
r249 74 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.1 $Y=3.33 $X2=4.23
+ $Y2=3.33
r250 73 112 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.36 $Y=3.33
+ $X2=4.56 $Y2=3.33
r251 73 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.36 $Y=3.33
+ $X2=4.23 $Y2=3.33
r252 69 72 41.1892 $w=2.68e-07 $l=9.65e-07 $layer=LI1_cond $X=15.08 $Y=1.985
+ $X2=15.08 $Y2=2.95
r253 67 162 3.14202 $w=2.7e-07 $l=1.15521e-07 $layer=LI1_cond $X=15.08 $Y=3.245
+ $X2=15.152 $Y2=3.33
r254 67 72 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.08 $Y=3.245
+ $X2=15.08 $Y2=2.95
r255 63 66 33.7002 $w=3.28e-07 $l=9.65e-07 $layer=LI1_cond $X=14.19 $Y=1.985
+ $X2=14.19 $Y2=2.95
r256 61 159 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.19 $Y=3.245
+ $X2=14.19 $Y2=3.33
r257 61 66 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=14.19 $Y=3.245
+ $X2=14.19 $Y2=2.95
r258 57 60 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=12.925 $Y=1.98
+ $X2=12.925 $Y2=2.445
r259 55 87 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=12.925 $Y=3.245
+ $X2=12.925 $Y2=3.33
r260 55 60 27.1163 $w=3.38e-07 $l=8e-07 $layer=LI1_cond $X=12.925 $Y=3.245
+ $X2=12.925 $Y2=2.445
r261 51 84 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=11.99 $Y=3.245
+ $X2=11.99 $Y2=3.33
r262 51 53 33.9084 $w=2.58e-07 $l=7.65e-07 $layer=LI1_cond $X=11.99 $Y=3.245
+ $X2=11.99 $Y2=2.48
r263 47 81 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=10.1 $Y=3.245
+ $X2=10.1 $Y2=3.33
r264 47 49 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=10.1 $Y=3.245
+ $X2=10.1 $Y2=2.67
r265 43 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=3.245
+ $X2=8.115 $Y2=3.33
r266 43 45 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=8.115 $Y=3.245
+ $X2=8.115 $Y2=2.735
r267 39 156 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=3.245
+ $X2=6.955 $Y2=3.33
r268 39 41 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=6.955 $Y=3.245
+ $X2=6.955 $Y2=2.735
r269 35 75 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.23 $Y=3.245
+ $X2=4.23 $Y2=3.33
r270 35 37 17.9515 $w=2.58e-07 $l=4.05e-07 $layer=LI1_cond $X=4.23 $Y=3.245
+ $X2=4.23 $Y2=2.84
r271 31 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r272 31 33 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.85
r273 10 72 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=14.91
+ $Y=1.835 $X2=15.05 $Y2=2.95
r274 10 69 400 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=14.91
+ $Y=1.835 $X2=15.05 $Y2=1.985
r275 9 66 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=14.065
+ $Y=1.835 $X2=14.19 $Y2=2.95
r276 9 63 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=14.065
+ $Y=1.835 $X2=14.19 $Y2=1.985
r277 8 60 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=12.745
+ $Y=1.835 $X2=12.885 $Y2=2.445
r278 8 57 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=12.745
+ $Y=1.835 $X2=12.93 $Y2=1.98
r279 7 53 300 $w=1.7e-07 $l=7.53392e-07 $layer=licon1_PDIFF $count=2 $X=11.79
+ $Y=1.835 $X2=12.025 $Y2=2.48
r280 6 49 600 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_PDIFF $count=1 $X=9.88
+ $Y=2.46 $X2=10.1 $Y2=2.67
r281 5 45 600 $w=1.7e-07 $l=5.72364e-07 $layer=licon1_PDIFF $count=1 $X=7.755
+ $Y=2.315 $X2=8.115 $Y2=2.735
r282 4 41 600 $w=1.7e-07 $l=5.18459e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=2.315 $X2=6.955 $Y2=2.735
r283 3 37 600 $w=1.7e-07 $l=9.6478e-07 $layer=licon1_PDIFF $count=1 $X=4.05
+ $Y=1.945 $X2=4.195 $Y2=2.84
r284 2 149 600 $w=1.7e-07 $l=8.3781e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.335 $X2=2.61 $Y2=3.07
r285 1 33 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.335 $X2=0.69 $Y2=2.85
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%A_268_467# 1 2 3 4 13 19 21 22 24 25 26 28
+ 29 32 33 34 37 40 44 45
c127 24 0 1.83654e-19 $X=2.605 $Y=1.195
c128 21 0 1.0849e-19 $X=2.52 $Y=0.79
r129 45 47 4.3277 $w=2.96e-07 $l=1.05e-07 $layer=LI1_cond $X=5.627 $Y=2.42
+ $X2=5.627 $Y2=2.525
r130 40 45 5.36356 $w=2.96e-07 $l=1.11781e-07 $layer=LI1_cond $X=5.565 $Y=2.335
+ $X2=5.627 $Y2=2.42
r131 40 44 67.7778 $w=1.78e-07 $l=1.1e-06 $layer=LI1_cond $X=5.565 $Y=2.335
+ $X2=5.565 $Y2=1.235
r132 35 44 7.48172 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=5.507 $Y=1.088
+ $X2=5.507 $Y2=1.235
r133 35 37 11.0556 $w=2.93e-07 $l=2.83e-07 $layer=LI1_cond $X=5.507 $Y=1.088
+ $X2=5.507 $Y2=0.805
r134 33 45 3.98214 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.475 $Y=2.42
+ $X2=5.627 $Y2=2.42
r135 33 34 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=5.475 $Y=2.42
+ $X2=3.93 $Y2=2.42
r136 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.845 $Y=2.505
+ $X2=3.93 $Y2=2.42
r137 31 32 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.845 $Y=2.505
+ $X2=3.845 $Y2=2.805
r138 30 42 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=2.9
+ $X2=3.145 $Y2=2.9
r139 29 32 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.76 $Y=2.9
+ $X2=3.845 $Y2=2.805
r140 29 30 30.9378 $w=1.88e-07 $l=5.3e-07 $layer=LI1_cond $X=3.76 $Y=2.9
+ $X2=3.23 $Y2=2.9
r141 27 28 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=3.145 $Y=1.365
+ $X2=3.145 $Y2=2.585
r142 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.06 $Y=1.28
+ $X2=3.145 $Y2=1.365
r143 25 26 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.06 $Y=1.28
+ $X2=2.69 $Y2=1.28
r144 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.605 $Y=1.195
+ $X2=2.69 $Y2=1.28
r145 23 24 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.605 $Y=0.875
+ $X2=2.605 $Y2=1.195
r146 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.52 $Y=0.79
+ $X2=2.605 $Y2=0.875
r147 21 22 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.52 $Y=0.79 $X2=2.22
+ $Y2=0.79
r148 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.095 $Y=0.705
+ $X2=2.22 $Y2=0.79
r149 17 19 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=2.095 $Y=0.705
+ $X2=2.095 $Y2=0.445
r150 13 42 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.145 $Y=2.695
+ $X2=3.145 $Y2=2.9
r151 13 28 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.145 $Y=2.695
+ $X2=3.145 $Y2=2.585
r152 13 15 77.0041 $w=2.18e-07 $l=1.47e-06 $layer=LI1_cond $X=3.06 $Y=2.695
+ $X2=1.59 $Y2=2.695
r153 4 47 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=5.53
+ $Y=2.315 $X2=5.655 $Y2=2.525
r154 3 15 600 $w=1.7e-07 $l=4.73788e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.335 $X2=1.59 $Y2=2.7
r155 2 37 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.595 $X2=5.525 $Y2=0.805
r156 1 19 182 $w=1.7e-07 $l=4.47856e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.235 $X2=2.055 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%Q_N 1 2 7 8 9 10 11 20 32 36
r29 36 37 5.41174 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.37 $Y=1.98
+ $X2=12.37 $Y2=1.815
r30 11 36 1.47406 $w=4.28e-07 $l=5.5e-08 $layer=LI1_cond $X=12.37 $Y=2.035
+ $X2=12.37 $Y2=1.98
r31 11 32 27.7449 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=12.437 $Y=2.12
+ $X2=12.437 $Y2=2.91
r32 10 37 5.66775 $w=3.03e-07 $l=1.5e-07 $layer=LI1_cond $X=12.307 $Y=1.665
+ $X2=12.307 $Y2=1.815
r33 9 10 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=12.307 $Y=1.295
+ $X2=12.307 $Y2=1.665
r34 8 9 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=12.307 $Y=0.925
+ $X2=12.307 $Y2=1.295
r35 7 8 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=12.307 $Y=0.555
+ $X2=12.307 $Y2=0.925
r36 7 20 4.72313 $w=3.03e-07 $l=1.25e-07 $layer=LI1_cond $X=12.307 $Y=0.555
+ $X2=12.307 $Y2=0.43
r37 2 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.315
+ $Y=1.835 $X2=12.455 $Y2=1.98
r38 2 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=12.315
+ $Y=1.835 $X2=12.455 $Y2=2.91
r39 1 20 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=12.165
+ $Y=0.245 $X2=12.305 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%Q 1 2 7 8 9 10 11 12 13 37
r23 13 34 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=14.65 $Y=2.775
+ $X2=14.65 $Y2=2.91
r24 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=14.65 $Y=2.405
+ $X2=14.65 $Y2=2.775
r25 11 12 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=14.65 $Y=1.96
+ $X2=14.65 $Y2=2.405
r26 10 11 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=14.65 $Y=1.665
+ $X2=14.65 $Y2=1.96
r27 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=14.65 $Y=1.295
+ $X2=14.65 $Y2=1.665
r28 9 43 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=14.65 $Y=1.295
+ $X2=14.65 $Y2=1.095
r29 8 43 7.92966 $w=6.63e-07 $l=1.7e-07 $layer=LI1_cond $X=14.442 $Y=0.925
+ $X2=14.442 $Y2=1.095
r30 7 8 6.65487 $w=6.63e-07 $l=3.7e-07 $layer=LI1_cond $X=14.442 $Y=0.555
+ $X2=14.442 $Y2=0.925
r31 7 37 2.42813 $w=6.63e-07 $l=1.35e-07 $layer=LI1_cond $X=14.442 $Y=0.555
+ $X2=14.442 $Y2=0.42
r32 2 34 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=14.48
+ $Y=1.835 $X2=14.62 $Y2=2.91
r33 2 11 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=14.48
+ $Y=1.835 $X2=14.62 $Y2=1.96
r34 1 37 45.5 $w=1.7e-07 $l=5.95357e-07 $layer=licon1_NDIFF $count=4 $X=14.11
+ $Y=0.235 $X2=14.62 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_2%VGND 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 57 63 67 71 73 75 78 79 81 82 84 85 87 88 90 91 92 116 127 131 136 142 145 148
+ 151 155
c174 49 0 1.0012e-19 $X=8.305 $Y=0.59
r175 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r176 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r177 149 152 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.68 $Y2=0
r178 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r179 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r180 142 143 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r181 140 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r182 140 152 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=13.68 $Y2=0
r183 139 140 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r184 137 151 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=13.94 $Y=0
+ $X2=13.797 $Y2=0
r185 137 139 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=13.94 $Y=0
+ $X2=14.64 $Y2=0
r186 136 154 4.14267 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=14.945 $Y=0
+ $X2=15.152 $Y2=0
r187 136 139 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=14.945 $Y=0
+ $X2=14.64 $Y2=0
r188 135 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r189 135 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r190 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r191 132 145 10.3577 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=11.985 $Y=0
+ $X2=11.767 $Y2=0
r192 132 134 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.985 $Y=0
+ $X2=12.24 $Y2=0
r193 131 148 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=12.63 $Y=0
+ $X2=12.797 $Y2=0
r194 131 134 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=12.63 $Y=0
+ $X2=12.24 $Y2=0
r195 130 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r196 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r197 127 145 10.3577 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=11.55 $Y=0
+ $X2=11.767 $Y2=0
r198 127 129 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.55 $Y=0
+ $X2=11.28 $Y2=0
r199 126 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r200 126 143 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=8.4 $Y2=0
r201 125 126 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r202 123 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.47 $Y=0
+ $X2=8.305 $Y2=0
r203 123 125 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=8.47 $Y=0
+ $X2=10.32 $Y2=0
r204 122 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r205 121 122 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r206 118 121 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r207 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r208 116 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.14 $Y=0
+ $X2=8.305 $Y2=0
r209 116 121 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.14 $Y=0
+ $X2=7.92 $Y2=0
r210 115 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r211 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r212 112 115 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r213 111 114 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r214 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r215 109 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r216 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r217 106 109 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.08 $Y2=0
r218 105 108 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r219 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r220 103 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.12 $Y2=0
r221 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r222 100 103 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=2.64 $Y2=0
r223 99 102 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r224 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r225 96 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r226 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r227 92 122 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=7.92 $Y2=0
r228 92 119 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=6.96 $Y2=0
r229 90 125 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=10.34 $Y=0 $X2=10.32
+ $Y2=0
r230 90 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.34 $Y=0
+ $X2=10.505 $Y2=0
r231 89 129 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=10.67 $Y=0
+ $X2=11.28 $Y2=0
r232 89 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.67 $Y=0
+ $X2=10.505 $Y2=0
r233 87 114 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.58 $Y=0 $X2=6.48
+ $Y2=0
r234 87 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.58 $Y=0 $X2=6.745
+ $Y2=0
r235 86 118 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.91 $Y=0 $X2=6.96
+ $Y2=0
r236 86 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.91 $Y=0 $X2=6.745
+ $Y2=0
r237 84 108 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.145 $Y=0
+ $X2=4.08 $Y2=0
r238 84 85 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.145 $Y=0 $X2=4.275
+ $Y2=0
r239 83 111 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.56 $Y2=0
r240 83 85 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.275
+ $Y2=0
r241 81 102 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.64
+ $Y2=0
r242 81 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.855
+ $Y2=0
r243 80 105 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=3.12
+ $Y2=0
r244 80 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=2.855
+ $Y2=0
r245 78 95 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.72
+ $Y2=0
r246 78 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.995
+ $Y2=0
r247 77 99 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.2
+ $Y2=0
r248 77 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=0.995
+ $Y2=0
r249 73 154 3.14202 $w=2.7e-07 $l=1.15521e-07 $layer=LI1_cond $X=15.08 $Y=0.085
+ $X2=15.152 $Y2=0
r250 73 75 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.08 $Y=0.085
+ $X2=15.08 $Y2=0.38
r251 69 151 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=13.797 $Y=0.085
+ $X2=13.797 $Y2=0
r252 69 71 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=13.797 $Y=0.085
+ $X2=13.797 $Y2=0.38
r253 68 148 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=12.965 $Y=0
+ $X2=12.797 $Y2=0
r254 67 151 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=13.655 $Y=0
+ $X2=13.797 $Y2=0
r255 67 68 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.655 $Y=0
+ $X2=12.965 $Y2=0
r256 63 65 18.9207 $w=3.33e-07 $l=5.5e-07 $layer=LI1_cond $X=12.797 $Y=0.39
+ $X2=12.797 $Y2=0.94
r257 61 148 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=12.797 $Y=0.085
+ $X2=12.797 $Y2=0
r258 61 63 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=12.797 $Y=0.085
+ $X2=12.797 $Y2=0.39
r259 57 59 11.6569 $w=4.33e-07 $l=4.4e-07 $layer=LI1_cond $X=11.767 $Y=0.39
+ $X2=11.767 $Y2=0.83
r260 55 145 1.70358 $w=4.35e-07 $l=8.5e-08 $layer=LI1_cond $X=11.767 $Y=0.085
+ $X2=11.767 $Y2=0
r261 55 57 8.08035 $w=4.33e-07 $l=3.05e-07 $layer=LI1_cond $X=11.767 $Y=0.085
+ $X2=11.767 $Y2=0.39
r262 51 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.505 $Y=0.085
+ $X2=10.505 $Y2=0
r263 51 53 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=10.505 $Y=0.085
+ $X2=10.505 $Y2=0.79
r264 47 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.305 $Y=0.085
+ $X2=8.305 $Y2=0
r265 47 49 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=8.305 $Y=0.085
+ $X2=8.305 $Y2=0.59
r266 43 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=0.085
+ $X2=6.745 $Y2=0
r267 43 45 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=6.745 $Y=0.085
+ $X2=6.745 $Y2=0.805
r268 39 85 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.275 $Y=0.085
+ $X2=4.275 $Y2=0
r269 39 41 21.0542 $w=2.58e-07 $l=4.75e-07 $layer=LI1_cond $X=4.275 $Y=0.085
+ $X2=4.275 $Y2=0.56
r270 35 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0
r271 35 37 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0.41
r272 31 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.995 $Y=0.085
+ $X2=0.995 $Y2=0
r273 31 33 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.995 $Y=0.085
+ $X2=0.995 $Y2=0.44
r274 10 75 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.91
+ $Y=0.235 $X2=15.05 $Y2=0.38
r275 9 71 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=13.695
+ $Y=0.235 $X2=13.82 $Y2=0.38
r276 8 65 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=12.595
+ $Y=0.245 $X2=12.735 $Y2=0.94
r277 8 63 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=12.595
+ $Y=0.245 $X2=12.83 $Y2=0.39
r278 7 59 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.665 $X2=11.715 $Y2=0.83
r279 7 57 182 $w=1.7e-07 $l=4.15331e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.665 $X2=11.875 $Y2=0.39
r280 6 53 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=10.365
+ $Y=0.595 $X2=10.505 $Y2=0.79
r281 5 49 182 $w=1.7e-07 $l=2.9749e-07 $layer=licon1_NDIFF $count=1 $X=8.01
+ $Y=0.595 $X2=8.305 $Y2=0.59
r282 4 45 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.605
+ $Y=0.595 $X2=6.745 $Y2=0.805
r283 3 41 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=4.185
+ $Y=0.365 $X2=4.31 $Y2=0.56
r284 2 37 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.855 $Y2=0.41
r285 1 33 182 $w=1.7e-07 $l=2.86356e-07 $layer=licon1_NDIFF $count=1 $X=0.8
+ $Y=0.235 $X2=0.995 $Y2=0.44
.ends

