* File: sky130_fd_sc_lp__ebufn_1.pxi.spice
* Created: Fri Aug 28 10:31:32 2020
* 
x_PM_SKY130_FD_SC_LP__EBUFN_1%A_105_263# N_A_105_263#_M1005_d
+ N_A_105_263#_M1004_d N_A_105_263#_M1007_g N_A_105_263#_M1003_g
+ N_A_105_263#_c_66_n N_A_105_263#_c_73_n N_A_105_263#_c_74_n
+ N_A_105_263#_c_75_n N_A_105_263#_c_76_n N_A_105_263#_c_77_n
+ N_A_105_263#_c_78_n N_A_105_263#_c_67_n N_A_105_263#_c_68_n
+ N_A_105_263#_c_69_n N_A_105_263#_c_70_n N_A_105_263#_c_80_n
+ N_A_105_263#_c_71_n PM_SKY130_FD_SC_LP__EBUFN_1%A_105_263#
x_PM_SKY130_FD_SC_LP__EBUFN_1%A_219_21# N_A_219_21#_M1002_s N_A_219_21#_M1001_s
+ N_A_219_21#_c_155_n N_A_219_21#_M1006_g N_A_219_21#_c_156_n
+ N_A_219_21#_c_157_n N_A_219_21#_c_158_n N_A_219_21#_c_159_n
+ N_A_219_21#_c_160_n PM_SKY130_FD_SC_LP__EBUFN_1%A_219_21#
x_PM_SKY130_FD_SC_LP__EBUFN_1%TE_B N_TE_B_M1000_g N_TE_B_c_195_n N_TE_B_c_196_n
+ N_TE_B_M1001_g N_TE_B_M1002_g TE_B N_TE_B_c_198_n N_TE_B_c_199_n
+ PM_SKY130_FD_SC_LP__EBUFN_1%TE_B
x_PM_SKY130_FD_SC_LP__EBUFN_1%A N_A_M1005_g N_A_M1004_g N_A_c_250_n N_A_c_255_n
+ A N_A_c_251_n N_A_c_252_n PM_SKY130_FD_SC_LP__EBUFN_1%A
x_PM_SKY130_FD_SC_LP__EBUFN_1%Z N_Z_M1003_s N_Z_M1007_s Z Z Z Z Z Z Z
+ N_Z_c_285_n N_Z_c_288_n Z PM_SKY130_FD_SC_LP__EBUFN_1%Z
x_PM_SKY130_FD_SC_LP__EBUFN_1%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_c_311_n
+ N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n VPWR N_VPWR_c_315_n
+ N_VPWR_c_316_n N_VPWR_c_310_n N_VPWR_c_318_n PM_SKY130_FD_SC_LP__EBUFN_1%VPWR
x_PM_SKY130_FD_SC_LP__EBUFN_1%VGND N_VGND_M1006_d N_VGND_M1002_d N_VGND_c_350_n
+ N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n N_VGND_c_354_n N_VGND_c_355_n
+ VGND N_VGND_c_356_n N_VGND_c_357_n PM_SKY130_FD_SC_LP__EBUFN_1%VGND
cc_1 VNB N_A_105_263#_M1007_g 5.24044e-19 $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.465
cc_2 VNB N_A_105_263#_c_66_n 0.0322538f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.54
cc_3 VNB N_A_105_263#_c_67_n 0.0262083f $X=-0.19 $Y=-0.245 $X2=3.67 $Y2=2.11
cc_4 VNB N_A_105_263#_c_68_n 0.0380388f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.48
cc_5 VNB N_A_105_263#_c_69_n 0.00794965f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.48
cc_6 VNB N_A_105_263#_c_70_n 0.0380365f $X=-0.19 $Y=-0.245 $X2=3.405 $Y2=0.87
cc_7 VNB N_A_105_263#_c_71_n 0.021392f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.315
cc_8 VNB N_A_219_21#_c_155_n 0.0186791f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.645
cc_9 VNB N_A_219_21#_c_156_n 0.0415516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_219_21#_c_157_n 0.012053f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.315
cc_11 VNB N_A_219_21#_c_158_n 0.0337425f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.785
cc_12 VNB N_A_219_21#_c_159_n 0.0132618f $X=-0.19 $Y=-0.245 $X2=1.69 $Y2=1.54
cc_13 VNB N_A_219_21#_c_160_n 0.0585697f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=2.905
cc_14 VNB N_TE_B_c_195_n 0.0433326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_TE_B_c_196_n 0.00493143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_TE_B_M1002_g 0.0251571f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.785
cc_17 VNB N_TE_B_c_198_n 0.0526695f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=2.99
cc_18 VNB N_TE_B_c_199_n 0.00310687f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=2.99
cc_19 VNB N_A_M1005_g 0.0289731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_c_250_n 0.0161592f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.315
cc_21 VNB N_A_c_251_n 0.0176768f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.625
cc_22 VNB N_A_c_252_n 0.00733039f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.905
cc_23 VNB Z 0.0260004f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.465
cc_24 VNB N_Z_c_285_n 0.0467718f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.48
cc_25 VNB N_VPWR_c_310_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.522 $Y2=2.195
cc_26 VNB N_VGND_c_350_n 0.0150353f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.465
cc_27 VNB N_VGND_c_351_n 0.0347654f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=0.785
cc_28 VNB N_VGND_c_352_n 0.0351624f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.625
cc_29 VNB N_VGND_c_353_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.905
cc_30 VNB N_VGND_c_354_n 0.0313519f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=2.99
cc_31 VNB N_VGND_c_355_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=2.28
cc_32 VNB N_VGND_c_356_n 0.0251917f $X=-0.19 $Y=-0.245 $X2=3.455 $Y2=2.275
cc_33 VNB N_VGND_c_357_n 0.246807f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.48
cc_34 VPB N_A_105_263#_M1007_g 0.0247909f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.465
cc_35 VPB N_A_105_263#_c_73_n 0.0238789f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.905
cc_36 VPB N_A_105_263#_c_74_n 0.022295f $X=-0.19 $Y=1.655 $X2=2.45 $Y2=2.99
cc_37 VPB N_A_105_263#_c_75_n 0.00353584f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=2.99
cc_38 VPB N_A_105_263#_c_76_n 0.00276053f $X=-0.19 $Y=1.655 $X2=2.535 $Y2=2.905
cc_39 VPB N_A_105_263#_c_77_n 0.00751042f $X=-0.19 $Y=1.655 $X2=3.29 $Y2=2.195
cc_40 VPB N_A_105_263#_c_78_n 0.00120748f $X=-0.19 $Y=1.655 $X2=2.62 $Y2=2.195
cc_41 VPB N_A_105_263#_c_67_n 0.0215851f $X=-0.19 $Y=1.655 $X2=3.67 $Y2=2.11
cc_42 VPB N_A_105_263#_c_80_n 0.0440363f $X=-0.19 $Y=1.655 $X2=3.455 $Y2=2.275
cc_43 VPB N_A_219_21#_c_159_n 0.00432912f $X=-0.19 $Y=1.655 $X2=1.69 $Y2=1.54
cc_44 VPB N_TE_B_M1000_g 0.0201857f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_TE_B_c_195_n 0.034951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_TE_B_c_196_n 0.00171595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_TE_B_M1001_g 0.0273718f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.465
cc_48 VPB N_TE_B_c_198_n 0.0446306f $X=-0.19 $Y=1.655 $X2=2.45 $Y2=2.99
cc_49 VPB N_TE_B_c_199_n 0.00307616f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=2.99
cc_50 VPB N_A_M1004_g 0.0297241f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.645
cc_51 VPB N_A_c_250_n 0.00878056f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.315
cc_52 VPB N_A_c_255_n 0.0168106f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=0.785
cc_53 VPB N_A_c_252_n 0.00524626f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.905
cc_54 VPB Z 0.00844535f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.465
cc_55 VPB Z 0.0501835f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.315
cc_56 VPB N_Z_c_288_n 0.0177785f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_311_n 0.0182969f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.465
cc_58 VPB N_VPWR_c_312_n 0.0175115f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.54
cc_59 VPB N_VPWR_c_313_n 0.031612f $X=-0.19 $Y=1.655 $X2=2.45 $Y2=2.99
cc_60 VPB N_VPWR_c_314_n 0.00632158f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=2.99
cc_61 VPB N_VPWR_c_315_n 0.0334466f $X=-0.19 $Y=1.655 $X2=3.29 $Y2=2.195
cc_62 VPB N_VPWR_c_316_n 0.0225667f $X=-0.19 $Y=1.655 $X2=3.67 $Y2=1.1
cc_63 VPB N_VPWR_c_310_n 0.0773255f $X=-0.19 $Y=1.655 $X2=3.522 $Y2=2.195
cc_64 VPB N_VPWR_c_318_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.315
cc_65 N_A_105_263#_c_66_n N_A_219_21#_c_155_n 0.00301952f $X=1.69 $Y=1.54 $X2=0
+ $Y2=0
cc_66 N_A_105_263#_c_68_n N_A_219_21#_c_155_n 0.0276468f $X=0.69 $Y=1.48 $X2=0
+ $Y2=0
cc_67 N_A_105_263#_c_71_n N_A_219_21#_c_157_n 0.0276468f $X=0.69 $Y=1.315 $X2=0
+ $Y2=0
cc_68 N_A_105_263#_c_66_n N_A_219_21#_c_159_n 0.0141516f $X=1.69 $Y=1.54 $X2=0
+ $Y2=0
cc_69 N_A_105_263#_c_73_n N_A_219_21#_c_159_n 0.0845765f $X=1.775 $Y=2.905 $X2=0
+ $Y2=0
cc_70 N_A_105_263#_c_74_n N_A_219_21#_c_159_n 0.0168878f $X=2.45 $Y=2.99 $X2=0
+ $Y2=0
cc_71 N_A_105_263#_c_78_n N_A_219_21#_c_159_n 0.00702791f $X=2.62 $Y=2.195 $X2=0
+ $Y2=0
cc_72 N_A_105_263#_c_73_n N_TE_B_M1000_g 0.00416382f $X=1.775 $Y=2.905 $X2=0
+ $Y2=0
cc_73 N_A_105_263#_c_66_n N_TE_B_c_195_n 0.0244499f $X=1.69 $Y=1.54 $X2=0 $Y2=0
cc_74 N_A_105_263#_c_73_n N_TE_B_c_195_n 0.00974534f $X=1.775 $Y=2.905 $X2=0
+ $Y2=0
cc_75 N_A_105_263#_M1007_g N_TE_B_c_196_n 0.0801807f $X=0.75 $Y=2.465 $X2=0
+ $Y2=0
cc_76 N_A_105_263#_c_66_n N_TE_B_c_196_n 0.00854499f $X=1.69 $Y=1.54 $X2=0 $Y2=0
cc_77 N_A_105_263#_c_68_n N_TE_B_c_196_n 0.00591602f $X=0.69 $Y=1.48 $X2=0 $Y2=0
cc_78 N_A_105_263#_c_73_n N_TE_B_M1001_g 0.0029121f $X=1.775 $Y=2.905 $X2=0
+ $Y2=0
cc_79 N_A_105_263#_c_74_n N_TE_B_M1001_g 0.00703402f $X=2.45 $Y=2.99 $X2=0 $Y2=0
cc_80 N_A_105_263#_c_76_n N_TE_B_M1001_g 0.00670669f $X=2.535 $Y=2.905 $X2=0
+ $Y2=0
cc_81 N_A_105_263#_c_78_n N_TE_B_M1001_g 0.00162743f $X=2.62 $Y=2.195 $X2=0
+ $Y2=0
cc_82 N_A_105_263#_c_66_n N_TE_B_c_198_n 4.72256e-19 $X=1.69 $Y=1.54 $X2=0 $Y2=0
cc_83 N_A_105_263#_c_73_n N_TE_B_c_198_n 0.00325876f $X=1.775 $Y=2.905 $X2=0
+ $Y2=0
cc_84 N_A_105_263#_c_77_n N_TE_B_c_198_n 0.00505125f $X=3.29 $Y=2.195 $X2=0
+ $Y2=0
cc_85 N_A_105_263#_c_78_n N_TE_B_c_198_n 0.00132244f $X=2.62 $Y=2.195 $X2=0
+ $Y2=0
cc_86 N_A_105_263#_c_77_n N_TE_B_c_199_n 0.0126538f $X=3.29 $Y=2.195 $X2=0 $Y2=0
cc_87 N_A_105_263#_c_78_n N_TE_B_c_199_n 0.015051f $X=2.62 $Y=2.195 $X2=0 $Y2=0
cc_88 N_A_105_263#_c_67_n N_A_M1005_g 0.00348663f $X=3.67 $Y=2.11 $X2=0 $Y2=0
cc_89 N_A_105_263#_c_70_n N_A_M1005_g 0.00703678f $X=3.405 $Y=0.87 $X2=0 $Y2=0
cc_90 N_A_105_263#_c_76_n N_A_M1004_g 0.00193708f $X=2.535 $Y=2.905 $X2=0 $Y2=0
cc_91 N_A_105_263#_c_77_n N_A_M1004_g 0.0144436f $X=3.29 $Y=2.195 $X2=0 $Y2=0
cc_92 N_A_105_263#_c_67_n N_A_M1004_g 0.00348663f $X=3.67 $Y=2.11 $X2=0 $Y2=0
cc_93 N_A_105_263#_c_80_n N_A_M1004_g 4.66927e-19 $X=3.455 $Y=2.275 $X2=0 $Y2=0
cc_94 N_A_105_263#_c_77_n N_A_c_255_n 0.00142599f $X=3.29 $Y=2.195 $X2=0 $Y2=0
cc_95 N_A_105_263#_c_80_n N_A_c_255_n 0.00335084f $X=3.455 $Y=2.275 $X2=0 $Y2=0
cc_96 N_A_105_263#_c_67_n N_A_c_251_n 0.00469931f $X=3.67 $Y=2.11 $X2=0 $Y2=0
cc_97 N_A_105_263#_c_70_n N_A_c_251_n 0.00398248f $X=3.405 $Y=0.87 $X2=0 $Y2=0
cc_98 N_A_105_263#_c_77_n N_A_c_252_n 0.022406f $X=3.29 $Y=2.195 $X2=0 $Y2=0
cc_99 N_A_105_263#_c_67_n N_A_c_252_n 0.0512207f $X=3.67 $Y=2.11 $X2=0 $Y2=0
cc_100 N_A_105_263#_c_70_n N_A_c_252_n 0.0149398f $X=3.405 $Y=0.87 $X2=0 $Y2=0
cc_101 N_A_105_263#_c_80_n N_A_c_252_n 0.0110804f $X=3.455 $Y=2.275 $X2=0 $Y2=0
cc_102 N_A_105_263#_M1007_g Z 0.00361456f $X=0.75 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_105_263#_c_68_n Z 0.00236386f $X=0.69 $Y=1.48 $X2=0 $Y2=0
cc_104 N_A_105_263#_c_69_n Z 0.0261014f $X=0.855 $Y=1.48 $X2=0 $Y2=0
cc_105 N_A_105_263#_c_71_n Z 0.00350258f $X=0.69 $Y=1.315 $X2=0 $Y2=0
cc_106 N_A_105_263#_M1007_g Z 0.0197637f $X=0.75 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_105_263#_c_68_n N_Z_c_285_n 0.00413786f $X=0.69 $Y=1.48 $X2=0 $Y2=0
cc_108 N_A_105_263#_c_69_n N_Z_c_285_n 0.01418f $X=0.855 $Y=1.48 $X2=0 $Y2=0
cc_109 N_A_105_263#_c_71_n N_Z_c_285_n 0.0161297f $X=0.69 $Y=1.315 $X2=0 $Y2=0
cc_110 N_A_105_263#_M1007_g N_Z_c_288_n 0.00554338f $X=0.75 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_105_263#_c_68_n N_Z_c_288_n 0.00349435f $X=0.69 $Y=1.48 $X2=0 $Y2=0
cc_112 N_A_105_263#_c_69_n N_Z_c_288_n 0.0145658f $X=0.855 $Y=1.48 $X2=0 $Y2=0
cc_113 N_A_105_263#_c_76_n N_VPWR_M1001_d 0.0100476f $X=2.535 $Y=2.905 $X2=0
+ $Y2=0
cc_114 N_A_105_263#_c_77_n N_VPWR_M1001_d 0.0119143f $X=3.29 $Y=2.195 $X2=0
+ $Y2=0
cc_115 N_A_105_263#_c_78_n N_VPWR_M1001_d 0.0013118f $X=2.62 $Y=2.195 $X2=0
+ $Y2=0
cc_116 N_A_105_263#_M1007_g N_VPWR_c_311_n 0.00485253f $X=0.75 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_105_263#_c_66_n N_VPWR_c_311_n 0.0263218f $X=1.69 $Y=1.54 $X2=0 $Y2=0
cc_118 N_A_105_263#_c_73_n N_VPWR_c_311_n 0.0879683f $X=1.775 $Y=2.905 $X2=0
+ $Y2=0
cc_119 N_A_105_263#_c_75_n N_VPWR_c_311_n 0.0150383f $X=1.86 $Y=2.99 $X2=0 $Y2=0
cc_120 N_A_105_263#_c_74_n N_VPWR_c_312_n 0.0150385f $X=2.45 $Y=2.99 $X2=0 $Y2=0
cc_121 N_A_105_263#_c_76_n N_VPWR_c_312_n 0.0351204f $X=2.535 $Y=2.905 $X2=0
+ $Y2=0
cc_122 N_A_105_263#_c_77_n N_VPWR_c_312_n 0.0219853f $X=3.29 $Y=2.195 $X2=0
+ $Y2=0
cc_123 N_A_105_263#_c_80_n N_VPWR_c_312_n 0.0135901f $X=3.455 $Y=2.275 $X2=0
+ $Y2=0
cc_124 N_A_105_263#_c_74_n N_VPWR_c_313_n 0.0501353f $X=2.45 $Y=2.99 $X2=0 $Y2=0
cc_125 N_A_105_263#_c_75_n N_VPWR_c_313_n 0.0121867f $X=1.86 $Y=2.99 $X2=0 $Y2=0
cc_126 N_A_105_263#_M1007_g N_VPWR_c_315_n 0.0054895f $X=0.75 $Y=2.465 $X2=0
+ $Y2=0
cc_127 N_A_105_263#_c_80_n N_VPWR_c_316_n 0.0115854f $X=3.455 $Y=2.275 $X2=0
+ $Y2=0
cc_128 N_A_105_263#_M1007_g N_VPWR_c_310_n 0.0110487f $X=0.75 $Y=2.465 $X2=0
+ $Y2=0
cc_129 N_A_105_263#_c_74_n N_VPWR_c_310_n 0.0287839f $X=2.45 $Y=2.99 $X2=0 $Y2=0
cc_130 N_A_105_263#_c_75_n N_VPWR_c_310_n 0.00660921f $X=1.86 $Y=2.99 $X2=0
+ $Y2=0
cc_131 N_A_105_263#_c_80_n N_VPWR_c_310_n 0.0150564f $X=3.455 $Y=2.275 $X2=0
+ $Y2=0
cc_132 N_A_105_263#_c_66_n N_VGND_c_350_n 0.0222877f $X=1.69 $Y=1.54 $X2=0 $Y2=0
cc_133 N_A_105_263#_c_71_n N_VGND_c_350_n 0.00323497f $X=0.69 $Y=1.315 $X2=0
+ $Y2=0
cc_134 N_A_105_263#_c_70_n N_VGND_c_351_n 0.0193955f $X=3.405 $Y=0.87 $X2=0
+ $Y2=0
cc_135 N_A_105_263#_c_71_n N_VGND_c_352_n 0.00438034f $X=0.69 $Y=1.315 $X2=0
+ $Y2=0
cc_136 N_A_105_263#_c_70_n N_VGND_c_356_n 0.00636446f $X=3.405 $Y=0.87 $X2=0
+ $Y2=0
cc_137 N_A_105_263#_c_70_n N_VGND_c_357_n 0.00977043f $X=3.405 $Y=0.87 $X2=0
+ $Y2=0
cc_138 N_A_105_263#_c_71_n N_VGND_c_357_n 0.00838285f $X=0.69 $Y=1.315 $X2=0
+ $Y2=0
cc_139 N_A_219_21#_c_159_n N_TE_B_c_195_n 0.0139283f $X=2.115 $Y=2.42 $X2=0
+ $Y2=0
cc_140 N_A_219_21#_c_155_n N_TE_B_c_196_n 0.00930485f $X=1.17 $Y=0.255 $X2=0
+ $Y2=0
cc_141 N_A_219_21#_c_159_n N_TE_B_M1001_g 0.0216267f $X=2.115 $Y=2.42 $X2=0
+ $Y2=0
cc_142 N_A_219_21#_c_158_n N_TE_B_M1002_g 0.00861458f $X=2.155 $Y=1.1 $X2=0
+ $Y2=0
cc_143 N_A_219_21#_c_159_n N_TE_B_M1002_g 0.0054718f $X=2.115 $Y=2.42 $X2=0
+ $Y2=0
cc_144 N_A_219_21#_c_160_n N_TE_B_M1002_g 0.0014464f $X=1.985 $Y=0.18 $X2=0
+ $Y2=0
cc_145 N_A_219_21#_c_158_n N_TE_B_c_198_n 0.00856211f $X=2.155 $Y=1.1 $X2=0
+ $Y2=0
cc_146 N_A_219_21#_c_159_n N_TE_B_c_198_n 0.0211991f $X=2.115 $Y=2.42 $X2=0
+ $Y2=0
cc_147 N_A_219_21#_c_158_n N_TE_B_c_199_n 0.0101731f $X=2.155 $Y=1.1 $X2=0 $Y2=0
cc_148 N_A_219_21#_c_159_n N_TE_B_c_199_n 0.0492328f $X=2.115 $Y=2.42 $X2=0
+ $Y2=0
cc_149 N_A_219_21#_c_155_n N_Z_c_285_n 0.00225454f $X=1.17 $Y=0.255 $X2=0 $Y2=0
cc_150 N_A_219_21#_c_155_n N_VGND_c_350_n 0.0217899f $X=1.17 $Y=0.255 $X2=0
+ $Y2=0
cc_151 N_A_219_21#_c_156_n N_VGND_c_350_n 0.0186694f $X=1.82 $Y=0.18 $X2=0 $Y2=0
cc_152 N_A_219_21#_c_157_n N_VGND_c_350_n 0.00363087f $X=1.245 $Y=0.18 $X2=0
+ $Y2=0
cc_153 N_A_219_21#_c_158_n N_VGND_c_350_n 0.0403315f $X=2.155 $Y=1.1 $X2=0 $Y2=0
cc_154 N_A_219_21#_c_159_n N_VGND_c_350_n 0.00495424f $X=2.115 $Y=2.42 $X2=0
+ $Y2=0
cc_155 N_A_219_21#_c_160_n N_VGND_c_350_n 0.00146315f $X=1.985 $Y=0.18 $X2=0
+ $Y2=0
cc_156 N_A_219_21#_c_158_n N_VGND_c_351_n 0.0347121f $X=2.155 $Y=1.1 $X2=0 $Y2=0
cc_157 N_A_219_21#_c_160_n N_VGND_c_351_n 0.00386118f $X=1.985 $Y=0.18 $X2=0
+ $Y2=0
cc_158 N_A_219_21#_c_157_n N_VGND_c_352_n 0.00486043f $X=1.245 $Y=0.18 $X2=0
+ $Y2=0
cc_159 N_A_219_21#_c_156_n N_VGND_c_354_n 0.0173548f $X=1.82 $Y=0.18 $X2=0 $Y2=0
cc_160 N_A_219_21#_c_158_n N_VGND_c_354_n 0.0325558f $X=2.155 $Y=1.1 $X2=0 $Y2=0
cc_161 N_A_219_21#_c_156_n N_VGND_c_357_n 0.0150893f $X=1.82 $Y=0.18 $X2=0 $Y2=0
cc_162 N_A_219_21#_c_157_n N_VGND_c_357_n 0.00972445f $X=1.245 $Y=0.18 $X2=0
+ $Y2=0
cc_163 N_A_219_21#_c_158_n N_VGND_c_357_n 0.0241216f $X=2.155 $Y=1.1 $X2=0 $Y2=0
cc_164 N_A_219_21#_c_160_n N_VGND_c_357_n 0.0101306f $X=1.985 $Y=0.18 $X2=0
+ $Y2=0
cc_165 N_TE_B_M1002_g N_A_M1005_g 0.0167532f $X=2.62 $Y=0.87 $X2=0 $Y2=0
cc_166 N_TE_B_M1001_g N_A_M1004_g 0.00890627f $X=2.33 $Y=2.45 $X2=0 $Y2=0
cc_167 N_TE_B_c_198_n N_A_c_251_n 0.0437135f $X=2.615 $Y=1.435 $X2=0 $Y2=0
cc_168 N_TE_B_c_199_n N_A_c_251_n 6.28879e-19 $X=2.615 $Y=1.435 $X2=0 $Y2=0
cc_169 N_TE_B_c_198_n N_A_c_252_n 0.00510719f $X=2.615 $Y=1.435 $X2=0 $Y2=0
cc_170 N_TE_B_c_199_n N_A_c_252_n 0.0437967f $X=2.615 $Y=1.435 $X2=0 $Y2=0
cc_171 N_TE_B_M1000_g N_Z_c_288_n 0.00355139f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_172 N_TE_B_M1000_g N_VPWR_c_311_n 0.0324505f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_173 N_TE_B_c_195_n N_VPWR_c_311_n 0.00471648f $X=2.255 $Y=1.63 $X2=0 $Y2=0
cc_174 N_TE_B_M1000_g N_VPWR_c_315_n 0.00486043f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_175 N_TE_B_M1000_g N_VPWR_c_310_n 0.00827383f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_176 N_TE_B_c_195_n N_VGND_c_350_n 0.00190137f $X=2.255 $Y=1.63 $X2=0 $Y2=0
cc_177 N_TE_B_M1002_g N_VGND_c_351_n 0.00456502f $X=2.62 $Y=0.87 $X2=0 $Y2=0
cc_178 N_TE_B_c_198_n N_VGND_c_351_n 0.00490468f $X=2.615 $Y=1.435 $X2=0 $Y2=0
cc_179 N_TE_B_c_199_n N_VGND_c_351_n 0.00338425f $X=2.615 $Y=1.435 $X2=0 $Y2=0
cc_180 N_TE_B_M1002_g N_VGND_c_354_n 0.00382459f $X=2.62 $Y=0.87 $X2=0 $Y2=0
cc_181 N_TE_B_M1002_g N_VGND_c_357_n 0.00459866f $X=2.62 $Y=0.87 $X2=0 $Y2=0
cc_182 N_A_M1004_g N_VPWR_c_312_n 0.00999043f $X=3.19 $Y=2.45 $X2=0 $Y2=0
cc_183 N_A_M1004_g N_VPWR_c_316_n 0.00435227f $X=3.19 $Y=2.45 $X2=0 $Y2=0
cc_184 N_A_M1004_g N_VPWR_c_310_n 0.00474762f $X=3.19 $Y=2.45 $X2=0 $Y2=0
cc_185 N_A_M1005_g N_VGND_c_351_n 0.00613347f $X=3.19 $Y=0.87 $X2=0 $Y2=0
cc_186 N_A_c_252_n N_VGND_c_351_n 0.00596356f $X=3.25 $Y=1.435 $X2=0 $Y2=0
cc_187 N_A_M1005_g N_VGND_c_356_n 0.00382459f $X=3.19 $Y=0.87 $X2=0 $Y2=0
cc_188 N_A_M1005_g N_VGND_c_357_n 0.00459866f $X=3.19 $Y=0.87 $X2=0 $Y2=0
cc_189 N_Z_c_288_n N_VPWR_c_311_n 0.0416688f $X=0.535 $Y=2 $X2=0 $Y2=0
cc_190 Z N_VPWR_c_315_n 0.0385824f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_191 N_Z_M1007_s N_VPWR_c_310_n 0.00231914f $X=0.39 $Y=1.835 $X2=0 $Y2=0
cc_192 Z N_VPWR_c_310_n 0.0220939f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_193 N_Z_c_285_n N_VGND_c_350_n 0.0265749f $X=0.565 $Y=0.51 $X2=0 $Y2=0
cc_194 N_Z_c_285_n N_VGND_c_352_n 0.0273846f $X=0.565 $Y=0.51 $X2=0 $Y2=0
cc_195 N_Z_c_285_n N_VGND_c_357_n 0.022222f $X=0.565 $Y=0.51 $X2=0 $Y2=0
cc_196 A_165_367# N_VPWR_c_310_n 0.010279f $X=0.825 $Y=1.835 $X2=3.6 $Y2=3.33
