* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor2_4 A B VGND VNB VPB VPWR X
M1000 VPWR A a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.1546e+12p pd=1.854e+07u as=2.4444e+12p ps=2.152e+07u
M1001 a_776_255# B a_1199_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=1.7262e+12p ps=1.534e+07u
M1002 VGND B a_776_255# VNB nshort w=840000u l=150000u
+  ad=2.6208e+12p pd=2.136e+07u as=9.408e+11p ps=8.96e+06u
M1003 VPWR B a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_27_367# a_776_255# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.16e+06u
M1006 VPWR A a_1199_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X B a_110_47# VNB nshort w=840000u l=150000u
+  ad=9.408e+11p pd=8.96e+06u as=9.408e+11p ps=8.96e+06u
M1008 a_776_255# A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_367# a_776_255# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_776_255# B a_1199_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_110_47# A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_776_255# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B a_776_255# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_110_47# B X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A a_776_255# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_776_255# A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X B a_110_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A a_110_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1199_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_776_255# a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1199_367# B a_776_255# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_776_255# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_367# B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_776_255# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1199_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_776_255# B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_776_255# B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND A a_110_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_776_255# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_27_367# B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_110_47# B X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND A a_776_255# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 X a_776_255# a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR A a_1199_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR A a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1199_367# B a_776_255# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_110_47# A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
