* NGSPICE file created from sky130_fd_sc_lp__o311a_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o311a_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR a_96_161# X VPB phighvt w=640000u l=150000u
+  ad=4.736e+11p pd=4.04e+06u as=1.696e+11p ps=1.81e+06u
M1001 a_96_161# C1 VPWR VPB phighvt w=640000u l=150000u
+  ad=3.68e+11p pd=3.71e+06u as=0p ps=0u
M1002 VGND a_96_161# X VNB nshort w=420000u l=150000u
+  ad=2.814e+11p pd=3.02e+06u as=2.541e+11p ps=2.05e+06u
M1003 a_270_481# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=1.92e+11p pd=1.88e+06u as=0p ps=0u
M1004 a_292_55# A3 VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=0p ps=0u
M1005 VGND A2 a_292_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_360_481# A2 a_270_481# VPB phighvt w=640000u l=150000u
+  ad=1.92e+11p pd=1.88e+06u as=0p ps=0u
M1007 a_96_161# A3 a_360_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_564_55# B1 a_292_55# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 VPWR B1 a_96_161# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_96_161# C1 a_564_55# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 a_292_55# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

