# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__ha_m
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__ha_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.050000 2.430000 1.380000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.030000 1.910000 3.290000 2.120000 ;
        RECT 2.960000 1.295000 3.290000 1.910000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.425000 0.470000 4.645000 2.860000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.470000 0.425000 2.490000 ;
        RECT 0.095000 2.490000 1.090000 2.860000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.605000  0.085000 0.795000 0.740000 ;
      RECT 0.605000  1.450000 0.775000 1.950000 ;
      RECT 0.605000  1.950000 1.850000 2.120000 ;
      RECT 0.975000  0.345000 1.300000 0.675000 ;
      RECT 0.975000  0.675000 1.145000 1.950000 ;
      RECT 1.270000  2.430000 1.480000 3.245000 ;
      RECT 1.325000  1.060000 1.495000 1.560000 ;
      RECT 1.325000  1.560000 2.780000 1.730000 ;
      RECT 1.540000  0.345000 1.750000 0.595000 ;
      RECT 1.540000  0.595000 2.770000 0.765000 ;
      RECT 1.680000  2.120000 1.850000 2.360000 ;
      RECT 1.680000  2.360000 2.125000 2.570000 ;
      RECT 1.990000  0.085000 2.320000 0.415000 ;
      RECT 2.560000  0.345000 2.770000 0.595000 ;
      RECT 2.610000  0.945000 3.800000 1.115000 ;
      RECT 2.610000  1.115000 2.780000 1.560000 ;
      RECT 2.790000  2.490000 3.120000 3.245000 ;
      RECT 3.050000  0.795000 3.800000 0.945000 ;
      RECT 3.470000  1.115000 3.800000 3.025000 ;
      RECT 3.995000  0.085000 4.185000 0.935000 ;
      RECT 3.995000  2.125000 4.185000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__ha_m
END LIBRARY
