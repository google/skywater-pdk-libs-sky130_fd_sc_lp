* File: sky130_fd_sc_lp__or4b_m.spice
* Created: Wed Sep  2 10:32:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4b_m.pex.spice"
.subckt sky130_fd_sc_lp__or4b_m  VNB VPB D_N C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_D_N_M1003_g N_A_38_125#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1005 N_A_215_125#_M1005_d N_A_38_125#_M1005_g N_VGND_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.7
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_C_M1006_g N_A_215_125#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.15855 AS=0.0588 PD=1.175 PS=0.7 NRD=15.708 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1002 N_A_215_125#_M1002_d N_B_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.15855 PD=0.7 PS=1.175 NRD=0 NRS=120 M=1 R=2.8 SA=75002
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_A_215_125#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0714 AS=0.0588 PD=0.76 PS=0.7 NRD=8.568 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_X_M1007_d N_A_215_125#_M1007_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0714 PD=1.37 PS=0.76 NRD=0 NRS=8.568 M=1 R=2.8 SA=75002.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_D_N_M1004_g N_A_38_125#_M1004_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_338_397# N_A_38_125#_M1000_g N_A_215_125#_M1000_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1008 A_410_397# N_C_M1008_g A_338_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 A_482_397# N_B_M1009_g A_410_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.9
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g A_482_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=42.1974 NRS=23.443 M=1 R=2.8 SA=75001.3
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_215_125#_M1001_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=9.3772 M=1 R=2.8 SA=75001.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__or4b_m.pxi.spice"
*
.ends
*
*
