* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__srsdfstp_1 CLK D SCD SCE SET_B SLEEP_B KAPWR VGND VNB VPB
+ VPWR Q
X0 a_1656_125# a_689_139# a_1728_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_2002_125# a_1972_99# a_2074_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_3466_403# a_1728_125# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_3466_403# a_1728_125# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_2216_99# a_2074_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_3466_403# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_3056_72# SLEEP_B a_3134_72# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_27_481# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_1336_97# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1728_125# a_659_113# a_1930_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_887_139# a_659_113# a_1132_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND a_659_113# a_689_139# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_3134_72# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1132_535# a_1068_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 VGND SLEEP_B a_3292_72# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1728_125# a_689_139# a_2862_414# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_2074_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR SCE a_213_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_1068_21# a_887_139# a_1336_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 KAPWR a_2216_99# a_2658_414# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 a_1541_125# a_659_113# a_1712_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_1712_451# a_659_113# a_1728_125# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 a_2463_119# a_1728_125# a_1972_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_3466_403# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_1930_125# a_1972_99# a_2002_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_2658_414# SET_B a_1728_125# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X26 a_659_113# CLK a_3056_72# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_887_139# a_689_139# a_996_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VGND a_1728_125# a_2463_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_111_119# SCE a_189_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VPWR a_887_139# a_1541_125# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X31 a_1541_125# a_689_139# a_1656_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 a_2862_414# a_1972_99# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X33 a_1068_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X34 a_275_119# a_339_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 VGND a_887_139# a_1541_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X36 a_1972_99# a_1728_125# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X37 KAPWR SLEEP_B a_2216_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X38 VPWR a_659_113# a_689_139# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X39 VGND SCD a_111_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VPWR a_887_139# a_1068_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X41 a_3292_72# SLEEP_B a_2216_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_189_119# a_339_93# a_27_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X43 a_189_119# a_689_139# a_887_139# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X44 a_996_73# a_1068_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 KAPWR CLK a_659_113# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X46 a_659_113# SLEEP_B KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X47 a_213_481# D a_189_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X48 a_339_93# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X49 a_189_119# D a_275_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X50 a_339_93# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X51 a_189_119# a_659_113# a_887_139# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
