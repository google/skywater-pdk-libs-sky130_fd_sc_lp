* File: sky130_fd_sc_lp__mux2i_1.pex.spice
* Created: Wed Sep  2 10:01:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2I_1%A0 3 7 9 13 14
c30 14 0 1.34632e-19 $X=0.505 $Y=1.51
r31 12 14 20.2947 $w=2.85e-07 $l=1.2e-07 $layer=POLY_cond $X=0.385 $Y=1.51
+ $X2=0.505 $Y2=1.51
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.51 $X2=0.385 $Y2=1.51
r33 9 13 4.63971 $w=3.83e-07 $l=1.55e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.51
r34 5 14 20.2947 $w=2.85e-07 $l=2.16852e-07 $layer=POLY_cond $X=0.625 $Y=1.675
+ $X2=0.505 $Y2=1.51
r35 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.625 $Y=1.675
+ $X2=0.625 $Y2=2.465
r36 1 14 17.7656 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.345
+ $X2=0.505 $Y2=1.51
r37 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.505 $Y=1.345
+ $X2=0.505 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_1%A1 3 7 9 12 13
c36 13 0 1.34632e-19 $X=1.145 $Y=1.51
c37 12 0 1.66137e-19 $X=1.145 $Y=1.51
r38 12 15 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=1.51 $X2=1.11
+ $Y2=1.675
r39 12 14 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=1.51 $X2=1.11
+ $Y2=1.345
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.145
+ $Y=1.51 $X2=1.145 $Y2=1.51
r41 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.145 $Y=1.665
+ $X2=1.145 $Y2=1.51
r42 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.105 $Y=2.465
+ $X2=1.105 $Y2=1.675
r43 3 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.985 $Y=0.785
+ $X2=0.985 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_1%A_304_237# 1 2 9 11 13 14 17 21 27 30 31 32
r67 30 31 3.84343 $w=2.4e-07 $l=9.44722e-08 $layer=LI1_cond $X=3.095 $Y=1.415
+ $X2=3.075 $Y2=1.5
r68 30 32 16.7628 $w=2.18e-07 $l=3.2e-07 $layer=LI1_cond $X=3.095 $Y=1.415
+ $X2=3.095 $Y2=1.095
r69 25 32 6.06832 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.115 $Y=0.965
+ $X2=3.115 $Y2=1.095
r70 25 27 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=3.115 $Y=0.965
+ $X2=3.115 $Y2=0.525
r71 21 23 38.3409 $w=2.58e-07 $l=8.65e-07 $layer=LI1_cond $X=3.075 $Y=2.045
+ $X2=3.075 $Y2=2.91
r72 19 31 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=1.585
+ $X2=3.075 $Y2=1.5
r73 19 21 20.3894 $w=2.58e-07 $l=4.6e-07 $layer=LI1_cond $X=3.075 $Y=1.585
+ $X2=3.075 $Y2=2.045
r74 17 33 11.0946 $w=3.91e-07 $l=9e-08 $layer=POLY_cond $X=1.685 $Y=1.425
+ $X2=1.595 $Y2=1.425
r75 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.685
+ $Y=1.5 $X2=1.685 $Y2=1.5
r76 14 31 2.60907 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.945 $Y=1.5
+ $X2=3.075 $Y2=1.5
r77 14 16 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=2.945 $Y=1.5
+ $X2=1.685 $Y2=1.5
r78 11 17 34.5166 $w=3.91e-07 $l=3.81576e-07 $layer=POLY_cond $X=1.965 $Y=1.185
+ $X2=1.685 $Y2=1.425
r79 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.965 $Y=1.185
+ $X2=1.965 $Y2=0.655
r80 7 33 25.3065 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.595 $Y=1.665
+ $X2=1.595 $Y2=1.425
r81 7 9 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.595 $Y=1.665 $X2=1.595
+ $Y2=2.465
r82 2 23 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.835 $X2=3.11 $Y2=2.91
r83 2 21 400 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.835 $X2=3.11 $Y2=2.045
r84 1 27 91 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=2 $X=3.025
+ $Y=0.345 $X2=3.15 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_1%S 1 3 6 8 9 12 15 19 20 24 26 28
r55 24 26 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=3.447 $Y=1.46
+ $X2=3.447 $Y2=1.295
r56 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.48
+ $Y=1.46 $X2=3.48 $Y2=1.46
r57 20 25 6.21713 $w=3.78e-07 $l=2.05e-07 $layer=LI1_cond $X=3.565 $Y=1.665
+ $X2=3.565 $Y2=1.46
r58 19 25 5.00403 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=3.565 $Y=1.295
+ $X2=3.565 $Y2=1.46
r59 16 18 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.215 $Y=1.65
+ $X2=2.395 $Y2=1.65
r60 15 26 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.365 $Y=0.765
+ $X2=3.365 $Y2=1.295
r61 12 28 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.325 $Y=2.465
+ $X2=3.325 $Y2=1.725
r62 9 18 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.47 $Y=1.65
+ $X2=2.395 $Y2=1.65
r63 8 28 32.8921 $w=3.95e-07 $l=7.5e-08 $layer=POLY_cond $X=3.447 $Y=1.65
+ $X2=3.447 $Y2=1.725
r64 8 24 26.7517 $w=3.95e-07 $l=1.9e-07 $layer=POLY_cond $X=3.447 $Y=1.65
+ $X2=3.447 $Y2=1.46
r65 8 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.25 $Y=1.65 $X2=2.47
+ $Y2=1.65
r66 4 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.395 $Y=1.575
+ $X2=2.395 $Y2=1.65
r67 4 6 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=2.395 $Y=1.575
+ $X2=2.395 $Y2=0.655
r68 1 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.215 $Y=1.725
+ $X2=2.215 $Y2=1.65
r69 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.215 $Y=1.725
+ $X2=2.215 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_1%A_52_367# 1 2 9 13 16 17 18 19 21 24
c50 13 0 1.66137e-19 $X=1.455 $Y=2.43
r51 19 26 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=1.985
+ $X2=2.445 $Y2=1.9
r52 19 21 35.5337 $w=2.98e-07 $l=9.25e-07 $layer=LI1_cond $X=2.445 $Y=1.985
+ $X2=2.445 $Y2=2.91
r53 17 26 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.295 $Y=1.9
+ $X2=2.445 $Y2=1.9
r54 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.295 $Y=1.9
+ $X2=1.625 $Y2=1.9
r55 15 18 6.9061 $w=1.67e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.54 $Y=1.985
+ $X2=1.625 $Y2=1.9
r56 15 16 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.54 $Y=1.985
+ $X2=1.54 $Y2=2.31
r57 14 24 2.15711 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=2.43
+ $X2=0.365 $Y2=2.43
r58 13 16 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.455 $Y=2.43
+ $X2=1.54 $Y2=2.31
r59 13 14 44.4171 $w=2.38e-07 $l=9.25e-07 $layer=LI1_cond $X=1.455 $Y=2.43
+ $X2=0.53 $Y2=2.43
r60 7 24 4.27425 $w=3e-07 $l=1.34164e-07 $layer=LI1_cond $X=0.335 $Y=2.31
+ $X2=0.365 $Y2=2.43
r61 7 9 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.335 $Y=2.31
+ $X2=0.335 $Y2=2.095
r62 2 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=1.98
r63 2 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=2.91
r64 1 24 300 $w=1.7e-07 $l=7.26137e-07 $layer=licon1_PDIFF $count=2 $X=0.26
+ $Y=1.835 $X2=0.41 $Y2=2.49
r65 1 9 600 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.835 $X2=0.385 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_1%Y 1 2 7 9 12 13 14
r30 14 17 19.013 $w=2.08e-07 $l=3.6e-07 $layer=LI1_cond $X=1.2 $Y=2.035 $X2=0.84
+ $Y2=2.035
r31 13 17 1.58442 $w=2.08e-07 $l=3e-08 $layer=LI1_cond $X=0.81 $Y=2.035 $X2=0.84
+ $Y2=2.035
r32 12 13 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.725 $Y=1.93
+ $X2=0.81 $Y2=2.035
r33 11 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.725 $Y=1.175
+ $X2=0.725 $Y2=1.93
r34 7 11 6.56923 $w=3.25e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.72 $Y=1
+ $X2=0.725 $Y2=1.175
r35 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.72 $Y=1 $X2=0.72
+ $Y2=0.68
r36 2 17 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=0.7
+ $Y=1.835 $X2=0.84 $Y2=2.035
r37 1 9 91 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=2 $X=0.58
+ $Y=0.365 $X2=0.72 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_1%VPWR 1 2 9 13 15 20 21 22 31 40
r39 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r40 37 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r41 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r44 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 31 39 4.69206 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.607 $Y2=3.33
r46 31 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 26 30 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 25 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 22 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 22 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 20 29 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.96 $Y2=3.33
r55 19 33 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=1.96 $Y2=3.33
r57 15 18 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=3.54 $Y=2.005
+ $X2=3.54 $Y2=2.95
r58 13 39 3.07411 $w=3.3e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.607 $Y2=3.33
r59 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.54 $Y2=2.95
r60 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.96 $Y=2.24 $X2=1.96
+ $Y2=2.95
r61 7 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=3.245 $X2=1.96
+ $Y2=3.33
r62 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=2.95
r63 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.835 $X2=3.54 $Y2=2.95
r64 2 15 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=3.4
+ $Y=1.835 $X2=3.54 $Y2=2.005
r65 1 12 400 $w=1.7e-07 $l=1.25163e-06 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.835 $X2=1.96 $Y2=2.95
r66 1 9 400 $w=1.7e-07 $l=5.30542e-07 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.835 $X2=1.96 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_1%A_29_73# 1 2 9 11 12 16
r25 11 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=0.34
+ $X2=1.75 $Y2=0.34
r26 11 12 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=1.585 $Y=0.34
+ $X2=0.385 $Y2=0.34
r27 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.245 $Y=0.425
+ $X2=0.385 $Y2=0.34
r28 7 9 3.49849 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=0.425
+ $X2=0.245 $Y2=0.51
r29 2 16 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.625
+ $Y=0.235 $X2=1.75 $Y2=0.38
r30 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.365 $X2=0.27 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_1%A_212_73# 1 2 9 11 12 15
r31 13 15 26.486 $w=2.83e-07 $l=6.55e-07 $layer=LI1_cond $X=2.632 $Y=1.075
+ $X2=2.632 $Y2=0.42
r32 11 13 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=2.49 $Y=1.16
+ $X2=2.632 $Y2=1.075
r33 11 12 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.49 $Y=1.16
+ $X2=1.385 $Y2=1.16
r34 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.22 $Y=1.075
+ $X2=1.385 $Y2=1.16
r35 7 9 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=1.22 $Y=1.075
+ $X2=1.22 $Y2=0.68
r36 2 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.47
+ $Y=0.235 $X2=2.61 $Y2=0.42
r37 1 9 91 $w=1.7e-07 $l=3.86814e-07 $layer=licon1_NDIFF $count=2 $X=1.06
+ $Y=0.365 $X2=1.22 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_1%VGND 1 2 9 11 13 15 17 22 28 32
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r37 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r39 26 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r40 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 23 28 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.195
+ $Y2=0
r42 23 25 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=3.12
+ $Y2=0
r43 22 31 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.627
+ $Y2=0
r44 22 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.12
+ $Y2=0
r45 19 20 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 17 28 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.195
+ $Y2=0
r47 17 19 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=2.085 $Y=0
+ $X2=0.24 $Y2=0
r48 15 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r49 15 20 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.24
+ $Y2=0
r50 11 31 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.627 $Y2=0
r51 11 13 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.58 $Y=0.085
+ $X2=3.58 $Y2=0.49
r52 7 28 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0
r53 7 9 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0.38
r54 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.44
+ $Y=0.345 $X2=3.58 $Y2=0.49
r55 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.04
+ $Y=0.235 $X2=2.18 $Y2=0.38
.ends

