* File: sky130_fd_sc_lp__dlrtp_1.pex.spice
* Created: Wed Sep  2 09:47:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRTP_1%D 2 5 9 10 11 12 13 18 20
c35 20 0 9.81893e-20 $X=0.677 $Y=0.88
c36 11 0 1.28937e-19 $X=0.72 $Y=0.925
r37 18 20 46.0284 $w=4.15e-07 $l=1.65e-07 $layer=POLY_cond $X=0.677 $Y=1.045
+ $X2=0.677 $Y2=0.88
r38 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.72
+ $Y=1.045 $X2=0.72 $Y2=1.045
r39 12 13 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.665
r40 12 19 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.045
r41 11 19 5.76222 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.745 $Y=0.925
+ $X2=0.745 $Y2=1.045
r42 9 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.585 $Y=0.56
+ $X2=0.585 $Y2=0.88
r43 5 10 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=0.545 $Y=2.64
+ $X2=0.545 $Y2=1.55
r44 2 10 51.6569 $w=4.15e-07 $l=2.07e-07 $layer=POLY_cond $X=0.677 $Y=1.343
+ $X2=0.677 $Y2=1.55
r45 1 18 5.62854 $w=4.15e-07 $l=4.2e-08 $layer=POLY_cond $X=0.677 $Y=1.087
+ $X2=0.677 $Y2=1.045
r46 1 2 34.3073 $w=4.15e-07 $l=2.56e-07 $layer=POLY_cond $X=0.677 $Y=1.087
+ $X2=0.677 $Y2=1.343
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%GATE 3 5 8 10 11 12 13 18 20
c42 20 0 1.28937e-19 $X=1.265 $Y=0.88
c43 11 0 9.81893e-20 $X=1.2 $Y=0.925
r44 18 20 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.265 $Y=1.045
+ $X2=1.265 $Y2=0.88
r45 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.27
+ $Y=1.045 $X2=1.27 $Y2=1.045
r46 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=1.295
+ $X2=1.205 $Y2=1.665
r47 12 19 8.47385 $w=3.38e-07 $l=2.5e-07 $layer=LI1_cond $X=1.205 $Y=1.295
+ $X2=1.205 $Y2=1.045
r48 11 19 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=1.205 $Y=0.925
+ $X2=1.205 $Y2=1.045
r49 8 10 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=1.17 $Y=2.64
+ $X2=1.17 $Y2=1.55
r50 5 10 47.1551 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=1.265 $Y=1.38
+ $X2=1.265 $Y2=1.55
r51 4 18 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=1.265 $Y=1.05
+ $X2=1.265 $Y2=1.045
r52 4 5 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=1.265 $Y=1.05 $X2=1.265
+ $Y2=1.38
r53 3 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.17 $Y=0.56 $X2=1.17
+ $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%A_249_70# 1 2 8 11 13 15 18 20 21 24 26 27
+ 30 34 36 39 43 48 50 59 60 68
c145 68 0 7.96279e-20 $X=2.43 $Y=0.93
c146 39 0 1.63114e-19 $X=3.74 $Y=1.175
c147 36 0 1.934e-19 $X=3.655 $Y=0.79
c148 26 0 1.17006e-19 $X=2.12 $Y=1.995
c149 24 0 1.54858e-19 $X=3.76 $Y=0.445
r150 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.85
+ $Y=1.34 $X2=3.85 $Y2=1.34
r151 56 59 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=3.74 $Y=1.305
+ $X2=3.85 $Y2=1.305
r152 54 68 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.41 $Y=0.93 $X2=2.43
+ $Y2=0.93
r153 54 65 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.41 $Y=0.93
+ $X2=2.195 $Y2=0.93
r154 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=0.93 $X2=2.41 $Y2=0.93
r155 50 53 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.41 $Y=0.79
+ $X2=2.41 $Y2=0.93
r156 46 48 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.44 $Y=2.57
+ $X2=1.635 $Y2=2.57
r157 41 43 8.47385 $w=3.38e-07 $l=2.5e-07 $layer=LI1_cond $X=1.385 $Y=0.5
+ $X2=1.635 $Y2=0.5
r158 39 56 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.74 $Y=1.175
+ $X2=3.74 $Y2=1.305
r159 38 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.74 $Y=0.875
+ $X2=3.74 $Y2=1.175
r160 37 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0.79
+ $X2=2.41 $Y2=0.79
r161 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.655 $Y=0.79
+ $X2=3.74 $Y2=0.875
r162 36 37 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=3.655 $Y=0.79
+ $X2=2.575 $Y2=0.79
r163 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.995 $X2=1.63 $Y2=1.995
r164 32 48 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.635 $Y=2.405
+ $X2=1.635 $Y2=2.57
r165 32 34 25.2626 $w=1.78e-07 $l=4.1e-07 $layer=LI1_cond $X=1.635 $Y=2.405
+ $X2=1.635 $Y2=1.995
r166 31 43 4.46199 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=1.635 $Y=0.67
+ $X2=1.635 $Y2=0.5
r167 31 34 81.6414 $w=1.78e-07 $l=1.325e-06 $layer=LI1_cond $X=1.635 $Y=0.67
+ $X2=1.635 $Y2=1.995
r168 30 60 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=3.85 $Y=1.515
+ $X2=3.85 $Y2=1.34
r169 29 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.85 $Y=1.175
+ $X2=3.85 $Y2=1.34
r170 26 35 85.682 $w=3.3e-07 $l=4.9e-07 $layer=POLY_cond $X=2.12 $Y=1.995
+ $X2=1.63 $Y2=1.995
r171 26 27 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.995
+ $X2=2.195 $Y2=1.995
r172 24 29 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.76 $Y=0.445
+ $X2=3.76 $Y2=1.175
r173 20 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.685 $Y=1.59
+ $X2=3.85 $Y2=1.515
r174 20 21 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.685 $Y=1.59
+ $X2=3.475 $Y2=1.59
r175 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.4 $Y=1.665
+ $X2=3.475 $Y2=1.59
r176 16 18 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.4 $Y=1.665
+ $X2=3.4 $Y2=2.685
r177 13 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=0.765
+ $X2=2.43 $Y2=0.93
r178 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.43 $Y=0.765
+ $X2=2.43 $Y2=0.445
r179 9 27 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=2.16
+ $X2=2.195 $Y2=1.995
r180 9 11 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.195 $Y=2.16
+ $X2=2.195 $Y2=2.685
r181 8 27 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.83
+ $X2=2.195 $Y2=1.995
r182 7 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.095
+ $X2=2.195 $Y2=0.93
r183 7 8 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=2.195 $Y=1.095
+ $X2=2.195 $Y2=1.83
r184 2 46 600 $w=1.7e-07 $l=3.33542e-07 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=2.32 $X2=1.44 $Y2=2.57
r185 1 41 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.245
+ $Y=0.35 $X2=1.385 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%A_41_464# 1 2 11 15 17 18 21 25 27 30 31 32
+ 34 35 37 38
c98 30 0 1.17006e-19 $X=1.1 $Y=2.905
r99 38 42 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=2.707 $Y=1.7
+ $X2=2.707 $Y2=1.535
r100 37 40 16.5175 $w=5.58e-07 $l=4.75e-07 $layer=LI1_cond $X=2.53 $Y=1.7
+ $X2=2.53 $Y2=2.175
r101 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.645
+ $Y=1.7 $X2=2.645 $Y2=1.7
r102 34 40 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.335 $Y=2.905
+ $X2=2.335 $Y2=2.175
r103 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.25 $Y=2.99
+ $X2=2.335 $Y2=2.905
r104 31 32 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=2.25 $Y=2.99
+ $X2=1.185 $Y2=2.99
r105 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.1 $Y=2.905
+ $X2=1.185 $Y2=2.99
r106 29 30 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.1 $Y=2.13
+ $X2=1.1 $Y2=2.905
r107 28 35 3.3199 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.455 $Y=2.045
+ $X2=0.31 $Y2=2.045
r108 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.015 $Y=2.045
+ $X2=1.1 $Y2=2.13
r109 27 28 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.015 $Y=2.045
+ $X2=0.455 $Y2=2.045
r110 23 35 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.31 $Y=2.13
+ $X2=0.31 $Y2=2.045
r111 23 25 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=0.31 $Y=2.13
+ $X2=0.31 $Y2=2.465
r112 19 35 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.31 $Y=1.96
+ $X2=0.31 $Y2=2.045
r113 19 21 55.8339 $w=2.88e-07 $l=1.405e-06 $layer=LI1_cond $X=0.31 $Y=1.96
+ $X2=0.31 $Y2=0.555
r114 17 18 45.2433 $w=4.55e-07 $l=1.5e-07 $layer=POLY_cond $X=2.797 $Y=2.055
+ $X2=2.797 $Y2=2.205
r115 15 18 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.04 $Y=2.685
+ $X2=3.04 $Y2=2.205
r116 11 42 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=2.86 $Y=0.445
+ $X2=2.86 $Y2=1.535
r117 7 38 7.57836 $w=4.55e-07 $l=6.2e-08 $layer=POLY_cond $X=2.707 $Y=1.762
+ $X2=2.707 $Y2=1.7
r118 7 17 35.8139 $w=4.55e-07 $l=2.93e-07 $layer=POLY_cond $X=2.707 $Y=1.762
+ $X2=2.707 $Y2=2.055
r119 2 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.205
+ $Y=2.32 $X2=0.33 $Y2=2.465
r120 1 21 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.35 $X2=0.37 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%A_371_473# 1 2 9 13 16 19 21 24 25 26 28 32
+ 34 35 38 41 43
c116 38 0 1.32117e-19 $X=3.31 $Y=1.14
c117 35 0 1.54858e-19 $X=3.075 $Y=1.205
c118 25 0 7.91208e-20 $X=3.88 $Y=2.99
c119 21 0 3.02476e-20 $X=2.99 $Y=1.28
r120 41 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=2.04
+ $X2=3.855 $Y2=2.205
r121 40 43 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=3.855 $Y=2.075
+ $X2=3.965 $Y2=2.075
r122 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.855
+ $Y=2.04 $X2=3.855 $Y2=2.04
r123 38 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.14
+ $X2=3.31 $Y2=0.975
r124 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.31
+ $Y=1.14 $X2=3.31 $Y2=1.14
r125 35 37 10.5404 $w=2.72e-07 $l=2.35e-07 $layer=LI1_cond $X=3.075 $Y=1.205
+ $X2=3.31 $Y2=1.205
r126 29 32 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=1.985 $Y=0.395
+ $X2=2.195 $Y2=0.395
r127 27 43 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.965 $Y=2.205
+ $X2=3.965 $Y2=2.075
r128 27 28 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.965 $Y=2.205
+ $X2=3.965 $Y2=2.905
r129 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.88 $Y=2.99
+ $X2=3.965 $Y2=2.905
r130 25 26 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.88 $Y=2.99
+ $X2=3.16 $Y2=2.99
r131 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.075 $Y=2.905
+ $X2=3.16 $Y2=2.99
r132 23 35 3.48705 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.075 $Y=1.365
+ $X2=3.075 $Y2=1.205
r133 23 24 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=3.075 $Y=1.365
+ $X2=3.075 $Y2=2.905
r134 22 34 1.59926 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=2.08 $Y=1.28
+ $X2=1.987 $Y2=1.28
r135 21 35 5.51876 $w=2.72e-07 $l=1.16619e-07 $layer=LI1_cond $X=2.99 $Y=1.28
+ $X2=3.075 $Y2=1.205
r136 21 22 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.99 $Y=1.28
+ $X2=2.08 $Y2=1.28
r137 17 34 4.86787 $w=1.82e-07 $l=8.5e-08 $layer=LI1_cond $X=1.987 $Y=1.365
+ $X2=1.987 $Y2=1.28
r138 17 19 72.2408 $w=1.83e-07 $l=1.205e-06 $layer=LI1_cond $X=1.987 $Y=1.365
+ $X2=1.987 $Y2=2.57
r139 16 34 4.86787 $w=1.82e-07 $l=8.59942e-08 $layer=LI1_cond $X=1.985 $Y=1.195
+ $X2=1.987 $Y2=1.28
r140 15 29 3.32261 $w=1.8e-07 $l=1.4e-07 $layer=LI1_cond $X=1.985 $Y=0.535
+ $X2=1.985 $Y2=0.395
r141 15 16 40.6667 $w=1.78e-07 $l=6.6e-07 $layer=LI1_cond $X=1.985 $Y=0.535
+ $X2=1.985 $Y2=1.195
r142 13 50 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.925 $Y=2.575
+ $X2=3.925 $Y2=2.205
r143 9 46 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.22 $Y=0.445
+ $X2=3.22 $Y2=0.975
r144 2 19 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=2.365 $X2=1.98 $Y2=2.57
r145 1 32 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.235 $X2=2.195 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%A_809_21# 1 2 7 9 14 18 22 26 28 31 35 38 39
+ 41 43 46 47 54 55 58
c123 46 0 3.37142e-20 $X=6.005 $Y=2.3
c124 39 0 1.35653e-19 $X=5.405 $Y=2.47
c125 26 0 1.63114e-19 $X=4.305 $Y=0.84
c126 14 0 7.91208e-20 $X=4.315 $Y=2.575
c127 7 0 1.934e-19 $X=4.12 $Y=0.765
r128 55 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.505
+ $X2=6.195 $Y2=1.67
r129 55 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.505
+ $X2=6.195 $Y2=1.34
r130 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.195
+ $Y=1.505 $X2=6.195 $Y2=1.505
r131 51 54 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.005 $Y=1.505
+ $X2=6.195 $Y2=1.505
r132 48 50 14.1648 $w=2.67e-07 $l=3.1e-07 $layer=LI1_cond $X=5.255 $Y=2.075
+ $X2=5.255 $Y2=2.385
r133 45 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.005 $Y=1.67
+ $X2=6.005 $Y2=1.505
r134 45 46 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.005 $Y=1.67
+ $X2=6.005 $Y2=2.3
r135 44 50 3.37873 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=5.555 $Y=2.385
+ $X2=5.255 $Y2=2.385
r136 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.92 $Y=2.385
+ $X2=6.005 $Y2=2.3
r137 43 44 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.92 $Y=2.385
+ $X2=5.555 $Y2=2.385
r138 39 50 3.63317 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=5.405 $Y=2.47
+ $X2=5.255 $Y2=2.385
r139 39 41 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=5.405 $Y=2.47
+ $X2=5.405 $Y2=2.91
r140 38 48 7.54419 $w=2.67e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.17 $Y=1.945
+ $X2=5.255 $Y2=2.075
r141 38 47 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.17 $Y=1.945
+ $X2=5.17 $Y2=1.165
r142 33 47 9.32938 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=5.065 $Y=0.975
+ $X2=5.065 $Y2=1.165
r143 33 35 14.1023 $w=3.78e-07 $l=4.65e-07 $layer=LI1_cond $X=5.065 $Y=0.975
+ $X2=5.065 $Y2=0.51
r144 31 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=2.04
+ $X2=4.395 $Y2=2.205
r145 31 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=2.04
+ $X2=4.395 $Y2=1.875
r146 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=2.04 $X2=4.395 $Y2=2.04
r147 28 48 0.877981 $w=2.6e-07 $l=1.7e-07 $layer=LI1_cond $X=5.085 $Y=2.075
+ $X2=5.255 $Y2=2.075
r148 28 30 30.5841 $w=2.58e-07 $l=6.9e-07 $layer=LI1_cond $X=5.085 $Y=2.075
+ $X2=4.395 $Y2=2.075
r149 24 26 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=4.12 $Y=0.84
+ $X2=4.305 $Y2=0.84
r150 22 62 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=6.14 $Y=2.465
+ $X2=6.14 $Y2=1.67
r151 18 61 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.105 $Y=0.785
+ $X2=6.105 $Y2=1.34
r152 14 59 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.315 $Y=2.575
+ $X2=4.315 $Y2=2.205
r153 10 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.305 $Y=0.915
+ $X2=4.305 $Y2=0.84
r154 10 58 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=4.305 $Y=0.915
+ $X2=4.305 $Y2=1.875
r155 7 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.12 $Y=0.765
+ $X2=4.12 $Y2=0.84
r156 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.12 $Y=0.765
+ $X2=4.12 $Y2=0.445
r157 2 50 600 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.835 $X2=5.42 $Y2=2.385
r158 2 41 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.835 $X2=5.42 $Y2=2.91
r159 1 35 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.865
+ $Y=0.365 $X2=4.99 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%A_659_47# 1 2 9 13 15 16 18 19 23 24 26 27
+ 28 34 37 39
c106 24 0 1.32117e-19 $X=3.51 $Y=1.69
r107 37 40 5.76222 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=4.725 $Y=1.5
+ $X2=4.725 $Y2=1.69
r108 37 39 8.5712 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=1.5
+ $X2=4.725 $Y2=1.335
r109 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.83
+ $Y=1.5 $X2=4.83 $Y2=1.5
r110 31 34 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.425 $Y=2.57
+ $X2=3.615 $Y2=2.57
r111 29 39 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.62 $Y=0.895
+ $X2=4.62 $Y2=1.335
r112 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.535 $Y=0.81
+ $X2=4.62 $Y2=0.895
r113 27 28 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.535 $Y=0.81
+ $X2=4.175 $Y2=0.81
r114 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.09 $Y=0.725
+ $X2=4.175 $Y2=0.81
r115 25 26 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.09 $Y=0.535
+ $X2=4.09 $Y2=0.725
r116 23 40 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.535 $Y=1.69
+ $X2=4.725 $Y2=1.69
r117 23 24 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=4.535 $Y=1.69
+ $X2=3.51 $Y2=1.69
r118 19 25 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.005 $Y=0.425
+ $X2=4.09 $Y2=0.535
r119 19 21 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=4.005 $Y=0.425
+ $X2=3.545 $Y2=0.425
r120 18 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=2.405
+ $X2=3.425 $Y2=2.57
r121 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.425 $Y=1.775
+ $X2=3.51 $Y2=1.69
r122 17 18 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.425 $Y=1.775
+ $X2=3.425 $Y2=2.405
r123 15 38 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=5.13 $Y=1.5 $X2=4.83
+ $Y2=1.5
r124 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.13 $Y=1.5
+ $X2=5.205 $Y2=1.5
r125 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.205 $Y=1.665
+ $X2=5.205 $Y2=1.5
r126 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.205 $Y=1.665
+ $X2=5.205 $Y2=2.465
r127 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.205 $Y=1.335
+ $X2=5.205 $Y2=1.5
r128 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.205 $Y=1.335
+ $X2=5.205 $Y2=0.785
r129 2 34 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=2.365 $X2=3.615 $Y2=2.57
r130 1 21 182 $w=1.7e-07 $l=3.29773e-07 $layer=licon1_NDIFF $count=1 $X=3.295
+ $Y=0.235 $X2=3.545 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%RESET_B 3 7 9 10 11 12 13 21 22 33
c48 21 0 1.69368e-19 $X=5.655 $Y=1.51
r49 33 42 3.08081 $w=1.78e-07 $l=5e-08 $layer=LI1_cond $X=5.515 $Y=1.295
+ $X2=5.515 $Y2=1.345
r50 22 34 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=5.582 $Y=1.51
+ $X2=5.582 $Y2=1.502
r51 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.655 $Y=1.51
+ $X2=5.655 $Y2=1.675
r52 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.655 $Y=1.51
+ $X2=5.655 $Y2=1.345
r53 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.655
+ $Y=1.51 $X2=5.655 $Y2=1.51
r54 12 13 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=5.582 $Y=1.665
+ $X2=5.582 $Y2=2.035
r55 12 22 5.67075 $w=3.13e-07 $l=1.55e-07 $layer=LI1_cond $X=5.582 $Y=1.665
+ $X2=5.582 $Y2=1.51
r56 11 34 5.12197 $w=3.13e-07 $l=1.4e-07 $layer=LI1_cond $X=5.582 $Y=1.362
+ $X2=5.582 $Y2=1.502
r57 11 42 2.72101 $w=3.13e-07 $l=1.7e-08 $layer=LI1_cond $X=5.582 $Y=1.362
+ $X2=5.582 $Y2=1.345
r58 11 33 1.10909 $w=1.78e-07 $l=1.8e-08 $layer=LI1_cond $X=5.515 $Y=1.277
+ $X2=5.515 $Y2=1.295
r59 10 11 21.6889 $w=1.78e-07 $l=3.52e-07 $layer=LI1_cond $X=5.515 $Y=0.925
+ $X2=5.515 $Y2=1.277
r60 9 10 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=5.515 $Y=0.555
+ $X2=5.515 $Y2=0.925
r61 7 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.635 $Y=2.465
+ $X2=5.635 $Y2=1.675
r62 3 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.565 $Y=0.785
+ $X2=5.565 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%VPWR 1 2 3 4 17 21 25 28 29 30 32 37 50 51
+ 54 57 64
r82 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r83 62 64 9.43299 $w=6.79e-07 $l=5.25e-07 $layer=LI1_cond $X=4.725 $Y=2.805
+ $X2=4.725 $Y2=3.33
r84 60 62 4.31222 $w=6.79e-07 $l=2.4e-07 $layer=LI1_cond $X=4.725 $Y=2.565
+ $X2=4.725 $Y2=2.805
r85 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r86 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r88 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r89 48 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r91 45 64 9.12129 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=5.085 $Y=3.33
+ $X2=4.725 $Y2=3.33
r92 45 47 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.085 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 44 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 41 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r96 40 43 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33 $X2=4.08
+ $Y2=3.33
r97 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r98 38 57 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.705 $Y2=3.33
r99 38 40 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.82 $Y=3.33 $X2=3.12
+ $Y2=3.33
r100 37 64 9.12129 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.725 $Y2=3.33
r101 37 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.08 $Y2=3.33
r102 36 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 33 54 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.845 $Y=3.33
+ $X2=0.75 $Y2=3.33
r106 33 35 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.845 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 32 57 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.59 $Y=3.33
+ $X2=2.705 $Y2=3.33
r108 32 35 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=2.59 $Y=3.33
+ $X2=1.2 $Y2=3.33
r109 30 44 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r110 30 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r111 28 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.725 $Y=3.33
+ $X2=5.52 $Y2=3.33
r112 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=3.33
+ $X2=5.89 $Y2=3.33
r113 27 50 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.055 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.055 $Y=3.33
+ $X2=5.89 $Y2=3.33
r115 23 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.89 $Y=3.245
+ $X2=5.89 $Y2=3.33
r116 23 25 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=5.89 $Y=3.245
+ $X2=5.89 $Y2=2.76
r117 19 57 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=3.245
+ $X2=2.705 $Y2=3.33
r118 19 21 36.8281 $w=2.28e-07 $l=7.35e-07 $layer=LI1_cond $X=2.705 $Y=3.245
+ $X2=2.705 $Y2=2.51
r119 15 54 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=3.245
+ $X2=0.75 $Y2=3.33
r120 15 17 45.5311 $w=1.88e-07 $l=7.8e-07 $layer=LI1_cond $X=0.75 $Y=3.245
+ $X2=0.75 $Y2=2.465
r121 4 25 600 $w=1.7e-07 $l=1.011e-06 $layer=licon1_PDIFF $count=1 $X=5.71
+ $Y=1.835 $X2=5.89 $Y2=2.76
r122 3 62 600 $w=1.7e-07 $l=7.89937e-07 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=2.365 $X2=4.99 $Y2=2.805
r123 3 60 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=2.365 $X2=4.53 $Y2=2.565
r124 2 21 300 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=2 $X=2.27
+ $Y=2.365 $X2=2.705 $Y2=2.51
r125 1 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.62
+ $Y=2.32 $X2=0.76 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%Q 1 2 9 13 14 15 16 23 33
r22 23 35 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=6.445 $Y=2.035
+ $X2=6.445 $Y2=2.015
r23 16 30 4.20486 $w=3.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.445 $Y=2.775
+ $X2=6.445 $Y2=2.91
r24 15 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.445 $Y=2.405
+ $X2=6.445 $Y2=2.775
r25 14 35 0.716383 $w=3.68e-07 $l=2.3e-08 $layer=LI1_cond $X=6.445 $Y=1.992
+ $X2=6.445 $Y2=2.015
r26 14 33 7.4687 $w=3.68e-07 $l=1.42e-07 $layer=LI1_cond $X=6.445 $Y=1.992
+ $X2=6.445 $Y2=1.85
r27 14 15 10.2163 $w=3.68e-07 $l=3.28e-07 $layer=LI1_cond $X=6.445 $Y=2.077
+ $X2=6.445 $Y2=2.405
r28 14 23 1.30818 $w=3.68e-07 $l=4.2e-08 $layer=LI1_cond $X=6.445 $Y=2.077
+ $X2=6.445 $Y2=2.035
r29 13 33 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.54 $Y=1.17 $X2=6.54
+ $Y2=1.85
r30 7 13 10.7251 $w=4.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.395 $Y=0.935
+ $X2=6.395 $Y2=1.17
r31 7 9 10.8156 $w=4.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.395 $Y=0.935
+ $X2=6.395 $Y2=0.51
r32 2 35 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=1.835 $X2=6.355 $Y2=2.015
r33 2 30 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=1.835 $X2=6.355 $Y2=2.91
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.18
+ $Y=0.365 $X2=6.32 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_1%VGND 1 2 3 4 17 21 25 29 32 33 34 36 44 57
+ 58 61 64 67
c88 36 0 7.96279e-20 $X=2.53 $Y=0
c89 21 0 3.02476e-20 $X=2.645 $Y=0.37
r90 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r91 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r92 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r93 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r94 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r95 55 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r96 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r97 52 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.47
+ $Y2=0
r98 52 54 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.595 $Y=0 $X2=5.52
+ $Y2=0
r99 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r100 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r101 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r102 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r103 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r104 45 64 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.67
+ $Y2=0
r105 45 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=3.12
+ $Y2=0
r106 44 67 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.345 $Y=0 $X2=4.47
+ $Y2=0
r107 44 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.345 $Y=0
+ $X2=4.08 $Y2=0
r108 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r109 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r110 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r111 40 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r112 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r113 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r114 37 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.88
+ $Y2=0
r115 37 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.2
+ $Y2=0
r116 36 64 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.67
+ $Y2=0
r117 36 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.16
+ $Y2=0
r118 34 51 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r119 34 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r120 32 54 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.775 $Y=0
+ $X2=5.52 $Y2=0
r121 32 33 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.775 $Y=0
+ $X2=5.882 $Y2=0
r122 31 57 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.99 $Y=0 $X2=6.48
+ $Y2=0
r123 31 33 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=5.99 $Y=0 $X2=5.882
+ $Y2=0
r124 27 33 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.882 $Y=0.085
+ $X2=5.882 $Y2=0
r125 27 29 22.7808 $w=2.13e-07 $l=4.25e-07 $layer=LI1_cond $X=5.882 $Y=0.085
+ $X2=5.882 $Y2=0.51
r126 23 67 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.47 $Y=0.085
+ $X2=4.47 $Y2=0
r127 23 25 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=4.47 $Y=0.085
+ $X2=4.47 $Y2=0.39
r128 19 64 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=0.085
+ $X2=2.67 $Y2=0
r129 19 21 11.7302 $w=2.78e-07 $l=2.85e-07 $layer=LI1_cond $X=2.67 $Y=0.085
+ $X2=2.67 $Y2=0.37
r130 15 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.88 $Y=0.085
+ $X2=0.88 $Y2=0
r131 15 17 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.88 $Y=0.085
+ $X2=0.88 $Y2=0.54
r132 4 29 91 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=2 $X=5.64
+ $Y=0.365 $X2=5.89 $Y2=0.51
r133 3 25 182 $w=1.7e-07 $l=3.02738e-07 $layer=licon1_NDIFF $count=1 $X=4.195
+ $Y=0.235 $X2=4.43 $Y2=0.39
r134 2 21 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=2.505
+ $Y=0.235 $X2=2.645 $Y2=0.37
r135 1 17 182 $w=1.7e-07 $l=3.00333e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.35 $X2=0.88 $Y2=0.54
.ends

