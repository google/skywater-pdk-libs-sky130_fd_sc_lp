* NGSPICE file created from sky130_fd_sc_lp__inputiso0p_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__inputiso0p_lp A SLEEP VGND VNB VPB VPWR X
M1000 a_432_489# A a_342_489# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.26e+11p ps=1.44e+06u
M1001 a_342_489# A a_340_93# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1002 VPWR SLEEP a_112_489# VPB phighvt w=420000u l=150000u
+  ad=4.83e+11p pd=4.6e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_602_93# a_342_489# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.759e+11p ps=3.47e+06u
M1004 X a_342_489# a_602_93# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 a_112_489# SLEEP a_27_93# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1006 VGND SLEEP a_112_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 a_340_93# a_27_93# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_602_367# a_342_489# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1009 X a_342_489# a_602_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1010 VPWR A a_432_489# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_270_489# a_27_93# VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1012 a_112_93# SLEEP a_27_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1013 a_342_489# a_27_93# a_270_489# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

