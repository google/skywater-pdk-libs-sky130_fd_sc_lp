* File: sky130_fd_sc_lp__o311ai_2.pxi.spice
* Created: Fri Aug 28 11:14:35 2020
* 
x_PM_SKY130_FD_SC_LP__O311AI_2%A1 N_A1_c_87_n N_A1_M1018_g N_A1_M1004_g
+ N_A1_c_89_n N_A1_M1019_g N_A1_M1012_g A1 A1 N_A1_c_92_n
+ PM_SKY130_FD_SC_LP__O311AI_2%A1
x_PM_SKY130_FD_SC_LP__O311AI_2%A2 N_A2_c_128_n N_A2_M1006_g N_A2_M1003_g
+ N_A2_c_130_n N_A2_M1017_g N_A2_M1015_g A2 A2 N_A2_c_133_n
+ PM_SKY130_FD_SC_LP__O311AI_2%A2
x_PM_SKY130_FD_SC_LP__O311AI_2%A3 N_A3_M1002_g N_A3_c_185_n N_A3_M1005_g
+ N_A3_M1014_g N_A3_c_186_n N_A3_M1016_g A3 A3 A3 N_A3_c_183_n N_A3_c_184_n A3
+ PM_SKY130_FD_SC_LP__O311AI_2%A3
x_PM_SKY130_FD_SC_LP__O311AI_2%B1 N_B1_c_233_n N_B1_M1000_g N_B1_c_237_n
+ N_B1_M1007_g N_B1_c_234_n N_B1_M1009_g N_B1_c_238_n N_B1_M1013_g B1 B1
+ N_B1_c_236_n PM_SKY130_FD_SC_LP__O311AI_2%B1
x_PM_SKY130_FD_SC_LP__O311AI_2%C1 N_C1_c_282_n N_C1_M1008_g N_C1_M1001_g
+ N_C1_c_284_n N_C1_M1011_g N_C1_M1010_g C1 N_C1_c_287_n
+ PM_SKY130_FD_SC_LP__O311AI_2%C1
x_PM_SKY130_FD_SC_LP__O311AI_2%A_35_367# N_A_35_367#_M1004_s N_A_35_367#_M1012_s
+ N_A_35_367#_M1015_s N_A_35_367#_c_330_n N_A_35_367#_c_326_n
+ N_A_35_367#_c_327_n N_A_35_367#_c_333_n N_A_35_367#_c_328_n
+ N_A_35_367#_c_335_n N_A_35_367#_c_329_n PM_SKY130_FD_SC_LP__O311AI_2%A_35_367#
x_PM_SKY130_FD_SC_LP__O311AI_2%VPWR N_VPWR_M1004_d N_VPWR_M1007_s N_VPWR_M1001_d
+ N_VPWR_c_374_n N_VPWR_c_375_n N_VPWR_c_376_n VPWR N_VPWR_c_377_n
+ N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_373_n N_VPWR_c_382_n
+ N_VPWR_c_383_n N_VPWR_c_384_n PM_SKY130_FD_SC_LP__O311AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O311AI_2%A_290_367# N_A_290_367#_M1003_d
+ N_A_290_367#_M1005_d N_A_290_367#_c_448_n N_A_290_367#_c_447_n
+ N_A_290_367#_c_451_n N_A_290_367#_c_455_n
+ PM_SKY130_FD_SC_LP__O311AI_2%A_290_367#
x_PM_SKY130_FD_SC_LP__O311AI_2%Y N_Y_M1008_s N_Y_M1011_s N_Y_M1005_s N_Y_M1016_s
+ N_Y_M1013_d N_Y_M1010_s N_Y_c_475_n N_Y_c_476_n N_Y_c_477_n N_Y_c_524_n
+ N_Y_c_490_n N_Y_c_528_n N_Y_c_501_n N_Y_c_471_n N_Y_c_472_n N_Y_c_478_n
+ N_Y_c_479_n N_Y_c_473_n N_Y_c_480_n Y Y PM_SKY130_FD_SC_LP__O311AI_2%Y
x_PM_SKY130_FD_SC_LP__O311AI_2%A_35_47# N_A_35_47#_M1018_s N_A_35_47#_M1019_s
+ N_A_35_47#_M1017_s N_A_35_47#_M1014_d N_A_35_47#_M1009_d N_A_35_47#_c_552_n
+ N_A_35_47#_c_553_n N_A_35_47#_c_557_n N_A_35_47#_c_592_p N_A_35_47#_c_561_n
+ N_A_35_47#_c_594_p N_A_35_47#_c_567_n N_A_35_47#_c_596_p N_A_35_47#_c_575_n
+ N_A_35_47#_c_565_n N_A_35_47#_c_572_n N_A_35_47#_c_573_n N_A_35_47#_c_554_n
+ PM_SKY130_FD_SC_LP__O311AI_2%A_35_47#
x_PM_SKY130_FD_SC_LP__O311AI_2%VGND N_VGND_M1018_d N_VGND_M1006_d N_VGND_M1002_s
+ N_VGND_c_615_n N_VGND_c_616_n N_VGND_c_617_n N_VGND_c_618_n VGND
+ N_VGND_c_619_n N_VGND_c_620_n N_VGND_c_621_n N_VGND_c_622_n N_VGND_c_623_n
+ PM_SKY130_FD_SC_LP__O311AI_2%VGND
x_PM_SKY130_FD_SC_LP__O311AI_2%A_710_47# N_A_710_47#_M1000_s N_A_710_47#_M1008_d
+ N_A_710_47#_c_683_n N_A_710_47#_c_689_n N_A_710_47#_c_685_n
+ PM_SKY130_FD_SC_LP__O311AI_2%A_710_47#
cc_1 VNB N_A1_c_87_n 0.0218823f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.185
cc_2 VNB N_A1_M1004_g 0.0100771f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.465
cc_3 VNB N_A1_c_89_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.185
cc_4 VNB N_A1_M1012_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.465
cc_5 VNB A1 0.0123156f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_A1_c_92_n 0.0557969f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.35
cc_7 VNB N_A2_c_128_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.185
cc_8 VNB N_A2_M1003_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.465
cc_9 VNB N_A2_c_130_n 0.0166069f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.185
cc_10 VNB N_A2_M1015_g 0.00767737f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.465
cc_11 VNB A2 0.00522773f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_A2_c_133_n 0.041537f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.35
cc_13 VNB N_A3_M1002_g 0.0237794f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.655
cc_14 VNB N_A3_M1014_g 0.0233235f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.655
cc_15 VNB A3 0.00650328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A3_c_183_n 0.0830025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_c_184_n 0.00738118f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.31
cc_18 VNB N_B1_c_233_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.185
cc_19 VNB N_B1_c_234_n 0.0199724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B1 0.00140291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_c_236_n 0.0896213f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.35
cc_22 VNB N_C1_c_282_n 0.0181493f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.185
cc_23 VNB N_C1_M1001_g 0.00123444f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.465
cc_24 VNB N_C1_c_284_n 0.0215832f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.185
cc_25 VNB N_C1_M1010_g 0.002325f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.465
cc_26 VNB C1 0.0164775f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_C1_c_287_n 0.0661667f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.35
cc_28 VNB N_A_35_367#_c_326_n 0.00318647f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_29 VNB N_A_35_367#_c_327_n 0.00439283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_35_367#_c_328_n 0.00732277f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.35
cc_31 VNB N_A_35_367#_c_329_n 0.00204018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_373_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_471_n 0.00751114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_472_n 0.0225638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_473_n 0.00485114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB Y 0.00446394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_35_47#_c_552_n 0.00767415f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_38 VNB N_A_35_47#_c_553_n 0.0224525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_35_47#_c_554_n 0.00416984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_615_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.465
cc_41 VNB N_VGND_c_616_n 3.16049e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_42 VNB N_VGND_c_617_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.35
cc_43 VNB N_VGND_c_618_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_619_n 0.0166487f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.35
cc_45 VNB N_VGND_c_620_n 0.0262476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_621_n 0.0685887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_622_n 0.29947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_623_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_710_47#_c_683_n 0.0145533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_A1_M1004_g 0.0232847f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.465
cc_51 VPB N_A1_M1012_g 0.018727f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_52 VPB N_A2_M1003_g 0.0189261f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.465
cc_53 VPB N_A2_M1015_g 0.0234838f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_54 VPB N_A3_c_185_n 0.0195571f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.465
cc_55 VPB N_A3_c_186_n 0.0153124f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_56 VPB N_A3_c_183_n 0.0103059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_B1_c_237_n 0.0174674f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.515
cc_58 VPB N_B1_c_238_n 0.0174674f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=0.655
cc_59 VPB N_B1_c_236_n 0.0252315f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.35
cc_60 VPB N_C1_M1001_g 0.0181089f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.465
cc_61 VPB N_C1_M1010_g 0.0248098f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_62 VPB N_A_35_367#_c_330_n 0.0498589f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_63 VPB N_A_35_367#_c_326_n 0.00559032f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_64 VPB N_A_35_367#_c_327_n 0.0054421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_35_367#_c_333_n 9.96097e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_35_367#_c_328_n 0.0073007f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=1.35
cc_67 VPB N_A_35_367#_c_335_n 0.00953236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_374_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_69 VPB N_VPWR_c_375_n 0.00205393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_376_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.945 $Y2=1.35
cc_71 VPB N_VPWR_c_377_n 0.0166359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_378_n 0.0658478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_379_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_380_n 0.0153759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_373_n 0.0492184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_382_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_383_n 0.0112045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_384_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_290_367#_c_447_n 0.0108768f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=2.465
cc_80 VPB N_Y_c_475_n 0.00805648f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.35
cc_81 VPB N_Y_c_476_n 0.0017678f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.35
cc_82 VPB N_Y_c_477_n 0.0034708f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=1.35
cc_83 VPB N_Y_c_478_n 0.0450352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_Y_c_479_n 0.00364055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_Y_c_480_n 0.0106959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB Y 6.40348e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 N_A1_c_89_n N_A2_c_128_n 0.0162674f $X=0.945 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_88 N_A1_M1012_g N_A2_M1003_g 0.0260572f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_89 A1 A2 0.0221081f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 N_A1_c_92_n A2 0.0019391f $X=0.945 $Y=1.35 $X2=0 $Y2=0
cc_91 A1 N_A2_c_133_n 2.15703e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_92 N_A1_c_92_n N_A2_c_133_n 0.0231498f $X=0.945 $Y=1.35 $X2=0 $Y2=0
cc_93 N_A1_M1004_g N_A_35_367#_c_330_n 0.0046421f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A1_M1004_g N_A_35_367#_c_326_n 0.0157274f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A1_M1012_g N_A_35_367#_c_326_n 0.0152957f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_96 A1 N_A_35_367#_c_326_n 0.0395983f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A1_c_92_n N_A_35_367#_c_326_n 0.00357126f $X=0.945 $Y=1.35 $X2=0 $Y2=0
cc_98 A1 N_A_35_367#_c_327_n 0.0203393f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A1_c_92_n N_A_35_367#_c_327_n 0.00308111f $X=0.945 $Y=1.35 $X2=0 $Y2=0
cc_100 N_A1_M1012_g N_A_35_367#_c_333_n 0.0014373f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A1_M1004_g N_VPWR_c_374_n 0.0194824f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A1_M1012_g N_VPWR_c_374_n 0.0186126f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A1_M1004_g N_VPWR_c_377_n 0.00486043f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A1_M1012_g N_VPWR_c_378_n 0.00486043f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A1_M1004_g N_VPWR_c_373_n 0.00921558f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A1_M1012_g N_VPWR_c_373_n 0.0082726f $X=0.945 $Y=2.465 $X2=0 $Y2=0
cc_107 A1 N_A_35_47#_c_552_n 0.0194145f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_108 N_A1_c_92_n N_A_35_47#_c_552_n 0.00275891f $X=0.945 $Y=1.35 $X2=0 $Y2=0
cc_109 N_A1_c_87_n N_A_35_47#_c_557_n 0.00974987f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_110 N_A1_c_89_n N_A_35_47#_c_557_n 0.010739f $X=0.945 $Y=1.185 $X2=0 $Y2=0
cc_111 A1 N_A_35_47#_c_557_n 0.0333975f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_112 N_A1_c_92_n N_A_35_47#_c_557_n 0.00224206f $X=0.945 $Y=1.35 $X2=0 $Y2=0
cc_113 N_A1_c_87_n N_VGND_c_615_n 0.0116902f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_114 N_A1_c_89_n N_VGND_c_615_n 0.0100168f $X=0.945 $Y=1.185 $X2=0 $Y2=0
cc_115 N_A1_c_89_n N_VGND_c_616_n 5.68743e-19 $X=0.945 $Y=1.185 $X2=0 $Y2=0
cc_116 N_A1_c_89_n N_VGND_c_617_n 0.00486043f $X=0.945 $Y=1.185 $X2=0 $Y2=0
cc_117 N_A1_c_87_n N_VGND_c_619_n 0.00486043f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_118 N_A1_c_87_n N_VGND_c_622_n 0.00551988f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_119 N_A1_c_89_n N_VGND_c_622_n 0.0045769f $X=0.945 $Y=1.185 $X2=0 $Y2=0
cc_120 N_A2_c_130_n N_A3_M1002_g 0.0140194f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_121 A2 N_A3_M1002_g 2.5054e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A2_c_133_n N_A3_M1002_g 0.0147373f $X=1.805 $Y=1.35 $X2=0 $Y2=0
cc_123 N_A2_M1015_g N_A3_c_183_n 0.00452632f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_124 A2 N_A3_c_184_n 0.0221103f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A2_c_133_n N_A3_c_184_n 0.00144554f $X=1.805 $Y=1.35 $X2=0 $Y2=0
cc_126 N_A2_M1003_g N_A_35_367#_c_333_n 0.0014373f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A2_M1003_g N_A_35_367#_c_328_n 0.0142932f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A2_M1015_g N_A_35_367#_c_328_n 0.0157274f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_129 A2 N_A_35_367#_c_328_n 0.0463087f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A2_c_133_n N_A_35_367#_c_328_n 0.00406421f $X=1.805 $Y=1.35 $X2=0 $Y2=0
cc_131 N_A2_M1015_g N_A_35_367#_c_335_n 0.00561046f $X=1.805 $Y=2.465 $X2=0
+ $Y2=0
cc_132 A2 N_A_35_367#_c_329_n 0.012044f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_133 N_A2_c_133_n N_A_35_367#_c_329_n 6.41898e-19 $X=1.805 $Y=1.35 $X2=0 $Y2=0
cc_134 N_A2_M1003_g N_VPWR_c_374_n 0.00141193f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A2_M1003_g N_VPWR_c_378_n 0.00547432f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A2_M1015_g N_VPWR_c_378_n 0.00357842f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A2_M1003_g N_VPWR_c_373_n 0.00990114f $X=1.375 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A2_M1015_g N_VPWR_c_373_n 0.00675085f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A2_M1003_g N_A_290_367#_c_448_n 0.0111073f $X=1.375 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A2_M1015_g N_A_290_367#_c_448_n 0.0171569f $X=1.805 $Y=2.465 $X2=0
+ $Y2=0
cc_141 N_A2_M1015_g N_A_290_367#_c_447_n 0.0125611f $X=1.805 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A2_M1003_g N_A_290_367#_c_451_n 0.00192258f $X=1.375 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A2_M1015_g N_A_290_367#_c_451_n 5.81207e-19 $X=1.805 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A2_M1015_g N_Y_c_477_n 5.12182e-19 $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A2_c_128_n N_A_35_47#_c_561_n 0.00974987f $X=1.375 $Y=1.185 $X2=0 $Y2=0
cc_146 N_A2_c_130_n N_A_35_47#_c_561_n 0.00974987f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_147 A2 N_A_35_47#_c_561_n 0.0393215f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A2_c_133_n N_A_35_47#_c_561_n 0.00224206f $X=1.805 $Y=1.35 $X2=0 $Y2=0
cc_149 A2 N_A_35_47#_c_565_n 0.0112582f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_150 N_A2_c_133_n N_A_35_47#_c_565_n 5.45826e-19 $X=1.805 $Y=1.35 $X2=0 $Y2=0
cc_151 N_A2_c_128_n N_VGND_c_615_n 5.68743e-19 $X=1.375 $Y=1.185 $X2=0 $Y2=0
cc_152 N_A2_c_128_n N_VGND_c_616_n 0.0100168f $X=1.375 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A2_c_130_n N_VGND_c_616_n 0.0101389f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_154 N_A2_c_128_n N_VGND_c_617_n 0.00486043f $X=1.375 $Y=1.185 $X2=0 $Y2=0
cc_155 N_A2_c_130_n N_VGND_c_620_n 0.00542663f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_156 N_A2_c_128_n N_VGND_c_622_n 0.0045769f $X=1.375 $Y=1.185 $X2=0 $Y2=0
cc_157 N_A2_c_130_n N_VGND_c_622_n 0.0046706f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_158 N_A3_M1014_g N_B1_c_233_n 0.0115767f $X=3.045 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A3_c_186_n N_B1_c_237_n 0.016684f $X=3.185 $Y=1.725 $X2=0 $Y2=0
cc_160 A3 B1 0.0209428f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_161 A3 N_B1_c_236_n 0.00241743f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_162 N_A3_c_183_n N_B1_c_236_n 0.0325869f $X=3.045 $Y=1.5 $X2=0 $Y2=0
cc_163 N_A3_c_183_n N_A_35_367#_c_328_n 0.00336688f $X=3.045 $Y=1.5 $X2=0 $Y2=0
cc_164 N_A3_c_184_n N_A_35_367#_c_328_n 0.0100227f $X=2.68 $Y=1.355 $X2=0 $Y2=0
cc_165 N_A3_c_185_n N_A_35_367#_c_335_n 2.69622e-19 $X=2.755 $Y=1.725 $X2=0
+ $Y2=0
cc_166 N_A3_c_186_n N_VPWR_c_375_n 0.00144469f $X=3.185 $Y=1.725 $X2=0 $Y2=0
cc_167 N_A3_c_185_n N_VPWR_c_378_n 0.00357842f $X=2.755 $Y=1.725 $X2=0 $Y2=0
cc_168 N_A3_c_186_n N_VPWR_c_378_n 0.00547432f $X=3.185 $Y=1.725 $X2=0 $Y2=0
cc_169 N_A3_c_185_n N_VPWR_c_373_n 0.00675085f $X=2.755 $Y=1.725 $X2=0 $Y2=0
cc_170 N_A3_c_186_n N_VPWR_c_373_n 0.00990114f $X=3.185 $Y=1.725 $X2=0 $Y2=0
cc_171 N_A3_c_185_n N_A_290_367#_c_447_n 0.0131508f $X=2.755 $Y=1.725 $X2=0
+ $Y2=0
cc_172 N_A3_c_186_n N_A_290_367#_c_447_n 0.00193114f $X=3.185 $Y=1.725 $X2=0
+ $Y2=0
cc_173 N_A3_c_185_n N_A_290_367#_c_455_n 0.0152352f $X=2.755 $Y=1.725 $X2=0
+ $Y2=0
cc_174 N_A3_c_186_n N_A_290_367#_c_455_n 0.00923485f $X=3.185 $Y=1.725 $X2=0
+ $Y2=0
cc_175 N_A3_c_183_n N_A_290_367#_c_455_n 5.58532e-19 $X=3.045 $Y=1.5 $X2=0 $Y2=0
cc_176 N_A3_c_185_n N_Y_c_476_n 0.0116329f $X=2.755 $Y=1.725 $X2=0 $Y2=0
cc_177 N_A3_c_186_n N_Y_c_476_n 0.010711f $X=3.185 $Y=1.725 $X2=0 $Y2=0
cc_178 A3 N_Y_c_476_n 0.0378926f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A3_c_183_n N_Y_c_476_n 0.0140789f $X=3.045 $Y=1.5 $X2=0 $Y2=0
cc_180 N_A3_c_184_n N_Y_c_476_n 0.00336833f $X=2.68 $Y=1.355 $X2=0 $Y2=0
cc_181 N_A3_c_183_n N_Y_c_477_n 0.00695035f $X=3.045 $Y=1.5 $X2=0 $Y2=0
cc_182 N_A3_c_184_n N_Y_c_477_n 0.0220761f $X=2.68 $Y=1.355 $X2=0 $Y2=0
cc_183 N_A3_M1002_g N_A_35_47#_c_567_n 0.0111176f $X=2.275 $Y=0.655 $X2=0 $Y2=0
cc_184 N_A3_M1014_g N_A_35_47#_c_567_n 0.011071f $X=3.045 $Y=0.655 $X2=0 $Y2=0
cc_185 A3 N_A_35_47#_c_567_n 0.0333436f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A3_c_183_n N_A_35_47#_c_567_n 0.0024569f $X=3.045 $Y=1.5 $X2=0 $Y2=0
cc_187 N_A3_c_184_n N_A_35_47#_c_567_n 0.0361529f $X=2.68 $Y=1.355 $X2=0 $Y2=0
cc_188 N_A3_c_184_n N_A_35_47#_c_572_n 0.00671683f $X=2.68 $Y=1.355 $X2=0 $Y2=0
cc_189 A3 N_A_35_47#_c_573_n 0.00272663f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A3_c_183_n N_A_35_47#_c_573_n 0.00181406f $X=3.045 $Y=1.5 $X2=0 $Y2=0
cc_191 N_A3_M1002_g N_VGND_c_616_n 5.51564e-19 $X=2.275 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A3_M1002_g N_VGND_c_620_n 0.0170615f $X=2.275 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A3_M1014_g N_VGND_c_620_n 0.0136347f $X=3.045 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A3_M1014_g N_VGND_c_621_n 0.00468308f $X=3.045 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A3_M1002_g N_VGND_c_622_n 0.00467065f $X=2.275 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A3_M1014_g N_VGND_c_622_n 0.00441586f $X=3.045 $Y=0.655 $X2=0 $Y2=0
cc_197 B1 N_C1_c_282_n 2.16322e-19 $X=3.995 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_198 N_B1_c_236_n N_C1_c_282_n 0.00384505f $X=3.975 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_199 N_B1_c_238_n N_C1_M1001_g 0.0169079f $X=4.425 $Y=1.725 $X2=0 $Y2=0
cc_200 N_B1_c_236_n N_C1_c_287_n 0.0169079f $X=3.975 $Y=1.35 $X2=0 $Y2=0
cc_201 N_B1_c_237_n N_VPWR_c_375_n 0.0182013f $X=3.615 $Y=1.725 $X2=0 $Y2=0
cc_202 N_B1_c_238_n N_VPWR_c_375_n 0.0169909f $X=4.425 $Y=1.725 $X2=0 $Y2=0
cc_203 N_B1_c_236_n N_VPWR_c_375_n 0.00268755f $X=3.975 $Y=1.35 $X2=0 $Y2=0
cc_204 N_B1_c_238_n N_VPWR_c_376_n 7.38487e-19 $X=4.425 $Y=1.725 $X2=0 $Y2=0
cc_205 N_B1_c_237_n N_VPWR_c_378_n 0.00486043f $X=3.615 $Y=1.725 $X2=0 $Y2=0
cc_206 N_B1_c_238_n N_VPWR_c_379_n 0.00486043f $X=4.425 $Y=1.725 $X2=0 $Y2=0
cc_207 N_B1_c_237_n N_VPWR_c_373_n 0.0082726f $X=3.615 $Y=1.725 $X2=0 $Y2=0
cc_208 N_B1_c_238_n N_VPWR_c_373_n 0.0082726f $X=4.425 $Y=1.725 $X2=0 $Y2=0
cc_209 N_B1_c_237_n N_Y_c_490_n 0.0119166f $X=3.615 $Y=1.725 $X2=0 $Y2=0
cc_210 N_B1_c_238_n N_Y_c_490_n 0.00807119f $X=4.425 $Y=1.725 $X2=0 $Y2=0
cc_211 B1 N_Y_c_490_n 0.053856f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_212 N_B1_c_236_n N_Y_c_490_n 0.0296281f $X=3.975 $Y=1.35 $X2=0 $Y2=0
cc_213 B1 N_Y_c_479_n 0.00190569f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_214 N_B1_c_236_n N_Y_c_479_n 0.0041154f $X=3.975 $Y=1.35 $X2=0 $Y2=0
cc_215 N_B1_c_234_n N_Y_c_473_n 7.59783e-19 $X=3.905 $Y=1.185 $X2=0 $Y2=0
cc_216 N_B1_c_234_n Y 0.00424849f $X=3.905 $Y=1.185 $X2=0 $Y2=0
cc_217 N_B1_c_238_n Y 0.00413046f $X=4.425 $Y=1.725 $X2=0 $Y2=0
cc_218 B1 Y 0.0283326f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_219 N_B1_c_236_n Y 0.0207017f $X=3.975 $Y=1.35 $X2=0 $Y2=0
cc_220 N_B1_c_233_n N_A_35_47#_c_575_n 0.0115355f $X=3.475 $Y=1.185 $X2=0 $Y2=0
cc_221 N_B1_c_234_n N_A_35_47#_c_575_n 0.01039f $X=3.905 $Y=1.185 $X2=0 $Y2=0
cc_222 B1 N_A_35_47#_c_575_n 0.0346481f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_223 N_B1_c_236_n N_A_35_47#_c_575_n 0.00263605f $X=3.975 $Y=1.35 $X2=0 $Y2=0
cc_224 B1 N_A_35_47#_c_554_n 0.0201095f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_225 N_B1_c_236_n N_A_35_47#_c_554_n 0.0065477f $X=3.975 $Y=1.35 $X2=0 $Y2=0
cc_226 N_B1_c_233_n N_VGND_c_620_n 0.00128107f $X=3.475 $Y=1.185 $X2=0 $Y2=0
cc_227 N_B1_c_233_n N_VGND_c_621_n 0.0054895f $X=3.475 $Y=1.185 $X2=0 $Y2=0
cc_228 N_B1_c_234_n N_VGND_c_621_n 0.00359361f $X=3.905 $Y=1.185 $X2=0 $Y2=0
cc_229 N_B1_c_233_n N_VGND_c_622_n 0.00631323f $X=3.475 $Y=1.185 $X2=0 $Y2=0
cc_230 N_B1_c_234_n N_VGND_c_622_n 0.00681249f $X=3.905 $Y=1.185 $X2=0 $Y2=0
cc_231 N_B1_c_234_n N_A_710_47#_c_683_n 0.0108881f $X=3.905 $Y=1.185 $X2=0 $Y2=0
cc_232 N_B1_c_233_n N_A_710_47#_c_685_n 0.00596801f $X=3.475 $Y=1.185 $X2=0
+ $Y2=0
cc_233 N_B1_c_234_n N_A_710_47#_c_685_n 0.010895f $X=3.905 $Y=1.185 $X2=0 $Y2=0
cc_234 N_C1_M1001_g N_VPWR_c_375_n 7.56945e-19 $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_235 N_C1_M1001_g N_VPWR_c_376_n 0.0149832f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_236 N_C1_M1010_g N_VPWR_c_376_n 0.0169864f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_237 N_C1_c_287_n N_VPWR_c_376_n 4.4534e-19 $X=5.47 $Y=1.46 $X2=0 $Y2=0
cc_238 N_C1_M1001_g N_VPWR_c_379_n 0.00486043f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_239 N_C1_M1010_g N_VPWR_c_380_n 0.00486043f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_240 N_C1_M1001_g N_VPWR_c_373_n 0.0082726f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_241 N_C1_M1010_g N_VPWR_c_373_n 0.00917987f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_242 N_C1_c_284_n N_Y_c_501_n 0.0136479f $X=5.285 $Y=1.295 $X2=0 $Y2=0
cc_243 C1 N_Y_c_501_n 0.00603379f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_244 C1 N_Y_c_471_n 0.0226827f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_245 N_C1_c_287_n N_Y_c_471_n 0.0014684f $X=5.47 $Y=1.46 $X2=0 $Y2=0
cc_246 N_C1_c_284_n N_Y_c_472_n 0.00149752f $X=5.285 $Y=1.295 $X2=0 $Y2=0
cc_247 N_C1_c_282_n N_Y_c_473_n 0.0120487f $X=4.855 $Y=1.295 $X2=0 $Y2=0
cc_248 N_C1_c_284_n N_Y_c_473_n 4.48476e-19 $X=5.285 $Y=1.295 $X2=0 $Y2=0
cc_249 N_C1_M1010_g N_Y_c_480_n 0.0159383f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_250 C1 N_Y_c_480_n 0.0301425f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_251 N_C1_c_287_n N_Y_c_480_n 0.00700691f $X=5.47 $Y=1.46 $X2=0 $Y2=0
cc_252 N_C1_c_282_n Y 0.00720244f $X=4.855 $Y=1.295 $X2=0 $Y2=0
cc_253 N_C1_M1001_g Y 0.0156639f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_254 N_C1_c_284_n Y 0.00571285f $X=5.285 $Y=1.295 $X2=0 $Y2=0
cc_255 N_C1_M1010_g Y 0.00268115f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_256 C1 Y 0.0271948f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_257 N_C1_c_287_n Y 0.0264077f $X=5.47 $Y=1.46 $X2=0 $Y2=0
cc_258 N_C1_c_282_n N_VGND_c_621_n 0.0029147f $X=4.855 $Y=1.295 $X2=0 $Y2=0
cc_259 N_C1_c_284_n N_VGND_c_621_n 0.00463152f $X=5.285 $Y=1.295 $X2=0 $Y2=0
cc_260 N_C1_c_282_n N_VGND_c_622_n 0.00428625f $X=4.855 $Y=1.295 $X2=0 $Y2=0
cc_261 N_C1_c_284_n N_VGND_c_622_n 0.00920454f $X=5.285 $Y=1.295 $X2=0 $Y2=0
cc_262 N_C1_c_282_n N_A_710_47#_c_683_n 0.0115438f $X=4.855 $Y=1.295 $X2=0 $Y2=0
cc_263 N_C1_c_284_n N_A_710_47#_c_683_n 0.00575349f $X=5.285 $Y=1.295 $X2=0
+ $Y2=0
cc_264 N_C1_c_284_n N_A_710_47#_c_689_n 0.00291499f $X=5.285 $Y=1.295 $X2=0
+ $Y2=0
cc_265 N_C1_c_287_n N_A_710_47#_c_689_n 3.20405e-19 $X=5.47 $Y=1.46 $X2=0 $Y2=0
cc_266 N_A_35_367#_c_326_n N_VPWR_c_374_n 0.0216087f $X=1.065 $Y=1.69 $X2=0
+ $Y2=0
cc_267 N_A_35_367#_c_330_n N_VPWR_c_377_n 0.0178111f $X=0.3 $Y=1.98 $X2=0 $Y2=0
cc_268 N_A_35_367#_c_333_n N_VPWR_c_378_n 0.0124525f $X=1.16 $Y=1.98 $X2=0 $Y2=0
cc_269 N_A_35_367#_M1004_s N_VPWR_c_373_n 0.00371702f $X=0.175 $Y=1.835 $X2=0
+ $Y2=0
cc_270 N_A_35_367#_M1012_s N_VPWR_c_373_n 0.00536646f $X=1.02 $Y=1.835 $X2=0
+ $Y2=0
cc_271 N_A_35_367#_M1015_s N_VPWR_c_373_n 0.0021598f $X=1.88 $Y=1.835 $X2=0
+ $Y2=0
cc_272 N_A_35_367#_c_330_n N_VPWR_c_373_n 0.0100304f $X=0.3 $Y=1.98 $X2=0 $Y2=0
cc_273 N_A_35_367#_c_333_n N_VPWR_c_373_n 0.00730901f $X=1.16 $Y=1.98 $X2=0
+ $Y2=0
cc_274 N_A_35_367#_c_328_n N_A_290_367#_c_448_n 0.0216087f $X=1.925 $Y=1.69
+ $X2=0 $Y2=0
cc_275 N_A_35_367#_M1015_s N_A_290_367#_c_447_n 0.00495471f $X=1.88 $Y=1.835
+ $X2=0 $Y2=0
cc_276 N_A_35_367#_c_335_n N_A_290_367#_c_447_n 0.0189128f $X=2.02 $Y=1.98 $X2=0
+ $Y2=0
cc_277 N_A_35_367#_c_335_n N_Y_c_475_n 0.0645801f $X=2.02 $Y=1.98 $X2=0 $Y2=0
cc_278 N_A_35_367#_c_328_n N_Y_c_477_n 0.00692503f $X=1.925 $Y=1.69 $X2=0 $Y2=0
cc_279 N_A_35_367#_c_335_n N_Y_c_477_n 0.00719825f $X=2.02 $Y=1.98 $X2=0 $Y2=0
cc_280 N_A_35_367#_c_327_n N_A_35_47#_c_552_n 7.84729e-19 $X=0.395 $Y=1.69 $X2=0
+ $Y2=0
cc_281 N_A_35_367#_c_326_n N_A_35_47#_c_557_n 0.00250493f $X=1.065 $Y=1.69 $X2=0
+ $Y2=0
cc_282 N_A_35_367#_c_329_n N_A_35_47#_c_565_n 0.00165326f $X=1.16 $Y=1.69 $X2=0
+ $Y2=0
cc_283 N_A_35_367#_c_328_n N_A_35_47#_c_572_n 0.00519785f $X=1.925 $Y=1.69 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_373_n N_A_290_367#_M1003_d 0.00223559f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_285 N_VPWR_c_373_n N_A_290_367#_M1005_d 0.00223559f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_286 N_VPWR_c_378_n N_A_290_367#_c_447_n 0.0821667f $X=3.665 $Y=3.33 $X2=0
+ $Y2=0
cc_287 N_VPWR_c_373_n N_A_290_367#_c_447_n 0.0507876f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_288 N_VPWR_c_378_n N_A_290_367#_c_451_n 0.0189946f $X=3.665 $Y=3.33 $X2=0
+ $Y2=0
cc_289 N_VPWR_c_373_n N_A_290_367#_c_451_n 0.0124451f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_373_n N_Y_M1005_s 0.0021598f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_291 N_VPWR_c_373_n N_Y_M1016_s 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_292 N_VPWR_c_373_n N_Y_M1013_d 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_293 N_VPWR_c_373_n N_Y_M1010_s 0.00371702f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_294 N_VPWR_c_378_n N_Y_c_524_n 0.0124525f $X=3.665 $Y=3.33 $X2=0 $Y2=0
cc_295 N_VPWR_c_373_n N_Y_c_524_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_296 N_VPWR_M1007_s N_Y_c_490_n 0.00580409f $X=3.69 $Y=1.835 $X2=0 $Y2=0
cc_297 N_VPWR_c_375_n N_Y_c_490_n 0.0479937f $X=3.83 $Y=2.12 $X2=0 $Y2=0
cc_298 N_VPWR_c_379_n N_Y_c_528_n 0.0124525f $X=4.905 $Y=3.33 $X2=0 $Y2=0
cc_299 N_VPWR_c_373_n N_Y_c_528_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_300 N_VPWR_c_380_n N_Y_c_478_n 0.0178111f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_301 N_VPWR_c_373_n N_Y_c_478_n 0.0100304f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_302 N_VPWR_M1001_d N_Y_c_480_n 2.87015e-19 $X=4.93 $Y=1.835 $X2=0 $Y2=0
cc_303 N_VPWR_c_376_n N_Y_c_480_n 0.00402765f $X=5.07 $Y=2.14 $X2=0 $Y2=0
cc_304 N_VPWR_M1001_d Y 0.00152714f $X=4.93 $Y=1.835 $X2=0 $Y2=0
cc_305 N_VPWR_c_376_n Y 0.0144316f $X=5.07 $Y=2.14 $X2=0 $Y2=0
cc_306 N_A_290_367#_c_447_n N_Y_M1005_s 0.00495471f $X=2.805 $Y=2.99 $X2=0 $Y2=0
cc_307 N_A_290_367#_c_447_n N_Y_c_475_n 0.0189128f $X=2.805 $Y=2.99 $X2=0 $Y2=0
cc_308 N_A_290_367#_M1005_d N_Y_c_476_n 0.00176461f $X=2.83 $Y=1.835 $X2=0 $Y2=0
cc_309 N_A_290_367#_c_455_n N_Y_c_476_n 0.0170776f $X=2.97 $Y=2.12 $X2=0 $Y2=0
cc_310 N_Y_c_479_n N_A_35_47#_c_573_n 0.00148174f $X=3.4 $Y=1.78 $X2=0 $Y2=0
cc_311 N_Y_c_473_n N_A_35_47#_c_554_n 0.0353114f $X=4.79 $Y=1.04 $X2=0 $Y2=0
cc_312 N_Y_c_472_n N_VGND_c_621_n 0.0127568f $X=5.5 $Y=0.5 $X2=0 $Y2=0
cc_313 N_Y_c_472_n N_VGND_c_622_n 0.0099985f $X=5.5 $Y=0.5 $X2=0 $Y2=0
cc_314 N_Y_c_501_n N_A_710_47#_M1008_d 8.3052e-19 $X=5.395 $Y=0.955 $X2=0 $Y2=0
cc_315 N_Y_c_473_n N_A_710_47#_M1008_d 0.00152714f $X=4.79 $Y=1.04 $X2=0 $Y2=0
cc_316 Y N_A_710_47#_M1008_d 0.0018839f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_317 N_Y_M1008_s N_A_710_47#_c_683_n 0.00258276f $X=4.515 $Y=0.345 $X2=0 $Y2=0
cc_318 N_Y_c_472_n N_A_710_47#_c_683_n 0.00415594f $X=5.5 $Y=0.5 $X2=0 $Y2=0
cc_319 N_Y_c_473_n N_A_710_47#_c_683_n 0.0266567f $X=4.79 $Y=1.04 $X2=0 $Y2=0
cc_320 N_Y_c_501_n N_A_710_47#_c_689_n 0.00315508f $X=5.395 $Y=0.955 $X2=0 $Y2=0
cc_321 N_Y_c_473_n N_A_710_47#_c_689_n 0.0120631f $X=4.79 $Y=1.04 $X2=0 $Y2=0
cc_322 N_A_35_47#_c_557_n N_VGND_M1018_d 0.00328155f $X=1.065 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_323 N_A_35_47#_c_561_n N_VGND_M1006_d 0.00328155f $X=1.925 $Y=0.93 $X2=0
+ $Y2=0
cc_324 N_A_35_47#_c_567_n N_VGND_M1002_s 0.012232f $X=3.17 $Y=0.93 $X2=0 $Y2=0
cc_325 N_A_35_47#_c_557_n N_VGND_c_615_n 0.016709f $X=1.065 $Y=0.93 $X2=0 $Y2=0
cc_326 N_A_35_47#_c_561_n N_VGND_c_616_n 0.016709f $X=1.925 $Y=0.93 $X2=0 $Y2=0
cc_327 N_A_35_47#_c_592_p N_VGND_c_617_n 0.0124525f $X=1.16 $Y=0.42 $X2=0 $Y2=0
cc_328 N_A_35_47#_c_553_n N_VGND_c_619_n 0.0178111f $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_329 N_A_35_47#_c_594_p N_VGND_c_620_n 0.015265f $X=2.035 $Y=0.42 $X2=0 $Y2=0
cc_330 N_A_35_47#_c_567_n N_VGND_c_620_n 0.0441491f $X=3.17 $Y=0.93 $X2=0 $Y2=0
cc_331 N_A_35_47#_c_596_p N_VGND_c_621_n 0.0122751f $X=3.26 $Y=0.42 $X2=0 $Y2=0
cc_332 N_A_35_47#_M1018_s N_VGND_c_622_n 0.00243868f $X=0.175 $Y=0.235 $X2=0
+ $Y2=0
cc_333 N_A_35_47#_M1019_s N_VGND_c_622_n 0.00280978f $X=1.02 $Y=0.235 $X2=0
+ $Y2=0
cc_334 N_A_35_47#_M1017_s N_VGND_c_622_n 0.00313145f $X=1.88 $Y=0.235 $X2=0
+ $Y2=0
cc_335 N_A_35_47#_M1014_d N_VGND_c_622_n 0.00284332f $X=3.12 $Y=0.235 $X2=0
+ $Y2=0
cc_336 N_A_35_47#_M1009_d N_VGND_c_622_n 0.00215176f $X=3.98 $Y=0.235 $X2=0
+ $Y2=0
cc_337 N_A_35_47#_c_553_n N_VGND_c_622_n 0.0100304f $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_338 N_A_35_47#_c_557_n N_VGND_c_622_n 0.0108383f $X=1.065 $Y=0.93 $X2=0 $Y2=0
cc_339 N_A_35_47#_c_592_p N_VGND_c_622_n 0.00730901f $X=1.16 $Y=0.42 $X2=0 $Y2=0
cc_340 N_A_35_47#_c_561_n N_VGND_c_622_n 0.0108383f $X=1.925 $Y=0.93 $X2=0 $Y2=0
cc_341 N_A_35_47#_c_594_p N_VGND_c_622_n 0.00886411f $X=2.035 $Y=0.42 $X2=0
+ $Y2=0
cc_342 N_A_35_47#_c_567_n N_VGND_c_622_n 0.0119704f $X=3.17 $Y=0.93 $X2=0 $Y2=0
cc_343 N_A_35_47#_c_596_p N_VGND_c_622_n 0.00711462f $X=3.26 $Y=0.42 $X2=0 $Y2=0
cc_344 N_A_35_47#_c_575_n N_VGND_c_622_n 0.00582354f $X=4.025 $Y=0.93 $X2=0
+ $Y2=0
cc_345 N_A_35_47#_c_575_n N_A_710_47#_M1000_s 0.00328155f $X=4.025 $Y=0.93
+ $X2=-0.19 $Y2=-0.245
cc_346 N_A_35_47#_M1009_d N_A_710_47#_c_683_n 0.00495471f $X=3.98 $Y=0.235 $X2=0
+ $Y2=0
cc_347 N_A_35_47#_c_575_n N_A_710_47#_c_683_n 0.00347435f $X=4.025 $Y=0.93 $X2=0
+ $Y2=0
cc_348 N_A_35_47#_c_554_n N_A_710_47#_c_683_n 0.0182319f $X=4.12 $Y=0.76 $X2=0
+ $Y2=0
cc_349 N_A_35_47#_c_575_n N_A_710_47#_c_685_n 0.0160582f $X=4.025 $Y=0.93 $X2=0
+ $Y2=0
cc_350 N_VGND_c_622_n N_A_710_47#_M1000_s 0.00225167f $X=5.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_351 N_VGND_c_621_n N_A_710_47#_c_683_n 0.0867598f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_622_n N_A_710_47#_c_683_n 0.0504013f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_621_n N_A_710_47#_c_685_n 0.0184793f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_c_622_n N_A_710_47#_c_685_n 0.0123776f $X=5.52 $Y=0 $X2=0 $Y2=0
