* File: sky130_fd_sc_lp__nand3b_4.spice
* Created: Wed Sep  2 10:04:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand3b_4.pex.spice"
.subckt sky130_fd_sc_lp__nand3b_4  VNB VPB A_N B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_N_M1013_g N_A_35_74#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_225_47#_M1000_d N_A_35_74#_M1000_g N_Y_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1010 N_A_225_47#_M1010_d N_A_35_74#_M1010_g N_Y_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1014 N_A_225_47#_M1010_d N_A_35_74#_M1014_g N_Y_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1025 N_A_225_47#_M1025_d N_A_35_74#_M1025_g N_Y_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1007 N_A_225_47#_M1025_d N_B_M1007_g N_A_652_47#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1008 N_A_225_47#_M1008_d N_B_M1008_g N_A_652_47#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1022 N_A_225_47#_M1008_d N_B_M1022_g N_A_652_47#_M1022_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1024 N_A_225_47#_M1024_d N_B_M1024_g N_A_652_47#_M1022_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_A_652_47#_M1002_d N_C_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1004 N_A_652_47#_M1002_d N_C_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1015 N_A_652_47#_M1015_d N_C_M1015_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1019 N_A_652_47#_M1015_d N_C_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_A_N_M1016_g N_A_35_74#_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.21735 AS=0.3339 PD=1.605 PS=3.05 NRD=8.5892 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.7 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A_35_74#_M1001_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.21735 PD=1.54 PS=1.605 NRD=0 NRS=1.5563 M=1 R=8.4 SA=75000.7
+ SB=75005.2 A=0.189 P=2.82 MULT=1
MM1009 N_Y_M1001_d N_A_35_74#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.8 A=0.189 P=2.82 MULT=1
MM1017 N_Y_M1017_d N_A_35_74#_M1017_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75004.4 A=0.189 P=2.82 MULT=1
MM1023 N_Y_M1017_d N_A_35_74#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1953 PD=1.54 PS=1.57 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75003.9
+ A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1023_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1953 PD=1.54 PS=1.57 NRD=0 NRS=4.6886 M=1 R=8.4 SA=75002.4
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1003_d N_B_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2268 PD=1.54 PS=1.62 NRD=0 NRS=5.4569 M=1 R=8.4 SA=75002.9
+ SB=75003 A=0.189 P=2.82 MULT=1
MM1012 N_Y_M1012_d N_B_M1012_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2268 PD=1.54 PS=1.62 NRD=0 NRS=7.0329 M=1 R=8.4 SA=75003.4
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1021 N_Y_M1012_d N_B_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.29295 PD=1.54 PS=1.725 NRD=0 NRS=12.4898 M=1 R=8.4 SA=75003.8
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1021_s N_C_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.29295 AS=0.1764 PD=1.725 PS=1.54 NRD=16.4101 NRS=0 M=1 R=8.4 SA=75004.4
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_C_M1011_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.9
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1011_d N_C_M1018_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1020 N_VPWR_M1020_d N_C_M1020_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=14.1367 P=18.89
*
.include "sky130_fd_sc_lp__nand3b_4.pxi.spice"
*
.ends
*
*
