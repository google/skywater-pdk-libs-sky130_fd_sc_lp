* File: sky130_fd_sc_lp__or4_1.spice
* Created: Fri Aug 28 11:24:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4_1.pex.spice"
.subckt sky130_fd_sc_lp__or4_1  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1003 N_A_40_480#_M1003_d N_D_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_C_M1001_g N_A_40_480#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0588 PD=1.04 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_40_480#_M1000_d N_B_M1000_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.1302 PD=0.72 PS=1.04 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_40_480#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0847 AS=0.063 PD=0.786667 PS=0.72 NRD=17.136 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_40_480#_M1009_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1694 PD=2.21 PS=1.57333 NRD=0 NRS=0 M=1 R=5.6 SA=75001.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 A_123_480# N_D_M1006_g N_A_40_480#_M1006_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1004 A_195_480# N_C_M1004_g A_123_480# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1005 A_267_480# N_B_M1005_g A_195_480# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75000.9
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g A_267_480# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.172725 AS=0.0441 PD=1.1875 PS=0.63 NRD=167.095 NRS=23.443 M=1 R=2.8
+ SA=75001.3 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1007 N_X_M1007_d N_A_40_480#_M1007_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.518175 PD=3.05 PS=3.5625 NRD=0 NRS=0 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__or4_1.pxi.spice"
*
.ends
*
*
