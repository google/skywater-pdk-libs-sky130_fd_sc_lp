* File: sky130_fd_sc_lp__or4bb_m.pxi.spice
* Created: Wed Sep  2 10:33:34 2020
* 
x_PM_SKY130_FD_SC_LP__OR4BB_M%C_N N_C_N_M1011_g N_C_N_M1010_g N_C_N_c_99_n
+ N_C_N_c_100_n N_C_N_c_101_n C_N C_N N_C_N_c_103_n
+ PM_SKY130_FD_SC_LP__OR4BB_M%C_N
x_PM_SKY130_FD_SC_LP__OR4BB_M%D_N N_D_N_M1006_g N_D_N_M1001_g D_N N_D_N_c_134_n
+ N_D_N_c_135_n PM_SKY130_FD_SC_LP__OR4BB_M%D_N
x_PM_SKY130_FD_SC_LP__OR4BB_M%A_196_530# N_A_196_530#_M1001_d
+ N_A_196_530#_M1006_d N_A_196_530#_c_167_n N_A_196_530#_c_177_n
+ N_A_196_530#_c_168_n N_A_196_530#_M1002_g N_A_196_530#_c_178_n
+ N_A_196_530#_M1004_g N_A_196_530#_c_169_n N_A_196_530#_c_170_n
+ N_A_196_530#_c_179_n N_A_196_530#_c_180_n N_A_196_530#_c_181_n
+ N_A_196_530#_c_171_n N_A_196_530#_c_172_n N_A_196_530#_c_173_n
+ N_A_196_530#_c_174_n N_A_196_530#_c_175_n N_A_196_530#_c_182_n
+ PM_SKY130_FD_SC_LP__OR4BB_M%A_196_530#
x_PM_SKY130_FD_SC_LP__OR4BB_M%A_27_530# N_A_27_530#_M1010_s N_A_27_530#_M1011_s
+ N_A_27_530#_c_238_n N_A_27_530#_M1005_g N_A_27_530#_M1009_g
+ N_A_27_530#_c_240_n N_A_27_530#_c_247_n N_A_27_530#_c_241_n
+ N_A_27_530#_c_242_n N_A_27_530#_c_243_n N_A_27_530#_c_244_n
+ PM_SKY130_FD_SC_LP__OR4BB_M%A_27_530#
x_PM_SKY130_FD_SC_LP__OR4BB_M%B N_B_M1007_g N_B_M1013_g N_B_c_314_n N_B_c_315_n
+ B N_B_c_316_n N_B_c_317_n PM_SKY130_FD_SC_LP__OR4BB_M%B
x_PM_SKY130_FD_SC_LP__OR4BB_M%A N_A_M1008_g N_A_M1003_g A A N_A_c_361_n
+ N_A_c_362_n PM_SKY130_FD_SC_LP__OR4BB_M%A
x_PM_SKY130_FD_SC_LP__OR4BB_M%A_336_439# N_A_336_439#_M1002_d
+ N_A_336_439#_M1013_d N_A_336_439#_M1004_s N_A_336_439#_M1000_g
+ N_A_336_439#_M1012_g N_A_336_439#_c_407_n N_A_336_439#_c_408_n
+ N_A_336_439#_c_417_n N_A_336_439#_c_409_n N_A_336_439#_c_418_n
+ N_A_336_439#_c_419_n N_A_336_439#_c_420_n N_A_336_439#_c_410_n
+ N_A_336_439#_c_421_n N_A_336_439#_c_411_n N_A_336_439#_c_412_n
+ N_A_336_439#_c_413_n N_A_336_439#_c_414_n N_A_336_439#_c_422_n
+ PM_SKY130_FD_SC_LP__OR4BB_M%A_336_439#
x_PM_SKY130_FD_SC_LP__OR4BB_M%VPWR N_VPWR_M1011_d N_VPWR_M1008_d N_VPWR_c_514_n
+ N_VPWR_c_515_n VPWR N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n
+ N_VPWR_c_513_n N_VPWR_c_520_n N_VPWR_c_521_n PM_SKY130_FD_SC_LP__OR4BB_M%VPWR
x_PM_SKY130_FD_SC_LP__OR4BB_M%X N_X_M1012_d N_X_M1000_d N_X_c_560_n X X X
+ PM_SKY130_FD_SC_LP__OR4BB_M%X
x_PM_SKY130_FD_SC_LP__OR4BB_M%VGND N_VGND_M1010_d N_VGND_M1002_s N_VGND_M1009_d
+ N_VGND_M1003_d N_VGND_c_578_n N_VGND_c_579_n N_VGND_c_580_n N_VGND_c_581_n
+ N_VGND_c_582_n N_VGND_c_583_n VGND N_VGND_c_584_n N_VGND_c_585_n
+ N_VGND_c_586_n N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n
+ PM_SKY130_FD_SC_LP__OR4BB_M%VGND
cc_1 VNB N_C_N_M1011_g 0.012749f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.86
cc_2 VNB N_C_N_c_99_n 0.0197225f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.775
cc_3 VNB N_C_N_c_100_n 0.0236573f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.28
cc_4 VNB N_C_N_c_101_n 0.0166257f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.445
cc_5 VNB C_N 0.0114808f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_C_N_c_103_n 0.0165017f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.94
cc_7 VNB N_D_N_M1001_g 0.0690113f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.455
cc_8 VNB N_A_196_530#_c_167_n 0.0132189f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.94
cc_9 VNB N_A_196_530#_c_168_n 0.020721f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_A_196_530#_c_169_n 0.0404689f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.94
cc_11 VNB N_A_196_530#_c_170_n 0.0175896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_196_530#_c_171_n 0.00195177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_196_530#_c_172_n 0.0092036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_196_530#_c_173_n 0.0105415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_196_530#_c_174_n 7.34898e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_196_530#_c_175_n 0.0303107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_530#_c_238_n 0.029944f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.455
cc_18 VNB N_A_27_530#_M1009_g 0.05067f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_19 VNB N_A_27_530#_c_240_n 0.0484712f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.94
cc_20 VNB N_A_27_530#_c_241_n 0.0329163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_530#_c_242_n 0.015658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_530#_c_243_n 0.0050149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_530#_c_244_n 0.00186192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_M1007_g 0.00512236f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.86
cc_25 VNB N_B_M1013_g 0.0231207f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.455
cc_26 VNB N_B_c_314_n 0.0193493f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.445
cc_27 VNB N_B_c_315_n 0.0150351f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_28 VNB N_B_c_316_n 0.0150011f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.94
cc_29 VNB N_B_c_317_n 0.0143579f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.94
cc_30 VNB N_A_M1003_g 0.0579184f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.455
cc_31 VNB N_A_336_439#_M1012_g 0.0356906f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.94
cc_32 VNB N_A_336_439#_c_407_n 0.0253576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_336_439#_c_408_n 0.0093778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_336_439#_c_409_n 0.00617348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_336_439#_c_410_n 0.00656093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_336_439#_c_411_n 0.00187503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_336_439#_c_412_n 0.0187513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_336_439#_c_413_n 0.00570334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_336_439#_c_414_n 0.00699662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_513_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_560_n 0.0168419f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.775
cc_42 VNB X 0.046742f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_43 VNB N_VGND_c_578_n 0.00527464f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.94
cc_44 VNB N_VGND_c_579_n 0.0207374f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.925
cc_45 VNB N_VGND_c_580_n 0.00436444f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.295
cc_46 VNB N_VGND_c_581_n 0.00286581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_582_n 0.0199325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_583_n 0.00484152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_584_n 0.0158991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_585_n 0.0186449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_586_n 0.233221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_587_n 0.0249743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_588_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_589_n 0.00521838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_590_n 0.00362723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VPB N_C_N_M1011_g 0.0710742f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.86
cc_57 VPB N_D_N_M1006_g 0.0298502f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.86
cc_58 VPB N_D_N_M1001_g 0.0197316f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.455
cc_59 VPB N_D_N_c_134_n 0.0303619f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_60 VPB N_D_N_c_135_n 0.0172887f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_61 VPB N_A_196_530#_c_167_n 0.0173993f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.94
cc_62 VPB N_A_196_530#_c_177_n 0.0260697f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.445
cc_63 VPB N_A_196_530#_c_178_n 0.0171603f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.94
cc_64 VPB N_A_196_530#_c_179_n 0.00561199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_196_530#_c_180_n 0.0248098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_196_530#_c_181_n 0.0450595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_196_530#_c_182_n 0.0401164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_27_530#_c_238_n 0.00823641f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.455
cc_69 VPB N_A_27_530#_M1005_g 0.04153f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.775
cc_70 VPB N_A_27_530#_c_247_n 0.0563644f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.925
cc_71 VPB N_A_27_530#_c_241_n 0.0226838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_27_530#_c_243_n 0.00629733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_27_530#_c_244_n 0.001516f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_B_M1007_g 0.0518206f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.86
cc_75 VPB N_A_M1008_g 0.018658f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.86
cc_76 VPB N_A_M1003_g 0.0136653f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.455
cc_77 VPB A 0.00294587f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.775
cc_78 VPB N_A_c_361_n 0.0293796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_c_362_n 0.0100645f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.94
cc_80 VPB N_A_336_439#_M1000_g 0.0552944f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_81 VPB N_A_336_439#_c_408_n 0.00899814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_336_439#_c_417_n 0.0127979f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.94
cc_83 VPB N_A_336_439#_c_418_n 0.00339305f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_336_439#_c_419_n 0.0102665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A_336_439#_c_420_n 0.00226891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_336_439#_c_421_n 0.016419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_336_439#_c_422_n 4.19818e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_514_n 0.0055417f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.775
cc_89 VPB N_VPWR_c_515_n 0.0192038f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_90 VPB N_VPWR_c_516_n 0.0188084f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.94
cc_91 VPB N_VPWR_c_517_n 0.0757171f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.94
cc_92 VPB N_VPWR_c_518_n 0.0194346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_513_n 0.0879711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_520_n 0.00362799f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_521_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB X 0.0653138f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_97 N_C_N_M1011_g N_D_N_M1001_g 0.0175663f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_98 N_C_N_c_99_n N_D_N_M1001_g 0.0147153f $X=0.54 $Y=0.775 $X2=0 $Y2=0
cc_99 C_N N_D_N_M1001_g 0.0141256f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_100 N_C_N_c_103_n N_D_N_M1001_g 0.0332003f $X=0.54 $Y=0.94 $X2=0 $Y2=0
cc_101 N_C_N_M1011_g N_D_N_c_134_n 0.0364452f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_102 N_C_N_M1011_g N_D_N_c_135_n 0.00478363f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_103 C_N N_A_196_530#_c_173_n 0.00724055f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_104 N_C_N_M1011_g N_A_27_530#_c_240_n 0.00643487f $X=0.475 $Y=2.86 $X2=0
+ $Y2=0
cc_105 N_C_N_c_99_n N_A_27_530#_c_240_n 0.00523038f $X=0.54 $Y=0.775 $X2=0 $Y2=0
cc_106 C_N N_A_27_530#_c_240_n 0.0483715f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_107 N_C_N_c_103_n N_A_27_530#_c_240_n 0.0163648f $X=0.54 $Y=0.94 $X2=0 $Y2=0
cc_108 N_C_N_M1011_g N_A_27_530#_c_247_n 0.0262494f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_109 N_C_N_M1011_g N_A_27_530#_c_241_n 0.0187224f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_110 N_C_N_c_101_n N_A_27_530#_c_241_n 0.00208215f $X=0.54 $Y=1.445 $X2=0
+ $Y2=0
cc_111 C_N N_A_27_530#_c_241_n 0.0266946f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_112 C_N N_A_27_530#_c_242_n 9.70106e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_113 N_C_N_c_103_n N_A_27_530#_c_242_n 0.0036613f $X=0.54 $Y=0.94 $X2=0 $Y2=0
cc_114 N_C_N_M1011_g N_VPWR_c_514_n 0.00281249f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_115 N_C_N_M1011_g N_VPWR_c_516_n 0.00560159f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_116 N_C_N_M1011_g N_VPWR_c_513_n 0.0113779f $X=0.475 $Y=2.86 $X2=0 $Y2=0
cc_117 N_C_N_c_99_n N_VGND_c_578_n 0.00279829f $X=0.54 $Y=0.775 $X2=0 $Y2=0
cc_118 C_N N_VGND_c_578_n 0.00655112f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_119 N_C_N_c_99_n N_VGND_c_586_n 0.00710295f $X=0.54 $Y=0.775 $X2=0 $Y2=0
cc_120 C_N N_VGND_c_586_n 0.00816365f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_121 N_C_N_c_99_n N_VGND_c_587_n 0.00575161f $X=0.54 $Y=0.775 $X2=0 $Y2=0
cc_122 N_C_N_c_103_n N_VGND_c_587_n 5.03641e-19 $X=0.54 $Y=0.94 $X2=0 $Y2=0
cc_123 N_D_N_M1001_g N_A_196_530#_c_169_n 0.0430706f $X=1.02 $Y=0.455 $X2=0
+ $Y2=0
cc_124 N_D_N_c_134_n N_A_196_530#_c_179_n 0.0132326f $X=0.995 $Y=2.17 $X2=0
+ $Y2=0
cc_125 N_D_N_c_135_n N_A_196_530#_c_179_n 0.00174014f $X=0.995 $Y=2.17 $X2=0
+ $Y2=0
cc_126 N_D_N_c_134_n N_A_196_530#_c_180_n 6.45436e-19 $X=0.995 $Y=2.17 $X2=0
+ $Y2=0
cc_127 N_D_N_c_135_n N_A_196_530#_c_180_n 0.0110324f $X=0.995 $Y=2.17 $X2=0
+ $Y2=0
cc_128 N_D_N_M1006_g N_A_196_530#_c_181_n 0.00520023f $X=0.905 $Y=2.86 $X2=0
+ $Y2=0
cc_129 N_D_N_M1001_g N_A_196_530#_c_171_n 0.00280541f $X=1.02 $Y=0.455 $X2=0
+ $Y2=0
cc_130 N_D_N_M1001_g N_A_196_530#_c_173_n 0.00344588f $X=1.02 $Y=0.455 $X2=0
+ $Y2=0
cc_131 N_D_N_M1001_g N_A_196_530#_c_174_n 0.00276459f $X=1.02 $Y=0.455 $X2=0
+ $Y2=0
cc_132 N_D_N_M1006_g N_A_196_530#_c_182_n 0.00937892f $X=0.905 $Y=2.86 $X2=0
+ $Y2=0
cc_133 N_D_N_c_135_n N_A_196_530#_c_182_n 0.0022663f $X=0.995 $Y=2.17 $X2=0
+ $Y2=0
cc_134 N_D_N_c_135_n N_A_27_530#_c_247_n 0.0370317f $X=0.995 $Y=2.17 $X2=0 $Y2=0
cc_135 N_D_N_M1001_g N_A_27_530#_c_241_n 0.0162379f $X=1.02 $Y=0.455 $X2=0 $Y2=0
cc_136 N_D_N_c_134_n N_A_27_530#_c_241_n 0.00436449f $X=0.995 $Y=2.17 $X2=0
+ $Y2=0
cc_137 N_D_N_c_135_n N_A_27_530#_c_241_n 0.038721f $X=0.995 $Y=2.17 $X2=0 $Y2=0
cc_138 N_D_N_c_135_n N_A_336_439#_c_417_n 0.0121789f $X=0.995 $Y=2.17 $X2=0
+ $Y2=0
cc_139 N_D_N_M1006_g N_VPWR_c_514_n 0.00271017f $X=0.905 $Y=2.86 $X2=0 $Y2=0
cc_140 N_D_N_c_135_n N_VPWR_c_514_n 0.011706f $X=0.995 $Y=2.17 $X2=0 $Y2=0
cc_141 N_D_N_M1006_g N_VPWR_c_517_n 0.00560159f $X=0.905 $Y=2.86 $X2=0 $Y2=0
cc_142 N_D_N_M1006_g N_VPWR_c_513_n 0.00707422f $X=0.905 $Y=2.86 $X2=0 $Y2=0
cc_143 N_D_N_c_135_n N_VPWR_c_513_n 0.00947836f $X=0.995 $Y=2.17 $X2=0 $Y2=0
cc_144 N_D_N_M1001_g N_VGND_c_578_n 0.00279829f $X=1.02 $Y=0.455 $X2=0 $Y2=0
cc_145 N_D_N_M1001_g N_VGND_c_579_n 0.00575161f $X=1.02 $Y=0.455 $X2=0 $Y2=0
cc_146 N_D_N_M1001_g N_VGND_c_580_n 0.00443498f $X=1.02 $Y=0.455 $X2=0 $Y2=0
cc_147 N_D_N_M1001_g N_VGND_c_586_n 0.0119749f $X=1.02 $Y=0.455 $X2=0 $Y2=0
cc_148 N_A_196_530#_c_167_n N_A_27_530#_c_238_n 0.00590096f $X=1.53 $Y=1.935
+ $X2=0 $Y2=0
cc_149 N_A_196_530#_c_170_n N_A_27_530#_c_238_n 0.0028398f $X=1.62 $Y=1.445
+ $X2=0 $Y2=0
cc_150 N_A_196_530#_c_174_n N_A_27_530#_c_238_n 3.01862e-19 $X=1.62 $Y=0.94
+ $X2=0 $Y2=0
cc_151 N_A_196_530#_c_167_n N_A_27_530#_M1005_g 0.00399091f $X=1.53 $Y=1.935
+ $X2=0 $Y2=0
cc_152 N_A_196_530#_c_177_n N_A_27_530#_M1005_g 0.0532928f $X=1.945 $Y=2.01
+ $X2=0 $Y2=0
cc_153 N_A_196_530#_c_168_n N_A_27_530#_M1009_g 0.0233344f $X=1.97 $Y=0.775
+ $X2=0 $Y2=0
cc_154 N_A_196_530#_c_172_n N_A_27_530#_M1009_g 3.70416e-19 $X=1.535 $Y=0.82
+ $X2=0 $Y2=0
cc_155 N_A_196_530#_c_174_n N_A_27_530#_M1009_g 0.00208693f $X=1.62 $Y=0.94
+ $X2=0 $Y2=0
cc_156 N_A_196_530#_c_175_n N_A_27_530#_M1009_g 0.0108569f $X=1.62 $Y=0.94 $X2=0
+ $Y2=0
cc_157 N_A_196_530#_c_167_n N_A_27_530#_c_241_n 0.0191719f $X=1.53 $Y=1.935
+ $X2=0 $Y2=0
cc_158 N_A_196_530#_c_177_n N_A_27_530#_c_241_n 0.0120164f $X=1.945 $Y=2.01
+ $X2=0 $Y2=0
cc_159 N_A_196_530#_c_170_n N_A_27_530#_c_241_n 0.00236232f $X=1.62 $Y=1.445
+ $X2=0 $Y2=0
cc_160 N_A_196_530#_c_174_n N_A_27_530#_c_241_n 0.0126388f $X=1.62 $Y=0.94 $X2=0
+ $Y2=0
cc_161 N_A_196_530#_c_167_n N_A_27_530#_c_244_n 9.39097e-19 $X=1.53 $Y=1.935
+ $X2=0 $Y2=0
cc_162 N_A_196_530#_c_170_n N_A_27_530#_c_244_n 2.98616e-19 $X=1.62 $Y=1.445
+ $X2=0 $Y2=0
cc_163 N_A_196_530#_c_174_n N_A_27_530#_c_244_n 0.00224942f $X=1.62 $Y=0.94
+ $X2=0 $Y2=0
cc_164 N_A_196_530#_c_177_n N_A_336_439#_c_417_n 0.00344897f $X=1.945 $Y=2.01
+ $X2=0 $Y2=0
cc_165 N_A_196_530#_c_178_n N_A_336_439#_c_417_n 0.0135989f $X=2.02 $Y=2.085
+ $X2=0 $Y2=0
cc_166 N_A_196_530#_c_180_n N_A_336_439#_c_417_n 0.00254755f $X=1.57 $Y=2.94
+ $X2=0 $Y2=0
cc_167 N_A_196_530#_c_182_n N_A_336_439#_c_417_n 0.00467798f $X=1.57 $Y=2.775
+ $X2=0 $Y2=0
cc_168 N_A_196_530#_c_168_n N_A_336_439#_c_413_n 0.00267426f $X=1.97 $Y=0.775
+ $X2=0 $Y2=0
cc_169 N_A_196_530#_c_172_n N_A_336_439#_c_413_n 0.00282742f $X=1.535 $Y=0.82
+ $X2=0 $Y2=0
cc_170 N_A_196_530#_c_178_n N_VPWR_c_517_n 0.00370896f $X=2.02 $Y=2.085 $X2=0
+ $Y2=0
cc_171 N_A_196_530#_c_180_n N_VPWR_c_517_n 0.0352571f $X=1.57 $Y=2.94 $X2=0
+ $Y2=0
cc_172 N_A_196_530#_c_181_n N_VPWR_c_517_n 0.00617531f $X=1.57 $Y=2.94 $X2=0
+ $Y2=0
cc_173 N_A_196_530#_c_178_n N_VPWR_c_513_n 0.00445256f $X=2.02 $Y=2.085 $X2=0
+ $Y2=0
cc_174 N_A_196_530#_c_180_n N_VPWR_c_513_n 0.0251483f $X=1.57 $Y=2.94 $X2=0
+ $Y2=0
cc_175 N_A_196_530#_c_181_n N_VPWR_c_513_n 0.00817244f $X=1.57 $Y=2.94 $X2=0
+ $Y2=0
cc_176 N_A_196_530#_c_169_n N_VGND_c_579_n 6.38144e-19 $X=1.97 $Y=0.85 $X2=0
+ $Y2=0
cc_177 N_A_196_530#_c_171_n N_VGND_c_579_n 0.00831344f $X=1.235 $Y=0.52 $X2=0
+ $Y2=0
cc_178 N_A_196_530#_c_172_n N_VGND_c_579_n 0.00481021f $X=1.535 $Y=0.82 $X2=0
+ $Y2=0
cc_179 N_A_196_530#_c_168_n N_VGND_c_580_n 0.00323623f $X=1.97 $Y=0.775 $X2=0
+ $Y2=0
cc_180 N_A_196_530#_c_169_n N_VGND_c_580_n 0.00625657f $X=1.97 $Y=0.85 $X2=0
+ $Y2=0
cc_181 N_A_196_530#_c_171_n N_VGND_c_580_n 0.00915916f $X=1.235 $Y=0.52 $X2=0
+ $Y2=0
cc_182 N_A_196_530#_c_172_n N_VGND_c_580_n 0.00434437f $X=1.535 $Y=0.82 $X2=0
+ $Y2=0
cc_183 N_A_196_530#_c_168_n N_VGND_c_581_n 7.74981e-19 $X=1.97 $Y=0.775 $X2=0
+ $Y2=0
cc_184 N_A_196_530#_c_168_n N_VGND_c_584_n 0.00585385f $X=1.97 $Y=0.775 $X2=0
+ $Y2=0
cc_185 N_A_196_530#_c_169_n N_VGND_c_584_n 5.32051e-19 $X=1.97 $Y=0.85 $X2=0
+ $Y2=0
cc_186 N_A_196_530#_M1001_d N_VGND_c_586_n 0.00355226f $X=1.095 $Y=0.245 $X2=0
+ $Y2=0
cc_187 N_A_196_530#_c_168_n N_VGND_c_586_n 0.0120255f $X=1.97 $Y=0.775 $X2=0
+ $Y2=0
cc_188 N_A_196_530#_c_169_n N_VGND_c_586_n 7.38536e-19 $X=1.97 $Y=0.85 $X2=0
+ $Y2=0
cc_189 N_A_196_530#_c_171_n N_VGND_c_586_n 0.00760397f $X=1.235 $Y=0.52 $X2=0
+ $Y2=0
cc_190 N_A_196_530#_c_172_n N_VGND_c_586_n 0.00868133f $X=1.535 $Y=0.82 $X2=0
+ $Y2=0
cc_191 N_A_27_530#_c_238_n N_B_M1007_g 0.0378751f $X=2.38 $Y=1.695 $X2=0 $Y2=0
cc_192 N_A_27_530#_c_244_n N_B_M1007_g 6.37062e-19 $X=2.29 $Y=1.53 $X2=0 $Y2=0
cc_193 N_A_27_530#_M1009_g N_B_M1013_g 0.0205467f $X=2.4 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A_27_530#_c_238_n N_B_c_314_n 0.0189458f $X=2.38 $Y=1.695 $X2=0 $Y2=0
cc_195 N_A_27_530#_c_238_n N_B_c_315_n 0.00311846f $X=2.38 $Y=1.695 $X2=0 $Y2=0
cc_196 N_A_27_530#_c_244_n N_B_c_315_n 4.74286e-19 $X=2.29 $Y=1.53 $X2=0 $Y2=0
cc_197 N_A_27_530#_M1009_g N_B_c_316_n 0.0189458f $X=2.4 $Y=0.445 $X2=0 $Y2=0
cc_198 N_A_27_530#_M1009_g N_B_c_317_n 0.0114328f $X=2.4 $Y=0.445 $X2=0 $Y2=0
cc_199 N_A_27_530#_c_244_n N_B_c_317_n 0.00889262f $X=2.29 $Y=1.53 $X2=0 $Y2=0
cc_200 N_A_27_530#_c_238_n N_A_336_439#_c_417_n 0.00149474f $X=2.38 $Y=1.695
+ $X2=0 $Y2=0
cc_201 N_A_27_530#_M1005_g N_A_336_439#_c_417_n 0.0210257f $X=2.38 $Y=2.405
+ $X2=0 $Y2=0
cc_202 N_A_27_530#_c_241_n N_A_336_439#_c_417_n 0.0222801f $X=2.205 $Y=1.71
+ $X2=0 $Y2=0
cc_203 N_A_27_530#_c_244_n N_A_336_439#_c_417_n 0.00760979f $X=2.29 $Y=1.53
+ $X2=0 $Y2=0
cc_204 N_A_27_530#_M1009_g N_A_336_439#_c_409_n 0.0141596f $X=2.4 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_A_27_530#_c_244_n N_A_336_439#_c_409_n 0.00239836f $X=2.29 $Y=1.53
+ $X2=0 $Y2=0
cc_206 N_A_27_530#_M1005_g N_A_336_439#_c_418_n 0.00675867f $X=2.38 $Y=2.405
+ $X2=0 $Y2=0
cc_207 N_A_27_530#_c_238_n N_A_336_439#_c_420_n 0.0021675f $X=2.38 $Y=1.695
+ $X2=0 $Y2=0
cc_208 N_A_27_530#_c_244_n N_A_336_439#_c_420_n 0.00669684f $X=2.29 $Y=1.53
+ $X2=0 $Y2=0
cc_209 N_A_27_530#_c_238_n N_A_336_439#_c_413_n 0.00272276f $X=2.38 $Y=1.695
+ $X2=0 $Y2=0
cc_210 N_A_27_530#_M1009_g N_A_336_439#_c_413_n 3.46155e-19 $X=2.4 $Y=0.445
+ $X2=0 $Y2=0
cc_211 N_A_27_530#_c_244_n N_A_336_439#_c_413_n 0.0027592f $X=2.29 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_27_530#_c_247_n N_VPWR_c_516_n 0.00999318f $X=0.26 $Y=2.795 $X2=0
+ $Y2=0
cc_213 N_A_27_530#_M1005_g N_VPWR_c_517_n 0.00370896f $X=2.38 $Y=2.405 $X2=0
+ $Y2=0
cc_214 N_A_27_530#_M1005_g N_VPWR_c_513_n 0.00445256f $X=2.38 $Y=2.405 $X2=0
+ $Y2=0
cc_215 N_A_27_530#_c_247_n N_VPWR_c_513_n 0.00941316f $X=0.26 $Y=2.795 $X2=0
+ $Y2=0
cc_216 N_A_27_530#_M1009_g N_VGND_c_581_n 0.00620585f $X=2.4 $Y=0.445 $X2=0
+ $Y2=0
cc_217 N_A_27_530#_M1009_g N_VGND_c_584_n 0.00408791f $X=2.4 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_A_27_530#_M1010_s N_VGND_c_586_n 0.00231734f $X=0.25 $Y=0.245 $X2=0
+ $Y2=0
cc_219 N_A_27_530#_M1009_g N_VGND_c_586_n 0.00477058f $X=2.4 $Y=0.445 $X2=0
+ $Y2=0
cc_220 N_A_27_530#_c_242_n N_VGND_c_586_n 0.0142319f $X=0.375 $Y=0.43 $X2=0
+ $Y2=0
cc_221 N_A_27_530#_c_242_n N_VGND_c_587_n 0.0229133f $X=0.375 $Y=0.43 $X2=0
+ $Y2=0
cc_222 N_B_M1007_g N_A_M1003_g 0.0149625f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_223 N_B_M1013_g N_A_M1003_g 0.0203905f $X=2.91 $Y=0.445 $X2=0 $Y2=0
cc_224 N_B_c_316_n N_A_M1003_g 0.0344824f $X=2.85 $Y=1.06 $X2=0 $Y2=0
cc_225 N_B_c_317_n N_A_M1003_g 5.71637e-19 $X=2.85 $Y=1.06 $X2=0 $Y2=0
cc_226 N_B_M1007_g A 0.0102124f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_227 N_B_M1007_g N_A_c_361_n 0.0613806f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_228 N_B_M1007_g N_A_c_362_n 0.00203786f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_229 N_B_M1007_g N_A_336_439#_c_417_n 0.00947252f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_230 N_B_M1013_g N_A_336_439#_c_409_n 0.0107961f $X=2.91 $Y=0.445 $X2=0 $Y2=0
cc_231 N_B_c_316_n N_A_336_439#_c_409_n 0.00510554f $X=2.85 $Y=1.06 $X2=0 $Y2=0
cc_232 N_B_c_317_n N_A_336_439#_c_409_n 0.0342561f $X=2.85 $Y=1.06 $X2=0 $Y2=0
cc_233 N_B_M1007_g N_A_336_439#_c_418_n 0.0079447f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_234 N_B_M1007_g N_A_336_439#_c_419_n 0.0101574f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_235 N_B_c_315_n N_A_336_439#_c_419_n 0.00142434f $X=2.85 $Y=1.565 $X2=0 $Y2=0
cc_236 N_B_c_317_n N_A_336_439#_c_419_n 0.0114648f $X=2.85 $Y=1.06 $X2=0 $Y2=0
cc_237 N_B_M1007_g N_A_336_439#_c_420_n 0.00269752f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_238 N_B_c_315_n N_A_336_439#_c_420_n 0.00381978f $X=2.85 $Y=1.565 $X2=0 $Y2=0
cc_239 N_B_c_317_n N_A_336_439#_c_420_n 0.0139705f $X=2.85 $Y=1.06 $X2=0 $Y2=0
cc_240 N_B_M1007_g N_A_336_439#_c_410_n 0.00192272f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_241 N_B_M1013_g N_A_336_439#_c_410_n 0.00195025f $X=2.91 $Y=0.445 $X2=0 $Y2=0
cc_242 N_B_c_315_n N_A_336_439#_c_410_n 0.00167619f $X=2.85 $Y=1.565 $X2=0 $Y2=0
cc_243 N_B_c_316_n N_A_336_439#_c_410_n 0.00324336f $X=2.85 $Y=1.06 $X2=0 $Y2=0
cc_244 N_B_c_317_n N_A_336_439#_c_410_n 0.0376138f $X=2.85 $Y=1.06 $X2=0 $Y2=0
cc_245 N_B_M1013_g N_A_336_439#_c_414_n 3.46474e-19 $X=2.91 $Y=0.445 $X2=0 $Y2=0
cc_246 N_B_M1007_g N_VPWR_c_517_n 0.00497279f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_247 N_B_M1007_g N_VPWR_c_513_n 0.00509887f $X=2.89 $Y=2.635 $X2=0 $Y2=0
cc_248 N_B_M1013_g N_VGND_c_581_n 0.00428262f $X=2.91 $Y=0.445 $X2=0 $Y2=0
cc_249 N_B_M1013_g N_VGND_c_582_n 0.0042361f $X=2.91 $Y=0.445 $X2=0 $Y2=0
cc_250 N_B_M1013_g N_VGND_c_586_n 0.00607497f $X=2.91 $Y=0.445 $X2=0 $Y2=0
cc_251 N_A_M1008_g N_A_336_439#_M1000_g 0.0152238f $X=3.25 $Y=2.635 $X2=0 $Y2=0
cc_252 N_A_M1003_g N_A_336_439#_M1000_g 0.00888894f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_253 A N_A_336_439#_M1000_g 0.00133901f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_254 N_A_c_361_n N_A_336_439#_M1000_g 0.0168826f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_255 N_A_c_362_n N_A_336_439#_M1000_g 0.00154828f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_256 N_A_M1003_g N_A_336_439#_M1012_g 0.0233804f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_257 A N_A_336_439#_c_417_n 0.0140468f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_258 N_A_c_362_n N_A_336_439#_c_417_n 0.0119407f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_259 N_A_M1003_g N_A_336_439#_c_418_n 4.96517e-19 $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_260 N_A_c_361_n N_A_336_439#_c_418_n 5.84301e-19 $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_261 N_A_c_362_n N_A_336_439#_c_418_n 0.0118708f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_262 N_A_c_361_n N_A_336_439#_c_419_n 5.72167e-19 $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_263 N_A_c_362_n N_A_336_439#_c_419_n 0.0119902f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_264 N_A_M1003_g N_A_336_439#_c_410_n 0.0215008f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_265 N_A_M1003_g N_A_336_439#_c_421_n 0.00576584f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_266 N_A_c_361_n N_A_336_439#_c_421_n 0.00220412f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_267 N_A_c_362_n N_A_336_439#_c_421_n 0.00979631f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_268 N_A_M1003_g N_A_336_439#_c_411_n 0.00178859f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_269 N_A_M1003_g N_A_336_439#_c_412_n 0.0395529f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_M1003_g N_A_336_439#_c_414_n 0.0117168f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_271 N_A_M1003_g N_A_336_439#_c_422_n 0.00519425f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_272 N_A_c_361_n N_A_336_439#_c_422_n 0.00208286f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_273 N_A_c_362_n N_A_336_439#_c_422_n 0.0131585f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_274 N_A_M1008_g N_VPWR_c_515_n 0.00480439f $X=3.25 $Y=2.635 $X2=0 $Y2=0
cc_275 A N_VPWR_c_515_n 0.0224028f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_276 N_A_c_361_n N_VPWR_c_515_n 7.92143e-19 $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_277 N_A_c_362_n N_VPWR_c_515_n 0.00725603f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_278 N_A_M1008_g N_VPWR_c_517_n 0.004712f $X=3.25 $Y=2.635 $X2=0 $Y2=0
cc_279 A N_VPWR_c_517_n 0.00570712f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_280 N_A_M1008_g N_VPWR_c_513_n 0.00509887f $X=3.25 $Y=2.635 $X2=0 $Y2=0
cc_281 A N_VPWR_c_513_n 0.00587701f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_282 A A_593_485# 0.00440771f $X=3.035 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_283 N_A_c_362_n X 0.0098176f $X=3.34 $Y=2.1 $X2=0 $Y2=0
cc_284 N_A_M1003_g N_VGND_c_582_n 0.00447054f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_285 N_A_M1003_g N_VGND_c_583_n 0.00629493f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_286 N_A_M1003_g N_VGND_c_586_n 0.00758342f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_287 N_A_336_439#_M1000_g N_VPWR_c_515_n 0.00417256f $X=3.825 $Y=2.635 $X2=0
+ $Y2=0
cc_288 N_A_336_439#_M1000_g N_VPWR_c_518_n 0.00497279f $X=3.825 $Y=2.635 $X2=0
+ $Y2=0
cc_289 N_A_336_439#_M1000_g N_VPWR_c_513_n 0.00509887f $X=3.825 $Y=2.635 $X2=0
+ $Y2=0
cc_290 N_A_336_439#_c_417_n N_VPWR_c_513_n 0.0408897f $X=2.685 $Y=2.34 $X2=0
+ $Y2=0
cc_291 N_A_336_439#_c_417_n A_419_439# 0.0020643f $X=2.685 $Y=2.34 $X2=-0.19
+ $Y2=-0.245
cc_292 N_A_336_439#_c_417_n A_491_439# 0.00541f $X=2.685 $Y=2.34 $X2=-0.19
+ $Y2=-0.245
cc_293 N_A_336_439#_M1012_g N_X_c_560_n 5.67952e-19 $X=3.845 $Y=0.445 $X2=0
+ $Y2=0
cc_294 N_A_336_439#_c_414_n N_X_c_560_n 0.00207433f $X=3.125 $Y=0.51 $X2=0 $Y2=0
cc_295 N_A_336_439#_M1000_g X 0.0236618f $X=3.825 $Y=2.635 $X2=0 $Y2=0
cc_296 N_A_336_439#_M1012_g X 0.0124105f $X=3.845 $Y=0.445 $X2=0 $Y2=0
cc_297 N_A_336_439#_c_408_n X 5.56488e-19 $X=3.79 $Y=1.695 $X2=0 $Y2=0
cc_298 N_A_336_439#_c_421_n X 0.0129667f $X=3.705 $Y=1.75 $X2=0 $Y2=0
cc_299 N_A_336_439#_c_411_n X 0.0437496f $X=3.79 $Y=1.19 $X2=0 $Y2=0
cc_300 N_A_336_439#_c_412_n X 0.0163644f $X=3.79 $Y=1.19 $X2=0 $Y2=0
cc_301 N_A_336_439#_c_409_n N_VGND_M1009_d 0.00256658f $X=3.02 $Y=0.71 $X2=0
+ $Y2=0
cc_302 N_A_336_439#_c_409_n N_VGND_c_581_n 0.0179938f $X=3.02 $Y=0.71 $X2=0
+ $Y2=0
cc_303 N_A_336_439#_c_409_n N_VGND_c_582_n 0.00319405f $X=3.02 $Y=0.71 $X2=0
+ $Y2=0
cc_304 N_A_336_439#_c_414_n N_VGND_c_582_n 0.0131793f $X=3.125 $Y=0.51 $X2=0
+ $Y2=0
cc_305 N_A_336_439#_M1012_g N_VGND_c_583_n 0.00297074f $X=3.845 $Y=0.445 $X2=0
+ $Y2=0
cc_306 N_A_336_439#_c_411_n N_VGND_c_583_n 6.50494e-19 $X=3.79 $Y=1.19 $X2=0
+ $Y2=0
cc_307 N_A_336_439#_c_412_n N_VGND_c_583_n 0.00285905f $X=3.79 $Y=1.19 $X2=0
+ $Y2=0
cc_308 N_A_336_439#_c_414_n N_VGND_c_583_n 0.014295f $X=3.125 $Y=0.51 $X2=0
+ $Y2=0
cc_309 N_A_336_439#_c_409_n N_VGND_c_584_n 0.00275886f $X=3.02 $Y=0.71 $X2=0
+ $Y2=0
cc_310 N_A_336_439#_c_413_n N_VGND_c_584_n 0.00749266f $X=2.185 $Y=0.53 $X2=0
+ $Y2=0
cc_311 N_A_336_439#_M1012_g N_VGND_c_585_n 0.00585385f $X=3.845 $Y=0.445 $X2=0
+ $Y2=0
cc_312 N_A_336_439#_M1002_d N_VGND_c_586_n 0.00370623f $X=2.045 $Y=0.235 $X2=0
+ $Y2=0
cc_313 N_A_336_439#_M1013_d N_VGND_c_586_n 0.00243781f $X=2.985 $Y=0.235 $X2=0
+ $Y2=0
cc_314 N_A_336_439#_M1012_g N_VGND_c_586_n 0.0118985f $X=3.845 $Y=0.445 $X2=0
+ $Y2=0
cc_315 N_A_336_439#_c_409_n N_VGND_c_586_n 0.0115767f $X=3.02 $Y=0.71 $X2=0
+ $Y2=0
cc_316 N_A_336_439#_c_413_n N_VGND_c_586_n 0.0074948f $X=2.185 $Y=0.53 $X2=0
+ $Y2=0
cc_317 N_A_336_439#_c_414_n N_VGND_c_586_n 0.0121309f $X=3.125 $Y=0.51 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_515_n X 0.00440091f $X=3.55 $Y=2.7 $X2=0 $Y2=0
cc_319 N_VPWR_c_518_n X 0.00997542f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_320 N_VPWR_c_513_n X 0.0101536f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_321 N_X_c_560_n N_VGND_c_585_n 0.0113196f $X=4.06 $Y=0.51 $X2=0 $Y2=0
cc_322 N_X_M1012_d N_VGND_c_586_n 0.0034811f $X=3.92 $Y=0.235 $X2=0 $Y2=0
cc_323 N_X_c_560_n N_VGND_c_586_n 0.00984396f $X=4.06 $Y=0.51 $X2=0 $Y2=0
