* File: sky130_fd_sc_lp__nor2_8.pex.spice
* Created: Wed Sep  2 10:07:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2_8%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 65 66 67 68 92
c142 63 0 1.22355e-19 $X=3.585 $Y=2.465
r143 91 92 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.155 $Y=1.51
+ $X2=3.585 $Y2=1.51
r144 90 91 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.725 $Y=1.51
+ $X2=3.155 $Y2=1.51
r145 89 90 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.295 $Y=1.51
+ $X2=2.725 $Y2=1.51
r146 87 89 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=2.025 $Y=1.51
+ $X2=2.295 $Y2=1.51
r147 87 88 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.025
+ $Y=1.51 $X2=2.025 $Y2=1.51
r148 85 87 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.865 $Y=1.51
+ $X2=2.025 $Y2=1.51
r149 84 88 11.0375 $w=3.53e-07 $l=3.4e-07 $layer=LI1_cond $X=1.685 $Y=1.592
+ $X2=2.025 $Y2=1.592
r150 83 85 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.685 $Y=1.51
+ $X2=1.865 $Y2=1.51
r151 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.685
+ $Y=1.51 $X2=1.685 $Y2=1.51
r152 81 83 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.435 $Y=1.51
+ $X2=1.685 $Y2=1.51
r153 79 81 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.345 $Y=1.51
+ $X2=1.435 $Y2=1.51
r154 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.345
+ $Y=1.51 $X2=1.345 $Y2=1.51
r155 76 79 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.005 $Y=1.51
+ $X2=1.345 $Y2=1.51
r156 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.005
+ $Y=1.51 $X2=1.005 $Y2=1.51
r157 73 76 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.575 $Y=1.51
+ $X2=1.005 $Y2=1.51
r158 68 88 4.38253 $w=3.53e-07 $l=1.35e-07 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=2.025 $Y2=1.592
r159 67 84 0.162316 $w=3.53e-07 $l=5e-09 $layer=LI1_cond $X=1.68 $Y=1.592
+ $X2=1.685 $Y2=1.592
r160 67 80 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=1.68 $Y=1.592
+ $X2=1.345 $Y2=1.592
r161 66 80 4.70716 $w=3.53e-07 $l=1.45e-07 $layer=LI1_cond $X=1.2 $Y=1.592
+ $X2=1.345 $Y2=1.592
r162 66 77 6.33032 $w=3.53e-07 $l=1.95e-07 $layer=LI1_cond $X=1.2 $Y=1.592
+ $X2=1.005 $Y2=1.592
r163 65 77 9.25201 $w=3.53e-07 $l=2.85e-07 $layer=LI1_cond $X=0.72 $Y=1.592
+ $X2=1.005 $Y2=1.592
r164 61 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=1.675
+ $X2=3.585 $Y2=1.51
r165 61 63 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.585 $Y=1.675
+ $X2=3.585 $Y2=2.465
r166 57 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=1.345
+ $X2=3.585 $Y2=1.51
r167 57 59 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.585 $Y=1.345
+ $X2=3.585 $Y2=0.745
r168 53 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.155 $Y=1.675
+ $X2=3.155 $Y2=1.51
r169 53 55 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.155 $Y=1.675
+ $X2=3.155 $Y2=2.465
r170 49 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.155 $Y=1.345
+ $X2=3.155 $Y2=1.51
r171 49 51 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.155 $Y=1.345
+ $X2=3.155 $Y2=0.745
r172 45 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.675
+ $X2=2.725 $Y2=1.51
r173 45 47 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.725 $Y=1.675
+ $X2=2.725 $Y2=2.465
r174 41 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.725 $Y=1.345
+ $X2=2.725 $Y2=1.51
r175 41 43 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.725 $Y=1.345
+ $X2=2.725 $Y2=0.745
r176 37 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.675
+ $X2=2.295 $Y2=1.51
r177 37 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.295 $Y=1.675
+ $X2=2.295 $Y2=2.465
r178 33 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.345
+ $X2=2.295 $Y2=1.51
r179 33 35 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.295 $Y=1.345
+ $X2=2.295 $Y2=0.745
r180 29 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.675
+ $X2=1.865 $Y2=1.51
r181 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.865 $Y=1.675
+ $X2=1.865 $Y2=2.465
r182 25 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.345
+ $X2=1.865 $Y2=1.51
r183 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.865 $Y=1.345
+ $X2=1.865 $Y2=0.745
r184 21 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.675
+ $X2=1.435 $Y2=1.51
r185 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.435 $Y=1.675
+ $X2=1.435 $Y2=2.465
r186 17 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.345
+ $X2=1.435 $Y2=1.51
r187 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.435 $Y=1.345
+ $X2=1.435 $Y2=0.745
r188 13 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.675
+ $X2=1.005 $Y2=1.51
r189 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.005 $Y=1.675
+ $X2=1.005 $Y2=2.465
r190 9 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.345
+ $X2=1.005 $Y2=1.51
r191 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.005 $Y=1.345
+ $X2=1.005 $Y2=0.745
r192 5 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.675
+ $X2=0.575 $Y2=1.51
r193 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.575 $Y=1.675
+ $X2=0.575 $Y2=2.465
r194 1 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.345
+ $X2=0.575 $Y2=1.51
r195 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.575 $Y=1.345 $X2=0.575
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_8%B 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 65 66 67 68 93
r151 91 93 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=6.665 $Y=1.51
+ $X2=7.025 $Y2=1.51
r152 91 92 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.665
+ $Y=1.51 $X2=6.665 $Y2=1.51
r153 89 91 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.595 $Y=1.51
+ $X2=6.665 $Y2=1.51
r154 87 89 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=6.325 $Y=1.51
+ $X2=6.595 $Y2=1.51
r155 87 88 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.325
+ $Y=1.51 $X2=6.325 $Y2=1.51
r156 85 87 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.165 $Y=1.51
+ $X2=6.325 $Y2=1.51
r157 83 85 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.985 $Y=1.51
+ $X2=6.165 $Y2=1.51
r158 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.985
+ $Y=1.51 $X2=5.985 $Y2=1.51
r159 81 83 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.735 $Y=1.51
+ $X2=5.985 $Y2=1.51
r160 80 84 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=5.645 $Y=1.587
+ $X2=5.985 $Y2=1.587
r161 79 81 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.645 $Y=1.51
+ $X2=5.735 $Y2=1.51
r162 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.645
+ $Y=1.51 $X2=5.645 $Y2=1.51
r163 77 79 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.305 $Y=1.51
+ $X2=5.645 $Y2=1.51
r164 76 77 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.875 $Y=1.51
+ $X2=5.305 $Y2=1.51
r165 75 76 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.445 $Y=1.51
+ $X2=4.875 $Y2=1.51
r166 73 75 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.015 $Y=1.51
+ $X2=4.445 $Y2=1.51
r167 68 92 10.4606 $w=3.23e-07 $l=2.95e-07 $layer=LI1_cond $X=6.96 $Y=1.587
+ $X2=6.665 $Y2=1.587
r168 67 92 6.56006 $w=3.23e-07 $l=1.85e-07 $layer=LI1_cond $X=6.48 $Y=1.587
+ $X2=6.665 $Y2=1.587
r169 67 88 5.49627 $w=3.23e-07 $l=1.55e-07 $layer=LI1_cond $X=6.48 $Y=1.587
+ $X2=6.325 $Y2=1.587
r170 66 88 11.5244 $w=3.23e-07 $l=3.25e-07 $layer=LI1_cond $X=6 $Y=1.587
+ $X2=6.325 $Y2=1.587
r171 66 84 0.531897 $w=3.23e-07 $l=1.5e-08 $layer=LI1_cond $X=6 $Y=1.587
+ $X2=5.985 $Y2=1.587
r172 65 80 4.43247 $w=3.23e-07 $l=1.25e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.645 $Y2=1.587
r173 61 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.675
+ $X2=7.025 $Y2=1.51
r174 61 63 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.025 $Y=1.675
+ $X2=7.025 $Y2=2.465
r175 57 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.345
+ $X2=7.025 $Y2=1.51
r176 57 59 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.025 $Y=1.345
+ $X2=7.025 $Y2=0.745
r177 53 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.675
+ $X2=6.595 $Y2=1.51
r178 53 55 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.595 $Y=1.675
+ $X2=6.595 $Y2=2.465
r179 49 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.345
+ $X2=6.595 $Y2=1.51
r180 49 51 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.595 $Y=1.345
+ $X2=6.595 $Y2=0.745
r181 45 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.165 $Y=1.675
+ $X2=6.165 $Y2=1.51
r182 45 47 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.165 $Y=1.675
+ $X2=6.165 $Y2=2.465
r183 41 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.165 $Y=1.345
+ $X2=6.165 $Y2=1.51
r184 41 43 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.165 $Y=1.345
+ $X2=6.165 $Y2=0.745
r185 37 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=1.675
+ $X2=5.735 $Y2=1.51
r186 37 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.735 $Y=1.675
+ $X2=5.735 $Y2=2.465
r187 33 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=1.345
+ $X2=5.735 $Y2=1.51
r188 33 35 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.735 $Y=1.345
+ $X2=5.735 $Y2=0.745
r189 29 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.675
+ $X2=5.305 $Y2=1.51
r190 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.305 $Y=1.675
+ $X2=5.305 $Y2=2.465
r191 25 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.345
+ $X2=5.305 $Y2=1.51
r192 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.305 $Y=1.345
+ $X2=5.305 $Y2=0.745
r193 21 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.875 $Y=1.675
+ $X2=4.875 $Y2=1.51
r194 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.875 $Y=1.675
+ $X2=4.875 $Y2=2.465
r195 17 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.875 $Y=1.345
+ $X2=4.875 $Y2=1.51
r196 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.875 $Y=1.345
+ $X2=4.875 $Y2=0.745
r197 13 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.675
+ $X2=4.445 $Y2=1.51
r198 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.445 $Y=1.675
+ $X2=4.445 $Y2=2.465
r199 9 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.345
+ $X2=4.445 $Y2=1.51
r200 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.445 $Y=1.345
+ $X2=4.445 $Y2=0.745
r201 5 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.675
+ $X2=4.015 $Y2=1.51
r202 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.015 $Y=1.675
+ $X2=4.015 $Y2=2.465
r203 1 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.345
+ $X2=4.015 $Y2=1.51
r204 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.015 $Y=1.345 $X2=4.015
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_8%A_47_367# 1 2 3 4 5 6 7 8 9 28 30 32 36 38 42
+ 44 48 50 53 56 60 62 66 68 72 74 78 83 85 86 94 95 96
r103 86 89 9.08914 $w=2.03e-07 $l=1.68e-07 $layer=LI1_cond $X=2.932 $Y=1.812
+ $X2=2.932 $Y2=1.98
r104 76 78 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=7.275 $Y=2.895
+ $X2=7.275 $Y2=2.425
r105 75 96 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.475 $Y=2.985
+ $X2=6.38 $Y2=2.985
r106 74 76 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=7.145 $Y=2.985
+ $X2=7.275 $Y2=2.895
r107 74 75 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.145 $Y=2.985
+ $X2=6.475 $Y2=2.985
r108 70 96 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=6.38 $Y=2.895 $X2=6.38
+ $Y2=2.985
r109 70 72 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=6.38 $Y=2.895
+ $X2=6.38 $Y2=2.425
r110 69 95 5.52892 $w=1.75e-07 $l=9.5e-08 $layer=LI1_cond $X=5.615 $Y=2.985
+ $X2=5.52 $Y2=2.985
r111 68 96 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.285 $Y=2.985
+ $X2=6.38 $Y2=2.985
r112 68 69 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=6.285 $Y=2.985
+ $X2=5.615 $Y2=2.985
r113 64 95 1.04816 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=5.52 $Y=2.895 $X2=5.52
+ $Y2=2.985
r114 64 66 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=5.52 $Y=2.895
+ $X2=5.52 $Y2=2.425
r115 63 94 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.755 $Y=2.99
+ $X2=4.66 $Y2=2.99
r116 62 95 5.52892 $w=1.75e-07 $l=9.74679e-08 $layer=LI1_cond $X=5.425 $Y=2.99
+ $X2=5.52 $Y2=2.985
r117 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.425 $Y=2.99
+ $X2=4.755 $Y2=2.99
r118 58 94 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=2.905
+ $X2=4.66 $Y2=2.99
r119 58 60 28.0191 $w=1.88e-07 $l=4.8e-07 $layer=LI1_cond $X=4.66 $Y=2.905
+ $X2=4.66 $Y2=2.425
r120 57 93 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.895 $Y=2.99
+ $X2=3.8 $Y2=2.99
r121 56 94 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.565 $Y=2.99
+ $X2=4.66 $Y2=2.99
r122 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.565 $Y=2.99
+ $X2=3.895 $Y2=2.99
r123 53 93 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=2.905 $X2=3.8
+ $Y2=2.99
r124 53 55 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=3.8 $Y=2.905
+ $X2=3.8 $Y2=1.98
r125 52 55 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=3.8 $Y=1.925
+ $X2=3.8 $Y2=1.98
r126 51 86 0.170324 $w=2.25e-07 $l=1.03e-07 $layer=LI1_cond $X=3.035 $Y=1.812
+ $X2=2.932 $Y2=1.812
r127 50 52 6.87974 $w=2.25e-07 $l=1.5331e-07 $layer=LI1_cond $X=3.705 $Y=1.812
+ $X2=3.8 $Y2=1.925
r128 50 51 34.3172 $w=2.23e-07 $l=6.7e-07 $layer=LI1_cond $X=3.705 $Y=1.812
+ $X2=3.035 $Y2=1.812
r129 48 91 19.8469 $w=1.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.94 $Y=2.45
+ $X2=2.94 $Y2=2.11
r130 45 85 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.175 $Y=2.025
+ $X2=2.08 $Y2=2.025
r131 44 91 4.67556 $w=2.03e-07 $l=8.5e-08 $layer=LI1_cond $X=2.932 $Y=2.025
+ $X2=2.932 $Y2=2.11
r132 44 89 2.43459 $w=2.03e-07 $l=4.5e-08 $layer=LI1_cond $X=2.932 $Y=2.025
+ $X2=2.932 $Y2=1.98
r133 44 45 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.83 $Y=2.025
+ $X2=2.175 $Y2=2.025
r134 40 85 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=2.11
+ $X2=2.08 $Y2=2.025
r135 40 42 46.6986 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=2.08 $Y=2.11 $X2=2.08
+ $Y2=2.91
r136 39 83 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.315 $Y=2.025
+ $X2=1.22 $Y2=2.025
r137 38 85 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.985 $Y=2.025
+ $X2=2.08 $Y2=2.025
r138 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.985 $Y=2.025
+ $X2=1.315 $Y2=2.025
r139 34 83 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.11
+ $X2=1.22 $Y2=2.025
r140 34 36 46.6986 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=1.22 $Y=2.11 $X2=1.22
+ $Y2=2.91
r141 33 81 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.455 $Y=2.025
+ $X2=0.32 $Y2=2.025
r142 32 83 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.125 $Y=2.025
+ $X2=1.22 $Y2=2.025
r143 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.125 $Y=2.025
+ $X2=0.455 $Y2=2.025
r144 28 81 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.32 $Y=2.11
+ $X2=0.32 $Y2=2.025
r145 28 30 34.1465 $w=2.68e-07 $l=8e-07 $layer=LI1_cond $X=0.32 $Y=2.11 $X2=0.32
+ $Y2=2.91
r146 9 78 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=7.1
+ $Y=1.835 $X2=7.24 $Y2=2.425
r147 8 72 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=6.24
+ $Y=1.835 $X2=6.38 $Y2=2.425
r148 7 66 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=5.38
+ $Y=1.835 $X2=5.52 $Y2=2.425
r149 6 60 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=4.52
+ $Y=1.835 $X2=4.66 $Y2=2.425
r150 5 93 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=1.835 $X2=3.8 $Y2=2.91
r151 5 55 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=1.835 $X2=3.8 $Y2=1.98
r152 4 89 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.835 $X2=2.94 $Y2=1.98
r153 4 48 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=2.8
+ $Y=1.835 $X2=2.94 $Y2=2.45
r154 3 85 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.08 $Y2=2.105
r155 3 42 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.08 $Y2=2.91
r156 2 83 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.22 $Y2=2.105
r157 2 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.22 $Y2=2.91
r158 1 81 400 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.835 $X2=0.36 $Y2=2.105
r159 1 30 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.835 $X2=0.36 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_8%VPWR 1 2 3 4 15 19 23 27 32 33 35 36 37 39 44
+ 60 61 64 67
r107 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 60 61 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 57 60 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r111 57 58 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r112 55 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r113 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 52 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.65 $Y2=3.33
r118 49 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 48 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r121 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r122 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.79 $Y2=3.33
r123 45 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.65 $Y2=3.33
r125 44 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 42 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r128 39 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.79 $Y2=3.33
r129 39 41 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r130 37 61 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=7.44 $Y2=3.33
r131 37 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r132 35 54 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=3.12 $Y2=3.33
r133 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=3.37 $Y2=3.33
r134 34 57 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.535 $Y=3.33
+ $X2=3.6 $Y2=3.33
r135 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.535 $Y=3.33
+ $X2=3.37 $Y2=3.33
r136 32 51 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=3.33
+ $X2=2.51 $Y2=3.33
r138 31 54 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.675 $Y=3.33
+ $X2=3.12 $Y2=3.33
r139 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=3.33
+ $X2=2.51 $Y2=3.33
r140 27 30 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.37 $Y=2.18
+ $X2=3.37 $Y2=2.95
r141 25 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.37 $Y=3.245
+ $X2=3.37 $Y2=3.33
r142 25 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.37 $Y=3.245
+ $X2=3.37 $Y2=2.95
r143 21 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=3.33
r144 21 23 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=2.365
r145 17 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=3.33
r146 17 19 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=2.365
r147 13 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=3.33
r148 13 15 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=2.365
r149 4 30 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.835 $X2=3.37 $Y2=2.95
r150 4 27 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.835 $X2=3.37 $Y2=2.18
r151 3 23 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=2.37
+ $Y=1.835 $X2=2.51 $Y2=2.365
r152 2 19 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=1.51
+ $Y=1.835 $X2=1.65 $Y2=2.365
r153 1 15 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=0.65
+ $Y=1.835 $X2=0.79 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_8%Y 1 2 3 4 5 6 7 8 9 10 11 12 39 41 42 45 47
+ 51 55 63 65 66 67 73 75 77 83 85 87 90 91 93 95 96 98 99 101 102 103 104 105
+ 113 119 123 128
c197 66 0 1.22355e-19 $X=5.245 $Y=1.17
r198 113 123 5.96046 $w=8.15e-07 $l=2.47386e-07 $layer=LI1_cond $X=4.065
+ $Y=1.347 $X2=4.08 $Y2=1.587
r199 105 128 12.8736 $w=8.15e-07 $l=8.6e-07 $layer=LI1_cond $X=4.23 $Y=1.587
+ $X2=5.09 $Y2=1.587
r200 105 123 0.523926 $w=8.15e-07 $l=3.5e-08 $layer=LI1_cond $X=4.115 $Y=1.587
+ $X2=4.08 $Y2=1.587
r201 105 119 39.0099 $w=2.18e-07 $l=7.4e-07 $layer=LI1_cond $X=4.23 $Y=1.21
+ $X2=4.23 $Y2=0.47
r202 105 113 1.46675 $w=2.73e-07 $l=3.5e-08 $layer=LI1_cond $X=4.03 $Y=1.347
+ $X2=4.065 $Y2=1.347
r203 104 105 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.347
+ $X2=4.03 $Y2=1.347
r204 95 103 6.49559 $w=2.73e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=1.347
+ $X2=3.12 $Y2=1.347
r205 95 96 3.75991 $w=2.75e-07 $l=9.5e-08 $layer=LI1_cond $X=3.275 $Y=1.347
+ $X2=3.37 $Y2=1.347
r206 94 104 5.65745 $w=2.73e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=1.347
+ $X2=3.6 $Y2=1.347
r207 94 96 3.75991 $w=2.75e-07 $l=9.5e-08 $layer=LI1_cond $X=3.465 $Y=1.347
+ $X2=3.37 $Y2=1.347
r208 92 103 21.5821 $w=2.73e-07 $l=5.15e-07 $layer=LI1_cond $X=2.605 $Y=1.347
+ $X2=3.12 $Y2=1.347
r209 92 93 4.52113 $w=2.22e-07 $l=3.54491e-07 $layer=LI1_cond $X=2.605 $Y=1.347
+ $X2=2.415 $Y2=1.075
r210 89 90 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.51 $Y=1.255
+ $X2=7.51 $Y2=1.92
r211 88 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=2.005
+ $X2=6.81 $Y2=2.005
r212 87 90 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.425 $Y=2.005
+ $X2=7.51 $Y2=1.92
r213 87 88 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.425 $Y=2.005
+ $X2=6.975 $Y2=2.005
r214 86 102 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.905 $Y=1.17
+ $X2=6.81 $Y2=1.17
r215 85 89 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.425 $Y=1.17
+ $X2=7.51 $Y2=1.255
r216 85 86 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.425 $Y=1.17
+ $X2=6.905 $Y2=1.17
r217 81 102 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.81 $Y=1.085
+ $X2=6.81 $Y2=1.17
r218 81 83 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=6.81 $Y=1.085
+ $X2=6.81 $Y2=0.47
r219 78 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=2.005
+ $X2=5.95 $Y2=2.005
r220 77 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=2.005
+ $X2=6.81 $Y2=2.005
r221 77 78 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.645 $Y=2.005
+ $X2=6.115 $Y2=2.005
r222 76 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.045 $Y=1.17
+ $X2=5.95 $Y2=1.17
r223 75 102 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.715 $Y=1.17
+ $X2=6.81 $Y2=1.17
r224 75 76 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.715 $Y=1.17
+ $X2=6.045 $Y2=1.17
r225 71 99 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=1.085
+ $X2=5.95 $Y2=1.17
r226 71 73 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=5.95 $Y=1.085
+ $X2=5.95 $Y2=0.47
r227 67 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=2.005
+ $X2=5.95 $Y2=2.005
r228 66 128 11.7564 $w=8.15e-07 $l=4.93654e-07 $layer=LI1_cond $X=5.255 $Y=2.005
+ $X2=5.09 $Y2=1.587
r229 66 67 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.255 $Y=2.005
+ $X2=5.785 $Y2=2.005
r230 65 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.855 $Y=1.17
+ $X2=5.95 $Y2=1.17
r231 65 66 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.855 $Y=1.17
+ $X2=5.245 $Y2=1.17
r232 61 128 9.59156 $w=1.9e-07 $l=5.02e-07 $layer=LI1_cond $X=5.09 $Y=1.085
+ $X2=5.09 $Y2=1.587
r233 61 63 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=5.09 $Y=1.085
+ $X2=5.09 $Y2=0.47
r234 53 96 2.70212 $w=1.9e-07 $l=1.37e-07 $layer=LI1_cond $X=3.37 $Y=1.21
+ $X2=3.37 $Y2=1.347
r235 53 55 43.1962 $w=1.88e-07 $l=7.4e-07 $layer=LI1_cond $X=3.37 $Y=1.21
+ $X2=3.37 $Y2=0.47
r236 49 93 1.91687 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=2.51 $Y=1.075
+ $X2=2.415 $Y2=1.075
r237 49 51 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=2.51 $Y=1.075
+ $X2=2.51 $Y2=0.47
r238 48 91 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.745 $Y=1.16
+ $X2=1.65 $Y2=1.16
r239 47 93 4.52113 $w=2.22e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=1.16
+ $X2=2.415 $Y2=1.075
r240 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.415 $Y=1.16
+ $X2=1.745 $Y2=1.16
r241 43 91 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=1.075
+ $X2=1.65 $Y2=1.16
r242 43 45 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=1.65 $Y=1.075
+ $X2=1.65 $Y2=0.48
r243 41 91 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.555 $Y=1.16
+ $X2=1.65 $Y2=1.16
r244 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.555 $Y=1.16
+ $X2=0.885 $Y2=1.16
r245 37 42 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.782 $Y=1.075
+ $X2=0.885 $Y2=1.16
r246 37 39 32.1907 $w=2.03e-07 $l=5.95e-07 $layer=LI1_cond $X=0.782 $Y=1.075
+ $X2=0.782 $Y2=0.48
r247 12 101 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=6.67
+ $Y=1.835 $X2=6.81 $Y2=2.04
r248 11 98 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=5.81
+ $Y=1.835 $X2=5.95 $Y2=2.04
r249 10 128 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.95
+ $Y=1.835 $X2=5.09 $Y2=1.98
r250 9 105 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.09
+ $Y=1.835 $X2=4.23 $Y2=1.98
r251 8 83 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.67
+ $Y=0.325 $X2=6.81 $Y2=0.47
r252 7 73 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.81
+ $Y=0.325 $X2=5.95 $Y2=0.47
r253 6 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.95
+ $Y=0.325 $X2=5.09 $Y2=0.47
r254 5 119 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.09
+ $Y=0.325 $X2=4.23 $Y2=0.47
r255 4 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.23
+ $Y=0.325 $X2=3.37 $Y2=0.47
r256 3 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.37
+ $Y=0.325 $X2=2.51 $Y2=0.47
r257 2 45 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.325 $X2=1.65 $Y2=0.48
r258 1 39 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.65
+ $Y=0.325 $X2=0.79 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_8%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 48
+ 52 56 60 64 67 68 69 70 72 73 74 75 76 77 79 84 96 110 115 118 121 124
r141 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r142 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r143 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r144 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r145 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r146 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r147 107 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r148 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r149 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r150 104 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r151 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r152 101 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=0
+ $X2=5.52 $Y2=0
r153 101 103 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.685 $Y=0 $X2=6
+ $Y2=0
r154 100 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r155 100 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r156 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r157 97 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=4.66 $Y2=0
r158 97 99 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=5.04 $Y2=0
r159 96 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=0
+ $X2=5.52 $Y2=0
r160 96 99 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.355 $Y=0
+ $X2=5.04 $Y2=0
r161 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r162 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r163 92 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r164 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r165 89 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.08 $Y2=0
r166 89 91 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.64 $Y2=0
r167 88 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r168 88 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r169 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r170 85 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=1.22 $Y2=0
r171 85 87 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r172 84 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=0
+ $X2=2.08 $Y2=0
r173 84 87 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=0
+ $X2=1.68 $Y2=0
r174 83 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r175 83 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r176 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r177 80 112 4.55932 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0
+ $X2=0.255 $Y2=0
r178 80 82 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.72
+ $Y2=0
r179 79 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=1.22 $Y2=0
r180 79 82 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r181 77 122 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.56 $Y2=0
r182 77 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r183 75 106 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.075 $Y=0
+ $X2=6.96 $Y2=0
r184 75 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.075 $Y=0 $X2=7.24
+ $Y2=0
r185 74 109 2.51176 $w=1.7e-07 $l=3.5e-08 $layer=LI1_cond $X=7.405 $Y=0 $X2=7.44
+ $Y2=0
r186 74 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.405 $Y=0 $X2=7.24
+ $Y2=0
r187 72 103 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.215 $Y=0 $X2=6
+ $Y2=0
r188 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.215 $Y=0 $X2=6.38
+ $Y2=0
r189 71 106 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.545 $Y=0
+ $X2=6.96 $Y2=0
r190 71 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.545 $Y=0 $X2=6.38
+ $Y2=0
r191 69 94 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.6
+ $Y2=0
r192 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.8
+ $Y2=0
r193 67 91 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=0
+ $X2=2.64 $Y2=0
r194 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.94
+ $Y2=0
r195 66 94 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.6
+ $Y2=0
r196 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=2.94
+ $Y2=0
r197 62 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0
r198 62 64 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=7.24 $Y=0.085
+ $X2=7.24 $Y2=0.47
r199 58 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.38 $Y=0.085
+ $X2=6.38 $Y2=0
r200 58 60 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=6.38 $Y=0.085
+ $X2=6.38 $Y2=0.47
r201 54 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.52 $Y2=0
r202 54 56 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.52 $Y2=0.47
r203 50 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.66 $Y2=0
r204 50 52 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.66 $Y2=0.47
r205 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=0 $X2=3.8
+ $Y2=0
r206 48 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=0
+ $X2=4.66 $Y2=0
r207 48 49 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.495 $Y=0
+ $X2=3.965 $Y2=0
r208 44 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=0.085 $X2=3.8
+ $Y2=0
r209 44 46 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.8 $Y=0.085
+ $X2=3.8 $Y2=0.47
r210 40 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0
r211 40 42 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0.47
r212 36 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0
r213 36 38 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0.45
r214 32 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r215 32 34 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.45
r216 28 112 3.1647 $w=3.25e-07 $l=1.27609e-07 $layer=LI1_cond $X=0.347 $Y=0.085
+ $X2=0.255 $Y2=0
r217 28 30 13.652 $w=3.23e-07 $l=3.85e-07 $layer=LI1_cond $X=0.347 $Y=0.085
+ $X2=0.347 $Y2=0.47
r218 9 64 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.1
+ $Y=0.325 $X2=7.24 $Y2=0.47
r219 8 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.24
+ $Y=0.325 $X2=6.38 $Y2=0.47
r220 7 56 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.38
+ $Y=0.325 $X2=5.52 $Y2=0.47
r221 6 52 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.52
+ $Y=0.325 $X2=4.66 $Y2=0.47
r222 5 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.66
+ $Y=0.325 $X2=3.8 $Y2=0.47
r223 4 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.8
+ $Y=0.325 $X2=2.94 $Y2=0.47
r224 3 38 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.94
+ $Y=0.325 $X2=2.08 $Y2=0.45
r225 2 34 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.08
+ $Y=0.325 $X2=1.22 $Y2=0.45
r226 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.225
+ $Y=0.325 $X2=0.35 $Y2=0.47
.ends

