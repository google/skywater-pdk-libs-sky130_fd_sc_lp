# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a2bb2oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a2bb2oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.805000 1.750000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.185000 1.385000 1.515000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.915000 1.210000 3.275000 1.760000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065000 1.200000 2.405000 1.750000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.569100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.450000 2.035000 2.745000 2.205000 ;
        RECT 1.450000 2.205000 1.775000 3.075000 ;
        RECT 1.950000 0.255000 2.150000 0.860000 ;
        RECT 1.950000 0.860000 2.745000 1.030000 ;
        RECT 2.575000 1.030000 2.745000 2.035000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.110000  0.085000 0.440000 1.040000 ;
      RECT 0.110000  1.920000 0.440000 3.245000 ;
      RECT 0.610000  0.255000 0.800000 0.845000 ;
      RECT 0.610000  0.845000 1.735000 1.015000 ;
      RECT 0.930000  1.920000 1.260000 3.075000 ;
      RECT 0.970000  0.085000 1.780000 0.675000 ;
      RECT 0.975000  1.695000 1.735000 1.865000 ;
      RECT 0.975000  1.865000 1.260000 1.920000 ;
      RECT 1.555000  1.015000 1.735000 1.200000 ;
      RECT 1.555000  1.200000 1.895000 1.515000 ;
      RECT 1.555000  1.515000 1.735000 1.695000 ;
      RECT 1.945000  2.375000 3.195000 2.545000 ;
      RECT 1.945000  2.545000 2.210000 3.075000 ;
      RECT 2.380000  2.715000 2.710000 3.245000 ;
      RECT 2.880000  2.545000 3.195000 3.075000 ;
      RECT 2.915000  1.930000 3.195000 2.375000 ;
      RECT 2.925000  0.085000 3.195000 1.040000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__a2bb2oi_1
END LIBRARY
