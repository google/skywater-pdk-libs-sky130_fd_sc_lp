* File: sky130_fd_sc_lp__einvn_8.spice
* Created: Fri Aug 28 10:33:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvn_8.pex.spice"
.subckt sky130_fd_sc_lp__einvn_8  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1023 N_A_110_57#_M1023_d N_TE_B_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_110_57#_M1004_g N_A_305_47#_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75006.6 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1004_d N_A_110_57#_M1012_g N_A_305_47#_M1012_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75006.2 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1014_d N_A_110_57#_M1014_g N_A_305_47#_M1012_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75005.8 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1014_d N_A_110_57#_M1016_g N_A_305_47#_M1016_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75005.3 A=0.126 P=1.98 MULT=1
MM1026 N_VGND_M1026_d N_A_110_57#_M1026_g N_A_305_47#_M1016_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75004.9 A=0.126 P=1.98 MULT=1
MM1027 N_VGND_M1026_d N_A_110_57#_M1027_g N_A_305_47#_M1027_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75004.5 A=0.126 P=1.98 MULT=1
MM1028 N_VGND_M1028_d N_A_110_57#_M1028_g N_A_305_47#_M1027_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1033 N_VGND_M1028_d N_A_110_57#_M1033_g N_A_305_47#_M1033_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1000 N_A_305_47#_M1033_s N_A_M1000_g N_Z_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1002 N_A_305_47#_M1002_d N_A_M1002_g N_Z_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.1
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1005 N_A_305_47#_M1002_d N_A_M1005_g N_Z_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.5
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1013 N_A_305_47#_M1013_d N_A_M1013_g N_Z_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.9
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1015 N_A_305_47#_M1013_d N_A_M1015_g N_Z_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.3
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1017 N_A_305_47#_M1017_d N_A_M1017_g N_Z_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.8
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1019 N_A_305_47#_M1017_d N_A_M1019_g N_Z_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1032 N_A_305_47#_M1032_d N_A_M1032_g N_Z_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_A_110_57#_M1010_d N_TE_B_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_TE_B_M1001_g N_A_305_367#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75006.6 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1001_d N_TE_B_M1006_g N_A_305_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75006.2 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_TE_B_M1011_g N_A_305_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75005.8 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1011_d N_TE_B_M1018_g N_A_305_367#_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75005.3 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_TE_B_M1022_g N_A_305_367#_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1024 N_VPWR_M1022_d N_TE_B_M1024_g N_A_305_367#_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1025_d N_TE_B_M1025_g N_A_305_367#_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1030 N_VPWR_M1025_d N_TE_B_M1030_g N_A_305_367#_M1030_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1003 N_A_305_367#_M1030_s N_A_M1003_g N_Z_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1007 N_A_305_367#_M1007_d N_A_M1007_g N_Z_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1008 N_A_305_367#_M1007_d N_A_M1008_g N_Z_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1009 N_A_305_367#_M1009_d N_A_M1009_g N_Z_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.9
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1020 N_A_305_367#_M1009_d N_A_M1020_g N_Z_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.3
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1021 N_A_305_367#_M1021_d N_A_M1021_g N_Z_M1020_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.8
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1029 N_A_305_367#_M1021_d N_A_M1029_g N_Z_M1029_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1031 N_A_305_367#_M1031_d N_A_M1031_g N_Z_M1029_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=17.7175 P=22.73
*
.include "sky130_fd_sc_lp__einvn_8.pxi.spice"
*
.ends
*
*
