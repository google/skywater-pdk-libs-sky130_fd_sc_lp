# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__mux4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.830000 1.175000 1.450000 2.175000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.155000 0.550000 2.175000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.400000 1.210000 5.880000 1.765000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.945000 1.080000 5.230000 1.765000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.990000 1.125000 3.650000 1.795000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.795000 1.355000 7.125000 1.865000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.725000 0.375000 9.995000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.095000  2.345000  1.735000 2.515000 ;
      RECT 0.095000  2.515000  0.355000 2.970000 ;
      RECT 0.125000  0.450000  0.385000 0.815000 ;
      RECT 0.125000  0.815000  1.225000 0.985000 ;
      RECT 0.525000  2.685000  0.855000 3.245000 ;
      RECT 0.555000  0.085000  0.885000 0.645000 ;
      RECT 1.025000  2.685000  1.285000 2.865000 ;
      RECT 1.025000  2.865000  2.665000 3.035000 ;
      RECT 1.055000  0.265000  2.225000 0.435000 ;
      RECT 1.055000  0.435000  1.225000 0.815000 ;
      RECT 1.395000  0.615000  1.725000 0.835000 ;
      RECT 1.395000  0.835000  2.075000 1.005000 ;
      RECT 1.475000  2.515000  1.735000 2.675000 ;
      RECT 1.895000  0.435000  2.225000 0.665000 ;
      RECT 1.905000  1.005000  2.075000 1.940000 ;
      RECT 1.905000  1.940000  2.305000 2.170000 ;
      RECT 1.905000  2.170000  2.235000 2.670000 ;
      RECT 2.255000  1.100000  2.820000 1.770000 ;
      RECT 2.405000  2.340000  2.665000 2.865000 ;
      RECT 2.560000  0.640000  2.820000 1.100000 ;
      RECT 2.650000  1.770000  2.820000 1.975000 ;
      RECT 2.650000  1.975000  4.435000 2.145000 ;
      RECT 2.885000  2.145000  3.175000 2.845000 ;
      RECT 2.990000  0.085000  3.320000 0.955000 ;
      RECT 3.345000  2.515000  3.645000 3.245000 ;
      RECT 3.510000  0.255000  5.220000 0.445000 ;
      RECT 3.510000  0.445000  3.805000 0.955000 ;
      RECT 3.955000  2.545000  4.205000 2.905000 ;
      RECT 3.955000  2.905000  5.115000 3.075000 ;
      RECT 3.975000  0.625000  4.200000 1.015000 ;
      RECT 3.975000  1.015000  4.775000 1.185000 ;
      RECT 4.175000  1.365000  4.435000 1.975000 ;
      RECT 4.370000  0.615000  4.700000 0.645000 ;
      RECT 4.370000  0.645000  6.160000 0.845000 ;
      RECT 4.385000  2.525000  4.775000 2.735000 ;
      RECT 4.605000  1.185000  4.775000 1.935000 ;
      RECT 4.605000  1.935000  6.615000 2.035000 ;
      RECT 4.605000  2.035000  7.600000 2.105000 ;
      RECT 4.605000  2.105000  4.775000 2.525000 ;
      RECT 4.890000  0.445000  5.220000 0.475000 ;
      RECT 4.945000  2.275000  6.005000 2.445000 ;
      RECT 4.945000  2.445000  5.115000 2.905000 ;
      RECT 5.285000  2.615000  5.535000 3.245000 ;
      RECT 5.390000  0.085000  5.720000 0.475000 ;
      RECT 5.705000  2.445000  6.005000 2.880000 ;
      RECT 5.890000  0.275000  6.160000 0.645000 ;
      RECT 6.225000  1.015000  7.250000 1.185000 ;
      RECT 6.225000  1.185000  6.555000 1.765000 ;
      RECT 6.410000  2.375000  6.750000 3.245000 ;
      RECT 6.445000  2.105000  7.600000 2.205000 ;
      RECT 6.490000  0.085000  6.820000 0.845000 ;
      RECT 6.920000  2.375000  7.250000 2.780000 ;
      RECT 6.920000  2.780000  7.650000 3.075000 ;
      RECT 7.000000  0.640000  7.250000 1.015000 ;
      RECT 7.430000  0.790000  7.710000 1.120000 ;
      RECT 7.430000  1.120000  7.600000 2.035000 ;
      RECT 7.430000  2.205000  7.600000 2.380000 ;
      RECT 7.430000  2.380000  8.850000 2.610000 ;
      RECT 7.780000  1.880000  8.050000 2.210000 ;
      RECT 7.880000  0.390000  8.910000 0.620000 ;
      RECT 7.880000  0.620000  8.050000 1.880000 ;
      RECT 8.220000  0.790000  8.445000 1.345000 ;
      RECT 8.220000  1.345000  9.555000 1.675000 ;
      RECT 8.220000  1.675000  8.440000 2.210000 ;
      RECT 8.610000  1.880000  8.850000 2.380000 ;
      RECT 8.615000  0.620000  8.910000 1.120000 ;
      RECT 9.225000  0.085000  9.555000 1.175000 ;
      RECT 9.225000  1.845000  9.555000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  1.950000 2.245000 2.120000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  1.950000 8.005000 2.120000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
    LAYER met1 ;
      RECT 2.015000 1.920000 2.305000 1.965000 ;
      RECT 2.015000 1.965000 8.065000 2.105000 ;
      RECT 2.015000 2.105000 2.305000 2.150000 ;
      RECT 7.775000 1.920000 8.065000 1.965000 ;
      RECT 7.775000 2.105000 8.065000 2.150000 ;
  END
END sky130_fd_sc_lp__mux4_1
END LIBRARY
