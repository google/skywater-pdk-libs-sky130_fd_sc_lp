# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a2bb2o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a2bb2o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 0.370000 1.295000 2.155000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.015000 1.925000 1.525000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.840000 3.755000 2.225000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.915000 0.280000 3.215000 2.225000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.255000 0.505000 1.095000 ;
        RECT 0.105000 1.095000 0.285000 1.815000 ;
        RECT 0.105000 1.815000 0.565000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.455000  1.345000 0.925000 1.645000 ;
      RECT 0.675000  0.085000 0.935000 1.095000 ;
      RECT 0.735000  2.665000 1.065000 3.245000 ;
      RECT 0.755000  1.645000 0.925000 2.325000 ;
      RECT 0.755000  2.325000 2.365000 2.495000 ;
      RECT 1.465000  0.280000 1.715000 0.665000 ;
      RECT 1.465000  0.665000 2.280000 0.835000 ;
      RECT 1.780000  1.705000 2.385000 1.875000 ;
      RECT 1.780000  1.875000 1.990000 2.145000 ;
      RECT 1.890000  0.085000 2.220000 0.495000 ;
      RECT 2.070000  2.495000 2.365000 3.020000 ;
      RECT 2.110000  0.835000 2.280000 1.005000 ;
      RECT 2.110000  1.005000 2.385000 1.705000 ;
      RECT 2.170000  2.055000 2.735000 2.225000 ;
      RECT 2.170000  2.225000 2.365000 2.325000 ;
      RECT 2.450000  0.280000 2.735000 0.675000 ;
      RECT 2.535000  2.395000 3.690000 2.565000 ;
      RECT 2.535000  2.565000 2.760000 3.020000 ;
      RECT 2.565000  0.675000 2.735000 2.055000 ;
      RECT 2.930000  2.735000 3.260000 3.245000 ;
      RECT 3.385000  0.085000 3.655000 0.610000 ;
      RECT 3.430000  2.565000 3.690000 3.020000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__a2bb2o_1
END LIBRARY
