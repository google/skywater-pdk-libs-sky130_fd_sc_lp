* File: sky130_fd_sc_lp__o21a_4.pxi.spice
* Created: Wed Sep  2 10:15:27 2020
* 
x_PM_SKY130_FD_SC_LP__O21A_4%A_90_23# N_A_90_23#_M1007_d N_A_90_23#_M1008_s
+ N_A_90_23#_M1006_s N_A_90_23#_M1001_g N_A_90_23#_M1002_g N_A_90_23#_M1003_g
+ N_A_90_23#_M1009_g N_A_90_23#_M1004_g N_A_90_23#_M1012_g N_A_90_23#_M1010_g
+ N_A_90_23#_M1018_g N_A_90_23#_c_193_p N_A_90_23#_c_102_n N_A_90_23#_c_103_n
+ N_A_90_23#_c_104_n N_A_90_23#_c_105_n N_A_90_23#_c_119_p N_A_90_23#_c_169_p
+ N_A_90_23#_c_131_p N_A_90_23#_c_184_p N_A_90_23#_c_122_p N_A_90_23#_c_106_n
+ N_A_90_23#_c_107_n N_A_90_23#_c_145_p N_A_90_23#_c_147_p N_A_90_23#_c_108_n
+ N_A_90_23#_c_109_n N_A_90_23#_c_110_n PM_SKY130_FD_SC_LP__O21A_4%A_90_23#
x_PM_SKY130_FD_SC_LP__O21A_4%B1 N_B1_M1008_g N_B1_M1007_g N_B1_M1017_g
+ N_B1_M1013_g B1 N_B1_c_256_n N_B1_c_253_n PM_SKY130_FD_SC_LP__O21A_4%B1
x_PM_SKY130_FD_SC_LP__O21A_4%A1 N_A1_M1016_g N_A1_M1000_g N_A1_M1019_g
+ N_A1_M1015_g N_A1_c_315_n N_A1_c_316_n N_A1_c_309_n N_A1_c_310_n N_A1_c_311_n
+ N_A1_c_318_n N_A1_c_312_n N_A1_c_358_p A1 A1 A1 PM_SKY130_FD_SC_LP__O21A_4%A1
x_PM_SKY130_FD_SC_LP__O21A_4%A2 N_A2_M1005_g N_A2_M1006_g N_A2_M1011_g
+ N_A2_M1014_g A2 N_A2_c_400_n N_A2_c_397_n PM_SKY130_FD_SC_LP__O21A_4%A2
x_PM_SKY130_FD_SC_LP__O21A_4%VPWR N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_M1018_d
+ N_VPWR_M1017_d N_VPWR_M1015_s N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_457_n
+ N_VPWR_c_497_n N_VPWR_c_458_n N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n
+ N_VPWR_c_462_n N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n VPWR
+ N_VPWR_c_466_n N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_454_n
+ PM_SKY130_FD_SC_LP__O21A_4%VPWR
x_PM_SKY130_FD_SC_LP__O21A_4%X N_X_M1001_d N_X_M1004_d N_X_M1002_s N_X_M1012_s
+ N_X_c_543_n N_X_c_548_n N_X_c_549_n N_X_c_593_p N_X_c_544_n N_X_c_581_n
+ N_X_c_550_n N_X_c_594_p N_X_c_585_n N_X_c_545_n N_X_c_551_n X X N_X_c_546_n X
+ PM_SKY130_FD_SC_LP__O21A_4%X
x_PM_SKY130_FD_SC_LP__O21A_4%A_792_367# N_A_792_367#_M1000_d
+ N_A_792_367#_M1014_d N_A_792_367#_c_601_n
+ PM_SKY130_FD_SC_LP__O21A_4%A_792_367#
x_PM_SKY130_FD_SC_LP__O21A_4%VGND N_VGND_M1001_s N_VGND_M1003_s N_VGND_M1010_s
+ N_VGND_M1016_s N_VGND_M1011_s N_VGND_c_613_n N_VGND_c_614_n N_VGND_c_615_n
+ N_VGND_c_616_n N_VGND_c_617_n N_VGND_c_618_n VGND N_VGND_c_619_n
+ N_VGND_c_620_n N_VGND_c_621_n N_VGND_c_622_n N_VGND_c_623_n N_VGND_c_624_n
+ N_VGND_c_625_n N_VGND_c_626_n N_VGND_c_627_n N_VGND_c_628_n
+ PM_SKY130_FD_SC_LP__O21A_4%VGND
x_PM_SKY130_FD_SC_LP__O21A_4%A_485_65# N_A_485_65#_M1007_s N_A_485_65#_M1013_s
+ N_A_485_65#_M1005_d N_A_485_65#_M1019_d N_A_485_65#_c_701_n
+ N_A_485_65#_c_702_n N_A_485_65#_c_703_n N_A_485_65#_c_723_n
+ N_A_485_65#_c_716_n N_A_485_65#_c_717_n N_A_485_65#_c_704_n
+ N_A_485_65#_c_705_n N_A_485_65#_c_706_n N_A_485_65#_c_707_n
+ PM_SKY130_FD_SC_LP__O21A_4%A_485_65#
cc_1 VNB N_A_90_23#_M1001_g 0.0258995f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.665
cc_2 VNB N_A_90_23#_M1003_g 0.0213923f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=0.665
cc_3 VNB N_A_90_23#_M1004_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=0.665
cc_4 VNB N_A_90_23#_M1010_g 0.0261293f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=0.665
cc_5 VNB N_A_90_23#_c_102_n 0.00250178f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.395
cc_6 VNB N_A_90_23#_c_103_n 4.09436e-19 $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.93
cc_7 VNB N_A_90_23#_c_104_n 0.0101734f $X=-0.19 $Y=-0.245 $X2=2.915 $Y2=1.16
cc_8 VNB N_A_90_23#_c_105_n 0.00844715f $X=-0.19 $Y=-0.245 $X2=2.345 $Y2=1.16
cc_9 VNB N_A_90_23#_c_106_n 0.0131278f $X=-0.19 $Y=-0.245 $X2=4.085 $Y2=1.16
cc_10 VNB N_A_90_23#_c_107_n 0.00309185f $X=-0.19 $Y=-0.245 $X2=4.175 $Y2=1.93
cc_11 VNB N_A_90_23#_c_108_n 0.00131117f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.49
cc_12 VNB N_A_90_23#_c_109_n 0.00341299f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.16
cc_13 VNB N_A_90_23#_c_110_n 0.091678f $X=-0.19 $Y=-0.245 $X2=2.135 $Y2=1.49
cc_14 VNB N_B1_M1007_g 0.0234455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_M1013_g 0.0202086f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.465
cc_16 VNB N_B1_c_253_n 0.0503038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_M1016_g 0.02165f $X=-0.19 $Y=-0.245 $X2=4.39 $Y2=1.835
cc_18 VNB N_A1_M1019_g 0.0261593f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.665
cc_19 VNB N_A1_c_309_n 0.0026956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_310_n 0.00849916f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=2.465
cc_21 VNB N_A1_c_311_n 0.0305967f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=2.465
cc_22 VNB N_A1_c_312_n 0.029017f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=0.665
cc_23 VNB N_A2_M1005_g 0.0200025f $X=-0.19 $Y=-0.245 $X2=4.39 $Y2=1.835
cc_24 VNB N_A2_M1011_g 0.0192547f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.665
cc_25 VNB N_A2_c_397_n 0.0316427f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=2.465
cc_26 VNB N_VPWR_c_454_n 0.243291f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=1.49
cc_27 VNB N_X_c_543_n 0.00169931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_544_n 0.00594953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_545_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=2.175 $Y2=1.49
cc_30 VNB N_X_c_546_n 0.0108425f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.49
cc_31 VNB X 0.0225881f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.395
cc_32 VNB N_VGND_c_613_n 0.0120364f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.465
cc_33 VNB N_VGND_c_614_n 0.0281524f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.325
cc_34 VNB N_VGND_c_615_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.655
cc_35 VNB N_VGND_c_616_n 0.00985637f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=1.325
cc_36 VNB N_VGND_c_617_n 0.00453441f $X=-0.19 $Y=-0.245 $X2=1.705 $Y2=1.655
cc_37 VNB N_VGND_c_618_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=1.325
cc_38 VNB N_VGND_c_619_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=2.135 $Y2=1.655
cc_39 VNB N_VGND_c_620_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.49
cc_40 VNB N_VGND_c_621_n 0.0413769f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=1.49
cc_41 VNB N_VGND_c_622_n 0.0136617f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.93
cc_42 VNB N_VGND_c_623_n 0.0196948f $X=-0.19 $Y=-0.245 $X2=2.78 $Y2=2.91
cc_43 VNB N_VGND_c_624_n 0.318433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_625_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=1.16
cc_45 VNB N_VGND_c_626_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=4.265 $Y2=2.035
cc_46 VNB N_VGND_c_627_n 0.0059779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_628_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=2.78 $Y2=2.095
cc_48 VNB N_A_485_65#_c_701_n 0.00398509f $X=-0.19 $Y=-0.245 $X2=0.845 $Y2=2.465
cc_49 VNB N_A_485_65#_c_702_n 0.00490999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_485_65#_c_703_n 0.00429866f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.325
cc_51 VNB N_A_485_65#_c_704_n 0.00184018f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=0.665
cc_52 VNB N_A_485_65#_c_705_n 0.0168011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_485_65#_c_706_n 0.00217937f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=1.325
cc_54 VNB N_A_485_65#_c_707_n 0.0316355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VPB N_A_90_23#_M1002_g 0.0229319f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.465
cc_56 VPB N_A_90_23#_M1009_g 0.0188632f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=2.465
cc_57 VPB N_A_90_23#_M1012_g 0.0188554f $X=-0.19 $Y=1.655 $X2=1.705 $Y2=2.465
cc_58 VPB N_A_90_23#_M1018_g 0.0187977f $X=-0.19 $Y=1.655 $X2=2.135 $Y2=2.465
cc_59 VPB N_A_90_23#_c_103_n 0.001335f $X=-0.19 $Y=1.655 $X2=2.26 $Y2=1.93
cc_60 VPB N_A_90_23#_c_107_n 0.00106287f $X=-0.19 $Y=1.655 $X2=4.175 $Y2=1.93
cc_61 VPB N_A_90_23#_c_110_n 0.0153801f $X=-0.19 $Y=1.655 $X2=2.135 $Y2=1.49
cc_62 VPB N_B1_M1008_g 0.0184362f $X=-0.19 $Y=1.655 $X2=4.39 $Y2=1.835
cc_63 VPB N_B1_M1017_g 0.0222091f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.665
cc_64 VPB N_B1_c_256_n 0.00919001f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=0.665
cc_65 VPB N_B1_c_253_n 0.0155346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A1_M1000_g 0.0226812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A1_M1015_g 0.0249717f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.465
cc_68 VPB N_A1_c_315_n 0.00214513f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=1.325
cc_69 VPB N_A1_c_316_n 0.00133672f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=0.665
cc_70 VPB N_A1_c_311_n 0.00752084f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=2.465
cc_71 VPB N_A1_c_318_n 0.00573302f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=0.665
cc_72 VPB N_A1_c_312_n 0.00792246f $X=-0.19 $Y=1.655 $X2=1.385 $Y2=0.665
cc_73 VPB N_A2_M1006_g 0.0181036f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A2_M1014_g 0.018668f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.465
cc_75 VPB N_A2_c_400_n 0.00258442f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=2.465
cc_76 VPB N_A2_c_397_n 0.00474859f $X=-0.19 $Y=1.655 $X2=1.275 $Y2=2.465
cc_77 VPB N_VPWR_c_455_n 0.0414999f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=1.325
cc_78 VPB N_VPWR_c_456_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.275 $Y2=2.465
cc_79 VPB N_VPWR_c_457_n 3.08929e-19 $X=-0.19 $Y=1.655 $X2=1.705 $Y2=1.655
cc_80 VPB N_VPWR_c_458_n 0.0137153f $X=-0.19 $Y=1.655 $X2=2.135 $Y2=1.655
cc_81 VPB N_VPWR_c_459_n 0.0561341f $X=-0.19 $Y=1.655 $X2=2.135 $Y2=2.465
cc_82 VPB N_VPWR_c_460_n 0.0169405f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.49
cc_83 VPB N_VPWR_c_461_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_462_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.045 $Y2=1.49
cc_85 VPB N_VPWR_c_463_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.045 $Y2=1.49
cc_86 VPB N_VPWR_c_464_n 0.0130339f $X=-0.19 $Y=1.655 $X2=2.26 $Y2=1.245
cc_87 VPB N_VPWR_c_465_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.26 $Y2=1.395
cc_88 VPB N_VPWR_c_466_n 0.0373044f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=0.68
cc_89 VPB N_VPWR_c_467_n 0.0129339f $X=-0.19 $Y=1.655 $X2=2.78 $Y2=2.015
cc_90 VPB N_VPWR_c_468_n 0.0149951f $X=-0.19 $Y=1.655 $X2=0.955 $Y2=1.49
cc_91 VPB N_VPWR_c_454_n 0.0637786f $X=-0.19 $Y=1.655 $X2=1.705 $Y2=1.49
cc_92 VPB N_X_c_548_n 0.00914439f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.465
cc_93 VPB N_X_c_549_n 0.0192979f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=2.465
cc_94 VPB N_X_c_550_n 0.00495564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_X_c_551_n 0.00144314f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.49
cc_96 VPB X 0.00576796f $X=-0.19 $Y=1.655 $X2=2.26 $Y2=1.395
cc_97 N_A_90_23#_M1018_g N_B1_M1008_g 0.0252333f $X=2.135 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_90_23#_c_119_p N_B1_M1008_g 0.0128856f $X=2.685 $Y=2.015 $X2=0 $Y2=0
cc_99 N_A_90_23#_c_102_n N_B1_M1007_g 0.00236876f $X=2.26 $Y=1.395 $X2=0 $Y2=0
cc_100 N_A_90_23#_c_104_n N_B1_M1007_g 0.0111609f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_90_23#_c_122_p N_B1_M1007_g 0.0112814f $X=3.08 $Y=0.68 $X2=0 $Y2=0
cc_102 N_A_90_23#_c_109_n N_B1_M1007_g 0.00169298f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_90_23#_c_110_n N_B1_M1007_g 2.84209e-19 $X=2.135 $Y=1.49 $X2=0 $Y2=0
cc_104 N_A_90_23#_c_122_p N_B1_M1013_g 0.00685613f $X=3.08 $Y=0.68 $X2=0 $Y2=0
cc_105 N_A_90_23#_c_106_n N_B1_M1013_g 0.0129877f $X=4.085 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_90_23#_c_109_n N_B1_M1013_g 0.00248676f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_90_23#_c_103_n N_B1_c_256_n 0.0138086f $X=2.26 $Y=1.93 $X2=0 $Y2=0
cc_108 N_A_90_23#_c_104_n N_B1_c_256_n 0.0283218f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_90_23#_c_119_p N_B1_c_256_n 0.0107813f $X=2.685 $Y=2.015 $X2=0 $Y2=0
cc_110 N_A_90_23#_c_131_p N_B1_c_256_n 0.0154121f $X=2.78 $Y=2.1 $X2=0 $Y2=0
cc_111 N_A_90_23#_c_108_n N_B1_c_256_n 0.0141599f $X=2.26 $Y=1.49 $X2=0 $Y2=0
cc_112 N_A_90_23#_c_109_n N_B1_c_256_n 0.0216405f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_90_23#_c_110_n N_B1_c_256_n 3.21781e-19 $X=2.135 $Y=1.49 $X2=0 $Y2=0
cc_114 N_A_90_23#_c_102_n N_B1_c_253_n 0.00112381f $X=2.26 $Y=1.395 $X2=0 $Y2=0
cc_115 N_A_90_23#_c_103_n N_B1_c_253_n 0.00476809f $X=2.26 $Y=1.93 $X2=0 $Y2=0
cc_116 N_A_90_23#_c_104_n N_B1_c_253_n 0.00876853f $X=2.915 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_90_23#_c_131_p N_B1_c_253_n 6.34959e-19 $X=2.78 $Y=2.1 $X2=0 $Y2=0
cc_118 N_A_90_23#_c_108_n N_B1_c_253_n 0.00223236f $X=2.26 $Y=1.49 $X2=0 $Y2=0
cc_119 N_A_90_23#_c_109_n N_B1_c_253_n 0.00271691f $X=3.08 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_90_23#_c_110_n N_B1_c_253_n 0.0252333f $X=2.135 $Y=1.49 $X2=0 $Y2=0
cc_121 N_A_90_23#_c_122_p N_A1_M1016_g 5.37284e-19 $X=3.08 $Y=0.68 $X2=0 $Y2=0
cc_122 N_A_90_23#_c_106_n N_A1_M1016_g 0.0113094f $X=4.085 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_90_23#_c_107_n N_A1_M1016_g 0.00206085f $X=4.175 $Y=1.93 $X2=0 $Y2=0
cc_124 N_A_90_23#_c_145_p N_A1_M1000_g 0.00144304f $X=4.265 $Y=2.035 $X2=0 $Y2=0
cc_125 N_A_90_23#_c_145_p N_A1_c_315_n 0.0164262f $X=4.265 $Y=2.035 $X2=0 $Y2=0
cc_126 N_A_90_23#_c_147_p N_A1_c_316_n 0.0116655f $X=4.53 $Y=2.035 $X2=0 $Y2=0
cc_127 N_A_90_23#_c_106_n N_A1_c_318_n 0.0236262f $X=4.085 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_90_23#_c_107_n N_A1_c_318_n 0.0369946f $X=4.175 $Y=1.93 $X2=0 $Y2=0
cc_129 N_A_90_23#_c_106_n N_A1_c_312_n 0.00660213f $X=4.085 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A_90_23#_c_107_n N_A1_c_312_n 0.00511448f $X=4.175 $Y=1.93 $X2=0 $Y2=0
cc_131 N_A_90_23#_M1006_s A1 0.0034413f $X=4.39 $Y=1.835 $X2=0 $Y2=0
cc_132 N_A_90_23#_c_145_p A1 0.00986534f $X=4.265 $Y=2.035 $X2=0 $Y2=0
cc_133 N_A_90_23#_c_147_p A1 0.0226703f $X=4.53 $Y=2.035 $X2=0 $Y2=0
cc_134 N_A_90_23#_c_106_n N_A2_M1005_g 0.00449426f $X=4.085 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_90_23#_c_107_n N_A2_M1005_g 0.00252571f $X=4.175 $Y=1.93 $X2=0 $Y2=0
cc_136 N_A_90_23#_c_107_n N_A2_M1006_g 0.0056656f $X=4.175 $Y=1.93 $X2=0 $Y2=0
cc_137 N_A_90_23#_c_145_p N_A2_M1006_g 0.00242641f $X=4.265 $Y=2.035 $X2=0 $Y2=0
cc_138 N_A_90_23#_c_147_p N_A2_M1006_g 0.00968336f $X=4.53 $Y=2.035 $X2=0 $Y2=0
cc_139 N_A_90_23#_c_107_n N_A2_M1011_g 4.46533e-19 $X=4.175 $Y=1.93 $X2=0 $Y2=0
cc_140 N_A_90_23#_c_107_n N_A2_M1014_g 7.02472e-19 $X=4.175 $Y=1.93 $X2=0 $Y2=0
cc_141 N_A_90_23#_c_147_p N_A2_M1014_g 0.00320127f $X=4.53 $Y=2.035 $X2=0 $Y2=0
cc_142 N_A_90_23#_c_107_n N_A2_c_400_n 0.0232646f $X=4.175 $Y=1.93 $X2=0 $Y2=0
cc_143 N_A_90_23#_c_147_p N_A2_c_400_n 0.0174347f $X=4.53 $Y=2.035 $X2=0 $Y2=0
cc_144 N_A_90_23#_c_107_n N_A2_c_397_n 0.0101549f $X=4.175 $Y=1.93 $X2=0 $Y2=0
cc_145 N_A_90_23#_c_147_p N_A2_c_397_n 5.72878e-19 $X=4.53 $Y=2.035 $X2=0 $Y2=0
cc_146 N_A_90_23#_c_103_n N_VPWR_M1018_d 0.00107328f $X=2.26 $Y=1.93 $X2=0 $Y2=0
cc_147 N_A_90_23#_c_119_p N_VPWR_M1018_d 0.00424436f $X=2.685 $Y=2.015 $X2=0
+ $Y2=0
cc_148 N_A_90_23#_c_169_p N_VPWR_M1018_d 8.52101e-19 $X=2.345 $Y=2.015 $X2=0
+ $Y2=0
cc_149 N_A_90_23#_M1002_g N_VPWR_c_455_n 0.0152824f $X=0.845 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_90_23#_M1009_g N_VPWR_c_455_n 7.27171e-19 $X=1.275 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_90_23#_M1002_g N_VPWR_c_456_n 7.27171e-19 $X=0.845 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_90_23#_M1009_g N_VPWR_c_456_n 0.0142189f $X=1.275 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A_90_23#_M1012_g N_VPWR_c_456_n 0.0142189f $X=1.705 $Y=2.465 $X2=0
+ $Y2=0
cc_154 N_A_90_23#_M1018_g N_VPWR_c_456_n 7.27171e-19 $X=2.135 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_90_23#_M1012_g N_VPWR_c_457_n 6.90148e-19 $X=1.705 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_90_23#_M1018_g N_VPWR_c_457_n 0.0147158f $X=2.135 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_90_23#_c_119_p N_VPWR_c_457_n 0.00890916f $X=2.685 $Y=2.015 $X2=0
+ $Y2=0
cc_158 N_A_90_23#_c_169_p N_VPWR_c_457_n 0.00897683f $X=2.345 $Y=2.015 $X2=0
+ $Y2=0
cc_159 N_A_90_23#_M1002_g N_VPWR_c_462_n 0.00486043f $X=0.845 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_90_23#_M1009_g N_VPWR_c_462_n 0.00486043f $X=1.275 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_90_23#_M1012_g N_VPWR_c_464_n 0.00486043f $X=1.705 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_90_23#_M1018_g N_VPWR_c_464_n 0.00486043f $X=2.135 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_90_23#_c_184_p N_VPWR_c_467_n 0.0124525f $X=2.78 $Y=2.91 $X2=0 $Y2=0
cc_164 N_A_90_23#_M1008_s N_VPWR_c_454_n 0.00536646f $X=2.64 $Y=1.835 $X2=0
+ $Y2=0
cc_165 N_A_90_23#_M1006_s N_VPWR_c_454_n 0.00231436f $X=4.39 $Y=1.835 $X2=0
+ $Y2=0
cc_166 N_A_90_23#_M1002_g N_VPWR_c_454_n 0.00824727f $X=0.845 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_90_23#_M1009_g N_VPWR_c_454_n 0.00824727f $X=1.275 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_90_23#_M1012_g N_VPWR_c_454_n 0.00824727f $X=1.705 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_90_23#_M1018_g N_VPWR_c_454_n 0.00824727f $X=2.135 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_90_23#_c_184_p N_VPWR_c_454_n 0.00730901f $X=2.78 $Y=2.91 $X2=0 $Y2=0
cc_171 N_A_90_23#_M1001_g N_X_c_543_n 0.0160841f $X=0.525 $Y=0.665 $X2=0 $Y2=0
cc_172 N_A_90_23#_c_193_p N_X_c_543_n 0.00867724f $X=2.175 $Y=1.49 $X2=0 $Y2=0
cc_173 N_A_90_23#_M1002_g N_X_c_548_n 0.015192f $X=0.845 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_90_23#_c_193_p N_X_c_548_n 0.0314885f $X=2.175 $Y=1.49 $X2=0 $Y2=0
cc_175 N_A_90_23#_c_110_n N_X_c_548_n 0.00911053f $X=2.135 $Y=1.49 $X2=0 $Y2=0
cc_176 N_A_90_23#_M1003_g N_X_c_544_n 0.0138332f $X=0.955 $Y=0.665 $X2=0 $Y2=0
cc_177 N_A_90_23#_M1004_g N_X_c_544_n 0.0135652f $X=1.385 $Y=0.665 $X2=0 $Y2=0
cc_178 N_A_90_23#_M1010_g N_X_c_544_n 0.00195123f $X=1.815 $Y=0.665 $X2=0 $Y2=0
cc_179 N_A_90_23#_c_193_p N_X_c_544_n 0.0625611f $X=2.175 $Y=1.49 $X2=0 $Y2=0
cc_180 N_A_90_23#_c_105_n N_X_c_544_n 0.00652734f $X=2.345 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_90_23#_c_110_n N_X_c_544_n 0.00582235f $X=2.135 $Y=1.49 $X2=0 $Y2=0
cc_182 N_A_90_23#_M1009_g N_X_c_550_n 0.0131657f $X=1.275 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_90_23#_M1012_g N_X_c_550_n 0.0129884f $X=1.705 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_90_23#_M1018_g N_X_c_550_n 6.42323e-19 $X=2.135 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_90_23#_c_193_p N_X_c_550_n 0.0617482f $X=2.175 $Y=1.49 $X2=0 $Y2=0
cc_186 N_A_90_23#_c_103_n N_X_c_550_n 0.00947169f $X=2.26 $Y=1.93 $X2=0 $Y2=0
cc_187 N_A_90_23#_c_110_n N_X_c_550_n 0.00548187f $X=2.135 $Y=1.49 $X2=0 $Y2=0
cc_188 N_A_90_23#_c_193_p N_X_c_545_n 0.0154426f $X=2.175 $Y=1.49 $X2=0 $Y2=0
cc_189 N_A_90_23#_c_110_n N_X_c_545_n 0.00262131f $X=2.135 $Y=1.49 $X2=0 $Y2=0
cc_190 N_A_90_23#_c_193_p N_X_c_551_n 0.0154426f $X=2.175 $Y=1.49 $X2=0 $Y2=0
cc_191 N_A_90_23#_c_110_n N_X_c_551_n 0.00296179f $X=2.135 $Y=1.49 $X2=0 $Y2=0
cc_192 N_A_90_23#_M1001_g X 0.0159287f $X=0.525 $Y=0.665 $X2=0 $Y2=0
cc_193 N_A_90_23#_M1002_g X 0.00274444f $X=0.845 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A_90_23#_c_193_p X 0.0155181f $X=2.175 $Y=1.49 $X2=0 $Y2=0
cc_195 N_A_90_23#_c_107_n N_A_792_367#_M1000_d 7.44237e-19 $X=4.175 $Y=1.93
+ $X2=-0.19 $Y2=-0.245
cc_196 N_A_90_23#_c_145_p N_A_792_367#_M1000_d 0.00285755f $X=4.265 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_197 N_A_90_23#_M1006_s N_A_792_367#_c_601_n 0.00366227f $X=4.39 $Y=1.835
+ $X2=0 $Y2=0
cc_198 N_A_90_23#_c_106_n N_VGND_M1016_s 0.00265361f $X=4.085 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_90_23#_M1001_g N_VGND_c_614_n 0.0120262f $X=0.525 $Y=0.665 $X2=0
+ $Y2=0
cc_200 N_A_90_23#_M1003_g N_VGND_c_614_n 6.10117e-19 $X=0.955 $Y=0.665 $X2=0
+ $Y2=0
cc_201 N_A_90_23#_M1001_g N_VGND_c_615_n 6.10117e-19 $X=0.525 $Y=0.665 $X2=0
+ $Y2=0
cc_202 N_A_90_23#_M1003_g N_VGND_c_615_n 0.0110386f $X=0.955 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_90_23#_M1004_g N_VGND_c_615_n 0.0110386f $X=1.385 $Y=0.665 $X2=0
+ $Y2=0
cc_204 N_A_90_23#_M1010_g N_VGND_c_615_n 6.10117e-19 $X=1.815 $Y=0.665 $X2=0
+ $Y2=0
cc_205 N_A_90_23#_M1004_g N_VGND_c_616_n 6.15775e-19 $X=1.385 $Y=0.665 $X2=0
+ $Y2=0
cc_206 N_A_90_23#_M1010_g N_VGND_c_616_n 0.0129f $X=1.815 $Y=0.665 $X2=0 $Y2=0
cc_207 N_A_90_23#_c_193_p N_VGND_c_616_n 0.00959752f $X=2.175 $Y=1.49 $X2=0
+ $Y2=0
cc_208 N_A_90_23#_c_105_n N_VGND_c_616_n 0.00178022f $X=2.345 $Y=1.16 $X2=0
+ $Y2=0
cc_209 N_A_90_23#_c_110_n N_VGND_c_616_n 0.00628361f $X=2.135 $Y=1.49 $X2=0
+ $Y2=0
cc_210 N_A_90_23#_M1001_g N_VGND_c_619_n 0.00477554f $X=0.525 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_90_23#_M1003_g N_VGND_c_619_n 0.00477554f $X=0.955 $Y=0.665 $X2=0
+ $Y2=0
cc_212 N_A_90_23#_M1004_g N_VGND_c_620_n 0.00477554f $X=1.385 $Y=0.665 $X2=0
+ $Y2=0
cc_213 N_A_90_23#_M1010_g N_VGND_c_620_n 0.00477554f $X=1.815 $Y=0.665 $X2=0
+ $Y2=0
cc_214 N_A_90_23#_M1001_g N_VGND_c_624_n 0.00825815f $X=0.525 $Y=0.665 $X2=0
+ $Y2=0
cc_215 N_A_90_23#_M1003_g N_VGND_c_624_n 0.00825815f $X=0.955 $Y=0.665 $X2=0
+ $Y2=0
cc_216 N_A_90_23#_M1004_g N_VGND_c_624_n 0.00825815f $X=1.385 $Y=0.665 $X2=0
+ $Y2=0
cc_217 N_A_90_23#_M1010_g N_VGND_c_624_n 0.00825815f $X=1.815 $Y=0.665 $X2=0
+ $Y2=0
cc_218 N_A_90_23#_c_104_n N_A_485_65#_M1007_s 0.00426494f $X=2.915 $Y=1.16
+ $X2=-0.19 $Y2=-0.245
cc_219 N_A_90_23#_c_106_n N_A_485_65#_M1013_s 0.00261503f $X=4.085 $Y=1.16 $X2=0
+ $Y2=0
cc_220 N_A_90_23#_M1010_g N_A_485_65#_c_701_n 8.83534e-19 $X=1.815 $Y=0.665
+ $X2=0 $Y2=0
cc_221 N_A_90_23#_c_104_n N_A_485_65#_c_701_n 0.0246174f $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_222 N_A_90_23#_M1007_d N_A_485_65#_c_702_n 0.00176461f $X=2.94 $Y=0.325 $X2=0
+ $Y2=0
cc_223 N_A_90_23#_c_104_n N_A_485_65#_c_702_n 0.00275981f $X=2.915 $Y=1.16 $X2=0
+ $Y2=0
cc_224 N_A_90_23#_c_122_p N_A_485_65#_c_702_n 0.0159249f $X=3.08 $Y=0.68 $X2=0
+ $Y2=0
cc_225 N_A_90_23#_c_106_n N_A_485_65#_c_702_n 0.00275981f $X=4.085 $Y=1.16 $X2=0
+ $Y2=0
cc_226 N_A_90_23#_c_106_n N_A_485_65#_c_716_n 0.0289875f $X=4.085 $Y=1.16 $X2=0
+ $Y2=0
cc_227 N_A_90_23#_c_106_n N_A_485_65#_c_717_n 0.0217959f $X=4.085 $Y=1.16 $X2=0
+ $Y2=0
cc_228 N_A_90_23#_c_106_n N_A_485_65#_c_706_n 0.0104705f $X=4.085 $Y=1.16 $X2=0
+ $Y2=0
cc_229 N_A_90_23#_c_107_n N_A_485_65#_c_706_n 7.75365e-19 $X=4.175 $Y=1.93 $X2=0
+ $Y2=0
cc_230 N_B1_M1013_g N_A1_M1016_g 0.0257574f $X=3.295 $Y=0.745 $X2=0 $Y2=0
cc_231 N_B1_c_256_n N_A1_M1000_g 4.85726e-19 $X=3.02 $Y=1.51 $X2=0 $Y2=0
cc_232 N_B1_M1017_g N_A1_c_315_n 0.00408523f $X=2.995 $Y=2.465 $X2=0 $Y2=0
cc_233 N_B1_c_256_n N_A1_c_315_n 0.00307247f $X=3.02 $Y=1.51 $X2=0 $Y2=0
cc_234 N_B1_c_256_n N_A1_c_318_n 0.00993482f $X=3.02 $Y=1.51 $X2=0 $Y2=0
cc_235 N_B1_c_253_n N_A1_c_318_n 0.00113931f $X=3.295 $Y=1.51 $X2=0 $Y2=0
cc_236 N_B1_c_256_n N_A1_c_312_n 6.77793e-19 $X=3.02 $Y=1.51 $X2=0 $Y2=0
cc_237 N_B1_c_253_n N_A1_c_312_n 0.0226543f $X=3.295 $Y=1.51 $X2=0 $Y2=0
cc_238 N_B1_M1008_g N_VPWR_c_457_n 0.0145295f $X=2.565 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B1_M1017_g N_VPWR_c_457_n 6.77251e-19 $X=2.995 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B1_M1017_g N_VPWR_c_497_n 0.0188239f $X=2.995 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B1_c_253_n N_VPWR_c_497_n 0.00550611f $X=3.295 $Y=1.51 $X2=0 $Y2=0
cc_242 N_B1_M1008_g N_VPWR_c_467_n 0.00486043f $X=2.565 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B1_M1017_g N_VPWR_c_467_n 0.00486043f $X=2.995 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B1_M1008_g N_VPWR_c_468_n 5.43889e-19 $X=2.565 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B1_M1017_g N_VPWR_c_468_n 0.00953603f $X=2.995 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B1_M1008_g N_VPWR_c_454_n 0.00824727f $X=2.565 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B1_M1017_g N_VPWR_c_454_n 0.00819843f $X=2.995 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B1_M1007_g N_VGND_c_616_n 0.00246418f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_249 N_B1_M1007_g N_VGND_c_621_n 0.00302501f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_250 N_B1_M1013_g N_VGND_c_621_n 0.00302501f $X=3.295 $Y=0.745 $X2=0 $Y2=0
cc_251 N_B1_M1007_g N_VGND_c_624_n 0.0048466f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_252 N_B1_M1013_g N_VGND_c_624_n 0.00442601f $X=3.295 $Y=0.745 $X2=0 $Y2=0
cc_253 N_B1_M1007_g N_A_485_65#_c_702_n 0.0127699f $X=2.865 $Y=0.745 $X2=0 $Y2=0
cc_254 N_B1_M1013_g N_A_485_65#_c_702_n 0.0115989f $X=3.295 $Y=0.745 $X2=0 $Y2=0
cc_255 N_A1_M1016_g N_A2_M1005_g 0.0308272f $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_256 N_A1_M1000_g N_A2_M1006_g 0.0326974f $X=3.885 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A1_c_315_n N_A2_M1006_g 0.00130469f $X=3.83 $Y=2.31 $X2=0 $Y2=0
cc_258 A1 N_A2_M1006_g 0.0111997f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_259 N_A1_M1019_g N_A2_M1011_g 0.0288889f $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_260 N_A1_M1015_g N_A2_M1014_g 0.0288889f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_261 A1 N_A2_M1014_g 0.0136241f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_262 N_A1_c_316_n N_A2_c_400_n 0.00820612f $X=5.04 $Y=2.31 $X2=0 $Y2=0
cc_263 N_A1_c_309_n N_A2_c_400_n 0.0172578f $X=5.125 $Y=1.535 $X2=0 $Y2=0
cc_264 N_A1_c_311_n N_A2_c_400_n 3.14489e-19 $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_265 A1 N_A2_c_400_n 0.00217636f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_266 N_A1_c_316_n N_A2_c_397_n 0.0095562f $X=5.04 $Y=2.31 $X2=0 $Y2=0
cc_267 N_A1_c_309_n N_A2_c_397_n 0.00176414f $X=5.125 $Y=1.535 $X2=0 $Y2=0
cc_268 N_A1_c_311_n N_A2_c_397_n 0.0288889f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_269 N_A1_c_318_n N_A2_c_397_n 3.2983e-19 $X=3.75 $Y=1.51 $X2=0 $Y2=0
cc_270 N_A1_c_312_n N_A2_c_397_n 0.0326974f $X=3.75 $Y=1.51 $X2=0 $Y2=0
cc_271 N_A1_c_315_n N_VPWR_M1017_d 0.00540748f $X=3.83 $Y=2.31 $X2=0 $Y2=0
cc_272 N_A1_c_358_p N_VPWR_M1017_d 0.00206053f $X=3.915 $Y=2.405 $X2=0 $Y2=0
cc_273 N_A1_M1000_g N_VPWR_c_497_n 0.011875f $X=3.885 $Y=2.465 $X2=0 $Y2=0
cc_274 N_A1_c_315_n N_VPWR_c_497_n 0.0293858f $X=3.83 $Y=2.31 $X2=0 $Y2=0
cc_275 N_A1_c_358_p N_VPWR_c_497_n 0.016181f $X=3.915 $Y=2.405 $X2=0 $Y2=0
cc_276 N_A1_M1015_g N_VPWR_c_459_n 0.00871805f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A1_c_316_n N_VPWR_c_459_n 0.0175042f $X=5.04 $Y=2.31 $X2=0 $Y2=0
cc_278 N_A1_c_310_n N_VPWR_c_459_n 0.0109957f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_279 N_A1_c_311_n N_VPWR_c_459_n 0.00323663f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_280 N_A1_M1000_g N_VPWR_c_466_n 0.00564095f $X=3.885 $Y=2.465 $X2=0 $Y2=0
cc_281 N_A1_M1015_g N_VPWR_c_466_n 0.00585385f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_282 N_A1_M1000_g N_VPWR_c_468_n 0.00931846f $X=3.885 $Y=2.465 $X2=0 $Y2=0
cc_283 N_A1_c_358_p N_VPWR_c_468_n 6.05013e-19 $X=3.915 $Y=2.405 $X2=0 $Y2=0
cc_284 N_A1_M1000_g N_VPWR_c_454_n 0.00524434f $X=3.885 $Y=2.465 $X2=0 $Y2=0
cc_285 N_A1_M1015_g N_VPWR_c_454_n 0.0110286f $X=5.175 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A1_c_316_n N_VPWR_c_454_n 0.00238129f $X=5.04 $Y=2.31 $X2=0 $Y2=0
cc_287 N_A1_c_358_p N_VPWR_c_454_n 0.00353718f $X=3.915 $Y=2.405 $X2=0 $Y2=0
cc_288 A1 N_VPWR_c_454_n 0.00378943f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_289 A1 N_A_792_367#_M1000_d 0.00541395f $X=4.955 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_290 N_A1_c_316_n N_A_792_367#_M1014_d 0.0060071f $X=5.04 $Y=2.31 $X2=0 $Y2=0
cc_291 A1 N_A_792_367#_M1014_d 0.00378934f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_292 N_A1_c_316_n N_A_792_367#_c_601_n 0.00725054f $X=5.04 $Y=2.31 $X2=0 $Y2=0
cc_293 A1 N_A_792_367#_c_601_n 0.0517563f $X=4.955 $Y=2.32 $X2=0 $Y2=0
cc_294 N_A1_M1016_g N_VGND_c_617_n 0.00332793f $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_295 N_A1_M1019_g N_VGND_c_618_n 0.0124972f $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_296 N_A1_M1016_g N_VGND_c_621_n 0.0035672f $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_297 N_A1_M1019_g N_VGND_c_623_n 0.00414769f $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_298 N_A1_M1016_g N_VGND_c_624_n 0.00509191f $X=3.805 $Y=0.745 $X2=0 $Y2=0
cc_299 N_A1_M1019_g N_VGND_c_624_n 0.00826786f $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_300 N_A1_M1016_g N_A_485_65#_c_702_n 0.00289145f $X=3.805 $Y=0.745 $X2=0
+ $Y2=0
cc_301 N_A1_M1016_g N_A_485_65#_c_723_n 0.00470958f $X=3.805 $Y=0.745 $X2=0
+ $Y2=0
cc_302 N_A1_M1016_g N_A_485_65#_c_716_n 0.00914313f $X=3.805 $Y=0.745 $X2=0
+ $Y2=0
cc_303 N_A1_M1016_g N_A_485_65#_c_717_n 7.31417e-19 $X=3.805 $Y=0.745 $X2=0
+ $Y2=0
cc_304 N_A1_M1019_g N_A_485_65#_c_705_n 0.0139982f $X=5.175 $Y=0.745 $X2=0 $Y2=0
cc_305 N_A1_c_309_n N_A_485_65#_c_705_n 0.0141511f $X=5.125 $Y=1.535 $X2=0 $Y2=0
cc_306 N_A1_c_310_n N_A_485_65#_c_705_n 0.0229279f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_307 N_A1_c_311_n N_A_485_65#_c_705_n 0.00457279f $X=5.265 $Y=1.51 $X2=0 $Y2=0
cc_308 N_A1_M1019_g N_A_485_65#_c_707_n 0.00354556f $X=5.175 $Y=0.745 $X2=0
+ $Y2=0
cc_309 N_A2_M1006_g N_VPWR_c_466_n 0.00373071f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_310 N_A2_M1014_g N_VPWR_c_466_n 0.00373071f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_311 N_A2_M1006_g N_VPWR_c_468_n 0.00144023f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_312 N_A2_M1006_g N_VPWR_c_454_n 0.00548684f $X=4.315 $Y=2.465 $X2=0 $Y2=0
cc_313 N_A2_M1014_g N_VPWR_c_454_n 0.00548684f $X=4.745 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A2_M1006_g N_A_792_367#_c_601_n 0.0122888f $X=4.315 $Y=2.465 $X2=0
+ $Y2=0
cc_315 N_A2_M1014_g N_A_792_367#_c_601_n 0.0123029f $X=4.745 $Y=2.465 $X2=0
+ $Y2=0
cc_316 N_A2_M1005_g N_VGND_c_617_n 0.00673865f $X=4.315 $Y=0.745 $X2=0 $Y2=0
cc_317 N_A2_M1011_g N_VGND_c_617_n 4.13439e-19 $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_318 N_A2_M1005_g N_VGND_c_618_n 5.515e-19 $X=4.315 $Y=0.745 $X2=0 $Y2=0
cc_319 N_A2_M1011_g N_VGND_c_618_n 0.0101667f $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_320 N_A2_M1005_g N_VGND_c_622_n 0.00305694f $X=4.315 $Y=0.745 $X2=0 $Y2=0
cc_321 N_A2_M1011_g N_VGND_c_622_n 0.00414769f $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_322 N_A2_M1005_g N_VGND_c_624_n 0.00391883f $X=4.315 $Y=0.745 $X2=0 $Y2=0
cc_323 N_A2_M1011_g N_VGND_c_624_n 0.00787505f $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_324 N_A2_M1005_g N_A_485_65#_c_723_n 6.08169e-19 $X=4.315 $Y=0.745 $X2=0
+ $Y2=0
cc_325 N_A2_M1005_g N_A_485_65#_c_716_n 0.014837f $X=4.315 $Y=0.745 $X2=0 $Y2=0
cc_326 N_A2_M1005_g N_A_485_65#_c_704_n 4.42052e-19 $X=4.315 $Y=0.745 $X2=0
+ $Y2=0
cc_327 N_A2_M1011_g N_A_485_65#_c_704_n 4.42052e-19 $X=4.745 $Y=0.745 $X2=0
+ $Y2=0
cc_328 N_A2_M1011_g N_A_485_65#_c_705_n 0.0144512f $X=4.745 $Y=0.745 $X2=0 $Y2=0
cc_329 N_A2_c_400_n N_A_485_65#_c_705_n 0.0108403f $X=4.61 $Y=1.51 $X2=0 $Y2=0
cc_330 N_A2_M1005_g N_A_485_65#_c_706_n 7.36763e-19 $X=4.315 $Y=0.745 $X2=0
+ $Y2=0
cc_331 N_A2_c_400_n N_A_485_65#_c_706_n 0.0151855f $X=4.61 $Y=1.51 $X2=0 $Y2=0
cc_332 N_A2_c_397_n N_A_485_65#_c_706_n 0.00256564f $X=4.745 $Y=1.51 $X2=0 $Y2=0
cc_333 N_VPWR_c_454_n N_X_M1002_s 0.00536646f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_334 N_VPWR_c_454_n N_X_M1012_s 0.00571434f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_335 N_VPWR_M1002_d N_X_c_548_n 0.00262981f $X=0.505 $Y=1.835 $X2=0 $Y2=0
cc_336 N_VPWR_c_455_n N_X_c_548_n 0.0220025f $X=0.63 $Y=2.18 $X2=0 $Y2=0
cc_337 N_VPWR_c_462_n N_X_c_581_n 0.0124525f $X=1.325 $Y=3.33 $X2=0 $Y2=0
cc_338 N_VPWR_c_454_n N_X_c_581_n 0.00730901f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_339 N_VPWR_M1009_d N_X_c_550_n 0.00176461f $X=1.35 $Y=1.835 $X2=0 $Y2=0
cc_340 N_VPWR_c_456_n N_X_c_550_n 0.0170777f $X=1.49 $Y=2.18 $X2=0 $Y2=0
cc_341 N_VPWR_c_464_n N_X_c_585_n 0.0120977f $X=2.185 $Y=3.33 $X2=0 $Y2=0
cc_342 N_VPWR_c_454_n N_X_c_585_n 0.00691495f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_343 N_VPWR_c_454_n N_A_792_367#_M1000_d 0.00253344f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_344 N_VPWR_c_454_n N_A_792_367#_M1014_d 0.00253292f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_466_n N_A_792_367#_c_601_n 0.0418796f $X=5.295 $Y=3.33 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_454_n N_A_792_367#_c_601_n 0.0376231f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_459_n N_A_485_65#_c_705_n 0.00505244f $X=5.39 $Y=1.98 $X2=0
+ $Y2=0
cc_348 N_X_c_543_n N_VGND_M1001_s 4.46468e-19 $X=0.645 $Y=1.14 $X2=-0.19
+ $Y2=-0.245
cc_349 N_X_c_546_n N_VGND_M1001_s 0.00196707f $X=0.217 $Y=1.225 $X2=-0.19
+ $Y2=-0.245
cc_350 N_X_c_544_n N_VGND_M1003_s 0.00176461f $X=1.505 $Y=1.14 $X2=0 $Y2=0
cc_351 N_X_c_543_n N_VGND_c_614_n 0.00524802f $X=0.645 $Y=1.14 $X2=0 $Y2=0
cc_352 N_X_c_546_n N_VGND_c_614_n 0.0185309f $X=0.217 $Y=1.225 $X2=0 $Y2=0
cc_353 N_X_c_544_n N_VGND_c_615_n 0.0170777f $X=1.505 $Y=1.14 $X2=0 $Y2=0
cc_354 N_X_c_593_p N_VGND_c_619_n 0.0124525f $X=0.74 $Y=0.42 $X2=0 $Y2=0
cc_355 N_X_c_594_p N_VGND_c_620_n 0.0124525f $X=1.6 $Y=0.42 $X2=0 $Y2=0
cc_356 N_X_M1001_d N_VGND_c_624_n 0.00536646f $X=0.6 $Y=0.245 $X2=0 $Y2=0
cc_357 N_X_M1004_d N_VGND_c_624_n 0.00536646f $X=1.46 $Y=0.245 $X2=0 $Y2=0
cc_358 N_X_c_593_p N_VGND_c_624_n 0.00730901f $X=0.74 $Y=0.42 $X2=0 $Y2=0
cc_359 N_X_c_594_p N_VGND_c_624_n 0.00730901f $X=1.6 $Y=0.42 $X2=0 $Y2=0
cc_360 N_VGND_c_616_n N_A_485_65#_c_701_n 0.0326426f $X=2.03 $Y=0.39 $X2=0 $Y2=0
cc_361 N_VGND_c_617_n N_A_485_65#_c_702_n 0.0100569f $X=4.09 $Y=0.45 $X2=0 $Y2=0
cc_362 N_VGND_c_621_n N_A_485_65#_c_702_n 0.0663614f $X=3.925 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_624_n N_A_485_65#_c_702_n 0.0368933f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_616_n N_A_485_65#_c_703_n 0.0125437f $X=2.03 $Y=0.39 $X2=0 $Y2=0
cc_365 N_VGND_c_621_n N_A_485_65#_c_703_n 0.0235489f $X=3.925 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_624_n N_A_485_65#_c_703_n 0.0128093f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_M1016_s N_A_485_65#_c_716_n 0.0051404f $X=3.88 $Y=0.325 $X2=0
+ $Y2=0
cc_368 N_VGND_c_617_n N_A_485_65#_c_716_n 0.0210125f $X=4.09 $Y=0.45 $X2=0 $Y2=0
cc_369 N_VGND_c_621_n N_A_485_65#_c_716_n 0.00196209f $X=3.925 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_622_n N_A_485_65#_c_716_n 0.00196761f $X=4.795 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_624_n N_A_485_65#_c_716_n 0.00906623f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_617_n N_A_485_65#_c_704_n 0.0105275f $X=4.09 $Y=0.45 $X2=0 $Y2=0
cc_373 N_VGND_c_618_n N_A_485_65#_c_704_n 0.0168617f $X=4.96 $Y=0.45 $X2=0 $Y2=0
cc_374 N_VGND_c_622_n N_A_485_65#_c_704_n 0.0102275f $X=4.795 $Y=0 $X2=0 $Y2=0
cc_375 N_VGND_c_624_n N_A_485_65#_c_704_n 0.00712543f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_376 N_VGND_M1011_s N_A_485_65#_c_705_n 0.00176461f $X=4.82 $Y=0.325 $X2=0
+ $Y2=0
cc_377 N_VGND_c_618_n N_A_485_65#_c_705_n 0.0170777f $X=4.96 $Y=0.45 $X2=0 $Y2=0
cc_378 N_VGND_c_618_n N_A_485_65#_c_707_n 0.0236511f $X=4.96 $Y=0.45 $X2=0 $Y2=0
cc_379 N_VGND_c_623_n N_A_485_65#_c_707_n 0.0140356f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_624_n N_A_485_65#_c_707_n 0.00977851f $X=5.52 $Y=0 $X2=0 $Y2=0
