* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 VPWR A2 a_511_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_77_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_63_367# C1 a_318_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_77_47# D1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND A2 a_813_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_813_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR A1 a_511_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_511_349# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR a_77_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 X a_77_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_511_349# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 X a_77_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_511_349# B1 a_318_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VGND B1 a_77_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_318_367# C1 a_63_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_63_367# D1 a_77_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_77_47# A1 a_813_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VGND D1 a_77_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_77_47# C1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 VGND a_77_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 X a_77_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 X a_77_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_318_367# B1 a_511_349# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 VGND C1 a_77_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 VGND a_77_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_77_47# D1 a_63_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_813_47# A1 a_77_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 VPWR a_77_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
