* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o22a_lp A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 VPWR A1 a_134_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_134_419# A2 a_232_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_30_173# B2 a_232_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_30_173# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_232_419# a_612_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_232_419# B1 a_30_173# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_232_419# B2 a_338_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_338_419# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VPWR a_232_419# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VGND A2 a_30_173# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_612_47# a_232_419# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
