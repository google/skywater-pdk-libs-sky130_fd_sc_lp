* File: sky130_fd_sc_lp__a41oi_lp.pxi.spice
* Created: Wed Sep  2 09:29:55 2020
* 
x_PM_SKY130_FD_SC_LP__A41OI_LP%A4 N_A4_M1003_g N_A4_M1010_g A4 A4 N_A4_c_72_n
+ PM_SKY130_FD_SC_LP__A41OI_LP%A4
x_PM_SKY130_FD_SC_LP__A41OI_LP%A3 N_A3_M1007_g N_A3_M1001_g A3 A3 N_A3_c_97_n
+ N_A3_c_98_n PM_SKY130_FD_SC_LP__A41OI_LP%A3
x_PM_SKY130_FD_SC_LP__A41OI_LP%A2 N_A2_M1009_g N_A2_M1002_g N_A2_c_136_n
+ N_A2_c_137_n A2 A2 A2 A2 N_A2_c_139_n PM_SKY130_FD_SC_LP__A41OI_LP%A2
x_PM_SKY130_FD_SC_LP__A41OI_LP%A1 N_A1_M1000_g N_A1_c_182_n N_A1_M1008_g
+ N_A1_c_183_n A1 A1 N_A1_c_185_n PM_SKY130_FD_SC_LP__A41OI_LP%A1
x_PM_SKY130_FD_SC_LP__A41OI_LP%B1 N_B1_c_221_n N_B1_M1005_g N_B1_c_222_n
+ N_B1_M1004_g N_B1_c_223_n N_B1_c_224_n N_B1_c_225_n N_B1_M1006_g N_B1_c_226_n
+ N_B1_c_227_n B1 B1 N_B1_c_229_n N_B1_c_230_n PM_SKY130_FD_SC_LP__A41OI_LP%B1
x_PM_SKY130_FD_SC_LP__A41OI_LP%A_27_409# N_A_27_409#_M1003_s N_A_27_409#_M1007_d
+ N_A_27_409#_M1008_d N_A_27_409#_c_274_n N_A_27_409#_c_275_n
+ N_A_27_409#_c_276_n N_A_27_409#_c_277_n N_A_27_409#_c_278_n
+ N_A_27_409#_c_279_n N_A_27_409#_c_280_n PM_SKY130_FD_SC_LP__A41OI_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__A41OI_LP%VPWR N_VPWR_M1003_d N_VPWR_M1002_d N_VPWR_c_328_n
+ N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n VPWR N_VPWR_c_332_n
+ N_VPWR_c_327_n N_VPWR_c_334_n PM_SKY130_FD_SC_LP__A41OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A41OI_LP%Y N_Y_M1000_d N_Y_M1004_d N_Y_c_368_n N_Y_c_369_n
+ N_Y_c_371_n N_Y_c_372_n N_Y_c_370_n Y N_Y_c_375_n
+ PM_SKY130_FD_SC_LP__A41OI_LP%Y
x_PM_SKY130_FD_SC_LP__A41OI_LP%VGND N_VGND_M1010_s N_VGND_M1006_d N_VGND_c_410_n
+ N_VGND_c_411_n N_VGND_c_412_n VGND N_VGND_c_413_n N_VGND_c_414_n
+ N_VGND_c_415_n N_VGND_c_416_n PM_SKY130_FD_SC_LP__A41OI_LP%VGND
cc_1 VNB N_A4_M1003_g 0.0447703f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_2 VNB N_A4_M1010_g 0.0246915f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.445
cc_3 VNB A4 0.0234322f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_4 VNB N_A4_c_72_n 0.0428322f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.975
cc_5 VNB N_A3_M1001_g 0.0523323f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.445
cc_6 VNB N_A3_c_97_n 0.0214009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A3_c_98_n 0.0177388f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.975
cc_8 VNB N_A2_M1009_g 0.0312488f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_9 VNB N_A2_c_136_n 0.0209095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_c_137_n 0.00185392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A2 0.0120812f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.975
cc_12 VNB N_A2_c_139_n 0.0153104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1000_g 0.0406925f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_14 VNB N_A1_c_182_n 0.00208309f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.81
cc_15 VNB N_A1_c_183_n 0.0234695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A1 0.00171029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_185_n 0.0165656f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.975
cc_18 VNB N_B1_c_221_n 0.0135266f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.14
cc_19 VNB N_B1_c_222_n 0.0223277f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.81
cc_20 VNB N_B1_c_223_n 0.00663733f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_21 VNB N_B1_c_224_n 0.00845382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_225_n 0.0177624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_c_226_n 0.00374626f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.975
cc_24 VNB N_B1_c_227_n 0.00768873f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.975
cc_25 VNB B1 0.00515302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B1_c_229_n 0.0163945f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.975
cc_27 VNB N_B1_c_230_n 0.0116351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_327_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_368_n 0.0197257f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.445
cc_30 VNB N_Y_c_369_n 0.00620767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_370_n 0.0336226f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.975
cc_32 VNB N_VGND_c_410_n 0.0177827f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_33 VNB N_VGND_c_411_n 0.0112965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_412_n 0.0162633f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.975
cc_35 VNB N_VGND_c_413_n 0.014713f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.975
cc_36 VNB N_VGND_c_414_n 0.0612975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_415_n 0.00511011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_416_n 0.19333f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A4_M1003_g 0.0496763f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_40 VPB N_A3_M1007_g 0.0316886f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_41 VPB N_A3_c_97_n 0.00911461f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A3_c_98_n 0.0115672f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.975
cc_43 VPB N_A2_M1002_g 0.0313463f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.445
cc_44 VPB N_A2_c_137_n 0.0105991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB A2 0.00175651f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.975
cc_46 VPB N_A1_c_182_n 0.0116001f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.81
cc_47 VPB N_A1_M1008_g 0.0313446f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.445
cc_48 VPB A1 7.45984e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B1_M1004_g 0.0359924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B1_c_226_n 0.0134868f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.975
cc_51 VPB B1 0.0020443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_27_409#_c_274_n 0.0374155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_27_409#_c_275_n 0.00254123f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.975
cc_54 VPB N_A_27_409#_c_276_n 0.010627f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.975
cc_55 VPB N_A_27_409#_c_277_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=0.975
cc_56 VPB N_A_27_409#_c_278_n 0.0164439f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.975
cc_57 VPB N_A_27_409#_c_279_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_27_409#_c_280_n 0.0090317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_328_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_329_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.975
cc_61 VPB N_VPWR_c_330_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.975
cc_62 VPB N_VPWR_c_331_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_332_n 0.0363846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_327_n 0.0552947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_334_n 0.0239038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_Y_c_371_n 0.0390561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_Y_c_372_n 0.0168327f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.975
cc_68 VPB N_Y_c_370_n 0.018132f $X=-0.19 $Y=1.655 $X2=0.775 $Y2=0.975
cc_69 N_A4_M1003_g N_A3_M1007_g 0.0319767f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_70 N_A4_M1003_g N_A3_M1001_g 0.0113064f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_71 N_A4_M1010_g N_A3_M1001_g 0.0561664f $X=0.775 $Y=0.445 $X2=0 $Y2=0
cc_72 A4 N_A3_M1001_g 0.00125176f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_73 N_A4_M1003_g N_A3_c_97_n 0.0181444f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_74 N_A4_M1003_g N_A3_c_98_n 0.0262765f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_75 A4 N_A3_c_98_n 0.036158f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_76 N_A4_c_72_n N_A3_c_98_n 0.0044625f $X=0.775 $Y=0.975 $X2=0 $Y2=0
cc_77 A4 A2 0.0102483f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_78 N_A4_M1003_g N_A_27_409#_c_274_n 0.0166777f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_79 N_A4_M1003_g N_A_27_409#_c_275_n 0.0179508f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_80 N_A4_M1003_g N_A_27_409#_c_276_n 0.00227038f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_81 N_A4_M1003_g N_A_27_409#_c_277_n 9.16417e-19 $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_82 N_A4_M1003_g N_VPWR_c_328_n 0.0186229f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_83 N_A4_M1003_g N_VPWR_c_327_n 0.014085f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_84 N_A4_M1003_g N_VPWR_c_334_n 0.00769046f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_85 N_A4_M1010_g N_VGND_c_410_n 0.0135345f $X=0.775 $Y=0.445 $X2=0 $Y2=0
cc_86 A4 N_VGND_c_410_n 0.0228504f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_87 N_A4_c_72_n N_VGND_c_410_n 0.00728544f $X=0.775 $Y=0.975 $X2=0 $Y2=0
cc_88 N_A4_M1010_g N_VGND_c_414_n 0.00486043f $X=0.775 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A4_M1010_g N_VGND_c_416_n 0.00492742f $X=0.775 $Y=0.445 $X2=0 $Y2=0
cc_90 A4 N_VGND_c_416_n 0.0146566f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_91 N_A3_M1001_g N_A2_M1009_g 0.0536938f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A3_M1007_g N_A2_M1002_g 0.0196643f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_93 N_A3_c_97_n N_A2_c_136_n 0.0209085f $X=1.075 $Y=1.615 $X2=0 $Y2=0
cc_94 N_A3_c_98_n N_A2_c_136_n 0.00113718f $X=1.075 $Y=1.615 $X2=0 $Y2=0
cc_95 N_A3_M1007_g N_A2_c_137_n 5.29533e-19 $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_96 N_A3_M1001_g A2 0.00925618f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A3_c_97_n A2 4.13429e-19 $X=1.075 $Y=1.615 $X2=0 $Y2=0
cc_98 N_A3_c_98_n A2 0.0221292f $X=1.075 $Y=1.615 $X2=0 $Y2=0
cc_99 N_A3_M1001_g N_A2_c_139_n 0.0209085f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A3_M1007_g N_A_27_409#_c_274_n 9.16417e-19 $X=1.075 $Y=2.545 $X2=0
+ $Y2=0
cc_101 N_A3_M1007_g N_A_27_409#_c_275_n 0.0179508f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_102 N_A3_c_97_n N_A_27_409#_c_275_n 8.85242e-19 $X=1.075 $Y=1.615 $X2=0 $Y2=0
cc_103 N_A3_c_98_n N_A_27_409#_c_275_n 0.0496958f $X=1.075 $Y=1.615 $X2=0 $Y2=0
cc_104 N_A3_c_98_n N_A_27_409#_c_276_n 0.0259457f $X=1.075 $Y=1.615 $X2=0 $Y2=0
cc_105 N_A3_M1007_g N_A_27_409#_c_277_n 0.0165176f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_106 N_A3_M1007_g N_A_27_409#_c_280_n 0.00164564f $X=1.075 $Y=2.545 $X2=0
+ $Y2=0
cc_107 N_A3_c_97_n N_A_27_409#_c_280_n 0.00107691f $X=1.075 $Y=1.615 $X2=0 $Y2=0
cc_108 N_A3_c_98_n N_A_27_409#_c_280_n 0.00492733f $X=1.075 $Y=1.615 $X2=0 $Y2=0
cc_109 N_A3_M1007_g N_VPWR_c_328_n 0.0175722f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_110 N_A3_M1007_g N_VPWR_c_329_n 8.63241e-19 $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_111 N_A3_M1007_g N_VPWR_c_330_n 0.00769046f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_112 N_A3_M1007_g N_VPWR_c_327_n 0.0134474f $X=1.075 $Y=2.545 $X2=0 $Y2=0
cc_113 N_A3_M1001_g N_VGND_c_410_n 0.00304577f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A3_M1001_g N_VGND_c_414_n 0.00585385f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A3_M1001_g N_VGND_c_416_n 0.0108184f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A2_M1009_g N_A1_M1000_g 0.0317578f $X=1.555 $Y=0.445 $X2=0 $Y2=0
cc_117 A2 N_A1_M1000_g 0.0118432f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_118 N_A2_c_137_n N_A1_c_182_n 0.0139741f $X=1.615 $Y=1.79 $X2=0 $Y2=0
cc_119 N_A2_M1002_g N_A1_M1008_g 0.0290426f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_120 N_A2_c_136_n N_A1_c_183_n 0.0139741f $X=1.615 $Y=1.625 $X2=0 $Y2=0
cc_121 A2 A1 0.0479466f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_122 N_A2_c_139_n A1 8.17732e-19 $X=1.615 $Y=1.285 $X2=0 $Y2=0
cc_123 N_A2_c_139_n N_A1_c_185_n 0.0139741f $X=1.615 $Y=1.285 $X2=0 $Y2=0
cc_124 N_A2_M1002_g N_A_27_409#_c_277_n 0.0166112f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_125 N_A2_M1002_g N_A_27_409#_c_278_n 0.0179678f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_126 N_A2_c_137_n N_A_27_409#_c_278_n 3.43978e-19 $X=1.615 $Y=1.79 $X2=0 $Y2=0
cc_127 A2 N_A_27_409#_c_278_n 0.0212958f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A2_M1002_g N_A_27_409#_c_279_n 9.20008e-19 $X=1.605 $Y=2.545 $X2=0
+ $Y2=0
cc_129 N_A2_M1002_g N_A_27_409#_c_280_n 0.00163378f $X=1.605 $Y=2.545 $X2=0
+ $Y2=0
cc_130 N_A2_c_137_n N_A_27_409#_c_280_n 2.25414e-19 $X=1.615 $Y=1.79 $X2=0 $Y2=0
cc_131 A2 N_A_27_409#_c_280_n 0.00449587f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_132 N_A2_M1002_g N_VPWR_c_328_n 8.63241e-19 $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_133 N_A2_M1002_g N_VPWR_c_329_n 0.017679f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_134 N_A2_M1002_g N_VPWR_c_330_n 0.00769046f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_135 N_A2_M1002_g N_VPWR_c_327_n 0.0134474f $X=1.605 $Y=2.545 $X2=0 $Y2=0
cc_136 A2 N_Y_c_369_n 0.0107107f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_137 N_A2_M1009_g N_Y_c_375_n 0.00124188f $X=1.555 $Y=0.445 $X2=0 $Y2=0
cc_138 A2 N_Y_c_375_n 0.0195547f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_139 N_A2_M1009_g N_VGND_c_414_n 0.00393362f $X=1.555 $Y=0.445 $X2=0 $Y2=0
cc_140 A2 N_VGND_c_414_n 0.00934799f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_141 N_A2_M1009_g N_VGND_c_416_n 0.00574526f $X=1.555 $Y=0.445 $X2=0 $Y2=0
cc_142 A2 N_VGND_c_416_n 0.0112118f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_143 A2 A_326_47# 0.00365071f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_144 N_A1_M1000_g N_B1_c_221_n 0.0186671f $X=2.065 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A1_c_183_n N_B1_c_222_n 0.0118132f $X=2.155 $Y=1.625 $X2=0 $Y2=0
cc_146 N_A1_M1008_g N_B1_M1004_g 0.0197328f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_147 N_A1_c_182_n N_B1_c_226_n 0.0118132f $X=2.155 $Y=1.79 $X2=0 $Y2=0
cc_148 A1 B1 0.0464033f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A1_c_185_n B1 0.00411324f $X=2.155 $Y=1.285 $X2=0 $Y2=0
cc_150 A1 N_B1_c_229_n 7.97216e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_151 N_A1_c_185_n N_B1_c_229_n 0.0118132f $X=2.155 $Y=1.285 $X2=0 $Y2=0
cc_152 N_A1_M1000_g N_B1_c_230_n 0.0014213f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_153 N_A1_M1008_g N_A_27_409#_c_277_n 9.03227e-19 $X=2.155 $Y=2.545 $X2=0
+ $Y2=0
cc_154 N_A1_c_182_n N_A_27_409#_c_278_n 5.7112e-19 $X=2.155 $Y=1.79 $X2=0 $Y2=0
cc_155 N_A1_M1008_g N_A_27_409#_c_278_n 0.0201488f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_156 A1 N_A_27_409#_c_278_n 0.0246384f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A1_M1008_g N_A_27_409#_c_279_n 0.0171582f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_158 N_A1_M1008_g N_VPWR_c_329_n 0.0158808f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_159 N_A1_M1008_g N_VPWR_c_332_n 0.00840515f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_160 N_A1_M1008_g N_VPWR_c_327_n 0.0146909f $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_161 N_A1_M1000_g N_Y_c_369_n 0.00699911f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_162 A1 N_Y_c_369_n 0.0229191f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A1_c_185_n N_Y_c_369_n 0.00138198f $X=2.155 $Y=1.285 $X2=0 $Y2=0
cc_164 N_A1_M1008_g N_Y_c_372_n 2.76452e-19 $X=2.155 $Y=2.545 $X2=0 $Y2=0
cc_165 N_A1_M1000_g N_Y_c_375_n 0.0121807f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A1_M1000_g N_VGND_c_414_n 0.00443991f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A1_M1000_g N_VGND_c_416_n 0.0077475f $X=2.065 $Y=0.445 $X2=0 $Y2=0
cc_168 N_B1_M1004_g N_A_27_409#_c_278_n 0.00446471f $X=2.685 $Y=2.545 $X2=0
+ $Y2=0
cc_169 B1 N_A_27_409#_c_278_n 0.00507306f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_170 N_B1_M1004_g N_A_27_409#_c_279_n 0.016587f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_171 N_B1_M1004_g N_VPWR_c_329_n 8.46437e-19 $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_172 N_B1_M1004_g N_VPWR_c_332_n 0.00826654f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_173 N_B1_M1004_g N_VPWR_c_327_n 0.0156126f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_174 N_B1_c_223_n N_Y_c_368_n 0.00754092f $X=2.78 $Y=0.805 $X2=0 $Y2=0
cc_175 N_B1_c_224_n N_Y_c_368_n 0.00576979f $X=2.57 $Y=0.805 $X2=0 $Y2=0
cc_176 N_B1_c_227_n N_Y_c_368_n 0.00684887f $X=2.855 $Y=0.805 $X2=0 $Y2=0
cc_177 B1 N_Y_c_368_n 0.0274862f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_178 N_B1_c_229_n N_Y_c_368_n 6.69339e-19 $X=2.725 $Y=1.285 $X2=0 $Y2=0
cc_179 N_B1_c_230_n N_Y_c_368_n 0.00534099f $X=2.745 $Y=1.12 $X2=0 $Y2=0
cc_180 N_B1_c_224_n N_Y_c_369_n 0.00194918f $X=2.57 $Y=0.805 $X2=0 $Y2=0
cc_181 N_B1_M1004_g N_Y_c_371_n 0.0143689f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_182 N_B1_M1004_g N_Y_c_372_n 0.00467277f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_183 N_B1_c_226_n N_Y_c_372_n 0.00244481f $X=2.745 $Y=1.79 $X2=0 $Y2=0
cc_184 B1 N_Y_c_372_n 0.00707451f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_185 N_B1_M1004_g N_Y_c_370_n 0.0071198f $X=2.685 $Y=2.545 $X2=0 $Y2=0
cc_186 B1 N_Y_c_370_n 0.0485299f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_187 N_B1_c_230_n N_Y_c_370_n 0.0231966f $X=2.745 $Y=1.12 $X2=0 $Y2=0
cc_188 N_B1_c_221_n N_Y_c_375_n 0.00881761f $X=2.495 $Y=0.73 $X2=0 $Y2=0
cc_189 N_B1_c_224_n N_Y_c_375_n 0.00234012f $X=2.57 $Y=0.805 $X2=0 $Y2=0
cc_190 N_B1_c_225_n N_Y_c_375_n 0.00157834f $X=2.855 $Y=0.73 $X2=0 $Y2=0
cc_191 N_B1_c_221_n N_VGND_c_412_n 0.00216659f $X=2.495 $Y=0.73 $X2=0 $Y2=0
cc_192 N_B1_c_225_n N_VGND_c_412_n 0.0119191f $X=2.855 $Y=0.73 $X2=0 $Y2=0
cc_193 N_B1_c_221_n N_VGND_c_414_n 0.00549284f $X=2.495 $Y=0.73 $X2=0 $Y2=0
cc_194 N_B1_c_223_n N_VGND_c_414_n 4.87571e-19 $X=2.78 $Y=0.805 $X2=0 $Y2=0
cc_195 N_B1_c_225_n N_VGND_c_414_n 0.00486043f $X=2.855 $Y=0.73 $X2=0 $Y2=0
cc_196 N_B1_c_221_n N_VGND_c_416_n 0.00601009f $X=2.495 $Y=0.73 $X2=0 $Y2=0
cc_197 N_B1_c_223_n N_VGND_c_416_n 6.51792e-19 $X=2.78 $Y=0.805 $X2=0 $Y2=0
cc_198 N_B1_c_225_n N_VGND_c_416_n 0.00426155f $X=2.855 $Y=0.73 $X2=0 $Y2=0
cc_199 N_A_27_409#_c_275_n N_VPWR_M1003_d 0.00180746f $X=1.175 $Y=2.055
+ $X2=-0.19 $Y2=1.655
cc_200 N_A_27_409#_c_278_n N_VPWR_M1002_d 0.00202522f $X=2.255 $Y=2.055 $X2=0
+ $Y2=0
cc_201 N_A_27_409#_c_274_n N_VPWR_c_328_n 0.0490886f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_202 N_A_27_409#_c_275_n N_VPWR_c_328_n 0.0163515f $X=1.175 $Y=2.055 $X2=0
+ $Y2=0
cc_203 N_A_27_409#_c_277_n N_VPWR_c_328_n 0.0490886f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_204 N_A_27_409#_c_277_n N_VPWR_c_329_n 0.0490886f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_205 N_A_27_409#_c_278_n N_VPWR_c_329_n 0.0164557f $X=2.255 $Y=2.055 $X2=0
+ $Y2=0
cc_206 N_A_27_409#_c_279_n N_VPWR_c_329_n 0.0454939f $X=2.42 $Y=2.19 $X2=0 $Y2=0
cc_207 N_A_27_409#_c_277_n N_VPWR_c_330_n 0.021949f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_208 N_A_27_409#_c_279_n N_VPWR_c_332_n 0.021949f $X=2.42 $Y=2.19 $X2=0 $Y2=0
cc_209 N_A_27_409#_c_274_n N_VPWR_c_327_n 0.0125808f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_210 N_A_27_409#_c_277_n N_VPWR_c_327_n 0.0124703f $X=1.34 $Y=2.19 $X2=0 $Y2=0
cc_211 N_A_27_409#_c_279_n N_VPWR_c_327_n 0.0124703f $X=2.42 $Y=2.19 $X2=0 $Y2=0
cc_212 N_A_27_409#_c_274_n N_VPWR_c_334_n 0.0220321f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_213 N_A_27_409#_c_278_n N_Y_c_372_n 0.00824572f $X=2.255 $Y=2.055 $X2=0 $Y2=0
cc_214 N_A_27_409#_c_279_n N_Y_c_372_n 0.0624161f $X=2.42 $Y=2.19 $X2=0 $Y2=0
cc_215 N_A_27_409#_c_278_n N_Y_c_370_n 0.00196599f $X=2.255 $Y=2.055 $X2=0 $Y2=0
cc_216 N_VPWR_c_332_n N_Y_c_371_n 0.0304602f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_217 N_VPWR_c_327_n N_Y_c_371_n 0.0174175f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_218 N_Y_c_368_n N_VGND_c_412_n 0.0238292f $X=3.07 $Y=0.855 $X2=0 $Y2=0
cc_219 N_Y_c_375_n N_VGND_c_412_n 0.0110361f $X=2.28 $Y=0.47 $X2=0 $Y2=0
cc_220 N_Y_c_375_n N_VGND_c_414_n 0.0223234f $X=2.28 $Y=0.47 $X2=0 $Y2=0
cc_221 N_Y_M1000_d N_VGND_c_416_n 0.0022543f $X=2.14 $Y=0.235 $X2=0 $Y2=0
cc_222 N_Y_c_368_n N_VGND_c_416_n 0.0158812f $X=3.07 $Y=0.855 $X2=0 $Y2=0
cc_223 N_Y_c_375_n N_VGND_c_416_n 0.0148533f $X=2.28 $Y=0.47 $X2=0 $Y2=0
cc_224 N_VGND_c_416_n A_170_47# 0.010279f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_225 N_VGND_c_416_n A_248_47# 0.00930162f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_226 N_VGND_c_416_n A_326_47# 0.00989122f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_227 N_VGND_c_416_n A_514_47# 0.00286135f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
