* File: sky130_fd_sc_lp__busdrivernovlp2_20.pxi.spice
* Created: Wed Sep  2 09:37:20 2020
* 
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%TE_B N_TE_B_M1052_g N_TE_B_c_376_n
+ N_TE_B_M1041_g N_TE_B_c_377_n N_TE_B_c_378_n N_TE_B_c_379_n N_TE_B_c_380_n
+ N_TE_B_M1024_g N_TE_B_c_381_n N_TE_B_c_382_n N_TE_B_M1049_g N_TE_B_M1018_g
+ N_TE_B_M1044_g N_TE_B_c_385_n N_TE_B_c_386_n N_TE_B_c_387_n N_TE_B_c_388_n
+ N_TE_B_c_389_n N_TE_B_c_390_n N_TE_B_c_391_n N_TE_B_c_435_p N_TE_B_c_392_n
+ N_TE_B_c_393_n N_TE_B_c_527_p N_TE_B_c_467_p N_TE_B_c_528_p N_TE_B_c_502_p
+ N_TE_B_c_394_n N_TE_B_c_477_p N_TE_B_c_395_n N_TE_B_c_396_n N_TE_B_c_397_n
+ N_TE_B_c_398_n TE_B N_TE_B_c_399_n N_TE_B_c_400_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%TE_B
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_27_367# N_A_27_367#_M1041_s
+ N_A_27_367#_M1052_s N_A_27_367#_c_588_n N_A_27_367#_M1015_g
+ N_A_27_367#_M1057_g N_A_27_367#_c_589_n N_A_27_367#_M1019_g
+ N_A_27_367#_c_579_n N_A_27_367#_c_580_n N_A_27_367#_M1035_g
+ N_A_27_367#_c_581_n N_A_27_367#_c_593_n N_A_27_367#_c_582_n
+ N_A_27_367#_c_583_n N_A_27_367#_c_584_n N_A_27_367#_c_585_n
+ N_A_27_367#_c_586_n N_A_27_367#_c_587_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_27_367#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_217_367# N_A_217_367#_M1020_d
+ N_A_217_367#_M1015_d N_A_217_367#_M1028_d N_A_217_367#_M1055_g
+ N_A_217_367#_c_684_n N_A_217_367#_c_685_n N_A_217_367#_M1038_g
+ N_A_217_367#_c_727_n N_A_217_367#_M1004_g N_A_217_367#_c_686_n
+ N_A_217_367#_c_687_n N_A_217_367#_c_730_n N_A_217_367#_M1008_g
+ N_A_217_367#_c_688_n N_A_217_367#_c_732_n N_A_217_367#_M1009_g
+ N_A_217_367#_c_689_n N_A_217_367#_c_734_n N_A_217_367#_M1012_g
+ N_A_217_367#_c_690_n N_A_217_367#_c_736_n N_A_217_367#_M1014_g
+ N_A_217_367#_c_691_n N_A_217_367#_c_738_n N_A_217_367#_M1016_g
+ N_A_217_367#_c_692_n N_A_217_367#_c_740_n N_A_217_367#_M1017_g
+ N_A_217_367#_c_693_n N_A_217_367#_c_742_n N_A_217_367#_M1022_g
+ N_A_217_367#_c_694_n N_A_217_367#_c_744_n N_A_217_367#_M1025_g
+ N_A_217_367#_c_695_n N_A_217_367#_c_746_n N_A_217_367#_M1026_g
+ N_A_217_367#_c_696_n N_A_217_367#_c_748_n N_A_217_367#_M1027_g
+ N_A_217_367#_c_697_n N_A_217_367#_c_750_n N_A_217_367#_M1032_g
+ N_A_217_367#_c_751_n N_A_217_367#_M1033_g N_A_217_367#_c_752_n
+ N_A_217_367#_M1036_g N_A_217_367#_c_753_n N_A_217_367#_M1037_g
+ N_A_217_367#_c_754_n N_A_217_367#_M1042_g N_A_217_367#_c_755_n
+ N_A_217_367#_M1048_g N_A_217_367#_c_756_n N_A_217_367#_M1050_g
+ N_A_217_367#_c_757_n N_A_217_367#_M1051_g N_A_217_367#_c_758_n
+ N_A_217_367#_M1053_g N_A_217_367#_c_698_n N_A_217_367#_c_699_n
+ N_A_217_367#_c_700_n N_A_217_367#_c_701_n N_A_217_367#_c_702_n
+ N_A_217_367#_c_703_n N_A_217_367#_c_704_n N_A_217_367#_c_705_n
+ N_A_217_367#_c_706_n N_A_217_367#_c_707_n N_A_217_367#_c_803_n
+ N_A_217_367#_c_808_n N_A_217_367#_c_769_n N_A_217_367#_c_770_n
+ N_A_217_367#_c_708_n N_A_217_367#_c_913_p N_A_217_367#_c_771_n
+ N_A_217_367#_c_772_n N_A_217_367#_c_709_n N_A_217_367#_c_710_n
+ N_A_217_367#_c_711_n N_A_217_367#_c_712_n N_A_217_367#_c_713_n
+ N_A_217_367#_c_714_n N_A_217_367#_c_715_n N_A_217_367#_c_716_n
+ N_A_217_367#_c_717_n N_A_217_367#_c_718_n N_A_217_367#_c_719_n
+ N_A_217_367#_c_720_n N_A_217_367#_c_721_n N_A_217_367#_c_722_n
+ N_A_217_367#_c_723_n N_A_217_367#_c_724_n N_A_217_367#_c_725_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_217_367#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_381_85# N_A_381_85#_M1055_d
+ N_A_381_85#_M1035_d N_A_381_85#_c_1185_n N_A_381_85#_c_1195_n
+ N_A_381_85#_M1007_g N_A_381_85#_c_1186_n N_A_381_85#_c_1197_n
+ N_A_381_85#_M1023_g N_A_381_85#_c_1187_n N_A_381_85#_c_1188_n
+ N_A_381_85#_c_1224_n N_A_381_85#_c_1189_n N_A_381_85#_c_1190_n
+ N_A_381_85#_c_1199_n N_A_381_85#_c_1200_n N_A_381_85#_c_1201_n
+ N_A_381_85#_c_1191_n N_A_381_85#_c_1192_n N_A_381_85#_c_1193_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_381_85#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_726_47# N_A_726_47#_M1024_d
+ N_A_726_47#_M1001_d N_A_726_47#_M1007_s N_A_726_47#_M1011_g
+ N_A_726_47#_M1000_g N_A_726_47#_M1005_g N_A_726_47#_M1006_g
+ N_A_726_47#_M1013_g N_A_726_47#_M1021_g N_A_726_47#_c_1305_n
+ N_A_726_47#_M1029_g N_A_726_47#_c_1306_n N_A_726_47#_M1034_g
+ N_A_726_47#_c_1307_n N_A_726_47#_M1040_g N_A_726_47#_c_1308_n
+ N_A_726_47#_M1043_g N_A_726_47#_c_1309_n N_A_726_47#_c_1310_n
+ N_A_726_47#_c_1311_n N_A_726_47#_M1046_g N_A_726_47#_c_1312_n
+ N_A_726_47#_c_1313_n N_A_726_47#_M1047_g N_A_726_47#_c_1314_n
+ N_A_726_47#_c_1315_n N_A_726_47#_M1054_g N_A_726_47#_c_1316_n
+ N_A_726_47#_c_1317_n N_A_726_47#_M1056_g N_A_726_47#_c_1318_n
+ N_A_726_47#_c_1319_n N_A_726_47#_M1058_g N_A_726_47#_c_1320_n
+ N_A_726_47#_c_1321_n N_A_726_47#_M1059_g N_A_726_47#_c_1322_n
+ N_A_726_47#_c_1323_n N_A_726_47#_c_1324_n N_A_726_47#_c_1325_n
+ N_A_726_47#_c_1326_n N_A_726_47#_c_1327_n N_A_726_47#_c_1328_n
+ N_A_726_47#_c_1357_n N_A_726_47#_c_1349_n N_A_726_47#_c_1434_n
+ N_A_726_47#_c_1329_n N_A_726_47#_c_1330_n N_A_726_47#_c_1331_n
+ N_A_726_47#_c_1332_n N_A_726_47#_c_1333_n N_A_726_47#_c_1334_n
+ N_A_726_47#_c_1335_n N_A_726_47#_c_1336_n N_A_726_47#_c_1337_n
+ N_A_726_47#_c_1338_n N_A_726_47#_c_1339_n N_A_726_47#_c_1340_n
+ N_A_726_47#_c_1341_n N_A_726_47#_c_1342_n N_A_726_47#_c_1343_n
+ N_A_726_47#_c_1344_n N_A_726_47#_c_1345_n N_A_726_47#_c_1346_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_726_47#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A N_A_M1030_g N_A_M1001_g N_A_c_1647_n
+ N_A_M1045_g N_A_M1010_g N_A_c_1636_n N_A_c_1637_n N_A_c_1650_n N_A_c_1651_n
+ N_A_c_1652_n N_A_c_1653_n N_A_c_1638_n N_A_c_1639_n N_A_M1002_g N_A_c_1656_n
+ N_A_M1028_g N_A_c_1641_n N_A_M1003_g N_A_c_1658_n N_A_M1031_g N_A_c_1643_n
+ N_A_c_1644_n A A N_A_c_1645_n A PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_1238_47# N_A_1238_47#_M1018_d
+ N_A_1238_47#_M1000_d N_A_1238_47#_M1020_g N_A_1238_47#_c_1795_n
+ N_A_1238_47#_c_1796_n N_A_1238_47#_M1039_g N_A_1238_47#_c_1807_n
+ N_A_1238_47#_c_1797_n N_A_1238_47#_c_1798_n N_A_1238_47#_c_1799_n
+ N_A_1238_47#_c_1804_n N_A_1238_47#_c_1800_n N_A_1238_47#_c_1805_n
+ N_A_1238_47#_c_1806_n N_A_1238_47#_c_1801_n N_A_1238_47#_c_1802_n
+ N_A_1238_47#_c_1803_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_1238_47#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%VPWR N_VPWR_M1052_d N_VPWR_M1019_s
+ N_VPWR_M1038_d N_VPWR_M1030_d N_VPWR_M1044_s N_VPWR_M1028_s N_VPWR_M1031_s
+ N_VPWR_M1008_d N_VPWR_M1012_d N_VPWR_M1016_d N_VPWR_M1022_d N_VPWR_M1026_d
+ N_VPWR_M1032_d N_VPWR_M1036_d N_VPWR_M1042_d N_VPWR_M1050_d N_VPWR_M1053_d
+ N_VPWR_c_1922_n N_VPWR_c_1923_n N_VPWR_c_1924_n N_VPWR_c_1925_n
+ N_VPWR_c_1926_n N_VPWR_c_1927_n N_VPWR_c_1928_n N_VPWR_c_1929_n
+ N_VPWR_c_1930_n N_VPWR_c_1931_n N_VPWR_c_1932_n N_VPWR_c_1933_n
+ N_VPWR_c_1934_n N_VPWR_c_1935_n N_VPWR_c_1936_n N_VPWR_c_1937_n
+ N_VPWR_c_1938_n N_VPWR_c_1939_n N_VPWR_c_1940_n N_VPWR_c_1941_n
+ N_VPWR_c_1942_n N_VPWR_c_1943_n N_VPWR_c_1944_n N_VPWR_c_1945_n
+ N_VPWR_c_1946_n N_VPWR_c_1947_n N_VPWR_c_1948_n N_VPWR_c_1949_n
+ N_VPWR_c_1950_n N_VPWR_c_1951_n N_VPWR_c_1952_n N_VPWR_c_1953_n
+ N_VPWR_c_1954_n N_VPWR_c_1955_n N_VPWR_c_1956_n N_VPWR_c_1957_n
+ N_VPWR_c_1958_n N_VPWR_c_1959_n VPWR N_VPWR_c_1960_n N_VPWR_c_1961_n
+ N_VPWR_c_1962_n N_VPWR_c_1963_n N_VPWR_c_1964_n N_VPWR_c_1965_n
+ N_VPWR_c_1966_n N_VPWR_c_1967_n N_VPWR_c_1968_n N_VPWR_c_1969_n
+ N_VPWR_c_1970_n N_VPWR_c_1971_n N_VPWR_c_1972_n N_VPWR_c_1921_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%VPWR
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_658_367# N_A_658_367#_M1007_d
+ N_A_658_367#_M1023_d N_A_658_367#_M1045_s N_A_658_367#_c_2236_n
+ N_A_658_367#_c_2195_n N_A_658_367#_c_2208_n N_A_658_367#_c_2196_n
+ N_A_658_367#_c_2212_n N_A_658_367#_c_2201_n N_A_658_367#_c_2197_n
+ N_A_658_367#_c_2214_n N_A_658_367#_c_2198_n
+ PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_658_367#
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%Z N_Z_M1005_s N_Z_M1006_s N_Z_M1021_s
+ N_Z_M1034_s N_Z_M1043_s N_Z_M1047_s N_Z_M1056_s N_Z_M1059_s N_Z_M1004_s
+ N_Z_M1009_s N_Z_M1014_s N_Z_M1017_s N_Z_M1025_s N_Z_M1027_s N_Z_M1033_s
+ N_Z_M1037_s N_Z_M1048_s N_Z_M1051_s N_Z_c_2258_n N_Z_c_2448_n N_Z_c_2262_n
+ N_Z_c_2250_n N_Z_c_2276_n Z N_Z_c_2251_n N_Z_c_2252_n N_Z_c_2253_n
+ N_Z_c_2254_n N_Z_c_2255_n N_Z_c_2256_n N_Z_c_2257_n N_Z_c_2337_n N_Z_c_2343_n
+ N_Z_c_2376_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%Z
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%VGND N_VGND_M1041_d N_VGND_M1024_s
+ N_VGND_M1049_s N_VGND_M1010_s N_VGND_M1011_d N_VGND_M1002_d N_VGND_M1005_d
+ N_VGND_M1013_d N_VGND_M1029_d N_VGND_M1040_d N_VGND_M1046_d N_VGND_M1054_d
+ N_VGND_M1058_d N_VGND_c_2515_n N_VGND_c_2516_n N_VGND_c_2517_n N_VGND_c_2518_n
+ N_VGND_c_2519_n N_VGND_c_2520_n N_VGND_c_2521_n N_VGND_c_2522_n
+ N_VGND_c_2523_n N_VGND_c_2524_n N_VGND_c_2525_n N_VGND_c_2526_n
+ N_VGND_c_2527_n N_VGND_c_2528_n N_VGND_c_2529_n N_VGND_c_2530_n
+ N_VGND_c_2531_n N_VGND_c_2532_n N_VGND_c_2533_n N_VGND_c_2534_n
+ N_VGND_c_2535_n N_VGND_c_2536_n N_VGND_c_2537_n N_VGND_c_2538_n
+ N_VGND_c_2539_n N_VGND_c_2540_n N_VGND_c_2541_n N_VGND_c_2542_n
+ N_VGND_c_2543_n N_VGND_c_2544_n VGND N_VGND_c_2545_n N_VGND_c_2546_n
+ N_VGND_c_2547_n N_VGND_c_2548_n N_VGND_c_2549_n N_VGND_c_2550_n
+ N_VGND_c_2551_n N_VGND_c_2552_n N_VGND_c_2553_n N_VGND_c_2554_n
+ N_VGND_c_2555_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%VGND
x_PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_1451_47# N_A_1451_47#_M1002_s
+ N_A_1451_47#_M1003_s N_A_1451_47#_M1039_s N_A_1451_47#_c_2767_n
+ N_A_1451_47#_c_2757_n N_A_1451_47#_c_2758_n N_A_1451_47#_c_2788_n
+ N_A_1451_47#_c_2789_n N_A_1451_47#_c_2762_n N_A_1451_47#_c_2759_n
+ N_A_1451_47#_c_2760_n PM_SKY130_FD_SC_LP__BUSDRIVERNOVLP2_20%A_1451_47#
cc_1 VNB N_TE_B_M1052_g 0.0206588f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.255
cc_2 VNB N_TE_B_c_376_n 0.0220037f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.955
cc_3 VNB N_TE_B_c_377_n 0.0175294f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=1.185
cc_4 VNB N_TE_B_c_378_n 0.0326205f $X=-0.19 $Y=-0.245 $X2=3.48 $Y2=1.26
cc_5 VNB N_TE_B_c_379_n 0.00838124f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=1.26
cc_6 VNB N_TE_B_c_380_n 0.0202044f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.185
cc_7 VNB N_TE_B_c_381_n 0.0211028f $X=-0.19 $Y=-0.245 $X2=3.91 $Y2=1.26
cc_8 VNB N_TE_B_c_382_n 0.0178456f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.185
cc_9 VNB N_TE_B_M1018_g 0.0332197f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.445
cc_10 VNB N_TE_B_M1044_g 0.018868f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=2.285
cc_11 VNB N_TE_B_c_385_n 0.0188663f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.935
cc_12 VNB N_TE_B_c_386_n 0.00514667f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.26
cc_13 VNB N_TE_B_c_387_n 0.0148477f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=1.08
cc_14 VNB N_TE_B_c_388_n 0.00255682f $X=-0.19 $Y=-0.245 $X2=1.655 $Y2=0.995
cc_15 VNB N_TE_B_c_389_n 0.0123515f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=0.35
cc_16 VNB N_TE_B_c_390_n 0.00235291f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=0.35
cc_17 VNB N_TE_B_c_391_n 0.00381153f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.435
cc_18 VNB N_TE_B_c_392_n 0.00287082f $X=-0.19 $Y=-0.245 $X2=3.335 $Y2=0.935
cc_19 VNB N_TE_B_c_393_n 0.00288925f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=0.935
cc_20 VNB N_TE_B_c_394_n 0.00180757f $X=-0.19 $Y=-0.245 $X2=5.815 $Y2=0.73
cc_21 VNB N_TE_B_c_395_n 0.00189697f $X=-0.19 $Y=-0.245 $X2=5.9 $Y2=0.995
cc_22 VNB N_TE_B_c_396_n 0.0541699f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.43
cc_23 VNB N_TE_B_c_397_n 0.00287105f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=1.16
cc_24 VNB N_TE_B_c_398_n 0.0371169f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=1.16
cc_25 VNB N_TE_B_c_399_n 0.0602824f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.16
cc_26 VNB N_TE_B_c_400_n 0.00340124f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.08
cc_27 VNB N_A_27_367#_M1057_g 0.0375773f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.185
cc_28 VNB N_A_27_367#_c_579_n 0.0158978f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.185
cc_29 VNB N_A_27_367#_c_580_n 0.0462521f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=0.655
cc_30 VNB N_A_27_367#_c_581_n 0.0377619f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=1.325
cc_31 VNB N_A_27_367#_c_582_n 0.0115318f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.935
cc_32 VNB N_A_27_367#_c_583_n 0.00985484f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.26
cc_33 VNB N_A_27_367#_c_584_n 0.00282795f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=1.08
cc_34 VNB N_A_27_367#_c_585_n 0.00844601f $X=-0.19 $Y=-0.245 $X2=1.655 $Y2=0.435
cc_35 VNB N_A_27_367#_c_586_n 0.0127763f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=0.35
cc_36 VNB N_A_27_367#_c_587_n 0.00264894f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=0.935
cc_37 VNB N_A_217_367#_M1055_g 0.0291401f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.185
cc_38 VNB N_A_217_367#_c_684_n 0.0388231f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=0.655
cc_39 VNB N_A_217_367#_c_685_n 0.00787644f $X=-0.19 $Y=-0.245 $X2=3.91 $Y2=1.26
cc_40 VNB N_A_217_367#_c_686_n 0.0103042f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=2.285
cc_41 VNB N_A_217_367#_c_687_n 0.00528518f $X=-0.19 $Y=-0.245 $X2=6.225
+ $Y2=2.285
cc_42 VNB N_A_217_367#_c_688_n 0.00532452f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.26
cc_43 VNB N_A_217_367#_c_689_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=0.35
cc_44 VNB N_A_217_367#_c_690_n 0.00536775f $X=-0.19 $Y=-0.245 $X2=2.805
+ $Y2=0.935
cc_45 VNB N_A_217_367#_c_691_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=0.435
cc_46 VNB N_A_217_367#_c_692_n 0.00536775f $X=-0.19 $Y=-0.245 $X2=5.9 $Y2=0.995
cc_47 VNB N_A_217_367#_c_693_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_217_367#_c_694_n 0.00536775f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_49 VNB N_A_217_367#_c_695_n 0.0051871f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.14
cc_50 VNB N_A_217_367#_c_696_n 0.00536775f $X=-0.19 $Y=-0.245 $X2=6.125
+ $Y2=0.995
cc_51 VNB N_A_217_367#_c_697_n 0.0075543f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.295
cc_52 VNB N_A_217_367#_c_698_n 0.00458719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_217_367#_c_699_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_217_367#_c_700_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_217_367#_c_701_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_217_367#_c_702_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_217_367#_c_703_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_217_367#_c_704_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_217_367#_c_705_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_217_367#_c_706_n 0.00287895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_217_367#_c_707_n 0.00385496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_217_367#_c_708_n 0.00269618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_217_367#_c_709_n 0.00781829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_217_367#_c_710_n 9.52526e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_217_367#_c_711_n 0.00101889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_217_367#_c_712_n 0.0124127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_217_367#_c_713_n 0.00181686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_217_367#_c_714_n 5.78534e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_217_367#_c_715_n 0.00344362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_217_367#_c_716_n 0.0164159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_217_367#_c_717_n 0.00865742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_217_367#_c_718_n 0.00272707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_217_367#_c_719_n 0.0206894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_217_367#_c_720_n 0.00173813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_217_367#_c_721_n 0.00173813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_217_367#_c_722_n 0.00173813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_217_367#_c_723_n 0.216896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_217_367#_c_724_n 0.0225506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_217_367#_c_725_n 0.00251871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_381_85#_c_1185_n 0.0122024f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.635
cc_81 VNB N_A_381_85#_c_1186_n 0.0136934f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.185
cc_82 VNB N_A_381_85#_c_1187_n 0.00359656f $X=-0.19 $Y=-0.245 $X2=3.985
+ $Y2=1.185
cc_83 VNB N_A_381_85#_c_1188_n 0.00555492f $X=-0.19 $Y=-0.245 $X2=6.115
+ $Y2=0.995
cc_84 VNB N_A_381_85#_c_1189_n 0.00823802f $X=-0.19 $Y=-0.245 $X2=6.225
+ $Y2=2.285
cc_85 VNB N_A_381_85#_c_1190_n 0.00245372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_381_85#_c_1191_n 0.00156675f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=0.35
cc_87 VNB N_A_381_85#_c_1192_n 0.00920877f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.435
cc_88 VNB N_A_381_85#_c_1193_n 0.0076243f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.85
cc_89 VNB N_A_726_47#_M1011_g 0.0336598f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.185
cc_90 VNB N_A_726_47#_M1005_g 0.023129f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.995
cc_91 VNB N_A_726_47#_M1006_g 0.0180558f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=1.325
cc_92 VNB N_A_726_47#_M1013_g 0.0180558f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.77
cc_93 VNB N_A_726_47#_M1021_g 0.0180558f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.08
cc_94 VNB N_A_726_47#_c_1305_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=1.655 $Y2=0.995
cc_95 VNB N_A_726_47#_c_1306_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.435
cc_96 VNB N_A_726_47#_c_1307_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=0.935
cc_97 VNB N_A_726_47#_c_1308_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=4.035 $Y2=0.35
cc_98 VNB N_A_726_47#_c_1309_n 0.0124835f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=0.645
cc_99 VNB N_A_726_47#_c_1310_n 0.175774f $X=-0.19 $Y=-0.245 $X2=5.815 $Y2=0.73
cc_100 VNB N_A_726_47#_c_1311_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=4.205 $Y2=0.73
cc_101 VNB N_A_726_47#_c_1312_n 0.0112546f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.35
cc_102 VNB N_A_726_47#_c_1313_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.43
cc_103 VNB N_A_726_47#_c_1314_n 0.0101163f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=1.16
cc_104 VNB N_A_726_47#_c_1315_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=1.16
cc_105 VNB N_A_726_47#_c_1316_n 0.0112546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_726_47#_c_1317_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_726_47#_c_1318_n 0.0101163f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.16
cc_108 VNB N_A_726_47#_c_1319_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.955
cc_109 VNB N_A_726_47#_c_1320_n 0.020322f $X=-0.19 $Y=-0.245 $X2=6.125 $Y2=1.325
cc_110 VNB N_A_726_47#_c_1321_n 0.0200313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_726_47#_c_1322_n 0.0233096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_726_47#_c_1323_n 0.00960202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_726_47#_c_1324_n 0.00578834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_726_47#_c_1325_n 0.00478657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_726_47#_c_1326_n 0.00478657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_726_47#_c_1327_n 0.00478657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_726_47#_c_1328_n 0.00478657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_726_47#_c_1329_n 0.0104357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_726_47#_c_1330_n 9.58006e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_726_47#_c_1331_n 0.0123812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_726_47#_c_1332_n 0.00490005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_726_47#_c_1333_n 0.00239286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_726_47#_c_1334_n 0.0231212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_726_47#_c_1335_n 0.0020192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_726_47#_c_1336_n 0.00112406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_726_47#_c_1337_n 0.013306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_726_47#_c_1338_n 0.0160487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_726_47#_c_1339_n 0.0108798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_726_47#_c_1340_n 0.0715275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_726_47#_c_1341_n 0.00922276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_726_47#_c_1342_n 0.00365776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_726_47#_c_1343_n 0.00365776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_726_47#_c_1344_n 0.00273005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_726_47#_c_1345_n 0.00273005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_726_47#_c_1346_n 0.00378122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_M1030_g 0.00900488f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.255
cc_137 VNB N_A_M1001_g 0.0305546f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.635
cc_138 VNB N_A_M1010_g 0.0285556f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=0.655
cc_139 VNB N_A_c_1636_n 0.0147362f $X=-0.19 $Y=-0.245 $X2=3.63 $Y2=1.26
cc_140 VNB N_A_c_1637_n 0.0539752f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.185
cc_141 VNB N_A_c_1638_n 0.012535f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=1.325
cc_142 VNB N_A_c_1639_n 0.0063278f $X=-0.19 $Y=-0.245 $X2=6.225 $Y2=2.285
cc_143 VNB N_A_M1002_g 0.0411809f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.77
cc_144 VNB N_A_c_1641_n 0.00496652f $X=-0.19 $Y=-0.245 $X2=1.655 $Y2=0.435
cc_145 VNB N_A_M1003_g 0.0330916f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.435
cc_146 VNB N_A_c_1643_n 0.00152826f $X=-0.19 $Y=-0.245 $X2=3.42 $Y2=0.85
cc_147 VNB N_A_c_1644_n 0.00437974f $X=-0.19 $Y=-0.245 $X2=4.035 $Y2=0.35
cc_148 VNB N_A_c_1645_n 0.00472961f $X=-0.19 $Y=-0.245 $X2=5.9 $Y2=1.16
cc_149 VNB N_A_1238_47#_c_1795_n 0.0257056f $X=-0.19 $Y=-0.245 $X2=3.48 $Y2=1.26
cc_150 VNB N_A_1238_47#_c_1796_n 0.0195693f $X=-0.19 $Y=-0.245 $X2=3.555
+ $Y2=1.185
cc_151 VNB N_A_1238_47#_c_1797_n 0.00940815f $X=-0.19 $Y=-0.245 $X2=3.985
+ $Y2=0.655
cc_152 VNB N_A_1238_47#_c_1798_n 0.00290084f $X=-0.19 $Y=-0.245 $X2=6.115
+ $Y2=0.995
cc_153 VNB N_A_1238_47#_c_1799_n 0.0102806f $X=-0.19 $Y=-0.245 $X2=6.225
+ $Y2=1.325
cc_154 VNB N_A_1238_47#_c_1800_n 0.00845788f $X=-0.19 $Y=-0.245 $X2=2.64
+ $Y2=0.935
cc_155 VNB N_A_1238_47#_c_1801_n 0.0025247f $X=-0.19 $Y=-0.245 $X2=2.64
+ $Y2=0.435
cc_156 VNB N_A_1238_47#_c_1802_n 0.0411758f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.85
cc_157 VNB N_A_1238_47#_c_1803_n 0.0177135f $X=-0.19 $Y=-0.245 $X2=3.335
+ $Y2=0.935
cc_158 VNB N_VPWR_c_1921_n 0.740851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_Z_c_2250_n 0.0203439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_Z_c_2251_n 0.00437785f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.08
cc_161 VNB N_Z_c_2252_n 0.00437785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_Z_c_2253_n 0.00437785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_Z_c_2254_n 0.00846135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_Z_c_2255_n 0.00549438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_Z_c_2256_n 0.00549438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_Z_c_2257_n 0.045274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2515_n 0.00995635f $X=-0.19 $Y=-0.245 $X2=3.42 $Y2=0.85
cc_168 VNB N_VGND_c_2516_n 0.00474148f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=0.645
cc_169 VNB N_VGND_c_2517_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=5.9 $Y2=0.995
cc_170 VNB N_VGND_c_2518_n 0.00487424f $X=-0.19 $Y=-0.245 $X2=5.9 $Y2=1.16
cc_171 VNB N_VGND_c_2519_n 0.00547112f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=1.16
cc_172 VNB N_VGND_c_2520_n 0.00238736f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0.43
cc_173 VNB N_VGND_c_2521_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.16
cc_174 VNB N_VGND_c_2522_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=6.125 $Y2=0.995
cc_175 VNB N_VGND_c_2523_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.08
cc_176 VNB N_VGND_c_2524_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2525_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2526_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2527_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2528_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2529_n 0.0216955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2530_n 0.00631443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2531_n 0.020053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2532_n 0.00516045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2533_n 0.0637743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_VGND_c_2534_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2535_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_VGND_c_2536_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_189 VNB N_VGND_c_2537_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_190 VNB N_VGND_c_2538_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_191 VNB N_VGND_c_2539_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_192 VNB N_VGND_c_2540_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_193 VNB N_VGND_c_2541_n 0.0185788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_194 VNB N_VGND_c_2542_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_195 VNB N_VGND_c_2543_n 0.018736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_196 VNB N_VGND_c_2544_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_197 VNB N_VGND_c_2545_n 0.0316002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_198 VNB N_VGND_c_2546_n 0.039312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_199 VNB N_VGND_c_2547_n 0.030281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_200 VNB N_VGND_c_2548_n 0.0198122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_201 VNB N_VGND_c_2549_n 0.0600283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_202 VNB N_VGND_c_2550_n 0.898453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_203 VNB N_VGND_c_2551_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_204 VNB N_VGND_c_2552_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_205 VNB N_VGND_c_2553_n 0.00510127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_206 VNB N_VGND_c_2554_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_207 VNB N_VGND_c_2555_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_208 VNB N_A_1451_47#_c_2757_n 0.00425653f $X=-0.19 $Y=-0.245 $X2=3.555
+ $Y2=1.185
cc_209 VNB N_A_1451_47#_c_2758_n 0.00119772f $X=-0.19 $Y=-0.245 $X2=3.555
+ $Y2=0.655
cc_210 VNB N_A_1451_47#_c_2759_n 0.00233608f $X=-0.19 $Y=-0.245 $X2=6.115
+ $Y2=0.445
cc_211 VNB N_A_1451_47#_c_2760_n 0.014871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_212 VPB N_TE_B_M1052_g 0.0268849f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.255
cc_213 VPB N_TE_B_M1044_g 0.0196873f $X=-0.19 $Y=1.655 $X2=6.225 $Y2=2.285
cc_214 VPB N_A_27_367#_c_588_n 0.0194767f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.635
cc_215 VPB N_A_27_367#_c_589_n 0.0171486f $X=-0.19 $Y=1.655 $X2=3.555 $Y2=0.655
cc_216 VPB N_A_27_367#_c_579_n 0.00897032f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=1.185
cc_217 VPB N_A_27_367#_c_580_n 0.0075659f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=0.655
cc_218 VPB N_A_27_367#_M1035_g 0.0388776f $X=-0.19 $Y=1.655 $X2=6.115 $Y2=0.445
cc_219 VPB N_A_27_367#_c_593_n 0.0403208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_27_367#_c_584_n 0.00700955f $X=-0.19 $Y=1.655 $X2=1.57 $Y2=1.08
cc_221 VPB N_A_27_367#_c_585_n 0.00476183f $X=-0.19 $Y=1.655 $X2=1.655 $Y2=0.435
cc_222 VPB N_A_27_367#_c_587_n 0.00272576f $X=-0.19 $Y=1.655 $X2=2.805 $Y2=0.935
cc_223 VPB N_A_217_367#_M1038_g 0.0339178f $X=-0.19 $Y=1.655 $X2=6.115 $Y2=0.995
cc_224 VPB N_A_217_367#_c_727_n 0.0198002f $X=-0.19 $Y=1.655 $X2=6.115 $Y2=0.445
cc_225 VPB N_A_217_367#_c_686_n 0.0049292f $X=-0.19 $Y=1.655 $X2=6.225 $Y2=2.285
cc_226 VPB N_A_217_367#_c_687_n 0.00311208f $X=-0.19 $Y=1.655 $X2=6.225
+ $Y2=2.285
cc_227 VPB N_A_217_367#_c_730_n 0.0155581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_217_367#_c_688_n 0.00544413f $X=-0.19 $Y=1.655 $X2=3.555 $Y2=1.26
cc_229 VPB N_A_217_367#_c_732_n 0.0155017f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=1.08
cc_230 VPB N_A_217_367#_c_689_n 0.0049292f $X=-0.19 $Y=1.655 $X2=2.475 $Y2=0.35
cc_231 VPB N_A_217_367#_c_734_n 0.0155111f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=0.435
cc_232 VPB N_A_217_367#_c_690_n 0.00544413f $X=-0.19 $Y=1.655 $X2=2.805
+ $Y2=0.935
cc_233 VPB N_A_217_367#_c_736_n 0.0155111f $X=-0.19 $Y=1.655 $X2=3.42 $Y2=0.85
cc_234 VPB N_A_217_367#_c_691_n 0.0049292f $X=-0.19 $Y=1.655 $X2=4.12 $Y2=0.435
cc_235 VPB N_A_217_367#_c_738_n 0.0155111f $X=-0.19 $Y=1.655 $X2=5.815 $Y2=0.73
cc_236 VPB N_A_217_367#_c_692_n 0.00544413f $X=-0.19 $Y=1.655 $X2=5.9 $Y2=0.995
cc_237 VPB N_A_217_367#_c_740_n 0.0155111f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=0.43
cc_238 VPB N_A_217_367#_c_693_n 0.0049292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_217_367#_c_742_n 0.0155111f $X=-0.19 $Y=1.655 $X2=6.115 $Y2=1.16
cc_240 VPB N_A_217_367#_c_694_n 0.00544413f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_241 VPB N_A_217_367#_c_744_n 0.0155111f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=0.43
cc_242 VPB N_A_217_367#_c_695_n 0.0049292f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.14
cc_243 VPB N_A_217_367#_c_746_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.16
cc_244 VPB N_A_217_367#_c_696_n 0.00544413f $X=-0.19 $Y=1.655 $X2=6.125
+ $Y2=0.995
cc_245 VPB N_A_217_367#_c_748_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.08
cc_246 VPB N_A_217_367#_c_697_n 0.0049292f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.295
cc_247 VPB N_A_217_367#_c_750_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_217_367#_c_751_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_217_367#_c_752_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_217_367#_c_753_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_217_367#_c_754_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_217_367#_c_755_n 0.0155111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_217_367#_c_756_n 0.0155152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_217_367#_c_757_n 0.0157552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_217_367#_c_758_n 0.0220709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_A_217_367#_c_698_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_217_367#_c_699_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_217_367#_c_700_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_217_367#_c_701_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_217_367#_c_702_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_217_367#_c_703_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_217_367#_c_704_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_217_367#_c_705_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_217_367#_c_706_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_217_367#_c_707_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_217_367#_c_769_n 0.00176583f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_217_367#_c_770_n 0.00147517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_217_367#_c_771_n 0.00476041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_217_367#_c_772_n 0.00180684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_217_367#_c_711_n 0.00291626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_217_367#_c_712_n 0.055471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_217_367#_c_714_n 4.18656e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_217_367#_c_715_n 0.00138281f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_A_217_367#_c_716_n 0.0160971f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_217_367#_c_717_n 0.0185751f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_217_367#_c_718_n 0.00431137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_A_217_367#_c_720_n 0.00187511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_A_217_367#_c_721_n 0.00187511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_217_367#_c_722_n 0.00187511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_A_217_367#_c_723_n 0.0534031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_A_217_367#_c_724_n 0.00353111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_A_217_367#_c_725_n 0.00286453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_A_381_85#_c_1185_n 0.0192899f $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.635
cc_284 VPB N_A_381_85#_c_1195_n 0.0190474f $X=-0.19 $Y=1.655 $X2=2.73 $Y2=1.185
cc_285 VPB N_A_381_85#_c_1186_n 0.00762556f $X=-0.19 $Y=1.655 $X2=3.555
+ $Y2=1.185
cc_286 VPB N_A_381_85#_c_1197_n 0.0169015f $X=-0.19 $Y=1.655 $X2=3.555 $Y2=0.655
cc_287 VPB N_A_381_85#_c_1187_n 0.00111435f $X=-0.19 $Y=1.655 $X2=3.985
+ $Y2=1.185
cc_288 VPB N_A_381_85#_c_1199_n 0.0271509f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=0.77
cc_289 VPB N_A_381_85#_c_1200_n 0.00216462f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=0.935
cc_290 VPB N_A_381_85#_c_1201_n 0.00351484f $X=-0.19 $Y=1.655 $X2=1.655
+ $Y2=0.435
cc_291 VPB N_A_381_85#_c_1193_n 0.0263483f $X=-0.19 $Y=1.655 $X2=2.64 $Y2=0.85
cc_292 VPB N_A_726_47#_M1000_g 0.0199761f $X=-0.19 $Y=1.655 $X2=3.63 $Y2=1.26
cc_293 VPB N_A_726_47#_c_1323_n 0.00665481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_A_726_47#_c_1349_n 8.73487e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_295 VPB N_A_726_47#_c_1331_n 8.88856e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_296 VPB N_A_726_47#_c_1339_n 0.00163717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_A_M1030_g 0.020105f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.255
cc_298 VPB N_A_c_1647_n 0.0173776f $X=-0.19 $Y=1.655 $X2=2.73 $Y2=1.185
cc_299 VPB N_A_c_1636_n 0.00568288f $X=-0.19 $Y=1.655 $X2=3.63 $Y2=1.26
cc_300 VPB N_A_c_1637_n 0.0127767f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=1.185
cc_301 VPB N_A_c_1650_n 0.0844944f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=0.655
cc_302 VPB N_A_c_1651_n 0.101846f $X=-0.19 $Y=1.655 $X2=6.115 $Y2=0.995
cc_303 VPB N_A_c_1652_n 0.0107356f $X=-0.19 $Y=1.655 $X2=6.115 $Y2=0.445
cc_304 VPB N_A_c_1653_n 0.0828094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_A_c_1638_n 0.00893085f $X=-0.19 $Y=1.655 $X2=6.225 $Y2=1.325
cc_306 VPB N_A_c_1639_n 0.00218133f $X=-0.19 $Y=1.655 $X2=6.225 $Y2=2.285
cc_307 VPB N_A_c_1656_n 0.0167171f $X=-0.19 $Y=1.655 $X2=3.555 $Y2=1.26
cc_308 VPB N_A_c_1641_n 0.00522816f $X=-0.19 $Y=1.655 $X2=1.655 $Y2=0.435
cc_309 VPB N_A_c_1658_n 0.0207545f $X=-0.19 $Y=1.655 $X2=3.335 $Y2=0.935
cc_310 VPB N_A_c_1643_n 0.00133723f $X=-0.19 $Y=1.655 $X2=3.42 $Y2=0.85
cc_311 VPB N_A_c_1644_n 0.00371853f $X=-0.19 $Y=1.655 $X2=4.035 $Y2=0.35
cc_312 VPB A 0.00331767f $X=-0.19 $Y=1.655 $X2=3.505 $Y2=0.35
cc_313 VPB N_A_c_1645_n 2.57446e-19 $X=-0.19 $Y=1.655 $X2=5.9 $Y2=1.16
cc_314 VPB N_A_1238_47#_c_1804_n 0.00221686f $X=-0.19 $Y=1.655 $X2=6.225
+ $Y2=2.285
cc_315 VPB N_A_1238_47#_c_1805_n 0.00860599f $X=-0.19 $Y=1.655 $X2=1.655
+ $Y2=0.435
cc_316 VPB N_A_1238_47#_c_1806_n 0.00465637f $X=-0.19 $Y=1.655 $X2=2.475
+ $Y2=0.35
cc_317 VPB N_VPWR_c_1922_n 0.0171007f $X=-0.19 $Y=1.655 $X2=5.9 $Y2=1.16
cc_318 VPB N_VPWR_c_1923_n 0.00516841f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_319 VPB N_VPWR_c_1924_n 0.0170611f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.14
cc_320 VPB N_VPWR_c_1925_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.93 $Y2=0.955
cc_321 VPB N_VPWR_c_1926_n 0.022125f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.08
cc_322 VPB N_VPWR_c_1927_n 0.0133128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_1928_n 0.00752604f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_1929_n 0.00238736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_1930_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_1931_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_1932_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_1933_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_1934_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_1935_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_1936_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_1937_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_1938_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_1939_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_1940_n 0.0108116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_336 VPB N_VPWR_c_1941_n 0.0352864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_337 VPB N_VPWR_c_1942_n 0.0489127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_338 VPB N_VPWR_c_1943_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_339 VPB N_VPWR_c_1944_n 0.0320257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_340 VPB N_VPWR_c_1945_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_341 VPB N_VPWR_c_1946_n 0.0194559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_342 VPB N_VPWR_c_1947_n 0.00356964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_343 VPB N_VPWR_c_1948_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_344 VPB N_VPWR_c_1949_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_345 VPB N_VPWR_c_1950_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_346 VPB N_VPWR_c_1951_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_347 VPB N_VPWR_c_1952_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_348 VPB N_VPWR_c_1953_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_349 VPB N_VPWR_c_1954_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_350 VPB N_VPWR_c_1955_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_351 VPB N_VPWR_c_1956_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_352 VPB N_VPWR_c_1957_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_353 VPB N_VPWR_c_1958_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_354 VPB N_VPWR_c_1959_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_355 VPB N_VPWR_c_1960_n 0.0207181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_356 VPB N_VPWR_c_1961_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_357 VPB N_VPWR_c_1962_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_358 VPB N_VPWR_c_1963_n 0.0226035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_359 VPB N_VPWR_c_1964_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_360 VPB N_VPWR_c_1965_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_361 VPB N_VPWR_c_1966_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_362 VPB N_VPWR_c_1967_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_363 VPB N_VPWR_c_1968_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_364 VPB N_VPWR_c_1969_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_365 VPB N_VPWR_c_1970_n 0.0128226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_366 VPB N_VPWR_c_1971_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_367 VPB N_VPWR_c_1972_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_368 VPB N_VPWR_c_1921_n 0.0833486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_369 VPB N_A_658_367#_c_2195_n 9.1862e-19 $X=-0.19 $Y=1.655 $X2=3.555
+ $Y2=1.185
cc_370 VPB N_A_658_367#_c_2196_n 0.00388039f $X=-0.19 $Y=1.655 $X2=3.985
+ $Y2=0.655
cc_371 VPB N_A_658_367#_c_2197_n 0.00370267f $X=-0.19 $Y=1.655 $X2=6.225
+ $Y2=2.285
cc_372 VPB N_A_658_367#_c_2198_n 0.00559171f $X=-0.19 $Y=1.655 $X2=2.475
+ $Y2=0.35
cc_373 N_TE_B_c_376_n N_A_27_367#_M1057_g 0.0187034f $X=0.93 $Y=0.955 $X2=0
+ $Y2=0
cc_374 N_TE_B_c_387_n N_A_27_367#_M1057_g 0.0174176f $X=1.57 $Y=1.08 $X2=0 $Y2=0
cc_375 N_TE_B_c_388_n N_A_27_367#_M1057_g 0.00496406f $X=1.655 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_TE_B_c_390_n N_A_27_367#_M1057_g 0.00103957f $X=1.74 $Y=0.35 $X2=0
+ $Y2=0
cc_377 N_TE_B_c_399_n N_A_27_367#_M1057_g 0.00512016f $X=0.67 $Y=1.16 $X2=0
+ $Y2=0
cc_378 N_TE_B_c_400_n N_A_27_367#_M1057_g 0.00142175f $X=0.67 $Y=1.08 $X2=0
+ $Y2=0
cc_379 N_TE_B_c_387_n N_A_27_367#_c_579_n 0.00371306f $X=1.57 $Y=1.08 $X2=0
+ $Y2=0
cc_380 N_TE_B_M1052_g N_A_27_367#_c_580_n 0.0269461f $X=0.48 $Y=2.255 $X2=0
+ $Y2=0
cc_381 N_TE_B_c_387_n N_A_27_367#_c_580_n 0.00426843f $X=1.57 $Y=1.08 $X2=0
+ $Y2=0
cc_382 N_TE_B_c_399_n N_A_27_367#_c_580_n 0.00167554f $X=0.67 $Y=1.16 $X2=0
+ $Y2=0
cc_383 N_TE_B_c_400_n N_A_27_367#_c_580_n 6.1328e-19 $X=0.67 $Y=1.08 $X2=0 $Y2=0
cc_384 N_TE_B_c_376_n N_A_27_367#_c_581_n 0.00309123f $X=0.93 $Y=0.955 $X2=0
+ $Y2=0
cc_385 N_TE_B_c_399_n N_A_27_367#_c_581_n 0.0184105f $X=0.67 $Y=1.16 $X2=0 $Y2=0
cc_386 N_TE_B_c_400_n N_A_27_367#_c_581_n 0.0244428f $X=0.67 $Y=1.08 $X2=0 $Y2=0
cc_387 N_TE_B_M1052_g N_A_27_367#_c_593_n 0.0173295f $X=0.48 $Y=2.255 $X2=0
+ $Y2=0
cc_388 N_TE_B_c_399_n N_A_27_367#_c_582_n 0.00553655f $X=0.67 $Y=1.16 $X2=0
+ $Y2=0
cc_389 N_TE_B_c_400_n N_A_27_367#_c_582_n 0.00323835f $X=0.67 $Y=1.08 $X2=0
+ $Y2=0
cc_390 N_TE_B_M1052_g N_A_27_367#_c_584_n 0.0138177f $X=0.48 $Y=2.255 $X2=0
+ $Y2=0
cc_391 N_TE_B_c_387_n N_A_27_367#_c_584_n 0.0094179f $X=1.57 $Y=1.08 $X2=0 $Y2=0
cc_392 N_TE_B_c_399_n N_A_27_367#_c_584_n 0.00215092f $X=0.67 $Y=1.16 $X2=0
+ $Y2=0
cc_393 N_TE_B_c_400_n N_A_27_367#_c_584_n 0.0251532f $X=0.67 $Y=1.08 $X2=0 $Y2=0
cc_394 N_TE_B_M1052_g N_A_27_367#_c_585_n 0.00507899f $X=0.48 $Y=2.255 $X2=0
+ $Y2=0
cc_395 N_TE_B_c_376_n N_A_27_367#_c_586_n 0.00547912f $X=0.93 $Y=0.955 $X2=0
+ $Y2=0
cc_396 N_TE_B_c_387_n N_A_27_367#_c_586_n 0.00232462f $X=1.57 $Y=1.08 $X2=0
+ $Y2=0
cc_397 N_TE_B_c_399_n N_A_27_367#_c_586_n 0.00719863f $X=0.67 $Y=1.16 $X2=0
+ $Y2=0
cc_398 N_TE_B_c_400_n N_A_27_367#_c_586_n 0.0205322f $X=0.67 $Y=1.08 $X2=0 $Y2=0
cc_399 N_TE_B_M1052_g N_A_27_367#_c_587_n 0.00104023f $X=0.48 $Y=2.255 $X2=0
+ $Y2=0
cc_400 N_TE_B_c_387_n N_A_27_367#_c_587_n 0.023957f $X=1.57 $Y=1.08 $X2=0 $Y2=0
cc_401 N_TE_B_c_400_n N_A_27_367#_c_587_n 0.0038595f $X=0.67 $Y=1.08 $X2=0 $Y2=0
cc_402 N_TE_B_c_387_n N_A_217_367#_M1055_g 0.0017106f $X=1.57 $Y=1.08 $X2=0
+ $Y2=0
cc_403 N_TE_B_c_388_n N_A_217_367#_M1055_g 0.00288045f $X=1.655 $Y=0.995 $X2=0
+ $Y2=0
cc_404 N_TE_B_c_389_n N_A_217_367#_M1055_g 0.0143986f $X=2.475 $Y=0.35 $X2=0
+ $Y2=0
cc_405 N_TE_B_c_435_p N_A_217_367#_M1055_g 9.729e-19 $X=2.64 $Y=0.85 $X2=0 $Y2=0
cc_406 N_TE_B_c_396_n N_A_217_367#_M1055_g 0.0104249f $X=2.64 $Y=0.43 $X2=0
+ $Y2=0
cc_407 N_TE_B_c_377_n N_A_217_367#_c_684_n 0.00453675f $X=2.73 $Y=1.185 $X2=0
+ $Y2=0
cc_408 N_TE_B_c_387_n N_A_217_367#_c_708_n 0.00757316f $X=1.57 $Y=1.08 $X2=0
+ $Y2=0
cc_409 N_TE_B_c_378_n N_A_217_367#_c_712_n 0.00429382f $X=3.48 $Y=1.26 $X2=0
+ $Y2=0
cc_410 N_TE_B_M1044_g N_A_217_367#_c_712_n 0.00945047f $X=6.225 $Y=2.285 $X2=0
+ $Y2=0
cc_411 N_TE_B_c_392_n N_A_217_367#_c_712_n 0.0126796f $X=3.335 $Y=0.935 $X2=0
+ $Y2=0
cc_412 N_TE_B_c_397_n N_A_217_367#_c_712_n 0.00270004f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_413 N_TE_B_c_398_n N_A_217_367#_c_712_n 0.00101921f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_414 N_TE_B_c_385_n N_A_217_367#_c_717_n 0.00107594f $X=2.64 $Y=0.935 $X2=0
+ $Y2=0
cc_415 N_TE_B_c_379_n N_A_217_367#_c_719_n 0.00453675f $X=2.805 $Y=1.26 $X2=0
+ $Y2=0
cc_416 N_TE_B_c_389_n N_A_381_85#_M1055_d 0.00642969f $X=2.475 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_417 N_TE_B_c_378_n N_A_381_85#_c_1185_n 0.0179855f $X=3.48 $Y=1.26 $X2=0
+ $Y2=0
cc_418 N_TE_B_c_392_n N_A_381_85#_c_1185_n 8.321e-19 $X=3.335 $Y=0.935 $X2=0
+ $Y2=0
cc_419 N_TE_B_c_381_n N_A_381_85#_c_1186_n 0.0179855f $X=3.91 $Y=1.26 $X2=0
+ $Y2=0
cc_420 N_TE_B_c_386_n N_A_381_85#_c_1187_n 0.0179855f $X=3.555 $Y=1.26 $X2=0
+ $Y2=0
cc_421 N_TE_B_c_377_n N_A_381_85#_c_1188_n 0.00483371f $X=2.73 $Y=1.185 $X2=0
+ $Y2=0
cc_422 N_TE_B_c_385_n N_A_381_85#_c_1188_n 3.56988e-19 $X=2.64 $Y=0.935 $X2=0
+ $Y2=0
cc_423 N_TE_B_c_387_n N_A_381_85#_c_1188_n 0.011083f $X=1.57 $Y=1.08 $X2=0 $Y2=0
cc_424 N_TE_B_c_388_n N_A_381_85#_c_1188_n 0.0152636f $X=1.655 $Y=0.995 $X2=0
+ $Y2=0
cc_425 N_TE_B_c_389_n N_A_381_85#_c_1188_n 0.0180114f $X=2.475 $Y=0.35 $X2=0
+ $Y2=0
cc_426 N_TE_B_c_435_p N_A_381_85#_c_1188_n 0.014099f $X=2.64 $Y=0.85 $X2=0 $Y2=0
cc_427 N_TE_B_c_393_n N_A_381_85#_c_1188_n 0.0114105f $X=2.805 $Y=0.935 $X2=0
+ $Y2=0
cc_428 N_TE_B_c_396_n N_A_381_85#_c_1188_n 0.00219292f $X=2.64 $Y=0.43 $X2=0
+ $Y2=0
cc_429 N_TE_B_c_378_n N_A_381_85#_c_1189_n 0.0125247f $X=3.48 $Y=1.26 $X2=0
+ $Y2=0
cc_430 N_TE_B_c_379_n N_A_381_85#_c_1189_n 0.00753428f $X=2.805 $Y=1.26 $X2=0
+ $Y2=0
cc_431 N_TE_B_c_385_n N_A_381_85#_c_1189_n 7.91308e-19 $X=2.64 $Y=0.935 $X2=0
+ $Y2=0
cc_432 N_TE_B_c_392_n N_A_381_85#_c_1189_n 0.012124f $X=3.335 $Y=0.935 $X2=0
+ $Y2=0
cc_433 N_TE_B_c_393_n N_A_381_85#_c_1189_n 0.0246488f $X=2.805 $Y=0.935 $X2=0
+ $Y2=0
cc_434 N_TE_B_c_378_n N_A_381_85#_c_1191_n 6.11732e-19 $X=3.48 $Y=1.26 $X2=0
+ $Y2=0
cc_435 N_TE_B_c_392_n N_A_381_85#_c_1191_n 0.00394155f $X=3.335 $Y=0.935 $X2=0
+ $Y2=0
cc_436 N_TE_B_c_379_n N_A_381_85#_c_1193_n 0.0179855f $X=2.805 $Y=1.26 $X2=0
+ $Y2=0
cc_437 N_TE_B_c_467_p N_A_726_47#_M1024_d 0.00340092f $X=4.035 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_438 N_TE_B_c_394_n N_A_726_47#_M1001_d 0.0111717f $X=5.815 $Y=0.73 $X2=0
+ $Y2=0
cc_439 N_TE_B_M1018_g N_A_726_47#_M1011_g 0.023235f $X=6.115 $Y=0.445 $X2=0
+ $Y2=0
cc_440 N_TE_B_M1044_g N_A_726_47#_M1000_g 0.0590987f $X=6.225 $Y=2.285 $X2=0
+ $Y2=0
cc_441 N_TE_B_M1044_g N_A_726_47#_c_1322_n 0.0209363f $X=6.225 $Y=2.285 $X2=0
+ $Y2=0
cc_442 N_TE_B_c_467_p N_A_726_47#_c_1357_n 0.012056f $X=4.035 $Y=0.35 $X2=0
+ $Y2=0
cc_443 N_TE_B_c_381_n N_A_726_47#_c_1349_n 4.71251e-19 $X=3.91 $Y=1.26 $X2=0
+ $Y2=0
cc_444 N_TE_B_c_382_n N_A_726_47#_c_1329_n 0.0120432f $X=3.985 $Y=1.185 $X2=0
+ $Y2=0
cc_445 N_TE_B_c_467_p N_A_726_47#_c_1329_n 0.00315383f $X=4.035 $Y=0.35 $X2=0
+ $Y2=0
cc_446 N_TE_B_c_394_n N_A_726_47#_c_1329_n 0.0721475f $X=5.815 $Y=0.73 $X2=0
+ $Y2=0
cc_447 N_TE_B_c_477_p N_A_726_47#_c_1329_n 0.00852929f $X=4.205 $Y=0.73 $X2=0
+ $Y2=0
cc_448 N_TE_B_c_380_n N_A_726_47#_c_1330_n 0.00292593f $X=3.555 $Y=1.185 $X2=0
+ $Y2=0
cc_449 N_TE_B_c_380_n N_A_726_47#_c_1331_n 4.53441e-19 $X=3.555 $Y=1.185 $X2=0
+ $Y2=0
cc_450 N_TE_B_c_381_n N_A_726_47#_c_1331_n 0.0188987f $X=3.91 $Y=1.26 $X2=0
+ $Y2=0
cc_451 N_TE_B_c_382_n N_A_726_47#_c_1331_n 4.53441e-19 $X=3.985 $Y=1.185 $X2=0
+ $Y2=0
cc_452 N_TE_B_M1044_g N_A_726_47#_c_1332_n 0.00218186f $X=6.225 $Y=2.285 $X2=0
+ $Y2=0
cc_453 N_TE_B_c_394_n N_A_726_47#_c_1332_n 0.0053601f $X=5.815 $Y=0.73 $X2=0
+ $Y2=0
cc_454 N_TE_B_c_395_n N_A_726_47#_c_1332_n 6.80643e-19 $X=5.9 $Y=0.995 $X2=0
+ $Y2=0
cc_455 N_TE_B_c_397_n N_A_726_47#_c_1332_n 0.022048f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_456 N_TE_B_c_398_n N_A_726_47#_c_1332_n 0.00310747f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_457 N_TE_B_M1044_g N_A_726_47#_c_1333_n 6.2539e-19 $X=6.225 $Y=2.285 $X2=0
+ $Y2=0
cc_458 N_TE_B_c_394_n N_A_726_47#_c_1333_n 0.00232506f $X=5.815 $Y=0.73 $X2=0
+ $Y2=0
cc_459 N_TE_B_c_397_n N_A_726_47#_c_1333_n 0.00135128f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_460 N_TE_B_M1044_g N_A_726_47#_c_1335_n 7.30184e-19 $X=6.225 $Y=2.285 $X2=0
+ $Y2=0
cc_461 N_TE_B_c_397_n N_A_726_47#_c_1335_n 0.00137254f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_462 N_TE_B_c_398_n N_A_726_47#_c_1335_n 7.57253e-19 $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_463 N_TE_B_c_397_n N_A_726_47#_c_1338_n 3.38888e-19 $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_464 N_TE_B_c_398_n N_A_726_47#_c_1338_n 0.0209363f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_465 N_TE_B_c_397_n N_A_726_47#_c_1339_n 0.0239976f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_466 N_TE_B_c_398_n N_A_726_47#_c_1339_n 0.0101228f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_467 N_TE_B_M1044_g N_A_726_47#_c_1346_n 9.13261e-19 $X=6.225 $Y=2.285 $X2=0
+ $Y2=0
cc_468 N_TE_B_c_394_n N_A_726_47#_c_1346_n 0.00978273f $X=5.815 $Y=0.73 $X2=0
+ $Y2=0
cc_469 N_TE_B_c_397_n N_A_726_47#_c_1346_n 0.0239396f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_470 N_TE_B_c_398_n N_A_726_47#_c_1346_n 8.16959e-19 $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_471 N_TE_B_c_382_n N_A_M1001_g 0.0180204f $X=3.985 $Y=1.185 $X2=0 $Y2=0
cc_472 N_TE_B_c_502_p N_A_M1001_g 0.0024976f $X=4.12 $Y=0.645 $X2=0 $Y2=0
cc_473 N_TE_B_c_394_n N_A_M1001_g 0.0139939f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_474 N_TE_B_M1018_g N_A_M1010_g 0.0140095f $X=6.115 $Y=0.445 $X2=0 $Y2=0
cc_475 N_TE_B_M1044_g N_A_M1010_g 0.00487788f $X=6.225 $Y=2.285 $X2=0 $Y2=0
cc_476 N_TE_B_c_394_n N_A_M1010_g 0.0139168f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_477 N_TE_B_c_395_n N_A_M1010_g 0.00337947f $X=5.9 $Y=0.995 $X2=0 $Y2=0
cc_478 N_TE_B_c_397_n N_A_M1010_g 8.71142e-19 $X=6.115 $Y=1.16 $X2=0 $Y2=0
cc_479 N_TE_B_c_398_n N_A_M1010_g 0.00685454f $X=6.115 $Y=1.16 $X2=0 $Y2=0
cc_480 N_TE_B_M1044_g N_A_c_1636_n 0.0280065f $X=6.225 $Y=2.285 $X2=0 $Y2=0
cc_481 N_TE_B_M1044_g N_A_c_1651_n 0.00894529f $X=6.225 $Y=2.285 $X2=0 $Y2=0
cc_482 N_TE_B_M1018_g N_A_1238_47#_c_1807_n 0.00706731f $X=6.115 $Y=0.445 $X2=0
+ $Y2=0
cc_483 N_TE_B_M1018_g N_A_1238_47#_c_1798_n 0.00438677f $X=6.115 $Y=0.445 $X2=0
+ $Y2=0
cc_484 N_TE_B_c_394_n N_A_1238_47#_c_1798_n 0.0140148f $X=5.815 $Y=0.73 $X2=0
+ $Y2=0
cc_485 N_TE_B_c_397_n N_A_1238_47#_c_1798_n 0.00363432f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_486 N_TE_B_c_398_n N_A_1238_47#_c_1798_n 0.00461974f $X=6.115 $Y=1.16 $X2=0
+ $Y2=0
cc_487 N_TE_B_M1044_g N_A_1238_47#_c_1805_n 0.00200968f $X=6.225 $Y=2.285 $X2=0
+ $Y2=0
cc_488 N_TE_B_M1044_g N_A_1238_47#_c_1806_n 4.74674e-19 $X=6.225 $Y=2.285 $X2=0
+ $Y2=0
cc_489 N_TE_B_M1052_g N_VPWR_c_1922_n 0.0094103f $X=0.48 $Y=2.255 $X2=0 $Y2=0
cc_490 N_TE_B_M1044_g N_VPWR_c_1926_n 0.0211184f $X=6.225 $Y=2.285 $X2=0 $Y2=0
cc_491 N_TE_B_c_397_n N_VPWR_c_1926_n 0.00554037f $X=6.115 $Y=1.16 $X2=0 $Y2=0
cc_492 N_TE_B_c_398_n N_VPWR_c_1926_n 0.00257503f $X=6.115 $Y=1.16 $X2=0 $Y2=0
cc_493 N_TE_B_M1052_g N_VPWR_c_1960_n 0.00385415f $X=0.48 $Y=2.255 $X2=0 $Y2=0
cc_494 N_TE_B_M1052_g N_VPWR_c_1921_n 0.0046122f $X=0.48 $Y=2.255 $X2=0 $Y2=0
cc_495 N_TE_B_M1044_g N_VPWR_c_1921_n 7.97988e-19 $X=6.225 $Y=2.285 $X2=0 $Y2=0
cc_496 N_TE_B_c_392_n N_VGND_M1024_s 0.0140174f $X=3.335 $Y=0.935 $X2=0 $Y2=0
cc_497 N_TE_B_c_527_p N_VGND_M1024_s 0.00491605f $X=3.42 $Y=0.85 $X2=0 $Y2=0
cc_498 N_TE_B_c_528_p N_VGND_M1024_s 0.00260983f $X=3.505 $Y=0.35 $X2=0 $Y2=0
cc_499 N_TE_B_c_467_p N_VGND_M1049_s 0.00257984f $X=4.035 $Y=0.35 $X2=0 $Y2=0
cc_500 N_TE_B_c_502_p N_VGND_M1049_s 0.00300067f $X=4.12 $Y=0.645 $X2=0 $Y2=0
cc_501 N_TE_B_c_394_n N_VGND_M1049_s 0.012805f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_502 N_TE_B_c_477_p N_VGND_M1049_s 9.936e-19 $X=4.205 $Y=0.73 $X2=0 $Y2=0
cc_503 N_TE_B_c_394_n N_VGND_M1010_s 0.01165f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_504 N_TE_B_c_395_n N_VGND_M1010_s 0.0024642f $X=5.9 $Y=0.995 $X2=0 $Y2=0
cc_505 N_TE_B_c_397_n N_VGND_M1010_s 8.11787e-19 $X=6.115 $Y=1.16 $X2=0 $Y2=0
cc_506 N_TE_B_c_376_n N_VGND_c_2515_n 0.00530389f $X=0.93 $Y=0.955 $X2=0 $Y2=0
cc_507 N_TE_B_c_387_n N_VGND_c_2515_n 0.0233617f $X=1.57 $Y=1.08 $X2=0 $Y2=0
cc_508 N_TE_B_c_390_n N_VGND_c_2515_n 0.0133632f $X=1.74 $Y=0.35 $X2=0 $Y2=0
cc_509 N_TE_B_c_380_n N_VGND_c_2516_n 0.00465534f $X=3.555 $Y=1.185 $X2=0 $Y2=0
cc_510 N_TE_B_c_391_n N_VGND_c_2516_n 0.0127796f $X=2.64 $Y=0.435 $X2=0 $Y2=0
cc_511 N_TE_B_c_435_p N_VGND_c_2516_n 0.0165658f $X=2.64 $Y=0.85 $X2=0 $Y2=0
cc_512 N_TE_B_c_392_n N_VGND_c_2516_n 0.0127692f $X=3.335 $Y=0.935 $X2=0 $Y2=0
cc_513 N_TE_B_c_527_p N_VGND_c_2516_n 0.0163238f $X=3.42 $Y=0.85 $X2=0 $Y2=0
cc_514 N_TE_B_c_528_p N_VGND_c_2516_n 0.013252f $X=3.505 $Y=0.35 $X2=0 $Y2=0
cc_515 N_TE_B_c_396_n N_VGND_c_2516_n 0.00316601f $X=2.64 $Y=0.43 $X2=0 $Y2=0
cc_516 N_TE_B_c_382_n N_VGND_c_2517_n 0.00315334f $X=3.985 $Y=1.185 $X2=0 $Y2=0
cc_517 N_TE_B_c_467_p N_VGND_c_2517_n 0.0138718f $X=4.035 $Y=0.35 $X2=0 $Y2=0
cc_518 N_TE_B_c_502_p N_VGND_c_2517_n 0.00216246f $X=4.12 $Y=0.645 $X2=0 $Y2=0
cc_519 N_TE_B_c_394_n N_VGND_c_2517_n 0.019543f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_520 N_TE_B_M1018_g N_VGND_c_2518_n 0.00538036f $X=6.115 $Y=0.445 $X2=0 $Y2=0
cc_521 N_TE_B_c_394_n N_VGND_c_2518_n 0.0240466f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_522 N_TE_B_M1018_g N_VGND_c_2519_n 0.00111032f $X=6.115 $Y=0.445 $X2=0 $Y2=0
cc_523 N_TE_B_c_394_n N_VGND_c_2529_n 0.0125599f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_524 N_TE_B_M1018_g N_VGND_c_2531_n 0.00549284f $X=6.115 $Y=0.445 $X2=0 $Y2=0
cc_525 N_TE_B_c_394_n N_VGND_c_2531_n 0.00195279f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_526 N_TE_B_c_376_n N_VGND_c_2545_n 0.00514022f $X=0.93 $Y=0.955 $X2=0 $Y2=0
cc_527 N_TE_B_c_389_n N_VGND_c_2546_n 0.0445118f $X=2.475 $Y=0.35 $X2=0 $Y2=0
cc_528 N_TE_B_c_390_n N_VGND_c_2546_n 0.0114622f $X=1.74 $Y=0.35 $X2=0 $Y2=0
cc_529 N_TE_B_c_391_n N_VGND_c_2546_n 0.0211073f $X=2.64 $Y=0.435 $X2=0 $Y2=0
cc_530 N_TE_B_c_396_n N_VGND_c_2546_n 0.00210642f $X=2.64 $Y=0.43 $X2=0 $Y2=0
cc_531 N_TE_B_c_380_n N_VGND_c_2547_n 0.0035993f $X=3.555 $Y=1.185 $X2=0 $Y2=0
cc_532 N_TE_B_c_382_n N_VGND_c_2547_n 0.0035993f $X=3.985 $Y=1.185 $X2=0 $Y2=0
cc_533 N_TE_B_c_467_p N_VGND_c_2547_n 0.0372962f $X=4.035 $Y=0.35 $X2=0 $Y2=0
cc_534 N_TE_B_c_528_p N_VGND_c_2547_n 0.00932233f $X=3.505 $Y=0.35 $X2=0 $Y2=0
cc_535 N_TE_B_c_394_n N_VGND_c_2547_n 0.00305828f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_536 N_TE_B_c_376_n N_VGND_c_2550_n 0.00528353f $X=0.93 $Y=0.955 $X2=0 $Y2=0
cc_537 N_TE_B_c_380_n N_VGND_c_2550_n 0.00682325f $X=3.555 $Y=1.185 $X2=0 $Y2=0
cc_538 N_TE_B_c_382_n N_VGND_c_2550_n 0.00612804f $X=3.985 $Y=1.185 $X2=0 $Y2=0
cc_539 N_TE_B_M1018_g N_VGND_c_2550_n 0.0109076f $X=6.115 $Y=0.445 $X2=0 $Y2=0
cc_540 N_TE_B_c_389_n N_VGND_c_2550_n 0.0274609f $X=2.475 $Y=0.35 $X2=0 $Y2=0
cc_541 N_TE_B_c_390_n N_VGND_c_2550_n 0.00657784f $X=1.74 $Y=0.35 $X2=0 $Y2=0
cc_542 N_TE_B_c_391_n N_VGND_c_2550_n 0.0125649f $X=2.64 $Y=0.435 $X2=0 $Y2=0
cc_543 N_TE_B_c_392_n N_VGND_c_2550_n 0.0129136f $X=3.335 $Y=0.935 $X2=0 $Y2=0
cc_544 N_TE_B_c_467_p N_VGND_c_2550_n 0.0250814f $X=4.035 $Y=0.35 $X2=0 $Y2=0
cc_545 N_TE_B_c_528_p N_VGND_c_2550_n 0.00646268f $X=3.505 $Y=0.35 $X2=0 $Y2=0
cc_546 N_TE_B_c_394_n N_VGND_c_2550_n 0.0335778f $X=5.815 $Y=0.73 $X2=0 $Y2=0
cc_547 N_TE_B_c_388_n A_303_85# 0.00144315f $X=1.655 $Y=0.995 $X2=-0.19
+ $Y2=-0.245
cc_548 N_A_27_367#_M1057_g N_A_217_367#_M1055_g 0.0492212f $X=1.44 $Y=0.635
+ $X2=0 $Y2=0
cc_549 N_A_27_367#_c_579_n N_A_217_367#_c_685_n 0.0146384f $X=1.875 $Y=1.64
+ $X2=0 $Y2=0
cc_550 N_A_27_367#_M1035_g N_A_217_367#_M1038_g 0.0275543f $X=1.95 $Y=2.675
+ $X2=0 $Y2=0
cc_551 N_A_27_367#_c_588_n N_A_217_367#_c_803_n 0.00215067f $X=1.01 $Y=1.715
+ $X2=0 $Y2=0
cc_552 N_A_27_367#_c_589_n N_A_217_367#_c_803_n 7.41524e-19 $X=1.44 $Y=1.715
+ $X2=0 $Y2=0
cc_553 N_A_27_367#_c_580_n N_A_217_367#_c_803_n 6.97554e-19 $X=1.515 $Y=1.64
+ $X2=0 $Y2=0
cc_554 N_A_27_367#_c_584_n N_A_217_367#_c_803_n 0.00177834f $X=1.085 $Y=1.675
+ $X2=0 $Y2=0
cc_555 N_A_27_367#_c_587_n N_A_217_367#_c_803_n 0.0207255f $X=1.25 $Y=1.51 $X2=0
+ $Y2=0
cc_556 N_A_27_367#_c_588_n N_A_217_367#_c_808_n 0.0105108f $X=1.01 $Y=1.715
+ $X2=0 $Y2=0
cc_557 N_A_27_367#_c_589_n N_A_217_367#_c_808_n 0.0119252f $X=1.44 $Y=1.715
+ $X2=0 $Y2=0
cc_558 N_A_27_367#_M1035_g N_A_217_367#_c_808_n 7.42189e-19 $X=1.95 $Y=2.675
+ $X2=0 $Y2=0
cc_559 N_A_27_367#_c_589_n N_A_217_367#_c_769_n 0.0141318f $X=1.44 $Y=1.715
+ $X2=0 $Y2=0
cc_560 N_A_27_367#_M1035_g N_A_217_367#_c_769_n 0.00463878f $X=1.95 $Y=2.675
+ $X2=0 $Y2=0
cc_561 N_A_27_367#_c_587_n N_A_217_367#_c_769_n 0.00164342f $X=1.25 $Y=1.51
+ $X2=0 $Y2=0
cc_562 N_A_27_367#_c_589_n N_A_217_367#_c_770_n 0.00462574f $X=1.44 $Y=1.715
+ $X2=0 $Y2=0
cc_563 N_A_27_367#_M1035_g N_A_217_367#_c_770_n 0.00238699f $X=1.95 $Y=2.675
+ $X2=0 $Y2=0
cc_564 N_A_27_367#_c_587_n N_A_217_367#_c_770_n 0.00276041f $X=1.25 $Y=1.51
+ $X2=0 $Y2=0
cc_565 N_A_27_367#_c_579_n N_A_217_367#_c_708_n 0.0103536f $X=1.875 $Y=1.64
+ $X2=0 $Y2=0
cc_566 N_A_27_367#_c_580_n N_A_217_367#_c_708_n 4.13742e-19 $X=1.515 $Y=1.64
+ $X2=0 $Y2=0
cc_567 N_A_27_367#_c_587_n N_A_217_367#_c_708_n 0.0126705f $X=1.25 $Y=1.51 $X2=0
+ $Y2=0
cc_568 N_A_27_367#_M1035_g N_A_217_367#_c_713_n 9.55876e-19 $X=1.95 $Y=2.675
+ $X2=0 $Y2=0
cc_569 N_A_27_367#_c_587_n N_A_217_367#_c_713_n 5.91484e-19 $X=1.25 $Y=1.51
+ $X2=0 $Y2=0
cc_570 N_A_27_367#_c_579_n N_A_217_367#_c_717_n 0.0207443f $X=1.875 $Y=1.64
+ $X2=0 $Y2=0
cc_571 N_A_27_367#_M1035_g N_A_217_367#_c_718_n 0.00165067f $X=1.95 $Y=2.675
+ $X2=0 $Y2=0
cc_572 N_A_27_367#_c_579_n N_A_217_367#_c_719_n 5.22753e-19 $X=1.875 $Y=1.64
+ $X2=0 $Y2=0
cc_573 N_A_27_367#_c_579_n N_A_217_367#_c_725_n 0.00590409f $X=1.875 $Y=1.64
+ $X2=0 $Y2=0
cc_574 N_A_27_367#_M1035_g N_A_217_367#_c_725_n 0.00602842f $X=1.95 $Y=2.675
+ $X2=0 $Y2=0
cc_575 N_A_27_367#_c_589_n N_A_381_85#_c_1224_n 2.24348e-19 $X=1.44 $Y=1.715
+ $X2=0 $Y2=0
cc_576 N_A_27_367#_M1035_g N_A_381_85#_c_1224_n 0.0102652f $X=1.95 $Y=2.675
+ $X2=0 $Y2=0
cc_577 N_A_27_367#_M1057_g N_A_381_85#_c_1190_n 0.0015948f $X=1.44 $Y=0.635
+ $X2=0 $Y2=0
cc_578 N_A_27_367#_c_587_n N_A_381_85#_c_1190_n 8.36512e-19 $X=1.25 $Y=1.51
+ $X2=0 $Y2=0
cc_579 N_A_27_367#_c_589_n N_A_381_85#_c_1200_n 4.66869e-19 $X=1.44 $Y=1.715
+ $X2=0 $Y2=0
cc_580 N_A_27_367#_M1035_g N_A_381_85#_c_1200_n 0.00559922f $X=1.95 $Y=2.675
+ $X2=0 $Y2=0
cc_581 N_A_27_367#_c_588_n N_VPWR_c_1922_n 0.00485573f $X=1.01 $Y=1.715 $X2=0
+ $Y2=0
cc_582 N_A_27_367#_c_593_n N_VPWR_c_1922_n 0.0506532f $X=0.265 $Y=1.98 $X2=0
+ $Y2=0
cc_583 N_A_27_367#_c_584_n N_VPWR_c_1922_n 0.0196257f $X=1.085 $Y=1.675 $X2=0
+ $Y2=0
cc_584 N_A_27_367#_c_589_n N_VPWR_c_1923_n 0.00349196f $X=1.44 $Y=1.715 $X2=0
+ $Y2=0
cc_585 N_A_27_367#_c_579_n N_VPWR_c_1923_n 7.09149e-19 $X=1.875 $Y=1.64 $X2=0
+ $Y2=0
cc_586 N_A_27_367#_M1035_g N_VPWR_c_1923_n 0.00714665f $X=1.95 $Y=2.675 $X2=0
+ $Y2=0
cc_587 N_A_27_367#_c_593_n N_VPWR_c_1960_n 0.00658678f $X=0.265 $Y=1.98 $X2=0
+ $Y2=0
cc_588 N_A_27_367#_c_588_n N_VPWR_c_1961_n 0.00549284f $X=1.01 $Y=1.715 $X2=0
+ $Y2=0
cc_589 N_A_27_367#_c_589_n N_VPWR_c_1961_n 0.00549284f $X=1.44 $Y=1.715 $X2=0
+ $Y2=0
cc_590 N_A_27_367#_M1035_g N_VPWR_c_1962_n 0.00549284f $X=1.95 $Y=2.675 $X2=0
+ $Y2=0
cc_591 N_A_27_367#_c_588_n N_VPWR_c_1921_n 0.0110929f $X=1.01 $Y=1.715 $X2=0
+ $Y2=0
cc_592 N_A_27_367#_c_589_n N_VPWR_c_1921_n 0.009987f $X=1.44 $Y=1.715 $X2=0
+ $Y2=0
cc_593 N_A_27_367#_M1035_g N_VPWR_c_1921_n 0.0101346f $X=1.95 $Y=2.675 $X2=0
+ $Y2=0
cc_594 N_A_27_367#_c_593_n N_VPWR_c_1921_n 0.00992454f $X=0.265 $Y=1.98 $X2=0
+ $Y2=0
cc_595 N_A_27_367#_M1057_g N_VGND_c_2515_n 0.00790149f $X=1.44 $Y=0.635 $X2=0
+ $Y2=0
cc_596 N_A_27_367#_c_586_n N_VGND_c_2515_n 0.0154542f $X=0.715 $Y=0.61 $X2=0
+ $Y2=0
cc_597 N_A_27_367#_c_582_n N_VGND_c_2545_n 0.00499037f $X=0.55 $Y=0.73 $X2=0
+ $Y2=0
cc_598 N_A_27_367#_c_583_n N_VGND_c_2545_n 0.00337272f $X=0.27 $Y=0.73 $X2=0
+ $Y2=0
cc_599 N_A_27_367#_c_586_n N_VGND_c_2545_n 0.011494f $X=0.715 $Y=0.61 $X2=0
+ $Y2=0
cc_600 N_A_27_367#_M1057_g N_VGND_c_2546_n 0.00447026f $X=1.44 $Y=0.635 $X2=0
+ $Y2=0
cc_601 N_A_27_367#_M1057_g N_VGND_c_2550_n 0.00443817f $X=1.44 $Y=0.635 $X2=0
+ $Y2=0
cc_602 N_A_27_367#_c_582_n N_VGND_c_2550_n 0.007933f $X=0.55 $Y=0.73 $X2=0 $Y2=0
cc_603 N_A_27_367#_c_583_n N_VGND_c_2550_n 0.00512101f $X=0.27 $Y=0.73 $X2=0
+ $Y2=0
cc_604 N_A_27_367#_c_586_n N_VGND_c_2550_n 0.0114702f $X=0.715 $Y=0.61 $X2=0
+ $Y2=0
cc_605 N_A_217_367#_c_712_n N_A_381_85#_c_1185_n 0.0118838f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_606 N_A_217_367#_c_712_n N_A_381_85#_c_1195_n 0.00361743f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_607 N_A_217_367#_c_712_n N_A_381_85#_c_1186_n 0.00641725f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_608 N_A_217_367#_c_712_n N_A_381_85#_c_1197_n 0.00556085f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_609 N_A_217_367#_c_712_n N_A_381_85#_c_1187_n 0.00134733f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_610 N_A_217_367#_M1055_g N_A_381_85#_c_1188_n 0.00912019f $X=1.83 $Y=0.635
+ $X2=0 $Y2=0
cc_611 N_A_217_367#_c_684_n N_A_381_85#_c_1188_n 0.00705911f $X=2.265 $Y=1.25
+ $X2=0 $Y2=0
cc_612 N_A_217_367#_M1038_g N_A_381_85#_c_1224_n 0.0161331f $X=2.38 $Y=2.675
+ $X2=0 $Y2=0
cc_613 N_A_217_367#_c_808_n N_A_381_85#_c_1224_n 8.98134e-19 $X=1.225 $Y=2.9
+ $X2=0 $Y2=0
cc_614 N_A_217_367#_c_684_n N_A_381_85#_c_1189_n 0.00949929f $X=2.265 $Y=1.25
+ $X2=0 $Y2=0
cc_615 N_A_217_367#_c_712_n N_A_381_85#_c_1189_n 0.0118074f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_616 N_A_217_367#_c_713_n N_A_381_85#_c_1189_n 0.00146502f $X=2.305 $Y=1.665
+ $X2=0 $Y2=0
cc_617 N_A_217_367#_c_717_n N_A_381_85#_c_1189_n 7.88491e-19 $X=2.4 $Y=1.74
+ $X2=0 $Y2=0
cc_618 N_A_217_367#_c_718_n N_A_381_85#_c_1189_n 0.0208595f $X=2.4 $Y=1.74 $X2=0
+ $Y2=0
cc_619 N_A_217_367#_c_719_n N_A_381_85#_c_1189_n 0.00436853f $X=2.4 $Y=1.575
+ $X2=0 $Y2=0
cc_620 N_A_217_367#_c_684_n N_A_381_85#_c_1190_n 0.00862767f $X=2.265 $Y=1.25
+ $X2=0 $Y2=0
cc_621 N_A_217_367#_c_713_n N_A_381_85#_c_1190_n 0.00650878f $X=2.305 $Y=1.665
+ $X2=0 $Y2=0
cc_622 N_A_217_367#_c_725_n N_A_381_85#_c_1190_n 0.0176716f $X=2.045 $Y=1.727
+ $X2=0 $Y2=0
cc_623 N_A_217_367#_M1038_g N_A_381_85#_c_1199_n 0.0131447f $X=2.38 $Y=2.675
+ $X2=0 $Y2=0
cc_624 N_A_217_367#_c_712_n N_A_381_85#_c_1199_n 0.0100972f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_625 N_A_217_367#_c_717_n N_A_381_85#_c_1199_n 0.00245042f $X=2.4 $Y=1.74
+ $X2=0 $Y2=0
cc_626 N_A_217_367#_c_718_n N_A_381_85#_c_1199_n 0.0154476f $X=2.4 $Y=1.74 $X2=0
+ $Y2=0
cc_627 N_A_217_367#_M1038_g N_A_381_85#_c_1200_n 0.00273924f $X=2.38 $Y=2.675
+ $X2=0 $Y2=0
cc_628 N_A_217_367#_c_808_n N_A_381_85#_c_1200_n 0.00398927f $X=1.225 $Y=2.9
+ $X2=0 $Y2=0
cc_629 N_A_217_367#_c_769_n N_A_381_85#_c_1200_n 0.0017045f $X=1.595 $Y=2.025
+ $X2=0 $Y2=0
cc_630 N_A_217_367#_c_713_n N_A_381_85#_c_1200_n 0.00242626f $X=2.305 $Y=1.665
+ $X2=0 $Y2=0
cc_631 N_A_217_367#_c_717_n N_A_381_85#_c_1200_n 0.00177873f $X=2.4 $Y=1.74
+ $X2=0 $Y2=0
cc_632 N_A_217_367#_c_718_n N_A_381_85#_c_1200_n 0.0219464f $X=2.4 $Y=1.74 $X2=0
+ $Y2=0
cc_633 N_A_217_367#_c_725_n N_A_381_85#_c_1200_n 0.00153198f $X=2.045 $Y=1.727
+ $X2=0 $Y2=0
cc_634 N_A_217_367#_M1038_g N_A_381_85#_c_1201_n 0.00551194f $X=2.38 $Y=2.675
+ $X2=0 $Y2=0
cc_635 N_A_217_367#_c_712_n N_A_381_85#_c_1191_n 0.0319293f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_636 N_A_217_367#_c_717_n N_A_381_85#_c_1191_n 5.22808e-19 $X=2.4 $Y=1.74
+ $X2=0 $Y2=0
cc_637 N_A_217_367#_c_718_n N_A_381_85#_c_1192_n 0.0190071f $X=2.4 $Y=1.74 $X2=0
+ $Y2=0
cc_638 N_A_217_367#_c_719_n N_A_381_85#_c_1192_n 0.00503139f $X=2.4 $Y=1.575
+ $X2=0 $Y2=0
cc_639 N_A_217_367#_c_712_n N_A_381_85#_c_1193_n 8.66966e-19 $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_640 N_A_217_367#_c_717_n N_A_381_85#_c_1193_n 0.0189135f $X=2.4 $Y=1.74 $X2=0
+ $Y2=0
cc_641 N_A_217_367#_c_718_n N_A_381_85#_c_1193_n 0.00123204f $X=2.4 $Y=1.74
+ $X2=0 $Y2=0
cc_642 N_A_217_367#_c_712_n N_A_726_47#_M1000_g 0.00625299f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_643 N_A_217_367#_c_697_n N_A_726_47#_c_1309_n 0.00461451f $X=13.745 $Y=1.65
+ $X2=0 $Y2=0
cc_644 N_A_217_367#_c_692_n N_A_726_47#_c_1310_n 0.131381f $X=11.595 $Y=1.65
+ $X2=0 $Y2=0
cc_645 N_A_217_367#_c_707_n N_A_726_47#_c_1310_n 0.00461451f $X=13.39 $Y=1.65
+ $X2=0 $Y2=0
cc_646 N_A_217_367#_c_716_n N_A_726_47#_c_1310_n 0.00288684f $X=16.965 $Y=1.665
+ $X2=0 $Y2=0
cc_647 N_A_217_367#_c_723_n N_A_726_47#_c_1310_n 3.5559e-19 $X=16.945 $Y=1.51
+ $X2=0 $Y2=0
cc_648 N_A_217_367#_c_720_n N_A_726_47#_c_1312_n 8.42755e-19 $X=14.025 $Y=1.51
+ $X2=0 $Y2=0
cc_649 N_A_217_367#_c_721_n N_A_726_47#_c_1316_n 8.42755e-19 $X=14.885 $Y=1.51
+ $X2=0 $Y2=0
cc_650 N_A_217_367#_c_722_n N_A_726_47#_c_1320_n 8.42755e-19 $X=15.745 $Y=1.51
+ $X2=0 $Y2=0
cc_651 N_A_217_367#_c_712_n N_A_726_47#_c_1323_n 0.0019964f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_652 N_A_217_367#_c_716_n N_A_726_47#_c_1324_n 0.00452657f $X=16.965 $Y=1.665
+ $X2=0 $Y2=0
cc_653 N_A_217_367#_c_723_n N_A_726_47#_c_1324_n 0.161543f $X=16.945 $Y=1.51
+ $X2=0 $Y2=0
cc_654 N_A_217_367#_c_712_n N_A_726_47#_c_1349_n 0.00461528f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_655 N_A_217_367#_c_712_n N_A_726_47#_c_1329_n 0.0351225f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_656 N_A_217_367#_c_712_n N_A_726_47#_c_1331_n 0.0228676f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_657 N_A_217_367#_c_712_n N_A_726_47#_c_1332_n 0.0518798f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_658 N_A_217_367#_c_712_n N_A_726_47#_c_1333_n 0.0243334f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_659 N_A_217_367#_c_698_n N_A_726_47#_c_1334_n 3.41113e-19 $X=9.52 $Y=1.65
+ $X2=0 $Y2=0
cc_660 N_A_217_367#_c_709_n N_A_726_47#_c_1334_n 0.0198902f $X=8.955 $Y=1.55
+ $X2=0 $Y2=0
cc_661 N_A_217_367#_c_710_n N_A_726_47#_c_1334_n 0.00901161f $X=8.85 $Y=0.815
+ $X2=0 $Y2=0
cc_662 N_A_217_367#_c_712_n N_A_726_47#_c_1334_n 0.18204f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_663 N_A_217_367#_c_714_n N_A_726_47#_c_1334_n 0.0341416f $X=9.33 $Y=1.665
+ $X2=0 $Y2=0
cc_664 N_A_217_367#_c_715_n N_A_726_47#_c_1334_n 0.00601005f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_665 N_A_217_367#_c_712_n N_A_726_47#_c_1335_n 0.0235513f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_666 N_A_217_367#_c_688_n N_A_726_47#_c_1336_n 0.00141799f $X=9.875 $Y=1.65
+ $X2=0 $Y2=0
cc_667 N_A_217_367#_c_709_n N_A_726_47#_c_1336_n 0.00207818f $X=8.955 $Y=1.55
+ $X2=0 $Y2=0
cc_668 N_A_217_367#_c_716_n N_A_726_47#_c_1336_n 0.367769f $X=16.965 $Y=1.665
+ $X2=0 $Y2=0
cc_669 N_A_217_367#_c_703_n N_A_726_47#_c_1337_n 0.00141799f $X=11.67 $Y=1.65
+ $X2=0 $Y2=0
cc_670 N_A_217_367#_c_712_n N_A_726_47#_c_1339_n 0.0191763f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_671 N_A_217_367#_c_698_n N_A_726_47#_c_1340_n 0.131381f $X=9.52 $Y=1.65 $X2=0
+ $Y2=0
cc_672 N_A_217_367#_c_709_n N_A_726_47#_c_1340_n 3.52385e-19 $X=8.955 $Y=1.55
+ $X2=0 $Y2=0
cc_673 N_A_217_367#_c_710_n N_A_726_47#_c_1340_n 9.57054e-19 $X=8.85 $Y=0.815
+ $X2=0 $Y2=0
cc_674 N_A_217_367#_c_716_n N_A_726_47#_c_1340_n 0.0029052f $X=16.965 $Y=1.665
+ $X2=0 $Y2=0
cc_675 N_A_217_367#_c_688_n N_A_726_47#_c_1341_n 0.00142857f $X=9.875 $Y=1.65
+ $X2=0 $Y2=0
cc_676 N_A_217_367#_c_709_n N_A_726_47#_c_1341_n 0.00494889f $X=8.955 $Y=1.55
+ $X2=0 $Y2=0
cc_677 N_A_217_367#_c_716_n N_A_726_47#_c_1341_n 8.68597e-19 $X=16.965 $Y=1.665
+ $X2=0 $Y2=0
cc_678 N_A_217_367#_c_690_n N_A_726_47#_c_1342_n 0.00329165f $X=10.735 $Y=1.65
+ $X2=0 $Y2=0
cc_679 N_A_217_367#_c_716_n N_A_726_47#_c_1342_n 0.00149426f $X=16.965 $Y=1.665
+ $X2=0 $Y2=0
cc_680 N_A_217_367#_c_692_n N_A_726_47#_c_1343_n 0.00329165f $X=11.595 $Y=1.65
+ $X2=0 $Y2=0
cc_681 N_A_217_367#_c_716_n N_A_726_47#_c_1343_n 0.00149426f $X=16.965 $Y=1.665
+ $X2=0 $Y2=0
cc_682 N_A_217_367#_c_694_n N_A_726_47#_c_1344_n 0.00329165f $X=12.455 $Y=1.65
+ $X2=0 $Y2=0
cc_683 N_A_217_367#_c_716_n N_A_726_47#_c_1344_n 0.00149426f $X=16.965 $Y=1.665
+ $X2=0 $Y2=0
cc_684 N_A_217_367#_c_696_n N_A_726_47#_c_1345_n 0.00329165f $X=13.315 $Y=1.65
+ $X2=0 $Y2=0
cc_685 N_A_217_367#_c_716_n N_A_726_47#_c_1345_n 0.00149426f $X=16.965 $Y=1.665
+ $X2=0 $Y2=0
cc_686 N_A_217_367#_c_712_n N_A_726_47#_c_1346_n 9.79329e-19 $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_687 N_A_217_367#_c_712_n N_A_M1030_g 0.00670447f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_688 N_A_217_367#_c_712_n N_A_c_1636_n 0.00450135f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_689 N_A_217_367#_c_712_n N_A_c_1637_n 0.00774925f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_690 N_A_217_367#_c_712_n N_A_c_1650_n 0.00662698f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_691 N_A_217_367#_c_913_p N_A_c_1653_n 0.00118389f $X=7.86 $Y=1.98 $X2=0 $Y2=0
cc_692 N_A_217_367#_c_772_n N_A_c_1653_n 5.07172e-19 $X=8.025 $Y=1.87 $X2=0
+ $Y2=0
cc_693 N_A_217_367#_c_712_n N_A_c_1653_n 5.21992e-19 $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_694 N_A_217_367#_c_712_n N_A_c_1638_n 0.00173802f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_695 N_A_217_367#_c_913_p N_A_c_1656_n 0.0154804f $X=7.86 $Y=1.98 $X2=0 $Y2=0
cc_696 N_A_217_367#_c_772_n N_A_c_1656_n 0.00389804f $X=8.025 $Y=1.87 $X2=0
+ $Y2=0
cc_697 N_A_217_367#_c_712_n N_A_c_1656_n 0.00552575f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_698 N_A_217_367#_c_772_n N_A_c_1641_n 0.00214316f $X=8.025 $Y=1.87 $X2=0
+ $Y2=0
cc_699 N_A_217_367#_c_712_n N_A_c_1641_n 0.00102431f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_700 N_A_217_367#_c_913_p N_A_c_1658_n 0.0197981f $X=7.86 $Y=1.98 $X2=0 $Y2=0
cc_701 N_A_217_367#_c_771_n N_A_c_1658_n 0.0131461f $X=8.87 $Y=1.87 $X2=0 $Y2=0
cc_702 N_A_217_367#_c_772_n N_A_c_1658_n 0.00132719f $X=8.025 $Y=1.87 $X2=0
+ $Y2=0
cc_703 N_A_217_367#_c_712_n N_A_c_1658_n 0.00148605f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_704 N_A_217_367#_c_712_n N_A_c_1644_n 0.00217226f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_705 N_A_217_367#_c_712_n A 0.00972116f $X=9.215 $Y=1.665 $X2=0 $Y2=0
cc_706 N_A_217_367#_c_712_n N_A_c_1645_n 0.0142287f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_707 N_A_217_367#_c_687_n N_A_1238_47#_c_1795_n 0.00729769f $X=9.165 $Y=1.65
+ $X2=0 $Y2=0
cc_708 N_A_217_367#_c_771_n N_A_1238_47#_c_1795_n 0.00384503f $X=8.87 $Y=1.87
+ $X2=0 $Y2=0
cc_709 N_A_217_367#_c_709_n N_A_1238_47#_c_1795_n 0.0118203f $X=8.955 $Y=1.55
+ $X2=0 $Y2=0
cc_710 N_A_217_367#_c_710_n N_A_1238_47#_c_1795_n 0.00637711f $X=8.85 $Y=0.815
+ $X2=0 $Y2=0
cc_711 N_A_217_367#_c_712_n N_A_1238_47#_c_1795_n 8.94762e-19 $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_712 N_A_217_367#_c_715_n N_A_1238_47#_c_1795_n 0.00202047f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_713 N_A_217_367#_c_709_n N_A_1238_47#_c_1796_n 0.00250732f $X=8.955 $Y=1.55
+ $X2=0 $Y2=0
cc_714 N_A_217_367#_c_710_n N_A_1238_47#_c_1796_n 0.00785494f $X=8.85 $Y=0.815
+ $X2=0 $Y2=0
cc_715 N_A_217_367#_c_772_n N_A_1238_47#_c_1804_n 0.00187397f $X=8.025 $Y=1.87
+ $X2=0 $Y2=0
cc_716 N_A_217_367#_c_712_n N_A_1238_47#_c_1804_n 0.0105874f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_717 N_A_217_367#_c_771_n N_A_1238_47#_c_1800_n 0.0389285f $X=8.87 $Y=1.87
+ $X2=0 $Y2=0
cc_718 N_A_217_367#_c_772_n N_A_1238_47#_c_1800_n 0.0212362f $X=8.025 $Y=1.87
+ $X2=0 $Y2=0
cc_719 N_A_217_367#_c_709_n N_A_1238_47#_c_1800_n 0.023582f $X=8.955 $Y=1.55
+ $X2=0 $Y2=0
cc_720 N_A_217_367#_c_712_n N_A_1238_47#_c_1800_n 0.0401558f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_721 N_A_217_367#_c_913_p N_A_1238_47#_c_1806_n 0.00187619f $X=7.86 $Y=1.98
+ $X2=0 $Y2=0
cc_722 N_A_217_367#_c_772_n N_A_1238_47#_c_1806_n 0.00369889f $X=8.025 $Y=1.87
+ $X2=0 $Y2=0
cc_723 N_A_217_367#_c_712_n N_A_1238_47#_c_1806_n 0.0144796f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_724 N_A_217_367#_c_712_n N_A_1238_47#_c_1801_n 0.00319242f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_725 N_A_217_367#_c_687_n N_A_1238_47#_c_1802_n 0.00113286f $X=9.165 $Y=1.65
+ $X2=0 $Y2=0
cc_726 N_A_217_367#_c_771_n N_A_1238_47#_c_1802_n 0.00591545f $X=8.87 $Y=1.87
+ $X2=0 $Y2=0
cc_727 N_A_217_367#_c_709_n N_A_1238_47#_c_1802_n 0.00174541f $X=8.955 $Y=1.55
+ $X2=0 $Y2=0
cc_728 N_A_217_367#_c_712_n N_A_1238_47#_c_1802_n 0.00345108f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_729 N_A_217_367#_c_709_n N_A_1238_47#_c_1803_n 0.00175618f $X=8.955 $Y=1.55
+ $X2=0 $Y2=0
cc_730 N_A_217_367#_c_710_n N_A_1238_47#_c_1803_n 0.00257664f $X=8.85 $Y=0.815
+ $X2=0 $Y2=0
cc_731 N_A_217_367#_c_769_n N_VPWR_M1019_s 0.00580291f $X=1.595 $Y=2.025 $X2=0
+ $Y2=0
cc_732 N_A_217_367#_c_770_n N_VPWR_M1019_s 0.00227514f $X=1.68 $Y=1.94 $X2=0
+ $Y2=0
cc_733 N_A_217_367#_c_771_n N_VPWR_M1031_s 0.0108206f $X=8.87 $Y=1.87 $X2=0
+ $Y2=0
cc_734 N_A_217_367#_c_711_n N_VPWR_M1031_s 0.00427649f $X=9.04 $Y=1.665 $X2=0
+ $Y2=0
cc_735 N_A_217_367#_c_769_n N_VPWR_c_1923_n 0.0161046f $X=1.595 $Y=2.025 $X2=0
+ $Y2=0
cc_736 N_A_217_367#_c_725_n N_VPWR_c_1923_n 0.00182541f $X=2.045 $Y=1.727 $X2=0
+ $Y2=0
cc_737 N_A_217_367#_M1038_g N_VPWR_c_1924_n 0.00449979f $X=2.38 $Y=2.675 $X2=0
+ $Y2=0
cc_738 N_A_217_367#_c_712_n N_VPWR_c_1926_n 0.0113983f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_739 N_A_217_367#_c_712_n N_VPWR_c_1927_n 0.00595261f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_740 N_A_217_367#_c_727_n N_VPWR_c_1928_n 0.0270394f $X=9.09 $Y=1.725 $X2=0
+ $Y2=0
cc_741 N_A_217_367#_c_771_n N_VPWR_c_1928_n 0.0484664f $X=8.87 $Y=1.87 $X2=0
+ $Y2=0
cc_742 N_A_217_367#_c_712_n N_VPWR_c_1928_n 0.00178515f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_743 N_A_217_367#_c_727_n N_VPWR_c_1929_n 0.00132485f $X=9.09 $Y=1.725 $X2=0
+ $Y2=0
cc_744 N_A_217_367#_c_730_n N_VPWR_c_1929_n 0.0138836f $X=9.52 $Y=1.725 $X2=0
+ $Y2=0
cc_745 N_A_217_367#_c_732_n N_VPWR_c_1929_n 0.00318602f $X=9.95 $Y=1.725 $X2=0
+ $Y2=0
cc_746 N_A_217_367#_c_734_n N_VPWR_c_1930_n 0.00315999f $X=10.38 $Y=1.725 $X2=0
+ $Y2=0
cc_747 N_A_217_367#_c_690_n N_VPWR_c_1930_n 0.0022751f $X=10.735 $Y=1.65 $X2=0
+ $Y2=0
cc_748 N_A_217_367#_c_736_n N_VPWR_c_1930_n 0.00315999f $X=10.81 $Y=1.725 $X2=0
+ $Y2=0
cc_749 N_A_217_367#_c_738_n N_VPWR_c_1931_n 0.00315999f $X=11.24 $Y=1.725 $X2=0
+ $Y2=0
cc_750 N_A_217_367#_c_692_n N_VPWR_c_1931_n 0.0022751f $X=11.595 $Y=1.65 $X2=0
+ $Y2=0
cc_751 N_A_217_367#_c_740_n N_VPWR_c_1931_n 0.00315999f $X=11.67 $Y=1.725 $X2=0
+ $Y2=0
cc_752 N_A_217_367#_c_740_n N_VPWR_c_1932_n 0.00549284f $X=11.67 $Y=1.725 $X2=0
+ $Y2=0
cc_753 N_A_217_367#_c_742_n N_VPWR_c_1932_n 0.00549284f $X=12.1 $Y=1.725 $X2=0
+ $Y2=0
cc_754 N_A_217_367#_c_742_n N_VPWR_c_1933_n 0.00315999f $X=12.1 $Y=1.725 $X2=0
+ $Y2=0
cc_755 N_A_217_367#_c_694_n N_VPWR_c_1933_n 0.0022751f $X=12.455 $Y=1.65 $X2=0
+ $Y2=0
cc_756 N_A_217_367#_c_744_n N_VPWR_c_1933_n 0.00315999f $X=12.53 $Y=1.725 $X2=0
+ $Y2=0
cc_757 N_A_217_367#_c_746_n N_VPWR_c_1934_n 0.00315999f $X=12.96 $Y=1.725 $X2=0
+ $Y2=0
cc_758 N_A_217_367#_c_696_n N_VPWR_c_1934_n 0.0022751f $X=13.315 $Y=1.65 $X2=0
+ $Y2=0
cc_759 N_A_217_367#_c_748_n N_VPWR_c_1934_n 0.00315999f $X=13.39 $Y=1.725 $X2=0
+ $Y2=0
cc_760 N_A_217_367#_c_750_n N_VPWR_c_1935_n 0.00315999f $X=13.82 $Y=1.725 $X2=0
+ $Y2=0
cc_761 N_A_217_367#_c_751_n N_VPWR_c_1935_n 0.00315999f $X=14.25 $Y=1.725 $X2=0
+ $Y2=0
cc_762 N_A_217_367#_c_720_n N_VPWR_c_1935_n 0.00309227f $X=14.025 $Y=1.51 $X2=0
+ $Y2=0
cc_763 N_A_217_367#_c_723_n N_VPWR_c_1935_n 6.2031e-19 $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_764 N_A_217_367#_c_752_n N_VPWR_c_1936_n 0.00315999f $X=14.68 $Y=1.725 $X2=0
+ $Y2=0
cc_765 N_A_217_367#_c_753_n N_VPWR_c_1936_n 0.00315999f $X=15.11 $Y=1.725 $X2=0
+ $Y2=0
cc_766 N_A_217_367#_c_721_n N_VPWR_c_1936_n 0.00309227f $X=14.885 $Y=1.51 $X2=0
+ $Y2=0
cc_767 N_A_217_367#_c_723_n N_VPWR_c_1936_n 6.2031e-19 $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_768 N_A_217_367#_c_754_n N_VPWR_c_1937_n 0.00315999f $X=15.54 $Y=1.725 $X2=0
+ $Y2=0
cc_769 N_A_217_367#_c_755_n N_VPWR_c_1937_n 0.00315999f $X=15.97 $Y=1.725 $X2=0
+ $Y2=0
cc_770 N_A_217_367#_c_722_n N_VPWR_c_1937_n 0.00309227f $X=15.745 $Y=1.51 $X2=0
+ $Y2=0
cc_771 N_A_217_367#_c_723_n N_VPWR_c_1937_n 6.2031e-19 $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_772 N_A_217_367#_c_755_n N_VPWR_c_1938_n 0.00549284f $X=15.97 $Y=1.725 $X2=0
+ $Y2=0
cc_773 N_A_217_367#_c_756_n N_VPWR_c_1938_n 0.00549284f $X=16.4 $Y=1.725 $X2=0
+ $Y2=0
cc_774 N_A_217_367#_c_756_n N_VPWR_c_1939_n 0.00315999f $X=16.4 $Y=1.725 $X2=0
+ $Y2=0
cc_775 N_A_217_367#_c_757_n N_VPWR_c_1939_n 0.00315999f $X=16.83 $Y=1.725 $X2=0
+ $Y2=0
cc_776 N_A_217_367#_c_723_n N_VPWR_c_1939_n 6.2031e-19 $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_777 N_A_217_367#_c_724_n N_VPWR_c_1939_n 0.00309227f $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_778 N_A_217_367#_c_758_n N_VPWR_c_1941_n 0.00651107f $X=17.26 $Y=1.725 $X2=0
+ $Y2=0
cc_779 N_A_217_367#_c_727_n N_VPWR_c_1946_n 0.00585385f $X=9.09 $Y=1.725 $X2=0
+ $Y2=0
cc_780 N_A_217_367#_c_730_n N_VPWR_c_1946_n 0.00486043f $X=9.52 $Y=1.725 $X2=0
+ $Y2=0
cc_781 N_A_217_367#_c_732_n N_VPWR_c_1948_n 0.00549284f $X=9.95 $Y=1.725 $X2=0
+ $Y2=0
cc_782 N_A_217_367#_c_734_n N_VPWR_c_1948_n 0.00549284f $X=10.38 $Y=1.725 $X2=0
+ $Y2=0
cc_783 N_A_217_367#_c_736_n N_VPWR_c_1950_n 0.00549284f $X=10.81 $Y=1.725 $X2=0
+ $Y2=0
cc_784 N_A_217_367#_c_738_n N_VPWR_c_1950_n 0.00549284f $X=11.24 $Y=1.725 $X2=0
+ $Y2=0
cc_785 N_A_217_367#_c_744_n N_VPWR_c_1952_n 0.00549284f $X=12.53 $Y=1.725 $X2=0
+ $Y2=0
cc_786 N_A_217_367#_c_746_n N_VPWR_c_1952_n 0.00549284f $X=12.96 $Y=1.725 $X2=0
+ $Y2=0
cc_787 N_A_217_367#_c_748_n N_VPWR_c_1954_n 0.00549284f $X=13.39 $Y=1.725 $X2=0
+ $Y2=0
cc_788 N_A_217_367#_c_750_n N_VPWR_c_1954_n 0.00549284f $X=13.82 $Y=1.725 $X2=0
+ $Y2=0
cc_789 N_A_217_367#_c_751_n N_VPWR_c_1956_n 0.00549284f $X=14.25 $Y=1.725 $X2=0
+ $Y2=0
cc_790 N_A_217_367#_c_752_n N_VPWR_c_1956_n 0.00549284f $X=14.68 $Y=1.725 $X2=0
+ $Y2=0
cc_791 N_A_217_367#_c_753_n N_VPWR_c_1958_n 0.00549284f $X=15.11 $Y=1.725 $X2=0
+ $Y2=0
cc_792 N_A_217_367#_c_754_n N_VPWR_c_1958_n 0.00549284f $X=15.54 $Y=1.725 $X2=0
+ $Y2=0
cc_793 N_A_217_367#_c_808_n N_VPWR_c_1961_n 0.0177952f $X=1.225 $Y=2.9 $X2=0
+ $Y2=0
cc_794 N_A_217_367#_M1038_g N_VPWR_c_1962_n 0.00549284f $X=2.38 $Y=2.675 $X2=0
+ $Y2=0
cc_795 N_A_217_367#_c_913_p N_VPWR_c_1964_n 0.0177952f $X=7.86 $Y=1.98 $X2=0
+ $Y2=0
cc_796 N_A_217_367#_c_757_n N_VPWR_c_1965_n 0.00549284f $X=16.83 $Y=1.725 $X2=0
+ $Y2=0
cc_797 N_A_217_367#_c_758_n N_VPWR_c_1965_n 0.00549284f $X=17.26 $Y=1.725 $X2=0
+ $Y2=0
cc_798 N_A_217_367#_M1015_d N_VPWR_c_1921_n 0.00223819f $X=1.085 $Y=1.835 $X2=0
+ $Y2=0
cc_799 N_A_217_367#_M1028_d N_VPWR_c_1921_n 0.00223819f $X=7.72 $Y=1.835 $X2=0
+ $Y2=0
cc_800 N_A_217_367#_M1038_g N_VPWR_c_1921_n 0.0111183f $X=2.38 $Y=2.675 $X2=0
+ $Y2=0
cc_801 N_A_217_367#_c_727_n N_VPWR_c_1921_n 0.0122727f $X=9.09 $Y=1.725 $X2=0
+ $Y2=0
cc_802 N_A_217_367#_c_730_n N_VPWR_c_1921_n 0.00824727f $X=9.52 $Y=1.725 $X2=0
+ $Y2=0
cc_803 N_A_217_367#_c_732_n N_VPWR_c_1921_n 0.00979325f $X=9.95 $Y=1.725 $X2=0
+ $Y2=0
cc_804 N_A_217_367#_c_734_n N_VPWR_c_1921_n 0.00979325f $X=10.38 $Y=1.725 $X2=0
+ $Y2=0
cc_805 N_A_217_367#_c_736_n N_VPWR_c_1921_n 0.00979325f $X=10.81 $Y=1.725 $X2=0
+ $Y2=0
cc_806 N_A_217_367#_c_738_n N_VPWR_c_1921_n 0.00979325f $X=11.24 $Y=1.725 $X2=0
+ $Y2=0
cc_807 N_A_217_367#_c_740_n N_VPWR_c_1921_n 0.00979325f $X=11.67 $Y=1.725 $X2=0
+ $Y2=0
cc_808 N_A_217_367#_c_742_n N_VPWR_c_1921_n 0.00979325f $X=12.1 $Y=1.725 $X2=0
+ $Y2=0
cc_809 N_A_217_367#_c_744_n N_VPWR_c_1921_n 0.00979325f $X=12.53 $Y=1.725 $X2=0
+ $Y2=0
cc_810 N_A_217_367#_c_746_n N_VPWR_c_1921_n 0.00979325f $X=12.96 $Y=1.725 $X2=0
+ $Y2=0
cc_811 N_A_217_367#_c_748_n N_VPWR_c_1921_n 0.00979325f $X=13.39 $Y=1.725 $X2=0
+ $Y2=0
cc_812 N_A_217_367#_c_750_n N_VPWR_c_1921_n 0.00979325f $X=13.82 $Y=1.725 $X2=0
+ $Y2=0
cc_813 N_A_217_367#_c_751_n N_VPWR_c_1921_n 0.00979325f $X=14.25 $Y=1.725 $X2=0
+ $Y2=0
cc_814 N_A_217_367#_c_752_n N_VPWR_c_1921_n 0.00979325f $X=14.68 $Y=1.725 $X2=0
+ $Y2=0
cc_815 N_A_217_367#_c_753_n N_VPWR_c_1921_n 0.00979325f $X=15.11 $Y=1.725 $X2=0
+ $Y2=0
cc_816 N_A_217_367#_c_754_n N_VPWR_c_1921_n 0.00979325f $X=15.54 $Y=1.725 $X2=0
+ $Y2=0
cc_817 N_A_217_367#_c_755_n N_VPWR_c_1921_n 0.00979325f $X=15.97 $Y=1.725 $X2=0
+ $Y2=0
cc_818 N_A_217_367#_c_756_n N_VPWR_c_1921_n 0.00979325f $X=16.4 $Y=1.725 $X2=0
+ $Y2=0
cc_819 N_A_217_367#_c_757_n N_VPWR_c_1921_n 0.00979325f $X=16.83 $Y=1.725 $X2=0
+ $Y2=0
cc_820 N_A_217_367#_c_758_n N_VPWR_c_1921_n 0.0107487f $X=17.26 $Y=1.725 $X2=0
+ $Y2=0
cc_821 N_A_217_367#_c_808_n N_VPWR_c_1921_n 0.0123247f $X=1.225 $Y=2.9 $X2=0
+ $Y2=0
cc_822 N_A_217_367#_c_913_p N_VPWR_c_1921_n 0.0123247f $X=7.86 $Y=1.98 $X2=0
+ $Y2=0
cc_823 N_A_217_367#_c_712_n N_A_658_367#_c_2195_n 0.00970332f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_824 N_A_217_367#_c_712_n N_A_658_367#_c_2196_n 0.0125894f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_825 N_A_217_367#_c_712_n N_A_658_367#_c_2201_n 0.0175686f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_826 N_A_217_367#_c_712_n N_A_658_367#_c_2197_n 0.010476f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_827 N_A_217_367#_c_686_n N_Z_c_2258_n 5.97954e-19 $X=9.445 $Y=1.65 $X2=0
+ $Y2=0
cc_828 N_A_217_367#_c_711_n N_Z_c_2258_n 2.13794e-19 $X=9.04 $Y=1.665 $X2=0
+ $Y2=0
cc_829 N_A_217_367#_c_714_n N_Z_c_2258_n 5.28259e-19 $X=9.33 $Y=1.665 $X2=0
+ $Y2=0
cc_830 N_A_217_367#_c_715_n N_Z_c_2258_n 0.0121334f $X=9.36 $Y=1.665 $X2=0 $Y2=0
cc_831 N_A_217_367#_c_730_n N_Z_c_2262_n 0.0107009f $X=9.52 $Y=1.725 $X2=0 $Y2=0
cc_832 N_A_217_367#_c_688_n N_Z_c_2262_n 0.00163567f $X=9.875 $Y=1.65 $X2=0
+ $Y2=0
cc_833 N_A_217_367#_c_732_n N_Z_c_2262_n 0.00988676f $X=9.95 $Y=1.725 $X2=0
+ $Y2=0
cc_834 N_A_217_367#_c_715_n N_Z_c_2262_n 0.00488282f $X=9.36 $Y=1.665 $X2=0
+ $Y2=0
cc_835 N_A_217_367#_c_716_n N_Z_c_2262_n 0.00527467f $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_836 N_A_217_367#_c_730_n N_Z_c_2250_n 0.00109027f $X=9.52 $Y=1.725 $X2=0
+ $Y2=0
cc_837 N_A_217_367#_c_732_n N_Z_c_2250_n 0.00608058f $X=9.95 $Y=1.725 $X2=0
+ $Y2=0
cc_838 N_A_217_367#_c_689_n N_Z_c_2250_n 0.0088652f $X=10.305 $Y=1.65 $X2=0
+ $Y2=0
cc_839 N_A_217_367#_c_734_n N_Z_c_2250_n 0.00573605f $X=10.38 $Y=1.725 $X2=0
+ $Y2=0
cc_840 N_A_217_367#_c_736_n N_Z_c_2250_n 6.8716e-19 $X=10.81 $Y=1.725 $X2=0
+ $Y2=0
cc_841 N_A_217_367#_c_699_n N_Z_c_2250_n 0.00326793f $X=9.95 $Y=1.65 $X2=0 $Y2=0
cc_842 N_A_217_367#_c_700_n N_Z_c_2250_n 0.00328496f $X=10.38 $Y=1.65 $X2=0
+ $Y2=0
cc_843 N_A_217_367#_c_715_n N_Z_c_2250_n 0.0034277f $X=9.36 $Y=1.665 $X2=0 $Y2=0
cc_844 N_A_217_367#_c_716_n N_Z_c_2250_n 0.0268554f $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_845 N_A_217_367#_c_730_n N_Z_c_2276_n 7.53173e-19 $X=9.52 $Y=1.725 $X2=0
+ $Y2=0
cc_846 N_A_217_367#_c_732_n N_Z_c_2276_n 0.0114517f $X=9.95 $Y=1.725 $X2=0 $Y2=0
cc_847 N_A_217_367#_c_734_n N_Z_c_2276_n 0.0110869f $X=10.38 $Y=1.725 $X2=0
+ $Y2=0
cc_848 N_A_217_367#_c_736_n N_Z_c_2276_n 6.42028e-19 $X=10.81 $Y=1.725 $X2=0
+ $Y2=0
cc_849 N_A_217_367#_c_734_n N_Z_c_2251_n 0.00191943f $X=10.38 $Y=1.725 $X2=0
+ $Y2=0
cc_850 N_A_217_367#_c_736_n N_Z_c_2251_n 0.0191846f $X=10.81 $Y=1.725 $X2=0
+ $Y2=0
cc_851 N_A_217_367#_c_691_n N_Z_c_2251_n 0.0088652f $X=11.165 $Y=1.65 $X2=0
+ $Y2=0
cc_852 N_A_217_367#_c_738_n N_Z_c_2251_n 0.0191874f $X=11.24 $Y=1.725 $X2=0
+ $Y2=0
cc_853 N_A_217_367#_c_740_n N_Z_c_2251_n 0.00191994f $X=11.67 $Y=1.725 $X2=0
+ $Y2=0
cc_854 N_A_217_367#_c_701_n N_Z_c_2251_n 0.00328496f $X=10.81 $Y=1.65 $X2=0
+ $Y2=0
cc_855 N_A_217_367#_c_702_n N_Z_c_2251_n 0.00328496f $X=11.24 $Y=1.65 $X2=0
+ $Y2=0
cc_856 N_A_217_367#_c_716_n N_Z_c_2251_n 0.0269783f $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_857 N_A_217_367#_c_738_n N_Z_c_2252_n 0.00191994f $X=11.24 $Y=1.725 $X2=0
+ $Y2=0
cc_858 N_A_217_367#_c_740_n N_Z_c_2252_n 0.0191874f $X=11.67 $Y=1.725 $X2=0
+ $Y2=0
cc_859 N_A_217_367#_c_693_n N_Z_c_2252_n 0.0088652f $X=12.025 $Y=1.65 $X2=0
+ $Y2=0
cc_860 N_A_217_367#_c_742_n N_Z_c_2252_n 0.0191874f $X=12.1 $Y=1.725 $X2=0 $Y2=0
cc_861 N_A_217_367#_c_744_n N_Z_c_2252_n 0.00191994f $X=12.53 $Y=1.725 $X2=0
+ $Y2=0
cc_862 N_A_217_367#_c_703_n N_Z_c_2252_n 0.00328496f $X=11.67 $Y=1.65 $X2=0
+ $Y2=0
cc_863 N_A_217_367#_c_704_n N_Z_c_2252_n 0.00328496f $X=12.1 $Y=1.65 $X2=0 $Y2=0
cc_864 N_A_217_367#_c_716_n N_Z_c_2252_n 0.0269783f $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_865 N_A_217_367#_c_742_n N_Z_c_2253_n 0.00191994f $X=12.1 $Y=1.725 $X2=0
+ $Y2=0
cc_866 N_A_217_367#_c_744_n N_Z_c_2253_n 0.0191874f $X=12.53 $Y=1.725 $X2=0
+ $Y2=0
cc_867 N_A_217_367#_c_695_n N_Z_c_2253_n 0.0088652f $X=12.885 $Y=1.65 $X2=0
+ $Y2=0
cc_868 N_A_217_367#_c_746_n N_Z_c_2253_n 0.0191874f $X=12.96 $Y=1.725 $X2=0
+ $Y2=0
cc_869 N_A_217_367#_c_748_n N_Z_c_2253_n 0.00191994f $X=13.39 $Y=1.725 $X2=0
+ $Y2=0
cc_870 N_A_217_367#_c_705_n N_Z_c_2253_n 0.00328496f $X=12.53 $Y=1.65 $X2=0
+ $Y2=0
cc_871 N_A_217_367#_c_706_n N_Z_c_2253_n 0.00328496f $X=12.96 $Y=1.65 $X2=0
+ $Y2=0
cc_872 N_A_217_367#_c_716_n N_Z_c_2253_n 0.0269783f $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_873 N_A_217_367#_c_746_n N_Z_c_2254_n 0.00191994f $X=12.96 $Y=1.725 $X2=0
+ $Y2=0
cc_874 N_A_217_367#_c_748_n N_Z_c_2254_n 0.0191874f $X=13.39 $Y=1.725 $X2=0
+ $Y2=0
cc_875 N_A_217_367#_c_697_n N_Z_c_2254_n 0.0109356f $X=13.745 $Y=1.65 $X2=0
+ $Y2=0
cc_876 N_A_217_367#_c_750_n N_Z_c_2254_n 0.0189797f $X=13.82 $Y=1.725 $X2=0
+ $Y2=0
cc_877 N_A_217_367#_c_751_n N_Z_c_2254_n 0.00182938f $X=14.25 $Y=1.725 $X2=0
+ $Y2=0
cc_878 N_A_217_367#_c_707_n N_Z_c_2254_n 0.00346539f $X=13.39 $Y=1.65 $X2=0
+ $Y2=0
cc_879 N_A_217_367#_c_716_n N_Z_c_2254_n 0.0295962f $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_880 N_A_217_367#_c_720_n N_Z_c_2254_n 0.0293538f $X=14.025 $Y=1.51 $X2=0
+ $Y2=0
cc_881 N_A_217_367#_c_723_n N_Z_c_2254_n 0.00807773f $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_882 N_A_217_367#_c_750_n N_Z_c_2255_n 0.00182938f $X=13.82 $Y=1.725 $X2=0
+ $Y2=0
cc_883 N_A_217_367#_c_751_n N_Z_c_2255_n 0.0189797f $X=14.25 $Y=1.725 $X2=0
+ $Y2=0
cc_884 N_A_217_367#_c_752_n N_Z_c_2255_n 0.0189797f $X=14.68 $Y=1.725 $X2=0
+ $Y2=0
cc_885 N_A_217_367#_c_753_n N_Z_c_2255_n 0.00182938f $X=15.11 $Y=1.725 $X2=0
+ $Y2=0
cc_886 N_A_217_367#_c_716_n N_Z_c_2255_n 0.0270023f $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_887 N_A_217_367#_c_720_n N_Z_c_2255_n 0.0285366f $X=14.025 $Y=1.51 $X2=0
+ $Y2=0
cc_888 N_A_217_367#_c_721_n N_Z_c_2255_n 0.0285366f $X=14.885 $Y=1.51 $X2=0
+ $Y2=0
cc_889 N_A_217_367#_c_723_n N_Z_c_2255_n 0.0256227f $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_890 N_A_217_367#_c_752_n N_Z_c_2256_n 0.00182938f $X=14.68 $Y=1.725 $X2=0
+ $Y2=0
cc_891 N_A_217_367#_c_753_n N_Z_c_2256_n 0.0189797f $X=15.11 $Y=1.725 $X2=0
+ $Y2=0
cc_892 N_A_217_367#_c_754_n N_Z_c_2256_n 0.0189797f $X=15.54 $Y=1.725 $X2=0
+ $Y2=0
cc_893 N_A_217_367#_c_755_n N_Z_c_2256_n 0.00182938f $X=15.97 $Y=1.725 $X2=0
+ $Y2=0
cc_894 N_A_217_367#_c_716_n N_Z_c_2256_n 0.0270023f $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_895 N_A_217_367#_c_721_n N_Z_c_2256_n 0.0285366f $X=14.885 $Y=1.51 $X2=0
+ $Y2=0
cc_896 N_A_217_367#_c_722_n N_Z_c_2256_n 0.0285366f $X=15.745 $Y=1.51 $X2=0
+ $Y2=0
cc_897 N_A_217_367#_c_723_n N_Z_c_2256_n 0.0256227f $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_898 N_A_217_367#_c_754_n N_Z_c_2257_n 0.00182938f $X=15.54 $Y=1.725 $X2=0
+ $Y2=0
cc_899 N_A_217_367#_c_755_n N_Z_c_2257_n 0.0189797f $X=15.97 $Y=1.725 $X2=0
+ $Y2=0
cc_900 N_A_217_367#_c_756_n N_Z_c_2257_n 0.019433f $X=16.4 $Y=1.725 $X2=0 $Y2=0
cc_901 N_A_217_367#_c_757_n N_Z_c_2257_n 0.00229336f $X=16.83 $Y=1.725 $X2=0
+ $Y2=0
cc_902 N_A_217_367#_c_716_n N_Z_c_2257_n 0.0352521f $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_903 N_A_217_367#_c_722_n N_Z_c_2257_n 0.0285366f $X=15.745 $Y=1.51 $X2=0
+ $Y2=0
cc_904 N_A_217_367#_c_723_n N_Z_c_2257_n 0.0304401f $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_905 N_A_217_367#_c_724_n N_Z_c_2257_n 0.0299743f $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_906 N_A_217_367#_c_756_n N_Z_c_2337_n 0.0012636f $X=16.4 $Y=1.725 $X2=0 $Y2=0
cc_907 N_A_217_367#_c_757_n N_Z_c_2337_n 0.0137496f $X=16.83 $Y=1.725 $X2=0
+ $Y2=0
cc_908 N_A_217_367#_c_758_n N_Z_c_2337_n 0.0249539f $X=17.26 $Y=1.725 $X2=0
+ $Y2=0
cc_909 N_A_217_367#_c_716_n N_Z_c_2337_n 7.67524e-19 $X=16.965 $Y=1.665 $X2=0
+ $Y2=0
cc_910 N_A_217_367#_c_723_n N_Z_c_2337_n 6.13936e-19 $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_911 N_A_217_367#_c_724_n N_Z_c_2337_n 0.0145361f $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_912 N_A_217_367#_c_727_n N_Z_c_2343_n 0.0077292f $X=9.09 $Y=1.725 $X2=0 $Y2=0
cc_913 N_A_217_367#_c_730_n N_Z_c_2343_n 0.00712149f $X=9.52 $Y=1.725 $X2=0
+ $Y2=0
cc_914 N_A_217_367#_c_688_n N_Z_c_2343_n 4.88914e-19 $X=9.875 $Y=1.65 $X2=0
+ $Y2=0
cc_915 N_A_217_367#_c_732_n N_Z_c_2343_n 0.00673785f $X=9.95 $Y=1.725 $X2=0
+ $Y2=0
cc_916 N_A_217_367#_c_734_n N_Z_c_2343_n 0.00810924f $X=10.38 $Y=1.725 $X2=0
+ $Y2=0
cc_917 N_A_217_367#_c_690_n N_Z_c_2343_n 4.88914e-19 $X=10.735 $Y=1.65 $X2=0
+ $Y2=0
cc_918 N_A_217_367#_c_736_n N_Z_c_2343_n 0.00811955f $X=10.81 $Y=1.725 $X2=0
+ $Y2=0
cc_919 N_A_217_367#_c_738_n N_Z_c_2343_n 0.00811955f $X=11.24 $Y=1.725 $X2=0
+ $Y2=0
cc_920 N_A_217_367#_c_692_n N_Z_c_2343_n 4.88914e-19 $X=11.595 $Y=1.65 $X2=0
+ $Y2=0
cc_921 N_A_217_367#_c_740_n N_Z_c_2343_n 0.00811955f $X=11.67 $Y=1.725 $X2=0
+ $Y2=0
cc_922 N_A_217_367#_c_742_n N_Z_c_2343_n 0.00811955f $X=12.1 $Y=1.725 $X2=0
+ $Y2=0
cc_923 N_A_217_367#_c_694_n N_Z_c_2343_n 4.88914e-19 $X=12.455 $Y=1.65 $X2=0
+ $Y2=0
cc_924 N_A_217_367#_c_744_n N_Z_c_2343_n 0.00811955f $X=12.53 $Y=1.725 $X2=0
+ $Y2=0
cc_925 N_A_217_367#_c_746_n N_Z_c_2343_n 0.00811955f $X=12.96 $Y=1.725 $X2=0
+ $Y2=0
cc_926 N_A_217_367#_c_696_n N_Z_c_2343_n 4.88914e-19 $X=13.315 $Y=1.65 $X2=0
+ $Y2=0
cc_927 N_A_217_367#_c_748_n N_Z_c_2343_n 0.00818091f $X=13.39 $Y=1.725 $X2=0
+ $Y2=0
cc_928 N_A_217_367#_c_750_n N_Z_c_2343_n 0.00820452f $X=13.82 $Y=1.725 $X2=0
+ $Y2=0
cc_929 N_A_217_367#_c_751_n N_Z_c_2343_n 0.00820452f $X=14.25 $Y=1.725 $X2=0
+ $Y2=0
cc_930 N_A_217_367#_c_752_n N_Z_c_2343_n 0.00820452f $X=14.68 $Y=1.725 $X2=0
+ $Y2=0
cc_931 N_A_217_367#_c_753_n N_Z_c_2343_n 0.00820452f $X=15.11 $Y=1.725 $X2=0
+ $Y2=0
cc_932 N_A_217_367#_c_754_n N_Z_c_2343_n 0.00820452f $X=15.54 $Y=1.725 $X2=0
+ $Y2=0
cc_933 N_A_217_367#_c_755_n N_Z_c_2343_n 0.00820452f $X=15.97 $Y=1.725 $X2=0
+ $Y2=0
cc_934 N_A_217_367#_c_756_n N_Z_c_2343_n 0.00820452f $X=16.4 $Y=1.725 $X2=0
+ $Y2=0
cc_935 N_A_217_367#_c_757_n N_Z_c_2343_n 0.00789246f $X=16.83 $Y=1.725 $X2=0
+ $Y2=0
cc_936 N_A_217_367#_c_758_n N_Z_c_2343_n 8.0075e-19 $X=17.26 $Y=1.725 $X2=0
+ $Y2=0
cc_937 N_A_217_367#_c_711_n N_Z_c_2343_n 0.00160508f $X=9.04 $Y=1.665 $X2=0
+ $Y2=0
cc_938 N_A_217_367#_c_712_n N_Z_c_2343_n 0.00456213f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_939 N_A_217_367#_c_714_n N_Z_c_2343_n 0.782868f $X=9.33 $Y=1.665 $X2=0 $Y2=0
cc_940 N_A_217_367#_c_715_n N_Z_c_2343_n 0.00249498f $X=9.36 $Y=1.665 $X2=0
+ $Y2=0
cc_941 N_A_217_367#_c_720_n N_Z_c_2343_n 8.62013e-19 $X=14.025 $Y=1.51 $X2=0
+ $Y2=0
cc_942 N_A_217_367#_c_721_n N_Z_c_2343_n 8.62013e-19 $X=14.885 $Y=1.51 $X2=0
+ $Y2=0
cc_943 N_A_217_367#_c_722_n N_Z_c_2343_n 8.62013e-19 $X=15.745 $Y=1.51 $X2=0
+ $Y2=0
cc_944 N_A_217_367#_c_724_n N_Z_c_2343_n 0.00404212f $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_945 N_A_217_367#_c_732_n N_Z_c_2376_n 4.0679e-19 $X=9.95 $Y=1.725 $X2=0 $Y2=0
cc_946 N_A_217_367#_c_734_n N_Z_c_2376_n 0.0023483f $X=10.38 $Y=1.725 $X2=0
+ $Y2=0
cc_947 N_A_217_367#_c_736_n N_Z_c_2376_n 6.12528e-19 $X=10.81 $Y=1.725 $X2=0
+ $Y2=0
cc_948 N_A_217_367#_M1055_g N_VGND_c_2515_n 2.363e-19 $X=1.83 $Y=0.635 $X2=0
+ $Y2=0
cc_949 N_A_217_367#_c_720_n N_VGND_c_2526_n 0.00626246f $X=14.025 $Y=1.51 $X2=0
+ $Y2=0
cc_950 N_A_217_367#_c_723_n N_VGND_c_2526_n 3.37033e-19 $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_951 N_A_217_367#_c_721_n N_VGND_c_2527_n 0.00626246f $X=14.885 $Y=1.51 $X2=0
+ $Y2=0
cc_952 N_A_217_367#_c_723_n N_VGND_c_2527_n 3.37033e-19 $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_953 N_A_217_367#_c_722_n N_VGND_c_2528_n 0.00626246f $X=15.745 $Y=1.51 $X2=0
+ $Y2=0
cc_954 N_A_217_367#_c_723_n N_VGND_c_2528_n 3.37033e-19 $X=16.945 $Y=1.51 $X2=0
+ $Y2=0
cc_955 N_A_217_367#_M1055_g N_VGND_c_2546_n 8.76173e-19 $X=1.83 $Y=0.635 $X2=0
+ $Y2=0
cc_956 N_A_217_367#_M1020_d N_VGND_c_2550_n 0.00289884f $X=8.63 $Y=0.235 $X2=0
+ $Y2=0
cc_957 N_A_217_367#_c_710_n N_A_1451_47#_c_2757_n 0.00760908f $X=8.85 $Y=0.815
+ $X2=0 $Y2=0
cc_958 N_A_217_367#_M1020_d N_A_1451_47#_c_2762_n 0.00503991f $X=8.63 $Y=0.235
+ $X2=0 $Y2=0
cc_959 N_A_217_367#_c_710_n N_A_1451_47#_c_2762_n 0.0208392f $X=8.85 $Y=0.815
+ $X2=0 $Y2=0
cc_960 N_A_217_367#_c_686_n N_A_1451_47#_c_2760_n 0.00162515f $X=9.445 $Y=1.65
+ $X2=0 $Y2=0
cc_961 N_A_217_367#_c_710_n N_A_1451_47#_c_2760_n 0.0351247f $X=8.85 $Y=0.815
+ $X2=0 $Y2=0
cc_962 N_A_217_367#_c_715_n N_A_1451_47#_c_2760_n 0.00580564f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_963 N_A_381_85#_c_1195_n N_A_726_47#_c_1349_n 0.00211934f $X=3.675 $Y=1.725
+ $X2=0 $Y2=0
cc_964 N_A_381_85#_c_1186_n N_A_726_47#_c_1349_n 0.00227601f $X=4.03 $Y=1.65
+ $X2=0 $Y2=0
cc_965 N_A_381_85#_c_1197_n N_A_726_47#_c_1349_n 9.04627e-19 $X=4.105 $Y=1.725
+ $X2=0 $Y2=0
cc_966 N_A_381_85#_c_1195_n N_A_726_47#_c_1434_n 0.0128321f $X=3.675 $Y=1.725
+ $X2=0 $Y2=0
cc_967 N_A_381_85#_c_1186_n N_A_726_47#_c_1329_n 0.0046664f $X=4.03 $Y=1.65
+ $X2=0 $Y2=0
cc_968 N_A_381_85#_c_1195_n N_A_726_47#_c_1331_n 0.00239164f $X=3.675 $Y=1.725
+ $X2=0 $Y2=0
cc_969 N_A_381_85#_c_1186_n N_A_726_47#_c_1331_n 0.00609215f $X=4.03 $Y=1.65
+ $X2=0 $Y2=0
cc_970 N_A_381_85#_c_1197_n N_A_726_47#_c_1331_n 0.00178591f $X=4.105 $Y=1.725
+ $X2=0 $Y2=0
cc_971 N_A_381_85#_c_1187_n N_A_726_47#_c_1331_n 0.00451524f $X=3.675 $Y=1.65
+ $X2=0 $Y2=0
cc_972 N_A_381_85#_c_1191_n N_A_726_47#_c_1331_n 0.00444864f $X=2.965 $Y=1.74
+ $X2=0 $Y2=0
cc_973 N_A_381_85#_c_1193_n N_A_726_47#_c_1331_n 3.49759e-19 $X=2.965 $Y=1.65
+ $X2=0 $Y2=0
cc_974 N_A_381_85#_c_1186_n N_A_M1030_g 0.033066f $X=4.03 $Y=1.65 $X2=0 $Y2=0
cc_975 N_A_381_85#_c_1199_n N_VPWR_c_1924_n 0.0196868f $X=2.8 $Y=2.17 $X2=0
+ $Y2=0
cc_976 N_A_381_85#_c_1197_n N_VPWR_c_1925_n 0.00110621f $X=4.105 $Y=1.725 $X2=0
+ $Y2=0
cc_977 N_A_381_85#_c_1195_n N_VPWR_c_1942_n 0.00359964f $X=3.675 $Y=1.725 $X2=0
+ $Y2=0
cc_978 N_A_381_85#_c_1197_n N_VPWR_c_1942_n 0.0035993f $X=4.105 $Y=1.725 $X2=0
+ $Y2=0
cc_979 N_A_381_85#_c_1224_n N_VPWR_c_1962_n 0.0177952f $X=2.165 $Y=2.4 $X2=0
+ $Y2=0
cc_980 N_A_381_85#_M1035_d N_VPWR_c_1921_n 0.00223819f $X=2.025 $Y=2.255 $X2=0
+ $Y2=0
cc_981 N_A_381_85#_c_1195_n N_VPWR_c_1921_n 0.00665257f $X=3.675 $Y=1.725 $X2=0
+ $Y2=0
cc_982 N_A_381_85#_c_1197_n N_VPWR_c_1921_n 0.00555902f $X=4.105 $Y=1.725 $X2=0
+ $Y2=0
cc_983 N_A_381_85#_c_1224_n N_VPWR_c_1921_n 0.0123247f $X=2.165 $Y=2.4 $X2=0
+ $Y2=0
cc_984 N_A_381_85#_c_1185_n N_A_658_367#_c_2195_n 0.0070413f $X=3.6 $Y=1.65
+ $X2=0 $Y2=0
cc_985 N_A_381_85#_c_1195_n N_A_658_367#_c_2195_n 0.00654151f $X=3.675 $Y=1.725
+ $X2=0 $Y2=0
cc_986 N_A_381_85#_c_1199_n N_A_658_367#_c_2195_n 0.0123436f $X=2.8 $Y=2.17
+ $X2=0 $Y2=0
cc_987 N_A_381_85#_c_1201_n N_A_658_367#_c_2195_n 0.0180063f $X=2.965 $Y=2.085
+ $X2=0 $Y2=0
cc_988 N_A_381_85#_c_1193_n N_A_658_367#_c_2195_n 7.45713e-19 $X=2.965 $Y=1.65
+ $X2=0 $Y2=0
cc_989 N_A_381_85#_c_1195_n N_A_658_367#_c_2208_n 0.0103737f $X=3.675 $Y=1.725
+ $X2=0 $Y2=0
cc_990 N_A_381_85#_c_1197_n N_A_658_367#_c_2208_n 0.011131f $X=4.105 $Y=1.725
+ $X2=0 $Y2=0
cc_991 N_A_381_85#_c_1195_n N_A_658_367#_c_2196_n 2.32852e-19 $X=3.675 $Y=1.725
+ $X2=0 $Y2=0
cc_992 N_A_381_85#_c_1197_n N_A_658_367#_c_2196_n 0.00686207f $X=4.105 $Y=1.725
+ $X2=0 $Y2=0
cc_993 N_A_381_85#_c_1195_n N_A_658_367#_c_2212_n 4.89844e-19 $X=3.675 $Y=1.725
+ $X2=0 $Y2=0
cc_994 N_A_381_85#_c_1197_n N_A_658_367#_c_2212_n 0.00652175f $X=4.105 $Y=1.725
+ $X2=0 $Y2=0
cc_995 N_A_381_85#_c_1197_n N_A_658_367#_c_2214_n 0.0017646f $X=4.105 $Y=1.725
+ $X2=0 $Y2=0
cc_996 N_A_726_47#_c_1331_n N_A_M1030_g 6.59265e-19 $X=3.83 $Y=1.815 $X2=0 $Y2=0
cc_997 N_A_726_47#_c_1329_n N_A_M1001_g 0.0137524f $X=5.435 $Y=1.08 $X2=0 $Y2=0
cc_998 N_A_726_47#_c_1333_n N_A_M1001_g 7.96608e-19 $X=5.665 $Y=1.295 $X2=0
+ $Y2=0
cc_999 N_A_726_47#_c_1346_n N_A_M1001_g 0.00127553f $X=5.535 $Y=1.08 $X2=0 $Y2=0
cc_1000 N_A_726_47#_c_1329_n N_A_M1010_g 0.00881192f $X=5.435 $Y=1.08 $X2=0
+ $Y2=0
cc_1001 N_A_726_47#_c_1333_n N_A_M1010_g 0.0035967f $X=5.665 $Y=1.295 $X2=0
+ $Y2=0
cc_1002 N_A_726_47#_c_1346_n N_A_M1010_g 0.00961967f $X=5.535 $Y=1.08 $X2=0
+ $Y2=0
cc_1003 N_A_726_47#_c_1332_n N_A_c_1636_n 0.00233995f $X=6.335 $Y=1.295 $X2=0
+ $Y2=0
cc_1004 N_A_726_47#_c_1333_n N_A_c_1636_n 5.78457e-19 $X=5.665 $Y=1.295 $X2=0
+ $Y2=0
cc_1005 N_A_726_47#_c_1346_n N_A_c_1636_n 0.00474286f $X=5.535 $Y=1.08 $X2=0
+ $Y2=0
cc_1006 N_A_726_47#_c_1329_n N_A_c_1637_n 0.008222f $X=5.435 $Y=1.08 $X2=0 $Y2=0
cc_1007 N_A_726_47#_c_1331_n N_A_c_1637_n 0.00526769f $X=3.83 $Y=1.815 $X2=0
+ $Y2=0
cc_1008 N_A_726_47#_c_1333_n N_A_c_1637_n 0.00129767f $X=5.665 $Y=1.295 $X2=0
+ $Y2=0
cc_1009 N_A_726_47#_c_1346_n N_A_c_1637_n 0.0021141f $X=5.535 $Y=1.08 $X2=0
+ $Y2=0
cc_1010 N_A_726_47#_M1000_g N_A_c_1651_n 0.00895007f $X=6.615 $Y=2.285 $X2=0
+ $Y2=0
cc_1011 N_A_726_47#_M1000_g N_A_c_1639_n 0.0242154f $X=6.615 $Y=2.285 $X2=0
+ $Y2=0
cc_1012 N_A_726_47#_c_1323_n N_A_c_1639_n 0.00586958f $X=6.675 $Y=1.665 $X2=0
+ $Y2=0
cc_1013 N_A_726_47#_c_1334_n N_A_M1002_g 0.00219247f $X=9.6 $Y=1.295 $X2=0 $Y2=0
cc_1014 N_A_726_47#_c_1338_n N_A_M1002_g 0.00574551f $X=6.675 $Y=1.16 $X2=0
+ $Y2=0
cc_1015 N_A_726_47#_c_1339_n N_A_M1002_g 2.52198e-19 $X=6.675 $Y=1.16 $X2=0
+ $Y2=0
cc_1016 N_A_726_47#_c_1334_n N_A_M1003_g 0.00188514f $X=9.6 $Y=1.295 $X2=0 $Y2=0
cc_1017 N_A_726_47#_c_1329_n N_A_c_1645_n 0.0231539f $X=5.435 $Y=1.08 $X2=0
+ $Y2=0
cc_1018 N_A_726_47#_c_1333_n N_A_c_1645_n 0.00181362f $X=5.665 $Y=1.295 $X2=0
+ $Y2=0
cc_1019 N_A_726_47#_c_1346_n N_A_c_1645_n 0.00378732f $X=5.535 $Y=1.08 $X2=0
+ $Y2=0
cc_1020 N_A_726_47#_c_1334_n N_A_1238_47#_c_1795_n 0.00791514f $X=9.6 $Y=1.295
+ $X2=0 $Y2=0
cc_1021 N_A_726_47#_c_1336_n N_A_1238_47#_c_1796_n 2.66194e-19 $X=9.715 $Y=1.295
+ $X2=0 $Y2=0
cc_1022 N_A_726_47#_c_1340_n N_A_1238_47#_c_1796_n 0.00927611f $X=10.305 $Y=1.2
+ $X2=0 $Y2=0
cc_1023 N_A_726_47#_c_1341_n N_A_1238_47#_c_1796_n 8.69935e-19 $X=9.745 $Y=1.2
+ $X2=0 $Y2=0
cc_1024 N_A_726_47#_M1011_g N_A_1238_47#_c_1797_n 0.0139025f $X=6.615 $Y=0.445
+ $X2=0 $Y2=0
cc_1025 N_A_726_47#_c_1334_n N_A_1238_47#_c_1797_n 0.00743058f $X=9.6 $Y=1.295
+ $X2=0 $Y2=0
cc_1026 N_A_726_47#_c_1335_n N_A_1238_47#_c_1797_n 6.0814e-19 $X=6.625 $Y=1.295
+ $X2=0 $Y2=0
cc_1027 N_A_726_47#_c_1338_n N_A_1238_47#_c_1797_n 0.00464128f $X=6.675 $Y=1.16
+ $X2=0 $Y2=0
cc_1028 N_A_726_47#_c_1339_n N_A_1238_47#_c_1797_n 0.0243351f $X=6.675 $Y=1.16
+ $X2=0 $Y2=0
cc_1029 N_A_726_47#_c_1332_n N_A_1238_47#_c_1798_n 0.00482518f $X=6.335 $Y=1.295
+ $X2=0 $Y2=0
cc_1030 N_A_726_47#_c_1335_n N_A_1238_47#_c_1798_n 0.00321557f $X=6.625 $Y=1.295
+ $X2=0 $Y2=0
cc_1031 N_A_726_47#_c_1339_n N_A_1238_47#_c_1798_n 0.00826268f $X=6.675 $Y=1.16
+ $X2=0 $Y2=0
cc_1032 N_A_726_47#_M1011_g N_A_1238_47#_c_1799_n 0.00516777f $X=6.615 $Y=0.445
+ $X2=0 $Y2=0
cc_1033 N_A_726_47#_c_1334_n N_A_1238_47#_c_1799_n 0.0120843f $X=9.6 $Y=1.295
+ $X2=0 $Y2=0
cc_1034 N_A_726_47#_c_1335_n N_A_1238_47#_c_1799_n 2.08724e-19 $X=6.625 $Y=1.295
+ $X2=0 $Y2=0
cc_1035 N_A_726_47#_c_1338_n N_A_1238_47#_c_1799_n 0.00115281f $X=6.675 $Y=1.16
+ $X2=0 $Y2=0
cc_1036 N_A_726_47#_c_1339_n N_A_1238_47#_c_1799_n 0.0199078f $X=6.675 $Y=1.16
+ $X2=0 $Y2=0
cc_1037 N_A_726_47#_M1000_g N_A_1238_47#_c_1804_n 0.00282137f $X=6.615 $Y=2.285
+ $X2=0 $Y2=0
cc_1038 N_A_726_47#_c_1339_n N_A_1238_47#_c_1804_n 0.00376523f $X=6.675 $Y=1.16
+ $X2=0 $Y2=0
cc_1039 N_A_726_47#_c_1334_n N_A_1238_47#_c_1800_n 0.0505095f $X=9.6 $Y=1.295
+ $X2=0 $Y2=0
cc_1040 N_A_726_47#_M1000_g N_A_1238_47#_c_1805_n 0.0143753f $X=6.615 $Y=2.285
+ $X2=0 $Y2=0
cc_1041 N_A_726_47#_M1000_g N_A_1238_47#_c_1806_n 0.00345929f $X=6.615 $Y=2.285
+ $X2=0 $Y2=0
cc_1042 N_A_726_47#_c_1323_n N_A_1238_47#_c_1806_n 0.00272372f $X=6.675 $Y=1.665
+ $X2=0 $Y2=0
cc_1043 N_A_726_47#_c_1339_n N_A_1238_47#_c_1806_n 0.0101998f $X=6.675 $Y=1.16
+ $X2=0 $Y2=0
cc_1044 N_A_726_47#_c_1322_n N_A_1238_47#_c_1801_n 0.00154624f $X=6.675 $Y=1.5
+ $X2=0 $Y2=0
cc_1045 N_A_726_47#_c_1334_n N_A_1238_47#_c_1801_n 0.00542805f $X=9.6 $Y=1.295
+ $X2=0 $Y2=0
cc_1046 N_A_726_47#_c_1335_n N_A_1238_47#_c_1801_n 2.37276e-19 $X=6.625 $Y=1.295
+ $X2=0 $Y2=0
cc_1047 N_A_726_47#_c_1339_n N_A_1238_47#_c_1801_n 0.0254125f $X=6.675 $Y=1.16
+ $X2=0 $Y2=0
cc_1048 N_A_726_47#_c_1334_n N_A_1238_47#_c_1802_n 0.0093209f $X=9.6 $Y=1.295
+ $X2=0 $Y2=0
cc_1049 N_A_726_47#_M1000_g N_VPWR_c_1926_n 0.00304014f $X=6.615 $Y=2.285 $X2=0
+ $Y2=0
cc_1050 N_A_726_47#_M1007_s N_VPWR_c_1921_n 0.00225465f $X=3.75 $Y=1.835 $X2=0
+ $Y2=0
cc_1051 N_A_726_47#_M1000_g N_VPWR_c_1921_n 9.49986e-19 $X=6.615 $Y=2.285 $X2=0
+ $Y2=0
cc_1052 N_A_726_47#_c_1349_n N_A_658_367#_c_2195_n 0.0629392f $X=3.83 $Y=1.96
+ $X2=0 $Y2=0
cc_1053 N_A_726_47#_M1007_s N_A_658_367#_c_2208_n 0.00340092f $X=3.75 $Y=1.835
+ $X2=0 $Y2=0
cc_1054 N_A_726_47#_c_1434_n N_A_658_367#_c_2208_n 0.0163574f $X=3.89 $Y=1.98
+ $X2=0 $Y2=0
cc_1055 N_A_726_47#_c_1349_n N_A_658_367#_c_2196_n 0.019167f $X=3.83 $Y=1.96
+ $X2=0 $Y2=0
cc_1056 N_A_726_47#_c_1329_n N_A_658_367#_c_2196_n 0.00423005f $X=5.435 $Y=1.08
+ $X2=0 $Y2=0
cc_1057 N_A_726_47#_c_1346_n N_A_658_367#_c_2197_n 0.00336301f $X=5.535 $Y=1.08
+ $X2=0 $Y2=0
cc_1058 N_A_726_47#_c_1340_n N_Z_c_2262_n 0.00154233f $X=10.305 $Y=1.2 $X2=0
+ $Y2=0
cc_1059 N_A_726_47#_c_1341_n N_Z_c_2262_n 0.00349691f $X=9.745 $Y=1.2 $X2=0
+ $Y2=0
cc_1060 N_A_726_47#_M1005_g N_Z_c_2250_n 0.0126545f $X=10.38 $Y=0.555 $X2=0
+ $Y2=0
cc_1061 N_A_726_47#_M1006_g N_Z_c_2250_n 6.57936e-19 $X=10.81 $Y=0.555 $X2=0
+ $Y2=0
cc_1062 N_A_726_47#_c_1310_n N_Z_c_2250_n 0.00440309f $X=13.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1063 N_A_726_47#_c_1337_n N_Z_c_2250_n 0.0353753f $X=13.185 $Y=1.295 $X2=0
+ $Y2=0
cc_1064 N_A_726_47#_c_1340_n N_Z_c_2250_n 0.0230572f $X=10.305 $Y=1.2 $X2=0
+ $Y2=0
cc_1065 N_A_726_47#_c_1341_n N_Z_c_2250_n 0.0256972f $X=9.745 $Y=1.2 $X2=0 $Y2=0
cc_1066 N_A_726_47#_c_1342_n N_Z_c_2250_n 0.0256972f $X=10.605 $Y=1.2 $X2=0
+ $Y2=0
cc_1067 N_A_726_47#_M1005_g N_Z_c_2251_n 6.57936e-19 $X=10.38 $Y=0.555 $X2=0
+ $Y2=0
cc_1068 N_A_726_47#_M1006_g N_Z_c_2251_n 0.0113519f $X=10.81 $Y=0.555 $X2=0
+ $Y2=0
cc_1069 N_A_726_47#_M1013_g N_Z_c_2251_n 0.0113519f $X=11.24 $Y=0.555 $X2=0
+ $Y2=0
cc_1070 N_A_726_47#_M1021_g N_Z_c_2251_n 6.57936e-19 $X=11.67 $Y=0.555 $X2=0
+ $Y2=0
cc_1071 N_A_726_47#_c_1310_n N_Z_c_2251_n 0.022527f $X=13.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1072 N_A_726_47#_c_1337_n N_Z_c_2251_n 0.0353753f $X=13.185 $Y=1.295 $X2=0
+ $Y2=0
cc_1073 N_A_726_47#_c_1342_n N_Z_c_2251_n 0.0256972f $X=10.605 $Y=1.2 $X2=0
+ $Y2=0
cc_1074 N_A_726_47#_c_1343_n N_Z_c_2251_n 0.0256972f $X=11.445 $Y=1.2 $X2=0
+ $Y2=0
cc_1075 N_A_726_47#_M1013_g N_Z_c_2252_n 6.57936e-19 $X=11.24 $Y=0.555 $X2=0
+ $Y2=0
cc_1076 N_A_726_47#_M1021_g N_Z_c_2252_n 0.0113519f $X=11.67 $Y=0.555 $X2=0
+ $Y2=0
cc_1077 N_A_726_47#_c_1305_n N_Z_c_2252_n 0.00987762f $X=12.1 $Y=0.985 $X2=0
+ $Y2=0
cc_1078 N_A_726_47#_c_1306_n N_Z_c_2252_n 5.10745e-19 $X=12.53 $Y=0.985 $X2=0
+ $Y2=0
cc_1079 N_A_726_47#_c_1310_n N_Z_c_2252_n 0.024478f $X=13.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1080 N_A_726_47#_c_1337_n N_Z_c_2252_n 0.0353753f $X=13.185 $Y=1.295 $X2=0
+ $Y2=0
cc_1081 N_A_726_47#_c_1343_n N_Z_c_2252_n 0.0256972f $X=11.445 $Y=1.2 $X2=0
+ $Y2=0
cc_1082 N_A_726_47#_c_1344_n N_Z_c_2252_n 0.0256972f $X=12.325 $Y=1.2 $X2=0
+ $Y2=0
cc_1083 N_A_726_47#_c_1305_n N_Z_c_2253_n 5.10745e-19 $X=12.1 $Y=0.985 $X2=0
+ $Y2=0
cc_1084 N_A_726_47#_c_1306_n N_Z_c_2253_n 0.00987762f $X=12.53 $Y=0.985 $X2=0
+ $Y2=0
cc_1085 N_A_726_47#_c_1307_n N_Z_c_2253_n 0.00987762f $X=12.96 $Y=0.985 $X2=0
+ $Y2=0
cc_1086 N_A_726_47#_c_1308_n N_Z_c_2253_n 5.10745e-19 $X=13.39 $Y=0.985 $X2=0
+ $Y2=0
cc_1087 N_A_726_47#_c_1310_n N_Z_c_2253_n 0.0265644f $X=13.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1088 N_A_726_47#_c_1337_n N_Z_c_2253_n 0.0353753f $X=13.185 $Y=1.295 $X2=0
+ $Y2=0
cc_1089 N_A_726_47#_c_1344_n N_Z_c_2253_n 0.0256972f $X=12.325 $Y=1.2 $X2=0
+ $Y2=0
cc_1090 N_A_726_47#_c_1345_n N_Z_c_2253_n 0.0256972f $X=13.185 $Y=1.2 $X2=0
+ $Y2=0
cc_1091 N_A_726_47#_c_1307_n N_Z_c_2254_n 5.10745e-19 $X=12.96 $Y=0.985 $X2=0
+ $Y2=0
cc_1092 N_A_726_47#_c_1308_n N_Z_c_2254_n 0.00987762f $X=13.39 $Y=0.985 $X2=0
+ $Y2=0
cc_1093 N_A_726_47#_c_1309_n N_Z_c_2254_n 0.0109356f $X=13.745 $Y=1.06 $X2=0
+ $Y2=0
cc_1094 N_A_726_47#_c_1310_n N_Z_c_2254_n 0.00980356f $X=13.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1095 N_A_726_47#_c_1311_n N_Z_c_2254_n 0.00987762f $X=13.82 $Y=0.985 $X2=0
+ $Y2=0
cc_1096 N_A_726_47#_c_1313_n N_Z_c_2254_n 5.10745e-19 $X=14.25 $Y=0.985 $X2=0
+ $Y2=0
cc_1097 N_A_726_47#_c_1324_n N_Z_c_2254_n 0.00446221f $X=13.82 $Y=1.06 $X2=0
+ $Y2=0
cc_1098 N_A_726_47#_c_1337_n N_Z_c_2254_n 0.00752419f $X=13.185 $Y=1.295 $X2=0
+ $Y2=0
cc_1099 N_A_726_47#_c_1345_n N_Z_c_2254_n 0.0257931f $X=13.185 $Y=1.2 $X2=0
+ $Y2=0
cc_1100 N_A_726_47#_c_1311_n N_Z_c_2255_n 5.10745e-19 $X=13.82 $Y=0.985 $X2=0
+ $Y2=0
cc_1101 N_A_726_47#_c_1313_n N_Z_c_2255_n 0.00987762f $X=14.25 $Y=0.985 $X2=0
+ $Y2=0
cc_1102 N_A_726_47#_c_1314_n N_Z_c_2255_n 0.0088652f $X=14.605 $Y=1.06 $X2=0
+ $Y2=0
cc_1103 N_A_726_47#_c_1315_n N_Z_c_2255_n 0.00987762f $X=14.68 $Y=0.985 $X2=0
+ $Y2=0
cc_1104 N_A_726_47#_c_1317_n N_Z_c_2255_n 5.10745e-19 $X=15.11 $Y=0.985 $X2=0
+ $Y2=0
cc_1105 N_A_726_47#_c_1325_n N_Z_c_2255_n 0.00428178f $X=14.25 $Y=1.06 $X2=0
+ $Y2=0
cc_1106 N_A_726_47#_c_1326_n N_Z_c_2255_n 0.00428178f $X=14.68 $Y=1.06 $X2=0
+ $Y2=0
cc_1107 N_A_726_47#_c_1315_n N_Z_c_2256_n 5.09252e-19 $X=14.68 $Y=0.985 $X2=0
+ $Y2=0
cc_1108 N_A_726_47#_c_1317_n N_Z_c_2256_n 0.00983119f $X=15.11 $Y=0.985 $X2=0
+ $Y2=0
cc_1109 N_A_726_47#_c_1318_n N_Z_c_2256_n 0.0088652f $X=15.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1110 N_A_726_47#_c_1319_n N_Z_c_2256_n 0.00983119f $X=15.54 $Y=0.985 $X2=0
+ $Y2=0
cc_1111 N_A_726_47#_c_1321_n N_Z_c_2256_n 5.09252e-19 $X=15.97 $Y=0.985 $X2=0
+ $Y2=0
cc_1112 N_A_726_47#_c_1327_n N_Z_c_2256_n 0.00428178f $X=15.11 $Y=1.06 $X2=0
+ $Y2=0
cc_1113 N_A_726_47#_c_1328_n N_Z_c_2256_n 0.00428178f $X=15.54 $Y=1.06 $X2=0
+ $Y2=0
cc_1114 N_A_726_47#_c_1319_n N_Z_c_2257_n 5.10745e-19 $X=15.54 $Y=0.985 $X2=0
+ $Y2=0
cc_1115 N_A_726_47#_c_1320_n N_Z_c_2257_n 0.00731f $X=15.895 $Y=1.06 $X2=0 $Y2=0
cc_1116 N_A_726_47#_c_1321_n N_Z_c_2257_n 0.010768f $X=15.97 $Y=0.985 $X2=0
+ $Y2=0
cc_1117 N_A_726_47#_c_1329_n N_VGND_M1049_s 0.00680998f $X=5.435 $Y=1.08 $X2=0
+ $Y2=0
cc_1118 N_A_726_47#_c_1346_n N_VGND_M1010_s 0.0019144f $X=5.535 $Y=1.08 $X2=0
+ $Y2=0
cc_1119 N_A_726_47#_M1011_g N_VGND_c_2519_n 0.00830301f $X=6.615 $Y=0.445 $X2=0
+ $Y2=0
cc_1120 N_A_726_47#_M1005_g N_VGND_c_2521_n 0.00271808f $X=10.38 $Y=0.555 $X2=0
+ $Y2=0
cc_1121 N_A_726_47#_M1006_g N_VGND_c_2521_n 0.00271808f $X=10.81 $Y=0.555 $X2=0
+ $Y2=0
cc_1122 N_A_726_47#_c_1310_n N_VGND_c_2521_n 7.91474e-19 $X=13.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1123 N_A_726_47#_c_1337_n N_VGND_c_2521_n 0.00100776f $X=13.185 $Y=1.295
+ $X2=0 $Y2=0
cc_1124 N_A_726_47#_c_1342_n N_VGND_c_2521_n 0.0130159f $X=10.605 $Y=1.2 $X2=0
+ $Y2=0
cc_1125 N_A_726_47#_M1013_g N_VGND_c_2522_n 0.00271808f $X=11.24 $Y=0.555 $X2=0
+ $Y2=0
cc_1126 N_A_726_47#_M1021_g N_VGND_c_2522_n 0.00271808f $X=11.67 $Y=0.555 $X2=0
+ $Y2=0
cc_1127 N_A_726_47#_c_1310_n N_VGND_c_2522_n 7.91474e-19 $X=13.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1128 N_A_726_47#_c_1337_n N_VGND_c_2522_n 0.00100776f $X=13.185 $Y=1.295
+ $X2=0 $Y2=0
cc_1129 N_A_726_47#_c_1343_n N_VGND_c_2522_n 0.0130159f $X=11.445 $Y=1.2 $X2=0
+ $Y2=0
cc_1130 N_A_726_47#_M1021_g N_VGND_c_2523_n 0.0054895f $X=11.67 $Y=0.555 $X2=0
+ $Y2=0
cc_1131 N_A_726_47#_c_1305_n N_VGND_c_2523_n 0.0054895f $X=12.1 $Y=0.985 $X2=0
+ $Y2=0
cc_1132 N_A_726_47#_c_1305_n N_VGND_c_2524_n 0.00271808f $X=12.1 $Y=0.985 $X2=0
+ $Y2=0
cc_1133 N_A_726_47#_c_1306_n N_VGND_c_2524_n 0.00271808f $X=12.53 $Y=0.985 $X2=0
+ $Y2=0
cc_1134 N_A_726_47#_c_1310_n N_VGND_c_2524_n 0.00254294f $X=13.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1135 N_A_726_47#_c_1337_n N_VGND_c_2524_n 0.00100776f $X=13.185 $Y=1.295
+ $X2=0 $Y2=0
cc_1136 N_A_726_47#_c_1344_n N_VGND_c_2524_n 0.0130158f $X=12.325 $Y=1.2 $X2=0
+ $Y2=0
cc_1137 N_A_726_47#_c_1307_n N_VGND_c_2525_n 0.00271808f $X=12.96 $Y=0.985 $X2=0
+ $Y2=0
cc_1138 N_A_726_47#_c_1308_n N_VGND_c_2525_n 0.00271808f $X=13.39 $Y=0.985 $X2=0
+ $Y2=0
cc_1139 N_A_726_47#_c_1310_n N_VGND_c_2525_n 0.00254294f $X=13.465 $Y=1.06 $X2=0
+ $Y2=0
cc_1140 N_A_726_47#_c_1337_n N_VGND_c_2525_n 0.00100776f $X=13.185 $Y=1.295
+ $X2=0 $Y2=0
cc_1141 N_A_726_47#_c_1345_n N_VGND_c_2525_n 0.0130158f $X=13.185 $Y=1.2 $X2=0
+ $Y2=0
cc_1142 N_A_726_47#_c_1311_n N_VGND_c_2526_n 0.00271808f $X=13.82 $Y=0.985 $X2=0
+ $Y2=0
cc_1143 N_A_726_47#_c_1312_n N_VGND_c_2526_n 0.0026233f $X=14.175 $Y=1.06 $X2=0
+ $Y2=0
cc_1144 N_A_726_47#_c_1313_n N_VGND_c_2526_n 0.00271808f $X=14.25 $Y=0.985 $X2=0
+ $Y2=0
cc_1145 N_A_726_47#_c_1315_n N_VGND_c_2527_n 0.00271808f $X=14.68 $Y=0.985 $X2=0
+ $Y2=0
cc_1146 N_A_726_47#_c_1316_n N_VGND_c_2527_n 0.0026233f $X=15.035 $Y=1.06 $X2=0
+ $Y2=0
cc_1147 N_A_726_47#_c_1317_n N_VGND_c_2527_n 0.00271808f $X=15.11 $Y=0.985 $X2=0
+ $Y2=0
cc_1148 N_A_726_47#_c_1319_n N_VGND_c_2528_n 0.00271808f $X=15.54 $Y=0.985 $X2=0
+ $Y2=0
cc_1149 N_A_726_47#_c_1320_n N_VGND_c_2528_n 0.0026233f $X=15.895 $Y=1.06 $X2=0
+ $Y2=0
cc_1150 N_A_726_47#_c_1321_n N_VGND_c_2528_n 0.00271808f $X=15.97 $Y=0.985 $X2=0
+ $Y2=0
cc_1151 N_A_726_47#_M1011_g N_VGND_c_2531_n 0.0038319f $X=6.615 $Y=0.445 $X2=0
+ $Y2=0
cc_1152 N_A_726_47#_M1005_g N_VGND_c_2533_n 0.0054895f $X=10.38 $Y=0.555 $X2=0
+ $Y2=0
cc_1153 N_A_726_47#_M1006_g N_VGND_c_2535_n 0.0054895f $X=10.81 $Y=0.555 $X2=0
+ $Y2=0
cc_1154 N_A_726_47#_M1013_g N_VGND_c_2535_n 0.0054895f $X=11.24 $Y=0.555 $X2=0
+ $Y2=0
cc_1155 N_A_726_47#_c_1306_n N_VGND_c_2537_n 0.0054895f $X=12.53 $Y=0.985 $X2=0
+ $Y2=0
cc_1156 N_A_726_47#_c_1307_n N_VGND_c_2537_n 0.0054895f $X=12.96 $Y=0.985 $X2=0
+ $Y2=0
cc_1157 N_A_726_47#_c_1308_n N_VGND_c_2539_n 0.0054895f $X=13.39 $Y=0.985 $X2=0
+ $Y2=0
cc_1158 N_A_726_47#_c_1311_n N_VGND_c_2539_n 0.0054895f $X=13.82 $Y=0.985 $X2=0
+ $Y2=0
cc_1159 N_A_726_47#_c_1313_n N_VGND_c_2541_n 0.0054895f $X=14.25 $Y=0.985 $X2=0
+ $Y2=0
cc_1160 N_A_726_47#_c_1315_n N_VGND_c_2541_n 0.0054895f $X=14.68 $Y=0.985 $X2=0
+ $Y2=0
cc_1161 N_A_726_47#_c_1317_n N_VGND_c_2543_n 0.00549117f $X=15.11 $Y=0.985 $X2=0
+ $Y2=0
cc_1162 N_A_726_47#_c_1319_n N_VGND_c_2543_n 0.00549117f $X=15.54 $Y=0.985 $X2=0
+ $Y2=0
cc_1163 N_A_726_47#_c_1321_n N_VGND_c_2549_n 0.0054895f $X=15.97 $Y=0.985 $X2=0
+ $Y2=0
cc_1164 N_A_726_47#_M1024_d N_VGND_c_2550_n 0.00225465f $X=3.63 $Y=0.235 $X2=0
+ $Y2=0
cc_1165 N_A_726_47#_M1001_d N_VGND_c_2550_n 0.00569151f $X=4.84 $Y=0.235 $X2=0
+ $Y2=0
cc_1166 N_A_726_47#_M1011_g N_VGND_c_2550_n 0.00470043f $X=6.615 $Y=0.445 $X2=0
+ $Y2=0
cc_1167 N_A_726_47#_M1005_g N_VGND_c_2550_n 0.0110927f $X=10.38 $Y=0.555 $X2=0
+ $Y2=0
cc_1168 N_A_726_47#_M1006_g N_VGND_c_2550_n 0.00979301f $X=10.81 $Y=0.555 $X2=0
+ $Y2=0
cc_1169 N_A_726_47#_M1013_g N_VGND_c_2550_n 0.00979301f $X=11.24 $Y=0.555 $X2=0
+ $Y2=0
cc_1170 N_A_726_47#_M1021_g N_VGND_c_2550_n 0.00979301f $X=11.67 $Y=0.555 $X2=0
+ $Y2=0
cc_1171 N_A_726_47#_c_1305_n N_VGND_c_2550_n 0.00979301f $X=12.1 $Y=0.985 $X2=0
+ $Y2=0
cc_1172 N_A_726_47#_c_1306_n N_VGND_c_2550_n 0.00979301f $X=12.53 $Y=0.985 $X2=0
+ $Y2=0
cc_1173 N_A_726_47#_c_1307_n N_VGND_c_2550_n 0.00979301f $X=12.96 $Y=0.985 $X2=0
+ $Y2=0
cc_1174 N_A_726_47#_c_1308_n N_VGND_c_2550_n 0.00979301f $X=13.39 $Y=0.985 $X2=0
+ $Y2=0
cc_1175 N_A_726_47#_c_1311_n N_VGND_c_2550_n 0.00979301f $X=13.82 $Y=0.985 $X2=0
+ $Y2=0
cc_1176 N_A_726_47#_c_1313_n N_VGND_c_2550_n 0.00979301f $X=14.25 $Y=0.985 $X2=0
+ $Y2=0
cc_1177 N_A_726_47#_c_1315_n N_VGND_c_2550_n 0.00979301f $X=14.68 $Y=0.985 $X2=0
+ $Y2=0
cc_1178 N_A_726_47#_c_1317_n N_VGND_c_2550_n 0.00979311f $X=15.11 $Y=0.985 $X2=0
+ $Y2=0
cc_1179 N_A_726_47#_c_1319_n N_VGND_c_2550_n 0.00979311f $X=15.54 $Y=0.985 $X2=0
+ $Y2=0
cc_1180 N_A_726_47#_c_1321_n N_VGND_c_2550_n 0.0110927f $X=15.97 $Y=0.985 $X2=0
+ $Y2=0
cc_1181 N_A_726_47#_M1011_g N_A_1451_47#_c_2767_n 0.00323073f $X=6.615 $Y=0.445
+ $X2=0 $Y2=0
cc_1182 N_A_726_47#_c_1334_n N_A_1451_47#_c_2757_n 0.0235872f $X=9.6 $Y=1.295
+ $X2=0 $Y2=0
cc_1183 N_A_726_47#_c_1334_n N_A_1451_47#_c_2758_n 0.00553971f $X=9.6 $Y=1.295
+ $X2=0 $Y2=0
cc_1184 N_A_726_47#_c_1334_n N_A_1451_47#_c_2760_n 0.00821049f $X=9.6 $Y=1.295
+ $X2=0 $Y2=0
cc_1185 N_A_726_47#_c_1340_n N_A_1451_47#_c_2760_n 6.57308e-19 $X=10.305 $Y=1.2
+ $X2=0 $Y2=0
cc_1186 N_A_726_47#_c_1341_n N_A_1451_47#_c_2760_n 0.0044621f $X=9.745 $Y=1.2
+ $X2=0 $Y2=0
cc_1187 N_A_M1010_g N_A_1238_47#_c_1807_n 7.99369e-19 $X=5.395 $Y=0.655 $X2=0
+ $Y2=0
cc_1188 N_A_M1002_g N_A_1238_47#_c_1797_n 8.94931e-19 $X=7.615 $Y=0.655 $X2=0
+ $Y2=0
cc_1189 N_A_M1002_g N_A_1238_47#_c_1799_n 0.00432636f $X=7.615 $Y=0.655 $X2=0
+ $Y2=0
cc_1190 N_A_c_1653_n N_A_1238_47#_c_1804_n 0.00422474f $X=7.125 $Y=3.075 $X2=0
+ $Y2=0
cc_1191 N_A_c_1639_n N_A_1238_47#_c_1804_n 0.00487705f $X=7.2 $Y=1.65 $X2=0
+ $Y2=0
cc_1192 N_A_c_1656_n N_A_1238_47#_c_1804_n 5.96015e-19 $X=7.645 $Y=1.725 $X2=0
+ $Y2=0
cc_1193 N_A_c_1638_n N_A_1238_47#_c_1800_n 0.0131505f $X=7.54 $Y=1.65 $X2=0
+ $Y2=0
cc_1194 N_A_c_1639_n N_A_1238_47#_c_1800_n 4.21068e-19 $X=7.2 $Y=1.65 $X2=0
+ $Y2=0
cc_1195 N_A_M1002_g N_A_1238_47#_c_1800_n 0.0147606f $X=7.615 $Y=0.655 $X2=0
+ $Y2=0
cc_1196 N_A_c_1641_n N_A_1238_47#_c_1800_n 0.00433481f $X=7.97 $Y=1.65 $X2=0
+ $Y2=0
cc_1197 N_A_M1003_g N_A_1238_47#_c_1800_n 0.0120019f $X=8.045 $Y=0.655 $X2=0
+ $Y2=0
cc_1198 N_A_c_1643_n N_A_1238_47#_c_1800_n 0.00440164f $X=7.63 $Y=1.65 $X2=0
+ $Y2=0
cc_1199 N_A_c_1644_n N_A_1238_47#_c_1800_n 0.00279845f $X=8.06 $Y=1.65 $X2=0
+ $Y2=0
cc_1200 N_A_c_1651_n N_A_1238_47#_c_1805_n 0.00542511f $X=7.05 $Y=3.15 $X2=0
+ $Y2=0
cc_1201 N_A_c_1653_n N_A_1238_47#_c_1805_n 0.010255f $X=7.125 $Y=3.075 $X2=0
+ $Y2=0
cc_1202 N_A_c_1653_n N_A_1238_47#_c_1806_n 0.0131697f $X=7.125 $Y=3.075 $X2=0
+ $Y2=0
cc_1203 N_A_c_1656_n N_A_1238_47#_c_1806_n 6.21675e-19 $X=7.645 $Y=1.725 $X2=0
+ $Y2=0
cc_1204 N_A_c_1639_n N_A_1238_47#_c_1801_n 0.00397919f $X=7.2 $Y=1.65 $X2=0
+ $Y2=0
cc_1205 N_A_M1003_g N_A_1238_47#_c_1802_n 0.0221307f $X=8.045 $Y=0.655 $X2=0
+ $Y2=0
cc_1206 N_A_c_1644_n N_A_1238_47#_c_1802_n 0.00196276f $X=8.06 $Y=1.65 $X2=0
+ $Y2=0
cc_1207 N_A_M1003_g N_A_1238_47#_c_1803_n 0.0219475f $X=8.045 $Y=0.655 $X2=0
+ $Y2=0
cc_1208 N_A_M1030_g N_VPWR_c_1925_n 0.0100794f $X=4.615 $Y=2.465 $X2=0 $Y2=0
cc_1209 N_A_c_1647_n N_VPWR_c_1925_n 0.0116849f $X=5.045 $Y=1.715 $X2=0 $Y2=0
cc_1210 N_A_c_1650_n N_VPWR_c_1925_n 0.00102654f $X=5.715 $Y=3.075 $X2=0 $Y2=0
cc_1211 N_A_c_1650_n N_VPWR_c_1926_n 0.0159523f $X=5.715 $Y=3.075 $X2=0 $Y2=0
cc_1212 N_A_c_1651_n N_VPWR_c_1926_n 0.0244686f $X=7.05 $Y=3.15 $X2=0 $Y2=0
cc_1213 N_A_c_1653_n N_VPWR_c_1927_n 0.0179948f $X=7.125 $Y=3.075 $X2=0 $Y2=0
cc_1214 N_A_c_1638_n N_VPWR_c_1927_n 0.00255175f $X=7.54 $Y=1.65 $X2=0 $Y2=0
cc_1215 N_A_c_1656_n N_VPWR_c_1927_n 0.00408079f $X=7.645 $Y=1.725 $X2=0 $Y2=0
cc_1216 N_A_c_1658_n N_VPWR_c_1928_n 0.0231672f $X=8.075 $Y=1.725 $X2=0 $Y2=0
cc_1217 N_A_M1030_g N_VPWR_c_1942_n 0.00486043f $X=4.615 $Y=2.465 $X2=0 $Y2=0
cc_1218 N_A_c_1651_n N_VPWR_c_1944_n 0.03343f $X=7.05 $Y=3.15 $X2=0 $Y2=0
cc_1219 N_A_c_1647_n N_VPWR_c_1963_n 0.00486043f $X=5.045 $Y=1.715 $X2=0 $Y2=0
cc_1220 N_A_c_1652_n N_VPWR_c_1963_n 0.00796123f $X=5.79 $Y=3.15 $X2=0 $Y2=0
cc_1221 N_A_c_1656_n N_VPWR_c_1964_n 0.00549284f $X=7.645 $Y=1.725 $X2=0 $Y2=0
cc_1222 N_A_c_1658_n N_VPWR_c_1964_n 0.00549284f $X=8.075 $Y=1.725 $X2=0 $Y2=0
cc_1223 N_A_M1030_g N_VPWR_c_1921_n 0.00482043f $X=4.615 $Y=2.465 $X2=0 $Y2=0
cc_1224 N_A_c_1647_n N_VPWR_c_1921_n 0.0051394f $X=5.045 $Y=1.715 $X2=0 $Y2=0
cc_1225 N_A_c_1651_n N_VPWR_c_1921_n 0.0466702f $X=7.05 $Y=3.15 $X2=0 $Y2=0
cc_1226 N_A_c_1652_n N_VPWR_c_1921_n 0.0105448f $X=5.79 $Y=3.15 $X2=0 $Y2=0
cc_1227 N_A_c_1656_n N_VPWR_c_1921_n 0.0100092f $X=7.645 $Y=1.725 $X2=0 $Y2=0
cc_1228 N_A_c_1658_n N_VPWR_c_1921_n 0.0113003f $X=8.075 $Y=1.725 $X2=0 $Y2=0
cc_1229 N_A_M1030_g N_A_658_367#_c_2196_n 0.00283516f $X=4.615 $Y=2.465 $X2=0
+ $Y2=0
cc_1230 A N_A_658_367#_c_2196_n 7.93802e-19 $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_1231 N_A_M1030_g N_A_658_367#_c_2201_n 0.0137188f $X=4.615 $Y=2.465 $X2=0
+ $Y2=0
cc_1232 N_A_c_1647_n N_A_658_367#_c_2201_n 0.0126676f $X=5.045 $Y=1.715 $X2=0
+ $Y2=0
cc_1233 N_A_c_1637_n N_A_658_367#_c_2201_n 0.00193941f $X=5.47 $Y=1.64 $X2=0
+ $Y2=0
cc_1234 A N_A_658_367#_c_2201_n 0.0106298f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_1235 N_A_c_1645_n N_A_658_367#_c_2201_n 9.91138e-19 $X=5.135 $Y=1.51 $X2=0
+ $Y2=0
cc_1236 N_A_c_1647_n N_A_658_367#_c_2197_n 0.00526545f $X=5.045 $Y=1.715 $X2=0
+ $Y2=0
cc_1237 N_A_c_1637_n N_A_658_367#_c_2197_n 0.00679431f $X=5.47 $Y=1.64 $X2=0
+ $Y2=0
cc_1238 N_A_c_1650_n N_A_658_367#_c_2197_n 0.00546871f $X=5.715 $Y=3.075 $X2=0
+ $Y2=0
cc_1239 N_A_c_1647_n N_A_658_367#_c_2198_n 0.00775858f $X=5.045 $Y=1.715 $X2=0
+ $Y2=0
cc_1240 N_A_c_1650_n N_A_658_367#_c_2198_n 0.00867389f $X=5.715 $Y=3.075 $X2=0
+ $Y2=0
cc_1241 N_A_M1001_g N_VGND_c_2517_n 0.0105661f $X=4.765 $Y=0.655 $X2=0 $Y2=0
cc_1242 N_A_M1010_g N_VGND_c_2517_n 0.00179115f $X=5.395 $Y=0.655 $X2=0 $Y2=0
cc_1243 N_A_M1010_g N_VGND_c_2518_n 0.00985574f $X=5.395 $Y=0.655 $X2=0 $Y2=0
cc_1244 N_A_M1002_g N_VGND_c_2519_n 0.00271318f $X=7.615 $Y=0.655 $X2=0 $Y2=0
cc_1245 N_A_M1002_g N_VGND_c_2520_n 0.00332744f $X=7.615 $Y=0.655 $X2=0 $Y2=0
cc_1246 N_A_M1003_g N_VGND_c_2520_n 0.0114807f $X=8.045 $Y=0.655 $X2=0 $Y2=0
cc_1247 N_A_M1001_g N_VGND_c_2529_n 0.00354752f $X=4.765 $Y=0.655 $X2=0 $Y2=0
cc_1248 N_A_M1010_g N_VGND_c_2529_n 0.00426565f $X=5.395 $Y=0.655 $X2=0 $Y2=0
cc_1249 N_A_M1003_g N_VGND_c_2533_n 0.00486043f $X=8.045 $Y=0.655 $X2=0 $Y2=0
cc_1250 N_A_M1002_g N_VGND_c_2548_n 0.00548839f $X=7.615 $Y=0.655 $X2=0 $Y2=0
cc_1251 N_A_M1001_g N_VGND_c_2550_n 0.00467942f $X=4.765 $Y=0.655 $X2=0 $Y2=0
cc_1252 N_A_M1010_g N_VGND_c_2550_n 0.00706722f $X=5.395 $Y=0.655 $X2=0 $Y2=0
cc_1253 N_A_M1002_g N_VGND_c_2550_n 0.0111559f $X=7.615 $Y=0.655 $X2=0 $Y2=0
cc_1254 N_A_M1003_g N_VGND_c_2550_n 0.0085771f $X=8.045 $Y=0.655 $X2=0 $Y2=0
cc_1255 N_A_M1002_g N_A_1451_47#_c_2767_n 0.0126834f $X=7.615 $Y=0.655 $X2=0
+ $Y2=0
cc_1256 N_A_M1003_g N_A_1451_47#_c_2767_n 6.64616e-19 $X=8.045 $Y=0.655 $X2=0
+ $Y2=0
cc_1257 N_A_M1002_g N_A_1451_47#_c_2757_n 0.0111208f $X=7.615 $Y=0.655 $X2=0
+ $Y2=0
cc_1258 N_A_c_1641_n N_A_1451_47#_c_2757_n 3.68268e-19 $X=7.97 $Y=1.65 $X2=0
+ $Y2=0
cc_1259 N_A_M1003_g N_A_1451_47#_c_2757_n 0.014649f $X=8.045 $Y=0.655 $X2=0
+ $Y2=0
cc_1260 N_A_c_1638_n N_A_1451_47#_c_2758_n 7.42231e-19 $X=7.54 $Y=1.65 $X2=0
+ $Y2=0
cc_1261 N_A_M1002_g N_A_1451_47#_c_2758_n 0.00345644f $X=7.615 $Y=0.655 $X2=0
+ $Y2=0
cc_1262 N_A_M1002_g N_A_1451_47#_c_2759_n 0.00206603f $X=7.615 $Y=0.655 $X2=0
+ $Y2=0
cc_1263 N_A_1238_47#_c_1805_n N_VPWR_c_1926_n 0.0224933f $X=6.83 $Y=2.01 $X2=0
+ $Y2=0
cc_1264 N_A_1238_47#_c_1806_n N_VPWR_c_1926_n 0.00552965f $X=7.105 $Y=1.93 $X2=0
+ $Y2=0
cc_1265 N_A_1238_47#_c_1800_n N_VPWR_c_1927_n 0.00375117f $X=8.525 $Y=1.44 $X2=0
+ $Y2=0
cc_1266 N_A_1238_47#_c_1805_n N_VPWR_c_1927_n 0.0318631f $X=6.83 $Y=2.01 $X2=0
+ $Y2=0
cc_1267 N_A_1238_47#_c_1805_n N_VPWR_c_1944_n 0.00703457f $X=6.83 $Y=2.01 $X2=0
+ $Y2=0
cc_1268 N_A_1238_47#_c_1805_n N_VPWR_c_1921_n 0.00887189f $X=6.83 $Y=2.01 $X2=0
+ $Y2=0
cc_1269 N_A_1238_47#_c_1797_n N_VGND_M1011_d 0.0025501f $X=7.02 $Y=0.73 $X2=0
+ $Y2=0
cc_1270 N_A_1238_47#_c_1807_n N_VGND_c_2518_n 0.0103102f $X=6.33 $Y=0.47 $X2=0
+ $Y2=0
cc_1271 N_A_1238_47#_c_1797_n N_VGND_c_2519_n 0.0196474f $X=7.02 $Y=0.73 $X2=0
+ $Y2=0
cc_1272 N_A_1238_47#_c_1803_n N_VGND_c_2520_n 0.00115093f $X=8.525 $Y=1.185
+ $X2=0 $Y2=0
cc_1273 N_A_1238_47#_c_1807_n N_VGND_c_2531_n 0.0191432f $X=6.33 $Y=0.47 $X2=0
+ $Y2=0
cc_1274 N_A_1238_47#_c_1797_n N_VGND_c_2531_n 0.00257363f $X=7.02 $Y=0.73 $X2=0
+ $Y2=0
cc_1275 N_A_1238_47#_c_1796_n N_VGND_c_2533_n 0.00359964f $X=9.065 $Y=1.185
+ $X2=0 $Y2=0
cc_1276 N_A_1238_47#_c_1803_n N_VGND_c_2533_n 0.0035993f $X=8.525 $Y=1.185 $X2=0
+ $Y2=0
cc_1277 N_A_1238_47#_c_1797_n N_VGND_c_2548_n 0.00362266f $X=7.02 $Y=0.73 $X2=0
+ $Y2=0
cc_1278 N_A_1238_47#_M1018_d N_VGND_c_2550_n 0.00297732f $X=6.19 $Y=0.235 $X2=0
+ $Y2=0
cc_1279 N_A_1238_47#_c_1796_n N_VGND_c_2550_n 0.00686121f $X=9.065 $Y=1.185
+ $X2=0 $Y2=0
cc_1280 N_A_1238_47#_c_1807_n N_VGND_c_2550_n 0.0125086f $X=6.33 $Y=0.47 $X2=0
+ $Y2=0
cc_1281 N_A_1238_47#_c_1797_n N_VGND_c_2550_n 0.0115093f $X=7.02 $Y=0.73 $X2=0
+ $Y2=0
cc_1282 N_A_1238_47#_c_1803_n N_VGND_c_2550_n 0.00576767f $X=8.525 $Y=1.185
+ $X2=0 $Y2=0
cc_1283 N_A_1238_47#_c_1797_n N_A_1451_47#_c_2767_n 0.0143078f $X=7.02 $Y=0.73
+ $X2=0 $Y2=0
cc_1284 N_A_1238_47#_c_1799_n N_A_1451_47#_c_2767_n 0.00817472f $X=7.105
+ $Y=1.275 $X2=0 $Y2=0
cc_1285 N_A_1238_47#_c_1800_n N_A_1451_47#_c_2757_n 0.0583494f $X=8.525 $Y=1.44
+ $X2=0 $Y2=0
cc_1286 N_A_1238_47#_c_1802_n N_A_1451_47#_c_2757_n 0.0032543f $X=8.525 $Y=1.26
+ $X2=0 $Y2=0
cc_1287 N_A_1238_47#_c_1803_n N_A_1451_47#_c_2757_n 0.00241546f $X=8.525
+ $Y=1.185 $X2=0 $Y2=0
cc_1288 N_A_1238_47#_c_1799_n N_A_1451_47#_c_2758_n 0.0140921f $X=7.105 $Y=1.275
+ $X2=0 $Y2=0
cc_1289 N_A_1238_47#_c_1800_n N_A_1451_47#_c_2758_n 0.0139193f $X=8.525 $Y=1.44
+ $X2=0 $Y2=0
cc_1290 N_A_1238_47#_c_1803_n N_A_1451_47#_c_2788_n 6.00691e-19 $X=8.525
+ $Y=1.185 $X2=0 $Y2=0
cc_1291 N_A_1238_47#_c_1796_n N_A_1451_47#_c_2789_n 9.2152e-19 $X=9.065 $Y=1.185
+ $X2=0 $Y2=0
cc_1292 N_A_1238_47#_c_1803_n N_A_1451_47#_c_2789_n 0.00806939f $X=8.525
+ $Y=1.185 $X2=0 $Y2=0
cc_1293 N_A_1238_47#_c_1796_n N_A_1451_47#_c_2762_n 0.0112699f $X=9.065 $Y=1.185
+ $X2=0 $Y2=0
cc_1294 N_A_1238_47#_c_1803_n N_A_1451_47#_c_2762_n 0.0110205f $X=8.525 $Y=1.185
+ $X2=0 $Y2=0
cc_1295 N_A_1238_47#_c_1796_n N_A_1451_47#_c_2760_n 0.00735376f $X=9.065
+ $Y=1.185 $X2=0 $Y2=0
cc_1296 N_VPWR_c_1921_n N_A_658_367#_M1007_d 0.00409662f $X=17.52 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_1297 N_VPWR_c_1921_n N_A_658_367#_M1023_d 0.0032464f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1298 N_VPWR_c_1921_n N_A_658_367#_M1045_s 0.00502036f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1299 N_VPWR_c_1924_n N_A_658_367#_c_2236_n 0.00598248f $X=2.595 $Y=2.6 $X2=0
+ $Y2=0
cc_1300 N_VPWR_c_1942_n N_A_658_367#_c_2236_n 0.0111659f $X=4.665 $Y=3.33 $X2=0
+ $Y2=0
cc_1301 N_VPWR_c_1921_n N_A_658_367#_c_2236_n 0.00656694f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1302 N_VPWR_c_1924_n N_A_658_367#_c_2195_n 0.0146001f $X=2.595 $Y=2.6 $X2=0
+ $Y2=0
cc_1303 N_VPWR_c_1942_n N_A_658_367#_c_2208_n 0.0534661f $X=4.665 $Y=3.33 $X2=0
+ $Y2=0
cc_1304 N_VPWR_c_1921_n N_A_658_367#_c_2208_n 0.0355256f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1305 N_VPWR_M1030_d N_A_658_367#_c_2201_n 0.0051181f $X=4.69 $Y=1.835 $X2=0
+ $Y2=0
cc_1306 N_VPWR_c_1925_n N_A_658_367#_c_2201_n 0.0159912f $X=4.83 $Y=2.895 $X2=0
+ $Y2=0
cc_1307 N_VPWR_c_1921_n N_A_658_367#_c_2201_n 0.0174331f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1308 N_VPWR_c_1926_n N_A_658_367#_c_2197_n 0.028739f $X=6.01 $Y=2.01 $X2=0
+ $Y2=0
cc_1309 N_VPWR_c_1925_n N_A_658_367#_c_2198_n 0.0171841f $X=4.83 $Y=2.895 $X2=0
+ $Y2=0
cc_1310 N_VPWR_c_1926_n N_A_658_367#_c_2198_n 0.0453411f $X=6.01 $Y=2.01 $X2=0
+ $Y2=0
cc_1311 N_VPWR_c_1963_n N_A_658_367#_c_2198_n 0.0164099f $X=5.845 $Y=3.33 $X2=0
+ $Y2=0
cc_1312 N_VPWR_c_1921_n N_A_658_367#_c_2198_n 0.0095959f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1313 N_VPWR_c_1921_n N_Z_M1004_s 0.00606379f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1314 N_VPWR_c_1921_n N_Z_M1009_s 0.00223819f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1315 N_VPWR_c_1921_n N_Z_M1014_s 0.00223819f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1316 N_VPWR_c_1921_n N_Z_M1017_s 0.00223819f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1317 N_VPWR_c_1921_n N_Z_M1025_s 0.00223819f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1318 N_VPWR_c_1921_n N_Z_M1027_s 0.00223819f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1319 N_VPWR_c_1921_n N_Z_M1033_s 0.00223819f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1320 N_VPWR_c_1921_n N_Z_M1037_s 0.00223819f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1321 N_VPWR_c_1921_n N_Z_M1048_s 0.00223819f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1322 N_VPWR_c_1921_n N_Z_M1051_s 0.00223819f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1323 N_VPWR_c_1928_n N_Z_c_2448_n 0.0245939f $X=8.37 $Y=2.27 $X2=0 $Y2=0
cc_1324 N_VPWR_c_1946_n N_Z_c_2448_n 0.0110337f $X=9.57 $Y=3.33 $X2=0 $Y2=0
cc_1325 N_VPWR_c_1921_n N_Z_c_2448_n 0.00648955f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1326 N_VPWR_M1008_d N_Z_c_2262_n 0.00278715f $X=9.595 $Y=1.835 $X2=0 $Y2=0
cc_1327 N_VPWR_c_1929_n N_Z_c_2262_n 0.0135053f $X=9.735 $Y=2.475 $X2=0 $Y2=0
cc_1328 N_VPWR_c_1948_n N_Z_c_2276_n 0.0177952f $X=10.51 $Y=3.33 $X2=0 $Y2=0
cc_1329 N_VPWR_c_1921_n N_Z_c_2276_n 0.0123247f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1330 N_VPWR_c_1950_n N_Z_c_2251_n 0.0177952f $X=11.37 $Y=3.33 $X2=0 $Y2=0
cc_1331 N_VPWR_c_1921_n N_Z_c_2251_n 0.0123247f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1332 N_VPWR_c_1932_n N_Z_c_2252_n 0.0177952f $X=12.23 $Y=3.33 $X2=0 $Y2=0
cc_1333 N_VPWR_c_1921_n N_Z_c_2252_n 0.0123247f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1334 N_VPWR_c_1952_n N_Z_c_2253_n 0.0177952f $X=13.09 $Y=3.33 $X2=0 $Y2=0
cc_1335 N_VPWR_c_1921_n N_Z_c_2253_n 0.0123247f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1336 N_VPWR_c_1954_n N_Z_c_2254_n 0.0177952f $X=13.95 $Y=3.33 $X2=0 $Y2=0
cc_1337 N_VPWR_c_1921_n N_Z_c_2254_n 0.0123247f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1338 N_VPWR_c_1956_n N_Z_c_2255_n 0.0177952f $X=14.81 $Y=3.33 $X2=0 $Y2=0
cc_1339 N_VPWR_c_1921_n N_Z_c_2255_n 0.0123247f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1340 N_VPWR_c_1958_n N_Z_c_2256_n 0.0177952f $X=15.67 $Y=3.33 $X2=0 $Y2=0
cc_1341 N_VPWR_c_1921_n N_Z_c_2256_n 0.0123247f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1342 N_VPWR_c_1938_n N_Z_c_2257_n 0.0177952f $X=16.53 $Y=3.33 $X2=0 $Y2=0
cc_1343 N_VPWR_c_1921_n N_Z_c_2257_n 0.0123247f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1344 N_VPWR_c_1965_n N_Z_c_2337_n 0.0177952f $X=17.39 $Y=3.33 $X2=0 $Y2=0
cc_1345 N_VPWR_c_1921_n N_Z_c_2337_n 0.0123247f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1346 N_VPWR_M1008_d N_Z_c_2343_n 0.00580551f $X=9.595 $Y=1.835 $X2=0 $Y2=0
cc_1347 N_VPWR_M1012_d N_Z_c_2343_n 0.00755348f $X=10.455 $Y=1.835 $X2=0 $Y2=0
cc_1348 N_VPWR_M1016_d N_Z_c_2343_n 0.00755348f $X=11.315 $Y=1.835 $X2=0 $Y2=0
cc_1349 N_VPWR_M1022_d N_Z_c_2343_n 0.00755348f $X=12.175 $Y=1.835 $X2=0 $Y2=0
cc_1350 N_VPWR_M1026_d N_Z_c_2343_n 0.00755348f $X=13.035 $Y=1.835 $X2=0 $Y2=0
cc_1351 N_VPWR_M1032_d N_Z_c_2343_n 0.00737217f $X=13.895 $Y=1.835 $X2=0 $Y2=0
cc_1352 N_VPWR_M1036_d N_Z_c_2343_n 0.00737217f $X=14.755 $Y=1.835 $X2=0 $Y2=0
cc_1353 N_VPWR_M1042_d N_Z_c_2343_n 0.00737217f $X=15.615 $Y=1.835 $X2=0 $Y2=0
cc_1354 N_VPWR_M1050_d N_Z_c_2343_n 0.00720066f $X=16.475 $Y=1.835 $X2=0 $Y2=0
cc_1355 N_VPWR_c_1928_n N_Z_c_2343_n 4.32939e-19 $X=8.37 $Y=2.27 $X2=0 $Y2=0
cc_1356 N_VPWR_c_1929_n N_Z_c_2343_n 0.00706262f $X=9.735 $Y=2.475 $X2=0 $Y2=0
cc_1357 N_VPWR_c_1930_n N_Z_c_2343_n 0.00945368f $X=10.595 $Y=2.455 $X2=0 $Y2=0
cc_1358 N_VPWR_c_1931_n N_Z_c_2343_n 0.00945368f $X=11.455 $Y=2.455 $X2=0 $Y2=0
cc_1359 N_VPWR_c_1933_n N_Z_c_2343_n 0.00945368f $X=12.315 $Y=2.455 $X2=0 $Y2=0
cc_1360 N_VPWR_c_1934_n N_Z_c_2343_n 0.00945368f $X=13.175 $Y=2.455 $X2=0 $Y2=0
cc_1361 N_VPWR_c_1935_n N_Z_c_2343_n 0.00607361f $X=14.035 $Y=2.455 $X2=0 $Y2=0
cc_1362 N_VPWR_c_1936_n N_Z_c_2343_n 0.00607361f $X=14.895 $Y=2.455 $X2=0 $Y2=0
cc_1363 N_VPWR_c_1937_n N_Z_c_2343_n 0.00607361f $X=15.755 $Y=2.455 $X2=0 $Y2=0
cc_1364 N_VPWR_c_1939_n N_Z_c_2343_n 0.00607361f $X=16.615 $Y=2.455 $X2=0 $Y2=0
cc_1365 N_Z_c_2252_n N_VGND_c_2523_n 0.0189236f $X=11.885 $Y=0.36 $X2=0 $Y2=0
cc_1366 N_Z_c_2250_n N_VGND_c_2533_n 0.0210192f $X=10.165 $Y=0.36 $X2=0 $Y2=0
cc_1367 N_Z_c_2251_n N_VGND_c_2535_n 0.0189236f $X=11.025 $Y=0.36 $X2=0 $Y2=0
cc_1368 N_Z_c_2253_n N_VGND_c_2537_n 0.0189236f $X=12.745 $Y=0.36 $X2=0 $Y2=0
cc_1369 N_Z_c_2254_n N_VGND_c_2539_n 0.0189236f $X=13.605 $Y=0.36 $X2=0 $Y2=0
cc_1370 N_Z_c_2255_n N_VGND_c_2541_n 0.0189236f $X=14.465 $Y=0.36 $X2=0 $Y2=0
cc_1371 N_Z_c_2256_n N_VGND_c_2543_n 0.0183421f $X=15.325 $Y=0.36 $X2=0 $Y2=0
cc_1372 N_Z_c_2257_n N_VGND_c_2549_n 0.0210192f $X=16.185 $Y=0.36 $X2=0 $Y2=0
cc_1373 N_Z_M1005_s N_VGND_c_2550_n 0.00231914f $X=10.02 $Y=0.235 $X2=0 $Y2=0
cc_1374 N_Z_M1006_s N_VGND_c_2550_n 0.00223559f $X=10.885 $Y=0.235 $X2=0 $Y2=0
cc_1375 N_Z_M1021_s N_VGND_c_2550_n 0.00223559f $X=11.745 $Y=0.235 $X2=0 $Y2=0
cc_1376 N_Z_M1034_s N_VGND_c_2550_n 0.00223559f $X=12.605 $Y=0.235 $X2=0 $Y2=0
cc_1377 N_Z_M1043_s N_VGND_c_2550_n 0.00223559f $X=13.465 $Y=0.235 $X2=0 $Y2=0
cc_1378 N_Z_M1047_s N_VGND_c_2550_n 0.00223559f $X=14.325 $Y=0.235 $X2=0 $Y2=0
cc_1379 N_Z_M1056_s N_VGND_c_2550_n 0.00223667f $X=15.185 $Y=0.235 $X2=0 $Y2=0
cc_1380 N_Z_M1059_s N_VGND_c_2550_n 0.00231914f $X=16.045 $Y=0.235 $X2=0 $Y2=0
cc_1381 N_Z_c_2250_n N_VGND_c_2550_n 0.0125689f $X=10.165 $Y=0.36 $X2=0 $Y2=0
cc_1382 N_Z_c_2251_n N_VGND_c_2550_n 0.0123859f $X=11.025 $Y=0.36 $X2=0 $Y2=0
cc_1383 N_Z_c_2252_n N_VGND_c_2550_n 0.0123859f $X=11.885 $Y=0.36 $X2=0 $Y2=0
cc_1384 N_Z_c_2253_n N_VGND_c_2550_n 0.0123859f $X=12.745 $Y=0.36 $X2=0 $Y2=0
cc_1385 N_Z_c_2254_n N_VGND_c_2550_n 0.0123859f $X=13.605 $Y=0.36 $X2=0 $Y2=0
cc_1386 N_Z_c_2255_n N_VGND_c_2550_n 0.0123859f $X=14.465 $Y=0.36 $X2=0 $Y2=0
cc_1387 N_Z_c_2256_n N_VGND_c_2550_n 0.0123555f $X=15.325 $Y=0.36 $X2=0 $Y2=0
cc_1388 N_Z_c_2257_n N_VGND_c_2550_n 0.0125689f $X=16.185 $Y=0.36 $X2=0 $Y2=0
cc_1389 N_Z_c_2250_n N_A_1451_47#_c_2760_n 0.0290655f $X=10.165 $Y=0.36 $X2=0
+ $Y2=0
cc_1390 N_VGND_c_2550_n N_A_1451_47#_M1002_s 0.0023412f $X=17.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1391 N_VGND_c_2550_n N_A_1451_47#_M1003_s 0.00480313f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1392 N_VGND_c_2550_n N_A_1451_47#_M1039_s 0.00253158f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1393 N_VGND_M1002_d N_A_1451_47#_c_2757_n 0.00180746f $X=7.69 $Y=0.235 $X2=0
+ $Y2=0
cc_1394 N_VGND_c_2520_n N_A_1451_47#_c_2757_n 0.0139831f $X=7.83 $Y=0.48 $X2=0
+ $Y2=0
cc_1395 N_VGND_c_2533_n N_A_1451_47#_c_2788_n 0.0197971f $X=10.51 $Y=0 $X2=0
+ $Y2=0
cc_1396 N_VGND_c_2550_n N_A_1451_47#_c_2788_n 0.0125699f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1397 N_VGND_c_2533_n N_A_1451_47#_c_2762_n 0.0375436f $X=10.51 $Y=0 $X2=0
+ $Y2=0
cc_1398 N_VGND_c_2550_n N_A_1451_47#_c_2762_n 0.0253849f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1399 N_VGND_c_2519_n N_A_1451_47#_c_2759_n 0.0113657f $X=6.84 $Y=0.38 $X2=0
+ $Y2=0
cc_1400 N_VGND_c_2548_n N_A_1451_47#_c_2759_n 0.0153859f $X=7.745 $Y=0 $X2=0
+ $Y2=0
cc_1401 N_VGND_c_2550_n N_A_1451_47#_c_2759_n 0.0119195f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1402 N_VGND_c_2533_n N_A_1451_47#_c_2760_n 0.0165434f $X=10.51 $Y=0 $X2=0
+ $Y2=0
cc_1403 N_VGND_c_2550_n N_A_1451_47#_c_2760_n 0.00967329f $X=17.52 $Y=0 $X2=0
+ $Y2=0
