* File: sky130_fd_sc_lp__a2bb2oi_1.pxi.spice
* Created: Fri Aug 28 09:56:38 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2OI_1%A1_N N_A1_N_M1003_g N_A1_N_M1005_g A1_N A1_N
+ N_A1_N_c_58_n N_A1_N_c_59_n PM_SKY130_FD_SC_LP__A2BB2OI_1%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_1%A2_N N_A2_N_c_82_n N_A2_N_M1008_g N_A2_N_c_83_n
+ N_A2_N_M1006_g A2_N PM_SKY130_FD_SC_LP__A2BB2OI_1%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_1%A_113_47# N_A_113_47#_M1003_d
+ N_A_113_47#_M1008_d N_A_113_47#_M1001_g N_A_113_47#_M1002_g
+ N_A_113_47#_c_174_p N_A_113_47#_c_131_n N_A_113_47#_c_126_n
+ N_A_113_47#_c_122_n N_A_113_47#_c_123_n N_A_113_47#_c_124_n
+ N_A_113_47#_c_116_n N_A_113_47#_c_117_n N_A_113_47#_c_118_n
+ N_A_113_47#_c_119_n N_A_113_47#_c_120_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_1%A_113_47#
x_PM_SKY130_FD_SC_LP__A2BB2OI_1%B2 N_B2_M1007_g N_B2_M1009_g B2 B2 N_B2_c_186_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_1%B2
x_PM_SKY130_FD_SC_LP__A2BB2OI_1%B1 N_B1_M1004_g N_B1_M1000_g B1 B1 N_B1_c_227_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_1%B1
x_PM_SKY130_FD_SC_LP__A2BB2OI_1%VPWR N_VPWR_M1005_s N_VPWR_M1009_d
+ N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_259_n
+ VPWR N_VPWR_c_260_n N_VPWR_c_254_n PM_SKY130_FD_SC_LP__A2BB2OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2OI_1%Y N_Y_M1001_d N_Y_M1002_s N_Y_c_306_n
+ N_Y_c_344_p N_Y_c_319_n N_Y_c_322_n N_Y_c_299_n N_Y_c_301_n Y Y
+ PM_SKY130_FD_SC_LP__A2BB2OI_1%Y
x_PM_SKY130_FD_SC_LP__A2BB2OI_1%A_381_367# N_A_381_367#_M1002_d
+ N_A_381_367#_M1000_d N_A_381_367#_c_352_n N_A_381_367#_c_353_n
+ N_A_381_367#_c_354_n N_A_381_367#_c_350_n N_A_381_367#_c_351_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_1%A_381_367#
x_PM_SKY130_FD_SC_LP__A2BB2OI_1%VGND N_VGND_M1003_s N_VGND_M1006_d
+ N_VGND_M1004_d N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n
+ VGND N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_1%VGND
cc_1 VNB N_A1_N_M1005_g 0.00640496f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=2.465
cc_2 VNB A1_N 0.0249249f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A1_N_c_58_n 0.0369149f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.375
cc_4 VNB N_A1_N_c_59_n 0.0214535f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.185
cc_5 VNB N_A2_N_c_82_n 0.0524722f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.185
cc_6 VNB N_A2_N_c_83_n 0.0195558f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.54
cc_7 VNB A2_N 0.00788829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_113_47#_M1002_g 0.00867823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_113_47#_c_116_n 0.00265633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_113_47#_c_117_n 0.0022716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_113_47#_c_118_n 0.0325233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_113_47#_c_119_n 0.00257608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_113_47#_c_120_n 0.018655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B2_M1007_g 0.0188303f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_15 VNB N_B2_M1009_g 0.00536644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB B2 0.00555619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B2_c_186_n 0.0313658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_M1004_g 0.0245313f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.655
cc_19 VNB N_B1_M1000_g 0.00623375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB B1 0.0235085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B1_c_227_n 0.0489198f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.375
cc_22 VNB N_VPWR_c_254_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_299_n 0.0039715f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.375
cc_24 VNB N_VGND_c_373_n 0.0108441f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_25 VNB N_VGND_c_374_n 0.0340274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_375_n 0.0126576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_376_n 0.0357914f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.375
cc_28 VNB N_VGND_c_377_n 0.0334572f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.48
cc_29 VNB N_VGND_c_378_n 0.0129339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_379_n 0.0157645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_380_n 0.190802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_A1_N_M1005_g 0.0244891f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=2.465
cc_33 VPB A1_N 0.0175471f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_34 VPB N_A2_N_c_82_n 0.0295483f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.185
cc_35 VPB N_A_113_47#_M1002_g 0.0239794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A_113_47#_c_122_n 0.00475187f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.54
cc_37 VPB N_A_113_47#_c_123_n 0.00911439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_113_47#_c_124_n 0.0172341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_113_47#_c_116_n 7.45301e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_B2_M1009_g 0.0207675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB B2 0.00349556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_B1_M1000_g 0.0256859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB B1 0.0108573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_255_n 0.0108182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_256_n 0.0484537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_257_n 0.00552868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_258_n 0.0516498f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.375
cc_48 VPB N_VPWR_c_259_n 0.0063159f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.185
cc_49 VPB N_VPWR_c_260_n 0.0197638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_254_n 0.0564846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_Y_c_299_n 0.00144614f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.375
cc_52 VPB N_Y_c_301_n 0.00191279f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.375
cc_53 VPB Y 0.00804254f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.54
cc_54 VPB N_A_381_367#_c_350_n 0.0171739f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.375
cc_55 VPB N_A_381_367#_c_351_n 0.0278252f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.54
cc_56 A1_N N_A2_N_c_82_n 0.00960535f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_57 N_A1_N_c_58_n N_A2_N_c_82_n 0.105228f $X=0.4 $Y=1.375 $X2=-0.19 $Y2=-0.245
cc_58 N_A1_N_c_59_n N_A2_N_c_83_n 0.0149993f $X=0.4 $Y=1.185 $X2=0 $Y2=0
cc_59 A1_N A2_N 0.0247656f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_60 N_A1_N_c_58_n A2_N 3.27212e-19 $X=0.4 $Y=1.375 $X2=0 $Y2=0
cc_61 A1_N N_A_113_47#_c_126_n 0.014492f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A1_N_M1005_g N_A_113_47#_c_122_n 4.87595e-19 $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_63 A1_N N_A_113_47#_c_122_n 0.00465617f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A1_N_M1005_g N_A_113_47#_c_123_n 0.00280141f $X=0.49 $Y=2.465 $X2=0
+ $Y2=0
cc_65 N_A1_N_M1005_g N_VPWR_c_256_n 0.029059f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_66 A1_N N_VPWR_c_256_n 0.0267909f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A1_N_c_58_n N_VPWR_c_256_n 7.65393e-19 $X=0.4 $Y=1.375 $X2=0 $Y2=0
cc_68 N_A1_N_M1005_g N_VPWR_c_258_n 0.00486043f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_69 N_A1_N_M1005_g N_VPWR_c_254_n 0.00827383f $X=0.49 $Y=2.465 $X2=0 $Y2=0
cc_70 A1_N N_VGND_c_374_n 0.0260006f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_A1_N_c_58_n N_VGND_c_374_n 0.00420175f $X=0.4 $Y=1.375 $X2=0 $Y2=0
cc_72 N_A1_N_c_59_n N_VGND_c_374_n 0.0156236f $X=0.4 $Y=1.185 $X2=0 $Y2=0
cc_73 N_A1_N_c_59_n N_VGND_c_378_n 0.00486043f $X=0.4 $Y=1.185 $X2=0 $Y2=0
cc_74 N_A1_N_c_59_n N_VGND_c_379_n 5.85381e-19 $X=0.4 $Y=1.185 $X2=0 $Y2=0
cc_75 N_A1_N_c_59_n N_VGND_c_380_n 0.0082726f $X=0.4 $Y=1.185 $X2=0 $Y2=0
cc_76 N_A2_N_c_82_n N_A_113_47#_M1002_g 0.00257977f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_77 N_A2_N_c_82_n N_A_113_47#_c_131_n 0.00219301f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_78 N_A2_N_c_83_n N_A_113_47#_c_131_n 0.0157505f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_79 A2_N N_A_113_47#_c_131_n 0.0283954f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A2_N_c_82_n N_A_113_47#_c_122_n 0.0178078f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_81 A2_N N_A_113_47#_c_122_n 0.0222787f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A2_N_c_82_n N_A_113_47#_c_123_n 0.0204471f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_83 N_A2_N_c_82_n N_A_113_47#_c_124_n 4.50292e-19 $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_84 A2_N N_A_113_47#_c_124_n 0.00917773f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A2_N_c_82_n N_A_113_47#_c_116_n 0.00334203f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_86 N_A2_N_c_82_n N_A_113_47#_c_118_n 0.0181945f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_87 A2_N N_A_113_47#_c_118_n 0.00113621f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A2_N_c_82_n N_A_113_47#_c_119_n 9.63909e-19 $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_89 N_A2_N_c_83_n N_A_113_47#_c_119_n 0.00387929f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_90 A2_N N_A_113_47#_c_119_n 0.0278944f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A2_N_c_82_n N_VPWR_c_256_n 0.00445595f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_92 N_A2_N_c_82_n N_VPWR_c_258_n 0.0054895f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_93 N_A2_N_c_82_n N_VPWR_c_254_n 0.0112391f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_94 N_A2_N_c_82_n N_Y_c_301_n 3.85331e-19 $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_95 N_A2_N_c_82_n Y 0.00172197f $X=0.88 $Y=1.725 $X2=0 $Y2=0
cc_96 N_A2_N_c_83_n N_VGND_c_374_n 6.16708e-19 $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_97 N_A2_N_c_83_n N_VGND_c_378_n 0.00486043f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_98 N_A2_N_c_83_n N_VGND_c_379_n 0.0131037f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_99 N_A2_N_c_83_n N_VGND_c_380_n 0.00455762f $X=0.92 $Y=1.185 $X2=0 $Y2=0
cc_100 N_A_113_47#_c_120_n N_B2_M1007_g 0.014916f $X=1.735 $Y=1.185 $X2=0 $Y2=0
cc_101 N_A_113_47#_M1002_g N_B2_M1009_g 0.0417522f $X=1.83 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_113_47#_c_124_n B2 0.003065f $X=1.555 $Y=1.78 $X2=0 $Y2=0
cc_103 N_A_113_47#_c_116_n B2 0.00900112f $X=1.645 $Y=1.695 $X2=0 $Y2=0
cc_104 N_A_113_47#_c_117_n B2 0.025042f $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_105 N_A_113_47#_c_118_n B2 0.00387454f $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_106 N_A_113_47#_c_117_n N_B2_c_186_n 3.25918e-19 $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_107 N_A_113_47#_c_118_n N_B2_c_186_n 0.0173002f $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_108 N_A_113_47#_c_122_n N_VPWR_c_256_n 0.00523904f $X=1.095 $Y=2.085 $X2=0
+ $Y2=0
cc_109 N_A_113_47#_c_123_n N_VPWR_c_256_n 0.031348f $X=1.095 $Y=2.95 $X2=0 $Y2=0
cc_110 N_A_113_47#_M1002_g N_VPWR_c_258_n 0.0055654f $X=1.83 $Y=2.465 $X2=0
+ $Y2=0
cc_111 N_A_113_47#_c_123_n N_VPWR_c_258_n 0.0210467f $X=1.095 $Y=2.95 $X2=0
+ $Y2=0
cc_112 N_A_113_47#_M1008_d N_VPWR_c_254_n 0.00215158f $X=0.955 $Y=1.835 $X2=0
+ $Y2=0
cc_113 N_A_113_47#_M1002_g N_VPWR_c_254_n 0.0114353f $X=1.83 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_113_47#_c_123_n N_VPWR_c_254_n 0.0125689f $X=1.095 $Y=2.95 $X2=0
+ $Y2=0
cc_115 N_A_113_47#_c_124_n N_Y_M1002_s 0.00253546f $X=1.555 $Y=1.78 $X2=0 $Y2=0
cc_116 N_A_113_47#_M1002_g N_Y_c_306_n 0.0132041f $X=1.83 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_113_47#_c_117_n N_Y_c_306_n 0.00338796f $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_118 N_A_113_47#_M1002_g N_Y_c_301_n 8.15255e-19 $X=1.83 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_113_47#_c_122_n N_Y_c_301_n 0.00410523f $X=1.095 $Y=2.085 $X2=0 $Y2=0
cc_120 N_A_113_47#_c_123_n N_Y_c_301_n 0.00977311f $X=1.095 $Y=2.95 $X2=0 $Y2=0
cc_121 N_A_113_47#_c_124_n N_Y_c_301_n 0.0215234f $X=1.555 $Y=1.78 $X2=0 $Y2=0
cc_122 N_A_113_47#_c_117_n N_Y_c_301_n 9.2046e-19 $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_123 N_A_113_47#_c_118_n N_Y_c_301_n 5.84327e-19 $X=1.73 $Y=1.35 $X2=0 $Y2=0
cc_124 N_A_113_47#_M1002_g Y 0.0103255f $X=1.83 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_113_47#_c_123_n Y 0.0668764f $X=1.095 $Y=2.95 $X2=0 $Y2=0
cc_126 N_A_113_47#_c_131_n N_VGND_M1006_d 0.0207784f $X=1.555 $Y=0.93 $X2=0
+ $Y2=0
cc_127 N_A_113_47#_c_119_n N_VGND_M1006_d 9.63639e-19 $X=1.725 $Y=1.2 $X2=0
+ $Y2=0
cc_128 N_A_113_47#_c_120_n N_VGND_c_377_n 0.00486043f $X=1.735 $Y=1.185 $X2=0
+ $Y2=0
cc_129 N_A_113_47#_c_174_p N_VGND_c_378_n 0.0124525f $X=0.705 $Y=0.42 $X2=0
+ $Y2=0
cc_130 N_A_113_47#_c_131_n N_VGND_c_379_n 0.0541574f $X=1.555 $Y=0.93 $X2=0
+ $Y2=0
cc_131 N_A_113_47#_c_117_n N_VGND_c_379_n 0.00106886f $X=1.73 $Y=1.35 $X2=0
+ $Y2=0
cc_132 N_A_113_47#_c_118_n N_VGND_c_379_n 5.94635e-19 $X=1.73 $Y=1.35 $X2=0
+ $Y2=0
cc_133 N_A_113_47#_c_120_n N_VGND_c_379_n 0.0146171f $X=1.735 $Y=1.185 $X2=0
+ $Y2=0
cc_134 N_A_113_47#_M1003_d N_VGND_c_380_n 0.00408812f $X=0.565 $Y=0.235 $X2=0
+ $Y2=0
cc_135 N_A_113_47#_c_174_p N_VGND_c_380_n 0.00730901f $X=0.705 $Y=0.42 $X2=0
+ $Y2=0
cc_136 N_A_113_47#_c_131_n N_VGND_c_380_n 0.00738659f $X=1.555 $Y=0.93 $X2=0
+ $Y2=0
cc_137 N_A_113_47#_c_120_n N_VGND_c_380_n 0.00822376f $X=1.735 $Y=1.185 $X2=0
+ $Y2=0
cc_138 N_B2_M1007_g N_B1_M1004_g 0.0329654f $X=2.26 $Y=0.655 $X2=0 $Y2=0
cc_139 N_B2_M1009_g N_B1_M1000_g 0.040305f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_140 B2 N_B1_M1000_g 5.52591e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_141 B2 N_B1_c_227_n 2.88683e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_142 N_B2_c_186_n N_B1_c_227_n 0.0172446f $X=2.31 $Y=1.375 $X2=0 $Y2=0
cc_143 N_B2_M1009_g N_VPWR_c_257_n 0.00540239f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_144 N_B2_M1009_g N_VPWR_c_258_n 0.0055654f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_145 N_B2_M1009_g N_VPWR_c_254_n 0.00637182f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_146 N_B2_M1009_g N_Y_c_306_n 0.0116934f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_147 B2 N_Y_c_306_n 0.0151805f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_148 N_B2_c_186_n N_Y_c_306_n 0.00205732f $X=2.31 $Y=1.375 $X2=0 $Y2=0
cc_149 N_B2_M1007_g N_Y_c_319_n 0.0105164f $X=2.26 $Y=0.655 $X2=0 $Y2=0
cc_150 B2 N_Y_c_319_n 0.0163287f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_151 N_B2_c_186_n N_Y_c_319_n 0.00298855f $X=2.31 $Y=1.375 $X2=0 $Y2=0
cc_152 B2 N_Y_c_322_n 0.00660675f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_153 N_B2_M1007_g N_Y_c_299_n 0.00339625f $X=2.26 $Y=0.655 $X2=0 $Y2=0
cc_154 N_B2_M1009_g N_Y_c_299_n 0.00636578f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_155 B2 N_Y_c_299_n 0.0423372f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B2_c_186_n N_Y_c_299_n 0.00215547f $X=2.31 $Y=1.375 $X2=0 $Y2=0
cc_157 N_B2_M1009_g Y 7.73936e-19 $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B2_M1009_g N_A_381_367#_c_352_n 0.0071006f $X=2.265 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_B2_M1009_g N_A_381_367#_c_353_n 0.00933636f $X=2.265 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_B2_M1009_g N_A_381_367#_c_354_n 5.65405e-19 $X=2.265 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_B2_M1009_g N_A_381_367#_c_351_n 5.91026e-19 $X=2.265 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_B2_M1007_g N_VGND_c_377_n 0.00585385f $X=2.26 $Y=0.655 $X2=0 $Y2=0
cc_163 N_B2_M1007_g N_VGND_c_379_n 0.00127567f $X=2.26 $Y=0.655 $X2=0 $Y2=0
cc_164 N_B2_M1007_g N_VGND_c_380_n 0.0067966f $X=2.26 $Y=0.655 $X2=0 $Y2=0
cc_165 N_B1_M1000_g N_VPWR_c_257_n 0.00364709f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_166 N_B1_M1000_g N_VPWR_c_260_n 0.00571722f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_167 N_B1_M1000_g N_VPWR_c_254_n 0.00736442f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_168 N_B1_M1000_g N_Y_c_306_n 0.0042002f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_169 N_B1_M1004_g N_Y_c_319_n 0.00530799f $X=2.79 $Y=0.655 $X2=0 $Y2=0
cc_170 N_B1_M1004_g N_Y_c_299_n 0.00864043f $X=2.79 $Y=0.655 $X2=0 $Y2=0
cc_171 N_B1_M1000_g N_Y_c_299_n 0.0146561f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_172 B1 N_Y_c_299_n 0.0404283f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_173 N_B1_c_227_n N_Y_c_299_n 0.00804595f $X=3.01 $Y=1.375 $X2=0 $Y2=0
cc_174 N_B1_M1000_g N_A_381_367#_c_352_n 4.10339e-19 $X=2.815 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_B1_M1000_g N_A_381_367#_c_353_n 0.0137932f $X=2.815 $Y=2.465 $X2=0
+ $Y2=0
cc_176 B1 N_A_381_367#_c_350_n 0.0238189f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_177 N_B1_c_227_n N_A_381_367#_c_350_n 0.00118142f $X=3.01 $Y=1.375 $X2=0
+ $Y2=0
cc_178 N_B1_M1000_g N_A_381_367#_c_351_n 0.00761777f $X=2.815 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_B1_M1004_g N_VGND_c_376_n 0.0205308f $X=2.79 $Y=0.655 $X2=0 $Y2=0
cc_180 B1 N_VGND_c_376_n 0.0232162f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_181 N_B1_c_227_n N_VGND_c_376_n 0.00197077f $X=3.01 $Y=1.375 $X2=0 $Y2=0
cc_182 N_B1_M1004_g N_VGND_c_377_n 0.00585385f $X=2.79 $Y=0.655 $X2=0 $Y2=0
cc_183 N_B1_M1004_g N_VGND_c_380_n 0.0111642f $X=2.79 $Y=0.655 $X2=0 $Y2=0
cc_184 N_VPWR_c_254_n A_113_367# 0.010279f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_185 N_VPWR_c_254_n N_Y_M1002_s 0.00215158f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_186 N_VPWR_M1009_d N_Y_c_306_n 0.00839356f $X=2.34 $Y=1.835 $X2=0 $Y2=0
cc_187 N_VPWR_M1009_d N_Y_c_299_n 0.00242173f $X=2.34 $Y=1.835 $X2=0 $Y2=0
cc_188 N_VPWR_c_258_n Y 0.0207058f $X=2.38 $Y=3.33 $X2=0 $Y2=0
cc_189 N_VPWR_c_254_n Y 0.0123974f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_190 N_VPWR_c_254_n N_A_381_367#_M1002_d 0.0036673f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_191 N_VPWR_c_254_n N_A_381_367#_M1000_d 0.00215158f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_258_n N_A_381_367#_c_352_n 0.0159044f $X=2.38 $Y=3.33 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_254_n N_A_381_367#_c_352_n 0.0100725f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_194 N_VPWR_M1009_d N_A_381_367#_c_353_n 0.00639101f $X=2.34 $Y=1.835 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_257_n N_A_381_367#_c_353_n 0.0226964f $X=2.545 $Y=2.83 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_254_n N_A_381_367#_c_353_n 0.0114824f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_260_n N_A_381_367#_c_351_n 0.0200252f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_254_n N_A_381_367#_c_351_n 0.0120553f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_199 N_Y_c_306_n N_A_381_367#_M1002_d 0.00668805f $X=2.575 $Y=2.12 $X2=-0.19
+ $Y2=-0.245
cc_200 N_Y_c_306_n N_A_381_367#_c_353_n 0.0307506f $X=2.575 $Y=2.12 $X2=0 $Y2=0
cc_201 N_Y_c_306_n N_A_381_367#_c_354_n 0.0154301f $X=2.575 $Y=2.12 $X2=0 $Y2=0
cc_202 N_Y_c_319_n N_VGND_c_376_n 0.0132054f $X=2.575 $Y=0.945 $X2=0 $Y2=0
cc_203 N_Y_c_299_n N_VGND_c_376_n 6.64331e-19 $X=2.66 $Y=2.035 $X2=0 $Y2=0
cc_204 N_Y_c_344_p N_VGND_c_377_n 0.0128073f $X=2.045 $Y=0.42 $X2=0 $Y2=0
cc_205 N_Y_M1001_d N_VGND_c_380_n 0.00402866f $X=1.905 $Y=0.235 $X2=0 $Y2=0
cc_206 N_Y_c_344_p N_VGND_c_380_n 0.00769778f $X=2.045 $Y=0.42 $X2=0 $Y2=0
cc_207 N_Y_c_319_n N_VGND_c_380_n 0.0196291f $X=2.575 $Y=0.945 $X2=0 $Y2=0
cc_208 N_Y_c_319_n A_467_47# 0.0106186f $X=2.575 $Y=0.945 $X2=-0.19 $Y2=-0.245
cc_209 N_Y_c_299_n A_467_47# 5.37627e-19 $X=2.66 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_210 N_VGND_c_380_n A_467_47# 0.00568775f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
