* File: sky130_fd_sc_lp__a32oi_2.spice
* Created: Wed Sep  2 09:28:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32oi_2.pex.spice"
.subckt sky130_fd_sc_lp__a32oi_2  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_B2_M1012_g N_A_43_65#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1012_d N_B2_M1013_g N_A_43_65#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_43_65#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1003_d N_B1_M1009_g N_A_43_65#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2814 PD=1.12 PS=2.35 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.5
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1007 N_Y_M1007_d N_A1_M1007_g N_A_509_65#_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2814 PD=1.12 PS=2.35 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.3
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1015 N_Y_M1007_d N_A1_M1015_g N_A_509_65#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_A_778_65#_M1004_d N_A2_M1004_g N_A_509_65#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1010 N_A_778_65#_M1004_d N_A2_M1010_g N_A_509_65#_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2814 PD=1.12 PS=2.35 NRD=0 NRS=9.996 M=1 R=5.6
+ SA=75001.6 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A3_M1006_g N_A_778_65#_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1017_d N_A3_M1017_g N_A_778_65#_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_B2_M1005_g N_A_43_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.2 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1005_d N_B2_M1011_g N_A_43_367#_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.8 A=0.189 P=2.82 MULT=1
MM1000 N_A_43_367#_M1011_s N_B1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1008 N_A_43_367#_M1008_d N_B1_M1008_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.32445 AS=0.1764 PD=1.775 PS=1.54 NRD=18.7544 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.9 A=0.189 P=2.82 MULT=1
MM1016 N_A_43_367#_M1008_d N_A1_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.32445 AS=0.45675 PD=1.775 PS=1.985 NRD=17.9664 NRS=0 M=1 R=8.4 SA=75002.1
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1019 N_A_43_367#_M1019_d N_A1_M1019_g N_VPWR_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.45675 PD=1.62 PS=1.985 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75003
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1002 N_A_43_367#_M1019_d N_A2_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.4095 PD=1.62 PS=1.91 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75003.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1018 N_A_43_367#_M1018_d N_A2_M1018_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.4095 PD=1.54 PS=1.91 NRD=0 NRS=0 M=1 R=8.4 SA=75004.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1001 N_A_43_367#_M1018_d N_A3_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_A_43_367#_M1014_d N_A3_M1014_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3463 P=16.97
*
.include "sky130_fd_sc_lp__a32oi_2.pxi.spice"
*
.ends
*
*
