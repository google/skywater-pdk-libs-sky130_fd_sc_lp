* File: sky130_fd_sc_lp__a21boi_0.pex.spice
* Created: Wed Sep  2 09:19:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BOI_0%B1_N 3 6 9 11 12 13 14 19
r37 19 21 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.84
+ $X2=0.597 $Y2=1.675
r38 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.84 $X2=0.63 $Y2=1.84
r39 13 14 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.712 $Y=2.035
+ $X2=0.712 $Y2=2.405
r40 13 20 5.9927 $w=3.73e-07 $l=1.95e-07 $layer=LI1_cond $X=0.712 $Y=2.035
+ $X2=0.712 $Y2=1.84
r41 12 20 5.37807 $w=3.73e-07 $l=1.75e-07 $layer=LI1_cond $X=0.712 $Y=1.665
+ $X2=0.712 $Y2=1.84
r42 9 11 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.475 $Y=2.77
+ $X2=0.475 $Y2=2.345
r43 6 11 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.597 $Y=2.148
+ $X2=0.597 $Y2=2.345
r44 5 19 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.597 $Y=1.872
+ $X2=0.597 $Y2=1.84
r45 5 6 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.597 $Y=1.872
+ $X2=0.597 $Y2=2.148
r46 3 21 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_0%A_27_47# 1 2 7 8 9 11 12 13 16 20 24 28 31
c65 8 0 1.6887e-19 $X=1.16 $Y=2.115
c66 7 0 1.73834e-19 $X=1.16 $Y=1.435
r67 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=0.93 $X2=0.925 $Y2=0.93
r68 26 31 1.34785 $w=6.15e-07 $l=1.43e-07 $layer=LI1_cond $X=0.38 $Y=1.087
+ $X2=0.237 $Y2=1.087
r69 26 28 10.5994 $w=6.13e-07 $l=5.45e-07 $layer=LI1_cond $X=0.38 $Y=1.087
+ $X2=0.925 $Y2=1.087
r70 22 31 9.54454 $w=2.72e-07 $l=3.13943e-07 $layer=LI1_cond $X=0.225 $Y=1.395
+ $X2=0.237 $Y2=1.087
r71 22 24 62.0546 $w=2.58e-07 $l=1.4e-06 $layer=LI1_cond $X=0.225 $Y=1.395
+ $X2=0.225 $Y2=2.795
r72 18 31 9.54454 $w=2.72e-07 $l=3.07e-07 $layer=LI1_cond $X=0.237 $Y=0.78
+ $X2=0.237 $Y2=1.087
r73 18 20 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=0.237 $Y=0.78
+ $X2=0.237 $Y2=0.445
r74 14 16 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.545 $Y=2.265 $X2=1.545
+ $Y2=2.735
r75 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.47 $Y=2.19
+ $X2=1.545 $Y2=2.265
r76 12 13 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=1.47 $Y=2.19
+ $X2=1.235 $Y2=2.19
r77 9 29 42.0031 $w=5.03e-07 $l=2.75409e-07 $layer=POLY_cond $X=1.245 $Y=0.765
+ $X2=1.04 $Y2=0.93
r78 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.245 $Y=0.765
+ $X2=1.245 $Y2=0.445
r79 8 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.16 $Y=2.115
+ $X2=1.235 $Y2=2.19
r80 7 29 74.5836 $w=5.03e-07 $l=5.61805e-07 $layer=POLY_cond $X=1.16 $Y=1.435
+ $X2=1.04 $Y2=0.93
r81 7 8 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.16 $Y=1.435 $X2=1.16
+ $Y2=2.115
r82 2 24 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.56 $X2=0.26 $Y2=2.795
r83 1 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_0%A1 3 5 7 9 10 11
c43 9 0 1.73834e-19 $X=2.16 $Y=0.925
c44 5 0 1.00938e-19 $X=1.975 $Y=1.875
c45 3 0 1.95047e-19 $X=1.675 $Y=0.445
r46 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.885
+ $Y=1.37 $X2=1.885 $Y2=1.37
r47 11 17 6.5952 $w=5.33e-07 $l=2.95e-07 $layer=LI1_cond $X=1.987 $Y=1.665
+ $X2=1.987 $Y2=1.37
r48 10 17 1.67675 $w=5.33e-07 $l=7.5e-08 $layer=LI1_cond $X=1.987 $Y=1.295
+ $X2=1.987 $Y2=1.37
r49 9 10 8.27194 $w=5.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.987 $Y=0.925
+ $X2=1.987 $Y2=1.295
r50 5 16 73.5676 $w=5.32e-07 $l=5.93709e-07 $layer=POLY_cond $X=1.975 $Y=1.875
+ $X2=1.782 $Y2=1.37
r51 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.975 $Y=1.875
+ $X2=1.975 $Y2=2.735
r52 1 16 43.2161 $w=5.32e-07 $l=2.17002e-07 $layer=POLY_cond $X=1.675 $Y=1.2
+ $X2=1.782 $Y2=1.37
r53 1 3 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.675 $Y=1.2
+ $X2=1.675 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_0%A2 3 5 6 9 13 14 15 16 21
c34 14 0 1.95047e-19 $X=2.64 $Y=0.925
r35 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.51
+ $Y=1.005 $X2=2.51 $Y2=1.005
r36 15 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=1.295
+ $X2=2.61 $Y2=1.665
r37 15 22 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.61 $Y=1.295
+ $X2=2.61 $Y2=1.005
r38 14 22 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=2.61 $Y=0.925 $X2=2.61
+ $Y2=1.005
r39 12 21 55.6971 $w=3.45e-07 $l=3.33e-07 $layer=POLY_cond $X=2.502 $Y=1.338
+ $X2=2.502 $Y2=1.005
r40 12 13 47.5363 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=2.502 $Y=1.338
+ $X2=2.502 $Y2=1.51
r41 11 21 6.69034 $w=3.45e-07 $l=4e-08 $layer=POLY_cond $X=2.502 $Y=0.965
+ $X2=2.502 $Y2=1.005
r42 9 13 628.138 $w=1.5e-07 $l=1.225e-06 $layer=POLY_cond $X=2.405 $Y=2.735
+ $X2=2.405 $Y2=1.51
r43 5 11 32.7621 $w=1.5e-07 $l=2.06116e-07 $layer=POLY_cond $X=2.33 $Y=0.89
+ $X2=2.502 $Y2=0.965
r44 5 6 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.33 $Y=0.89 $X2=2.11
+ $Y2=0.89
r45 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.035 $Y=0.815
+ $X2=2.11 $Y2=0.89
r46 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.035 $Y=0.815
+ $X2=2.035 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_0%VPWR 1 2 9 13 15 17 22 29 30 33 36
r37 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 27 36 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.187 $Y2=3.33
r42 27 29 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.32 $Y=3.33 $X2=2.64
+ $Y2=3.33
r43 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r46 23 25 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 22 36 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.055 $Y=3.33
+ $X2=2.187 $Y2=3.33
r48 22 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.055 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r52 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 11 36 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.187 $Y=3.245
+ $X2=2.187 $Y2=3.33
r56 11 13 29.3547 $w=2.63e-07 $l=6.75e-07 $layer=LI1_cond $X=2.187 $Y=3.245
+ $X2=2.187 $Y2=2.57
r57 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r58 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.795
r59 2 13 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=2.415 $X2=2.19 $Y2=2.57
r60 1 9 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.56 $X2=0.69 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_0%Y 1 2 10 13 14 15 16 32
r36 16 27 5.97049 $w=4.13e-07 $l=2.15e-07 $layer=LI1_cond $X=1.277 $Y=2.775
+ $X2=1.277 $Y2=2.56
r37 15 27 4.30431 $w=4.13e-07 $l=1.55e-07 $layer=LI1_cond $X=1.277 $Y=2.405
+ $X2=1.277 $Y2=2.56
r38 14 15 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.277 $Y=2.035
+ $X2=1.277 $Y2=2.405
r39 14 21 7.30343 $w=4.13e-07 $l=2.63e-07 $layer=LI1_cond $X=1.277 $Y=2.035
+ $X2=1.277 $Y2=1.772
r40 13 21 2.97136 $w=4.13e-07 $l=1.07e-07 $layer=LI1_cond $X=1.277 $Y=1.665
+ $X2=1.277 $Y2=1.772
r41 13 32 6.90831 $w=4.13e-07 $l=1e-07 $layer=LI1_cond $X=1.277 $Y=1.665
+ $X2=1.277 $Y2=1.565
r42 12 32 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.4 $Y=0.61 $X2=1.4
+ $Y2=1.565
r43 10 12 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=0.445
+ $X2=1.47 $Y2=0.61
r44 2 27 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.205
+ $Y=2.415 $X2=1.33 $Y2=2.56
r45 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.32
+ $Y=0.235 $X2=1.46 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_0%A_324_483# 1 2 9 11 12 15
c24 12 0 1.6887e-19 $X=1.885 $Y=2.14
c25 11 0 1.00938e-19 $X=2.49 $Y=2.14
r26 13 15 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=2.637 $Y=2.225
+ $X2=2.637 $Y2=2.56
r27 11 13 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=2.49 $Y=2.14
+ $X2=2.637 $Y2=2.225
r28 11 12 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.49 $Y=2.14
+ $X2=1.885 $Y2=2.14
r29 7 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.77 $Y=2.225
+ $X2=1.885 $Y2=2.14
r30 7 9 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.77 $Y=2.225
+ $X2=1.77 $Y2=2.56
r31 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=2.415 $X2=2.62 $Y2=2.56
r32 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.62
+ $Y=2.415 $X2=1.76 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_0%VGND 1 2 9 11 13 18 25 26 36
r35 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r36 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r37 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.25
+ $Y2=0
r39 23 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.64
+ $Y2=0
r40 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r41 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 19 21 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.145 $Y=0 $X2=1.2
+ $Y2=0
r43 18 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.25
+ $Y2=0
r44 18 21 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=1.2
+ $Y2=0
r45 16 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r46 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 13 33 8.94546 $w=5.93e-07 $l=4.45e-07 $layer=LI1_cond $X=0.847 $Y=0
+ $X2=0.847 $Y2=0.445
r48 13 19 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=0.847 $Y=0 $X2=1.145
+ $Y2=0
r49 13 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r50 13 15 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r51 11 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r52 11 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r53 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=0.085 $X2=2.25
+ $Y2=0
r54 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.25 $Y=0.085 $X2=2.25
+ $Y2=0.445
r55 2 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.11
+ $Y=0.235 $X2=2.25 $Y2=0.445
r56 1 33 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=1.03 $Y2=0.445
.ends

