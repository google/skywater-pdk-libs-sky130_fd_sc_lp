* NGSPICE file created from sky130_fd_sc_lp__o32ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_489_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=6.678e+11p pd=6.1e+06u as=3.78e+11p ps=3.12e+06u
M1001 a_76_69# B2 Y VNB nshort w=840000u l=150000u
+  ad=7.098e+11p pd=6.73e+06u as=2.772e+11p ps=2.34e+06u
M1002 VGND A1 a_76_69# VNB nshort w=840000u l=150000u
+  ad=7.434e+11p pd=5.13e+06u as=0p ps=0u
M1003 VGND A3 a_76_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_159_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1005 Y B2 a_159_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=8.694e+11p pd=3.9e+06u as=0p ps=0u
M1006 a_399_367# A3 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=3.78e+11p pd=3.12e+06u as=0p ps=0u
M1007 a_76_69# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_489_367# A2 a_399_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_76_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

