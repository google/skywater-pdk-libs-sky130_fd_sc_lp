* File: sky130_fd_sc_lp__srsdfrtn_1.spice
* Created: Fri Aug 28 11:33:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__srsdfrtn_1.pex.spice"
.subckt sky130_fd_sc_lp__srsdfrtn_1  VNB VPB SCE D SCD RESET_B CLK_N SLEEP_B
+ VPWR KAPWR Q VGND
* 
* VGND	VGND
* Q	Q
* KAPWR	KAPWR
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* CLK_N	CLK_N
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_SCE_M1001_g N_A_27_55#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.1155 PD=1.38 PS=1.39 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_A_305_97#_M1023_d N_SCE_M1023_g N_noxref_30_M1023_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1155 PD=0.7 PS=1.39 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1040 noxref_31 N_D_M1040_g N_A_305_97#_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 N_noxref_32_M1003_d N_A_27_55#_M1003_g noxref_31 VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_noxref_30_M1022_d N_SCD_M1022_g N_noxref_32_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_742_63#_M1018_g N_A_666_89#_M1018_s VNB NSHORT L=0.15
+ W=0.42 AD=0.09275 AS=0.3513 PD=0.975 PS=3.02 NRD=0 NRS=223.26 M=1 R=2.8
+ SA=75000.3 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1028 N_noxref_32_M1028_d N_RESET_B_M1028_g N_VGND_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.09275 PD=1.41 PS=0.975 NRD=0 NRS=47.376 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1041 N_A_1113_419#_M1041_d N_A_742_63#_M1041_g N_A_1009_107#_M1041_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.3054 PD=0.7 PS=2.68 NRD=0 NRS=192.036 M=1
+ R=2.8 SA=75000.3 SB=75001 A=0.063 P=1.14 MULT=1
MM1045 A_1201_215# N_A_666_89#_M1045_g N_A_1113_419#_M1041_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1034 N_A_305_97#_M1034_d N_A_666_89#_M1034_g A_1201_215# VNB NSHORT L=0.15
+ W=0.42 AD=0.1155 AS=0.0441 PD=1.39 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 A_1373_77# N_A_1343_51#_M1035_g N_A_1009_107#_M1035_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0525 AS=0.1239 PD=0.67 PS=1.43 NRD=19.992 NRS=2.856 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_A_1453_77#_M1012_d N_A_1343_51#_M1012_g A_1373_77# VNB NSHORT L=0.15
+ W=0.42 AD=0.1155 AS=0.0525 PD=1.39 PS=0.67 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_1453_77#_M1007_d N_RESET_B_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1866 PD=0.7 PS=1.8 NRD=0 NRS=31.428 M=1 R=2.8 SA=75000.3
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_A_1724_21#_M1027_g N_A_1453_77#_M1007_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001 A=0.063 P=1.14 MULT=1
MM1048 A_1840_47# N_A_1113_419#_M1048_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1032 N_A_1343_51#_M1032_d N_A_1113_419#_M1032_g A_1840_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1038 A_2198_97# N_CLK_N_M1038_g N_A_742_63#_M1038_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.2666 PD=0.66 PS=2.32 NRD=18.564 NRS=165.636 M=1 R=2.8
+ SA=75000.3 SB=75002 A=0.063 P=1.14 MULT=1
MM1039 A_2276_97# N_SLEEP_B_M1039_g A_2198_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0504 PD=0.63 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75000.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1043 N_VGND_M1043_d N_SLEEP_B_M1043_g A_2276_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.15785 AS=0.0441 PD=1.28 PS=0.63 NRD=91.656 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1006 A_2480_97# N_SLEEP_B_M1006_g N_VGND_M1043_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.15785 PD=0.66 PS=1.28 NRD=18.564 NRS=91.656 M=1 R=2.8
+ SA=75001.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_A_1724_21#_M1020_d N_SLEEP_B_M1020_g A_2480_97# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75002.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1044 N_A_2717_427#_M1044_d N_A_742_63#_M1044_g N_A_1343_51#_M1044_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.151547 AS=0.2048 PD=1.29208 PS=1.92 NRD=6.552 NRS=6.552 M=1
+ R=4.26667 SA=75000.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1013 A_2879_99# N_A_666_89#_M1013_g N_A_2717_427#_M1044_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0994528 PD=0.63 PS=0.847925 NRD=14.28 NRS=32.856 M=1
+ R=2.8 SA=75000.8 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1002 A_2951_99# N_A_666_89#_M1002_g A_2879_99# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0441 PD=0.66 PS=0.63 NRD=18.564 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1051 N_VGND_M1051_d N_A_2999_73#_M1051_g A_2951_99# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 A_3115_99# N_RESET_B_M1008_g N_VGND_M1051_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_2999_73#_M1009_d N_A_2717_427#_M1009_g A_3115_99# VNB NSHORT L=0.15
+ W=0.42 AD=0.168 AS=0.0504 PD=1.64 PS=0.66 NRD=32.856 NRS=18.564 M=1 R=2.8
+ SA=75002.4 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_A_2717_427#_M1036_g N_A_3368_57#_M1036_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0952 AS=0.1197 PD=0.823333 PS=1.41 NRD=32.856 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1033 N_Q_M1033_d N_A_3368_57#_M1033_g N_VGND_M1036_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1904 PD=2.25 PS=1.64667 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_SCE_M1016_g N_A_27_55#_M1016_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=21.5321 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1025 A_247_491# N_SCE_M1025_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.112 PD=0.88 PS=0.99 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1026 N_A_305_97#_M1026_d N_D_M1026_g A_247_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.1
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1004 A_411_491# N_A_27_55#_M1004_g N_A_305_97#_M1026_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1568 AS=0.0896 PD=1.13 PS=0.92 NRD=58.4696 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1052 N_VPWR_M1052_d N_SCD_M1052_g A_411_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1568 PD=1.85 PS=1.13 NRD=0 NRS=58.4696 M=1 R=4.26667 SA=75002.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1021 N_VPWR_M1021_d N_A_742_63#_M1021_g N_A_666_89#_M1021_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.208 AS=0.1824 PD=1.29 PS=1.85 NRD=113.886 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1049 N_A_305_97#_M1049_d N_RESET_B_M1049_g N_VPWR_M1021_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.138023 AS=0.208 PD=1.24981 PS=1.29 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001 SB=75002 A=0.096 P=1.58 MULT=1
MM1000 A_1041_419# N_A_742_63#_M1000_g N_A_305_97#_M1049_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0905774 PD=0.63 PS=0.820189 NRD=23.443 NRS=56.2829 M=1
+ R=2.8 SA=75001.6 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1037 N_A_1113_419#_M1037_d N_A_742_63#_M1037_g A_1041_419# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0979606 AS=0.0441 PD=0.825211 PS=0.63 NRD=53.9386 NRS=23.443 M=1
+ R=2.8 SA=75001.9 SB=75002 A=0.063 P=1.14 MULT=1
MM1053 A_1242_419# N_A_666_89#_M1053_g N_A_1113_419#_M1037_d VPB PHIGHVT L=0.25
+ W=1 AD=0.2575 AS=0.233239 PD=1.515 PS=1.96479 NRD=39.8728 NRS=0 M=1 R=4
+ SA=125001 SB=125001 A=0.25 P=2.5 MULT=1
MM1010 N_KAPWR_M1010_d N_A_1343_51#_M1010_g A_1242_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.65 AS=0.2575 PD=3.3 PS=1.515 NRD=75.8253 NRS=39.8728 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1011 A_1682_341# N_RESET_B_M1011_g N_A_1113_419#_M1011_s VPB PHIGHVT L=0.25
+ W=1 AD=0.105 AS=0.265 PD=1.21 PS=2.53 NRD=9.8303 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1014 N_KAPWR_M1014_d N_A_1724_21#_M1014_g A_1682_341# VPB PHIGHVT L=0.25 W=1
+ AD=0.257612 AS=0.105 PD=1.735 PS=1.21 NRD=39.9122 NRS=9.8303 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1029 N_A_1343_51#_M1029_d N_A_1113_419#_M1029_g N_KAPWR_M1014_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.38375 AS=0.257612 PD=2.91 PS=1.735 NRD=19.6803 NRS=39.9122 M=1
+ R=4 SA=125001 SB=125000 A=0.25 P=2.5 MULT=1
MM1042 N_A_742_63#_M1042_d N_CLK_N_M1042_g N_KAPWR_M1042_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1019 N_KAPWR_M1019_d N_SLEEP_B_M1019_g N_A_742_63#_M1042_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.130888 AS=0.0896 PD=1.07317 PS=0.92 NRD=29.2348 NRS=0 M=1
+ R=4.26667 SA=75000.6 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1017 N_A_1724_21#_M1017_d N_SLEEP_B_M1017_g N_KAPWR_M1019_d VPB PHIGHVT L=0.25
+ W=1 AD=0.265 AS=0.204512 PD=2.53 PS=1.67683 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1050 A_2645_427# N_A_742_63#_M1050_g N_A_2562_427#_M1050_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1030 N_A_2717_427#_M1030_d N_A_742_63#_M1030_g A_2645_427# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0896 AS=0.0441 PD=0.81 PS=0.63 NRD=44.5417 NRS=23.443 M=1 R=2.8
+ SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1015 N_A_1343_51#_M1015_d N_A_666_89#_M1015_g N_A_2717_427#_M1030_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.4494 AS=0.1792 PD=2.75 PS=1.62 NRD=58.6272 NRS=0
+ M=1 R=5.6 SA=75000.6 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1031 N_VPWR_M1031_d N_A_2999_73#_M1031_g N_A_2562_427#_M1031_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_A_2999_73#_M1005_d N_RESET_B_M1005_g N_VPWR_M1031_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1046 N_VPWR_M1046_d N_A_2717_427#_M1046_g N_A_2999_73#_M1005_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1134 AS=0.0588 PD=1.38 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1047 N_VPWR_M1047_d N_A_2717_427#_M1047_g N_A_3368_57#_M1047_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.140429 AS=0.176 PD=1.10821 PS=1.83 NRD=33.0763 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1024 N_Q_M1024_d N_A_3368_57#_M1024_g N_VPWR_M1047_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3465 AS=0.276471 PD=3.07 PS=2.18179 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX54_noxref VNB VPB NWDIODE A=34.6584 P=42.18
c_192 VNB 0 2.94065e-19 $X=0 $Y=0
c_361 VPB 0 1.47946e-19 $X=0 $Y=3.085
c_3074 A_1373_77# 0 2.87822e-20 $X=6.865 $Y=0.385
*
.include "sky130_fd_sc_lp__srsdfrtn_1.pxi.spice"
*
.ends
*
*
