# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xor2_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__xor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.210000 1.765000 1.555000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.455000 1.725000 ;
        RECT 0.085000 1.725000 2.115000 1.895000 ;
        RECT 1.935000 1.345000 2.115000 1.725000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.846300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.040000 0.595000 2.455000 1.165000 ;
        RECT 2.285000 1.165000 2.455000 1.570000 ;
        RECT 2.285000 1.570000 2.735000 1.750000 ;
        RECT 2.505000 1.750000 2.735000 1.795000 ;
        RECT 2.505000 1.795000 2.835000 2.065000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.170000  0.085000 0.430000 1.040000 ;
      RECT 0.170000  2.065000 2.110000 2.235000 ;
      RECT 0.170000  2.235000 0.500000 3.075000 ;
      RECT 0.600000  0.335000 0.860000 0.870000 ;
      RECT 0.600000  0.870000 1.870000 1.040000 ;
      RECT 0.990000  2.405000 1.270000 3.245000 ;
      RECT 1.030000  0.085000 1.360000 0.700000 ;
      RECT 1.440000  2.405000 1.770000 2.575000 ;
      RECT 1.440000  2.575000 3.265000 2.745000 ;
      RECT 1.440000  2.745000 1.770000 3.075000 ;
      RECT 1.700000  0.255000 2.795000 0.425000 ;
      RECT 1.700000  0.425000 1.870000 0.870000 ;
      RECT 1.940000  2.235000 3.235000 2.405000 ;
      RECT 1.965000  2.915000 2.295000 3.245000 ;
      RECT 2.625000  0.425000 2.795000 1.230000 ;
      RECT 2.625000  1.230000 3.235000 1.400000 ;
      RECT 2.905000  1.400000 3.235000 1.625000 ;
      RECT 2.935000  2.745000 3.265000 2.925000 ;
      RECT 2.965000  0.085000 3.215000 1.060000 ;
      RECT 3.065000  1.625000 3.235000 2.235000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__xor2_1
