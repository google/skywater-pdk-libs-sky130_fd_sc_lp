* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_113_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=1.932e+12p pd=1.804e+07u as=1.6212e+12p ps=1.562e+07u
M1001 a_457_367# A2 a_30_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.4112e+12p pd=1.232e+07u as=1.7262e+12p ps=1.534e+07u
M1002 a_113_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=2.1168e+12p pd=1.848e+07u as=2.4318e+12p ps=2.15e+07u
M1004 Y C1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_30_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_113_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1166_65# C1 Y VNB nshort w=840000u l=150000u
+  ad=1.2432e+12p pd=1.136e+07u as=6.3e+11p ps=4.86e+06u
M1009 a_113_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1166_65# B1 a_113_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_113_47# B1 a_1166_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1166_65# C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_30_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A3 a_457_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A2 a_113_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A1 a_113_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y C1 a_1166_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_113_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_30_367# A2 a_457_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A3 a_457_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y C1 a_1166_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_113_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_30_367# A2 a_457_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND A3 a_113_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A1 a_30_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND A1 a_113_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_113_47# B1 a_1166_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A1 a_30_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_457_367# A3 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Y B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Y C1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1166_65# B1 a_113_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_457_367# A2 a_30_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_457_367# A3 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND A3 a_113_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND A2 a_113_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
