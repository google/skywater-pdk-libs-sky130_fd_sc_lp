* NGSPICE file created from sky130_fd_sc_lp__o2111a_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VGND A2 a_517_49# VNB nshort w=840000u l=150000u
+  ad=4.578e+11p pd=4.45e+06u as=7.434e+11p ps=5.13e+06u
M1001 a_80_21# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=8.442e+11p pd=6.38e+06u as=2.3562e+12p ps=1.13e+07u
M1002 a_409_49# C1 a_337_49# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=1.764e+11p ps=2.1e+06u
M1003 VGND a_80_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1004 a_517_49# B1 a_409_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_337_49# D1 a_80_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1006 VPWR C1 a_80_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_685_367# A2 a_80_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1008 VPWR A1 a_685_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_517_49# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_80_21# D1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_80_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

