* File: sky130_fd_sc_lp__xor3_1.pex.spice
* Created: Fri Aug 28 11:37:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XOR3_1%A_86_305# 1 2 3 4 15 19 21 23 24 26 29 31 34
+ 38 39 45 46 49
c103 39 0 1.65079e-19 $X=0.595 $Y=1.69
r104 49 51 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=1.05
+ $X2=4.405 $Y2=1.215
r105 46 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.485 $Y=1.905
+ $X2=4.485 $Y2=1.215
r106 45 47 19.647 $w=6.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.23 $Y=2.07
+ $X2=4.23 $Y2=2.745
r107 45 46 10.6764 $w=6.78e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=2.07
+ $X2=4.23 $Y2=1.905
r108 39 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.69
+ $X2=0.595 $Y2=1.855
r109 39 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.69
+ $X2=0.595 $Y2=1.525
r110 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.69 $X2=0.595 $Y2=1.69
r111 34 47 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.975 $Y=2.895
+ $X2=3.975 $Y2=2.745
r112 32 43 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=2.98
+ $X2=1.605 $Y2=2.98
r113 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.89 $Y=2.98
+ $X2=3.975 $Y2=2.895
r114 31 32 138.31 $w=1.68e-07 $l=2.12e-06 $layer=LI1_cond $X=3.89 $Y=2.98
+ $X2=1.77 $Y2=2.98
r115 27 41 5.50001 $w=2.69e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.565 $Y=1.845
+ $X2=1.605 $Y2=1.93
r116 27 29 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.565 $Y=1.845
+ $X2=1.565 $Y2=1.08
r117 24 43 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=2.895
+ $X2=1.605 $Y2=2.98
r118 24 26 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.605 $Y=2.895
+ $X2=1.605 $Y2=2.2
r119 23 41 9.69525 $w=3.3e-07 $l=2.5e-07 $layer=LI1_cond $X=1.605 $Y=2.18
+ $X2=1.605 $Y2=1.93
r120 23 26 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=1.605 $Y=2.18
+ $X2=1.605 $Y2=2.2
r121 22 38 10.0619 $w=2.91e-07 $l=3.15595e-07 $layer=LI1_cond $X=0.79 $Y=1.93
+ $X2=0.615 $Y2=1.69
r122 21 41 3.42229 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.44 $Y=1.93
+ $X2=1.605 $Y2=1.93
r123 21 22 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.44 $Y=1.93
+ $X2=0.79 $Y2=1.93
r124 19 53 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.655 $Y=0.905
+ $X2=0.655 $Y2=1.525
r125 15 54 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=0.57 $Y=2.555
+ $X2=0.57 $Y2=1.855
r126 4 45 300 $w=1.7e-07 $l=6.4591e-07 $layer=licon1_PDIFF $count=2 $X=3.495
+ $Y=1.885 $X2=4.055 $Y2=2.07
r127 3 43 600 $w=1.7e-07 $l=9.12318e-07 $layer=licon1_PDIFF $count=1 $X=1.465
+ $Y=2.055 $X2=1.605 $Y2=2.9
r128 3 26 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.465
+ $Y=2.055 $X2=1.605 $Y2=2.2
r129 2 49 182 $w=1.7e-07 $l=5.83095e-07 $layer=licon1_NDIFF $count=1 $X=4.03
+ $Y=0.625 $X2=4.405 $Y2=1.05
r130 1 29 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.425
+ $Y=0.585 $X2=1.565 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%A 1 3 6 8 15
c39 8 0 1.65079e-19 $X=1.2 $Y=1.295
c40 6 0 1.42935e-19 $X=1.39 $Y=2.555
r41 14 15 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.35 $Y=1.5 $X2=1.39
+ $Y2=1.5
r42 11 14 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.135 $Y=1.5
+ $X2=1.35 $Y2=1.5
r43 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.135
+ $Y=1.5 $X2=1.135 $Y2=1.5
r44 8 12 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.135 $Y=1.295
+ $X2=1.135 $Y2=1.5
r45 4 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.665
+ $X2=1.39 $Y2=1.5
r46 4 6 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=1.39 $Y=1.665 $X2=1.39
+ $Y2=2.555
r47 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.335
+ $X2=1.35 $Y2=1.5
r48 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.35 $Y=1.335 $X2=1.35
+ $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%A_474_313# 1 2 9 13 15 16 19 21 25 30 33 34
+ 37 44 45 46
c101 34 0 1.8437e-19 $X=4.06 $Y=0.7
c102 19 0 1.2352e-19 $X=3.42 $Y=2.305
r103 45 50 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=4.025 $Y=1.56
+ $X2=4.025 $Y2=1.655
r104 45 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.56
+ $X2=4.025 $Y2=1.395
r105 44 46 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.025 $Y=1.56
+ $X2=4.025 $Y2=1.395
r106 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.025
+ $Y=1.56 $X2=4.025 $Y2=1.56
r107 39 41 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=4.955 $Y=1.93
+ $X2=4.955 $Y2=2.9
r108 37 39 49.555 $w=2.48e-07 $l=1.075e-06 $layer=LI1_cond $X=4.955 $Y=0.855
+ $X2=4.955 $Y2=1.93
r109 35 37 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=4.955 $Y=0.785
+ $X2=4.955 $Y2=0.855
r110 33 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.83 $Y=0.7
+ $X2=4.955 $Y2=0.785
r111 33 34 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.83 $Y=0.7
+ $X2=4.06 $Y2=0.7
r112 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.975 $Y=0.785
+ $X2=4.06 $Y2=0.7
r113 31 46 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.975 $Y=0.785
+ $X2=3.975 $Y2=1.395
r114 27 29 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.445 $Y=1.64
+ $X2=2.595 $Y2=1.64
r115 25 49 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.955 $Y=0.945
+ $X2=3.955 $Y2=1.395
r116 22 30 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=3.495 $Y=1.655
+ $X2=3.42 $Y2=1.655
r117 21 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.86 $Y=1.655
+ $X2=4.025 $Y2=1.655
r118 21 22 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=3.86 $Y=1.655
+ $X2=3.495 $Y2=1.655
r119 17 30 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.42 $Y=1.745
+ $X2=3.42 $Y2=1.655
r120 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.42 $Y=1.745
+ $X2=3.42 $Y2=2.305
r121 16 29 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.67 $Y=1.64
+ $X2=2.595 $Y2=1.64
r122 15 30 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=3.345 $Y=1.64
+ $X2=3.42 $Y2=1.655
r123 15 16 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.345 $Y=1.64
+ $X2=2.67 $Y2=1.64
r124 11 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.595 $Y=1.565
+ $X2=2.595 $Y2=1.64
r125 11 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.595 $Y=1.565
+ $X2=2.595 $Y2=1.015
r126 7 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.445 $Y=1.715
+ $X2=2.445 $Y2=1.64
r127 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.445 $Y=1.715
+ $X2=2.445 $Y2=2.375
r128 2 41 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=4.85
+ $Y=1.785 $X2=4.995 $Y2=2.9
r129 2 39 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.85
+ $Y=1.785 $X2=4.995 $Y2=1.93
r130 1 37 182 $w=1.7e-07 $l=6.88694e-07 $layer=licon1_NDIFF $count=1 $X=4.85
+ $Y=0.235 $X2=4.995 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%B 3 7 9 10 11 12 15 17 21 23 26 28 31 33 36
+ 38 39 40 41 44 46
c121 46 0 2.0478e-20 $X=5.425 $Y=1.35
c122 26 0 4.68776e-20 $X=4.7 $Y=1.185
c123 21 0 4.21924e-20 $X=3.295 $Y=0.905
c124 7 0 1.76189e-20 $X=2.05 $Y=0.905
c125 3 0 9.95914e-20 $X=1.935 $Y=2.475
r126 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.425
+ $Y=1.35 $X2=5.425 $Y2=1.35
r127 43 46 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.21 $Y=1.35
+ $X2=5.425 $Y2=1.35
r128 43 44 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.21 $Y=1.35
+ $X2=5.135 $Y2=1.35
r129 41 47 3.26812 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=5.52 $Y=1.347
+ $X2=5.425 $Y2=1.347
r130 34 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.515
+ $X2=5.21 $Y2=1.35
r131 34 36 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=5.21 $Y=1.515
+ $X2=5.21 $Y2=2.415
r132 31 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.185
+ $X2=5.21 $Y2=1.35
r133 31 33 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.21 $Y=1.185
+ $X2=5.21 $Y2=0.655
r134 30 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.775 $Y=1.26
+ $X2=4.7 $Y2=1.26
r135 30 44 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.775 $Y=1.26
+ $X2=5.135 $Y2=1.26
r136 27 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.7 $Y=1.335
+ $X2=4.7 $Y2=1.26
r137 27 28 887.085 $w=1.5e-07 $l=1.73e-06 $layer=POLY_cond $X=4.7 $Y=1.335
+ $X2=4.7 $Y2=3.065
r138 26 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.7 $Y=1.185
+ $X2=4.7 $Y2=1.26
r139 25 26 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=4.7 $Y=0.255
+ $X2=4.7 $Y2=1.185
r140 24 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.37 $Y=0.18
+ $X2=3.295 $Y2=0.18
r141 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.625 $Y=0.18
+ $X2=4.7 $Y2=0.255
r142 23 24 643.521 $w=1.5e-07 $l=1.255e-06 $layer=POLY_cond $X=4.625 $Y=0.18
+ $X2=3.37 $Y2=0.18
r143 19 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.295 $Y=0.255
+ $X2=3.295 $Y2=0.18
r144 19 21 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.295 $Y=0.255
+ $X2=3.295 $Y2=0.905
r145 18 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.95 $Y=3.14
+ $X2=2.875 $Y2=3.14
r146 17 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.625 $Y=3.14
+ $X2=4.7 $Y2=3.065
r147 17 18 858.883 $w=1.5e-07 $l=1.675e-06 $layer=POLY_cond $X=4.625 $Y=3.14
+ $X2=2.95 $Y2=3.14
r148 13 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=3.065
+ $X2=2.875 $Y2=3.14
r149 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.875 $Y=3.065
+ $X2=2.875 $Y2=2.375
r150 11 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.22 $Y=0.18
+ $X2=3.295 $Y2=0.18
r151 11 12 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=3.22 $Y=0.18
+ $X2=2.125 $Y2=0.18
r152 9 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.8 $Y=3.14
+ $X2=2.875 $Y2=3.14
r153 9 10 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.8 $Y=3.14 $X2=2.01
+ $Y2=3.14
r154 5 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.05 $Y=0.255
+ $X2=2.125 $Y2=0.18
r155 5 7 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.05 $Y=0.255
+ $X2=2.05 $Y2=0.905
r156 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.935 $Y=3.065
+ $X2=2.01 $Y2=3.14
r157 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.935 $Y=3.065
+ $X2=1.935 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%A_1263_295# 1 2 9 13 15 16 19 22 23 25 28 33
+ 34 35
r73 34 35 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=8.15 $Y=2.245
+ $X2=8.15 $Y2=1.125
r74 33 34 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=8.065 $Y=2.41
+ $X2=8.065 $Y2=2.245
r75 26 35 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=8.19 $Y=1 $X2=8.19
+ $Y2=1.125
r76 26 28 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=8.19 $Y=1 $X2=8.19
+ $Y2=0.895
r77 24 33 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=8.065 $Y=2.415
+ $X2=8.065 $Y2=2.41
r78 24 25 16.2698 $w=3.38e-07 $l=4.8e-07 $layer=LI1_cond $X=8.065 $Y=2.415
+ $X2=8.065 $Y2=2.895
r79 22 25 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=7.895 $Y=2.98
+ $X2=8.065 $Y2=2.895
r80 22 23 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=7.895 $Y=2.98
+ $X2=6.645 $Y2=2.98
r81 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.48
+ $Y=1.64 $X2=6.48 $Y2=1.64
r82 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.48 $Y=2.895
+ $X2=6.645 $Y2=2.98
r83 17 19 43.8278 $w=3.28e-07 $l=1.255e-06 $layer=LI1_cond $X=6.48 $Y=2.895
+ $X2=6.48 $Y2=1.64
r84 15 20 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=6.665 $Y=1.64
+ $X2=6.48 $Y2=1.64
r85 15 16 5.03009 $w=3.3e-07 $l=9.2e-08 $layer=POLY_cond $X=6.665 $Y=1.64
+ $X2=6.757 $Y2=1.64
r86 11 16 37.0704 $w=1.5e-07 $l=1.73767e-07 $layer=POLY_cond $X=6.775 $Y=1.805
+ $X2=6.757 $Y2=1.64
r87 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.775 $Y=1.805
+ $X2=6.775 $Y2=2.385
r88 7 16 37.0704 $w=1.5e-07 $l=1.73292e-07 $layer=POLY_cond $X=6.74 $Y=1.475
+ $X2=6.757 $Y2=1.64
r89 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.74 $Y=1.475 $X2=6.74
+ $Y2=0.955
r90 2 33 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=7.835
+ $Y=1.915 $X2=7.98 $Y2=2.41
r91 1 28 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.005
+ $Y=0.685 $X2=8.15 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%C 1 3 6 8 9 12 16 19 21
r68 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.375
+ $Y=1.55 $X2=7.375 $Y2=1.55
r69 24 26 26.0127 $w=3.15e-07 $l=1.7e-07 $layer=POLY_cond $X=7.205 $Y=1.55
+ $X2=7.375 $Y2=1.55
r70 23 24 5.35556 $w=3.15e-07 $l=3.5e-08 $layer=POLY_cond $X=7.17 $Y=1.55
+ $X2=7.205 $Y2=1.55
r71 21 27 9.3293 $w=3.13e-07 $l=2.55e-07 $layer=LI1_cond $X=7.377 $Y=1.295
+ $X2=7.377 $Y2=1.55
r72 18 19 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=8.195 $Y=1.46
+ $X2=8.365 $Y2=1.46
r73 14 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.365 $Y=1.385
+ $X2=8.365 $Y2=1.46
r74 14 16 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=8.365 $Y=1.385
+ $X2=8.365 $Y2=0.895
r75 10 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.195 $Y=1.535
+ $X2=8.195 $Y2=1.46
r76 10 12 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=8.195 $Y=1.535
+ $X2=8.195 $Y2=2.235
r77 9 26 38.5363 $w=3.15e-07 $l=2.05122e-07 $layer=POLY_cond $X=7.54 $Y=1.46
+ $X2=7.375 $Y2=1.55
r78 8 18 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.12 $Y=1.46
+ $X2=8.195 $Y2=1.46
r79 8 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.12 $Y=1.46 $X2=7.54
+ $Y2=1.46
r80 4 24 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.205 $Y=1.715
+ $X2=7.205 $Y2=1.55
r81 4 6 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.205 $Y=1.715
+ $X2=7.205 $Y2=2.385
r82 1 23 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.17 $Y=1.385
+ $X2=7.17 $Y2=1.55
r83 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.17 $Y=1.385 $X2=7.17
+ $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%A_1363_127# 1 2 9 13 17 21 25 29 30 33 36 37
+ 42
r78 41 42 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.99 $Y=1.47 $X2=9.06
+ $Y2=1.47
r79 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r80 33 47 6.71605 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6.99 $Y=2.035
+ $X2=6.99 $Y2=1.92
r81 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=2.035
+ $X2=6.96 $Y2=2.035
r82 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=2.035
+ $X2=6.96 $Y2=2.035
r83 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=8.88 $Y2=2.035
r84 29 30 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=7.105 $Y2=2.035
r85 28 37 20.9535 $w=2.18e-07 $l=4e-07 $layer=LI1_cond $X=8.9 $Y=1.635 $X2=8.9
+ $Y2=2.035
r86 26 41 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=8.845 $Y=1.47
+ $X2=8.99 $Y2=1.47
r87 25 28 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.845 $Y=1.47
+ $X2=8.845 $Y2=1.635
r88 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.845
+ $Y=1.47 $X2=8.845 $Y2=1.47
r89 21 47 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.955 $Y=1.13
+ $X2=6.955 $Y2=1.92
r90 15 33 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=6.99 $Y=2.085 $X2=6.99
+ $Y2=2.035
r91 15 17 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.99 $Y=2.085
+ $X2=6.99 $Y2=2.11
r92 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.06 $Y=1.635
+ $X2=9.06 $Y2=1.47
r93 11 13 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=9.06 $Y=1.635
+ $X2=9.06 $Y2=2.465
r94 7 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.99 $Y=1.305
+ $X2=8.99 $Y2=1.47
r95 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.99 $Y=1.305 $X2=8.99
+ $Y2=0.685
r96 2 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.85
+ $Y=1.965 $X2=6.99 $Y2=2.11
r97 1 21 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=6.815
+ $Y=0.635 $X2=6.955 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%A_42_411# 1 2 3 4 17 19 22 23 24 27 29 33 34
+ 40 41 42 43
c83 27 0 1.2352e-19 $X=2.66 $Y=2.2
c84 23 0 9.95914e-20 $X=2.495 $Y=1.51
r85 40 41 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.2
+ $X2=0.265 $Y2=2.035
r86 38 41 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.175 $Y=1.245
+ $X2=0.175 $Y2=2.035
r87 37 38 17.7387 $w=5.13e-07 $l=5.15e-07 $layer=LI1_cond $X=0.347 $Y=0.73
+ $X2=0.347 $Y2=1.245
r88 34 37 1.85799 $w=5.13e-07 $l=8e-08 $layer=LI1_cond $X=0.347 $Y=0.65
+ $X2=0.347 $Y2=0.73
r89 33 42 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.74 $Y=1.425
+ $X2=2.66 $Y2=1.51
r90 33 43 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.74 $Y=1.425
+ $X2=2.74 $Y2=1.245
r91 29 43 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=2.832 $Y=1.068
+ $X2=2.832 $Y2=1.245
r92 29 31 4.74254 $w=3.55e-07 $l=1.38e-07 $layer=LI1_cond $X=2.832 $Y=1.068
+ $X2=2.832 $Y2=0.93
r93 25 42 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=1.595
+ $X2=2.66 $Y2=1.51
r94 25 27 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=2.66 $Y=1.595
+ $X2=2.66 $Y2=2.2
r95 23 42 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=1.51
+ $X2=2.66 $Y2=1.51
r96 23 24 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.495 $Y=1.51 $X2=2
+ $Y2=1.51
r97 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.915 $Y=1.425
+ $X2=2 $Y2=1.51
r98 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.915 $Y=0.735
+ $X2=1.915 $Y2=1.425
r99 20 34 7.34265 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=0.605 $Y=0.65
+ $X2=0.347 $Y2=0.65
r100 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.83 $Y=0.65
+ $X2=1.915 $Y2=0.735
r101 19 20 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=1.83 $Y=0.65
+ $X2=0.605 $Y2=0.65
r102 15 40 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.265 $Y=2.21
+ $X2=0.265 $Y2=2.2
r103 15 17 22.7196 $w=3.48e-07 $l=6.9e-07 $layer=LI1_cond $X=0.265 $Y=2.21
+ $X2=0.265 $Y2=2.9
r104 4 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.52
+ $Y=2.055 $X2=2.66 $Y2=2.2
r105 3 40 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=2.055 $X2=0.355 $Y2=2.2
r106 3 17 400 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=2.055 $X2=0.355 $Y2=2.9
r107 2 31 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=2.67
+ $Y=0.805 $X2=2.925 $Y2=0.93
r108 1 37 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.295
+ $Y=0.585 $X2=0.44 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%VPWR 1 2 3 12 16 22 27 28 29 31 36 49 50 53
+ 56
r74 56 57 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r77 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r78 47 57 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=5.52 $Y2=3.33
r79 46 47 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r80 44 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=3.33
+ $X2=5.425 $Y2=3.33
r81 44 46 183.326 $w=1.68e-07 $l=2.81e-06 $layer=LI1_cond $X=5.59 $Y=3.33
+ $X2=8.4 $Y2=3.33
r82 43 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r83 42 43 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 39 42 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 39 40 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r87 37 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.785 $Y2=3.33
r88 37 39 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=3.33 $X2=1.2
+ $Y2=3.33
r89 36 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=3.33
+ $X2=5.425 $Y2=3.33
r90 36 42 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=3.33
+ $X2=5.04 $Y2=3.33
r91 34 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r92 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r93 31 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.785 $Y2=3.33
r94 31 33 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.24 $Y2=3.33
r95 29 43 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.04 $Y2=3.33
r96 29 40 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=4.8 $Y=3.33 $X2=1.2
+ $Y2=3.33
r97 27 46 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=8.44 $Y=3.33 $X2=8.4
+ $Y2=3.33
r98 27 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=3.33
+ $X2=8.525 $Y2=3.33
r99 26 49 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.61 $Y=3.33
+ $X2=9.36 $Y2=3.33
r100 26 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.61 $Y=3.33
+ $X2=8.525 $Y2=3.33
r101 22 25 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=8.525 $Y=1.98
+ $X2=8.525 $Y2=2.95
r102 20 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=3.245
+ $X2=8.525 $Y2=3.33
r103 20 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.525 $Y=3.245
+ $X2=8.525 $Y2=2.95
r104 16 19 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=5.425 $Y=1.93
+ $X2=5.425 $Y2=2.9
r105 14 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=3.245
+ $X2=5.425 $Y2=3.33
r106 14 19 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=5.425 $Y=3.245
+ $X2=5.425 $Y2=2.9
r107 10 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r108 10 12 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.36
r109 3 25 400 $w=1.7e-07 $l=1.15549e-06 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=1.915 $X2=8.525 $Y2=2.95
r110 3 22 400 $w=1.7e-07 $l=2.85657e-07 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=1.915 $X2=8.525 $Y2=1.98
r111 2 19 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.785 $X2=5.425 $Y2=2.9
r112 2 16 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.785 $X2=5.425 $Y2=1.93
r113 1 12 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=0.645
+ $Y=2.055 $X2=0.785 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%A_402_411# 1 2 3 4 15 17 18 22 23 24 26 27 28
+ 30 31 32 35 41 42
c129 28 0 4.68776e-20 $X=5.43 $Y=0.86
c130 15 0 1.60554e-19 $X=2.15 $Y=2.2
r131 41 42 8.72283 $w=3.78e-07 $l=1.7e-07 $layer=LI1_cond $X=7.61 $Y=1.895
+ $X2=7.61 $Y2=2.065
r132 37 41 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=7.8 $Y=0.435
+ $X2=7.8 $Y2=1.895
r133 35 42 1.36474 $w=3.78e-07 $l=4.5e-08 $layer=LI1_cond $X=7.525 $Y=2.11
+ $X2=7.525 $Y2=2.065
r134 31 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.715 $Y=0.35
+ $X2=7.8 $Y2=0.435
r135 31 32 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=7.715 $Y=0.35
+ $X2=6.34 $Y2=0.35
r136 30 40 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.215 $Y=0.775
+ $X2=6.215 $Y2=0.86
r137 29 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.215 $Y=0.435
+ $X2=6.34 $Y2=0.35
r138 29 30 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=6.215 $Y=0.435
+ $X2=6.215 $Y2=0.775
r139 27 40 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.09 $Y=0.86
+ $X2=6.215 $Y2=0.86
r140 27 28 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.09 $Y=0.86
+ $X2=5.43 $Y2=0.86
r141 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.345 $Y=0.775
+ $X2=5.43 $Y2=0.86
r142 25 26 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.345 $Y=0.435
+ $X2=5.345 $Y2=0.775
r143 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.26 $Y=0.35
+ $X2=5.345 $Y2=0.435
r144 23 24 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=5.26 $Y=0.35
+ $X2=3.71 $Y2=0.35
r145 20 22 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=3.625 $Y=2.545
+ $X2=3.625 $Y2=0.73
r146 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=0.435
+ $X2=3.71 $Y2=0.35
r147 19 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.625 $Y=0.435
+ $X2=3.625 $Y2=0.73
r148 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.54 $Y=2.63
+ $X2=3.625 $Y2=2.545
r149 17 18 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=3.54 $Y=2.63
+ $X2=2.315 $Y2=2.63
r150 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.15 $Y=2.545
+ $X2=2.315 $Y2=2.63
r151 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.15 $Y=2.545
+ $X2=2.15 $Y2=2.2
r152 4 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.28
+ $Y=1.965 $X2=7.42 $Y2=2.11
r153 3 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.01
+ $Y=2.055 $X2=2.15 $Y2=2.2
r154 2 40 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.11
+ $Y=0.635 $X2=6.255 $Y2=0.78
r155 1 22 91 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=2 $X=3.37
+ $Y=0.585 $X2=3.625 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%A_425_117# 1 2 3 4 15 19 20 23 24 26 27 28 30
+ 35 36 39 42 43 49
c114 35 0 6.26704e-20 $X=5.855 $Y=2.035
r115 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=2.035 $X2=6
+ $Y2=2.035
r116 39 49 8.66137 $w=3.53e-07 $l=1.7e-07 $layer=LI1_cond $X=3.182 $Y=2.035
+ $X2=3.182 $Y2=1.865
r117 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=2.035
+ $X2=3.12 $Y2=2.035
r118 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=2.035
+ $X2=3.12 $Y2=2.035
r119 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.855 $Y=2.035
+ $X2=6 $Y2=2.035
r120 35 36 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=5.855 $Y=2.035
+ $X2=3.265 $Y2=2.035
r121 30 33 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=7.345 $Y=0.7
+ $X2=7.345 $Y2=0.805
r122 29 43 34.1123 $w=2.48e-07 $l=7.4e-07 $layer=LI1_cond $X=6.01 $Y=1.295
+ $X2=6.01 $Y2=2.035
r123 27 30 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.22 $Y=0.7
+ $X2=7.345 $Y2=0.7
r124 27 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.22 $Y=0.7
+ $X2=6.69 $Y2=0.7
r125 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.605 $Y=0.785
+ $X2=6.69 $Y2=0.7
r126 25 26 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.605 $Y=0.785
+ $X2=6.605 $Y2=1.125
r127 24 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.135 $Y=1.21
+ $X2=6.01 $Y2=1.295
r128 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.52 $Y=1.21
+ $X2=6.605 $Y2=1.125
r129 23 24 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.52 $Y=1.21
+ $X2=6.135 $Y2=1.21
r130 21 49 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=3.275 $Y=0.435
+ $X2=3.275 $Y2=1.865
r131 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.19 $Y=0.35
+ $X2=3.275 $Y2=0.435
r132 19 20 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.19 $Y=0.35
+ $X2=2.43 $Y2=0.35
r133 15 17 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=2.305 $Y=0.73
+ $X2=2.305 $Y2=1.08
r134 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.305 $Y=0.435
+ $X2=2.43 $Y2=0.35
r135 13 15 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.305 $Y=0.435
+ $X2=2.305 $Y2=0.73
r136 4 43 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.905
+ $Y=1.965 $X2=6.05 $Y2=2.11
r137 3 39 600 $w=1.7e-07 $l=2.83417e-07 $layer=licon1_PDIFF $count=1 $X=2.95
+ $Y=2.055 $X2=3.205 $Y2=2.115
r138 2 33 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=7.245
+ $Y=0.635 $X2=7.385 $Y2=0.805
r139 1 17 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=2.125
+ $Y=0.585 $X2=2.265 $Y2=1.08
r140 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.125
+ $Y=0.585 $X2=2.265 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%X 1 2 7 8 9 10 11 12 13 24 45
r17 22 45 0.45038 $w=4.33e-07 $l=1.7e-08 $layer=LI1_cond $X=9.257 $Y=0.908
+ $X2=9.257 $Y2=0.925
r18 13 42 5.05457 $w=2.83e-07 $l=1.25e-07 $layer=LI1_cond $X=9.332 $Y=2.775
+ $X2=9.332 $Y2=2.9
r19 12 13 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=9.332 $Y=2.405
+ $X2=9.332 $Y2=2.775
r20 11 12 17.1856 $w=2.83e-07 $l=4.25e-07 $layer=LI1_cond $X=9.332 $Y=1.98
+ $X2=9.332 $Y2=2.405
r21 10 11 12.7375 $w=2.83e-07 $l=3.15e-07 $layer=LI1_cond $X=9.332 $Y=1.665
+ $X2=9.332 $Y2=1.98
r22 9 10 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=9.332 $Y=1.295
+ $X2=9.332 $Y2=1.665
r23 9 47 6.87422 $w=2.83e-07 $l=1.7e-07 $layer=LI1_cond $X=9.332 $Y=1.295
+ $X2=9.332 $Y2=1.125
r24 8 47 5.7677 $w=4.33e-07 $l=1.66e-07 $layer=LI1_cond $X=9.257 $Y=0.959
+ $X2=9.257 $Y2=1.125
r25 8 45 0.90076 $w=4.33e-07 $l=3.4e-08 $layer=LI1_cond $X=9.257 $Y=0.959
+ $X2=9.257 $Y2=0.925
r26 8 22 0.90076 $w=4.33e-07 $l=3.4e-08 $layer=LI1_cond $X=9.257 $Y=0.874
+ $X2=9.257 $Y2=0.908
r27 7 8 8.45125 $w=4.33e-07 $l=3.19e-07 $layer=LI1_cond $X=9.257 $Y=0.555
+ $X2=9.257 $Y2=0.874
r28 7 24 3.31162 $w=4.33e-07 $l=1.25e-07 $layer=LI1_cond $X=9.257 $Y=0.555
+ $X2=9.257 $Y2=0.43
r29 2 42 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=9.135
+ $Y=1.835 $X2=9.275 $Y2=2.9
r30 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.135
+ $Y=1.835 $X2=9.275 $Y2=1.98
r31 1 24 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=9.065
+ $Y=0.265 $X2=9.205 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_1%VGND 1 2 3 12 16 20 21 28 29 31 32 33 52 53
r69 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r70 50 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r71 49 50 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r72 47 50 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6 $Y=0 $X2=8.4
+ $Y2=0
r73 46 49 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.4 $Y2=0
r74 46 47 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r75 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r76 43 44 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r77 40 43 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.52
+ $Y2=0
r78 40 41 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r79 37 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r80 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r81 33 44 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.52
+ $Y2=0
r82 33 41 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=1.2
+ $Y2=0
r83 31 49 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=8.53 $Y=0 $X2=8.4
+ $Y2=0
r84 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.53 $Y=0 $X2=8.695
+ $Y2=0
r85 30 52 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=8.86 $Y=0 $X2=9.36
+ $Y2=0
r86 30 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.86 $Y=0 $X2=8.695
+ $Y2=0
r87 28 43 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.52
+ $Y2=0
r88 28 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.61 $Y=0 $X2=5.735
+ $Y2=0
r89 27 46 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.86 $Y=0 $X2=6
+ $Y2=0
r90 27 29 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.86 $Y=0 $X2=5.735
+ $Y2=0
r91 23 40 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.2
+ $Y2=0
r92 21 36 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.72
+ $Y2=0
r93 20 25 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.95
+ $Y2=0.3
r94 20 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.115
+ $Y2=0
r95 20 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r96 16 18 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=8.695 $Y=0.41
+ $X2=8.695 $Y2=0.96
r97 14 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.695 $Y=0.085
+ $X2=8.695 $Y2=0
r98 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.695 $Y=0.085
+ $X2=8.695 $Y2=0.41
r99 10 29 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0.085
+ $X2=5.735 $Y2=0
r100 10 12 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=5.735 $Y=0.085
+ $X2=5.735 $Y2=0.405
r101 3 18 182 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_NDIFF $count=1 $X=8.44
+ $Y=0.685 $X2=8.695 $Y2=0.96
r102 3 16 182 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_NDIFF $count=1 $X=8.44
+ $Y=0.685 $X2=8.695 $Y2=0.41
r103 2 12 182 $w=1.7e-07 $l=4.87647e-07 $layer=licon1_NDIFF $count=1 $X=5.285
+ $Y=0.235 $X2=5.695 $Y2=0.405
r104 1 25 182 $w=1.7e-07 $l=3.79374e-07 $layer=licon1_NDIFF $count=1 $X=0.73
+ $Y=0.585 $X2=0.95 $Y2=0.3
.ends

