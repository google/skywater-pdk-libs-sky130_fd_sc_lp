* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4_lp A B C D VGND VNB VPB VPWR X
M1000 VGND A a_646_167# VNB nshort w=420000u l=150000u
+  ad=3.549e+11p pd=4.21e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_154_419# D a_27_47# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=2.85e+11p ps=2.57e+06u
M1002 a_804_167# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1003 a_646_167# A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.906e+11p ps=4.38e+06u
M1004 a_114_47# D a_27_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 a_272_47# C VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1006 a_27_47# C a_272_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_366_419# B a_252_419# VPB phighvt w=1e+06u l=250000u
+  ad=1.21e+12p pd=4.42e+06u as=3.2e+11p ps=2.64e+06u
M1008 X a_27_47# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=5.65e+11p ps=3.13e+06u
M1009 a_252_419# C a_154_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_47# B a_465_185# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.5225e+11p ps=1.67e+06u
M1011 a_465_185# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_366_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_27_47# a_804_167# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1014 VGND D a_114_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
