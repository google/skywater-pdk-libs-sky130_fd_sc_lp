* File: sky130_fd_sc_lp__clkinvlp_16.spice
* Created: Wed Sep  2 09:41:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkinvlp_16.pex.spice"
.subckt sky130_fd_sc_lp__clkinvlp_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_A_M1025_g A_268_67# VNB NSHORT L=0.15 W=0.55 AD=0.14575
+ AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.2
+ SB=75007.7 A=0.0825 P=1.4 MULT=1
MM1001 A_268_67# N_A_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.5 SB=75007.3
+ A=0.0825 P=1.4 MULT=1
MM1005 A_426_67# N_A_M1005_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75001 SB=75006.9
+ A=0.0825 P=1.4 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g A_426_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001.3
+ SB=75006.5 A=0.0825 P=1.4 MULT=1
MM1010 N_VGND_M1004_d N_A_M1010_g A_1058_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001.8
+ SB=75006.1 A=0.0825 P=1.4 MULT=1
MM1006 A_1058_67# N_A_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75002.1 SB=75005.7
+ A=0.0825 P=1.4 MULT=1
MM1008 A_1532_67# N_A_M1008_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75002.6 SB=75005.3
+ A=0.0825 P=1.4 MULT=1
MM1031 N_VGND_M1031_d N_A_M1031_g A_1532_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75002.9
+ SB=75004.9 A=0.0825 P=1.4 MULT=1
MM1015 N_VGND_M1031_d N_A_M1015_g A_1216_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75003.3
+ SB=75004.5 A=0.0825 P=1.4 MULT=1
MM1013 A_1216_67# N_A_M1013_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75003.7 SB=75004.1
+ A=0.0825 P=1.4 MULT=1
MM1014 A_110_67# N_A_M1014_g N_Y_M1013_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75004.1 SB=75003.7
+ A=0.0825 P=1.4 MULT=1
MM1024 N_VGND_M1024_d N_A_M1024_g A_110_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75004.5
+ SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1019 N_VGND_M1024_d N_A_M1019_g A_584_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75004.9
+ SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1018 A_584_67# N_A_M1018_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75005.3 SB=75002.6
+ A=0.0825 P=1.4 MULT=1
MM1020 A_742_67# N_A_M1020_g N_Y_M1018_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75005.7 SB=75002.1
+ A=0.0825 P=1.4 MULT=1
MM1027 N_VGND_M1027_d N_A_M1027_g A_742_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75006.1
+ SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1026 N_VGND_M1027_d N_A_M1026_g A_1374_67# VNB NSHORT L=0.15 W=0.55 AD=0.077
+ AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75006.5
+ SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1028 A_1374_67# N_A_M1028_g N_Y_M1028_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75006.9 SB=75001
+ A=0.0825 P=1.4 MULT=1
MM1032 A_900_67# N_A_M1032_g N_Y_M1028_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75007.3 SB=75000.5
+ A=0.0825 P=1.4 MULT=1
MM1033 N_VGND_M1033_d N_A_M1033_g A_900_67# VNB NSHORT L=0.15 W=0.55 AD=0.14575
+ AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75007.7
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125008 A=0.25 P=2.5
+ MULT=1
MM1002 N_Y_M1000_d N_A_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125008 A=0.25 P=2.5
+ MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VPWR_M1002_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125007 A=0.25 P=2.5
+ MULT=1
MM1007 N_Y_M1003_d N_A_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125006 A=0.25 P=2.5
+ MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VPWR_M1007_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125006 A=0.25 P=2.5
+ MULT=1
MM1011 N_Y_M1009_d N_A_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125005 A=0.25 P=2.5
+ MULT=1
MM1012 N_Y_M1012_d N_A_M1012_g N_VPWR_M1011_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125005 A=0.25 P=2.5
+ MULT=1
MM1016 N_Y_M1012_d N_A_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125004 A=0.25 P=2.5
+ MULT=1
MM1017 N_Y_M1017_d N_A_M1017_g N_VPWR_M1016_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125004 A=0.25 P=2.5
+ MULT=1
MM1021 N_Y_M1017_d N_A_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125005 SB=125003 A=0.25 P=2.5
+ MULT=1
MM1022 N_Y_M1022_d N_A_M1022_g N_VPWR_M1021_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125005 SB=125003 A=0.25 P=2.5
+ MULT=1
MM1023 N_Y_M1022_d N_A_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125006 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1029 N_Y_M1029_d N_A_M1029_g N_VPWR_M1023_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125006 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1030 N_Y_M1029_d N_A_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125007 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1034 N_Y_M1034_d N_A_M1034_g N_VPWR_M1030_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125008 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1035 N_Y_M1034_d N_A_M1035_g N_VPWR_M1035_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 M=1 R=4 SA=125008 SB=125000 A=0.25 P=2.5
+ MULT=1
DX36_noxref VNB VPB NWDIODE A=17.7175 P=22.73
*
.include "sky130_fd_sc_lp__clkinvlp_16.pxi.spice"
*
.ends
*
*
