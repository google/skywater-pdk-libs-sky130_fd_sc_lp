* File: sky130_fd_sc_lp__o2bb2a_2.pxi.spice
* Created: Wed Sep  2 10:21:28 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2A_2%B1 N_B1_M1004_g N_B1_M1001_g N_B1_c_91_n
+ N_B1_c_92_n B1 N_B1_c_94_n PM_SKY130_FD_SC_LP__O2BB2A_2%B1
x_PM_SKY130_FD_SC_LP__O2BB2A_2%B2 N_B2_M1010_g N_B2_M1003_g N_B2_c_120_n
+ N_B2_c_121_n B2 N_B2_c_123_n PM_SKY130_FD_SC_LP__O2BB2A_2%B2
x_PM_SKY130_FD_SC_LP__O2BB2A_2%A_300_21# N_A_300_21#_M1011_s N_A_300_21#_M1000_d
+ N_A_300_21#_M1009_g N_A_300_21#_M1007_g N_A_300_21#_c_158_n
+ N_A_300_21#_c_159_n N_A_300_21#_c_160_n N_A_300_21#_c_161_n
+ N_A_300_21#_c_162_n N_A_300_21#_c_163_n PM_SKY130_FD_SC_LP__O2BB2A_2%A_300_21#
x_PM_SKY130_FD_SC_LP__O2BB2A_2%A2_N N_A2_N_M1000_g N_A2_N_c_227_n N_A2_N_M1011_g
+ N_A2_N_c_228_n N_A2_N_c_229_n A2_N A2_N PM_SKY130_FD_SC_LP__O2BB2A_2%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2A_2%A1_N N_A1_N_M1008_g N_A1_N_M1012_g A1_N A1_N A1_N
+ N_A1_N_c_273_n PM_SKY130_FD_SC_LP__O2BB2A_2%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2A_2%A_222_367# N_A_222_367#_M1009_d
+ N_A_222_367#_M1010_d N_A_222_367#_c_313_n N_A_222_367#_M1002_g
+ N_A_222_367#_M1005_g N_A_222_367#_c_315_n N_A_222_367#_M1006_g
+ N_A_222_367#_M1013_g N_A_222_367#_c_324_n N_A_222_367#_c_317_n
+ N_A_222_367#_c_326_n N_A_222_367#_c_318_n N_A_222_367#_c_319_n
+ N_A_222_367#_c_327_n N_A_222_367#_c_328_n N_A_222_367#_c_329_n
+ N_A_222_367#_c_330_n N_A_222_367#_c_331_n N_A_222_367#_c_332_n
+ N_A_222_367#_c_320_n N_A_222_367#_c_334_n N_A_222_367#_c_321_n
+ PM_SKY130_FD_SC_LP__O2BB2A_2%A_222_367#
x_PM_SKY130_FD_SC_LP__O2BB2A_2%VPWR N_VPWR_M1001_s N_VPWR_M1007_d N_VPWR_M1008_d
+ N_VPWR_M1013_d N_VPWR_c_441_n N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n
+ N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n N_VPWR_c_449_n
+ VPWR N_VPWR_c_450_n N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_440_n
+ PM_SKY130_FD_SC_LP__O2BB2A_2%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2A_2%X N_X_M1002_d N_X_M1005_s X X X X X X X
+ N_X_c_498_n PM_SKY130_FD_SC_LP__O2BB2A_2%X
x_PM_SKY130_FD_SC_LP__O2BB2A_2%A_67_47# N_A_67_47#_M1004_s N_A_67_47#_M1003_d
+ N_A_67_47#_c_515_n N_A_67_47#_c_516_n N_A_67_47#_c_517_n N_A_67_47#_c_533_p
+ PM_SKY130_FD_SC_LP__O2BB2A_2%A_67_47#
x_PM_SKY130_FD_SC_LP__O2BB2A_2%VGND N_VGND_M1004_d N_VGND_M1012_d N_VGND_M1006_s
+ N_VGND_c_539_n N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n N_VGND_c_543_n
+ N_VGND_c_544_n VGND N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n
+ N_VGND_c_548_n PM_SKY130_FD_SC_LP__O2BB2A_2%VGND
cc_1 VNB N_B1_M1004_g 0.0375506f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.445
cc_2 VNB N_B1_c_91_n 0.0249397f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.5
cc_3 VNB N_B1_c_92_n 0.0114369f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.665
cc_4 VNB B1 0.030001f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_B1_c_94_n 0.0168101f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.16
cc_6 VNB N_B2_M1003_g 0.0276322f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.155
cc_7 VNB N_B2_c_120_n 0.0208296f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.5
cc_8 VNB N_B2_c_121_n 0.0095707f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.665
cc_9 VNB B2 0.00409202f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_B2_c_123_n 0.0148583f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.16
cc_11 VNB N_A_300_21#_M1009_g 0.0532367f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.16
cc_12 VNB N_A_300_21#_c_158_n 0.00834365f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.16
cc_13 VNB N_A_300_21#_c_159_n 0.00587424f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.16
cc_14 VNB N_A_300_21#_c_160_n 0.0372922f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.33
cc_15 VNB N_A_300_21#_c_161_n 0.0161608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_300_21#_c_162_n 0.00137076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_300_21#_c_163_n 0.00359215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_N_M1000_g 0.0295232f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.445
cc_19 VNB N_A2_N_c_227_n 0.0195565f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.665
cc_20 VNB N_A2_N_c_228_n 0.0471324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_N_c_229_n 0.0343663f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.16
cc_22 VNB A2_N 0.0121392f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.5
cc_23 VNB N_A1_N_M1008_g 0.00899951f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.445
cc_24 VNB N_A1_N_M1012_g 0.0402948f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.155
cc_25 VNB A1_N 0.00499604f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.16
cc_26 VNB N_A1_N_c_273_n 0.0403041f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.33
cc_27 VNB N_A_222_367#_c_313_n 0.0174094f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.155
cc_28 VNB N_A_222_367#_M1005_g 0.00782487f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.665
cc_29 VNB N_A_222_367#_c_315_n 0.0210923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_222_367#_M1013_g 0.0106048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_222_367#_c_317_n 0.00304537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_222_367#_c_318_n 0.00636643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_222_367#_c_319_n 0.00715909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_222_367#_c_320_n 0.003711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_222_367#_c_321_n 0.0705678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_440_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_498_n 0.00186095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_67_47#_c_515_n 0.0144956f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.16
cc_39 VNB N_A_67_47#_c_516_n 0.018162f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.5
cc_40 VNB N_A_67_47#_c_517_n 0.0135259f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.665
cc_41 VNB N_VGND_c_539_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.665
cc_42 VNB N_VGND_c_540_n 0.00635104f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.16
cc_43 VNB N_VGND_c_541_n 0.0132265f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.33
cc_44 VNB N_VGND_c_542_n 0.0468913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_543_n 0.0215789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_544_n 0.00436274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_545_n 0.0614829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_546_n 0.0156522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_547_n 0.00532666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_548_n 0.27183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_B1_M1001_g 0.0264754f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.155
cc_52 VPB N_B1_c_92_n 0.0053729f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.665
cc_53 VPB B1 0.00405683f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_54 VPB N_B2_M1010_g 0.0219278f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.445
cc_55 VPB N_B2_c_121_n 0.00615906f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.665
cc_56 VPB N_A_300_21#_M1007_g 0.0253973f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_57 VPB N_A_300_21#_c_158_n 2.50584e-19 $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.16
cc_58 VPB N_A_300_21#_c_160_n 0.0121555f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.33
cc_59 VPB N_A_300_21#_c_162_n 0.00504408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A2_N_M1000_g 0.0249785f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.445
cc_61 VPB N_A1_N_M1008_g 0.0219638f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.445
cc_62 VPB N_A_222_367#_M1005_g 0.0225271f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.665
cc_63 VPB N_A_222_367#_M1013_g 0.0265092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_222_367#_c_324_n 0.00811869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_222_367#_c_317_n 0.0010595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_222_367#_c_326_n 0.00703609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_222_367#_c_327_n 0.00232732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_222_367#_c_328_n 0.0181513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_222_367#_c_329_n 0.00375904f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_222_367#_c_330_n 0.00214544f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_222_367#_c_331_n 0.00783938f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_222_367#_c_332_n 8.88701e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_222_367#_c_320_n 3.34066e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_222_367#_c_334_n 0.00791998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_441_n 0.0822738f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.16
cc_76 VPB N_VPWR_c_442_n 0.0447718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_443_n 0.0173732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_444_n 0.0132006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_445_n 0.0626262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_446_n 0.0115308f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_447_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_448_n 0.0381228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_449_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_450_n 0.0335824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_451_n 0.0156522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_452_n 0.00587781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_440_n 0.10815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_X_c_498_n 0.00127418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 N_B1_M1001_g N_B2_M1010_g 0.0242591f $X=0.675 $Y=2.155 $X2=0 $Y2=0
cc_90 N_B1_M1004_g N_B2_M1003_g 0.0218185f $X=0.675 $Y=0.445 $X2=0 $Y2=0
cc_91 N_B1_c_91_n N_B2_c_120_n 0.0242591f $X=0.585 $Y=1.5 $X2=0 $Y2=0
cc_92 N_B1_c_92_n N_B2_c_121_n 0.0242591f $X=0.585 $Y=1.665 $X2=0 $Y2=0
cc_93 B1 B2 0.0537867f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B1_c_94_n B2 6.4208e-19 $X=0.585 $Y=1.16 $X2=0 $Y2=0
cc_95 B1 N_B2_c_123_n 0.00425212f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_96 N_B1_c_94_n N_B2_c_123_n 0.0242591f $X=0.585 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B1_M1001_g N_VPWR_c_441_n 0.0165606f $X=0.675 $Y=2.155 $X2=0 $Y2=0
cc_98 N_B1_c_92_n N_VPWR_c_441_n 0.00465857f $X=0.585 $Y=1.665 $X2=0 $Y2=0
cc_99 B1 N_VPWR_c_441_n 0.0150592f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B1_M1001_g N_VPWR_c_448_n 0.00259749f $X=0.675 $Y=2.155 $X2=0 $Y2=0
cc_101 N_B1_M1001_g N_VPWR_c_440_n 0.00344639f $X=0.675 $Y=2.155 $X2=0 $Y2=0
cc_102 N_B1_M1004_g N_A_67_47#_c_516_n 0.0133491f $X=0.675 $Y=0.445 $X2=0 $Y2=0
cc_103 B1 N_A_67_47#_c_516_n 0.0208624f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B1_c_94_n N_A_67_47#_c_516_n 6.46979e-19 $X=0.585 $Y=1.16 $X2=0 $Y2=0
cc_105 B1 N_A_67_47#_c_517_n 0.0135046f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B1_c_94_n N_A_67_47#_c_517_n 0.00413223f $X=0.585 $Y=1.16 $X2=0 $Y2=0
cc_107 N_B1_M1004_g N_VGND_c_539_n 0.00783675f $X=0.675 $Y=0.445 $X2=0 $Y2=0
cc_108 N_B1_M1004_g N_VGND_c_543_n 0.00413026f $X=0.675 $Y=0.445 $X2=0 $Y2=0
cc_109 N_B1_M1004_g N_VGND_c_548_n 0.00597133f $X=0.675 $Y=0.445 $X2=0 $Y2=0
cc_110 N_B2_M1003_g N_A_300_21#_M1009_g 0.0223674f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_111 B2 N_A_300_21#_M1009_g 0.00196327f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B2_c_123_n N_A_300_21#_M1009_g 0.0216864f $X=1.125 $Y=1.16 $X2=0 $Y2=0
cc_113 N_B2_M1010_g N_A_300_21#_M1007_g 0.00891457f $X=1.035 $Y=2.155 $X2=0
+ $Y2=0
cc_114 N_B2_c_120_n N_A_300_21#_c_158_n 0.0216864f $X=1.125 $Y=1.5 $X2=0 $Y2=0
cc_115 N_B2_M1010_g N_A_222_367#_c_324_n 6.17434e-19 $X=1.035 $Y=2.155 $X2=0
+ $Y2=0
cc_116 N_B2_M1010_g N_A_222_367#_c_317_n 0.00156713f $X=1.035 $Y=2.155 $X2=0
+ $Y2=0
cc_117 N_B2_c_120_n N_A_222_367#_c_317_n 0.00145353f $X=1.125 $Y=1.5 $X2=0 $Y2=0
cc_118 B2 N_A_222_367#_c_317_n 0.0394426f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_119 B2 N_A_222_367#_c_318_n 0.0142472f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B2_c_123_n N_A_222_367#_c_318_n 5.69795e-19 $X=1.125 $Y=1.16 $X2=0
+ $Y2=0
cc_121 N_B2_M1010_g N_A_222_367#_c_334_n 0.00182441f $X=1.035 $Y=2.155 $X2=0
+ $Y2=0
cc_122 N_B2_c_121_n N_A_222_367#_c_334_n 0.00397127f $X=1.125 $Y=1.665 $X2=0
+ $Y2=0
cc_123 B2 N_A_222_367#_c_334_n 0.0122788f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_124 N_B2_M1010_g N_VPWR_c_441_n 0.00235915f $X=1.035 $Y=2.155 $X2=0 $Y2=0
cc_125 N_B2_M1010_g N_VPWR_c_448_n 0.00312414f $X=1.035 $Y=2.155 $X2=0 $Y2=0
cc_126 N_B2_M1010_g N_VPWR_c_440_n 0.00410284f $X=1.035 $Y=2.155 $X2=0 $Y2=0
cc_127 N_B2_M1003_g N_A_67_47#_c_516_n 0.0116186f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_128 B2 N_A_67_47#_c_516_n 0.0224506f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B2_c_123_n N_A_67_47#_c_516_n 0.00550373f $X=1.125 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B2_M1003_g N_VGND_c_539_n 0.00685255f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_131 N_B2_M1003_g N_VGND_c_545_n 0.00413026f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_132 N_B2_M1003_g N_VGND_c_548_n 0.00484119f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_133 N_A_300_21#_c_160_n N_A2_N_M1000_g 0.0123987f $X=1.98 $Y=1.5 $X2=0 $Y2=0
cc_134 N_A_300_21#_c_161_n N_A2_N_M1000_g 0.00921333f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_135 N_A_300_21#_c_162_n N_A2_N_M1000_g 0.00488559f $X=2.77 $Y=1.98 $X2=0
+ $Y2=0
cc_136 N_A_300_21#_c_163_n N_A2_N_M1000_g 0.0163935f $X=2.662 $Y=1.46 $X2=0
+ $Y2=0
cc_137 N_A_300_21#_c_161_n N_A2_N_c_227_n 0.0112986f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_138 N_A_300_21#_M1009_g N_A2_N_c_228_n 0.00840288f $X=1.575 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A_300_21#_c_159_n N_A2_N_c_228_n 0.00752705f $X=2.47 $Y=1.46 $X2=0
+ $Y2=0
cc_140 N_A_300_21#_c_160_n N_A2_N_c_228_n 0.00574503f $X=1.98 $Y=1.5 $X2=0 $Y2=0
cc_141 N_A_300_21#_c_161_n N_A2_N_c_228_n 0.00527364f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_142 N_A_300_21#_c_161_n N_A2_N_c_229_n 0.0232289f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_143 N_A_300_21#_c_159_n A2_N 0.0144488f $X=2.47 $Y=1.46 $X2=0 $Y2=0
cc_144 N_A_300_21#_c_160_n A2_N 2.90291e-19 $X=1.98 $Y=1.5 $X2=0 $Y2=0
cc_145 N_A_300_21#_c_161_n A2_N 0.0589414f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_300_21#_c_162_n N_A1_N_M1008_g 0.00243271f $X=2.77 $Y=1.98 $X2=0
+ $Y2=0
cc_147 N_A_300_21#_c_161_n N_A1_N_M1012_g 0.0018902f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_148 N_A_300_21#_c_161_n A1_N 0.0676925f $X=2.635 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_300_21#_c_163_n A1_N 0.0147233f $X=2.662 $Y=1.46 $X2=0 $Y2=0
cc_150 N_A_300_21#_c_161_n N_A1_N_c_273_n 0.00127769f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_151 N_A_300_21#_c_163_n N_A1_N_c_273_n 0.00275397f $X=2.662 $Y=1.46 $X2=0
+ $Y2=0
cc_152 N_A_300_21#_M1007_g N_A_222_367#_c_324_n 0.0204804f $X=1.575 $Y=2.155
+ $X2=0 $Y2=0
cc_153 N_A_300_21#_M1009_g N_A_222_367#_c_317_n 0.00934294f $X=1.575 $Y=0.445
+ $X2=0 $Y2=0
cc_154 N_A_300_21#_M1007_g N_A_222_367#_c_317_n 0.00498533f $X=1.575 $Y=2.155
+ $X2=0 $Y2=0
cc_155 N_A_300_21#_c_158_n N_A_222_367#_c_317_n 0.0120248f $X=1.575 $Y=1.5 $X2=0
+ $Y2=0
cc_156 N_A_300_21#_c_159_n N_A_222_367#_c_317_n 0.0189661f $X=2.47 $Y=1.46 $X2=0
+ $Y2=0
cc_157 N_A_300_21#_c_159_n N_A_222_367#_c_326_n 0.0507459f $X=2.47 $Y=1.46 $X2=0
+ $Y2=0
cc_158 N_A_300_21#_c_160_n N_A_222_367#_c_326_n 0.0128567f $X=1.98 $Y=1.5 $X2=0
+ $Y2=0
cc_159 N_A_300_21#_c_162_n N_A_222_367#_c_326_n 0.0101967f $X=2.77 $Y=1.98 $X2=0
+ $Y2=0
cc_160 N_A_300_21#_c_163_n N_A_222_367#_c_326_n 0.00220674f $X=2.662 $Y=1.46
+ $X2=0 $Y2=0
cc_161 N_A_300_21#_M1009_g N_A_222_367#_c_318_n 0.0124737f $X=1.575 $Y=0.445
+ $X2=0 $Y2=0
cc_162 N_A_300_21#_c_159_n N_A_222_367#_c_318_n 0.0058875f $X=2.47 $Y=1.46 $X2=0
+ $Y2=0
cc_163 N_A_300_21#_c_160_n N_A_222_367#_c_318_n 0.00617576f $X=1.98 $Y=1.5 $X2=0
+ $Y2=0
cc_164 N_A_300_21#_c_161_n N_A_222_367#_c_318_n 0.00254815f $X=2.635 $Y=0.445
+ $X2=0 $Y2=0
cc_165 N_A_300_21#_M1009_g N_A_222_367#_c_319_n 0.00826593f $X=1.575 $Y=0.445
+ $X2=0 $Y2=0
cc_166 N_A_300_21#_c_161_n N_A_222_367#_c_319_n 0.00218763f $X=2.635 $Y=0.445
+ $X2=0 $Y2=0
cc_167 N_A_300_21#_M1007_g N_A_222_367#_c_327_n 0.00119967f $X=1.575 $Y=2.155
+ $X2=0 $Y2=0
cc_168 N_A_300_21#_c_162_n N_A_222_367#_c_327_n 0.019289f $X=2.77 $Y=1.98 $X2=0
+ $Y2=0
cc_169 N_A_300_21#_c_162_n N_A_222_367#_c_328_n 0.0147685f $X=2.77 $Y=1.98 $X2=0
+ $Y2=0
cc_170 N_A_300_21#_c_162_n N_A_222_367#_c_330_n 0.0206927f $X=2.77 $Y=1.98 $X2=0
+ $Y2=0
cc_171 N_A_300_21#_c_162_n N_A_222_367#_c_332_n 0.012381f $X=2.77 $Y=1.98 $X2=0
+ $Y2=0
cc_172 N_A_300_21#_c_162_n N_A_222_367#_c_320_n 0.00303848f $X=2.77 $Y=1.98
+ $X2=0 $Y2=0
cc_173 N_A_300_21#_c_163_n N_A_222_367#_c_320_n 0.00237376f $X=2.662 $Y=1.46
+ $X2=0 $Y2=0
cc_174 N_A_300_21#_M1007_g N_A_222_367#_c_334_n 0.0071237f $X=1.575 $Y=2.155
+ $X2=0 $Y2=0
cc_175 N_A_300_21#_M1007_g N_VPWR_c_442_n 0.0064334f $X=1.575 $Y=2.155 $X2=0
+ $Y2=0
cc_176 N_A_300_21#_M1007_g N_VPWR_c_448_n 0.00312414f $X=1.575 $Y=2.155 $X2=0
+ $Y2=0
cc_177 N_A_300_21#_M1007_g N_VPWR_c_440_n 0.00410284f $X=1.575 $Y=2.155 $X2=0
+ $Y2=0
cc_178 N_A_300_21#_M1009_g N_A_67_47#_c_516_n 0.00150647f $X=1.575 $Y=0.445
+ $X2=0 $Y2=0
cc_179 N_A_300_21#_M1009_g N_VGND_c_539_n 0.00119572f $X=1.575 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_300_21#_c_161_n N_VGND_c_540_n 0.00595779f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_181 N_A_300_21#_M1009_g N_VGND_c_545_n 0.00585385f $X=1.575 $Y=0.445 $X2=0
+ $Y2=0
cc_182 N_A_300_21#_c_161_n N_VGND_c_545_n 0.021367f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_183 N_A_300_21#_M1011_s N_VGND_c_548_n 0.00216892f $X=2.51 $Y=0.235 $X2=0
+ $Y2=0
cc_184 N_A_300_21#_M1009_g N_VGND_c_548_n 0.0124078f $X=1.575 $Y=0.445 $X2=0
+ $Y2=0
cc_185 N_A_300_21#_c_161_n N_VGND_c_548_n 0.0143313f $X=2.635 $Y=0.445 $X2=0
+ $Y2=0
cc_186 N_A2_N_c_227_n N_A1_N_M1012_g 0.0498038f $X=2.85 $Y=0.765 $X2=0 $Y2=0
cc_187 N_A2_N_c_229_n N_A1_N_M1012_g 0.00510271f $X=2.555 $Y=0.915 $X2=0 $Y2=0
cc_188 N_A2_N_M1000_g A1_N 2.52419e-19 $X=2.555 $Y=2.155 $X2=0 $Y2=0
cc_189 N_A2_N_c_227_n A1_N 0.00268783f $X=2.85 $Y=0.765 $X2=0 $Y2=0
cc_190 N_A2_N_c_229_n A1_N 6.12914e-19 $X=2.555 $Y=0.915 $X2=0 $Y2=0
cc_191 N_A2_N_M1000_g N_A1_N_c_273_n 0.0307692f $X=2.555 $Y=2.155 $X2=0 $Y2=0
cc_192 N_A2_N_c_229_n N_A1_N_c_273_n 9.98312e-19 $X=2.555 $Y=0.915 $X2=0 $Y2=0
cc_193 N_A2_N_M1000_g N_A_222_367#_c_326_n 0.00593682f $X=2.555 $Y=2.155 $X2=0
+ $Y2=0
cc_194 N_A2_N_c_228_n N_A_222_367#_c_326_n 2.22939e-19 $X=2.48 $Y=0.93 $X2=0
+ $Y2=0
cc_195 N_A2_N_M1000_g N_A_222_367#_c_318_n 4.02953e-19 $X=2.555 $Y=2.155 $X2=0
+ $Y2=0
cc_196 N_A2_N_c_228_n N_A_222_367#_c_318_n 9.16933e-19 $X=2.48 $Y=0.93 $X2=0
+ $Y2=0
cc_197 A2_N N_A_222_367#_c_318_n 0.00785203f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_198 N_A2_N_c_228_n N_A_222_367#_c_319_n 0.0020885f $X=2.48 $Y=0.93 $X2=0
+ $Y2=0
cc_199 A2_N N_A_222_367#_c_319_n 0.0500617f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_200 N_A2_N_M1000_g N_A_222_367#_c_327_n 0.0194725f $X=2.555 $Y=2.155 $X2=0
+ $Y2=0
cc_201 N_A2_N_M1000_g N_A_222_367#_c_328_n 0.00629772f $X=2.555 $Y=2.155 $X2=0
+ $Y2=0
cc_202 N_A2_N_M1000_g N_A_222_367#_c_330_n 5.47226e-19 $X=2.555 $Y=2.155 $X2=0
+ $Y2=0
cc_203 N_A2_N_M1000_g N_VPWR_c_442_n 0.0026354f $X=2.555 $Y=2.155 $X2=0 $Y2=0
cc_204 N_A2_N_M1000_g N_VPWR_c_450_n 2.17715e-19 $X=2.555 $Y=2.155 $X2=0 $Y2=0
cc_205 N_A2_N_c_227_n N_VGND_c_545_n 0.00468185f $X=2.85 $Y=0.765 $X2=0 $Y2=0
cc_206 N_A2_N_c_228_n N_VGND_c_545_n 0.00471202f $X=2.48 $Y=0.93 $X2=0 $Y2=0
cc_207 A2_N N_VGND_c_545_n 0.0106094f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_208 N_A2_N_c_227_n N_VGND_c_548_n 0.00928792f $X=2.85 $Y=0.765 $X2=0 $Y2=0
cc_209 N_A2_N_c_228_n N_VGND_c_548_n 0.00469115f $X=2.48 $Y=0.93 $X2=0 $Y2=0
cc_210 A2_N N_VGND_c_548_n 0.00863123f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_211 N_A1_N_M1012_g N_A_222_367#_c_313_n 0.0195557f $X=3.21 $Y=0.445 $X2=0
+ $Y2=0
cc_212 A1_N N_A_222_367#_c_313_n 0.0010168f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_213 N_A1_N_M1008_g N_A_222_367#_M1005_g 0.00849696f $X=2.985 $Y=2.155 $X2=0
+ $Y2=0
cc_214 N_A1_N_M1008_g N_A_222_367#_c_327_n 5.0589e-19 $X=2.985 $Y=2.155 $X2=0
+ $Y2=0
cc_215 N_A1_N_M1008_g N_A_222_367#_c_328_n 0.00582977f $X=2.985 $Y=2.155 $X2=0
+ $Y2=0
cc_216 N_A1_N_M1008_g N_A_222_367#_c_330_n 0.0192257f $X=2.985 $Y=2.155 $X2=0
+ $Y2=0
cc_217 A1_N N_A_222_367#_c_331_n 0.00227977f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_218 N_A1_N_c_273_n N_A_222_367#_c_331_n 0.00231634f $X=3.21 $Y=1.35 $X2=0
+ $Y2=0
cc_219 N_A1_N_M1008_g N_A_222_367#_c_332_n 0.00556971f $X=2.985 $Y=2.155 $X2=0
+ $Y2=0
cc_220 A1_N N_A_222_367#_c_332_n 0.0150437f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_221 N_A1_N_c_273_n N_A_222_367#_c_332_n 0.00114102f $X=3.21 $Y=1.35 $X2=0
+ $Y2=0
cc_222 N_A1_N_M1008_g N_A_222_367#_c_320_n 0.00152908f $X=2.985 $Y=2.155 $X2=0
+ $Y2=0
cc_223 A1_N N_A_222_367#_c_320_n 0.0166783f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_224 N_A1_N_c_273_n N_A_222_367#_c_320_n 0.00122371f $X=3.21 $Y=1.35 $X2=0
+ $Y2=0
cc_225 A1_N N_A_222_367#_c_321_n 0.00123535f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_226 N_A1_N_c_273_n N_A_222_367#_c_321_n 0.0217704f $X=3.21 $Y=1.35 $X2=0
+ $Y2=0
cc_227 N_A1_N_M1008_g N_VPWR_c_443_n 0.00185967f $X=2.985 $Y=2.155 $X2=0 $Y2=0
cc_228 N_A1_N_M1008_g N_VPWR_c_450_n 2.35436e-19 $X=2.985 $Y=2.155 $X2=0 $Y2=0
cc_229 N_A1_N_M1012_g N_VGND_c_540_n 0.0108425f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_230 A1_N N_VGND_c_540_n 0.0415804f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_231 N_A1_N_M1012_g N_VGND_c_545_n 0.00462105f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_232 A1_N N_VGND_c_545_n 0.00510013f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_233 N_A1_N_M1012_g N_VGND_c_548_n 0.00768096f $X=3.21 $Y=0.445 $X2=0 $Y2=0
cc_234 A1_N N_VGND_c_548_n 0.00660835f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_235 A1_N A_585_47# 0.00228524f $X=3.035 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_236 N_A_222_367#_c_326_n N_VPWR_M1007_d 0.016829f $X=2.325 $Y=1.84 $X2=0
+ $Y2=0
cc_237 N_A_222_367#_c_327_n N_VPWR_M1007_d 0.00673251f $X=2.41 $Y=2.665 $X2=0
+ $Y2=0
cc_238 N_A_222_367#_c_330_n N_VPWR_M1008_d 0.00691935f $X=3.12 $Y=2.665 $X2=0
+ $Y2=0
cc_239 N_A_222_367#_c_331_n N_VPWR_M1008_d 0.00990497f $X=3.495 $Y=1.77 $X2=0
+ $Y2=0
cc_240 N_A_222_367#_c_324_n N_VPWR_c_441_n 0.00974231f $X=1.305 $Y=1.98 $X2=0
+ $Y2=0
cc_241 N_A_222_367#_c_324_n N_VPWR_c_442_n 0.0186408f $X=1.305 $Y=1.98 $X2=0
+ $Y2=0
cc_242 N_A_222_367#_c_326_n N_VPWR_c_442_n 0.0266856f $X=2.325 $Y=1.84 $X2=0
+ $Y2=0
cc_243 N_A_222_367#_c_327_n N_VPWR_c_442_n 0.0440661f $X=2.41 $Y=2.665 $X2=0
+ $Y2=0
cc_244 N_A_222_367#_c_329_n N_VPWR_c_442_n 0.0150385f $X=2.495 $Y=2.75 $X2=0
+ $Y2=0
cc_245 N_A_222_367#_M1005_g N_VPWR_c_443_n 0.0173688f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_246 N_A_222_367#_M1013_g N_VPWR_c_443_n 8.49233e-19 $X=4.225 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_A_222_367#_c_328_n N_VPWR_c_443_n 0.0151624f $X=3.035 $Y=2.75 $X2=0
+ $Y2=0
cc_248 N_A_222_367#_c_330_n N_VPWR_c_443_n 0.0498641f $X=3.12 $Y=2.665 $X2=0
+ $Y2=0
cc_249 N_A_222_367#_c_331_n N_VPWR_c_443_n 0.0267628f $X=3.495 $Y=1.77 $X2=0
+ $Y2=0
cc_250 N_A_222_367#_c_321_n N_VPWR_c_443_n 7.7289e-19 $X=4.225 $Y=1.35 $X2=0
+ $Y2=0
cc_251 N_A_222_367#_M1013_g N_VPWR_c_445_n 0.00720926f $X=4.225 $Y=2.465 $X2=0
+ $Y2=0
cc_252 N_A_222_367#_c_328_n N_VPWR_c_450_n 0.0184403f $X=3.035 $Y=2.75 $X2=0
+ $Y2=0
cc_253 N_A_222_367#_c_329_n N_VPWR_c_450_n 0.00476346f $X=2.495 $Y=2.75 $X2=0
+ $Y2=0
cc_254 N_A_222_367#_M1005_g N_VPWR_c_451_n 0.00486043f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_255 N_A_222_367#_M1013_g N_VPWR_c_451_n 0.00533769f $X=4.225 $Y=2.465 $X2=0
+ $Y2=0
cc_256 N_A_222_367#_M1005_g N_VPWR_c_440_n 0.00824727f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_A_222_367#_M1013_g N_VPWR_c_440_n 0.0104368f $X=4.225 $Y=2.465 $X2=0
+ $Y2=0
cc_258 N_A_222_367#_c_324_n N_VPWR_c_440_n 0.020087f $X=1.305 $Y=1.98 $X2=0
+ $Y2=0
cc_259 N_A_222_367#_c_328_n N_VPWR_c_440_n 0.0228785f $X=3.035 $Y=2.75 $X2=0
+ $Y2=0
cc_260 N_A_222_367#_c_329_n N_VPWR_c_440_n 0.00570745f $X=2.495 $Y=2.75 $X2=0
+ $Y2=0
cc_261 N_A_222_367#_c_313_n N_X_c_498_n 0.00339384f $X=3.795 $Y=1.185 $X2=0
+ $Y2=0
cc_262 N_A_222_367#_M1005_g N_X_c_498_n 0.00301993f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_263 N_A_222_367#_c_315_n N_X_c_498_n 0.0157796f $X=4.225 $Y=1.185 $X2=0 $Y2=0
cc_264 N_A_222_367#_M1013_g N_X_c_498_n 0.0318546f $X=4.225 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A_222_367#_c_331_n N_X_c_498_n 0.0132472f $X=3.495 $Y=1.77 $X2=0 $Y2=0
cc_266 N_A_222_367#_c_320_n N_X_c_498_n 0.0367766f $X=3.66 $Y=1.35 $X2=0 $Y2=0
cc_267 N_A_222_367#_c_321_n N_X_c_498_n 0.0309552f $X=4.225 $Y=1.35 $X2=0 $Y2=0
cc_268 N_A_222_367#_c_318_n N_A_67_47#_c_516_n 0.00207487f $X=1.777 $Y=0.995
+ $X2=0 $Y2=0
cc_269 N_A_222_367#_c_319_n N_A_67_47#_c_516_n 0.0145852f $X=1.79 $Y=0.445 $X2=0
+ $Y2=0
cc_270 N_A_222_367#_c_313_n N_VGND_c_540_n 0.018226f $X=3.795 $Y=1.185 $X2=0
+ $Y2=0
cc_271 N_A_222_367#_c_315_n N_VGND_c_540_n 7.52068e-19 $X=4.225 $Y=1.185 $X2=0
+ $Y2=0
cc_272 N_A_222_367#_c_331_n N_VGND_c_540_n 0.00278385f $X=3.495 $Y=1.77 $X2=0
+ $Y2=0
cc_273 N_A_222_367#_c_320_n N_VGND_c_540_n 0.0189748f $X=3.66 $Y=1.35 $X2=0
+ $Y2=0
cc_274 N_A_222_367#_c_321_n N_VGND_c_540_n 0.00160017f $X=4.225 $Y=1.35 $X2=0
+ $Y2=0
cc_275 N_A_222_367#_c_315_n N_VGND_c_542_n 0.00663461f $X=4.225 $Y=1.185 $X2=0
+ $Y2=0
cc_276 N_A_222_367#_c_319_n N_VGND_c_545_n 0.0127882f $X=1.79 $Y=0.445 $X2=0
+ $Y2=0
cc_277 N_A_222_367#_c_313_n N_VGND_c_546_n 0.00486043f $X=3.795 $Y=1.185 $X2=0
+ $Y2=0
cc_278 N_A_222_367#_c_315_n N_VGND_c_546_n 0.00533769f $X=4.225 $Y=1.185 $X2=0
+ $Y2=0
cc_279 N_A_222_367#_M1009_d N_VGND_c_548_n 0.003281f $X=1.65 $Y=0.235 $X2=0
+ $Y2=0
cc_280 N_A_222_367#_c_313_n N_VGND_c_548_n 0.00824727f $X=3.795 $Y=1.185 $X2=0
+ $Y2=0
cc_281 N_A_222_367#_c_315_n N_VGND_c_548_n 0.0104368f $X=4.225 $Y=1.185 $X2=0
+ $Y2=0
cc_282 N_A_222_367#_c_319_n N_VGND_c_548_n 0.00896147f $X=1.79 $Y=0.445 $X2=0
+ $Y2=0
cc_283 N_VPWR_c_440_n N_X_M1005_s 0.00380103f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_284 N_VPWR_c_445_n N_X_c_498_n 0.0466048f $X=4.44 $Y=1.98 $X2=0 $Y2=0
cc_285 N_VPWR_c_451_n N_X_c_498_n 0.0163698f $X=4.355 $Y=3.33 $X2=0 $Y2=0
cc_286 N_VPWR_c_440_n N_X_c_498_n 0.0101905f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_287 N_X_c_498_n N_VGND_c_542_n 0.0313225f $X=4.01 $Y=0.42 $X2=0 $Y2=0
cc_288 N_X_c_498_n N_VGND_c_546_n 0.0163698f $X=4.01 $Y=0.42 $X2=0 $Y2=0
cc_289 N_X_M1002_d N_VGND_c_548_n 0.00380103f $X=3.87 $Y=0.235 $X2=0 $Y2=0
cc_290 N_X_c_498_n N_VGND_c_548_n 0.0101905f $X=4.01 $Y=0.42 $X2=0 $Y2=0
cc_291 N_A_67_47#_c_516_n N_VGND_c_539_n 0.02044f $X=1.245 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A_67_47#_c_515_n N_VGND_c_543_n 0.0157295f $X=0.46 $Y=0.445 $X2=0 $Y2=0
cc_293 N_A_67_47#_c_516_n N_VGND_c_543_n 0.00268101f $X=1.245 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_67_47#_c_516_n N_VGND_c_545_n 0.00268101f $X=1.245 $Y=0.74 $X2=0
+ $Y2=0
cc_295 N_A_67_47#_c_533_p N_VGND_c_545_n 0.012276f $X=1.36 $Y=0.445 $X2=0 $Y2=0
cc_296 N_A_67_47#_M1004_s N_VGND_c_548_n 0.00225688f $X=0.335 $Y=0.235 $X2=0
+ $Y2=0
cc_297 N_A_67_47#_M1003_d N_VGND_c_548_n 0.00273173f $X=1.22 $Y=0.235 $X2=0
+ $Y2=0
cc_298 N_A_67_47#_c_515_n N_VGND_c_548_n 0.0106102f $X=0.46 $Y=0.445 $X2=0 $Y2=0
cc_299 N_A_67_47#_c_516_n N_VGND_c_548_n 0.00958291f $X=1.245 $Y=0.74 $X2=0
+ $Y2=0
cc_300 N_A_67_47#_c_533_p N_VGND_c_548_n 0.00927439f $X=1.36 $Y=0.445 $X2=0
+ $Y2=0
cc_301 N_VGND_c_548_n A_585_47# 0.00535573f $X=4.56 $Y=0 $X2=-0.19 $Y2=-0.245
