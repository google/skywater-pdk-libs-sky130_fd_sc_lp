* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a22oi_0 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 a_45_405# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=5.408e+11p pd=5.53e+06u as=1.792e+11p ps=1.84e+06u
M1001 VGND A2 a_307_47# VNB nshort w=420000u l=150000u
+  ad=2.457e+11p pd=2.85e+06u as=8.82e+10p ps=1.26e+06u
M1002 VPWR A1 a_45_405# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B1 a_121_47# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=8.82e+10p ps=1.26e+06u
M1004 Y B2 a_45_405# VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1005 a_45_405# B1 Y VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_121_47# B2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_307_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
