* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor2_lp A B VNB VPB Y
X0 Y B a_294_112# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_294_112# B VNB SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VNB A a_130_112# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_130_490# B Y w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_130_112# A Y SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPB A a_130_490# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
