* File: sky130_fd_sc_lp__einvn_8.pex.spice
* Created: Wed Sep  2 09:51:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVN_8%A_110_57# 1 2 7 8 9 11 12 14 16 17 19 21 22
+ 24 26 27 29 31 32 34 36 37 39 41 42 44 46 48 49 50 51 52 53 54 57 61 69 70
c142 42 0 7.28141e-20 $X=4.8 $Y=1.265
c143 37 0 1.4515e-19 $X=4.37 $Y=1.265
c144 27 0 1.4515e-19 $X=3.51 $Y=1.265
c145 17 0 1.4515e-19 $X=2.65 $Y=1.265
c146 7 0 1.99871e-19 $X=1.79 $Y=1.265
r147 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=0.83 $X2=1.15 $Y2=0.83
r148 61 63 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=1.15 $Y=1.98
+ $X2=1.15 $Y2=2.91
r149 59 69 1.48468 $w=3.3e-07 $l=1.88e-07 $layer=LI1_cond $X=1.15 $Y=1.04
+ $X2=1.15 $Y2=0.852
r150 59 61 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=1.15 $Y=1.04
+ $X2=1.15 $Y2=1.98
r151 55 69 14.1366 $w=3.73e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.852
+ $X2=1.15 $Y2=0.852
r152 55 57 12.4113 $w=2.08e-07 $l=2.35e-07 $layer=LI1_cond $X=0.69 $Y=0.665
+ $X2=0.69 $Y2=0.43
r153 47 70 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.15 $Y=1.185
+ $X2=1.15 $Y2=0.83
r154 44 46 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.875 $Y=1.185
+ $X2=4.875 $Y2=0.655
r155 43 54 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=4.52 $Y=1.265
+ $X2=4.445 $Y2=1.265
r156 42 44 26.9672 $w=1.6e-07 $l=1.11355e-07 $layer=POLY_cond $X=4.8 $Y=1.265
+ $X2=4.875 $Y2=1.185
r157 42 43 129.769 $w=1.6e-07 $l=2.8e-07 $layer=POLY_cond $X=4.8 $Y=1.265
+ $X2=4.52 $Y2=1.265
r158 39 54 6.22635 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=4.445 $Y=1.185
+ $X2=4.445 $Y2=1.265
r159 39 41 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.445 $Y=1.185
+ $X2=4.445 $Y2=0.655
r160 38 53 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=4.09 $Y=1.265
+ $X2=4.015 $Y2=1.265
r161 37 54 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=4.37 $Y=1.265
+ $X2=4.445 $Y2=1.265
r162 37 38 129.769 $w=1.6e-07 $l=2.8e-07 $layer=POLY_cond $X=4.37 $Y=1.265
+ $X2=4.09 $Y2=1.265
r163 34 53 6.22635 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=4.015 $Y=1.185
+ $X2=4.015 $Y2=1.265
r164 34 36 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.015 $Y=1.185
+ $X2=4.015 $Y2=0.655
r165 33 52 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=3.66 $Y=1.265
+ $X2=3.585 $Y2=1.265
r166 32 53 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=3.94 $Y=1.265
+ $X2=4.015 $Y2=1.265
r167 32 33 129.769 $w=1.6e-07 $l=2.8e-07 $layer=POLY_cond $X=3.94 $Y=1.265
+ $X2=3.66 $Y2=1.265
r168 29 52 6.22635 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=3.585 $Y=1.185
+ $X2=3.585 $Y2=1.265
r169 29 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.585 $Y=1.185
+ $X2=3.585 $Y2=0.655
r170 28 51 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=3.23 $Y=1.265
+ $X2=3.155 $Y2=1.265
r171 27 52 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=3.51 $Y=1.265
+ $X2=3.585 $Y2=1.265
r172 27 28 129.769 $w=1.6e-07 $l=2.8e-07 $layer=POLY_cond $X=3.51 $Y=1.265
+ $X2=3.23 $Y2=1.265
r173 24 51 6.22635 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=3.155 $Y=1.185
+ $X2=3.155 $Y2=1.265
r174 24 26 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.155 $Y=1.185
+ $X2=3.155 $Y2=0.655
r175 23 50 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=2.8 $Y=1.265
+ $X2=2.725 $Y2=1.265
r176 22 51 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=3.08 $Y=1.265
+ $X2=3.155 $Y2=1.265
r177 22 23 129.769 $w=1.6e-07 $l=2.8e-07 $layer=POLY_cond $X=3.08 $Y=1.265
+ $X2=2.8 $Y2=1.265
r178 19 50 6.22635 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=2.725 $Y=1.185
+ $X2=2.725 $Y2=1.265
r179 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.725 $Y=1.185
+ $X2=2.725 $Y2=0.655
r180 18 49 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=1.265
+ $X2=2.295 $Y2=1.265
r181 17 50 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=2.65 $Y=1.265
+ $X2=2.725 $Y2=1.265
r182 17 18 129.769 $w=1.6e-07 $l=2.8e-07 $layer=POLY_cond $X=2.65 $Y=1.265
+ $X2=2.37 $Y2=1.265
r183 14 49 6.22635 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=2.295 $Y=1.185
+ $X2=2.295 $Y2=1.265
r184 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.295 $Y=1.185
+ $X2=2.295 $Y2=0.655
r185 13 48 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=1.94 $Y=1.265
+ $X2=1.865 $Y2=1.265
r186 12 49 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=2.22 $Y=1.265
+ $X2=2.295 $Y2=1.265
r187 12 13 129.769 $w=1.6e-07 $l=2.8e-07 $layer=POLY_cond $X=2.22 $Y=1.265
+ $X2=1.94 $Y2=1.265
r188 9 48 6.22635 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=1.865 $Y=1.185
+ $X2=1.865 $Y2=1.265
r189 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.865 $Y=1.185
+ $X2=1.865 $Y2=0.655
r190 8 47 31.3783 $w=1.6e-07 $l=2.0106e-07 $layer=POLY_cond $X=1.315 $Y=1.265
+ $X2=1.15 $Y2=1.185
r191 7 48 19.3363 $w=1.6e-07 $l=7.5e-08 $layer=POLY_cond $X=1.79 $Y=1.265
+ $X2=1.865 $Y2=1.265
r192 7 8 220.144 $w=1.6e-07 $l=4.75e-07 $layer=POLY_cond $X=1.79 $Y=1.265
+ $X2=1.315 $Y2=1.265
r193 2 63 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=2.91
r194 2 61 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=1.98
r195 1 55 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.285 $X2=0.69 $Y2=0.875
r196 1 57 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.285 $X2=0.69 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_8%TE_B 3 5 7 8 9 10 12 13 15 17 18 20 22 23 25
+ 27 28 30 32 33 35 37 38 40 42 43 45 47 48 49 50 51 52 53 54 55 57 58 59 69 73
c160 43 0 1.19405e-19 $X=4.8 $Y=1.64
r161 71 85 2.72196 $w=3.1e-07 $l=2.18e-07 $layer=LI1_cond $X=0.26 $Y=1.645
+ $X2=0.26 $Y2=1.427
r162 71 73 0.743512 $w=3.08e-07 $l=2e-08 $layer=LI1_cond $X=0.26 $Y=1.645
+ $X2=0.26 $Y2=1.665
r163 69 85 9.27253 $w=4.33e-07 $l=3.5e-07 $layer=LI1_cond $X=0.61 $Y=1.427
+ $X2=0.26 $Y2=1.427
r164 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.46 $X2=0.61 $Y2=1.46
r165 66 68 17.7787 $w=3.66e-07 $l=1.35e-07 $layer=POLY_cond $X=0.475 $Y=1.51
+ $X2=0.61 $Y2=1.51
r166 58 59 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.775
r167 57 58 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.035
+ $X2=0.26 $Y2=2.405
r168 55 85 0.529859 $w=4.33e-07 $l=2e-08 $layer=LI1_cond $X=0.24 $Y=1.427
+ $X2=0.26 $Y2=1.427
r169 55 57 12.5653 $w=3.08e-07 $l=3.38e-07 $layer=LI1_cond $X=0.26 $Y=1.697
+ $X2=0.26 $Y2=2.035
r170 55 73 1.18962 $w=3.08e-07 $l=3.2e-08 $layer=LI1_cond $X=0.26 $Y=1.697
+ $X2=0.26 $Y2=1.665
r171 45 47 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.875 $Y=1.725
+ $X2=4.875 $Y2=2.465
r172 44 54 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.52 $Y=1.64
+ $X2=4.445 $Y2=1.64
r173 43 45 27.0678 $w=1.7e-07 $l=1.16619e-07 $layer=POLY_cond $X=4.8 $Y=1.64
+ $X2=4.875 $Y2=1.725
r174 43 44 118.386 $w=1.7e-07 $l=2.8e-07 $layer=POLY_cond $X=4.8 $Y=1.64
+ $X2=4.52 $Y2=1.64
r175 40 54 7.09928 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=4.445 $Y=1.725
+ $X2=4.445 $Y2=1.64
r176 40 42 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.445 $Y=1.725
+ $X2=4.445 $Y2=2.465
r177 39 53 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.09 $Y=1.64
+ $X2=4.015 $Y2=1.64
r178 38 54 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=4.37 $Y=1.64
+ $X2=4.445 $Y2=1.64
r179 38 39 118.386 $w=1.7e-07 $l=2.8e-07 $layer=POLY_cond $X=4.37 $Y=1.64
+ $X2=4.09 $Y2=1.64
r180 35 53 7.09928 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=4.015 $Y=1.725
+ $X2=4.015 $Y2=1.64
r181 35 37 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.015 $Y=1.725
+ $X2=4.015 $Y2=2.465
r182 34 52 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.66 $Y=1.64
+ $X2=3.585 $Y2=1.64
r183 33 53 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.94 $Y=1.64
+ $X2=4.015 $Y2=1.64
r184 33 34 118.386 $w=1.7e-07 $l=2.8e-07 $layer=POLY_cond $X=3.94 $Y=1.64
+ $X2=3.66 $Y2=1.64
r185 30 52 7.09928 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=3.585 $Y=1.725
+ $X2=3.585 $Y2=1.64
r186 30 32 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.585 $Y=1.725
+ $X2=3.585 $Y2=2.465
r187 29 51 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.23 $Y=1.64
+ $X2=3.155 $Y2=1.64
r188 28 52 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.51 $Y=1.64
+ $X2=3.585 $Y2=1.64
r189 28 29 118.386 $w=1.7e-07 $l=2.8e-07 $layer=POLY_cond $X=3.51 $Y=1.64
+ $X2=3.23 $Y2=1.64
r190 25 51 7.09928 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=3.155 $Y=1.725
+ $X2=3.155 $Y2=1.64
r191 25 27 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.155 $Y=1.725
+ $X2=3.155 $Y2=2.465
r192 24 50 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.8 $Y=1.64
+ $X2=2.725 $Y2=1.64
r193 23 51 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=3.08 $Y=1.64
+ $X2=3.155 $Y2=1.64
r194 23 24 118.386 $w=1.7e-07 $l=2.8e-07 $layer=POLY_cond $X=3.08 $Y=1.64
+ $X2=2.8 $Y2=1.64
r195 20 50 7.09928 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=2.725 $Y=1.725
+ $X2=2.725 $Y2=1.64
r196 20 22 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.725 $Y=1.725
+ $X2=2.725 $Y2=2.465
r197 19 49 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=1.64
+ $X2=2.295 $Y2=1.64
r198 18 50 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.65 $Y=1.64
+ $X2=2.725 $Y2=1.64
r199 18 19 118.386 $w=1.7e-07 $l=2.8e-07 $layer=POLY_cond $X=2.65 $Y=1.64
+ $X2=2.37 $Y2=1.64
r200 15 49 7.09928 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=2.295 $Y=1.725
+ $X2=2.295 $Y2=1.64
r201 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.295 $Y=1.725
+ $X2=2.295 $Y2=2.465
r202 14 48 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.94 $Y=1.64
+ $X2=1.865 $Y2=1.64
r203 13 49 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=2.22 $Y=1.64
+ $X2=2.295 $Y2=1.64
r204 13 14 118.386 $w=1.7e-07 $l=2.8e-07 $layer=POLY_cond $X=2.22 $Y=1.64
+ $X2=1.94 $Y2=1.64
r205 10 48 7.09928 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.865 $Y=1.725
+ $X2=1.865 $Y2=1.64
r206 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.865 $Y=1.725
+ $X2=1.865 $Y2=2.465
r207 8 48 18.3685 $w=1.7e-07 $l=7.5e-08 $layer=POLY_cond $X=1.79 $Y=1.64
+ $X2=1.865 $Y2=1.64
r208 8 9 338.246 $w=1.7e-07 $l=8e-07 $layer=POLY_cond $X=1.79 $Y=1.64 $X2=0.99
+ $Y2=1.64
r209 5 9 23.8115 $w=3.66e-07 $l=1.16619e-07 $layer=POLY_cond $X=0.915 $Y=1.725
+ $X2=0.99 $Y2=1.64
r210 5 68 40.1667 $w=3.66e-07 $l=3.98246e-07 $layer=POLY_cond $X=0.915 $Y=1.725
+ $X2=0.61 $Y2=1.51
r211 5 7 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.915 $Y=1.725
+ $X2=0.915 $Y2=2.465
r212 1 66 23.7042 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=1.51
r213 1 3 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=0.705
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_8%A 1 3 6 8 10 13 15 17 20 22 24 27 29 31 34
+ 36 38 41 43 45 48 50 52 55 57 58 72
c140 58 0 7.28141e-20 $X=6 $Y=1.295
r141 71 72 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.885 $Y=1.35
+ $X2=8.315 $Y2=1.35
r142 70 71 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.455 $Y=1.35
+ $X2=7.885 $Y2=1.35
r143 69 70 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.025 $Y=1.35
+ $X2=7.455 $Y2=1.35
r144 68 69 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.595 $Y=1.35
+ $X2=7.025 $Y2=1.35
r145 67 68 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.165 $Y=1.35
+ $X2=6.595 $Y2=1.35
r146 65 67 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=5.85 $Y=1.35
+ $X2=6.165 $Y2=1.35
r147 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.85
+ $Y=1.35 $X2=5.85 $Y2=1.35
r148 63 65 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.735 $Y=1.35
+ $X2=5.85 $Y2=1.35
r149 61 63 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.305 $Y=1.35
+ $X2=5.735 $Y2=1.35
r150 58 66 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6 $Y=1.35 $X2=5.85
+ $Y2=1.35
r151 57 66 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.52 $Y=1.35
+ $X2=5.85 $Y2=1.35
r152 53 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.315 $Y=1.515
+ $X2=8.315 $Y2=1.35
r153 53 55 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.315 $Y=1.515
+ $X2=8.315 $Y2=2.465
r154 50 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.315 $Y=1.185
+ $X2=8.315 $Y2=1.35
r155 50 52 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.315 $Y=1.185
+ $X2=8.315 $Y2=0.655
r156 46 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.885 $Y=1.515
+ $X2=7.885 $Y2=1.35
r157 46 48 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.885 $Y=1.515
+ $X2=7.885 $Y2=2.465
r158 43 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.885 $Y=1.185
+ $X2=7.885 $Y2=1.35
r159 43 45 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.885 $Y=1.185
+ $X2=7.885 $Y2=0.655
r160 39 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.455 $Y=1.515
+ $X2=7.455 $Y2=1.35
r161 39 41 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.455 $Y=1.515
+ $X2=7.455 $Y2=2.465
r162 36 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.455 $Y=1.185
+ $X2=7.455 $Y2=1.35
r163 36 38 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.455 $Y=1.185
+ $X2=7.455 $Y2=0.655
r164 32 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.515
+ $X2=7.025 $Y2=1.35
r165 32 34 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.025 $Y=1.515
+ $X2=7.025 $Y2=2.465
r166 29 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.185
+ $X2=7.025 $Y2=1.35
r167 29 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.025 $Y=1.185
+ $X2=7.025 $Y2=0.655
r168 25 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.515
+ $X2=6.595 $Y2=1.35
r169 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.595 $Y=1.515
+ $X2=6.595 $Y2=2.465
r170 22 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.185
+ $X2=6.595 $Y2=1.35
r171 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.595 $Y=1.185
+ $X2=6.595 $Y2=0.655
r172 18 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.165 $Y=1.515
+ $X2=6.165 $Y2=1.35
r173 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.165 $Y=1.515
+ $X2=6.165 $Y2=2.465
r174 15 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.165 $Y=1.185
+ $X2=6.165 $Y2=1.35
r175 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.165 $Y=1.185
+ $X2=6.165 $Y2=0.655
r176 11 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=1.515
+ $X2=5.735 $Y2=1.35
r177 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.735 $Y=1.515
+ $X2=5.735 $Y2=2.465
r178 8 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=1.185
+ $X2=5.735 $Y2=1.35
r179 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.735 $Y=1.185
+ $X2=5.735 $Y2=0.655
r180 4 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.515
+ $X2=5.305 $Y2=1.35
r181 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.305 $Y=1.515
+ $X2=5.305 $Y2=2.465
r182 1 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.185
+ $X2=5.305 $Y2=1.35
r183 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.305 $Y=1.185
+ $X2=5.305 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_8%VPWR 1 2 3 4 5 18 24 30 36 40 44 49 50 51 52
+ 53 55 60 77 78 81 84 87
r128 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 77 78 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r131 75 78 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=8.88 $Y2=3.33
r132 74 77 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=8.88 $Y2=3.33
r133 74 75 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r134 72 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=3.33
+ $X2=4.66 $Y2=3.33
r135 72 74 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.825 $Y=3.33
+ $X2=5.04 $Y2=3.33
r136 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r137 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r138 68 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r139 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r140 65 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.08 $Y2=3.33
r141 65 67 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.64 $Y2=3.33
r142 64 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r143 64 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r144 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r145 61 81 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.7 $Y2=3.33
r146 61 63 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r147 60 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=2.08 $Y2=3.33
r148 60 63 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r149 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r150 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r151 55 81 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.7 $Y2=3.33
r152 55 57 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.24 $Y2=3.33
r153 53 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r154 53 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r155 53 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r156 51 70 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.635 $Y=3.33
+ $X2=3.6 $Y2=3.33
r157 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=3.33
+ $X2=3.8 $Y2=3.33
r158 49 67 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.64 $Y2=3.33
r159 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.94 $Y2=3.33
r160 48 70 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=3.6 $Y2=3.33
r161 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=2.94 $Y2=3.33
r162 44 47 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=4.66 $Y=2.18
+ $X2=4.66 $Y2=2.95
r163 42 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=3.245
+ $X2=4.66 $Y2=3.33
r164 42 47 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.66 $Y=3.245
+ $X2=4.66 $Y2=2.95
r165 41 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=3.8 $Y2=3.33
r166 40 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=3.33
+ $X2=4.66 $Y2=3.33
r167 40 41 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.495 $Y=3.33
+ $X2=3.965 $Y2=3.33
r168 36 39 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.8 $Y=2.18 $X2=3.8
+ $Y2=2.95
r169 34 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=3.245 $X2=3.8
+ $Y2=3.33
r170 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.8 $Y=3.245
+ $X2=3.8 $Y2=2.95
r171 30 33 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.94 $Y=2.18
+ $X2=2.94 $Y2=2.95
r172 28 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=3.245
+ $X2=2.94 $Y2=3.33
r173 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.94 $Y=3.245
+ $X2=2.94 $Y2=2.95
r174 24 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.08 $Y=2.18
+ $X2=2.08 $Y2=2.95
r175 22 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=3.33
r176 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=2.95
r177 18 21 51.2294 $w=2.08e-07 $l=9.7e-07 $layer=LI1_cond $X=0.7 $Y=1.98 $X2=0.7
+ $Y2=2.95
r178 16 81 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=3.245
+ $X2=0.7 $Y2=3.33
r179 16 21 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=3.245
+ $X2=0.7 $Y2=2.95
r180 5 47 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.835 $X2=4.66 $Y2=2.95
r181 5 44 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.835 $X2=4.66 $Y2=2.18
r182 4 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=1.835 $X2=3.8 $Y2=2.95
r183 4 36 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=1.835 $X2=3.8 $Y2=2.18
r184 3 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.835 $X2=2.94 $Y2=2.95
r185 3 30 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=2.8
+ $Y=1.835 $X2=2.94 $Y2=2.18
r186 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.08 $Y2=2.95
r187 2 24 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=1.835 $X2=2.08 $Y2=2.18
r188 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.7 $Y2=2.95
r189 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.7 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_8%A_305_367# 1 2 3 4 5 6 7 8 9 30 34 35 38 42
+ 46 50 54 58 61 64 68 72 76 80 84 88 90 92 94 95 96 99 100 101
c129 96 0 1.4515e-19 $X=4.23 $Y=1.8
c130 95 0 1.4515e-19 $X=3.37 $Y=1.8
c131 94 0 1.4515e-19 $X=2.51 $Y=1.8
c132 35 0 1.99871e-19 $X=1.745 $Y=1.8
r133 90 103 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.565 $Y=2.905
+ $X2=8.565 $Y2=2.99
r134 90 92 40.5571 $w=2.58e-07 $l=9.15e-07 $layer=LI1_cond $X=8.565 $Y=2.905
+ $X2=8.565 $Y2=1.99
r135 89 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.765 $Y=2.99
+ $X2=7.67 $Y2=2.99
r136 88 103 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.435 $Y=2.99
+ $X2=8.565 $Y2=2.99
r137 88 89 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.435 $Y=2.99
+ $X2=7.765 $Y2=2.99
r138 84 87 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=7.67 $Y=2.22
+ $X2=7.67 $Y2=2.9
r139 82 101 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=2.905
+ $X2=7.67 $Y2=2.99
r140 82 87 0.291866 $w=1.88e-07 $l=5e-09 $layer=LI1_cond $X=7.67 $Y=2.905
+ $X2=7.67 $Y2=2.9
r141 81 100 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.905 $Y=2.99
+ $X2=6.81 $Y2=2.99
r142 80 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.575 $Y=2.99
+ $X2=7.67 $Y2=2.99
r143 80 81 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.575 $Y=2.99
+ $X2=6.905 $Y2=2.99
r144 76 79 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=6.81 $Y=2.22
+ $X2=6.81 $Y2=2.9
r145 74 100 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.81 $Y=2.905
+ $X2=6.81 $Y2=2.99
r146 74 79 0.291866 $w=1.88e-07 $l=5e-09 $layer=LI1_cond $X=6.81 $Y=2.905
+ $X2=6.81 $Y2=2.9
r147 73 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.045 $Y=2.99
+ $X2=5.95 $Y2=2.99
r148 72 100 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.715 $Y=2.99
+ $X2=6.81 $Y2=2.99
r149 72 73 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.715 $Y=2.99
+ $X2=6.045 $Y2=2.99
r150 68 71 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=5.95 $Y=2.22
+ $X2=5.95 $Y2=2.9
r151 66 99 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=2.905
+ $X2=5.95 $Y2=2.99
r152 66 71 0.291866 $w=1.88e-07 $l=5e-09 $layer=LI1_cond $X=5.95 $Y=2.905
+ $X2=5.95 $Y2=2.9
r153 65 98 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.185 $Y=2.99
+ $X2=5.09 $Y2=2.99
r154 64 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.855 $Y=2.99
+ $X2=5.95 $Y2=2.99
r155 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.855 $Y=2.99
+ $X2=5.185 $Y2=2.99
r156 61 98 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=2.905
+ $X2=5.09 $Y2=2.99
r157 61 63 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=5.09 $Y=2.905
+ $X2=5.09 $Y2=1.98
r158 60 63 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=5.09 $Y=1.925
+ $X2=5.09 $Y2=1.98
r159 59 96 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.325 $Y=1.8
+ $X2=4.23 $Y2=1.8
r160 58 60 6.98266 $w=2.5e-07 $l=1.65831e-07 $layer=LI1_cond $X=4.995 $Y=1.8
+ $X2=5.09 $Y2=1.925
r161 58 59 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=4.995 $Y=1.8
+ $X2=4.325 $Y2=1.8
r162 54 56 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=4.23 $Y=1.98
+ $X2=4.23 $Y2=2.91
r163 52 96 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=4.23 $Y=1.925
+ $X2=4.23 $Y2=1.8
r164 52 54 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=4.23 $Y=1.925
+ $X2=4.23 $Y2=1.98
r165 51 95 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=3.465 $Y=1.8
+ $X2=3.37 $Y2=1.8
r166 50 96 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.135 $Y=1.8
+ $X2=4.23 $Y2=1.8
r167 50 51 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=4.135 $Y=1.8
+ $X2=3.465 $Y2=1.8
r168 46 48 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.37 $Y=1.98
+ $X2=3.37 $Y2=2.91
r169 44 95 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.37 $Y=1.925
+ $X2=3.37 $Y2=1.8
r170 44 46 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=3.37 $Y=1.925
+ $X2=3.37 $Y2=1.98
r171 43 94 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=2.605 $Y=1.8
+ $X2=2.51 $Y2=1.8
r172 42 95 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=3.275 $Y=1.8
+ $X2=3.37 $Y2=1.8
r173 42 43 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.275 $Y=1.8
+ $X2=2.605 $Y2=1.8
r174 38 40 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.51 $Y=1.98
+ $X2=2.51 $Y2=2.91
r175 36 94 2.34704 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=2.51 $Y=1.925
+ $X2=2.51 $Y2=1.8
r176 36 38 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=2.51 $Y=1.925
+ $X2=2.51 $Y2=1.98
r177 34 94 4.08801 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=2.415 $Y=1.8
+ $X2=2.51 $Y2=1.8
r178 34 35 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.415 $Y=1.8
+ $X2=1.745 $Y2=1.8
r179 30 32 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=1.615 $Y=1.98
+ $X2=1.615 $Y2=2.91
r180 28 35 6.8199 $w=2.5e-07 $l=1.82071e-07 $layer=LI1_cond $X=1.615 $Y=1.925
+ $X2=1.745 $Y2=1.8
r181 28 30 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=1.615 $Y=1.925
+ $X2=1.615 $Y2=1.98
r182 9 103 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.39
+ $Y=1.835 $X2=8.53 $Y2=2.91
r183 9 92 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=8.39
+ $Y=1.835 $X2=8.53 $Y2=1.99
r184 8 87 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=7.53
+ $Y=1.835 $X2=7.67 $Y2=2.9
r185 8 84 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=7.53
+ $Y=1.835 $X2=7.67 $Y2=2.22
r186 7 79 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=6.67
+ $Y=1.835 $X2=6.81 $Y2=2.9
r187 7 76 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=6.67
+ $Y=1.835 $X2=6.81 $Y2=2.22
r188 6 71 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=1.835 $X2=5.95 $Y2=2.9
r189 6 68 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=1.835 $X2=5.95 $Y2=2.22
r190 5 98 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.835 $X2=5.09 $Y2=2.91
r191 5 63 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.835 $X2=5.09 $Y2=1.98
r192 4 56 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.09
+ $Y=1.835 $X2=4.23 $Y2=2.91
r193 4 54 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.09
+ $Y=1.835 $X2=4.23 $Y2=1.98
r194 3 48 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.835 $X2=3.37 $Y2=2.91
r195 3 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.835 $X2=3.37 $Y2=1.98
r196 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.835 $X2=2.51 $Y2=2.91
r197 2 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.835 $X2=2.51 $Y2=1.98
r198 1 32 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.835 $X2=1.65 $Y2=2.91
r199 1 30 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.835 $X2=1.65 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_8%Z 1 2 3 4 5 6 7 8 31 33 34 37 41 45 49 53 55
+ 56 57 58 59 60 79
c85 34 0 1.19405e-19 $X=5.685 $Y=1.78
r86 59 79 2.97561 $w=7.38e-07 $l=1.8e-07 $layer=LI1_cond $X=7.92 $Y=1.282
+ $X2=8.1 $Y2=1.282
r87 59 60 9.67097 $w=1.7e-07 $l=3.83e-07 $layer=LI1_cond $X=7.92 $Y=1.282
+ $X2=7.92 $Y2=1.665
r88 57 59 7.93496 $w=7.38e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.282
+ $X2=7.92 $Y2=1.282
r89 57 58 9.67097 $w=1.7e-07 $l=3.83e-07 $layer=LI1_cond $X=7.44 $Y=1.282
+ $X2=7.44 $Y2=1.665
r90 55 56 9.67097 $w=1.7e-07 $l=3.83e-07 $layer=LI1_cond $X=6.96 $Y=1.282
+ $X2=6.96 $Y2=1.665
r91 55 68 9.58808 $w=7.38e-07 $l=5.8e-07 $layer=LI1_cond $X=6.96 $Y=1.282
+ $X2=6.38 $Y2=1.282
r92 51 79 0.247967 $w=7.38e-07 $l=1.5e-08 $layer=LI1_cond $X=8.115 $Y=1.282
+ $X2=8.1 $Y2=1.282
r93 51 53 19.9058 $w=2.18e-07 $l=3.8e-07 $layer=LI1_cond $X=8.115 $Y=1.14
+ $X2=8.115 $Y2=0.76
r94 47 79 5.47063 $w=3.3e-07 $l=5.93e-07 $layer=LI1_cond $X=8.1 $Y=1.875 $X2=8.1
+ $Y2=1.282
r95 47 49 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=8.1 $Y=1.875
+ $X2=8.1 $Y2=1.98
r96 43 57 3.30623 $w=7.38e-07 $l=2e-07 $layer=LI1_cond $X=7.24 $Y=1.282 $X2=7.44
+ $Y2=1.282
r97 43 55 4.62873 $w=7.38e-07 $l=2.8e-07 $layer=LI1_cond $X=7.24 $Y=1.282
+ $X2=6.96 $Y2=1.282
r98 43 45 22.1818 $w=1.88e-07 $l=3.8e-07 $layer=LI1_cond $X=7.24 $Y=1.14
+ $X2=7.24 $Y2=0.76
r99 39 43 5.47063 $w=3.3e-07 $l=5.93e-07 $layer=LI1_cond $X=7.24 $Y=1.875
+ $X2=7.24 $Y2=1.282
r100 39 41 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.24 $Y=1.875
+ $X2=7.24 $Y2=1.98
r101 35 68 5.47063 $w=3.3e-07 $l=5.93e-07 $layer=LI1_cond $X=6.38 $Y=1.875
+ $X2=6.38 $Y2=1.282
r102 35 37 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=6.38 $Y=1.875
+ $X2=6.38 $Y2=1.98
r103 33 68 5.12165 $w=7.38e-07 $l=4.65994e-07 $layer=LI1_cond $X=6.305 $Y=0.852
+ $X2=6.38 $Y2=1.282
r104 33 34 30.9378 $w=1.88e-07 $l=5.3e-07 $layer=LI1_cond $X=6.215 $Y=1.78
+ $X2=5.685 $Y2=1.78
r105 29 34 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=5.52 $Y=1.875
+ $X2=5.685 $Y2=1.78
r106 29 31 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=5.52 $Y=1.875
+ $X2=5.52 $Y2=1.98
r107 27 33 27.8359 $w=3.23e-07 $l=7.85e-07 $layer=LI1_cond $X=5.52 $Y=0.852
+ $X2=6.305 $Y2=0.852
r108 8 49 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.96
+ $Y=1.835 $X2=8.1 $Y2=1.98
r109 7 41 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.1
+ $Y=1.835 $X2=7.24 $Y2=1.98
r110 6 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.24
+ $Y=1.835 $X2=6.38 $Y2=1.98
r111 5 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=5.38
+ $Y=1.835 $X2=5.52 $Y2=1.98
r112 4 53 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=7.96
+ $Y=0.235 $X2=8.1 $Y2=0.76
r113 3 45 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=7.1
+ $Y=0.235 $X2=7.24 $Y2=0.76
r114 2 68 182 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_NDIFF $count=1 $X=6.24
+ $Y=0.235 $X2=6.38 $Y2=0.855
r115 1 27 182 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_NDIFF $count=1 $X=5.38
+ $Y=0.235 $X2=5.52 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_8%VGND 1 2 3 4 5 16 18 22 26 30 32 36 39 40 42
+ 43 44 45 46 66 67 73
r117 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r118 66 67 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r119 64 67 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=8.88
+ $Y2=0
r120 63 66 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=8.88
+ $Y2=0
r121 63 64 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r122 61 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.79 $Y=0 $X2=4.66
+ $Y2=0
r123 61 63 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.79 $Y=0 $X2=5.04
+ $Y2=0
r124 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r125 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r126 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r127 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r128 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r129 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r130 51 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r131 50 53 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r132 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r133 48 70 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r134 48 50 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.72
+ $Y2=0
r135 46 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r136 46 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r137 46 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r138 44 59 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.6
+ $Y2=0
r139 44 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.8
+ $Y2=0
r140 42 56 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.64
+ $Y2=0
r141 42 43 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.81 $Y=0 $X2=2.94
+ $Y2=0
r142 41 59 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=3.6
+ $Y2=0
r143 41 43 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=2.94
+ $Y2=0
r144 39 53 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=1.68
+ $Y2=0
r145 39 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=2.08
+ $Y2=0
r146 38 56 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.64
+ $Y2=0
r147 38 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.08
+ $Y2=0
r148 34 73 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.66 $Y2=0
r149 34 36 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=4.66 $Y=0.085
+ $X2=4.66 $Y2=0.38
r150 33 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.93 $Y=0 $X2=3.8
+ $Y2=0
r151 32 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.66
+ $Y2=0
r152 32 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=3.93
+ $Y2=0
r153 28 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=0.085
+ $X2=3.8 $Y2=0
r154 28 30 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.8 $Y=0.085
+ $X2=3.8 $Y2=0.38
r155 24 43 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0
r156 24 26 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.94 $Y=0.085
+ $X2=2.94 $Y2=0.38
r157 20 40 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0
r158 20 22 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0.38
r159 16 70 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=0.085
+ $X2=0.195 $Y2=0
r160 16 18 13.4777 $w=2.93e-07 $l=3.45e-07 $layer=LI1_cond $X=0.242 $Y=0.085
+ $X2=0.242 $Y2=0.43
r161 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.52
+ $Y=0.235 $X2=4.66 $Y2=0.38
r162 4 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.66
+ $Y=0.235 $X2=3.8 $Y2=0.38
r163 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.8
+ $Y=0.235 $X2=2.94 $Y2=0.38
r164 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.94
+ $Y=0.235 $X2=2.08 $Y2=0.38
r165 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.285 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_8%A_305_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 52 55 56 62 66 70 72 73 74 78 80
r153 68 70 0.192074 $w=2.98e-07 $l=5e-09 $layer=LI1_cond $X=8.545 $Y=0.425
+ $X2=8.545 $Y2=0.43
r154 67 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.835 $Y=0.34
+ $X2=7.67 $Y2=0.34
r155 66 68 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=8.395 $Y=0.34
+ $X2=8.545 $Y2=0.425
r156 66 67 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.395 $Y=0.34
+ $X2=7.835 $Y2=0.34
r157 63 78 7.19657 $w=2.17e-07 $l=1.87029e-07 $layer=LI1_cond $X=6.975 $Y=0.34
+ $X2=6.81 $Y2=0.387
r158 62 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.505 $Y=0.34
+ $X2=7.67 $Y2=0.34
r159 62 63 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.505 $Y=0.34
+ $X2=6.975 $Y2=0.34
r160 57 76 3.15837 $w=2.65e-07 $l=1.13e-07 $layer=LI1_cond $X=5.185 $Y=0.387
+ $X2=5.072 $Y2=0.387
r161 57 59 33.2686 $w=2.63e-07 $l=7.65e-07 $layer=LI1_cond $X=5.185 $Y=0.387
+ $X2=5.95 $Y2=0.387
r162 56 78 7.19657 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=0.387
+ $X2=6.81 $Y2=0.387
r163 56 59 30.2244 $w=2.63e-07 $l=6.95e-07 $layer=LI1_cond $X=6.645 $Y=0.387
+ $X2=5.95 $Y2=0.387
r164 53 55 17.1586 $w=2.23e-07 $l=3.35e-07 $layer=LI1_cond $X=5.072 $Y=1.285
+ $X2=5.072 $Y2=0.95
r165 52 76 3.71737 $w=2.25e-07 $l=1.33e-07 $layer=LI1_cond $X=5.072 $Y=0.52
+ $X2=5.072 $Y2=0.387
r166 52 55 22.0245 $w=2.23e-07 $l=4.3e-07 $layer=LI1_cond $X=5.072 $Y=0.52
+ $X2=5.072 $Y2=0.95
r167 51 74 5.92271 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=4.36 $Y=1.395
+ $X2=4.23 $Y2=1.395
r168 50 53 6.81761 $w=2.2e-07 $l=1.57683e-07 $layer=LI1_cond $X=4.96 $Y=1.395
+ $X2=5.072 $Y2=1.285
r169 50 51 31.4303 $w=2.18e-07 $l=6e-07 $layer=LI1_cond $X=4.96 $Y=1.395
+ $X2=4.36 $Y2=1.395
r170 46 74 0.748496 $w=2.6e-07 $l=1.1e-07 $layer=LI1_cond $X=4.23 $Y=1.285
+ $X2=4.23 $Y2=1.395
r171 46 48 38.3409 $w=2.58e-07 $l=8.65e-07 $layer=LI1_cond $X=4.23 $Y=1.285
+ $X2=4.23 $Y2=0.42
r172 45 73 5.92271 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=3.5 $Y=1.395
+ $X2=3.37 $Y2=1.395
r173 44 74 5.92271 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=4.1 $Y=1.395
+ $X2=4.23 $Y2=1.395
r174 44 45 31.4303 $w=2.18e-07 $l=6e-07 $layer=LI1_cond $X=4.1 $Y=1.395 $X2=3.5
+ $Y2=1.395
r175 40 73 0.748496 $w=2.6e-07 $l=1.1e-07 $layer=LI1_cond $X=3.37 $Y=1.285
+ $X2=3.37 $Y2=1.395
r176 40 42 38.3409 $w=2.58e-07 $l=8.65e-07 $layer=LI1_cond $X=3.37 $Y=1.285
+ $X2=3.37 $Y2=0.42
r177 39 72 5.92271 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=1.395
+ $X2=2.51 $Y2=1.395
r178 38 73 5.92271 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=3.24 $Y=1.395
+ $X2=3.37 $Y2=1.395
r179 38 39 31.4303 $w=2.18e-07 $l=6e-07 $layer=LI1_cond $X=3.24 $Y=1.395
+ $X2=2.64 $Y2=1.395
r180 34 72 0.748496 $w=2.6e-07 $l=1.1e-07 $layer=LI1_cond $X=2.51 $Y=1.285
+ $X2=2.51 $Y2=1.395
r181 34 36 38.3409 $w=2.58e-07 $l=8.65e-07 $layer=LI1_cond $X=2.51 $Y=1.285
+ $X2=2.51 $Y2=0.42
r182 32 72 5.92271 $w=2.2e-07 $l=1.3e-07 $layer=LI1_cond $X=2.38 $Y=1.395
+ $X2=2.51 $Y2=1.395
r183 32 33 31.4303 $w=2.18e-07 $l=6e-07 $layer=LI1_cond $X=2.38 $Y=1.395
+ $X2=1.78 $Y2=1.395
r184 28 33 7.00622 $w=2.2e-07 $l=1.95407e-07 $layer=LI1_cond $X=1.632 $Y=1.285
+ $X2=1.78 $Y2=1.395
r185 28 30 33.792 $w=2.93e-07 $l=8.65e-07 $layer=LI1_cond $X=1.632 $Y=1.285
+ $X2=1.632 $Y2=0.42
r186 9 70 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=8.39
+ $Y=0.235 $X2=8.53 $Y2=0.43
r187 8 80 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=7.53
+ $Y=0.235 $X2=7.67 $Y2=0.395
r188 7 78 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=6.67
+ $Y=0.235 $X2=6.81 $Y2=0.385
r189 6 59 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=5.81
+ $Y=0.235 $X2=5.95 $Y2=0.42
r190 5 76 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.95
+ $Y=0.235 $X2=5.09 $Y2=0.42
r191 5 55 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=4.95
+ $Y=0.235 $X2=5.09 $Y2=0.95
r192 4 48 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.09
+ $Y=0.235 $X2=4.23 $Y2=0.42
r193 3 42 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.23
+ $Y=0.235 $X2=3.37 $Y2=0.42
r194 2 36 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.37
+ $Y=0.235 $X2=2.51 $Y2=0.42
r195 1 30 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=1.525
+ $Y=0.235 $X2=1.65 $Y2=0.42
.ends

