* File: sky130_fd_sc_lp__decapkapwr_6.pxi.spice
* Created: Wed Sep  2 09:42:40 2020
* 
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_6%VGND N_VGND_M1001_s N_VGND_c_25_n
+ N_VGND_c_26_n N_VGND_c_27_n N_VGND_c_28_n N_VGND_c_29_n N_VGND_c_30_n
+ N_VGND_c_31_n VGND N_VGND_M1000_g N_VGND_c_32_n N_VGND_c_33_n
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_6%VGND
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_6%KAPWR N_KAPWR_M1000_s N_KAPWR_c_57_n
+ N_KAPWR_c_58_n N_KAPWR_c_67_n N_KAPWR_c_55_n N_KAPWR_c_56_n N_KAPWR_c_61_n
+ N_KAPWR_c_62_n KAPWR N_KAPWR_M1001_g N_KAPWR_c_63_n
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_6%KAPWR
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_6%VPWR VPWR N_VPWR_c_91_n VPWR
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_6%VPWR
cc_1 VNB N_VGND_c_25_n 0.012758f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.085
cc_2 VNB N_VGND_c_26_n 0.0651019f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.38
cc_3 VNB N_VGND_c_27_n 0.00211035f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.77
cc_4 VNB N_VGND_c_28_n 4.97259e-19 $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.77
cc_5 VNB N_VGND_c_29_n 0.0193278f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.77
cc_6 VNB N_VGND_c_30_n 0.0105251f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.085
cc_7 VNB N_VGND_c_31_n 0.0400716f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.405
cc_8 VNB N_VGND_c_32_n 0.0598957f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=0
cc_9 VNB N_VGND_c_33_n 0.170588f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0
cc_10 VNB N_KAPWR_c_55_n 0.016303f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.77
cc_11 VNB N_KAPWR_c_56_n 0.216628f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.77
cc_12 VNB VPWR 0.123877f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=0.235
cc_13 VPB N_VGND_c_27_n 0.0140672f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.77
cc_14 VPB N_VGND_c_28_n 0.00874558f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.77
cc_15 VPB N_VGND_c_29_n 0.222599f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.77
cc_16 VPB N_KAPWR_c_57_n 0.00922717f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.085
cc_17 VPB N_KAPWR_c_58_n 0.023615f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.38
cc_18 VPB N_KAPWR_c_55_n 8.77427e-19 $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.77
cc_19 VPB N_KAPWR_c_56_n 0.0211573f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.77
cc_20 VPB N_KAPWR_c_61_n 0.00961815f $X=-0.19 $Y=1.655 $X2=2.615 $Y2=1.085
cc_21 VPB N_KAPWR_c_62_n 0.0486658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_KAPWR_c_63_n 0.0254524f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=0
cc_23 VPB VPWR 0.0430575f $X=-0.19 $Y=1.655 $X2=0.21 $Y2=0.235
cc_24 VPB N_VPWR_c_91_n 0.0756674f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=1.605
cc_25 N_VGND_c_29_n N_KAPWR_c_57_n 0.00685959f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_26 N_VGND_c_27_n N_KAPWR_c_58_n 0.0205458f $X=0.5 $Y=1.77 $X2=0 $Y2=0
cc_27 N_VGND_c_29_n N_KAPWR_c_58_n 0.0280564f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_28 N_VGND_c_29_n N_KAPWR_c_67_n 0.117197f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_29 N_VGND_c_28_n N_KAPWR_c_55_n 0.0024823f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_30 N_VGND_c_29_n N_KAPWR_c_55_n 0.0064509f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_31 N_VGND_c_31_n N_KAPWR_c_55_n 0.0246728f $X=2.615 $Y=0.405 $X2=0 $Y2=0
cc_32 N_VGND_c_26_n N_KAPWR_c_56_n 0.0654854f $X=0.335 $Y=0.38 $X2=0 $Y2=0
cc_33 N_VGND_c_28_n N_KAPWR_c_56_n 0.00473507f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_34 N_VGND_c_29_n N_KAPWR_c_56_n 0.127834f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_35 N_VGND_c_31_n N_KAPWR_c_56_n 0.0532165f $X=2.615 $Y=0.405 $X2=0 $Y2=0
cc_36 N_VGND_c_32_n N_KAPWR_c_56_n 0.0760645f $X=2.45 $Y=0 $X2=0 $Y2=0
cc_37 N_VGND_c_33_n N_KAPWR_c_56_n 0.120027f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_38 N_VGND_c_29_n N_KAPWR_c_61_n 0.00738552f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_39 N_VGND_c_29_n N_KAPWR_c_62_n 0.0443938f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_40 N_VGND_c_29_n N_KAPWR_c_63_n 0.0972887f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_41 N_VGND_c_29_n VPWR 0.0458048f $X=0.915 $Y=1.77 $X2=-0.19 $Y2=-0.245
cc_42 N_VGND_c_29_n N_VPWR_c_91_n 0.0524183f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_43 N_KAPWR_M1000_s VPWR 0.00234386f $X=0.135 $Y=2.095 $X2=-0.19 $Y2=-0.245
cc_44 N_KAPWR_c_57_n VPWR 0.00306712f $X=0.26 $Y=2.675 $X2=-0.19 $Y2=-0.245
cc_45 N_KAPWR_c_67_n VPWR 0.0106097f $X=2.385 $Y=2.81 $X2=-0.19 $Y2=-0.245
cc_46 N_KAPWR_c_61_n VPWR 0.00338053f $X=2.567 $Y=2.675 $X2=-0.19 $Y2=-0.245
cc_47 N_KAPWR_c_63_n VPWR 0.290153f $X=2.665 $Y=2.81 $X2=-0.19 $Y2=-0.245
cc_48 N_KAPWR_c_57_n N_VPWR_c_91_n 0.0212079f $X=0.26 $Y=2.675 $X2=0 $Y2=0
cc_49 N_KAPWR_c_67_n N_VPWR_c_91_n 0.0690021f $X=2.385 $Y=2.81 $X2=0 $Y2=0
cc_50 N_KAPWR_c_61_n N_VPWR_c_91_n 0.0236354f $X=2.567 $Y=2.675 $X2=0 $Y2=0
cc_51 N_KAPWR_c_63_n N_VPWR_c_91_n 0.00579034f $X=2.665 $Y=2.81 $X2=0 $Y2=0
