* File: sky130_fd_sc_lp__sdfxtp_1.spice
* Created: Fri Aug 28 11:30:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfxtp_1.pex.spice"
.subckt sky130_fd_sc_lp__sdfxtp_1  VNB VPB D SCE SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* SCE	SCE
* D	D
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_SCE_M1017_g N_A_78_123#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1010 A_247_123# N_A_78_123#_M1010_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1006 N_A_319_123#_M1006_d N_D_M1006_g A_247_123# VNB NSHORT L=0.15 W=0.42
+ AD=0.12075 AS=0.0441 PD=0.995 PS=0.63 NRD=84.276 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1031 A_464_123# N_SCE_M1031_g N_A_319_123#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.12075 PD=0.63 PS=0.995 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_SCD_M1016_g A_464_123# VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.0441 PD=0.73 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_628_123#_M1009_d N_CLK_M1009_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0651 PD=1.37 PS=0.73 NRD=0 NRS=8.568 M=1 R=2.8
+ SA=75002.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_823_47#_M1004_d N_A_628_123#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_1051_125#_M1018_d N_A_628_123#_M1018_g N_A_319_123#_M1018_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1012 A_1137_125# N_A_823_47#_M1012_g N_A_1051_125#_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_A_1201_99#_M1030_g A_1137_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.15017 AS=0.0672 PD=1.00642 PS=0.74 NRD=28.56 NRS=30 M=1 R=2.8 SA=75001.1
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_1201_99#_M1003_d N_A_1051_125#_M1003_g N_VGND_M1030_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.179079 AS=0.22883 PD=1.43698 PS=1.53358 NRD=15.936
+ NRS=47.808 M=1 R=4.26667 SA=75001.4 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1014 N_A_1459_449#_M1014_d N_A_823_47#_M1014_g N_A_1201_99#_M1003_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.12915 AS=0.117521 PD=1.035 PS=0.943019 NRD=95.712
+ NRS=64.224 M=1 R=2.8 SA=75001.3 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1025 A_1664_65# N_A_628_123#_M1025_g N_A_1459_449#_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.12915 PD=0.63 PS=1.035 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_1657_383#_M1026_g A_1664_65# VNB NSHORT L=0.15 W=0.42
+ AD=0.0855057 AS=0.0441 PD=0.80434 PS=0.63 NRD=27.852 NRS=14.28 M=1 R=2.8
+ SA=75002.4 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_A_1657_383#_M1000_d N_A_1459_449#_M1000_g N_VGND_M1026_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.130294 PD=1.81 PS=1.22566 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75002 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1019 N_Q_M1019_d N_A_1657_383#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1020 N_VPWR_M1020_d N_SCE_M1020_g N_A_78_123#_M1020_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1152 AS=0.1696 PD=1 PS=1.81 NRD=10.7562 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1023 A_283_491# N_SCE_M1023_g N_VPWR_M1020_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1152 PD=0.85 PS=1 NRD=15.3857 NRS=13.8491 M=1 R=4.26667
+ SA=75000.7 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1028 N_A_319_123#_M1028_d N_D_M1028_g A_283_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.1
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1011 A_441_491# N_A_78_123#_M1011_g N_A_319_123#_M1028_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=32.308 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_SCD_M1007_g A_441_491# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1008 AS=0.1024 PD=0.955 PS=0.96 NRD=7.683 NRS=32.308 M=1 R=4.26667
+ SA=75002 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1027 N_A_628_123#_M1027_d N_CLK_M1027_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1008 PD=1.81 PS=0.955 NRD=0 NRS=3.0732 M=1 R=4.26667
+ SA=75002.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_A_823_47#_M1024_d N_A_628_123#_M1024_g N_VPWR_M1024_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.32 AS=0.192 PD=2.28 PS=1.88 NRD=72.3187 NRS=10.7562 M=1
+ R=4.26667 SA=75000.2 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1002 N_A_1051_125#_M1002_d N_A_823_47#_M1002_g N_A_319_123#_M1002_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1029 A_1157_449# N_A_628_123#_M1029_g N_A_1051_125#_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0462 AS=0.0588 PD=0.64 PS=0.7 NRD=25.7873 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1015 N_VPWR_M1015_d N_A_1201_99#_M1015_g A_1157_449# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.140133 AS=0.0462 PD=1.00667 PS=0.64 NRD=130.69 NRS=25.7873 M=1 R=2.8
+ SA=75001 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_1201_99#_M1013_d N_A_1051_125#_M1013_g N_VPWR_M1015_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.280267 PD=1.12 PS=2.01333 NRD=0 NRS=19.9167 M=1
+ R=5.6 SA=75001 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1008 N_A_1459_449#_M1008_d N_A_628_123#_M1008_g N_A_1201_99#_M1013_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2464 AS=0.1176 PD=1.96 PS=1.12 NRD=79.7259 NRS=0
+ M=1 R=5.6 SA=75001.4 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1021 A_1615_495# N_A_823_47#_M1021_g N_A_1459_449#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0756 AS=0.1232 PD=0.78 PS=0.98 NRD=58.6272 NRS=4.6886 M=1 R=2.8
+ SA=75002.1 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1022_d N_A_1657_383#_M1022_g A_1615_495# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1064 AS=0.0756 PD=0.876667 PS=0.78 NRD=92.6294 NRS=58.6272 M=1
+ R=2.8 SA=75002.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_A_1657_383#_M1001_d N_A_1459_449#_M1001_g N_VPWR_M1022_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.2128 PD=2.21 PS=1.75333 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_Q_M1005_d N_A_1657_383#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=20.4031 P=25.61
c_218 VPB 0 6.83332e-20 $X=0 $Y=3.085
c_1519 A_1157_449# 0 6.8524e-20 $X=5.785 $Y=2.245
*
.include "sky130_fd_sc_lp__sdfxtp_1.pxi.spice"
*
.ends
*
*
