* NGSPICE file created from sky130_fd_sc_lp__or4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
M1000 a_276_47# A VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=1.0133e+12p ps=8.83e+06u
M1001 VGND a_462_351# a_276_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_276_403# A VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.316e+11p ps=7.72e+06u
M1003 VGND C_N a_40_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 a_348_403# B a_276_403# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 X a_276_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1006 VGND B a_276_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR C_N a_40_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 VGND a_276_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 a_462_351# D_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1010 a_276_47# a_40_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_462_351# D_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1012 a_420_403# a_40_47# a_348_403# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1013 VPWR a_276_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_276_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_276_47# a_462_351# a_420_403# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

