* File: sky130_fd_sc_lp__o21a_m.pex.spice
* Created: Wed Sep  2 10:15:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21A_M%A_80_23# 1 2 9 11 13 16 18 21 23 24 25 27 28
+ 31 34 37 41 44
r75 38 41 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.33 $Y=2.82 $X2=1.41
+ $Y2=2.82
r76 37 44 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=0.94
+ $X2=0.577 $Y2=0.775
r77 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=0.94 $X2=0.59 $Y2=0.94
r78 34 38 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.33 $Y=2.715
+ $X2=1.33 $Y2=2.82
r79 33 34 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.33 $Y=2.47
+ $X2=1.33 $Y2=2.715
r80 29 31 6.8658 $w=2.08e-07 $l=1.3e-07 $layer=LI1_cond $X=1.21 $Y=0.775
+ $X2=1.21 $Y2=0.645
r81 27 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.245 $Y=2.385
+ $X2=1.33 $Y2=2.47
r82 27 28 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.245 $Y=2.385
+ $X2=0.675 $Y2=2.385
r83 26 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=0.86
+ $X2=0.59 $Y2=0.86
r84 25 29 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.105 $Y=0.86
+ $X2=1.21 $Y2=0.775
r85 25 26 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.105 $Y=0.86
+ $X2=0.675 $Y2=0.86
r86 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.59 $Y=2.3
+ $X2=0.675 $Y2=2.385
r87 23 36 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.59 $Y=0.945
+ $X2=0.59 $Y2=0.86
r88 23 24 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=0.59 $Y=0.945
+ $X2=0.59 $Y2=2.3
r89 19 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.475 $Y=2.195
+ $X2=0.765 $Y2=2.195
r90 14 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.765 $Y=2.27
+ $X2=0.765 $Y2=2.195
r91 14 16 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.765 $Y=2.27
+ $X2=0.765 $Y2=2.885
r92 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.12
+ $X2=0.475 $Y2=2.195
r93 13 18 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.475 $Y=2.12
+ $X2=0.475 $Y2=1.445
r94 11 18 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.577 $Y=1.268
+ $X2=0.577 $Y2=1.445
r95 10 37 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.577 $Y=0.952
+ $X2=0.577 $Y2=0.94
r96 10 11 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.577 $Y=0.952
+ $X2=0.577 $Y2=1.268
r97 9 44 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.455
+ $X2=0.475 $Y2=0.775
r98 2 41 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.27
+ $Y=2.675 $X2=1.41 $Y2=2.82
r99 1 31 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.37 $X2=1.21 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_M%B1 3 7 12 13 14 15 16 21
c49 3 0 1.78534e-19 $X=1.195 $Y=2.885
r50 15 16 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.172 $Y=1.665
+ $X2=1.172 $Y2=2.035
r51 14 15 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.172 $Y=1.295
+ $X2=1.172 $Y2=1.665
r52 14 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.145
+ $Y=1.375 $X2=1.145 $Y2=1.375
r53 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.145 $Y=1.715
+ $X2=1.145 $Y2=1.375
r54 12 13 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.715
+ $X2=1.145 $Y2=1.88
r55 5 21 64.8846 $w=2.08e-07 $l=4.539e-07 $layer=POLY_cond $X=1.425 $Y=1.04
+ $X2=1.145 $Y2=1.375
r56 5 7 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.425 $Y=1.04
+ $X2=1.425 $Y2=0.58
r57 3 13 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.195 $Y=2.885
+ $X2=1.195 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_M%A2 2 5 9 11 12 13 14 15 21
c50 21 0 1.44993e-19 $X=1.715 $Y=1.595
c51 12 0 1.94558e-19 $X=1.68 $Y=1.295
r52 21 23 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.595
+ $X2=1.74 $Y2=1.43
r53 14 15 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=1.697 $Y=2.035
+ $X2=1.697 $Y2=2.405
r54 13 14 23.8049 $w=2.03e-07 $l=4.4e-07 $layer=LI1_cond $X=1.697 $Y=1.595
+ $X2=1.697 $Y2=2.035
r55 13 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.715
+ $Y=1.595 $X2=1.715 $Y2=1.595
r56 12 13 16.2306 $w=2.03e-07 $l=3e-07 $layer=LI1_cond $X=1.697 $Y=1.295
+ $X2=1.697 $Y2=1.595
r57 9 23 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.855 $Y=0.58
+ $X2=1.855 $Y2=1.43
r58 5 11 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.625 $Y=2.885
+ $X2=1.625 $Y2=2.1
r59 2 11 48.9106 $w=3.8e-07 $l=1.9e-07 $layer=POLY_cond $X=1.74 $Y=1.91 $X2=1.74
+ $Y2=2.1
r60 1 21 3.65891 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.74 $Y=1.62 $X2=1.74
+ $Y2=1.595
r61 1 2 42.4433 $w=3.8e-07 $l=2.9e-07 $layer=POLY_cond $X=1.74 $Y=1.62 $X2=1.74
+ $Y2=1.91
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_M%A1 3 6 9 13 17 18 19 20 21 22 28
c37 9 0 1.94558e-19 $X=2.285 $Y=0.58
r38 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.335
+ $Y=1.595 $X2=2.335 $Y2=1.595
r39 21 22 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.247 $Y=2.035
+ $X2=2.247 $Y2=2.405
r40 20 21 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.247 $Y=1.665
+ $X2=2.247 $Y2=2.035
r41 20 29 2.33829 $w=3.43e-07 $l=7e-08 $layer=LI1_cond $X=2.247 $Y=1.665
+ $X2=2.247 $Y2=1.595
r42 19 29 10.0212 $w=3.43e-07 $l=3e-07 $layer=LI1_cond $X=2.247 $Y=1.295
+ $X2=2.247 $Y2=1.595
r43 17 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.335 $Y=1.935
+ $X2=2.335 $Y2=1.595
r44 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.935
+ $X2=2.335 $Y2=2.1
r45 16 28 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.43
+ $X2=2.335 $Y2=1.595
r46 11 13 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.985 $Y=2.415
+ $X2=2.245 $Y2=2.415
r47 9 16 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=2.285 $Y=0.58
+ $X2=2.285 $Y2=1.43
r48 6 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.245 $Y=2.34
+ $X2=2.245 $Y2=2.415
r49 6 18 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.245 $Y=2.34
+ $X2=2.245 $Y2=2.1
r50 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.985 $Y=2.49
+ $X2=1.985 $Y2=2.415
r51 1 3 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.985 $Y=2.49
+ $X2=1.985 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_M%X 1 2 9 12 13 14 15 16 24 36
c22 36 0 1.78534e-19 $X=0.55 $Y=2.82
r23 16 24 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.24 $Y=2.82
+ $X2=0.24 $Y2=2.715
r24 16 36 9.21118 $w=3.53e-07 $l=2.25e-07 $layer=LI1_cond $X=0.325 $Y=2.82
+ $X2=0.55 $Y2=2.82
r25 16 24 0.848128 $w=1.68e-07 $l=1.3e-08 $layer=LI1_cond $X=0.24 $Y=2.702
+ $X2=0.24 $Y2=2.715
r26 15 16 19.3765 $w=1.68e-07 $l=2.97e-07 $layer=LI1_cond $X=0.24 $Y=2.405
+ $X2=0.24 $Y2=2.702
r27 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.405
r28 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r29 12 13 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r30 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.24 $Y=0.595 $X2=0.24
+ $Y2=1.295
r31 9 11 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=0.43
+ $X2=0.26 $Y2=0.595
r32 2 36 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.425
+ $Y=2.675 $X2=0.55 $Y2=2.82
r33 1 9 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.245 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_M%VPWR 1 2 9 13 16 17 18 24 30 31 34
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.2 $Y2=3.33
r41 28 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.2 $Y2=3.33
r45 24 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 18 22 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 16 21 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.98 $Y2=3.33
r51 15 26 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.98 $Y2=3.33
r53 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=3.245 $X2=2.2
+ $Y2=3.33
r54 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.2 $Y=3.245
+ $X2=2.2 $Y2=2.95
r55 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.98 $Y=3.245 $X2=0.98
+ $Y2=3.33
r56 7 9 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.98 $Y=3.245 $X2=0.98
+ $Y2=2.95
r57 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.06
+ $Y=2.675 $X2=2.2 $Y2=2.95
r58 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.84
+ $Y=2.675 $X2=0.98 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_M%VGND 1 2 9 13 16 17 18 20 30 31 34
r38 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r41 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r42 25 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.69
+ $Y2=0
r43 25 27 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.68
+ $Y2=0
r44 23 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r45 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 20 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.69
+ $Y2=0
r47 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r48 18 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r49 18 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r50 16 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=1.68
+ $Y2=0
r51 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=2.07
+ $Y2=0
r52 15 30 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.64
+ $Y2=0
r53 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.07
+ $Y2=0
r54 11 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0.085
+ $X2=2.07 $Y2=0
r55 11 13 22.71 $w=2.08e-07 $l=4.3e-07 $layer=LI1_cond $X=2.07 $Y=0.085 $X2=2.07
+ $Y2=0.515
r56 7 34 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r57 7 9 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.39
r58 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.37 $X2=2.07 $Y2=0.515
r59 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.245 $X2=0.69 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O21A_M%A_300_74# 1 2 9 11 12 15
c23 11 0 1.44993e-19 $X=2.395 $Y=0.945
r24 13 15 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.5 $Y=0.86 $X2=2.5
+ $Y2=0.645
r25 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.395 $Y=0.945
+ $X2=2.5 $Y2=0.86
r26 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.395 $Y=0.945
+ $X2=1.745 $Y2=0.945
r27 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.64 $Y=0.86
+ $X2=1.745 $Y2=0.945
r28 7 9 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.64 $Y=0.86 $X2=1.64
+ $Y2=0.645
r29 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.37 $X2=2.5 $Y2=0.645
r30 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.645
.ends

