* File: sky130_fd_sc_lp__o41a_2.spice
* Created: Wed Sep  2 10:27:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41a_2.pex.spice"
.subckt sky130_fd_sc_lp__o41a_2  VNB VPB B1 A4 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_102_53#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A_102_53#_M1011_g N_X_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_465_49#_M1004_d N_B1_M1004_g N_A_102_53#_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1365 AS=0.2226 PD=1.165 PS=2.21 NRD=6.42 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75002.2 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_A4_M1010_g N_A_465_49#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1617 AS=0.1365 PD=1.225 PS=1.165 NRD=7.848 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1006 N_A_465_49#_M1006_d N_A3_M1006_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1617 PD=1.12 PS=1.225 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001.2
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A2_M1012_g N_A_465_49#_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1176 PD=1.23 PS=1.12 NRD=8.568 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1002 N_A_465_49#_M1002_d N_A1_M1002_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=7.14 M=1 R=5.6 SA=75002.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_102_53#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.8 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A_102_53#_M1013_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.53865 AS=0.1764 PD=2.115 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1007 N_A_102_53#_M1007_d N_B1_M1007_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.53865 PD=1.88 PS=2.115 NRD=0 NRS=29.9637 M=1 R=8.4 SA=75001.6
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1008 A_573_367# N_A4_M1008_g N_A_102_53#_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3906 PD=1.47 PS=1.88 NRD=7.8012 NRS=17.7103 M=1 R=8.4
+ SA=75002.4 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1009 A_645_367# N_A3_M1009_g A_573_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75002.8
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1001 A_753_367# N_A2_M1001_g A_645_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.2457 PD=1.65 PS=1.65 NRD=21.8867 NRS=21.8867 M=1 R=8.4 SA=75003.3
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g A_753_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3402 AS=0.2457 PD=3.06 PS=1.65 NRD=0.7683 NRS=21.8867 M=1 R=8.4
+ SA=75003.8 SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
c_73 VPB 0 1.52271e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o41a_2.pxi.spice"
*
.ends
*
*
