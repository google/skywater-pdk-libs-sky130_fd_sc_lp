* File: sky130_fd_sc_lp__a21bo_4.pxi.spice
* Created: Wed Sep  2 09:18:53 2020
* 
x_PM_SKY130_FD_SC_LP__A21BO_4%B1_N N_B1_N_M1013_g N_B1_N_M1021_g B1_N B1_N
+ N_B1_N_c_116_n PM_SKY130_FD_SC_LP__A21BO_4%B1_N
x_PM_SKY130_FD_SC_LP__A21BO_4%A_188_315# N_A_188_315#_M1005_d
+ N_A_188_315#_M1012_d N_A_188_315#_M1004_d N_A_188_315#_c_163_n
+ N_A_188_315#_M1000_g N_A_188_315#_c_149_n N_A_188_315#_c_150_n
+ N_A_188_315#_M1001_g N_A_188_315#_c_166_n N_A_188_315#_M1003_g
+ N_A_188_315#_M1011_g N_A_188_315#_M1009_g N_A_188_315#_M1018_g
+ N_A_188_315#_M1016_g N_A_188_315#_M1019_g N_A_188_315#_c_157_n
+ N_A_188_315#_c_158_n N_A_188_315#_c_159_n N_A_188_315#_c_160_n
+ N_A_188_315#_c_248_p N_A_188_315#_c_161_n N_A_188_315#_c_274_p
+ N_A_188_315#_c_162_n N_A_188_315#_c_292_p N_A_188_315#_c_181_p
+ PM_SKY130_FD_SC_LP__A21BO_4%A_188_315#
x_PM_SKY130_FD_SC_LP__A21BO_4%A_42_47# N_A_42_47#_M1013_s N_A_42_47#_M1021_s
+ N_A_42_47#_M1005_g N_A_42_47#_M1004_g N_A_42_47#_M1020_g N_A_42_47#_M1017_g
+ N_A_42_47#_c_297_n N_A_42_47#_c_298_n N_A_42_47#_c_299_n N_A_42_47#_c_307_n
+ N_A_42_47#_c_308_n N_A_42_47#_c_309_n N_A_42_47#_c_300_n N_A_42_47#_c_301_n
+ N_A_42_47#_c_311_n N_A_42_47#_c_302_n N_A_42_47#_c_313_n N_A_42_47#_c_314_n
+ PM_SKY130_FD_SC_LP__A21BO_4%A_42_47#
x_PM_SKY130_FD_SC_LP__A21BO_4%A2 N_A2_M1008_g N_A2_M1002_g N_A2_M1007_g
+ N_A2_M1010_g N_A2_c_401_n N_A2_c_402_n N_A2_c_403_n N_A2_c_404_n N_A2_c_405_n
+ N_A2_c_406_n A2 A2 A2 PM_SKY130_FD_SC_LP__A21BO_4%A2
x_PM_SKY130_FD_SC_LP__A21BO_4%A1 N_A1_M1012_g N_A1_M1006_g N_A1_M1014_g
+ N_A1_M1015_g A1 N_A1_c_487_n N_A1_c_488_n PM_SKY130_FD_SC_LP__A21BO_4%A1
x_PM_SKY130_FD_SC_LP__A21BO_4%VPWR N_VPWR_M1021_d N_VPWR_M1003_d N_VPWR_M1016_d
+ N_VPWR_M1008_d N_VPWR_M1015_s N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n
+ N_VPWR_c_539_n N_VPWR_c_540_n VPWR N_VPWR_c_541_n N_VPWR_c_542_n
+ N_VPWR_c_543_n N_VPWR_c_544_n N_VPWR_c_545_n N_VPWR_c_546_n N_VPWR_c_535_n
+ N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n
+ PM_SKY130_FD_SC_LP__A21BO_4%VPWR
x_PM_SKY130_FD_SC_LP__A21BO_4%X N_X_M1001_d N_X_M1018_d N_X_M1000_s N_X_M1009_s
+ N_X_c_627_n N_X_c_628_n N_X_c_629_n N_X_c_688_p N_X_c_630_n N_X_c_659_n
+ N_X_c_631_n X X X X X N_X_c_640_n X PM_SKY130_FD_SC_LP__A21BO_4%X
x_PM_SKY130_FD_SC_LP__A21BO_4%A_645_367# N_A_645_367#_M1004_s
+ N_A_645_367#_M1017_s N_A_645_367#_M1006_d N_A_645_367#_M1010_s
+ N_A_645_367#_c_734_n N_A_645_367#_c_702_n N_A_645_367#_c_697_n
+ N_A_645_367#_c_694_n N_A_645_367#_c_714_n N_A_645_367#_c_719_n
+ N_A_645_367#_c_695_n N_A_645_367#_c_727_n N_A_645_367#_c_696_n
+ PM_SKY130_FD_SC_LP__A21BO_4%A_645_367#
x_PM_SKY130_FD_SC_LP__A21BO_4%VGND N_VGND_M1013_d N_VGND_M1011_s N_VGND_M1019_s
+ N_VGND_M1020_s N_VGND_M1007_s N_VGND_c_748_n N_VGND_c_749_n N_VGND_c_750_n
+ N_VGND_c_751_n N_VGND_c_752_n N_VGND_c_753_n N_VGND_c_754_n N_VGND_c_755_n
+ VGND N_VGND_c_756_n N_VGND_c_757_n N_VGND_c_758_n N_VGND_c_759_n
+ N_VGND_c_760_n N_VGND_c_761_n PM_SKY130_FD_SC_LP__A21BO_4%VGND
x_PM_SKY130_FD_SC_LP__A21BO_4%A_908_47# N_A_908_47#_M1002_d N_A_908_47#_M1014_s
+ N_A_908_47#_c_837_n N_A_908_47#_c_840_n N_A_908_47#_c_835_n
+ PM_SKY130_FD_SC_LP__A21BO_4%A_908_47#
cc_1 VNB N_B1_N_M1013_g 0.0234932f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.655
cc_2 VNB N_B1_N_M1021_g 0.00689566f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_3 VNB B1_N 0.00802562f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_B1_N_c_116_n 0.0365322f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.375
cc_5 VNB N_A_188_315#_c_149_n 0.00552439f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.375
cc_6 VNB N_A_188_315#_c_150_n 0.00862475f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.375
cc_7 VNB N_A_188_315#_M1001_g 0.0227508f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.54
cc_8 VNB N_A_188_315#_M1011_g 0.019692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_188_315#_M1009_g 0.00249126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_188_315#_M1018_g 0.0198398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_188_315#_M1016_g 0.00296861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_188_315#_M1019_g 0.0248264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_188_315#_c_157_n 0.00516705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_188_315#_c_158_n 0.0878725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_188_315#_c_159_n 0.00262086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_188_315#_c_160_n 0.00870979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_188_315#_c_161_n 0.00175198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_188_315#_c_162_n 0.0150795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_42_47#_M1005_g 0.0289725f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_A_42_47#_M1020_g 0.0238784f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.54
cc_21 VNB N_A_42_47#_c_297_n 0.0381372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_42_47#_c_298_n 0.0296411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_42_47#_c_299_n 0.0261174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_42_47#_c_300_n 0.00313077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_42_47#_c_301_n 0.0071071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_42_47#_c_302_n 0.0296283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A2_M1008_g 0.00144794f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.655
cc_28 VNB N_A2_M1002_g 0.0225597f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_29 VNB N_A2_M1007_g 0.0346167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A2_c_401_n 3.0309e-19 $X=-0.19 $Y=-0.245 $X2=0.622 $Y2=1.295
cc_31 VNB N_A2_c_402_n 8.23343e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_c_403_n 0.0284647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A2_c_404_n 0.0047115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_c_405_n 0.0204126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_c_406_n 0.0292907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A1_M1012_g 0.0237827f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.655
cc_37 VNB N_A1_M1014_g 0.0247591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A1_c_487_n 9.48006e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A1_c_488_n 0.0333185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_535_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_627_n 0.00655255f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.375
cc_42 VNB N_X_c_628_n 0.00119648f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.375
cc_43 VNB N_X_c_629_n 0.00160619f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.21
cc_44 VNB N_X_c_630_n 0.00516594f $X=-0.19 $Y=-0.245 $X2=0.622 $Y2=1.375
cc_45 VNB N_X_c_631_n 0.00147023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_748_n 0.00183337f $X=-0.19 $Y=-0.245 $X2=0.622 $Y2=1.295
cc_47 VNB N_VGND_c_749_n 3.10897e-19 $X=-0.19 $Y=-0.245 $X2=0.622 $Y2=1.665
cc_48 VNB N_VGND_c_750_n 0.0129657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_751_n 0.00274299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_752_n 0.0109324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_753_n 0.0441559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_754_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_755_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_756_n 0.0170099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_757_n 0.0289278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_758_n 0.036822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_759_n 0.010461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_760_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_761_n 0.308537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_908_47#_c_835_n 0.00278917f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.21
cc_61 VPB N_B1_N_M1021_g 0.0235722f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_62 VPB B1_N 0.00400287f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_63 VPB N_A_188_315#_c_163_n 0.0156976f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_64 VPB N_A_188_315#_c_149_n 0.00250514f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.375
cc_65 VPB N_A_188_315#_c_150_n 0.00248781f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.375
cc_66 VPB N_A_188_315#_c_166_n 0.0156464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_188_315#_M1009_g 0.0192708f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_188_315#_M1016_g 0.0234401f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_188_315#_c_158_n 0.00414427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_42_47#_M1004_g 0.0214827f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.375
cc_71 VPB N_A_42_47#_M1017_g 0.0183672f $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.375
cc_72 VPB N_A_42_47#_c_297_n 0.0166607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_42_47#_c_298_n 0.0067831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_42_47#_c_307_n 0.0111174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_42_47#_c_308_n 0.0180306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_42_47#_c_309_n 0.0116754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_42_47#_c_300_n 6.56038e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_42_47#_c_311_n 0.00790378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_42_47#_c_302_n 0.0128993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_42_47#_c_313_n 0.0322095f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_42_47#_c_314_n 0.00979504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A2_M1008_g 0.0196855f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.655
cc_83 VPB N_A2_M1010_g 0.0256101f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.375
cc_84 VPB N_A2_c_401_n 0.00141571f $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.295
cc_85 VPB N_A2_c_402_n 0.0031284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A2_c_406_n 0.00640735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A1_M1006_g 0.0190578f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_88 VPB N_A1_M1015_g 0.0183785f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.375
cc_89 VPB N_A1_c_487_n 0.00260829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A1_c_488_n 0.00490381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_536_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.295
cc_92 VPB N_VPWR_c_537_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.665
cc_93 VPB N_VPWR_c_538_n 0.00985867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_539_n 0.00218438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_540_n 4.06069e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_541_n 0.0178885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_542_n 0.0147084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_543_n 0.0147084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_544_n 0.0456136f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_545_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_546_n 0.0156941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_535_n 0.0578448f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_548_n 0.0043699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_549_n 0.0043699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_550_n 0.00510963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_551_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_552_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_X_c_627_n 7.28369e-19 $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.375
cc_109 VPB X 0.0160709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_645_367#_c_694_n 0.0035501f $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.375
cc_111 VPB N_A_645_367#_c_695_n 0.02445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_645_367#_c_696_n 0.0305687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 N_B1_N_M1021_g N_A_188_315#_c_150_n 0.0565306f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_114 B1_N N_A_188_315#_c_150_n 0.00143467f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B1_N_M1013_g N_A_188_315#_M1001_g 0.00561591f $X=0.55 $Y=0.655 $X2=0
+ $Y2=0
cc_116 N_B1_N_c_116_n N_A_188_315#_M1001_g 0.00523253f $X=0.535 $Y=1.375 $X2=0
+ $Y2=0
cc_117 N_B1_N_M1021_g N_A_188_315#_c_158_n 4.89192e-19 $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_B1_N_M1021_g N_A_42_47#_c_308_n 0.0112766f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_119 B1_N N_A_42_47#_c_308_n 0.00425075f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B1_N_c_116_n N_A_42_47#_c_301_n 0.00233061f $X=0.535 $Y=1.375 $X2=0
+ $Y2=0
cc_121 B1_N N_A_42_47#_c_311_n 0.00113248f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B1_N_c_116_n N_A_42_47#_c_311_n 0.00255949f $X=0.535 $Y=1.375 $X2=0
+ $Y2=0
cc_123 N_B1_N_M1013_g N_A_42_47#_c_302_n 0.00404367f $X=0.55 $Y=0.655 $X2=0
+ $Y2=0
cc_124 N_B1_N_M1021_g N_A_42_47#_c_302_n 0.00514311f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_125 B1_N N_A_42_47#_c_302_n 0.0435564f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B1_N_c_116_n N_A_42_47#_c_302_n 0.00804797f $X=0.535 $Y=1.375 $X2=0
+ $Y2=0
cc_127 N_B1_N_M1021_g N_VPWR_c_536_n 0.0100126f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_128 N_B1_N_M1021_g N_VPWR_c_541_n 0.00486043f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_129 N_B1_N_M1021_g N_VPWR_c_535_n 0.00545839f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_130 N_B1_N_M1013_g N_X_c_627_n 4.76559e-19 $X=0.55 $Y=0.655 $X2=0 $Y2=0
cc_131 N_B1_N_M1021_g N_X_c_627_n 4.93753e-19 $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_132 B1_N N_X_c_627_n 0.0406448f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_133 N_B1_N_c_116_n N_X_c_627_n 9.89993e-19 $X=0.535 $Y=1.375 $X2=0 $Y2=0
cc_134 N_B1_N_M1013_g N_X_c_629_n 0.00376834f $X=0.55 $Y=0.655 $X2=0 $Y2=0
cc_135 N_B1_N_M1021_g X 7.19541e-19 $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_136 N_B1_N_M1021_g N_X_c_640_n 0.0067709f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_137 B1_N N_X_c_640_n 0.0118622f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_138 N_B1_N_M1013_g N_VGND_c_748_n 0.0131393f $X=0.55 $Y=0.655 $X2=0 $Y2=0
cc_139 B1_N N_VGND_c_748_n 0.00895776f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B1_N_c_116_n N_VGND_c_748_n 2.89261e-19 $X=0.535 $Y=1.375 $X2=0 $Y2=0
cc_141 N_B1_N_M1013_g N_VGND_c_756_n 0.00486043f $X=0.55 $Y=0.655 $X2=0 $Y2=0
cc_142 N_B1_N_M1013_g N_VGND_c_761_n 0.00924348f $X=0.55 $Y=0.655 $X2=0 $Y2=0
cc_143 N_A_188_315#_c_159_n N_A_42_47#_M1005_g 0.00380729f $X=2.735 $Y=1.355
+ $X2=0 $Y2=0
cc_144 N_A_188_315#_c_160_n N_A_42_47#_M1005_g 0.019859f $X=3.615 $Y=1.08 $X2=0
+ $Y2=0
cc_145 N_A_188_315#_c_161_n N_A_42_47#_M1005_g 0.00510287f $X=3.78 $Y=1.97 $X2=0
+ $Y2=0
cc_146 N_A_188_315#_c_161_n N_A_42_47#_M1004_g 0.0156957f $X=3.78 $Y=1.97 $X2=0
+ $Y2=0
cc_147 N_A_188_315#_c_161_n N_A_42_47#_M1020_g 0.00563734f $X=3.78 $Y=1.97 $X2=0
+ $Y2=0
cc_148 N_A_188_315#_c_162_n N_A_42_47#_M1020_g 0.0104133f $X=5.015 $Y=1.08 $X2=0
+ $Y2=0
cc_149 N_A_188_315#_c_181_p N_A_42_47#_M1020_g 0.00541858f $X=3.78 $Y=1.08 $X2=0
+ $Y2=0
cc_150 N_A_188_315#_c_161_n N_A_42_47#_M1017_g 0.0137855f $X=3.78 $Y=1.97 $X2=0
+ $Y2=0
cc_151 N_A_188_315#_M1016_g N_A_42_47#_c_297_n 0.00189802f $X=2.305 $Y=2.465
+ $X2=0 $Y2=0
cc_152 N_A_188_315#_c_157_n N_A_42_47#_c_297_n 0.00144247f $X=2.65 $Y=1.445
+ $X2=0 $Y2=0
cc_153 N_A_188_315#_c_158_n N_A_42_47#_c_297_n 0.017407f $X=2.53 $Y=1.44 $X2=0
+ $Y2=0
cc_154 N_A_188_315#_c_160_n N_A_42_47#_c_297_n 0.00924173f $X=3.615 $Y=1.08
+ $X2=0 $Y2=0
cc_155 N_A_188_315#_c_161_n N_A_42_47#_c_298_n 0.0253617f $X=3.78 $Y=1.97 $X2=0
+ $Y2=0
cc_156 N_A_188_315#_c_162_n N_A_42_47#_c_298_n 0.00164242f $X=5.015 $Y=1.08
+ $X2=0 $Y2=0
cc_157 N_A_188_315#_c_163_n N_A_42_47#_c_308_n 0.0116049f $X=1.015 $Y=1.725
+ $X2=0 $Y2=0
cc_158 N_A_188_315#_c_166_n N_A_42_47#_c_308_n 0.011669f $X=1.445 $Y=1.725 $X2=0
+ $Y2=0
cc_159 N_A_188_315#_M1009_g N_A_42_47#_c_308_n 0.011669f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_188_315#_M1016_g N_A_42_47#_c_308_n 0.0136563f $X=2.305 $Y=2.465
+ $X2=0 $Y2=0
cc_161 N_A_188_315#_M1016_g N_A_42_47#_c_309_n 0.00402661f $X=2.305 $Y=2.465
+ $X2=0 $Y2=0
cc_162 N_A_188_315#_c_161_n N_A_42_47#_c_309_n 0.00532256f $X=3.78 $Y=1.97 $X2=0
+ $Y2=0
cc_163 N_A_188_315#_M1016_g N_A_42_47#_c_300_n 0.001012f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_188_315#_c_157_n N_A_42_47#_c_300_n 0.0151783f $X=2.65 $Y=1.445 $X2=0
+ $Y2=0
cc_165 N_A_188_315#_c_158_n N_A_42_47#_c_300_n 6.13035e-19 $X=2.53 $Y=1.44 $X2=0
+ $Y2=0
cc_166 N_A_188_315#_c_159_n N_A_42_47#_c_300_n 7.13863e-19 $X=2.735 $Y=1.355
+ $X2=0 $Y2=0
cc_167 N_A_188_315#_c_160_n N_A_42_47#_c_300_n 0.0247317f $X=3.615 $Y=1.08 $X2=0
+ $Y2=0
cc_168 N_A_188_315#_c_161_n N_A_42_47#_c_300_n 0.0264895f $X=3.78 $Y=1.97 $X2=0
+ $Y2=0
cc_169 N_A_188_315#_M1016_g N_A_42_47#_c_314_n 0.00391125f $X=2.305 $Y=2.465
+ $X2=0 $Y2=0
cc_170 N_A_188_315#_c_160_n N_A_42_47#_c_314_n 0.00314223f $X=3.615 $Y=1.08
+ $X2=0 $Y2=0
cc_171 N_A_188_315#_c_161_n N_A2_M1008_g 6.37827e-19 $X=3.78 $Y=1.97 $X2=0 $Y2=0
cc_172 N_A_188_315#_c_161_n N_A2_M1002_g 6.50897e-19 $X=3.78 $Y=1.97 $X2=0 $Y2=0
cc_173 N_A_188_315#_c_162_n N_A2_M1002_g 0.0146745f $X=5.015 $Y=1.08 $X2=0 $Y2=0
cc_174 N_A_188_315#_c_161_n N_A2_c_401_n 0.00475538f $X=3.78 $Y=1.97 $X2=0 $Y2=0
cc_175 N_A_188_315#_c_161_n N_A2_c_403_n 5.40555e-19 $X=3.78 $Y=1.97 $X2=0 $Y2=0
cc_176 N_A_188_315#_c_162_n N_A2_c_403_n 0.00439476f $X=5.015 $Y=1.08 $X2=0
+ $Y2=0
cc_177 N_A_188_315#_c_161_n N_A2_c_404_n 0.0126614f $X=3.78 $Y=1.97 $X2=0 $Y2=0
cc_178 N_A_188_315#_c_162_n N_A2_c_404_n 0.0267435f $X=5.015 $Y=1.08 $X2=0 $Y2=0
cc_179 N_A_188_315#_c_162_n N_A1_M1012_g 0.0141226f $X=5.015 $Y=1.08 $X2=0 $Y2=0
cc_180 N_A_188_315#_c_162_n N_A1_M1014_g 0.00280684f $X=5.015 $Y=1.08 $X2=0
+ $Y2=0
cc_181 N_A_188_315#_c_162_n N_A1_c_487_n 0.024394f $X=5.015 $Y=1.08 $X2=0 $Y2=0
cc_182 N_A_188_315#_c_162_n N_A1_c_488_n 7.69325e-19 $X=5.015 $Y=1.08 $X2=0
+ $Y2=0
cc_183 N_A_188_315#_c_163_n N_VPWR_c_536_n 0.0109552f $X=1.015 $Y=1.725 $X2=0
+ $Y2=0
cc_184 N_A_188_315#_c_166_n N_VPWR_c_536_n 0.00156061f $X=1.445 $Y=1.725 $X2=0
+ $Y2=0
cc_185 N_A_188_315#_c_163_n N_VPWR_c_537_n 0.00156061f $X=1.015 $Y=1.725 $X2=0
+ $Y2=0
cc_186 N_A_188_315#_c_166_n N_VPWR_c_537_n 0.0109982f $X=1.445 $Y=1.725 $X2=0
+ $Y2=0
cc_187 N_A_188_315#_M1009_g N_VPWR_c_537_n 0.0109982f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_188_315#_M1016_g N_VPWR_c_537_n 0.00156061f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_A_188_315#_M1009_g N_VPWR_c_538_n 0.00156061f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A_188_315#_M1016_g N_VPWR_c_538_n 0.012276f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A_188_315#_c_163_n N_VPWR_c_542_n 0.00486043f $X=1.015 $Y=1.725 $X2=0
+ $Y2=0
cc_192 N_A_188_315#_c_166_n N_VPWR_c_542_n 0.00486043f $X=1.445 $Y=1.725 $X2=0
+ $Y2=0
cc_193 N_A_188_315#_M1009_g N_VPWR_c_543_n 0.00486043f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_A_188_315#_M1016_g N_VPWR_c_543_n 0.00486043f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_188_315#_M1004_d N_VPWR_c_535_n 0.00225186f $X=3.64 $Y=1.835 $X2=0
+ $Y2=0
cc_196 N_A_188_315#_c_163_n N_VPWR_c_535_n 0.00451441f $X=1.015 $Y=1.725 $X2=0
+ $Y2=0
cc_197 N_A_188_315#_c_166_n N_VPWR_c_535_n 0.00451441f $X=1.445 $Y=1.725 $X2=0
+ $Y2=0
cc_198 N_A_188_315#_M1009_g N_VPWR_c_535_n 0.00451441f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A_188_315#_M1016_g N_VPWR_c_535_n 0.00451441f $X=2.305 $Y=2.465 $X2=0
+ $Y2=0
cc_200 N_A_188_315#_c_163_n N_X_c_627_n 0.00178848f $X=1.015 $Y=1.725 $X2=0
+ $Y2=0
cc_201 N_A_188_315#_c_149_n N_X_c_627_n 0.00635392f $X=1.245 $Y=1.65 $X2=0 $Y2=0
cc_202 N_A_188_315#_c_150_n N_X_c_627_n 0.0044673f $X=1.09 $Y=1.65 $X2=0 $Y2=0
cc_203 N_A_188_315#_M1001_g N_X_c_627_n 0.00845388f $X=1.32 $Y=0.655 $X2=0 $Y2=0
cc_204 N_A_188_315#_c_166_n N_X_c_627_n 0.00146658f $X=1.445 $Y=1.725 $X2=0
+ $Y2=0
cc_205 N_A_188_315#_M1009_g N_X_c_627_n 3.97256e-19 $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_206 N_A_188_315#_c_157_n N_X_c_627_n 0.0136179f $X=2.65 $Y=1.445 $X2=0 $Y2=0
cc_207 N_A_188_315#_c_149_n N_X_c_628_n 0.00148775f $X=1.245 $Y=1.65 $X2=0 $Y2=0
cc_208 N_A_188_315#_M1001_g N_X_c_628_n 0.0153272f $X=1.32 $Y=0.655 $X2=0 $Y2=0
cc_209 N_A_188_315#_c_157_n N_X_c_628_n 0.00631231f $X=2.65 $Y=1.445 $X2=0 $Y2=0
cc_210 N_A_188_315#_M1011_g N_X_c_630_n 0.0134504f $X=1.75 $Y=0.655 $X2=0 $Y2=0
cc_211 N_A_188_315#_M1018_g N_X_c_630_n 0.0132657f $X=2.18 $Y=0.655 $X2=0 $Y2=0
cc_212 N_A_188_315#_M1019_g N_X_c_630_n 0.00106524f $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_213 N_A_188_315#_c_157_n N_X_c_630_n 0.0588634f $X=2.65 $Y=1.445 $X2=0 $Y2=0
cc_214 N_A_188_315#_c_158_n N_X_c_630_n 0.00583384f $X=2.53 $Y=1.44 $X2=0 $Y2=0
cc_215 N_A_188_315#_c_159_n N_X_c_630_n 7.72671e-19 $X=2.735 $Y=1.355 $X2=0
+ $Y2=0
cc_216 N_A_188_315#_c_248_p N_X_c_630_n 0.0141411f $X=2.82 $Y=1.08 $X2=0 $Y2=0
cc_217 N_A_188_315#_M1019_g N_X_c_659_n 0.00562295f $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_218 N_A_188_315#_c_248_p N_X_c_659_n 7.52334e-19 $X=2.82 $Y=1.08 $X2=0 $Y2=0
cc_219 N_A_188_315#_c_157_n N_X_c_631_n 0.0147416f $X=2.65 $Y=1.445 $X2=0 $Y2=0
cc_220 N_A_188_315#_c_158_n N_X_c_631_n 0.00298081f $X=2.53 $Y=1.44 $X2=0 $Y2=0
cc_221 N_A_188_315#_c_163_n X 0.00745999f $X=1.015 $Y=1.725 $X2=0 $Y2=0
cc_222 N_A_188_315#_c_149_n X 0.00311899f $X=1.245 $Y=1.65 $X2=0 $Y2=0
cc_223 N_A_188_315#_c_166_n X 0.01563f $X=1.445 $Y=1.725 $X2=0 $Y2=0
cc_224 N_A_188_315#_M1009_g X 0.01563f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A_188_315#_M1016_g X 0.0191489f $X=2.305 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A_188_315#_c_157_n X 0.0749742f $X=2.65 $Y=1.445 $X2=0 $Y2=0
cc_227 N_A_188_315#_c_158_n X 0.0137879f $X=2.53 $Y=1.44 $X2=0 $Y2=0
cc_228 N_A_188_315#_c_163_n N_X_c_640_n 0.00755263f $X=1.015 $Y=1.725 $X2=0
+ $Y2=0
cc_229 N_A_188_315#_M1004_d N_A_645_367#_c_697_n 0.00332344f $X=3.64 $Y=1.835
+ $X2=0 $Y2=0
cc_230 N_A_188_315#_c_161_n N_A_645_367#_c_697_n 0.0159805f $X=3.78 $Y=1.97
+ $X2=0 $Y2=0
cc_231 N_A_188_315#_c_161_n N_A_645_367#_c_694_n 0.0200659f $X=3.78 $Y=1.97
+ $X2=0 $Y2=0
cc_232 N_A_188_315#_c_162_n N_A_645_367#_c_694_n 0.00554531f $X=5.015 $Y=1.08
+ $X2=0 $Y2=0
cc_233 N_A_188_315#_c_160_n N_VGND_M1019_s 0.00780768f $X=3.615 $Y=1.08 $X2=0
+ $Y2=0
cc_234 N_A_188_315#_c_248_p N_VGND_M1019_s 7.47232e-19 $X=2.82 $Y=1.08 $X2=0
+ $Y2=0
cc_235 N_A_188_315#_c_162_n N_VGND_M1020_s 0.00261503f $X=5.015 $Y=1.08 $X2=0
+ $Y2=0
cc_236 N_A_188_315#_M1001_g N_VGND_c_748_n 0.0111663f $X=1.32 $Y=0.655 $X2=0
+ $Y2=0
cc_237 N_A_188_315#_M1011_g N_VGND_c_748_n 6.28067e-19 $X=1.75 $Y=0.655 $X2=0
+ $Y2=0
cc_238 N_A_188_315#_M1001_g N_VGND_c_749_n 6.11179e-19 $X=1.32 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_A_188_315#_M1011_g N_VGND_c_749_n 0.010086f $X=1.75 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_188_315#_M1018_g N_VGND_c_749_n 0.0101197f $X=2.18 $Y=0.655 $X2=0
+ $Y2=0
cc_241 N_A_188_315#_M1019_g N_VGND_c_749_n 6.05913e-19 $X=2.62 $Y=0.655 $X2=0
+ $Y2=0
cc_242 N_A_188_315#_c_274_p N_VGND_c_750_n 0.0124525f $X=3.74 $Y=0.42 $X2=0
+ $Y2=0
cc_243 N_A_188_315#_c_162_n N_VGND_c_751_n 0.0218003f $X=5.015 $Y=1.08 $X2=0
+ $Y2=0
cc_244 N_A_188_315#_M1001_g N_VGND_c_754_n 0.00486043f $X=1.32 $Y=0.655 $X2=0
+ $Y2=0
cc_245 N_A_188_315#_M1011_g N_VGND_c_754_n 0.00486043f $X=1.75 $Y=0.655 $X2=0
+ $Y2=0
cc_246 N_A_188_315#_M1018_g N_VGND_c_757_n 0.00549879f $X=2.18 $Y=0.655 $X2=0
+ $Y2=0
cc_247 N_A_188_315#_M1019_g N_VGND_c_757_n 0.0168168f $X=2.62 $Y=0.655 $X2=0
+ $Y2=0
cc_248 N_A_188_315#_c_160_n N_VGND_c_757_n 0.048368f $X=3.615 $Y=1.08 $X2=0
+ $Y2=0
cc_249 N_A_188_315#_c_248_p N_VGND_c_757_n 0.00798224f $X=2.82 $Y=1.08 $X2=0
+ $Y2=0
cc_250 N_A_188_315#_M1005_d N_VGND_c_761_n 0.00536646f $X=3.6 $Y=0.235 $X2=0
+ $Y2=0
cc_251 N_A_188_315#_M1012_d N_VGND_c_761_n 0.00225186f $X=4.97 $Y=0.235 $X2=0
+ $Y2=0
cc_252 N_A_188_315#_M1001_g N_VGND_c_761_n 0.00824727f $X=1.32 $Y=0.655 $X2=0
+ $Y2=0
cc_253 N_A_188_315#_M1011_g N_VGND_c_761_n 0.00824727f $X=1.75 $Y=0.655 $X2=0
+ $Y2=0
cc_254 N_A_188_315#_M1018_g N_VGND_c_761_n 0.00827314f $X=2.18 $Y=0.655 $X2=0
+ $Y2=0
cc_255 N_A_188_315#_M1019_g N_VGND_c_761_n 0.00827319f $X=2.62 $Y=0.655 $X2=0
+ $Y2=0
cc_256 N_A_188_315#_c_274_p N_VGND_c_761_n 0.00730901f $X=3.74 $Y=0.42 $X2=0
+ $Y2=0
cc_257 N_A_188_315#_c_162_n N_A_908_47#_M1002_d 0.00176461f $X=5.015 $Y=1.08
+ $X2=-0.19 $Y2=-0.245
cc_258 N_A_188_315#_M1012_d N_A_908_47#_c_837_n 0.00332344f $X=4.97 $Y=0.235
+ $X2=0 $Y2=0
cc_259 N_A_188_315#_c_162_n N_A_908_47#_c_837_n 0.0031163f $X=5.015 $Y=1.08
+ $X2=0 $Y2=0
cc_260 N_A_188_315#_c_292_p N_A_908_47#_c_837_n 0.0124648f $X=5.11 $Y=0.76 $X2=0
+ $Y2=0
cc_261 N_A_188_315#_c_162_n N_A_908_47#_c_840_n 0.0168339f $X=5.015 $Y=1.08
+ $X2=0 $Y2=0
cc_262 N_A_188_315#_c_162_n N_A_908_47#_c_835_n 0.00137291f $X=5.015 $Y=1.08
+ $X2=0 $Y2=0
cc_263 N_A_42_47#_c_298_n N_A2_M1008_g 0.0209742f $X=3.995 $Y=1.51 $X2=0 $Y2=0
cc_264 N_A_42_47#_M1020_g N_A2_M1002_g 0.0256319f $X=3.955 $Y=0.655 $X2=0 $Y2=0
cc_265 N_A_42_47#_c_298_n N_A2_c_401_n 5.87646e-19 $X=3.995 $Y=1.51 $X2=0 $Y2=0
cc_266 N_A_42_47#_M1020_g N_A2_c_403_n 0.00261228f $X=3.955 $Y=0.655 $X2=0 $Y2=0
cc_267 N_A_42_47#_c_298_n N_A2_c_403_n 0.0186929f $X=3.995 $Y=1.51 $X2=0 $Y2=0
cc_268 N_A_42_47#_c_298_n N_A2_c_404_n 0.0012199f $X=3.995 $Y=1.51 $X2=0 $Y2=0
cc_269 N_A_42_47#_c_308_n N_VPWR_M1021_d 0.00350222f $X=2.905 $Y=2.455 $X2=-0.19
+ $Y2=-0.245
cc_270 N_A_42_47#_c_308_n N_VPWR_M1003_d 0.00350222f $X=2.905 $Y=2.455 $X2=0
+ $Y2=0
cc_271 N_A_42_47#_c_308_n N_VPWR_M1016_d 0.00517872f $X=2.905 $Y=2.455 $X2=0
+ $Y2=0
cc_272 N_A_42_47#_c_308_n N_VPWR_c_536_n 0.0166744f $X=2.905 $Y=2.455 $X2=0
+ $Y2=0
cc_273 N_A_42_47#_c_308_n N_VPWR_c_537_n 0.0166744f $X=2.905 $Y=2.455 $X2=0
+ $Y2=0
cc_274 N_A_42_47#_c_308_n N_VPWR_c_538_n 0.0214848f $X=2.905 $Y=2.455 $X2=0
+ $Y2=0
cc_275 N_A_42_47#_M1017_g N_VPWR_c_539_n 0.00109252f $X=3.995 $Y=2.465 $X2=0
+ $Y2=0
cc_276 N_A_42_47#_c_313_n N_VPWR_c_541_n 0.0257002f $X=0.37 $Y=2.495 $X2=0 $Y2=0
cc_277 N_A_42_47#_M1004_g N_VPWR_c_544_n 0.00357877f $X=3.565 $Y=2.465 $X2=0
+ $Y2=0
cc_278 N_A_42_47#_M1017_g N_VPWR_c_544_n 0.00357877f $X=3.995 $Y=2.465 $X2=0
+ $Y2=0
cc_279 N_A_42_47#_M1021_s N_VPWR_c_535_n 0.00246126f $X=0.245 $Y=1.835 $X2=0
+ $Y2=0
cc_280 N_A_42_47#_M1004_g N_VPWR_c_535_n 0.00665089f $X=3.565 $Y=2.465 $X2=0
+ $Y2=0
cc_281 N_A_42_47#_M1017_g N_VPWR_c_535_n 0.00537654f $X=3.995 $Y=2.465 $X2=0
+ $Y2=0
cc_282 N_A_42_47#_c_308_n N_VPWR_c_535_n 0.058646f $X=2.905 $Y=2.455 $X2=0 $Y2=0
cc_283 N_A_42_47#_c_313_n N_VPWR_c_535_n 0.0141073f $X=0.37 $Y=2.495 $X2=0 $Y2=0
cc_284 N_A_42_47#_c_308_n N_X_M1000_s 0.00488146f $X=2.905 $Y=2.455 $X2=0 $Y2=0
cc_285 N_A_42_47#_c_308_n N_X_M1009_s 0.00496259f $X=2.905 $Y=2.455 $X2=0 $Y2=0
cc_286 N_A_42_47#_c_308_n X 0.00861686f $X=2.905 $Y=2.455 $X2=0 $Y2=0
cc_287 N_A_42_47#_c_308_n X 0.0923053f $X=2.905 $Y=2.455 $X2=0 $Y2=0
cc_288 N_A_42_47#_c_314_n X 0.0326324f $X=3.112 $Y=1.875 $X2=0 $Y2=0
cc_289 N_A_42_47#_c_308_n N_X_c_640_n 0.0180752f $X=2.905 $Y=2.455 $X2=0 $Y2=0
cc_290 N_A_42_47#_c_314_n N_A_645_367#_M1004_s 0.00225602f $X=3.112 $Y=1.875
+ $X2=-0.19 $Y2=-0.245
cc_291 N_A_42_47#_c_297_n N_A_645_367#_c_702_n 0.00464136f $X=3.45 $Y=1.51 $X2=0
+ $Y2=0
cc_292 N_A_42_47#_c_308_n N_A_645_367#_c_702_n 0.0142846f $X=2.905 $Y=2.455
+ $X2=0 $Y2=0
cc_293 N_A_42_47#_c_309_n N_A_645_367#_c_702_n 0.0242923f $X=2.99 $Y=2.37 $X2=0
+ $Y2=0
cc_294 N_A_42_47#_c_314_n N_A_645_367#_c_702_n 0.00646238f $X=3.112 $Y=1.875
+ $X2=0 $Y2=0
cc_295 N_A_42_47#_M1004_g N_A_645_367#_c_697_n 0.0114565f $X=3.565 $Y=2.465
+ $X2=0 $Y2=0
cc_296 N_A_42_47#_M1017_g N_A_645_367#_c_697_n 0.0114565f $X=3.995 $Y=2.465
+ $X2=0 $Y2=0
cc_297 N_A_42_47#_M1017_g N_A_645_367#_c_694_n 5.21778e-19 $X=3.995 $Y=2.465
+ $X2=0 $Y2=0
cc_298 N_A_42_47#_M1005_g N_VGND_c_750_n 0.00487821f $X=3.525 $Y=0.655 $X2=0
+ $Y2=0
cc_299 N_A_42_47#_M1020_g N_VGND_c_750_n 0.00486043f $X=3.955 $Y=0.655 $X2=0
+ $Y2=0
cc_300 N_A_42_47#_M1005_g N_VGND_c_751_n 6.11179e-19 $X=3.525 $Y=0.655 $X2=0
+ $Y2=0
cc_301 N_A_42_47#_M1020_g N_VGND_c_751_n 0.0101096f $X=3.955 $Y=0.655 $X2=0
+ $Y2=0
cc_302 N_A_42_47#_c_299_n N_VGND_c_756_n 0.023546f $X=0.335 $Y=0.42 $X2=0 $Y2=0
cc_303 N_A_42_47#_M1005_g N_VGND_c_757_n 0.0116428f $X=3.525 $Y=0.655 $X2=0
+ $Y2=0
cc_304 N_A_42_47#_M1020_g N_VGND_c_757_n 6.26872e-19 $X=3.955 $Y=0.655 $X2=0
+ $Y2=0
cc_305 N_A_42_47#_M1013_s N_VGND_c_761_n 0.00371702f $X=0.21 $Y=0.235 $X2=0
+ $Y2=0
cc_306 N_A_42_47#_M1005_g N_VGND_c_761_n 0.00824731f $X=3.525 $Y=0.655 $X2=0
+ $Y2=0
cc_307 N_A_42_47#_M1020_g N_VGND_c_761_n 0.00824727f $X=3.955 $Y=0.655 $X2=0
+ $Y2=0
cc_308 N_A_42_47#_c_299_n N_VGND_c_761_n 0.0131407f $X=0.335 $Y=0.42 $X2=0 $Y2=0
cc_309 N_A2_M1002_g N_A1_M1012_g 0.0235613f $X=4.465 $Y=0.655 $X2=0 $Y2=0
cc_310 N_A2_c_403_n N_A1_M1012_g 0.0216583f $X=4.445 $Y=1.46 $X2=0 $Y2=0
cc_311 N_A2_c_404_n N_A1_M1012_g 0.00222012f $X=4.56 $Y=1.48 $X2=0 $Y2=0
cc_312 A2 N_A1_M1006_g 0.0135148f $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_313 N_A2_M1007_g N_A1_M1014_g 0.029101f $X=5.755 $Y=0.655 $X2=0 $Y2=0
cc_314 N_A2_c_405_n N_A1_M1014_g 0.00305366f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_315 N_A2_M1010_g N_A1_M1015_g 0.029101f $X=5.755 $Y=2.465 $X2=0 $Y2=0
cc_316 A2 N_A1_M1015_g 0.0146927f $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_317 N_A2_c_401_n N_A1_c_487_n 0.00808075f $X=4.56 $Y=1.94 $X2=0 $Y2=0
cc_318 N_A2_c_402_n N_A1_c_487_n 0.00964898f $X=5.55 $Y=1.94 $X2=0 $Y2=0
cc_319 N_A2_c_403_n N_A1_c_487_n 2.92617e-19 $X=4.445 $Y=1.46 $X2=0 $Y2=0
cc_320 N_A2_c_404_n N_A1_c_487_n 0.0166287f $X=4.56 $Y=1.48 $X2=0 $Y2=0
cc_321 N_A2_c_405_n N_A1_c_487_n 0.0250397f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_322 N_A2_c_406_n N_A1_c_487_n 2.50566e-19 $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_323 A2 N_A1_c_487_n 0.0243849f $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_324 N_A2_M1008_g N_A1_c_488_n 0.0446586f $X=4.425 $Y=2.465 $X2=0 $Y2=0
cc_325 N_A2_c_401_n N_A1_c_488_n 0.00460666f $X=4.56 $Y=1.94 $X2=0 $Y2=0
cc_326 N_A2_c_402_n N_A1_c_488_n 0.00310497f $X=5.55 $Y=1.94 $X2=0 $Y2=0
cc_327 N_A2_c_406_n N_A1_c_488_n 0.029101f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_328 A2 N_A1_c_488_n 5.53026e-19 $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_329 N_A2_c_401_n N_VPWR_M1008_d 0.0021661f $X=4.56 $Y=1.94 $X2=0 $Y2=0
cc_330 A2 N_VPWR_M1008_d 0.00574419f $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_331 N_A2_c_402_n N_VPWR_M1015_s 0.00247598f $X=5.55 $Y=1.94 $X2=0 $Y2=0
cc_332 N_A2_M1008_g N_VPWR_c_539_n 0.0116435f $X=4.425 $Y=2.465 $X2=0 $Y2=0
cc_333 N_A2_M1010_g N_VPWR_c_540_n 0.0122401f $X=5.755 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A2_M1008_g N_VPWR_c_544_n 0.00486043f $X=4.425 $Y=2.465 $X2=0 $Y2=0
cc_335 N_A2_M1010_g N_VPWR_c_546_n 0.00486043f $X=5.755 $Y=2.465 $X2=0 $Y2=0
cc_336 N_A2_M1008_g N_VPWR_c_535_n 0.0082726f $X=4.425 $Y=2.465 $X2=0 $Y2=0
cc_337 N_A2_M1010_g N_VPWR_c_535_n 0.00918921f $X=5.755 $Y=2.465 $X2=0 $Y2=0
cc_338 A2 N_A_645_367#_M1006_d 0.00333747f $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_339 N_A2_M1008_g N_A_645_367#_c_694_n 5.21778e-19 $X=4.425 $Y=2.465 $X2=0
+ $Y2=0
cc_340 N_A2_c_401_n N_A_645_367#_c_694_n 0.00637253f $X=4.56 $Y=1.94 $X2=0 $Y2=0
cc_341 N_A2_c_403_n N_A_645_367#_c_694_n 5.59096e-19 $X=4.445 $Y=1.46 $X2=0
+ $Y2=0
cc_342 N_A2_c_404_n N_A_645_367#_c_694_n 0.00200627f $X=4.56 $Y=1.48 $X2=0 $Y2=0
cc_343 N_A2_M1008_g N_A_645_367#_c_714_n 0.0142935f $X=4.425 $Y=2.465 $X2=0
+ $Y2=0
cc_344 N_A2_c_401_n N_A_645_367#_c_714_n 0.00874961f $X=4.56 $Y=1.94 $X2=0 $Y2=0
cc_345 N_A2_c_403_n N_A_645_367#_c_714_n 2.37977e-19 $X=4.445 $Y=1.46 $X2=0
+ $Y2=0
cc_346 N_A2_c_404_n N_A_645_367#_c_714_n 0.00337393f $X=4.56 $Y=1.48 $X2=0 $Y2=0
cc_347 A2 N_A_645_367#_c_714_n 0.0187491f $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_348 N_A2_M1010_g N_A_645_367#_c_719_n 0.0143943f $X=5.755 $Y=2.465 $X2=0
+ $Y2=0
cc_349 N_A2_c_402_n N_A_645_367#_c_719_n 0.0131194f $X=5.55 $Y=1.94 $X2=0 $Y2=0
cc_350 N_A2_c_405_n N_A_645_367#_c_719_n 0.00383255f $X=5.845 $Y=1.51 $X2=0
+ $Y2=0
cc_351 A2 N_A_645_367#_c_719_n 0.0101781f $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_352 N_A2_M1010_g N_A_645_367#_c_695_n 0.00118035f $X=5.755 $Y=2.465 $X2=0
+ $Y2=0
cc_353 N_A2_c_402_n N_A_645_367#_c_695_n 0.00152757f $X=5.55 $Y=1.94 $X2=0 $Y2=0
cc_354 N_A2_c_405_n N_A_645_367#_c_695_n 0.0145803f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_355 N_A2_c_406_n N_A_645_367#_c_695_n 0.00419966f $X=5.845 $Y=1.51 $X2=0
+ $Y2=0
cc_356 A2 N_A_645_367#_c_727_n 0.0135577f $X=5.435 $Y=1.95 $X2=0 $Y2=0
cc_357 N_A2_M1002_g N_VGND_c_751_n 0.00610432f $X=4.465 $Y=0.655 $X2=0 $Y2=0
cc_358 N_A2_M1007_g N_VGND_c_753_n 0.00840623f $X=5.755 $Y=0.655 $X2=0 $Y2=0
cc_359 N_A2_c_405_n N_VGND_c_753_n 0.0104826f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_360 N_A2_c_406_n N_VGND_c_753_n 0.00115467f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_361 N_A2_M1002_g N_VGND_c_758_n 0.00547432f $X=4.465 $Y=0.655 $X2=0 $Y2=0
cc_362 N_A2_M1007_g N_VGND_c_758_n 0.00577794f $X=5.755 $Y=0.655 $X2=0 $Y2=0
cc_363 N_A2_M1002_g N_VGND_c_761_n 0.0101107f $X=4.465 $Y=0.655 $X2=0 $Y2=0
cc_364 N_A2_M1007_g N_VGND_c_761_n 0.0113461f $X=5.755 $Y=0.655 $X2=0 $Y2=0
cc_365 N_A2_M1002_g N_A_908_47#_c_840_n 0.00649214f $X=4.465 $Y=0.655 $X2=0
+ $Y2=0
cc_366 N_A2_M1007_g N_A_908_47#_c_835_n 0.00910838f $X=5.755 $Y=0.655 $X2=0
+ $Y2=0
cc_367 N_A2_c_405_n N_A_908_47#_c_835_n 0.0168511f $X=5.845 $Y=1.51 $X2=0 $Y2=0
cc_368 N_A1_M1006_g N_VPWR_c_539_n 0.00243207f $X=4.895 $Y=2.465 $X2=0 $Y2=0
cc_369 N_A1_M1006_g N_VPWR_c_540_n 5.9204e-19 $X=4.895 $Y=2.465 $X2=0 $Y2=0
cc_370 N_A1_M1015_g N_VPWR_c_540_n 0.0106448f $X=5.325 $Y=2.465 $X2=0 $Y2=0
cc_371 N_A1_M1006_g N_VPWR_c_545_n 0.00585385f $X=4.895 $Y=2.465 $X2=0 $Y2=0
cc_372 N_A1_M1015_g N_VPWR_c_545_n 0.00486043f $X=5.325 $Y=2.465 $X2=0 $Y2=0
cc_373 N_A1_M1006_g N_VPWR_c_535_n 0.0107716f $X=4.895 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A1_M1015_g N_VPWR_c_535_n 0.00824727f $X=5.325 $Y=2.465 $X2=0 $Y2=0
cc_375 N_A1_M1006_g N_A_645_367#_c_714_n 0.013172f $X=4.895 $Y=2.465 $X2=0 $Y2=0
cc_376 N_A1_M1015_g N_A_645_367#_c_719_n 0.0122129f $X=5.325 $Y=2.465 $X2=0
+ $Y2=0
cc_377 N_A1_M1012_g N_VGND_c_758_n 0.00357842f $X=4.895 $Y=0.655 $X2=0 $Y2=0
cc_378 N_A1_M1014_g N_VGND_c_758_n 0.00357877f $X=5.325 $Y=0.655 $X2=0 $Y2=0
cc_379 N_A1_M1012_g N_VGND_c_761_n 0.00537652f $X=4.895 $Y=0.655 $X2=0 $Y2=0
cc_380 N_A1_M1014_g N_VGND_c_761_n 0.00537654f $X=5.325 $Y=0.655 $X2=0 $Y2=0
cc_381 N_A1_M1012_g N_A_908_47#_c_837_n 0.0083305f $X=4.895 $Y=0.655 $X2=0 $Y2=0
cc_382 N_A1_M1014_g N_A_908_47#_c_837_n 0.012237f $X=5.325 $Y=0.655 $X2=0 $Y2=0
cc_383 N_A1_M1012_g N_A_908_47#_c_840_n 0.00634543f $X=4.895 $Y=0.655 $X2=0
+ $Y2=0
cc_384 N_A1_M1014_g N_A_908_47#_c_840_n 5.12214e-19 $X=5.325 $Y=0.655 $X2=0
+ $Y2=0
cc_385 N_A1_M1014_g N_A_908_47#_c_835_n 6.89974e-19 $X=5.325 $Y=0.655 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_535_n N_X_M1000_s 0.00389913f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_387 N_VPWR_c_535_n N_X_M1009_s 0.00389913f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_388 N_VPWR_M1003_d X 0.0018161f $X=1.52 $Y=1.835 $X2=0 $Y2=0
cc_389 N_VPWR_M1016_d X 0.00398813f $X=2.38 $Y=1.835 $X2=0 $Y2=0
cc_390 N_VPWR_M1021_d N_X_c_640_n 0.0059201f $X=0.66 $Y=1.835 $X2=0 $Y2=0
cc_391 N_VPWR_c_535_n N_A_645_367#_M1004_s 0.00284736f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_392 N_VPWR_c_535_n N_A_645_367#_M1017_s 0.00376627f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_393 N_VPWR_c_535_n N_A_645_367#_M1006_d 0.00397496f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_394 N_VPWR_c_535_n N_A_645_367#_M1010_s 0.00371702f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_395 N_VPWR_c_538_n N_A_645_367#_c_734_n 0.00623131f $X=2.52 $Y=2.875 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_544_n N_A_645_367#_c_734_n 0.0136445f $X=4.475 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_535_n N_A_645_367#_c_734_n 0.00777554f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_398 N_VPWR_c_538_n N_A_645_367#_c_702_n 0.00652289f $X=2.52 $Y=2.875 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_544_n N_A_645_367#_c_697_n 0.0486406f $X=4.475 $Y=3.33 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_535_n N_A_645_367#_c_697_n 0.0310522f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_401 N_VPWR_M1008_d N_A_645_367#_c_714_n 0.00433179f $X=4.5 $Y=1.835 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_539_n N_A_645_367#_c_714_n 0.0185459f $X=4.64 $Y=2.75 $X2=0
+ $Y2=0
cc_403 N_VPWR_M1015_s N_A_645_367#_c_719_n 0.00352922f $X=5.4 $Y=1.835 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_540_n N_A_645_367#_c_719_n 0.0170777f $X=5.54 $Y=2.75 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_545_n N_A_645_367#_c_727_n 0.0138717f $X=5.375 $Y=3.33 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_535_n N_A_645_367#_c_727_n 0.00886411f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_407 N_VPWR_c_546_n N_A_645_367#_c_696_n 0.0178111f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_408 N_VPWR_c_535_n N_A_645_367#_c_696_n 0.0100304f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_409 N_X_c_628_n N_VGND_M1013_d 2.33864e-19 $X=1.44 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_410 N_X_c_629_n N_VGND_M1013_d 0.00327847f $X=1.165 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_411 N_X_c_630_n N_VGND_M1011_s 0.00180746f $X=2.3 $Y=1.09 $X2=0 $Y2=0
cc_412 N_X_c_628_n N_VGND_c_748_n 0.00362085f $X=1.44 $Y=1.09 $X2=0 $Y2=0
cc_413 N_X_c_629_n N_VGND_c_748_n 0.0153275f $X=1.165 $Y=1.09 $X2=0 $Y2=0
cc_414 N_X_c_630_n N_VGND_c_749_n 0.0163515f $X=2.3 $Y=1.09 $X2=0 $Y2=0
cc_415 N_X_c_688_p N_VGND_c_754_n 0.0124525f $X=1.535 $Y=0.42 $X2=0 $Y2=0
cc_416 N_X_c_659_n N_VGND_c_757_n 0.0532148f $X=2.395 $Y=0.42 $X2=0 $Y2=0
cc_417 N_X_M1001_d N_VGND_c_761_n 0.00536646f $X=1.395 $Y=0.235 $X2=0 $Y2=0
cc_418 N_X_M1018_d N_VGND_c_761_n 0.00614263f $X=2.255 $Y=0.235 $X2=0 $Y2=0
cc_419 N_X_c_688_p N_VGND_c_761_n 0.00730901f $X=1.535 $Y=0.42 $X2=0 $Y2=0
cc_420 N_X_c_659_n N_VGND_c_761_n 0.00692023f $X=2.395 $Y=0.42 $X2=0 $Y2=0
cc_421 N_VGND_c_761_n N_A_908_47#_M1002_d 0.00223559f $X=6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_422 N_VGND_c_761_n N_A_908_47#_M1014_s 0.00223561f $X=6 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_758_n N_A_908_47#_c_837_n 0.0326395f $X=5.855 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_761_n N_A_908_47#_c_837_n 0.0208532f $X=6 $Y=0 $X2=0 $Y2=0
cc_425 N_VGND_c_758_n N_A_908_47#_c_840_n 0.0188708f $X=5.855 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_761_n N_A_908_47#_c_840_n 0.0123968f $X=6 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_753_n N_A_908_47#_c_835_n 0.0248279f $X=5.97 $Y=0.38 $X2=0 $Y2=0
cc_428 N_VGND_c_758_n N_A_908_47#_c_835_n 0.0147831f $X=5.855 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_761_n N_A_908_47#_c_835_n 0.00962336f $X=6 $Y=0 $X2=0 $Y2=0
