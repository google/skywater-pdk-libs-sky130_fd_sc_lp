* File: sky130_fd_sc_lp__nor4b_1.spice
* Created: Fri Aug 28 10:58:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4b_1.pex.spice"
.subckt sky130_fd_sc_lp__nor4b_1  VNB VPB D_N A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_D_N_M1005_g N_A_80_131#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0917 AS=0.1113 PD=0.82 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84 AD=0.1365
+ AS=0.1834 PD=1.165 PS=1.64 NRD=6.42 NRS=7.848 M=1 R=5.6 SA=75000.5 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.84 AD=0.1617
+ AS=0.1365 PD=1.225 PS=1.165 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.9 SB=75001.2
+ A=0.126 P=1.98 MULT=1
MM1008 N_Y_M1008_d N_C_M1008_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1617 PD=1.12 PS=1.225 NRD=0 NRS=7.848 M=1 R=5.6 SA=75001.5 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_80_131#_M1004_g N_Y_M1008_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_D_N_M1009_g N_A_80_131#_M1009_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0966 AS=0.1113 PD=0.825 PS=1.37 NRD=82.0702 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1001 A_271_367# N_A_M1001_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.2898 PD=1.47 PS=2.475 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.4 SB=75001.7
+ A=0.189 P=2.82 MULT=1
MM1003 A_343_367# N_B_M1003_g A_271_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75000.7
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1007 A_451_367# N_C_M1007_g A_343_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.2457 PD=1.65 PS=1.65 NRD=21.8867 NRS=21.8867 M=1 R=8.4 SA=75001.3
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1000 N_Y_M1000_d N_A_80_131#_M1000_g A_451_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.378 AS=0.2457 PD=3.12 PS=1.65 NRD=5.4569 NRS=21.8867 M=1 R=8.4 SA=75001.8
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__nor4b_1.pxi.spice"
*
.ends
*
*
