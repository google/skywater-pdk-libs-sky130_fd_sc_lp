* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlrbn_lp D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
X0 VGND GATE_N a_272_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_68# D a_114_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_27_68# a_758_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_451_419# a_252_396# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_1277_153# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_952_305# a_796_419# a_1277_153# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1861_76# a_1617_76# Q_N VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_796_419# a_952_305# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VGND a_952_305# a_1435_153# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_27_68# a_698_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_796_419# a_252_396# a_904_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 VPWR a_1617_76# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_698_419# a_451_419# a_796_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_904_419# a_952_305# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 a_1703_76# a_952_305# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_451_419# a_252_396# a_542_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_950_47# a_952_305# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_1617_76# a_1861_76# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_68# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X19 VPWR a_952_305# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 a_272_68# GATE_N a_252_396# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1617_76# a_952_305# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_758_47# a_252_396# a_796_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_1435_153# a_952_305# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_542_47# a_252_396# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_796_419# a_451_419# a_950_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_952_305# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 VPWR GATE_N a_252_396# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X28 a_1617_76# a_952_305# a_1703_76# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_114_68# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
