* File: sky130_fd_sc_lp__mux2i_lp.spice
* Created: Wed Sep  2 10:01:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2i_lp.pex.spice"
.subckt sky130_fd_sc_lp__mux2i_lp  VNB VPB S A1 A0 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1001 A_114_49# N_S_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_A1_M1008_g A_114_49# VNB NSHORT L=0.15 W=0.42 AD=0.1419
+ AS=0.0504 PD=1.17 PS=0.66 NRD=80.808 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1005 A_324_49# N_A0_M1005_g N_Y_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1419 PD=0.66 PS=1.17 NRD=18.564 NRS=80.808 M=1 R=2.8 SA=75001.3
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_365_255#_M1006_g A_324_49# VNB NSHORT L=0.15 W=0.42
+ AD=0.08085 AS=0.0504 PD=0.805 PS=0.66 NRD=21.42 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 A_509_49# N_S_M1003_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.08085 PD=0.66 PS=0.805 NRD=18.564 NRS=8.568 M=1 R=2.8 SA=75002.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_365_255#_M1004_d N_S_M1004_g A_509_49# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 A_125_527# N_S_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A0_M1002_g A_125_527# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75000.6 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1009 A_289_527# N_A1_M1009_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0798
+ AS=0.0588 PD=0.8 PS=0.7 NRD=63.3158 NRS=0 M=1 R=2.8 SA=75001 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_365_255#_M1007_g A_289_527# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.08925 AS=0.0798 PD=0.845 PS=0.8 NRD=68.0044 NRS=63.3158 M=1 R=2.8
+ SA=75001.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 A_510_527# N_S_M1011_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.08925 PD=0.63 PS=0.845 NRD=23.443 NRS=0 M=1 R=2.8 SA=75002.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_365_255#_M1000_d N_S_M1000_g A_510_527# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__mux2i_lp.pxi.spice"
*
.ends
*
*
