* File: sky130_fd_sc_lp__isobufsrc_1.spice
* Created: Fri Aug 28 10:41:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__isobufsrc_1.pex.spice"
.subckt sky130_fd_sc_lp__isobufsrc_1  VNB VPB A SLEEP VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_79_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1036 AS=0.1113 PD=0.863333 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_SLEEP_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2072 PD=1.12 PS=1.72667 NRD=0 NRS=12.492 M=1 R=5.6 SA=75000.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A_79_47#_M1001_g N_X_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_79_47#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0966 AS=0.1113 PD=0.825 PS=1.37 NRD=82.0702 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1005 A_283_367# N_SLEEP_M1005_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.2898 PD=1.47 PS=2.475 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1000 N_X_M1000_d N_A_79_47#_M1000_g A_283_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.6174 AS=0.1323 PD=3.5 PS=1.47 NRD=14.8341 NRS=7.8012 M=1 R=8.4 SA=75000.7
+ SB=75000.4 A=0.189 P=2.82 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__isobufsrc_1.pxi.spice"
*
.ends
*
*
