* File: sky130_fd_sc_lp__a32o_m.pex.spice
* Created: Fri Aug 28 10:01:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32O_M%A_84_153# 1 2 11 14 16 17 18 20 25 27 30 31
+ 36 38 40
c89 16 0 1.80904e-19 $X=0.51 $Y=0.765
r90 34 36 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=2.57 $Y=2.05 $X2=2.65
+ $Y2=2.05
r91 31 41 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.5
+ $X2=0.587 $Y2=1.665
r92 31 40 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.5
+ $X2=0.587 $Y2=1.335
r93 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.5 $X2=0.59 $Y2=1.5
r94 27 36 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.65 $Y=1.945
+ $X2=2.65 $Y2=2.05
r95 26 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=1.505
+ $X2=2.65 $Y2=1.42
r96 26 27 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.65 $Y=1.505
+ $X2=2.65 $Y2=1.945
r97 25 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=1.335
+ $X2=2.65 $Y2=1.42
r98 24 25 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.65 $Y=0.585
+ $X2=2.65 $Y2=1.335
r99 20 24 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.565 $Y=0.48
+ $X2=2.65 $Y2=0.585
r100 20 22 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=2.565 $Y=0.48
+ $X2=2.29 $Y2=0.48
r101 19 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=1.42
+ $X2=0.59 $Y2=1.42
r102 18 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=1.42
+ $X2=2.65 $Y2=1.42
r103 18 19 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=2.565 $Y=1.42
+ $X2=0.675 $Y2=1.42
r104 17 40 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.495 $Y=0.915
+ $X2=0.495 $Y2=1.335
r105 16 17 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.51 $Y=0.765
+ $X2=0.51 $Y2=0.915
r106 14 41 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.555 $Y=2.135
+ $X2=0.555 $Y2=1.665
r107 11 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.525 $Y=0.445
+ $X2=0.525 $Y2=0.765
r108 2 34 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.925 $X2=2.57 $Y2=2.05
r109 1 22 182 $w=1.7e-07 $l=3.51781e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.235 $X2=2.29 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_M%A3 3 6 8 11 12 13
c37 6 0 2.66518e-19 $X=1.065 $Y=2.135
r38 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=0.93
+ $X2=0.975 $Y2=1.095
r39 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=0.93
+ $X2=0.975 $Y2=0.765
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=0.93 $X2=0.975 $Y2=0.93
r41 8 12 16.161 $w=1.73e-07 $l=2.55e-07 $layer=LI1_cond $X=0.72 $Y=0.927
+ $X2=0.975 $Y2=0.927
r42 6 14 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.065 $Y=2.135
+ $X2=1.065 $Y2=1.095
r43 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.065 $Y=0.445
+ $X2=1.065 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_M%A2 3 6 8 9 13 15
r34 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=0.93
+ $X2=1.515 $Y2=1.095
r35 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=0.93
+ $X2=1.515 $Y2=0.765
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.515
+ $Y=0.93 $X2=1.515 $Y2=0.93
r37 9 14 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=1.557 $Y=0.925
+ $X2=1.557 $Y2=0.93
r38 8 9 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.557 $Y=0.555
+ $X2=1.557 $Y2=0.925
r39 6 16 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.495 $Y=2.135
+ $X2=1.495 $Y2=1.095
r40 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.425 $Y=0.445
+ $X2=1.425 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_M%A1 3 7 10 11 12 15 17
r44 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.055 $Y=0.93
+ $X2=2.055 $Y2=1.095
r45 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.055 $Y=0.93
+ $X2=2.055 $Y2=0.765
r46 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=0.93 $X2=2.055 $Y2=0.93
r47 12 16 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.16 $Y=0.93
+ $X2=2.055 $Y2=0.93
r48 10 11 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.945 $Y=1.335
+ $X2=1.945 $Y2=1.485
r49 10 18 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.965 $Y=1.335
+ $X2=1.965 $Y2=1.095
r50 7 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.965 $Y=0.445
+ $X2=1.965 $Y2=0.765
r51 3 11 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.925 $Y=2.135
+ $X2=1.925 $Y2=1.485
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_M%B1 4 7 11 13 14 15 16 17 24
c47 17 0 1.64219e-19 $X=3.12 $Y=2.775
c48 4 0 2.98451e-19 $X=2.355 $Y=2.135
r49 24 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=2.88
+ $X2=2.265 $Y2=2.715
r50 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.265
+ $Y=2.88 $X2=2.265 $Y2=2.88
r51 16 17 20.1154 $w=2.73e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=2.827
+ $X2=3.12 $Y2=2.827
r52 16 25 15.7151 $w=2.73e-07 $l=3.75e-07 $layer=LI1_cond $X=2.64 $Y=2.827
+ $X2=2.265 $Y2=2.827
r53 15 25 4.40024 $w=2.73e-07 $l=1.05e-07 $layer=LI1_cond $X=2.16 $Y=2.827
+ $X2=2.265 $Y2=2.827
r54 14 15 20.1154 $w=2.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.827
+ $X2=2.16 $Y2=2.827
r55 13 14 20.1154 $w=2.73e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.827
+ $X2=1.68 $Y2=2.827
r56 9 11 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.355 $Y=1.38
+ $X2=2.505 $Y2=1.38
r57 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=1.305
+ $X2=2.505 $Y2=1.38
r58 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.505 $Y=1.305
+ $X2=2.505 $Y2=0.445
r59 4 26 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.355 $Y=2.135
+ $X2=2.355 $Y2=2.715
r60 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.355 $Y=1.455
+ $X2=2.355 $Y2=1.38
r61 1 4 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.355 $Y=1.455
+ $X2=2.355 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_M%B2 1 3 6 9 12 16 18 19 20 21 26
c38 19 0 1.11231e-19 $X=3.12 $Y=0.925
r39 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=1.295
+ $X2=3.105 $Y2=1.665
r40 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.105 $Y=0.925
+ $X2=3.105 $Y2=1.295
r41 19 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.005 $X2=3.09 $Y2=1.005
r42 17 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.09 $Y=1.345
+ $X2=3.09 $Y2=1.005
r43 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.345
+ $X2=3.09 $Y2=1.51
r44 16 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.09 $Y=0.99
+ $X2=3.09 $Y2=1.005
r45 15 16 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.022 $Y=0.84
+ $X2=3.022 $Y2=0.99
r46 10 12 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.785 $Y=1.74 $X2=3
+ $Y2=1.74
r47 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3 $Y=1.665 $X2=3
+ $Y2=1.74
r48 9 18 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=3 $Y=1.665 $X2=3
+ $Y2=1.51
r49 6 15 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.865 $Y=0.445
+ $X2=2.865 $Y2=0.84
r50 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.785 $Y=1.815
+ $X2=2.785 $Y2=1.74
r51 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.785 $Y=1.815
+ $X2=2.785 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_M%X 1 2 9 16 18
c14 9 0 1.80904e-19 $X=0.29 $Y=0.495
r15 13 18 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.24 $Y=1.905
+ $X2=0.24 $Y2=0.925
r16 12 16 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.24 $Y=2.07 $X2=0.34
+ $Y2=2.07
r17 12 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=2.07
+ $X2=0.24 $Y2=1.905
r18 11 18 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.24 $Y=0.66
+ $X2=0.24 $Y2=0.925
r19 9 11 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=0.495
+ $X2=0.275 $Y2=0.66
r20 2 16 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.925 $X2=0.34 $Y2=2.07
r21 1 9 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_M%VPWR 1 2 9 12 13 17 19 20 22 32 33 36
c28 13 0 1.8722e-19 $X=1.625 $Y=2.42
r29 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r31 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r33 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r34 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=0.77 $Y2=3.33
r35 27 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=1.2 $Y2=3.33
r36 25 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.77 $Y2=3.33
r39 22 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 20 33 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 20 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 15 17 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.72 $Y=2.335
+ $X2=1.72 $Y2=2.2
r43 14 19 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=2.42
+ $X2=0.77 $Y2=2.42
r44 13 15 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.625 $Y=2.42
+ $X2=1.72 $Y2=2.335
r45 13 14 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.625 $Y=2.42
+ $X2=0.935 $Y2=2.42
r46 12 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=3.33
r47 11 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=2.505
+ $X2=0.77 $Y2=2.42
r48 11 12 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=0.77 $Y=2.505
+ $X2=0.77 $Y2=3.245
r49 7 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=2.335 $X2=0.77
+ $Y2=2.42
r50 7 9 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.77 $Y=2.335
+ $X2=0.77 $Y2=2.05
r51 2 17 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.925 $X2=1.71 $Y2=2.2
r52 1 9 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.925 $X2=0.77 $Y2=2.05
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_M%A_228_385# 1 2 3 10 15 16 17 20 22
c36 10 0 1.023e-19 $X=2.035 $Y=1.77
r37 22 25 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.28 $Y=1.77 $X2=1.28
+ $Y2=2.05
r38 18 20 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=3.02 $Y=2.335
+ $X2=3.02 $Y2=2.2
r39 16 18 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.915 $Y=2.42
+ $X2=3.02 $Y2=2.335
r40 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.915 $Y=2.42
+ $X2=2.225 $Y2=2.42
r41 13 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.13 $Y=2.335
+ $X2=2.225 $Y2=2.42
r42 13 15 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=2.13 $Y=2.335
+ $X2=2.13 $Y2=2.2
r43 12 15 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=2.13 $Y=1.855
+ $X2=2.13 $Y2=2.2
r44 11 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=1.77
+ $X2=1.28 $Y2=1.77
r45 10 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.035 $Y=1.77
+ $X2=2.13 $Y2=1.855
r46 10 11 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.035 $Y=1.77
+ $X2=1.445 $Y2=1.77
r47 3 20 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.925 $X2=3.02 $Y2=2.2
r48 2 15 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.925 $X2=2.14 $Y2=2.2
r49 1 25 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.925 $X2=1.28 $Y2=2.05
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_M%VGND 1 2 9 11 13 15 17 22 31 35
r50 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r51 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r53 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r55 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r56 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r57 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.74
+ $Y2=0
r58 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.2
+ $Y2=0
r59 22 34 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r60 22 28 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r61 20 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r62 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.74
+ $Y2=0
r64 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.24
+ $Y2=0
r65 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r66 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r67 11 34 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r68 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.38
r69 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0
r70 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.38
r71 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.38
r72 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.38
.ends

