* File: sky130_fd_sc_lp__a221o_0.pxi.spice
* Created: Fri Aug 28 09:52:21 2020
* 
x_PM_SKY130_FD_SC_LP__A221O_0%A_72_312# N_A_72_312#_M1005_d N_A_72_312#_M1010_d
+ N_A_72_312#_M1011_d N_A_72_312#_M1000_g N_A_72_312#_M1003_g N_A_72_312#_c_96_n
+ N_A_72_312#_c_97_n N_A_72_312#_c_84_n N_A_72_312#_c_98_n N_A_72_312#_c_85_n
+ N_A_72_312#_c_86_n N_A_72_312#_c_87_n N_A_72_312#_c_88_n N_A_72_312#_c_89_n
+ N_A_72_312#_c_90_n N_A_72_312#_c_91_n N_A_72_312#_c_101_n N_A_72_312#_c_102_n
+ N_A_72_312#_c_92_n N_A_72_312#_c_93_n N_A_72_312#_c_103_n N_A_72_312#_c_94_n
+ PM_SKY130_FD_SC_LP__A221O_0%A_72_312#
x_PM_SKY130_FD_SC_LP__A221O_0%A2 N_A2_M1001_g N_A2_M1009_g N_A2_c_207_n
+ N_A2_c_208_n A2 N_A2_c_210_n PM_SKY130_FD_SC_LP__A221O_0%A2
x_PM_SKY130_FD_SC_LP__A221O_0%A1 N_A1_M1007_g N_A1_M1005_g N_A1_c_252_n
+ N_A1_c_253_n N_A1_c_259_n N_A1_c_254_n A1 A1 N_A1_c_256_n
+ PM_SKY130_FD_SC_LP__A221O_0%A1
x_PM_SKY130_FD_SC_LP__A221O_0%B1 N_B1_c_298_n N_B1_M1004_g N_B1_M1002_g B1 B1
+ N_B1_c_301_n PM_SKY130_FD_SC_LP__A221O_0%B1
x_PM_SKY130_FD_SC_LP__A221O_0%B2 N_B2_M1006_g N_B2_M1008_g B2 N_B2_c_336_n
+ N_B2_c_337_n PM_SKY130_FD_SC_LP__A221O_0%B2
x_PM_SKY130_FD_SC_LP__A221O_0%C1 N_C1_M1010_g N_C1_M1011_g C1 N_C1_c_372_n
+ PM_SKY130_FD_SC_LP__A221O_0%C1
x_PM_SKY130_FD_SC_LP__A221O_0%X N_X_M1003_s N_X_M1000_s N_X_c_405_n N_X_c_401_n
+ X X X N_X_c_403_n X PM_SKY130_FD_SC_LP__A221O_0%X
x_PM_SKY130_FD_SC_LP__A221O_0%VPWR N_VPWR_M1000_d N_VPWR_M1007_d N_VPWR_c_427_n
+ N_VPWR_c_428_n VPWR N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_426_n
+ N_VPWR_c_432_n N_VPWR_c_433_n PM_SKY130_FD_SC_LP__A221O_0%VPWR
x_PM_SKY130_FD_SC_LP__A221O_0%A_216_484# N_A_216_484#_M1001_d
+ N_A_216_484#_M1002_d N_A_216_484#_c_467_n N_A_216_484#_c_468_n
+ N_A_216_484#_c_469_n N_A_216_484#_c_474_n
+ PM_SKY130_FD_SC_LP__A221O_0%A_216_484#
x_PM_SKY130_FD_SC_LP__A221O_0%A_409_429# N_A_409_429#_M1002_s
+ N_A_409_429#_M1008_d N_A_409_429#_c_504_n N_A_409_429#_c_505_n
+ N_A_409_429#_c_506_n N_A_409_429#_c_507_n
+ PM_SKY130_FD_SC_LP__A221O_0%A_409_429#
x_PM_SKY130_FD_SC_LP__A221O_0%VGND N_VGND_M1003_d N_VGND_M1006_d N_VGND_c_529_n
+ N_VGND_c_530_n N_VGND_c_531_n N_VGND_c_532_n VGND N_VGND_c_533_n
+ N_VGND_c_534_n N_VGND_c_535_n PM_SKY130_FD_SC_LP__A221O_0%VGND
cc_1 VNB N_A_72_312#_M1003_g 0.0669341f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_2 VNB N_A_72_312#_c_84_n 0.00260186f $X=-0.19 $Y=-0.245 $X2=0.557 $Y2=1.677
cc_3 VNB N_A_72_312#_c_85_n 0.0144839f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.725
cc_4 VNB N_A_72_312#_c_86_n 0.0127524f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.81
cc_5 VNB N_A_72_312#_c_87_n 0.00184249f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.81
cc_6 VNB N_A_72_312#_c_88_n 0.00449019f $X=-0.19 $Y=-0.245 $X2=2.44 $Y2=0.445
cc_7 VNB N_A_72_312#_c_89_n 0.00358743f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=0.445
cc_8 VNB N_A_72_312#_c_90_n 0.00503997f $X=-0.19 $Y=-0.245 $X2=3.01 $Y2=0.73
cc_9 VNB N_A_72_312#_c_91_n 0.00655347f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=1.845
cc_10 VNB N_A_72_312#_c_92_n 0.0101943f $X=-0.19 $Y=-0.245 $X2=3.427 $Y2=0.645
cc_11 VNB N_A_72_312#_c_93_n 0.0143202f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=0.445
cc_12 VNB N_A_72_312#_c_94_n 0.0114771f $X=-0.19 $Y=-0.245 $X2=0.557 $Y2=1.56
cc_13 VNB N_A2_M1009_g 0.0275802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_207_n 0.0191971f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.74
cc_15 VNB N_A2_c_208_n 0.00920083f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.74
cc_16 VNB A2 0.00953157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_210_n 0.0148245f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_18 VNB N_A1_M1005_g 0.0278806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_252_n 0.0200048f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.23
cc_20 VNB N_A1_c_253_n 0.00301004f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.74
cc_21 VNB N_A1_c_254_n 0.0183575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB A1 0.0100717f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.725
cc_23 VNB N_A1_c_256_n 0.0177117f $X=-0.19 $Y=-0.245 $X2=0.557 $Y2=1.725
cc_24 VNB N_B1_c_298_n 0.0569452f $X=-0.19 $Y=-0.245 $X2=3.27 $Y2=0.235
cc_25 VNB N_B1_M1004_g 0.0230911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB B1 0.00398293f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.74
cc_27 VNB N_B1_c_301_n 0.0195778f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_28 VNB N_B2_M1006_g 0.0306371f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=2.145
cc_29 VNB N_B2_M1008_g 0.0138057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B2_c_336_n 0.0303478f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.74
cc_31 VNB N_B2_c_337_n 0.00730499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_C1_M1010_g 0.0380833f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=2.145
cc_33 VNB C1 0.0310147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_C1_c_372_n 0.0701232f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.74
cc_35 VNB N_X_c_401_n 0.0125155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB X 0.0359437f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.56
cc_37 VNB N_X_c_403_n 0.0137263f $X=-0.19 $Y=-0.245 $X2=3.01 $Y2=0.73
cc_38 VNB X 0.00878251f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=1.845
cc_39 VNB N_VPWR_c_426_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.81
cc_40 VNB N_VGND_c_529_n 0.00549375f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.74
cc_41 VNB N_VGND_c_530_n 0.00557617f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_42 VNB N_VGND_c_531_n 0.0416322f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.725
cc_43 VNB N_VGND_c_532_n 0.00631504f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.56
cc_44 VNB N_VGND_c_533_n 0.0219951f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.81
cc_45 VNB N_VGND_c_534_n 0.216558f $X=-0.19 $Y=-0.245 $X2=2.44 $Y2=0.445
cc_46 VNB N_VGND_c_535_n 0.0262785f $X=-0.19 $Y=-0.245 $X2=2.08 $Y2=0.445
cc_47 VPB N_A_72_312#_M1000_g 0.0245699f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_48 VPB N_A_72_312#_c_96_n 0.0257754f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.065
cc_49 VPB N_A_72_312#_c_97_n 0.0174687f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.23
cc_50 VPB N_A_72_312#_c_98_n 0.00146717f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.725
cc_51 VPB N_A_72_312#_c_85_n 0.0053288f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.725
cc_52 VPB N_A_72_312#_c_91_n 0.00322883f $X=-0.19 $Y=1.655 $X2=3.1 $Y2=1.845
cc_53 VPB N_A_72_312#_c_101_n 0.0127995f $X=-0.19 $Y=1.655 $X2=3.455 $Y2=1.93
cc_54 VPB N_A_72_312#_c_102_n 0.00322899f $X=-0.19 $Y=1.655 $X2=3.19 $Y2=1.93
cc_55 VPB N_A_72_312#_c_103_n 0.0340608f $X=-0.19 $Y=1.655 $X2=3.55 $Y2=2.29
cc_56 VPB N_A2_M1001_g 0.0516403f $X=-0.19 $Y=1.655 $X2=3.41 $Y2=2.145
cc_57 VPB N_A2_c_208_n 0.00660201f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_58 VPB N_A1_M1007_g 0.0374148f $X=-0.19 $Y=1.655 $X2=3.41 $Y2=2.145
cc_59 VPB N_A1_c_253_n 0.0162133f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_60 VPB N_A1_c_259_n 0.0175186f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.445
cc_61 VPB N_B1_c_298_n 0.0126836f $X=-0.19 $Y=1.655 $X2=3.27 $Y2=0.235
cc_62 VPB N_B1_M1002_g 0.0368249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_B2_M1008_g 0.0369157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_C1_M1011_g 0.0473306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB C1 0.00297379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_C1_c_372_n 0.00991458f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_67 VPB N_X_c_405_n 0.0366995f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_68 VPB N_X_c_401_n 0.035457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_427_n 0.0158871f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_70 VPB N_VPWR_c_428_n 0.0164339f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.445
cc_71 VPB N_VPWR_c_429_n 0.0164391f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.56
cc_72 VPB N_VPWR_c_430_n 0.0531529f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=0.81
cc_73 VPB N_VPWR_c_426_n 0.07787f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.81
cc_74 VPB N_VPWR_c_432_n 0.0244252f $X=-0.19 $Y=1.655 $X2=2.08 $Y2=0.445
cc_75 VPB N_VPWR_c_433_n 0.00564836f $X=-0.19 $Y=1.655 $X2=2.61 $Y2=0.73
cc_76 VPB N_A_216_484#_c_467_n 0.0135888f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_216_484#_c_468_n 0.0319547f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_78 VPB N_A_216_484#_c_469_n 0.00382651f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_79 VPB N_A_409_429#_c_504_n 0.0117577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_409_429#_c_505_n 0.0192652f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_81 VPB N_A_409_429#_c_506_n 0.00423633f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.74
cc_82 VPB N_A_409_429#_c_507_n 0.00101327f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.445
cc_83 N_A_72_312#_M1000_g N_A2_M1001_g 0.0130196f $X=0.555 $Y=2.74 $X2=0 $Y2=0
cc_84 N_A_72_312#_c_84_n N_A2_M1001_g 0.00228974f $X=0.557 $Y=1.677 $X2=0 $Y2=0
cc_85 N_A_72_312#_c_85_n N_A2_M1001_g 0.0292727f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_86 N_A_72_312#_M1003_g N_A2_M1009_g 0.0222137f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_72_312#_c_86_n N_A2_M1009_g 0.00972633f $X=1.2 $Y=0.81 $X2=0 $Y2=0
cc_88 N_A_72_312#_c_88_n N_A2_M1009_g 2.92591e-19 $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_72_312#_c_89_n N_A2_M1009_g 0.0112362f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_90 N_A_72_312#_c_94_n N_A2_M1009_g 0.00164599f $X=0.557 $Y=1.56 $X2=0 $Y2=0
cc_91 N_A_72_312#_c_84_n N_A2_c_208_n 4.1922e-19 $X=0.557 $Y=1.677 $X2=0 $Y2=0
cc_92 N_A_72_312#_c_85_n N_A2_c_208_n 0.00685375f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_93 N_A_72_312#_M1003_g A2 6.17778e-19 $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_72_312#_c_86_n A2 0.0230109f $X=1.2 $Y=0.81 $X2=0 $Y2=0
cc_95 N_A_72_312#_c_89_n A2 0.0142303f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_72_312#_c_94_n A2 0.0341406f $X=0.557 $Y=1.56 $X2=0 $Y2=0
cc_97 N_A_72_312#_M1003_g N_A2_c_210_n 0.0307431f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_72_312#_c_86_n N_A2_c_210_n 0.00513626f $X=1.2 $Y=0.81 $X2=0 $Y2=0
cc_99 N_A_72_312#_c_94_n N_A2_c_210_n 0.00296442f $X=0.557 $Y=1.56 $X2=0 $Y2=0
cc_100 N_A_72_312#_c_88_n N_A1_M1005_g 0.012803f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A_72_312#_c_89_n N_A1_M1005_g 0.00595778f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_102 N_A_72_312#_c_88_n A1 0.0177597f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_103 N_A_72_312#_c_89_n A1 0.00410836f $X=1.37 $Y=0.445 $X2=0 $Y2=0
cc_104 N_A_72_312#_c_88_n N_A1_c_256_n 0.00104374f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_72_312#_c_88_n N_B1_M1004_g 0.0178772f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_72_312#_c_88_n B1 0.0135958f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_72_312#_c_88_n N_B1_c_301_n 0.00149776f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_72_312#_c_88_n N_B2_M1006_g 0.0105193f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_72_312#_c_90_n N_B2_M1006_g 0.0096451f $X=3.01 $Y=0.73 $X2=0 $Y2=0
cc_110 N_A_72_312#_c_91_n N_B2_M1006_g 0.00452057f $X=3.1 $Y=1.845 $X2=0 $Y2=0
cc_111 N_A_72_312#_c_102_n N_B2_M1008_g 0.00156042f $X=3.19 $Y=1.93 $X2=0 $Y2=0
cc_112 N_A_72_312#_c_90_n N_B2_c_336_n 0.00536414f $X=3.01 $Y=0.73 $X2=0 $Y2=0
cc_113 N_A_72_312#_c_91_n N_B2_c_336_n 0.00823322f $X=3.1 $Y=1.845 $X2=0 $Y2=0
cc_114 N_A_72_312#_c_88_n N_B2_c_337_n 0.00790909f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_72_312#_c_90_n N_B2_c_337_n 0.013615f $X=3.01 $Y=0.73 $X2=0 $Y2=0
cc_116 N_A_72_312#_c_91_n N_B2_c_337_n 0.0405267f $X=3.1 $Y=1.845 $X2=0 $Y2=0
cc_117 N_A_72_312#_c_88_n N_C1_M1010_g 4.72572e-19 $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_118 N_A_72_312#_c_91_n N_C1_M1010_g 0.00969233f $X=3.1 $Y=1.845 $X2=0 $Y2=0
cc_119 N_A_72_312#_c_92_n N_C1_M1010_g 0.0155664f $X=3.427 $Y=0.645 $X2=0 $Y2=0
cc_120 N_A_72_312#_c_91_n N_C1_M1011_g 0.00439376f $X=3.1 $Y=1.845 $X2=0 $Y2=0
cc_121 N_A_72_312#_c_101_n N_C1_M1011_g 0.018657f $X=3.455 $Y=1.93 $X2=0 $Y2=0
cc_122 N_A_72_312#_c_103_n N_C1_M1011_g 0.00400853f $X=3.55 $Y=2.29 $X2=0 $Y2=0
cc_123 N_A_72_312#_c_91_n C1 0.0488536f $X=3.1 $Y=1.845 $X2=0 $Y2=0
cc_124 N_A_72_312#_c_101_n C1 0.0295574f $X=3.455 $Y=1.93 $X2=0 $Y2=0
cc_125 N_A_72_312#_c_92_n C1 0.0163584f $X=3.427 $Y=0.645 $X2=0 $Y2=0
cc_126 N_A_72_312#_c_91_n N_C1_c_372_n 0.018229f $X=3.1 $Y=1.845 $X2=0 $Y2=0
cc_127 N_A_72_312#_c_101_n N_C1_c_372_n 0.00815254f $X=3.455 $Y=1.93 $X2=0 $Y2=0
cc_128 N_A_72_312#_c_92_n N_C1_c_372_n 0.00925866f $X=3.427 $Y=0.645 $X2=0 $Y2=0
cc_129 N_A_72_312#_M1000_g N_X_c_405_n 8.31719e-19 $X=0.555 $Y=2.74 $X2=0 $Y2=0
cc_130 N_A_72_312#_c_97_n N_X_c_405_n 0.00411556f $X=0.525 $Y=2.23 $X2=0 $Y2=0
cc_131 N_A_72_312#_c_98_n N_X_c_405_n 0.00293724f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_132 N_A_72_312#_M1000_g N_X_c_401_n 0.00557933f $X=0.555 $Y=2.74 $X2=0 $Y2=0
cc_133 N_A_72_312#_M1003_g N_X_c_401_n 0.00112021f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_134 N_A_72_312#_c_84_n N_X_c_401_n 0.0491882f $X=0.557 $Y=1.677 $X2=0 $Y2=0
cc_135 N_A_72_312#_c_85_n N_X_c_401_n 0.0164925f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_136 N_A_72_312#_c_94_n N_X_c_401_n 0.0101928f $X=0.557 $Y=1.56 $X2=0 $Y2=0
cc_137 N_A_72_312#_M1003_g X 0.00944256f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_138 N_A_72_312#_c_87_n X 0.014748f $X=0.675 $Y=0.81 $X2=0 $Y2=0
cc_139 N_A_72_312#_c_94_n X 0.0382518f $X=0.557 $Y=1.56 $X2=0 $Y2=0
cc_140 N_A_72_312#_M1003_g N_X_c_403_n 0.00346132f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A_72_312#_c_87_n N_X_c_403_n 0.00206954f $X=0.675 $Y=0.81 $X2=0 $Y2=0
cc_142 N_A_72_312#_M1000_g N_VPWR_c_427_n 0.00301473f $X=0.555 $Y=2.74 $X2=0
+ $Y2=0
cc_143 N_A_72_312#_c_97_n N_VPWR_c_427_n 9.86952e-19 $X=0.525 $Y=2.23 $X2=0
+ $Y2=0
cc_144 N_A_72_312#_c_98_n N_VPWR_c_427_n 0.00249633f $X=0.525 $Y=1.725 $X2=0
+ $Y2=0
cc_145 N_A_72_312#_c_103_n N_VPWR_c_430_n 0.00653432f $X=3.55 $Y=2.29 $X2=0
+ $Y2=0
cc_146 N_A_72_312#_M1000_g N_VPWR_c_426_n 0.0112317f $X=0.555 $Y=2.74 $X2=0
+ $Y2=0
cc_147 N_A_72_312#_c_103_n N_VPWR_c_426_n 0.00842003f $X=3.55 $Y=2.29 $X2=0
+ $Y2=0
cc_148 N_A_72_312#_M1000_g N_VPWR_c_432_n 0.00550375f $X=0.555 $Y=2.74 $X2=0
+ $Y2=0
cc_149 N_A_72_312#_c_98_n N_A_216_484#_c_467_n 0.0105339f $X=0.525 $Y=1.725
+ $X2=0 $Y2=0
cc_150 N_A_72_312#_c_91_n N_A_216_484#_c_468_n 0.00386331f $X=3.1 $Y=1.845 $X2=0
+ $Y2=0
cc_151 N_A_72_312#_c_102_n N_A_216_484#_c_468_n 0.00795763f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_152 N_A_72_312#_c_98_n N_A_216_484#_c_469_n 0.0071287f $X=0.525 $Y=1.725
+ $X2=0 $Y2=0
cc_153 N_A_72_312#_c_102_n N_A_216_484#_c_474_n 0.00408414f $X=3.19 $Y=1.93
+ $X2=0 $Y2=0
cc_154 N_A_72_312#_c_103_n N_A_216_484#_c_474_n 0.00395446f $X=3.55 $Y=2.29
+ $X2=0 $Y2=0
cc_155 N_A_72_312#_c_101_n N_A_409_429#_c_507_n 0.00497828f $X=3.455 $Y=1.93
+ $X2=0 $Y2=0
cc_156 N_A_72_312#_c_102_n N_A_409_429#_c_507_n 0.0165005f $X=3.19 $Y=1.93 $X2=0
+ $Y2=0
cc_157 N_A_72_312#_c_103_n N_A_409_429#_c_507_n 0.0232498f $X=3.55 $Y=2.29 $X2=0
+ $Y2=0
cc_158 N_A_72_312#_c_90_n N_VGND_M1006_d 0.00228741f $X=3.01 $Y=0.73 $X2=0 $Y2=0
cc_159 N_A_72_312#_c_92_n N_VGND_M1006_d 5.42526e-19 $X=3.427 $Y=0.645 $X2=0
+ $Y2=0
cc_160 N_A_72_312#_M1003_g N_VGND_c_529_n 0.00498814f $X=0.585 $Y=0.445 $X2=0
+ $Y2=0
cc_161 N_A_72_312#_c_86_n N_VGND_c_529_n 0.0245582f $X=1.2 $Y=0.81 $X2=0 $Y2=0
cc_162 N_A_72_312#_c_90_n N_VGND_c_530_n 0.021074f $X=3.01 $Y=0.73 $X2=0 $Y2=0
cc_163 N_A_72_312#_c_86_n N_VGND_c_531_n 0.00235592f $X=1.2 $Y=0.81 $X2=0 $Y2=0
cc_164 N_A_72_312#_c_88_n N_VGND_c_531_n 0.0628771f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A_72_312#_c_89_n N_VGND_c_531_n 0.00837801f $X=1.37 $Y=0.445 $X2=0
+ $Y2=0
cc_166 N_A_72_312#_c_90_n N_VGND_c_531_n 0.00238193f $X=3.01 $Y=0.73 $X2=0 $Y2=0
cc_167 N_A_72_312#_c_92_n N_VGND_c_533_n 0.00260208f $X=3.427 $Y=0.645 $X2=0
+ $Y2=0
cc_168 N_A_72_312#_c_93_n N_VGND_c_533_n 0.0157815f $X=3.41 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_72_312#_M1005_d N_VGND_c_534_n 0.00518052f $X=1.59 $Y=0.235 $X2=0
+ $Y2=0
cc_170 N_A_72_312#_M1010_d N_VGND_c_534_n 0.00220958f $X=3.27 $Y=0.235 $X2=0
+ $Y2=0
cc_171 N_A_72_312#_M1003_g N_VGND_c_534_n 0.00743784f $X=0.585 $Y=0.445 $X2=0
+ $Y2=0
cc_172 N_A_72_312#_c_86_n N_VGND_c_534_n 0.00618208f $X=1.2 $Y=0.81 $X2=0 $Y2=0
cc_173 N_A_72_312#_c_87_n N_VGND_c_534_n 0.00338644f $X=0.675 $Y=0.81 $X2=0
+ $Y2=0
cc_174 N_A_72_312#_c_88_n N_VGND_c_534_n 0.0451312f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_175 N_A_72_312#_c_89_n N_VGND_c_534_n 0.00629885f $X=1.37 $Y=0.445 $X2=0
+ $Y2=0
cc_176 N_A_72_312#_c_90_n N_VGND_c_534_n 0.00565529f $X=3.01 $Y=0.73 $X2=0 $Y2=0
cc_177 N_A_72_312#_c_92_n N_VGND_c_534_n 0.00408341f $X=3.427 $Y=0.645 $X2=0
+ $Y2=0
cc_178 N_A_72_312#_c_93_n N_VGND_c_534_n 0.0110631f $X=3.41 $Y=0.445 $X2=0 $Y2=0
cc_179 N_A_72_312#_M1003_g N_VGND_c_535_n 0.00425274f $X=0.585 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_72_312#_c_86_n N_VGND_c_535_n 5.92998e-19 $X=1.2 $Y=0.81 $X2=0 $Y2=0
cc_181 N_A_72_312#_c_87_n N_VGND_c_535_n 0.00209494f $X=0.675 $Y=0.81 $X2=0
+ $Y2=0
cc_182 N_A_72_312#_c_88_n A_246_47# 0.00145479f $X=2.44 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_72_312#_c_89_n A_246_47# 0.00212597f $X=1.37 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_72_312#_c_88_n A_474_47# 0.00357715f $X=2.44 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A2_M1009_g N_A1_M1005_g 0.0246053f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A2_c_207_n N_A1_c_252_n 0.0246053f $X=1.065 $Y=1.5 $X2=0 $Y2=0
cc_187 N_A2_M1001_g N_A1_c_253_n 0.00819952f $X=1.005 $Y=2.74 $X2=0 $Y2=0
cc_188 N_A2_M1001_g N_A1_c_259_n 0.024502f $X=1.005 $Y=2.74 $X2=0 $Y2=0
cc_189 N_A2_c_208_n N_A1_c_254_n 0.0246053f $X=1.065 $Y=1.665 $X2=0 $Y2=0
cc_190 N_A2_M1009_g A1 9.72558e-19 $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_191 A2 A1 0.0418529f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A2_c_210_n A1 4.50775e-19 $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_193 A2 N_A1_c_256_n 0.00414812f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A2_c_210_n N_A1_c_256_n 0.0246053f $X=1.065 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A2_M1001_g N_VPWR_c_427_n 0.00177492f $X=1.005 $Y=2.74 $X2=0 $Y2=0
cc_196 N_A2_M1001_g N_VPWR_c_429_n 0.00550375f $X=1.005 $Y=2.74 $X2=0 $Y2=0
cc_197 N_A2_M1001_g N_VPWR_c_426_n 0.0104172f $X=1.005 $Y=2.74 $X2=0 $Y2=0
cc_198 N_A2_M1001_g N_A_216_484#_c_467_n 0.00814125f $X=1.005 $Y=2.74 $X2=0
+ $Y2=0
cc_199 A2 N_A_216_484#_c_468_n 7.88607e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_200 N_A2_M1001_g N_A_216_484#_c_469_n 0.00248817f $X=1.005 $Y=2.74 $X2=0
+ $Y2=0
cc_201 N_A2_c_208_n N_A_216_484#_c_469_n 0.00390321f $X=1.065 $Y=1.665 $X2=0
+ $Y2=0
cc_202 A2 N_A_216_484#_c_469_n 0.0228155f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A2_M1009_g N_VGND_c_529_n 0.0050379f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_204 N_A2_M1009_g N_VGND_c_531_n 0.00424336f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A2_M1009_g N_VGND_c_534_n 0.00612198f $X=1.155 $Y=0.445 $X2=0 $Y2=0
cc_206 N_A1_c_252_n N_B1_c_298_n 0.0180191f $X=1.62 $Y=1.425 $X2=0 $Y2=0
cc_207 N_A1_c_253_n N_B1_c_298_n 0.00435082f $X=1.515 $Y=1.905 $X2=0 $Y2=0
cc_208 N_A1_c_254_n N_B1_c_298_n 0.0025806f $X=1.62 $Y=1.605 $X2=0 $Y2=0
cc_209 A1 N_B1_c_298_n 0.00109745f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_210 N_A1_M1005_g N_B1_M1004_g 0.00741301f $X=1.515 $Y=0.445 $X2=0 $Y2=0
cc_211 A1 B1 0.0516466f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_212 N_A1_c_256_n B1 6.49729e-19 $X=1.635 $Y=1.1 $X2=0 $Y2=0
cc_213 N_A1_M1005_g N_B1_c_301_n 0.00227833f $X=1.515 $Y=0.445 $X2=0 $Y2=0
cc_214 A1 N_B1_c_301_n 0.00407286f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_215 N_A1_c_256_n N_B1_c_301_n 0.0180191f $X=1.635 $Y=1.1 $X2=0 $Y2=0
cc_216 A1 N_B2_c_337_n 0.002386f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_217 N_A1_M1007_g N_VPWR_c_428_n 0.00386163f $X=1.435 $Y=2.74 $X2=0 $Y2=0
cc_218 N_A1_c_259_n N_VPWR_c_428_n 0.00174455f $X=1.515 $Y=1.98 $X2=0 $Y2=0
cc_219 N_A1_M1007_g N_VPWR_c_429_n 0.00550375f $X=1.435 $Y=2.74 $X2=0 $Y2=0
cc_220 N_A1_M1007_g N_VPWR_c_426_n 0.0114216f $X=1.435 $Y=2.74 $X2=0 $Y2=0
cc_221 N_A1_c_259_n N_A_216_484#_c_467_n 0.00918611f $X=1.515 $Y=1.98 $X2=0
+ $Y2=0
cc_222 N_A1_c_253_n N_A_216_484#_c_468_n 0.0111776f $X=1.515 $Y=1.905 $X2=0
+ $Y2=0
cc_223 N_A1_c_259_n N_A_216_484#_c_468_n 0.0121385f $X=1.515 $Y=1.98 $X2=0 $Y2=0
cc_224 N_A1_c_254_n N_A_216_484#_c_468_n 0.00144471f $X=1.62 $Y=1.605 $X2=0
+ $Y2=0
cc_225 A1 N_A_216_484#_c_468_n 0.0232012f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_226 N_A1_M1007_g N_A_409_429#_c_504_n 0.00512799f $X=1.435 $Y=2.74 $X2=0
+ $Y2=0
cc_227 N_A1_M1005_g N_VGND_c_531_n 0.00363059f $X=1.515 $Y=0.445 $X2=0 $Y2=0
cc_228 N_A1_M1005_g N_VGND_c_534_n 0.00596462f $X=1.515 $Y=0.445 $X2=0 $Y2=0
cc_229 N_B1_M1004_g N_B2_M1006_g 0.0402178f $X=2.295 $Y=0.445 $X2=0 $Y2=0
cc_230 B1 N_B2_M1006_g 0.00111454f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_231 N_B1_c_298_n N_B2_M1008_g 0.0362757f $X=2.19 $Y=1.33 $X2=0 $Y2=0
cc_232 B1 N_B2_c_336_n 3.05971e-19 $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_233 N_B1_c_301_n N_B2_c_336_n 0.0402178f $X=2.175 $Y=1.005 $X2=0 $Y2=0
cc_234 N_B1_c_298_n N_B2_c_337_n 0.00461423f $X=2.19 $Y=1.33 $X2=0 $Y2=0
cc_235 B1 N_B2_c_337_n 0.0291124f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_236 N_B1_M1002_g N_VPWR_c_428_n 7.86472e-19 $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B1_M1002_g N_VPWR_c_430_n 6.36823e-19 $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B1_c_298_n N_A_216_484#_c_468_n 0.00694611f $X=2.19 $Y=1.33 $X2=0 $Y2=0
cc_239 N_B1_M1002_g N_A_216_484#_c_468_n 0.020021f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_240 B1 N_A_216_484#_c_468_n 0.0140557f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_241 N_B1_M1002_g N_A_216_484#_c_474_n 0.016689f $X=2.405 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B1_M1002_g N_A_409_429#_c_504_n 0.0037363f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_243 N_B1_M1002_g N_A_409_429#_c_505_n 0.00895017f $X=2.405 $Y=2.465 $X2=0
+ $Y2=0
cc_244 N_B1_M1004_g N_VGND_c_531_n 0.00363059f $X=2.295 $Y=0.445 $X2=0 $Y2=0
cc_245 N_B1_M1004_g N_VGND_c_534_n 0.00596462f $X=2.295 $Y=0.445 $X2=0 $Y2=0
cc_246 N_B2_M1006_g N_C1_M1010_g 0.0217404f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_247 N_B2_M1008_g N_C1_M1011_g 0.0257186f $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B2_c_336_n N_C1_c_372_n 0.0372142f $X=2.745 $Y=1.215 $X2=0 $Y2=0
cc_249 N_B2_c_337_n N_C1_c_372_n 4.7794e-19 $X=2.745 $Y=1.215 $X2=0 $Y2=0
cc_250 N_B2_M1008_g N_VPWR_c_430_n 6.36823e-19 $X=2.835 $Y=2.465 $X2=0 $Y2=0
cc_251 N_B2_M1008_g N_A_216_484#_c_468_n 0.00434687f $X=2.835 $Y=2.465 $X2=0
+ $Y2=0
cc_252 N_B2_c_336_n N_A_216_484#_c_468_n 8.91778e-19 $X=2.745 $Y=1.215 $X2=0
+ $Y2=0
cc_253 N_B2_c_337_n N_A_216_484#_c_468_n 0.0234627f $X=2.745 $Y=1.215 $X2=0
+ $Y2=0
cc_254 N_B2_M1008_g N_A_216_484#_c_474_n 0.0122237f $X=2.835 $Y=2.465 $X2=0
+ $Y2=0
cc_255 N_B2_M1008_g N_A_409_429#_c_505_n 0.00889096f $X=2.835 $Y=2.465 $X2=0
+ $Y2=0
cc_256 N_B2_M1008_g N_A_409_429#_c_507_n 0.00498904f $X=2.835 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_B2_M1006_g N_VGND_c_530_n 0.00444512f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_258 N_B2_M1006_g N_VGND_c_531_n 0.00415306f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_259 N_B2_M1006_g N_VGND_c_534_n 0.00590165f $X=2.655 $Y=0.445 $X2=0 $Y2=0
cc_260 N_C1_M1011_g N_VPWR_c_430_n 0.00393989f $X=3.335 $Y=2.465 $X2=0 $Y2=0
cc_261 N_C1_M1011_g N_VPWR_c_426_n 0.00410091f $X=3.335 $Y=2.465 $X2=0 $Y2=0
cc_262 N_C1_M1011_g N_A_216_484#_c_474_n 4.87801e-19 $X=3.335 $Y=2.465 $X2=0
+ $Y2=0
cc_263 N_C1_M1011_g N_A_409_429#_c_505_n 0.0010503f $X=3.335 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_C1_M1011_g N_A_409_429#_c_507_n 0.0129833f $X=3.335 $Y=2.465 $X2=0
+ $Y2=0
cc_265 N_C1_c_372_n N_A_409_429#_c_507_n 2.98189e-19 $X=3.445 $Y=1.16 $X2=0
+ $Y2=0
cc_266 N_C1_M1010_g N_VGND_c_530_n 0.00334823f $X=3.195 $Y=0.445 $X2=0 $Y2=0
cc_267 N_C1_M1010_g N_VGND_c_533_n 0.00426565f $X=3.195 $Y=0.445 $X2=0 $Y2=0
cc_268 N_C1_M1010_g N_VGND_c_534_n 0.00713854f $X=3.195 $Y=0.445 $X2=0 $Y2=0
cc_269 N_X_c_405_n N_VPWR_c_427_n 0.00274452f $X=0.34 $Y=2.565 $X2=0 $Y2=0
cc_270 N_X_c_405_n N_VPWR_c_426_n 0.0148886f $X=0.34 $Y=2.565 $X2=0 $Y2=0
cc_271 N_X_c_405_n N_VPWR_c_432_n 0.0274478f $X=0.34 $Y=2.565 $X2=0 $Y2=0
cc_272 N_X_M1003_s N_VGND_c_534_n 0.0021695f $X=0.245 $Y=0.235 $X2=0 $Y2=0
cc_273 N_X_c_403_n N_VGND_c_534_n 0.0165448f $X=0.37 $Y=0.445 $X2=0 $Y2=0
cc_274 N_X_c_403_n N_VGND_c_535_n 0.0237759f $X=0.37 $Y=0.445 $X2=0 $Y2=0
cc_275 N_VPWR_c_427_n N_A_216_484#_c_467_n 0.00265959f $X=0.79 $Y=2.565 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_428_n N_A_216_484#_c_467_n 0.00267021f $X=1.65 $Y=2.565 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_429_n N_A_216_484#_c_467_n 0.0181367f $X=1.52 $Y=3.33 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_426_n N_A_216_484#_c_467_n 0.00983606f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_428_n N_A_216_484#_c_468_n 0.0124288f $X=1.65 $Y=2.565 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_428_n N_A_409_429#_c_504_n 0.0380441f $X=1.65 $Y=2.565 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_430_n N_A_409_429#_c_505_n 0.0667586f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_282 N_VPWR_c_426_n N_A_409_429#_c_505_n 0.0380121f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_283 N_VPWR_c_428_n N_A_409_429#_c_506_n 0.0137896f $X=1.65 $Y=2.565 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_430_n N_A_409_429#_c_506_n 0.0200723f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_285 N_VPWR_c_426_n N_A_409_429#_c_506_n 0.0108858f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_286 N_A_216_484#_c_467_n N_A_409_429#_c_504_n 0.00824056f $X=1.22 $Y=2.545
+ $X2=0 $Y2=0
cc_287 N_A_216_484#_c_468_n N_A_409_429#_c_504_n 0.0225468f $X=2.455 $Y=1.87
+ $X2=0 $Y2=0
cc_288 N_A_216_484#_c_474_n N_A_409_429#_c_504_n 0.0228787f $X=2.62 $Y=2.27
+ $X2=0 $Y2=0
cc_289 N_A_216_484#_c_474_n N_A_409_429#_c_505_n 0.0205115f $X=2.62 $Y=2.27
+ $X2=0 $Y2=0
cc_290 N_VGND_c_534_n A_246_47# 0.0016882f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_291 N_VGND_c_534_n A_474_47# 0.0016882f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
