# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrbn_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrbn_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.090000 0.835000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.402600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.510000 0.745000 7.875000 1.180000 ;
        RECT 7.510000 1.180000 8.055000 1.205000 ;
        RECT 7.705000 1.205000 8.055000 3.065000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.402600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.380000 1.850000 9.970000 2.890000 ;
        RECT 9.640000 0.360000 9.970000 0.820000 ;
        RECT 9.800000 0.820000 9.970000 1.850000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.335000 1.605000 6.665000 2.520000 ;
    END
  END RESET_B
  PIN GATE_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.085000 0.960000 1.500000 1.780000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
        RECT 0.905000  0.085000  1.235000 0.780000 ;
        RECT 3.045000  0.085000  3.375000 0.675000 ;
        RECT 5.345000  0.085000  5.675000 0.425000 ;
        RECT 6.720000  0.085000  7.050000 1.075000 ;
        RECT 8.850000  0.085000  9.180000 0.820000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
        RECT 9.275000 -0.085000 9.445000 0.085000 ;
        RECT 9.755000 -0.085000 9.925000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.080000 3.415000 ;
        RECT 0.705000 2.740000  1.035000 3.245000 ;
        RECT 3.015000 2.405000  3.265000 3.245000 ;
        RECT 4.985000 2.385000  5.315000 3.245000 ;
        RECT 7.195000 2.075000  7.525000 3.245000 ;
        RECT 8.850000 1.850000  9.180000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
        RECT 9.275000 3.245000 9.445000 3.415000 ;
        RECT 9.755000 3.245000 9.925000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.320000 0.445000 0.780000 ;
      RECT 0.090000 0.780000 0.260000 1.960000 ;
      RECT 0.090000 1.960000 0.505000 2.390000 ;
      RECT 0.090000 2.390000 1.385000 2.560000 ;
      RECT 0.090000 2.560000 0.505000 3.000000 ;
      RECT 1.215000 2.560000 1.385000 2.895000 ;
      RECT 1.215000 2.895000 2.835000 3.065000 ;
      RECT 1.235000 1.960000 1.965000 2.210000 ;
      RECT 1.695000 0.320000 1.965000 1.960000 ;
      RECT 1.695000 2.210000 1.965000 2.630000 ;
      RECT 2.145000 0.265000 2.585000 0.675000 ;
      RECT 2.145000 0.675000 2.315000 1.705000 ;
      RECT 2.145000 1.705000 3.045000 1.875000 ;
      RECT 2.145000 1.875000 2.485000 2.715000 ;
      RECT 2.495000 0.855000 4.360000 1.025000 ;
      RECT 2.495000 1.025000 2.695000 1.525000 ;
      RECT 2.665000 2.055000 3.490000 2.225000 ;
      RECT 2.665000 2.225000 2.835000 2.895000 ;
      RECT 2.875000 1.255000 3.850000 1.425000 ;
      RECT 2.875000 1.425000 3.045000 1.705000 ;
      RECT 3.225000 1.605000 3.490000 2.055000 ;
      RECT 3.680000 1.425000 4.770000 1.595000 ;
      RECT 3.680000 1.595000 4.030000 1.755000 ;
      RECT 3.965000 2.035000 5.645000 2.205000 ;
      RECT 3.965000 2.205000 4.295000 3.065000 ;
      RECT 4.030000 1.025000 4.360000 1.185000 ;
      RECT 4.295000 0.265000 4.710000 0.605000 ;
      RECT 4.295000 0.605000 6.185000 0.675000 ;
      RECT 4.540000 0.675000 6.185000 0.775000 ;
      RECT 4.600000 0.955000 4.930000 1.285000 ;
      RECT 4.600000 1.285000 4.770000 1.425000 ;
      RECT 4.965000 1.525000 5.295000 1.855000 ;
      RECT 5.125000 0.955000 6.260000 1.205000 ;
      RECT 5.125000 1.205000 5.295000 1.525000 ;
      RECT 5.475000 1.565000 5.890000 1.895000 ;
      RECT 5.475000 1.895000 5.645000 2.035000 ;
      RECT 5.825000 2.075000 6.155000 2.700000 ;
      RECT 5.825000 2.700000 7.015000 2.870000 ;
      RECT 5.825000 2.870000 6.155000 3.065000 ;
      RECT 5.855000 0.325000 6.185000 0.605000 ;
      RECT 6.090000 1.205000 6.260000 1.255000 ;
      RECT 6.090000 1.255000 7.330000 1.425000 ;
      RECT 6.845000 1.425000 7.330000 1.625000 ;
      RECT 6.845000 1.625000 7.015000 2.700000 ;
      RECT 8.060000 0.360000 8.405000 0.820000 ;
      RECT 8.235000 0.820000 8.405000 1.000000 ;
      RECT 8.235000 1.000000 9.485000 1.170000 ;
      RECT 8.235000 1.170000 8.650000 2.890000 ;
      RECT 9.155000 1.170000 9.485000 1.670000 ;
  END
END sky130_fd_sc_lp__dlrbn_lp
