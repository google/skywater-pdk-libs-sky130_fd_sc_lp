* File: sky130_fd_sc_lp__o2111ai_0.spice
* Created: Fri Aug 28 11:00:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111ai_0.pex.spice"
.subckt sky130_fd_sc_lp__o2111ai_0  VNB VPB D1 C1 B1 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1006 A_195_47# N_D1_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.2541 PD=0.63 PS=2.05 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.5 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1007 A_267_47# N_C1_M1007_g A_195_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.9 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_339_47#_M1009_d N_B1_M1009_g A_267_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0441 PD=1.04 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_339_47#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1302 PD=0.7 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_339_47#_M1004_d N_A1_M1004_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_D1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_C1_M1000_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.3072 AS=0.0896 PD=1.6 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1056 AS=0.3072 PD=0.97 PS=1.6 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1005 A_520_465# N_A2_M1005_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.1056 PD=0.85 PS=0.97 NRD=15.3857 NRS=15.3857 M=1 R=4.26667 SA=75002.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_520_465# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75002.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o2111ai_0.pxi.spice"
*
.ends
*
*
