* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__invlp_8 A VGND VNB VPB VPWR Y
X0 Y A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_114_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_114_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_114_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 Y A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_114_367# A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_114_367# A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VPWR A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_114_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 Y A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_114_53# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_114_53# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_114_367# A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Y A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_114_53# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 Y A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_114_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VPWR A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 a_114_367# A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_114_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 Y A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VGND A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 Y A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 VPWR A a_114_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VGND A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X28 a_114_53# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 a_114_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 a_114_53# A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X31 Y A a_114_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
