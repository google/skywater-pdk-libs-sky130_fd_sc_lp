# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__mux4_m
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__mux4_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.315000 1.160000 4.645000 1.490000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.470000 3.235000 1.980000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 1.485000 1.285000 2.860000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.365000 1.470000 2.725000 1.980000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 0.265000 0.675000 0.435000 ;
        RECT 0.155000 0.435000 0.325000 0.640000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.795000 0.840000 7.125000 1.355000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.795000 0.345000 8.005000 2.945000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 8.160000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 8.350000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.315000  0.820000 0.700000 1.135000 ;
      RECT 0.315000  1.135000 1.825000 1.305000 ;
      RECT 0.315000  1.305000 0.525000 2.625000 ;
      RECT 0.745000  2.425000 0.935000 3.245000 ;
      RECT 0.880000  0.085000 1.210000 0.880000 ;
      RECT 1.520000  0.275000 2.525000 0.445000 ;
      RECT 1.520000  0.445000 1.690000 1.135000 ;
      RECT 1.520000  1.305000 1.825000 1.830000 ;
      RECT 1.760000  2.175000 3.175000 2.345000 ;
      RECT 1.760000  2.345000 2.005000 2.625000 ;
      RECT 1.870000  0.625000 2.175000 0.955000 ;
      RECT 2.005000  0.955000 2.175000 2.175000 ;
      RECT 2.355000  0.445000 2.525000 1.100000 ;
      RECT 2.355000  1.100000 3.695000 1.270000 ;
      RECT 2.495000  2.525000 2.825000 3.245000 ;
      RECT 2.705000  0.085000 2.895000 0.920000 ;
      RECT 3.005000  2.345000 3.175000 2.745000 ;
      RECT 3.005000  2.745000 4.395000 2.915000 ;
      RECT 3.415000  0.710000 4.045000 0.920000 ;
      RECT 3.525000  1.270000 3.695000 1.880000 ;
      RECT 3.570000  2.355000 4.045000 2.565000 ;
      RECT 3.875000  0.920000 4.045000 1.725000 ;
      RECT 3.875000  1.725000 5.445000 1.895000 ;
      RECT 3.875000  1.895000 4.045000 2.355000 ;
      RECT 4.225000  2.075000 5.095000 2.245000 ;
      RECT 4.225000  2.245000 4.395000 2.745000 ;
      RECT 4.265000  0.085000 4.475000 0.940000 ;
      RECT 4.575000  2.425000 4.745000 3.245000 ;
      RECT 4.925000  2.245000 5.095000 2.805000 ;
      RECT 4.925000  2.805000 6.595000 2.975000 ;
      RECT 5.255000  0.965000 5.445000 1.725000 ;
      RECT 5.275000  1.895000 5.445000 2.625000 ;
      RECT 5.590000  0.265000 7.145000 0.435000 ;
      RECT 5.625000  0.615000 6.595000 0.785000 ;
      RECT 5.625000  0.785000 5.795000 2.805000 ;
      RECT 5.975000  0.965000 6.165000 1.535000 ;
      RECT 5.975000  1.535000 7.615000 1.705000 ;
      RECT 5.975000  1.705000 6.165000 2.625000 ;
      RECT 6.345000  1.885000 7.145000 2.055000 ;
      RECT 6.385000  0.785000 6.595000 1.165000 ;
      RECT 6.385000  2.425000 6.595000 2.805000 ;
      RECT 6.935000  0.435000 7.145000 0.595000 ;
      RECT 6.935000  2.055000 7.145000 2.945000 ;
      RECT 7.365000  2.745000 7.575000 3.245000 ;
      RECT 7.385000  0.085000 7.575000 0.545000 ;
      RECT 7.445000  1.190000 7.615000 1.535000 ;
      RECT 7.445000  1.705000 7.615000 1.860000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__mux4_m
END LIBRARY
