* File: sky130_fd_sc_lp__o22ai_4.pex.spice
* Created: Wed Sep  2 10:20:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22AI_4%A1 3 7 11 15 19 23 27 31 33 42 43 49 50 52
+ 53 54 55 56 57 73
c133 52 0 1.60411e-19 $X=3.385 $Y=2.035
r134 72 73 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.365 $Y=1.46
+ $X2=1.38 $Y2=1.46
r135 69 70 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.935 $Y=1.46
+ $X2=0.95 $Y2=1.46
r136 66 67 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.505 $Y=1.46
+ $X2=0.52 $Y2=1.46
r137 56 57 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=2.035
+ $X2=3.12 $Y2=2.035
r138 55 56 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.035
+ $X2=2.64 $Y2=2.035
r139 54 55 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=2.16 $Y2=2.035
r140 54 78 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=1.455 $Y2=2.035
r141 53 78 6.18617 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.24 $Y=2.035
+ $X2=1.455 $Y2=2.035
r142 52 57 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=2.035
+ $X2=3.12 $Y2=2.035
r143 50 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=1.44
+ $X2=3.55 $Y2=1.605
r144 50 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.55 $Y=1.44
+ $X2=3.55 $Y2=1.275
r145 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.44 $X2=3.55 $Y2=1.44
r146 46 72 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=1.46
+ $X2=1.365 $Y2=1.46
r147 46 70 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.29 $Y=1.46
+ $X2=0.95 $Y2=1.46
r148 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.29
+ $Y=1.46 $X2=1.29 $Y2=1.46
r149 43 53 7.01894 $w=5.98e-07 $l=3.2e-07 $layer=LI1_cond $X=1.24 $Y=1.63
+ $X2=1.24 $Y2=1.95
r150 43 45 2.87101 $w=4.3e-07 $l=1.43e-07 $layer=LI1_cond $X=1.24 $Y=1.63
+ $X2=1.24 $Y2=1.487
r151 42 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=1.95
+ $X2=3.385 $Y2=2.035
r152 41 49 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.47 $Y=1.525 $X2=3.47
+ $Y2=1.435
r153 41 42 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.47 $Y=1.525
+ $X2=3.47 $Y2=1.95
r154 40 69 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=0.61 $Y=1.46
+ $X2=0.935 $Y2=1.46
r155 40 67 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.61 $Y=1.46 $X2=0.52
+ $Y2=1.46
r156 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.46 $X2=0.61 $Y2=1.46
r157 36 66 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.505 $Y2=1.46
r158 35 39 13.7484 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.27 $Y=1.487
+ $X2=0.61 $Y2=1.487
r159 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.46 $X2=0.27 $Y2=1.46
r160 33 45 4.31656 $w=2.85e-07 $l=2.15e-07 $layer=LI1_cond $X=1.025 $Y=1.487
+ $X2=1.24 $Y2=1.487
r161 33 39 16.7812 $w=2.83e-07 $l=4.15e-07 $layer=LI1_cond $X=1.025 $Y=1.487
+ $X2=0.61 $Y2=1.487
r162 31 77 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.53 $Y=2.465
+ $X2=3.53 $Y2=1.605
r163 27 76 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.515 $Y=0.655
+ $X2=3.515 $Y2=1.275
r164 21 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.625
+ $X2=1.38 $Y2=1.46
r165 21 23 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.38 $Y=1.625
+ $X2=1.38 $Y2=2.465
r166 17 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.365 $Y=1.295
+ $X2=1.365 $Y2=1.46
r167 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.365 $Y=1.295
+ $X2=1.365 $Y2=0.655
r168 13 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.625
+ $X2=0.95 $Y2=1.46
r169 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.95 $Y=1.625
+ $X2=0.95 $Y2=2.465
r170 9 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.295
+ $X2=0.935 $Y2=1.46
r171 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.935 $Y=1.295
+ $X2=0.935 $Y2=0.655
r172 5 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.625
+ $X2=0.52 $Y2=1.46
r173 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.52 $Y=1.625
+ $X2=0.52 $Y2=2.465
r174 1 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.295
+ $X2=0.505 $Y2=1.46
r175 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.505 $Y=1.295
+ $X2=0.505 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_4%A2 3 7 11 15 19 23 27 31 33 34 35 51
c85 51 0 6.80066e-20 $X=3.085 $Y=1.51
r86 51 52 2.20427 $w=3.28e-07 $l=1.5e-08 $layer=POLY_cond $X=3.085 $Y=1.51
+ $X2=3.1 $Y2=1.51
r87 49 51 13.2256 $w=3.28e-07 $l=9e-08 $layer=POLY_cond $X=2.995 $Y=1.51
+ $X2=3.085 $Y2=1.51
r88 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.995
+ $Y=1.51 $X2=2.995 $Y2=1.51
r89 47 49 47.7591 $w=3.28e-07 $l=3.25e-07 $layer=POLY_cond $X=2.67 $Y=1.51
+ $X2=2.995 $Y2=1.51
r90 46 47 2.20427 $w=3.28e-07 $l=1.5e-08 $layer=POLY_cond $X=2.655 $Y=1.51
+ $X2=2.67 $Y2=1.51
r91 45 46 60.9848 $w=3.28e-07 $l=4.15e-07 $layer=POLY_cond $X=2.24 $Y=1.51
+ $X2=2.655 $Y2=1.51
r92 44 45 2.20427 $w=3.28e-07 $l=1.5e-08 $layer=POLY_cond $X=2.225 $Y=1.51
+ $X2=2.24 $Y2=1.51
r93 42 44 36.7378 $w=3.28e-07 $l=2.5e-07 $layer=POLY_cond $X=1.975 $Y=1.51
+ $X2=2.225 $Y2=1.51
r94 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.975
+ $Y=1.51 $X2=1.975 $Y2=1.51
r95 40 42 24.247 $w=3.28e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.51
+ $X2=1.975 $Y2=1.51
r96 39 40 2.20427 $w=3.28e-07 $l=1.5e-08 $layer=POLY_cond $X=1.795 $Y=1.51
+ $X2=1.81 $Y2=1.51
r97 35 50 3.55692 $w=4.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.12 $Y=1.547
+ $X2=2.995 $Y2=1.547
r98 34 50 10.1017 $w=4.03e-07 $l=3.55e-07 $layer=LI1_cond $X=2.64 $Y=1.547
+ $X2=2.995 $Y2=1.547
r99 33 34 13.6586 $w=4.03e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.547
+ $X2=2.64 $Y2=1.547
r100 33 43 5.26425 $w=4.03e-07 $l=1.85e-07 $layer=LI1_cond $X=2.16 $Y=1.547
+ $X2=1.975 $Y2=1.547
r101 29 52 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.1 $Y=1.675
+ $X2=3.1 $Y2=1.51
r102 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.1 $Y=1.675
+ $X2=3.1 $Y2=2.465
r103 25 51 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.345
+ $X2=3.085 $Y2=1.51
r104 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.085 $Y=1.345
+ $X2=3.085 $Y2=0.655
r105 21 47 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.675
+ $X2=2.67 $Y2=1.51
r106 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.67 $Y=1.675
+ $X2=2.67 $Y2=2.465
r107 17 46 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.655 $Y=1.345
+ $X2=2.655 $Y2=1.51
r108 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.655 $Y=1.345
+ $X2=2.655 $Y2=0.655
r109 13 45 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.24 $Y=1.675
+ $X2=2.24 $Y2=1.51
r110 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.24 $Y=1.675
+ $X2=2.24 $Y2=2.465
r111 9 44 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.345
+ $X2=2.225 $Y2=1.51
r112 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.225 $Y=1.345
+ $X2=2.225 $Y2=0.655
r113 5 40 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.675
+ $X2=1.81 $Y2=1.51
r114 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.81 $Y=1.675
+ $X2=1.81 $Y2=2.465
r115 1 39 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.345
+ $X2=1.795 $Y2=1.51
r116 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.795 $Y=1.345
+ $X2=1.795 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_4%B1 3 7 11 15 19 23 27 30 32 36 37 39 40 41
+ 56 59 61 62 69 71
c125 56 0 1.55509e-19 $X=4.86 $Y=1.44
c126 30 0 1.08593e-19 $X=7.04 $Y=2.465
c127 7 0 2.60081e-19 $X=4.03 $Y=2.465
r128 56 57 4.46296 $w=3.24e-07 $l=3e-08 $layer=POLY_cond $X=4.86 $Y=1.44
+ $X2=4.89 $Y2=1.44
r129 55 61 3.01408 $w=3.23e-07 $l=8.5e-08 $layer=LI1_cond $X=4.8 $Y=1.372
+ $X2=4.885 $Y2=1.372
r130 54 56 8.92593 $w=3.24e-07 $l=6e-08 $layer=POLY_cond $X=4.8 $Y=1.44 $X2=4.86
+ $Y2=1.44
r131 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.8
+ $Y=1.44 $X2=4.8 $Y2=1.44
r132 52 54 50.5802 $w=3.24e-07 $l=3.4e-07 $layer=POLY_cond $X=4.46 $Y=1.44
+ $X2=4.8 $Y2=1.44
r133 51 52 4.46296 $w=3.24e-07 $l=3e-08 $layer=POLY_cond $X=4.43 $Y=1.44
+ $X2=4.46 $Y2=1.44
r134 50 62 1.5099 $w=3.25e-07 $l=3.7e-08 $layer=LI1_cond $X=4.12 $Y=1.372
+ $X2=4.157 $Y2=1.372
r135 50 69 1.64865 $w=2.96e-07 $l=4e-08 $layer=LI1_cond $X=4.12 $Y=1.372
+ $X2=4.08 $Y2=1.372
r136 49 51 46.1173 $w=3.24e-07 $l=3.1e-07 $layer=POLY_cond $X=4.12 $Y=1.44
+ $X2=4.43 $Y2=1.44
r137 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.12
+ $Y=1.44 $X2=4.12 $Y2=1.44
r138 47 49 13.3889 $w=3.24e-07 $l=9e-08 $layer=POLY_cond $X=4.03 $Y=1.44
+ $X2=4.12 $Y2=1.44
r139 46 47 4.46296 $w=3.24e-07 $l=3e-08 $layer=POLY_cond $X=4 $Y=1.44 $X2=4.03
+ $Y2=1.44
r140 41 61 3.69742 $w=2.38e-07 $l=7.7e-08 $layer=LI1_cond $X=5.005 $Y=1.295
+ $X2=5.005 $Y2=1.372
r141 41 71 9.84378 $w=2.38e-07 $l=2.05e-07 $layer=LI1_cond $X=5.005 $Y=1.295
+ $X2=5.005 $Y2=1.09
r142 40 55 8.51035 $w=3.23e-07 $l=2.4e-07 $layer=LI1_cond $X=4.56 $Y=1.372
+ $X2=4.8 $Y2=1.372
r143 39 69 0.164865 $w=2.96e-07 $l=4e-09 $layer=LI1_cond $X=4.076 $Y=1.372
+ $X2=4.08 $Y2=1.372
r144 39 40 14.1485 $w=3.23e-07 $l=3.99e-07 $layer=LI1_cond $X=4.161 $Y=1.372
+ $X2=4.56 $Y2=1.372
r145 39 62 0.141839 $w=3.23e-07 $l=4e-09 $layer=LI1_cond $X=4.161 $Y=1.372
+ $X2=4.157 $Y2=1.372
r146 37 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.1 $Y=1.35
+ $X2=7.1 $Y2=1.515
r147 37 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.1 $Y=1.35
+ $X2=7.1 $Y2=1.185
r148 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.1
+ $Y=1.35 $X2=7.1 $Y2=1.35
r149 34 36 7.61047 $w=2.63e-07 $l=1.75e-07 $layer=LI1_cond $X=7.062 $Y=1.175
+ $X2=7.062 $Y2=1.35
r150 33 71 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.125 $Y=1.09
+ $X2=5.005 $Y2=1.09
r151 32 34 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=6.93 $Y=1.09
+ $X2=7.062 $Y2=1.175
r152 32 33 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=6.93 $Y=1.09
+ $X2=5.125 $Y2=1.09
r153 30 60 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.04 $Y=2.465
+ $X2=7.04 $Y2=1.515
r154 27 59 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.01 $Y=0.655
+ $X2=7.01 $Y2=1.185
r155 21 57 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.605
+ $X2=4.89 $Y2=1.44
r156 21 23 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.89 $Y=1.605
+ $X2=4.89 $Y2=2.465
r157 17 56 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.86 $Y=1.275
+ $X2=4.86 $Y2=1.44
r158 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=4.86 $Y=1.275
+ $X2=4.86 $Y2=0.655
r159 13 52 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.46 $Y=1.605
+ $X2=4.46 $Y2=1.44
r160 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.46 $Y=1.605
+ $X2=4.46 $Y2=2.465
r161 9 51 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.43 $Y=1.275
+ $X2=4.43 $Y2=1.44
r162 9 11 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=4.43 $Y=1.275
+ $X2=4.43 $Y2=0.655
r163 5 47 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.03 $Y=1.605
+ $X2=4.03 $Y2=1.44
r164 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.03 $Y=1.605
+ $X2=4.03 $Y2=2.465
r165 1 46 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4 $Y=1.275 $X2=4
+ $Y2=1.44
r166 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=4 $Y=1.275 $X2=4
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_4%B2 3 7 11 15 19 23 27 31 40 43 52 57
c88 52 0 1.55509e-19 $X=5.81 $Y=1.44
c89 40 0 1.08593e-19 $X=6.49 $Y=1.44
r90 56 57 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.58 $Y=1.44 $X2=6.61
+ $Y2=1.44
r91 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.81
+ $Y=1.44 $X2=5.81 $Y2=1.44
r92 49 51 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.75 $Y=1.44 $X2=5.81
+ $Y2=1.44
r93 48 49 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.72 $Y=1.44 $X2=5.75
+ $Y2=1.44
r94 47 48 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=5.32 $Y=1.44 $X2=5.72
+ $Y2=1.44
r95 45 47 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.29 $Y=1.44 $X2=5.32
+ $Y2=1.44
r96 43 52 8.36451 $w=3.08e-07 $l=2.25e-07 $layer=LI1_cond $X=5.965 $Y=1.665
+ $X2=5.965 $Y2=1.44
r97 41 56 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.49 $Y=1.44 $X2=6.58
+ $Y2=1.44
r98 41 54 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=6.49 $Y=1.44 $X2=6.18
+ $Y2=1.44
r99 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.49
+ $Y=1.44 $X2=6.49 $Y2=1.44
r100 38 54 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.15 $Y=1.44 $X2=6.18
+ $Y2=1.44
r101 38 51 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.15 $Y=1.44
+ $X2=5.81 $Y2=1.44
r102 37 40 19.8469 $w=1.88e-07 $l=3.4e-07 $layer=LI1_cond $X=6.15 $Y=1.44
+ $X2=6.49 $Y2=1.44
r103 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.15
+ $Y=1.44 $X2=6.15 $Y2=1.44
r104 35 52 3.60126 $w=1.9e-07 $l=1.55e-07 $layer=LI1_cond $X=6.12 $Y=1.44
+ $X2=5.965 $Y2=1.44
r105 35 37 1.7512 $w=1.88e-07 $l=3e-08 $layer=LI1_cond $X=6.12 $Y=1.44 $X2=6.15
+ $Y2=1.44
r106 29 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.61 $Y=1.605
+ $X2=6.61 $Y2=1.44
r107 29 31 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.61 $Y=1.605
+ $X2=6.61 $Y2=2.465
r108 25 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.58 $Y=1.275
+ $X2=6.58 $Y2=1.44
r109 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.58 $Y=1.275
+ $X2=6.58 $Y2=0.655
r110 21 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.18 $Y=1.605
+ $X2=6.18 $Y2=1.44
r111 21 23 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.18 $Y=1.605
+ $X2=6.18 $Y2=2.465
r112 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.15 $Y=1.275
+ $X2=6.15 $Y2=1.44
r113 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.15 $Y=1.275
+ $X2=6.15 $Y2=0.655
r114 13 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.75 $Y=1.605
+ $X2=5.75 $Y2=1.44
r115 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.75 $Y=1.605
+ $X2=5.75 $Y2=2.465
r116 9 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.72 $Y=1.275
+ $X2=5.72 $Y2=1.44
r117 9 11 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.72 $Y=1.275
+ $X2=5.72 $Y2=0.655
r118 5 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.32 $Y=1.605
+ $X2=5.32 $Y2=1.44
r119 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.32 $Y=1.605
+ $X2=5.32 $Y2=2.465
r120 1 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.29 $Y=1.275
+ $X2=5.29 $Y2=1.44
r121 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.29 $Y=1.275
+ $X2=5.29 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_4%VPWR 1 2 3 4 5 16 18 24 28 30 34 36 38 42 43
+ 44 46 58 70 73 77
r108 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r109 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r110 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r111 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r112 65 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r113 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r114 62 65 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 62 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 61 64 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r117 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r118 59 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=3.33
+ $X2=4.675 $Y2=3.33
r119 59 61 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.84 $Y=3.33 $X2=5.04
+ $Y2=3.33
r120 58 76 4.4922 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=7.09 $Y=3.33
+ $X2=7.385 $Y2=3.33
r121 58 64 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.09 $Y=3.33
+ $X2=6.96 $Y2=3.33
r122 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r123 54 57 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r124 54 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 53 56 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r126 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 51 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.33 $Y=3.33
+ $X2=1.165 $Y2=3.33
r128 51 53 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.33 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 50 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r131 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r132 47 67 4.32199 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=3.33
+ $X2=0.215 $Y2=3.33
r133 47 49 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 46 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=1.165
+ $Y2=3.33
r135 46 49 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r136 44 74 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r137 44 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r138 42 56 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.65 $Y=3.33 $X2=3.6
+ $Y2=3.33
r139 42 43 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.65 $Y=3.33
+ $X2=3.805 $Y2=3.33
r140 38 41 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=7.255 $Y=2.19
+ $X2=7.255 $Y2=2.95
r141 36 76 3.27398 $w=3.3e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.255 $Y=3.245
+ $X2=7.385 $Y2=3.33
r142 36 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.255 $Y=3.245
+ $X2=7.255 $Y2=2.95
r143 32 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.675 $Y=3.245
+ $X2=4.675 $Y2=3.33
r144 32 34 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=4.675 $Y=3.245
+ $X2=4.675 $Y2=2.515
r145 31 43 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.96 $Y=3.33
+ $X2=3.805 $Y2=3.33
r146 30 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.51 $Y=3.33
+ $X2=4.675 $Y2=3.33
r147 30 31 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.51 $Y=3.33
+ $X2=3.96 $Y2=3.33
r148 26 43 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=3.245
+ $X2=3.805 $Y2=3.33
r149 26 28 16.3573 $w=3.08e-07 $l=4.4e-07 $layer=LI1_cond $X=3.805 $Y=3.245
+ $X2=3.805 $Y2=2.805
r150 22 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=3.245
+ $X2=1.165 $Y2=3.33
r151 22 24 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.165 $Y=3.245
+ $X2=1.165 $Y2=2.795
r152 18 21 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=0.285 $Y=1.98
+ $X2=0.285 $Y2=2.95
r153 16 67 3.11585 $w=2.9e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.215 $Y2=3.33
r154 16 21 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.285 $Y2=2.95
r155 5 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.115
+ $Y=1.835 $X2=7.255 $Y2=2.95
r156 5 38 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=7.115
+ $Y=1.835 $X2=7.255 $Y2=2.19
r157 4 34 300 $w=1.7e-07 $l=7.46726e-07 $layer=licon1_PDIFF $count=2 $X=4.535
+ $Y=1.835 $X2=4.675 $Y2=2.515
r158 3 28 600 $w=1.7e-07 $l=1.05847e-06 $layer=licon1_PDIFF $count=1 $X=3.605
+ $Y=1.835 $X2=3.79 $Y2=2.805
r159 2 24 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.835 $X2=1.165 $Y2=2.795
r160 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.835 $X2=0.305 $Y2=2.95
r161 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.835 $X2=0.305 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_4%A_119_367# 1 2 3 4 15 19 21 22 27 30
c41 27 0 9.96699e-20 $X=3.315 $Y=2.915
r42 25 27 34.7755 $w=2.83e-07 $l=8.6e-07 $layer=LI1_cond $X=2.455 $Y=2.932
+ $X2=3.315 $Y2=2.932
r43 23 34 2.93074 $w=2.85e-07 $l=1e-07 $layer=LI1_cond $X=1.7 $Y=2.932 $X2=1.6
+ $Y2=2.932
r44 23 25 30.5296 $w=2.83e-07 $l=7.55e-07 $layer=LI1_cond $X=1.7 $Y=2.932
+ $X2=2.455 $Y2=2.932
r45 22 34 4.16165 $w=2e-07 $l=1.42e-07 $layer=LI1_cond $X=1.6 $Y=2.79 $X2=1.6
+ $Y2=2.932
r46 21 32 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=2.46 $X2=1.6
+ $Y2=2.375
r47 21 22 18.3 $w=1.98e-07 $l=3.3e-07 $layer=LI1_cond $X=1.6 $Y=2.46 $X2=1.6
+ $Y2=2.79
r48 20 30 2.64776 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.855 $Y=2.375
+ $X2=0.727 $Y2=2.375
r49 19 32 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.5 $Y=2.375 $X2=1.6
+ $Y2=2.375
r50 19 20 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.5 $Y=2.375
+ $X2=0.855 $Y2=2.375
r51 13 30 3.80849 $w=2.42e-07 $l=8.5e-08 $layer=LI1_cond $X=0.727 $Y=2.29
+ $X2=0.727 $Y2=2.375
r52 13 15 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.727 $Y=2.29
+ $X2=0.727 $Y2=1.98
r53 4 27 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=3.175
+ $Y=1.835 $X2=3.315 $Y2=2.915
r54 3 25 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.835 $X2=2.455 $Y2=2.915
r55 2 34 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.455
+ $Y=1.835 $X2=1.595 $Y2=2.91
r56 2 32 600 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=1 $X=1.455
+ $Y=1.835 $X2=1.595 $Y2=2.455
r57 1 30 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.835 $X2=0.735 $Y2=2.44
r58 1 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.835 $X2=0.735 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_4%Y 1 2 3 4 5 6 7 8 29 32 33 34 35 43 45 47 49
+ 51 53 56 58 59 68 69 73 81 83
r148 73 81 1.22538 $w=3.93e-07 $l=4.2e-08 $layer=LI1_cond $X=4.518 $Y=0.842
+ $X2=4.56 $Y2=0.842
r149 69 83 7.02476 $w=3.93e-07 $l=1.34e-07 $layer=LI1_cond $X=4.581 $Y=0.842
+ $X2=4.715 $Y2=0.842
r150 69 81 0.612691 $w=3.93e-07 $l=2.1e-08 $layer=LI1_cond $X=4.581 $Y=0.842
+ $X2=4.56 $Y2=0.842
r151 69 73 0.641867 $w=3.93e-07 $l=2.2e-08 $layer=LI1_cond $X=4.496 $Y=0.842
+ $X2=4.518 $Y2=0.842
r152 69 78 8.19839 $w=3.93e-07 $l=2.81e-07 $layer=LI1_cond $X=4.496 $Y=0.842
+ $X2=4.215 $Y2=0.842
r153 68 78 3.93873 $w=3.93e-07 $l=1.35e-07 $layer=LI1_cond $X=4.08 $Y=0.842
+ $X2=4.215 $Y2=0.842
r154 66 67 1.44746 $w=2.95e-07 $l=3.5e-08 $layer=LI1_cond $X=6.395 $Y=1.98
+ $X2=6.395 $Y2=2.015
r155 64 66 7.85763 $w=2.95e-07 $l=1.9e-07 $layer=LI1_cond $X=6.395 $Y=1.79
+ $X2=6.395 $Y2=1.98
r156 62 63 1.44746 $w=2.95e-07 $l=3.5e-08 $layer=LI1_cond $X=5.535 $Y=1.98
+ $X2=5.535 $Y2=2.015
r157 60 62 7.85763 $w=2.95e-07 $l=1.9e-07 $layer=LI1_cond $X=5.535 $Y=1.79
+ $X2=5.535 $Y2=1.98
r158 58 59 8.12648 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=2.455
+ $X2=3.05 $Y2=2.455
r159 55 56 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=7.45 $Y=0.835
+ $X2=7.45 $Y2=1.705
r160 54 64 3.96227 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.56 $Y=1.79
+ $X2=6.395 $Y2=1.79
r161 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.365 $Y=1.79
+ $X2=7.45 $Y2=1.705
r162 53 54 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=7.365 $Y=1.79
+ $X2=6.56 $Y2=1.79
r163 49 67 3.30767 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.395 $Y=2.1
+ $X2=6.395 $Y2=2.015
r164 49 51 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=6.395 $Y=2.1
+ $X2=6.395 $Y2=2.615
r165 48 63 3.96227 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.7 $Y=2.015
+ $X2=5.535 $Y2=2.015
r166 47 67 3.96227 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=2.015
+ $X2=6.395 $Y2=2.015
r167 47 48 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.23 $Y=2.015
+ $X2=5.7 $Y2=2.015
r168 43 63 3.30767 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=2.1
+ $X2=5.535 $Y2=2.015
r169 43 45 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=5.535 $Y=2.1
+ $X2=5.535 $Y2=2.615
r170 40 42 50.201 $w=1.88e-07 $l=8.6e-07 $layer=LI1_cond $X=5.935 $Y=0.74
+ $X2=6.795 $Y2=0.74
r171 38 40 50.201 $w=1.88e-07 $l=8.6e-07 $layer=LI1_cond $X=5.075 $Y=0.74
+ $X2=5.935 $Y2=0.74
r172 38 83 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=5.075 $Y=0.74
+ $X2=4.715 $Y2=0.74
r173 35 55 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.365 $Y=0.74
+ $X2=7.45 $Y2=0.835
r174 35 42 33.2727 $w=1.88e-07 $l=5.7e-07 $layer=LI1_cond $X=7.365 $Y=0.74
+ $X2=6.795 $Y2=0.74
r175 33 60 3.96227 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.37 $Y=1.79
+ $X2=5.535 $Y2=1.79
r176 33 34 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=5.37 $Y=1.79
+ $X2=3.96 $Y2=1.79
r177 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.875 $Y=1.875
+ $X2=3.96 $Y2=1.79
r178 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.875 $Y=1.875
+ $X2=3.875 $Y2=2.29
r179 29 32 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.79 $Y=2.38
+ $X2=3.875 $Y2=2.29
r180 29 59 45.596 $w=1.78e-07 $l=7.4e-07 $layer=LI1_cond $X=3.79 $Y=2.38
+ $X2=3.05 $Y2=2.38
r181 27 58 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.025 $Y=2.455
+ $X2=2.885 $Y2=2.455
r182 8 66 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=1.835 $X2=6.395 $Y2=1.98
r183 8 51 600 $w=1.7e-07 $l=8.47113e-07 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=1.835 $X2=6.395 $Y2=2.615
r184 7 62 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=1.835 $X2=5.535 $Y2=1.98
r185 7 45 600 $w=1.7e-07 $l=8.47113e-07 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=1.835 $X2=5.535 $Y2=2.615
r186 6 58 600 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.835 $X2=2.885 $Y2=2.455
r187 5 27 600 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=1 $X=1.885
+ $Y=1.835 $X2=2.025 $Y2=2.455
r188 4 42 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.235 $X2=6.795 $Y2=0.74
r189 3 40 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.235 $X2=5.935 $Y2=0.74
r190 2 38 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=4.935
+ $Y=0.235 $X2=5.075 $Y2=0.74
r191 1 78 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=4.075
+ $Y=0.235 $X2=4.215 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_4%A_821_367# 1 2 3 4 13 15 17 19 23 24 27 29
+ 31 33 39
r37 31 41 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.825 $Y=2.905
+ $X2=6.825 $Y2=2.99
r38 31 33 40.5694 $w=1.88e-07 $l=6.95e-07 $layer=LI1_cond $X=6.825 $Y=2.905
+ $X2=6.825 $Y2=2.21
r39 30 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.06 $Y=2.99
+ $X2=5.965 $Y2=2.99
r40 29 41 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.73 $Y=2.99
+ $X2=6.825 $Y2=2.99
r41 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.73 $Y=2.99
+ $X2=6.06 $Y2=2.99
r42 25 39 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.965 $Y=2.905
+ $X2=5.965 $Y2=2.99
r43 25 27 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=5.965 $Y=2.905
+ $X2=5.965 $Y2=2.435
r44 23 39 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.87 $Y=2.99
+ $X2=5.965 $Y2=2.99
r45 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.87 $Y=2.99 $X2=5.2
+ $Y2=2.99
r46 20 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.105 $Y=2.905
+ $X2=5.2 $Y2=2.99
r47 20 22 0.291866 $w=1.88e-07 $l=5e-09 $layer=LI1_cond $X=5.105 $Y=2.905
+ $X2=5.105 $Y2=2.9
r48 19 38 3.31928 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=5.105 $Y=2.225
+ $X2=5.105 $Y2=2.135
r49 19 22 39.4019 $w=1.88e-07 $l=6.75e-07 $layer=LI1_cond $X=5.105 $Y=2.225
+ $X2=5.105 $Y2=2.9
r50 18 36 3.69874 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=4.34 $Y=2.135
+ $X2=4.235 $Y2=2.135
r51 17 38 3.50369 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.01 $Y=2.135
+ $X2=5.105 $Y2=2.135
r52 17 18 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=5.01 $Y=2.135
+ $X2=4.34 $Y2=2.135
r53 13 36 3.17035 $w=2.1e-07 $l=9e-08 $layer=LI1_cond $X=4.235 $Y=2.225
+ $X2=4.235 $Y2=2.135
r54 13 15 36.1775 $w=2.08e-07 $l=6.85e-07 $layer=LI1_cond $X=4.235 $Y=2.225
+ $X2=4.235 $Y2=2.91
r55 4 41 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.685
+ $Y=1.835 $X2=6.825 $Y2=2.91
r56 4 33 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=6.685
+ $Y=1.835 $X2=6.825 $Y2=2.21
r57 3 27 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=5.825
+ $Y=1.835 $X2=5.965 $Y2=2.435
r58 2 38 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.835 $X2=5.105 $Y2=2.21
r59 2 22 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.835 $X2=5.105 $Y2=2.9
r60 1 36 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.835 $X2=4.245 $Y2=2.21
r61 1 15 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.835 $X2=4.245 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_4%A_33_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38 42
+ 44 48 50 52 53 62 64 65 66
c94 50 0 6.80066e-20 $X=3.635 $Y=1.09
r95 60 62 45.05 $w=2.18e-07 $l=8.6e-07 $layer=LI1_cond $X=6.365 $Y=0.365
+ $X2=7.225 $Y2=0.365
r96 58 60 45.05 $w=2.18e-07 $l=8.6e-07 $layer=LI1_cond $X=5.505 $Y=0.365
+ $X2=6.365 $Y2=0.365
r97 56 58 45.05 $w=2.18e-07 $l=8.6e-07 $layer=LI1_cond $X=4.645 $Y=0.365
+ $X2=5.505 $Y2=0.365
r98 54 68 3.10749 $w=2.2e-07 $l=9e-08 $layer=LI1_cond $X=3.815 $Y=0.365
+ $X2=3.725 $Y2=0.365
r99 54 56 43.4785 $w=2.18e-07 $l=8.3e-07 $layer=LI1_cond $X=3.815 $Y=0.365
+ $X2=4.645 $Y2=0.365
r100 52 68 3.79804 $w=1.8e-07 $l=1.1e-07 $layer=LI1_cond $X=3.725 $Y=0.475
+ $X2=3.725 $Y2=0.365
r101 52 53 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=3.725 $Y=0.475
+ $X2=3.725 $Y2=1.005
r102 51 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.965 $Y=1.09
+ $X2=2.87 $Y2=1.09
r103 50 53 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.635 $Y=1.09
+ $X2=3.725 $Y2=1.005
r104 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.635 $Y=1.09
+ $X2=2.965 $Y2=1.09
r105 46 66 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.005
+ $X2=2.87 $Y2=1.09
r106 46 48 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=2.87 $Y=1.005
+ $X2=2.87 $Y2=0.42
r107 45 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.105 $Y=1.09
+ $X2=2.01 $Y2=1.09
r108 44 66 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.775 $Y=1.09
+ $X2=2.87 $Y2=1.09
r109 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.775 $Y=1.09
+ $X2=2.105 $Y2=1.09
r110 40 65 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=1.005
+ $X2=2.01 $Y2=1.09
r111 40 42 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=2.01 $Y=1.005
+ $X2=2.01 $Y2=0.42
r112 39 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.245 $Y=1.09
+ $X2=1.15 $Y2=1.09
r113 38 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.915 $Y=1.09
+ $X2=2.01 $Y2=1.09
r114 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.915 $Y=1.09
+ $X2=1.245 $Y2=1.09
r115 34 64 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=1.005
+ $X2=1.15 $Y2=1.09
r116 34 36 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=1.15 $Y=1.005
+ $X2=1.15 $Y2=0.42
r117 32 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.055 $Y=1.09
+ $X2=1.15 $Y2=1.09
r118 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.055 $Y=1.09
+ $X2=0.385 $Y2=1.09
r119 28 33 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.255 $Y=1.005
+ $X2=0.385 $Y2=1.09
r120 28 30 25.93 $w=2.58e-07 $l=5.85e-07 $layer=LI1_cond $X=0.255 $Y=1.005
+ $X2=0.255 $Y2=0.42
r121 9 62 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=7.085
+ $Y=0.235 $X2=7.225 $Y2=0.37
r122 8 60 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=6.225
+ $Y=0.235 $X2=6.365 $Y2=0.37
r123 7 58 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=5.365
+ $Y=0.235 $X2=5.505 $Y2=0.37
r124 6 56 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=4.505
+ $Y=0.235 $X2=4.645 $Y2=0.37
r125 5 68 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.59
+ $Y=0.235 $X2=3.73 $Y2=0.42
r126 4 48 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.73
+ $Y=0.235 $X2=2.87 $Y2=0.42
r127 3 42 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.235 $X2=2.01 $Y2=0.42
r128 2 36 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.01
+ $Y=0.235 $X2=1.15 $Y2=0.42
r129 1 30 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 40 59 60 63
r96 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 59 60 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r98 56 59 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=7.44
+ $Y2=0
r99 56 57 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r100 54 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r101 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r102 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r103 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r104 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r105 48 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r106 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r107 45 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.72
+ $Y2=0
r108 45 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.2
+ $Y2=0
r109 43 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r110 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r111 40 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.72
+ $Y2=0
r112 40 42 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0
+ $X2=0.24 $Y2=0
r113 38 60 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=7.44
+ $Y2=0
r114 38 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r115 36 53 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.12
+ $Y2=0
r116 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.3
+ $Y2=0
r117 35 56 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.6
+ $Y2=0
r118 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=0 $X2=3.3
+ $Y2=0
r119 33 50 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.275 $Y=0
+ $X2=2.16 $Y2=0
r120 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.44
+ $Y2=0
r121 32 53 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.605 $Y=0
+ $X2=3.12 $Y2=0
r122 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.605 $Y=0 $X2=2.44
+ $Y2=0
r123 30 47 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.2
+ $Y2=0
r124 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.58
+ $Y2=0
r125 29 50 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.745 $Y=0
+ $X2=2.16 $Y2=0
r126 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.58
+ $Y2=0
r127 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=0.085 $X2=3.3
+ $Y2=0
r128 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.3 $Y=0.085
+ $X2=3.3 $Y2=0.38
r129 21 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.44 $Y=0.085
+ $X2=2.44 $Y2=0
r130 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.44 $Y=0.085
+ $X2=2.44 $Y2=0.38
r131 17 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0
r132 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.58 $Y=0.085
+ $X2=1.58 $Y2=0.38
r133 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0
r134 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.72 $Y=0.085
+ $X2=0.72 $Y2=0.38
r135 4 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.16
+ $Y=0.235 $X2=3.3 $Y2=0.38
r136 3 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.3
+ $Y=0.235 $X2=2.44 $Y2=0.38
r137 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.44
+ $Y=0.235 $X2=1.58 $Y2=0.38
r138 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.58
+ $Y=0.235 $X2=0.72 $Y2=0.38
.ends

