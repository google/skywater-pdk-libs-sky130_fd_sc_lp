* File: sky130_fd_sc_lp__o21bai_lp.spice
* Created: Fri Aug 28 11:07:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21bai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o21bai_lp  VNB VPB A1 A2 B1_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1_N	B1_N
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A1_M1003_g N_A_28_110#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.09135 AS=0.1197 PD=0.855 PS=1.41 NRD=24.276 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_28_110#_M1006_d N_A2_M1006_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.09135 PD=0.7 PS=0.855 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A_288_21#_M1004_g N_A_28_110#_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_516_47# N_B1_N_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_288_21#_M1008_d N_B1_N_M1008_g A_516_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_140_413# N_A1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.25 W=1 AD=0.105
+ AS=0.285 PD=1.21 PS=2.57 NRD=9.8303 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1000 N_Y_M1000_d N_A2_M1000_g A_140_413# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=9.8303 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_A_288_21#_M1005_g N_Y_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.27 AS=0.14 PD=1.605 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1001 N_A_288_21#_M1001_d N_B1_N_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.27 PD=2.57 PS=1.605 NRD=0 NRS=51.2003 M=1 R=4 SA=125002
+ SB=125000 A=0.25 P=2.5 MULT=1
DX9_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o21bai_lp.pxi.spice"
*
.ends
*
*
