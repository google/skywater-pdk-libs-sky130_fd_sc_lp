* File: sky130_fd_sc_lp__dfxtp_1.pxi.spice
* Created: Wed Sep  2 09:45:07 2020
* 
x_PM_SKY130_FD_SC_LP__DFXTP_1%CLK N_CLK_c_151_n N_CLK_M1002_g N_CLK_M1021_g
+ N_CLK_c_153_n N_CLK_c_154_n N_CLK_c_159_n CLK CLK CLK CLK N_CLK_c_156_n
+ PM_SKY130_FD_SC_LP__DFXTP_1%CLK
x_PM_SKY130_FD_SC_LP__DFXTP_1%D N_D_M1023_g N_D_c_183_n N_D_M1018_g D D
+ N_D_c_185_n PM_SKY130_FD_SC_LP__DFXTP_1%D
x_PM_SKY130_FD_SC_LP__DFXTP_1%A_217_413# N_A_217_413#_M1011_s
+ N_A_217_413#_M1012_s N_A_217_413#_M1004_g N_A_217_413#_M1016_g
+ N_A_217_413#_M1009_g N_A_217_413#_c_225_n N_A_217_413#_c_226_n
+ N_A_217_413#_M1003_g N_A_217_413#_c_235_n N_A_217_413#_c_228_n
+ N_A_217_413#_c_237_n N_A_217_413#_c_238_n N_A_217_413#_c_239_n
+ N_A_217_413#_c_240_n N_A_217_413#_c_229_n N_A_217_413#_c_230_n
+ N_A_217_413#_c_243_n N_A_217_413#_c_244_n N_A_217_413#_c_260_p
+ N_A_217_413#_c_268_p N_A_217_413#_c_231_n N_A_217_413#_c_232_n
+ N_A_217_413#_c_246_n N_A_217_413#_c_247_n
+ PM_SKY130_FD_SC_LP__DFXTP_1%A_217_413#
x_PM_SKY130_FD_SC_LP__DFXTP_1%A_668_137# N_A_668_137#_M1005_d
+ N_A_668_137#_M1000_d N_A_668_137#_M1008_g N_A_668_137#_M1022_g
+ N_A_668_137#_c_392_n N_A_668_137#_c_387_n N_A_668_137#_c_394_n
+ N_A_668_137#_c_395_n N_A_668_137#_c_388_n N_A_668_137#_c_389_n
+ N_A_668_137#_c_390_n PM_SKY130_FD_SC_LP__DFXTP_1%A_668_137#
x_PM_SKY130_FD_SC_LP__DFXTP_1%A_526_413# N_A_526_413#_M1020_d
+ N_A_526_413#_M1004_d N_A_526_413#_M1000_g N_A_526_413#_c_460_n
+ N_A_526_413#_M1005_g N_A_526_413#_c_461_n N_A_526_413#_c_462_n
+ N_A_526_413#_c_463_n N_A_526_413#_c_464_n N_A_526_413#_c_465_n
+ PM_SKY130_FD_SC_LP__DFXTP_1%A_526_413#
x_PM_SKY130_FD_SC_LP__DFXTP_1%A_110_70# N_A_110_70#_M1002_d N_A_110_70#_M1021_d
+ N_A_110_70#_c_532_n N_A_110_70#_c_533_n N_A_110_70#_M1012_g
+ N_A_110_70#_M1011_g N_A_110_70#_c_550_n N_A_110_70#_c_551_n
+ N_A_110_70#_c_536_n N_A_110_70#_c_537_n N_A_110_70#_M1020_g
+ N_A_110_70#_c_539_n N_A_110_70#_M1019_g N_A_110_70#_c_553_n
+ N_A_110_70#_M1001_g N_A_110_70#_M1017_g N_A_110_70#_c_541_n
+ N_A_110_70#_c_542_n N_A_110_70#_c_555_n N_A_110_70#_c_543_n
+ N_A_110_70#_c_544_n N_A_110_70#_c_545_n N_A_110_70#_c_546_n
+ N_A_110_70#_c_547_n N_A_110_70#_c_548_n PM_SKY130_FD_SC_LP__DFXTP_1%A_110_70#
x_PM_SKY130_FD_SC_LP__DFXTP_1%A_1158_93# N_A_1158_93#_M1010_d
+ N_A_1158_93#_M1014_d N_A_1158_93#_M1013_g N_A_1158_93#_M1006_g
+ N_A_1158_93#_c_673_n N_A_1158_93#_M1007_g N_A_1158_93#_M1015_g
+ N_A_1158_93#_c_675_n N_A_1158_93#_c_676_n N_A_1158_93#_c_683_n
+ N_A_1158_93#_c_684_n N_A_1158_93#_c_677_n N_A_1158_93#_c_724_p
+ PM_SKY130_FD_SC_LP__DFXTP_1%A_1158_93#
x_PM_SKY130_FD_SC_LP__DFXTP_1%A_957_379# N_A_957_379#_M1009_d
+ N_A_957_379#_M1001_d N_A_957_379#_c_744_n N_A_957_379#_M1010_g
+ N_A_957_379#_c_745_n N_A_957_379#_M1014_g N_A_957_379#_c_753_n
+ N_A_957_379#_c_754_n N_A_957_379#_c_747_n N_A_957_379#_c_748_n
+ N_A_957_379#_c_763_n N_A_957_379#_c_749_n N_A_957_379#_c_750_n
+ N_A_957_379#_c_751_n PM_SKY130_FD_SC_LP__DFXTP_1%A_957_379#
x_PM_SKY130_FD_SC_LP__DFXTP_1%VPWR N_VPWR_M1021_s N_VPWR_M1012_d N_VPWR_M1022_d
+ N_VPWR_M1006_d N_VPWR_M1015_s N_VPWR_c_823_n N_VPWR_c_824_n N_VPWR_c_825_n
+ N_VPWR_c_826_n N_VPWR_c_827_n N_VPWR_c_828_n N_VPWR_c_829_n VPWR
+ N_VPWR_c_830_n N_VPWR_c_831_n N_VPWR_c_832_n N_VPWR_c_833_n N_VPWR_c_822_n
+ N_VPWR_c_835_n N_VPWR_c_836_n N_VPWR_c_837_n N_VPWR_c_838_n
+ PM_SKY130_FD_SC_LP__DFXTP_1%VPWR
x_PM_SKY130_FD_SC_LP__DFXTP_1%A_440_413# N_A_440_413#_M1018_d
+ N_A_440_413#_M1023_d N_A_440_413#_c_909_n N_A_440_413#_c_915_n
+ PM_SKY130_FD_SC_LP__DFXTP_1%A_440_413#
x_PM_SKY130_FD_SC_LP__DFXTP_1%Q N_Q_M1007_d N_Q_M1015_d Q Q Q Q Q Q Q
+ N_Q_c_932_n PM_SKY130_FD_SC_LP__DFXTP_1%Q
x_PM_SKY130_FD_SC_LP__DFXTP_1%VGND N_VGND_M1002_s N_VGND_M1011_d N_VGND_M1008_d
+ N_VGND_M1013_d N_VGND_M1007_s N_VGND_c_945_n N_VGND_c_946_n N_VGND_c_947_n
+ N_VGND_c_948_n N_VGND_c_949_n N_VGND_c_950_n N_VGND_c_951_n N_VGND_c_952_n
+ VGND N_VGND_c_953_n N_VGND_c_954_n N_VGND_c_955_n N_VGND_c_956_n
+ N_VGND_c_957_n N_VGND_c_958_n N_VGND_c_959_n N_VGND_c_960_n
+ PM_SKY130_FD_SC_LP__DFXTP_1%VGND
cc_1 VNB N_CLK_c_151_n 0.0238663f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.428
cc_2 VNB N_CLK_M1002_g 0.0298841f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.56
cc_3 VNB N_CLK_c_153_n 0.0233222f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.625
cc_4 VNB N_CLK_c_154_n 0.00191994f $X=-0.19 $Y=-0.245 $X2=0.442 $Y2=1.865
cc_5 VNB CLK 0.0333978f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_CLK_c_156_n 0.0241522f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.12
cc_7 VNB N_D_c_183_n 0.0176548f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.955
cc_8 VNB D 8.19434e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_D_c_185_n 0.0336948f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_A_217_413#_M1016_g 0.0261195f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.625
cc_11 VNB N_A_217_413#_M1009_g 0.0222728f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_12 VNB N_A_217_413#_c_225_n 0.0265877f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_13 VNB N_A_217_413#_c_226_n 0.0493576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_217_413#_M1003_g 0.00635817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_217_413#_c_228_n 0.00673757f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.12
cc_16 VNB N_A_217_413#_c_229_n 0.00370634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_217_413#_c_230_n 0.0194662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_217_413#_c_231_n 0.00927833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_217_413#_c_232_n 8.97215e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_668_137#_M1008_g 0.0182157f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.015
cc_21 VNB N_A_668_137#_c_387_n 0.028107f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_668_137#_c_388_n 0.0035417f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.12
cc_23 VNB N_A_668_137#_c_389_n 0.00782974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_668_137#_c_390_n 0.00423454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_526_413#_c_460_n 0.016459f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_26 VNB N_A_526_413#_c_461_n 0.00640517f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_27 VNB N_A_526_413#_c_462_n 0.00932044f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_A_526_413#_c_463_n 3.7538e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_29 VNB N_A_526_413#_c_464_n 0.00132469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_526_413#_c_465_n 0.0350039f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.12
cc_31 VNB N_A_110_70#_c_532_n 0.0165114f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.56
cc_32 VNB N_A_110_70#_c_533_n 0.0172546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_110_70#_M1012_g 0.00188361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_110_70#_M1011_g 0.0530929f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_35 VNB N_A_110_70#_c_536_n 0.0675572f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_36 VNB N_A_110_70#_c_537_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_110_70#_M1020_g 0.0558156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_110_70#_c_539_n 0.219718f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.12
cc_39 VNB N_A_110_70#_M1017_g 0.036525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_110_70#_c_541_n 0.0098012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_110_70#_c_542_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_110_70#_c_543_n 0.00997866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_110_70#_c_544_n 0.00149064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_110_70#_c_545_n 4.58581e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_110_70#_c_546_n 0.00747554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_110_70#_c_547_n 0.0456571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_110_70#_c_548_n 0.00991919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1158_93#_M1013_g 0.0340924f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.015
cc_49 VNB N_A_1158_93#_c_673_n 0.090302f $X=-0.19 $Y=-0.245 $X2=0.442 $Y2=2.015
cc_50 VNB N_A_1158_93#_M1007_g 0.0259655f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_51 VNB N_A_1158_93#_c_675_n 0.00275628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1158_93#_c_676_n 0.0266436f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.12
cc_53 VNB N_A_1158_93#_c_677_n 0.021192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_957_379#_c_744_n 0.0208806f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.56
cc_55 VNB N_A_957_379#_c_745_n 0.038646f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_56 VNB N_A_957_379#_M1014_g 0.0106522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_957_379#_c_747_n 0.00219706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_957_379#_c_748_n 0.0251145f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.12
cc_59 VNB N_A_957_379#_c_749_n 0.00372729f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.12
cc_60 VNB N_A_957_379#_c_750_n 0.00158418f $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=1.295
cc_61 VNB N_A_957_379#_c_751_n 0.00101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VPWR_c_822_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_440_413#_c_909_n 0.00396641f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=2.015
cc_64 VNB N_Q_c_932_n 0.0627574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_945_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_66 VNB N_VGND_c_946_n 0.0216486f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_67 VNB N_VGND_c_947_n 0.0180213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_948_n 0.033463f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.12
cc_69 VNB N_VGND_c_949_n 0.00994046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_950_n 0.0218065f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_71 VNB N_VGND_c_951_n 0.037664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_952_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_953_n 0.0465304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_954_n 0.0509501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_955_n 0.029584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_956_n 0.0170439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_957_n 0.445046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_958_n 0.00892233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_959_n 0.00620692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_960_n 0.00509721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VPB N_CLK_M1021_g 0.0406496f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_82 VPB N_CLK_c_154_n 0.0138368f $X=-0.19 $Y=1.655 $X2=0.442 $Y2=1.865
cc_83 VPB N_CLK_c_159_n 0.0138993f $X=-0.19 $Y=1.655 $X2=0.442 $Y2=2.015
cc_84 VPB CLK 0.0228521f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_85 VPB N_D_M1023_g 0.0329331f $X=-0.19 $Y=1.655 $X2=0.41 $Y2=1.625
cc_86 VPB D 0.00518963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_D_c_185_n 0.011109f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_88 VPB N_A_217_413#_M1004_g 0.01916f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.015
cc_89 VPB N_A_217_413#_M1003_g 0.0280698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_217_413#_c_235_n 0.00954858f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=0.955
cc_91 VPB N_A_217_413#_c_228_n 0.0031914f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.12
cc_92 VPB N_A_217_413#_c_237_n 0.00521658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_217_413#_c_238_n 8.11598e-19 $X=-0.19 $Y=1.655 $X2=0.255 $Y2=2.035
cc_94 VPB N_A_217_413#_c_239_n 0.0102507f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_217_413#_c_240_n 0.00354423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_217_413#_c_229_n 0.00226955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_217_413#_c_230_n 0.0409852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_217_413#_c_243_n 0.0180602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_217_413#_c_244_n 0.00106916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_217_413#_c_232_n 0.00278921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_217_413#_c_246_n 0.00367817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_217_413#_c_247_n 0.00172351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_668_137#_M1022_g 0.0309257f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.625
cc_104 VPB N_A_668_137#_c_392_n 0.00328532f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_105 VPB N_A_668_137#_c_387_n 0.00808173f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_106 VPB N_A_668_137#_c_394_n 0.00698716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_668_137#_c_395_n 0.00152477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_668_137#_c_389_n 0.00471064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_526_413#_M1000_g 0.0232885f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.015
cc_110 VPB N_A_526_413#_c_461_n 0.00609526f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_111 VPB N_A_526_413#_c_464_n 0.00137469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_526_413#_c_465_n 0.00916022f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.12
cc_113 VPB N_A_110_70#_M1012_g 0.0545267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_110_70#_c_550_n 0.121792f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_115 VPB N_A_110_70#_c_551_n 0.012806f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_116 VPB N_A_110_70#_M1019_g 0.0568313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_110_70#_c_553_n 0.106086f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.12
cc_118 VPB N_A_110_70#_M1001_g 0.0430955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_110_70#_c_555_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_110_70#_c_545_n 0.0166044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_1158_93#_M1006_g 0.0220194f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.625
cc_122 VPB N_A_1158_93#_c_673_n 0.0237626f $X=-0.19 $Y=1.655 $X2=0.442 $Y2=2.015
cc_123 VPB N_A_1158_93#_M1015_g 0.0281399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_1158_93#_c_675_n 0.00394115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_1158_93#_c_676_n 0.0122435f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.12
cc_126 VPB N_A_1158_93#_c_683_n 0.0226189f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=0.955
cc_127 VPB N_A_1158_93#_c_684_n 0.00292334f $X=-0.19 $Y=1.655 $X2=0.255
+ $Y2=1.295
cc_128 VPB N_A_1158_93#_c_677_n 0.0100883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_957_379#_M1014_g 0.0301161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_957_379#_c_753_n 0.00174205f $X=-0.19 $Y=1.655 $X2=0.442
+ $Y2=1.865
cc_131 VPB N_A_957_379#_c_754_n 0.010665f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_132 VPB N_A_957_379#_c_749_n 0.00490387f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.12
cc_133 VPB N_VPWR_c_823_n 0.0112117f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_134 VPB N_VPWR_c_824_n 0.0367112f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_135 VPB N_VPWR_c_825_n 0.0140122f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_826_n 0.0105843f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.12
cc_137 VPB N_VPWR_c_827_n 0.0577143f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_138 VPB N_VPWR_c_828_n 0.0370362f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_139 VPB N_VPWR_c_829_n 0.0333637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_830_n 0.0301921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_831_n 0.05209f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_832_n 0.0280568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_833_n 0.0170439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_822_n 0.120957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_835_n 0.00297041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_836_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_837_n 0.00728331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_838_n 0.00574453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_440_413#_c_909_n 0.00643717f $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=2.015
cc_150 VPB N_Q_c_932_n 0.0577091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 N_CLK_c_151_n N_A_110_70#_c_533_n 0.0209128f $X=0.352 $Y=1.428 $X2=0
+ $Y2=0
cc_152 N_CLK_M1002_g N_A_110_70#_c_543_n 0.00268035f $X=0.475 $Y=0.56 $X2=0
+ $Y2=0
cc_153 CLK N_A_110_70#_c_543_n 0.103091f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_154 N_CLK_c_151_n N_A_110_70#_c_544_n 0.00268035f $X=0.352 $Y=1.428 $X2=0
+ $Y2=0
cc_155 N_CLK_c_154_n N_A_110_70#_c_545_n 0.0049069f $X=0.442 $Y=1.865 $X2=0
+ $Y2=0
cc_156 N_CLK_c_159_n N_A_110_70#_c_545_n 0.0140524f $X=0.442 $Y=2.015 $X2=0
+ $Y2=0
cc_157 N_CLK_c_156_n N_A_110_70#_c_546_n 0.00268035f $X=0.32 $Y=1.12 $X2=0 $Y2=0
cc_158 CLK N_A_110_70#_c_547_n 5.10822e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_159 N_CLK_c_156_n N_A_110_70#_c_547_n 0.0209128f $X=0.32 $Y=1.12 $X2=0 $Y2=0
cc_160 N_CLK_c_153_n N_A_110_70#_c_548_n 0.00268035f $X=0.352 $Y=1.625 $X2=0
+ $Y2=0
cc_161 N_CLK_M1021_g N_VPWR_c_824_n 0.0154699f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_162 N_CLK_c_153_n N_VPWR_c_824_n 5.05536e-19 $X=0.352 $Y=1.625 $X2=0 $Y2=0
cc_163 N_CLK_c_159_n N_VPWR_c_824_n 3.62213e-19 $X=0.442 $Y=2.015 $X2=0 $Y2=0
cc_164 CLK N_VPWR_c_824_n 0.0305153f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_165 N_CLK_M1021_g N_VPWR_c_830_n 0.00396895f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_166 N_CLK_M1021_g N_VPWR_c_822_n 0.00796233f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_167 N_CLK_M1002_g N_VGND_c_946_n 0.0138885f $X=0.475 $Y=0.56 $X2=0 $Y2=0
cc_168 CLK N_VGND_c_946_n 0.0266998f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_169 N_CLK_c_156_n N_VGND_c_946_n 0.00130362f $X=0.32 $Y=1.12 $X2=0 $Y2=0
cc_170 N_CLK_M1002_g N_VGND_c_951_n 0.00396895f $X=0.475 $Y=0.56 $X2=0 $Y2=0
cc_171 N_CLK_M1002_g N_VGND_c_957_n 0.00796233f $X=0.475 $Y=0.56 $X2=0 $Y2=0
cc_172 CLK N_VGND_c_957_n 0.0015796f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_173 N_D_c_185_n N_A_217_413#_M1016_g 0.00196236f $X=2.195 $Y=1.51 $X2=0 $Y2=0
cc_174 N_D_M1023_g N_A_217_413#_c_228_n 8.3456e-19 $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_175 D N_A_217_413#_c_228_n 0.0443895f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_176 N_D_M1023_g N_A_217_413#_c_237_n 0.00523336f $X=2.125 $Y=2.275 $X2=0
+ $Y2=0
cc_177 D N_A_217_413#_c_237_n 0.0424013f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_178 N_D_c_185_n N_A_217_413#_c_237_n 0.00128172f $X=2.195 $Y=1.51 $X2=0 $Y2=0
cc_179 N_D_M1023_g N_A_217_413#_c_238_n 0.011771f $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_180 N_D_M1023_g N_A_217_413#_c_239_n 0.00765926f $X=2.125 $Y=2.275 $X2=0
+ $Y2=0
cc_181 N_D_M1023_g N_A_217_413#_c_240_n 4.783e-19 $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_182 N_D_M1023_g N_A_217_413#_c_229_n 6.67736e-19 $X=2.125 $Y=2.275 $X2=0
+ $Y2=0
cc_183 N_D_M1023_g N_A_217_413#_c_230_n 0.020723f $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_184 N_D_c_185_n N_A_217_413#_c_230_n 0.00649961f $X=2.195 $Y=1.51 $X2=0 $Y2=0
cc_185 N_D_c_183_n N_A_526_413#_c_461_n 6.78917e-19 $X=2.195 $Y=1.345 $X2=0
+ $Y2=0
cc_186 N_D_M1023_g N_A_110_70#_M1012_g 0.0132019f $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_187 D N_A_110_70#_M1012_g 0.00158863f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_188 N_D_c_185_n N_A_110_70#_M1012_g 0.00163056f $X=2.195 $Y=1.51 $X2=0 $Y2=0
cc_189 N_D_c_183_n N_A_110_70#_M1011_g 0.0115108f $X=2.195 $Y=1.345 $X2=0 $Y2=0
cc_190 D N_A_110_70#_M1011_g 0.00804897f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_191 N_D_c_185_n N_A_110_70#_M1011_g 0.0181691f $X=2.195 $Y=1.51 $X2=0 $Y2=0
cc_192 N_D_M1023_g N_A_110_70#_c_550_n 0.00299967f $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_193 N_D_c_183_n N_A_110_70#_c_536_n 0.00484404f $X=2.195 $Y=1.345 $X2=0 $Y2=0
cc_194 N_D_c_183_n N_A_110_70#_M1020_g 0.0125781f $X=2.195 $Y=1.345 $X2=0 $Y2=0
cc_195 D N_A_110_70#_c_541_n 0.00460904f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_196 N_D_M1023_g N_VPWR_c_825_n 8.93275e-19 $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_197 N_D_M1023_g N_A_440_413#_c_909_n 0.00576621f $X=2.125 $Y=2.275 $X2=0
+ $Y2=0
cc_198 N_D_c_183_n N_A_440_413#_c_909_n 0.00272437f $X=2.195 $Y=1.345 $X2=0
+ $Y2=0
cc_199 D N_A_440_413#_c_909_n 0.0427757f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_200 N_D_c_185_n N_A_440_413#_c_909_n 0.00947916f $X=2.195 $Y=1.51 $X2=0 $Y2=0
cc_201 N_D_c_183_n N_A_440_413#_c_915_n 0.00554147f $X=2.195 $Y=1.345 $X2=0
+ $Y2=0
cc_202 D N_VGND_M1011_d 0.0064005f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_203 N_D_c_183_n N_VGND_c_947_n 0.00688977f $X=2.195 $Y=1.345 $X2=0 $Y2=0
cc_204 D N_VGND_c_947_n 0.0292282f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_205 N_D_c_185_n N_VGND_c_947_n 0.00121913f $X=2.195 $Y=1.51 $X2=0 $Y2=0
cc_206 N_D_c_183_n N_VGND_c_957_n 9.72468e-19 $X=2.195 $Y=1.345 $X2=0 $Y2=0
cc_207 N_A_217_413#_c_260_p N_A_668_137#_M1000_d 0.00744487f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_208 N_A_217_413#_M1016_g N_A_668_137#_M1008_g 0.0509957f $X=3.055 $Y=1.025
+ $X2=0 $Y2=0
cc_209 N_A_217_413#_c_230_n N_A_668_137#_M1022_g 0.00258153f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_210 N_A_217_413#_c_243_n N_A_668_137#_M1022_g 3.10585e-19 $X=3.325 $Y=2.742
+ $X2=0 $Y2=0
cc_211 N_A_217_413#_c_244_n N_A_668_137#_M1022_g 0.00284341f $X=3.41 $Y=2.605
+ $X2=0 $Y2=0
cc_212 N_A_217_413#_c_260_p N_A_668_137#_M1022_g 0.0113527f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_213 N_A_217_413#_M1016_g N_A_668_137#_c_392_n 2.9947e-19 $X=3.055 $Y=1.025
+ $X2=0 $Y2=0
cc_214 N_A_217_413#_M1016_g N_A_668_137#_c_387_n 0.00954449f $X=3.055 $Y=1.025
+ $X2=0 $Y2=0
cc_215 N_A_217_413#_c_268_p N_A_668_137#_c_387_n 3.68875e-19 $X=3.495 $Y=2.37
+ $X2=0 $Y2=0
cc_216 N_A_217_413#_c_260_p N_A_668_137#_c_394_n 0.0403677f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_217 N_A_217_413#_c_260_p N_A_668_137#_c_395_n 0.0114121f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_218 N_A_217_413#_c_268_p N_A_668_137#_c_395_n 0.00856116f $X=3.495 $Y=2.37
+ $X2=0 $Y2=0
cc_219 N_A_217_413#_M1009_g N_A_668_137#_c_388_n 0.00186293f $X=4.815 $Y=0.805
+ $X2=0 $Y2=0
cc_220 N_A_217_413#_c_226_n N_A_668_137#_c_389_n 0.00240493f $X=5.175 $Y=1.46
+ $X2=0 $Y2=0
cc_221 N_A_217_413#_c_260_p N_A_668_137#_c_389_n 0.0136682f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_222 N_A_217_413#_c_231_n N_A_668_137#_c_389_n 0.0214511f $X=4.845 $Y=1.595
+ $X2=0 $Y2=0
cc_223 N_A_217_413#_c_232_n N_A_668_137#_c_389_n 0.0285888f $X=4.845 $Y=2.285
+ $X2=0 $Y2=0
cc_224 N_A_217_413#_c_226_n N_A_668_137#_c_390_n 0.00186293f $X=5.175 $Y=1.46
+ $X2=0 $Y2=0
cc_225 N_A_217_413#_c_231_n N_A_668_137#_c_390_n 0.00375266f $X=4.845 $Y=1.595
+ $X2=0 $Y2=0
cc_226 N_A_217_413#_c_229_n N_A_526_413#_M1004_d 0.00410748f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_227 N_A_217_413#_c_243_n N_A_526_413#_M1000_g 9.97658e-19 $X=3.325 $Y=2.742
+ $X2=0 $Y2=0
cc_228 N_A_217_413#_c_260_p N_A_526_413#_M1000_g 0.0124199f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_229 N_A_217_413#_c_232_n N_A_526_413#_M1000_g 6.74093e-19 $X=4.845 $Y=2.285
+ $X2=0 $Y2=0
cc_230 N_A_217_413#_M1009_g N_A_526_413#_c_460_n 0.00883626f $X=4.815 $Y=0.805
+ $X2=0 $Y2=0
cc_231 N_A_217_413#_M1004_g N_A_526_413#_c_461_n 0.00154777f $X=2.555 $Y=2.275
+ $X2=0 $Y2=0
cc_232 N_A_217_413#_M1016_g N_A_526_413#_c_461_n 0.00746291f $X=3.055 $Y=1.025
+ $X2=0 $Y2=0
cc_233 N_A_217_413#_c_229_n N_A_526_413#_c_461_n 0.0632465f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_234 N_A_217_413#_c_230_n N_A_526_413#_c_461_n 0.0126492f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_235 N_A_217_413#_c_243_n N_A_526_413#_c_461_n 0.0164036f $X=3.325 $Y=2.742
+ $X2=0 $Y2=0
cc_236 N_A_217_413#_M1016_g N_A_526_413#_c_463_n 0.0123879f $X=3.055 $Y=1.025
+ $X2=0 $Y2=0
cc_237 N_A_217_413#_c_229_n N_A_526_413#_c_463_n 7.89851e-19 $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_238 N_A_217_413#_c_230_n N_A_526_413#_c_463_n 0.00503429f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_239 N_A_217_413#_c_226_n N_A_526_413#_c_465_n 0.00895651f $X=5.175 $Y=1.46
+ $X2=0 $Y2=0
cc_240 N_A_217_413#_c_228_n N_A_110_70#_c_532_n 0.012356f $X=1.325 $Y=1.02 $X2=0
+ $Y2=0
cc_241 N_A_217_413#_c_246_n N_A_110_70#_c_533_n 0.00494261f $X=1.045 $Y=2.045
+ $X2=0 $Y2=0
cc_242 N_A_217_413#_c_235_n N_A_110_70#_M1012_g 2.3258e-19 $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_243 N_A_217_413#_c_228_n N_A_110_70#_M1012_g 0.0120997f $X=1.325 $Y=1.02
+ $X2=0 $Y2=0
cc_244 N_A_217_413#_c_237_n N_A_110_70#_M1012_g 0.0123887f $X=1.905 $Y=2.045
+ $X2=0 $Y2=0
cc_245 N_A_217_413#_c_238_n N_A_110_70#_M1012_g 0.00167042f $X=1.99 $Y=2.605
+ $X2=0 $Y2=0
cc_246 N_A_217_413#_c_246_n N_A_110_70#_M1012_g 0.00586086f $X=1.045 $Y=2.045
+ $X2=0 $Y2=0
cc_247 N_A_217_413#_c_228_n N_A_110_70#_M1011_g 0.00211455f $X=1.325 $Y=1.02
+ $X2=0 $Y2=0
cc_248 N_A_217_413#_M1004_g N_A_110_70#_c_550_n 0.00299962f $X=2.555 $Y=2.275
+ $X2=0 $Y2=0
cc_249 N_A_217_413#_c_239_n N_A_110_70#_c_550_n 0.00817803f $X=2.595 $Y=2.742
+ $X2=0 $Y2=0
cc_250 N_A_217_413#_c_240_n N_A_110_70#_c_550_n 0.00349153f $X=2.075 $Y=2.742
+ $X2=0 $Y2=0
cc_251 N_A_217_413#_c_243_n N_A_110_70#_c_550_n 0.00663475f $X=3.325 $Y=2.742
+ $X2=0 $Y2=0
cc_252 N_A_217_413#_c_247_n N_A_110_70#_c_550_n 0.00359829f $X=2.685 $Y=2.742
+ $X2=0 $Y2=0
cc_253 N_A_217_413#_M1016_g N_A_110_70#_M1020_g 0.0133385f $X=3.055 $Y=1.025
+ $X2=0 $Y2=0
cc_254 N_A_217_413#_c_229_n N_A_110_70#_M1020_g 7.93057e-19 $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_255 N_A_217_413#_c_230_n N_A_110_70#_M1020_g 0.0106665f $X=2.69 $Y=1.74 $X2=0
+ $Y2=0
cc_256 N_A_217_413#_M1016_g N_A_110_70#_c_539_n 0.0042755f $X=3.055 $Y=1.025
+ $X2=0 $Y2=0
cc_257 N_A_217_413#_M1009_g N_A_110_70#_c_539_n 0.0104164f $X=4.815 $Y=0.805
+ $X2=0 $Y2=0
cc_258 N_A_217_413#_M1004_g N_A_110_70#_M1019_g 0.0074843f $X=2.555 $Y=2.275
+ $X2=0 $Y2=0
cc_259 N_A_217_413#_c_229_n N_A_110_70#_M1019_g 0.00194944f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_260 N_A_217_413#_c_243_n N_A_110_70#_M1019_g 0.0240991f $X=3.325 $Y=2.742
+ $X2=0 $Y2=0
cc_261 N_A_217_413#_c_244_n N_A_110_70#_M1019_g 0.00349413f $X=3.41 $Y=2.605
+ $X2=0 $Y2=0
cc_262 N_A_217_413#_c_268_p N_A_110_70#_M1019_g 0.00349056f $X=3.495 $Y=2.37
+ $X2=0 $Y2=0
cc_263 N_A_217_413#_c_243_n N_A_110_70#_c_553_n 0.00164948f $X=3.325 $Y=2.742
+ $X2=0 $Y2=0
cc_264 N_A_217_413#_c_260_p N_A_110_70#_c_553_n 0.00811928f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_265 N_A_217_413#_c_226_n N_A_110_70#_M1001_g 0.00287639f $X=5.175 $Y=1.46
+ $X2=0 $Y2=0
cc_266 N_A_217_413#_M1003_g N_A_110_70#_M1001_g 0.00712119f $X=5.505 $Y=2.105
+ $X2=0 $Y2=0
cc_267 N_A_217_413#_c_260_p N_A_110_70#_M1001_g 0.0189825f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_268 N_A_217_413#_c_232_n N_A_110_70#_M1001_g 0.0139123f $X=4.845 $Y=2.285
+ $X2=0 $Y2=0
cc_269 N_A_217_413#_M1009_g N_A_110_70#_M1017_g 0.0115228f $X=4.815 $Y=0.805
+ $X2=0 $Y2=0
cc_270 N_A_217_413#_c_225_n N_A_110_70#_M1017_g 0.00831117f $X=5.43 $Y=1.46
+ $X2=0 $Y2=0
cc_271 N_A_217_413#_c_228_n N_A_110_70#_c_541_n 0.00336852f $X=1.325 $Y=1.02
+ $X2=0 $Y2=0
cc_272 N_A_217_413#_c_237_n N_A_110_70#_c_541_n 0.00297883f $X=1.905 $Y=2.045
+ $X2=0 $Y2=0
cc_273 N_A_217_413#_c_228_n N_A_110_70#_c_543_n 0.00505542f $X=1.325 $Y=1.02
+ $X2=0 $Y2=0
cc_274 N_A_217_413#_c_235_n N_A_110_70#_c_545_n 0.0349691f $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_275 N_A_217_413#_c_228_n N_A_110_70#_c_545_n 0.0148107f $X=1.325 $Y=1.02
+ $X2=0 $Y2=0
cc_276 N_A_217_413#_c_246_n N_A_110_70#_c_545_n 0.00965767f $X=1.045 $Y=2.045
+ $X2=0 $Y2=0
cc_277 N_A_217_413#_c_228_n N_A_110_70#_c_546_n 0.0517311f $X=1.325 $Y=1.02
+ $X2=0 $Y2=0
cc_278 N_A_217_413#_c_228_n N_A_110_70#_c_547_n 0.00457503f $X=1.325 $Y=1.02
+ $X2=0 $Y2=0
cc_279 N_A_217_413#_c_225_n N_A_1158_93#_M1013_g 0.0321291f $X=5.43 $Y=1.46
+ $X2=0 $Y2=0
cc_280 N_A_217_413#_c_226_n N_A_1158_93#_M1013_g 0.00235011f $X=5.175 $Y=1.46
+ $X2=0 $Y2=0
cc_281 N_A_217_413#_c_225_n N_A_1158_93#_c_684_n 0.00123406f $X=5.43 $Y=1.46
+ $X2=0 $Y2=0
cc_282 N_A_217_413#_M1003_g N_A_1158_93#_c_677_n 0.0321291f $X=5.505 $Y=2.105
+ $X2=0 $Y2=0
cc_283 N_A_217_413#_c_260_p N_A_957_379#_M1001_d 0.00565152f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_284 N_A_217_413#_c_232_n N_A_957_379#_M1001_d 0.00376738f $X=4.845 $Y=2.285
+ $X2=0 $Y2=0
cc_285 N_A_217_413#_c_226_n N_A_957_379#_c_753_n 0.00339564f $X=5.175 $Y=1.46
+ $X2=0 $Y2=0
cc_286 N_A_217_413#_c_232_n N_A_957_379#_c_753_n 0.0295062f $X=4.845 $Y=2.285
+ $X2=0 $Y2=0
cc_287 N_A_217_413#_c_260_p N_A_957_379#_c_754_n 0.0136604f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_288 N_A_217_413#_M1009_g N_A_957_379#_c_747_n 0.00140583f $X=4.815 $Y=0.805
+ $X2=0 $Y2=0
cc_289 N_A_217_413#_c_225_n N_A_957_379#_c_748_n 0.00483947f $X=5.43 $Y=1.46
+ $X2=0 $Y2=0
cc_290 N_A_217_413#_M1009_g N_A_957_379#_c_763_n 0.00390483f $X=4.815 $Y=0.805
+ $X2=0 $Y2=0
cc_291 N_A_217_413#_c_225_n N_A_957_379#_c_763_n 0.00133249f $X=5.43 $Y=1.46
+ $X2=0 $Y2=0
cc_292 N_A_217_413#_c_226_n N_A_957_379#_c_763_n 0.00567047f $X=5.175 $Y=1.46
+ $X2=0 $Y2=0
cc_293 N_A_217_413#_c_231_n N_A_957_379#_c_763_n 0.00286778f $X=4.845 $Y=1.595
+ $X2=0 $Y2=0
cc_294 N_A_217_413#_c_225_n N_A_957_379#_c_749_n 0.0143831f $X=5.43 $Y=1.46
+ $X2=0 $Y2=0
cc_295 N_A_217_413#_c_226_n N_A_957_379#_c_749_n 0.00122868f $X=5.175 $Y=1.46
+ $X2=0 $Y2=0
cc_296 N_A_217_413#_M1003_g N_A_957_379#_c_749_n 0.0147705f $X=5.505 $Y=2.105
+ $X2=0 $Y2=0
cc_297 N_A_217_413#_c_231_n N_A_957_379#_c_749_n 0.0216921f $X=4.845 $Y=1.595
+ $X2=0 $Y2=0
cc_298 N_A_217_413#_c_232_n N_A_957_379#_c_749_n 0.0150398f $X=4.845 $Y=2.285
+ $X2=0 $Y2=0
cc_299 N_A_217_413#_M1009_g N_A_957_379#_c_750_n 0.00123789f $X=4.815 $Y=0.805
+ $X2=0 $Y2=0
cc_300 N_A_217_413#_c_225_n N_A_957_379#_c_750_n 8.13702e-19 $X=5.43 $Y=1.46
+ $X2=0 $Y2=0
cc_301 N_A_217_413#_c_226_n N_A_957_379#_c_750_n 0.00148399f $X=5.175 $Y=1.46
+ $X2=0 $Y2=0
cc_302 N_A_217_413#_c_231_n N_A_957_379#_c_750_n 0.00813903f $X=4.845 $Y=1.595
+ $X2=0 $Y2=0
cc_303 N_A_217_413#_c_237_n N_VPWR_M1012_d 0.00904105f $X=1.905 $Y=2.045 $X2=0
+ $Y2=0
cc_304 N_A_217_413#_c_238_n N_VPWR_M1012_d 0.00413223f $X=1.99 $Y=2.605 $X2=0
+ $Y2=0
cc_305 N_A_217_413#_c_260_p N_VPWR_M1022_d 0.00734754f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_306 N_A_217_413#_c_235_n N_VPWR_c_825_n 7.2147e-19 $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_307 N_A_217_413#_c_237_n N_VPWR_c_825_n 0.0144005f $X=1.905 $Y=2.045 $X2=0
+ $Y2=0
cc_308 N_A_217_413#_c_238_n N_VPWR_c_825_n 0.0227504f $X=1.99 $Y=2.605 $X2=0
+ $Y2=0
cc_309 N_A_217_413#_c_240_n N_VPWR_c_825_n 0.0235372f $X=2.075 $Y=2.742 $X2=0
+ $Y2=0
cc_310 N_A_217_413#_c_243_n N_VPWR_c_826_n 0.0158898f $X=3.325 $Y=2.742 $X2=0
+ $Y2=0
cc_311 N_A_217_413#_c_260_p N_VPWR_c_826_n 0.0240018f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_312 N_A_217_413#_c_235_n N_VPWR_c_830_n 0.00618524f $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_313 N_A_217_413#_c_239_n N_VPWR_c_831_n 0.0153947f $X=2.595 $Y=2.742 $X2=0
+ $Y2=0
cc_314 N_A_217_413#_c_240_n N_VPWR_c_831_n 0.00538918f $X=2.075 $Y=2.742 $X2=0
+ $Y2=0
cc_315 N_A_217_413#_c_243_n N_VPWR_c_831_n 0.0212904f $X=3.325 $Y=2.742 $X2=0
+ $Y2=0
cc_316 N_A_217_413#_c_247_n N_VPWR_c_831_n 0.00570619f $X=2.685 $Y=2.742 $X2=0
+ $Y2=0
cc_317 N_A_217_413#_M1003_g N_VPWR_c_822_n 0.00373935f $X=5.505 $Y=2.105 $X2=0
+ $Y2=0
cc_318 N_A_217_413#_c_235_n N_VPWR_c_822_n 0.00902036f $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_319 N_A_217_413#_c_239_n N_VPWR_c_822_n 0.0152988f $X=2.595 $Y=2.742 $X2=0
+ $Y2=0
cc_320 N_A_217_413#_c_240_n N_VPWR_c_822_n 0.00520658f $X=2.075 $Y=2.742 $X2=0
+ $Y2=0
cc_321 N_A_217_413#_c_243_n N_VPWR_c_822_n 0.0211706f $X=3.325 $Y=2.742 $X2=0
+ $Y2=0
cc_322 N_A_217_413#_c_247_n N_VPWR_c_822_n 0.00551285f $X=2.685 $Y=2.742 $X2=0
+ $Y2=0
cc_323 N_A_217_413#_M1016_g N_A_440_413#_c_909_n 8.31225e-19 $X=3.055 $Y=1.025
+ $X2=0 $Y2=0
cc_324 N_A_217_413#_c_237_n N_A_440_413#_c_909_n 0.0111246f $X=1.905 $Y=2.045
+ $X2=0 $Y2=0
cc_325 N_A_217_413#_c_239_n N_A_440_413#_c_909_n 0.0146898f $X=2.595 $Y=2.742
+ $X2=0 $Y2=0
cc_326 N_A_217_413#_c_229_n N_A_440_413#_c_909_n 0.0479278f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_327 N_A_217_413#_c_230_n N_A_440_413#_c_909_n 0.00377014f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_328 N_A_217_413#_c_230_n N_A_440_413#_c_915_n 0.00168196f $X=2.69 $Y=1.74
+ $X2=0 $Y2=0
cc_329 N_A_217_413#_c_268_p A_666_413# 9.64975e-19 $X=3.495 $Y=2.37 $X2=-0.19
+ $Y2=-0.245
cc_330 N_A_217_413#_M1016_g N_VGND_c_957_n 9.72468e-19 $X=3.055 $Y=1.025 $X2=0
+ $Y2=0
cc_331 N_A_217_413#_M1009_g N_VGND_c_957_n 9.39239e-19 $X=4.815 $Y=0.805 $X2=0
+ $Y2=0
cc_332 N_A_217_413#_c_228_n N_VGND_c_957_n 0.00885308f $X=1.325 $Y=1.02 $X2=0
+ $Y2=0
cc_333 N_A_668_137#_M1022_g N_A_526_413#_M1000_g 0.0246912f $X=3.615 $Y=2.275
+ $X2=0 $Y2=0
cc_334 N_A_668_137#_c_392_n N_A_526_413#_M1000_g 0.00305791f $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_335 N_A_668_137#_c_387_n N_A_526_413#_M1000_g 6.0939e-19 $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_336 N_A_668_137#_c_394_n N_A_526_413#_M1000_g 0.0136122f $X=4.41 $Y=1.985
+ $X2=0 $Y2=0
cc_337 N_A_668_137#_c_389_n N_A_526_413#_M1000_g 0.00518709f $X=4.495 $Y=1.855
+ $X2=0 $Y2=0
cc_338 N_A_668_137#_c_388_n N_A_526_413#_c_460_n 0.00351765f $X=4.57 $Y=0.74
+ $X2=0 $Y2=0
cc_339 N_A_668_137#_M1008_g N_A_526_413#_c_461_n 0.00390112f $X=3.415 $Y=1.025
+ $X2=0 $Y2=0
cc_340 N_A_668_137#_M1022_g N_A_526_413#_c_461_n 8.19233e-19 $X=3.615 $Y=2.275
+ $X2=0 $Y2=0
cc_341 N_A_668_137#_c_392_n N_A_526_413#_c_461_n 0.0269081f $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_342 N_A_668_137#_c_387_n N_A_526_413#_c_461_n 0.00104456f $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_343 N_A_668_137#_c_395_n N_A_526_413#_c_461_n 0.0151687f $X=3.7 $Y=1.985
+ $X2=0 $Y2=0
cc_344 N_A_668_137#_M1008_g N_A_526_413#_c_462_n 0.0169027f $X=3.415 $Y=1.025
+ $X2=0 $Y2=0
cc_345 N_A_668_137#_c_392_n N_A_526_413#_c_462_n 0.0257346f $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_346 N_A_668_137#_c_387_n N_A_526_413#_c_462_n 0.00583405f $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_347 N_A_668_137#_c_394_n N_A_526_413#_c_462_n 0.00925836f $X=4.41 $Y=1.985
+ $X2=0 $Y2=0
cc_348 N_A_668_137#_c_390_n N_A_526_413#_c_462_n 0.00327951f $X=4.547 $Y=1.245
+ $X2=0 $Y2=0
cc_349 N_A_668_137#_M1008_g N_A_526_413#_c_463_n 0.0013871f $X=3.415 $Y=1.025
+ $X2=0 $Y2=0
cc_350 N_A_668_137#_M1008_g N_A_526_413#_c_464_n 0.00189344f $X=3.415 $Y=1.025
+ $X2=0 $Y2=0
cc_351 N_A_668_137#_c_392_n N_A_526_413#_c_464_n 0.0113761f $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_352 N_A_668_137#_c_387_n N_A_526_413#_c_464_n 0.00145067f $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_353 N_A_668_137#_c_394_n N_A_526_413#_c_464_n 0.0196341f $X=4.41 $Y=1.985
+ $X2=0 $Y2=0
cc_354 N_A_668_137#_c_389_n N_A_526_413#_c_464_n 0.0297561f $X=4.495 $Y=1.855
+ $X2=0 $Y2=0
cc_355 N_A_668_137#_M1008_g N_A_526_413#_c_465_n 5.40088e-19 $X=3.415 $Y=1.025
+ $X2=0 $Y2=0
cc_356 N_A_668_137#_c_392_n N_A_526_413#_c_465_n 9.36413e-19 $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_357 N_A_668_137#_c_387_n N_A_526_413#_c_465_n 0.0141651f $X=3.535 $Y=1.53
+ $X2=0 $Y2=0
cc_358 N_A_668_137#_c_394_n N_A_526_413#_c_465_n 0.00638897f $X=4.41 $Y=1.985
+ $X2=0 $Y2=0
cc_359 N_A_668_137#_c_390_n N_A_526_413#_c_465_n 0.00351765f $X=4.547 $Y=1.245
+ $X2=0 $Y2=0
cc_360 N_A_668_137#_M1008_g N_A_110_70#_c_539_n 0.00495681f $X=3.415 $Y=1.025
+ $X2=0 $Y2=0
cc_361 N_A_668_137#_c_388_n N_A_110_70#_c_539_n 0.00553555f $X=4.57 $Y=0.74
+ $X2=0 $Y2=0
cc_362 N_A_668_137#_M1022_g N_A_110_70#_M1019_g 0.0412139f $X=3.615 $Y=2.275
+ $X2=0 $Y2=0
cc_363 N_A_668_137#_c_395_n N_A_110_70#_M1019_g 0.00124224f $X=3.7 $Y=1.985
+ $X2=0 $Y2=0
cc_364 N_A_668_137#_M1022_g N_A_110_70#_c_553_n 0.00391504f $X=3.615 $Y=2.275
+ $X2=0 $Y2=0
cc_365 N_A_668_137#_c_389_n N_A_110_70#_M1001_g 0.00225297f $X=4.495 $Y=1.855
+ $X2=0 $Y2=0
cc_366 N_A_668_137#_c_390_n N_A_110_70#_M1001_g 0.00163028f $X=4.547 $Y=1.245
+ $X2=0 $Y2=0
cc_367 N_A_668_137#_c_388_n N_A_957_379#_c_747_n 0.00463468f $X=4.57 $Y=0.74
+ $X2=0 $Y2=0
cc_368 N_A_668_137#_c_390_n N_A_957_379#_c_750_n 0.00278978f $X=4.547 $Y=1.245
+ $X2=0 $Y2=0
cc_369 N_A_668_137#_c_394_n N_VPWR_M1022_d 0.00437482f $X=4.41 $Y=1.985 $X2=0
+ $Y2=0
cc_370 N_A_668_137#_M1022_g N_VPWR_c_822_n 9.7053e-19 $X=3.615 $Y=2.275 $X2=0
+ $Y2=0
cc_371 N_A_668_137#_c_395_n A_666_413# 0.00106188f $X=3.7 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_372 N_A_668_137#_M1008_g N_VGND_c_948_n 0.00987181f $X=3.415 $Y=1.025 $X2=0
+ $Y2=0
cc_373 N_A_668_137#_c_388_n N_VGND_c_948_n 0.00164866f $X=4.57 $Y=0.74 $X2=0
+ $Y2=0
cc_374 N_A_668_137#_c_388_n N_VGND_c_954_n 0.00628238f $X=4.57 $Y=0.74 $X2=0
+ $Y2=0
cc_375 N_A_668_137#_M1008_g N_VGND_c_957_n 9.72468e-19 $X=3.415 $Y=1.025 $X2=0
+ $Y2=0
cc_376 N_A_668_137#_c_388_n N_VGND_c_957_n 0.00757207f $X=4.57 $Y=0.74 $X2=0
+ $Y2=0
cc_377 N_A_526_413#_c_461_n N_A_110_70#_M1020_g 7.35428e-19 $X=3.03 $Y=2.27
+ $X2=0 $Y2=0
cc_378 N_A_526_413#_c_463_n N_A_110_70#_M1020_g 4.35816e-19 $X=3.155 $Y=1.19
+ $X2=0 $Y2=0
cc_379 N_A_526_413#_c_460_n N_A_110_70#_c_539_n 0.0104164f $X=4.325 $Y=1.345
+ $X2=0 $Y2=0
cc_380 N_A_526_413#_c_463_n N_A_110_70#_c_539_n 0.00436181f $X=3.155 $Y=1.19
+ $X2=0 $Y2=0
cc_381 N_A_526_413#_c_461_n N_A_110_70#_M1019_g 0.00159149f $X=3.03 $Y=2.27
+ $X2=0 $Y2=0
cc_382 N_A_526_413#_c_462_n N_A_110_70#_M1019_g 0.00375567f $X=3.98 $Y=1.19
+ $X2=0 $Y2=0
cc_383 N_A_526_413#_M1000_g N_A_110_70#_c_553_n 0.0100858f $X=4.2 $Y=2.315 $X2=0
+ $Y2=0
cc_384 N_A_526_413#_M1000_g N_A_110_70#_M1001_g 0.0314706f $X=4.2 $Y=2.315 $X2=0
+ $Y2=0
cc_385 N_A_526_413#_M1000_g N_VPWR_c_826_n 0.00752351f $X=4.2 $Y=2.315 $X2=0
+ $Y2=0
cc_386 N_A_526_413#_M1000_g N_VPWR_c_822_n 9.39239e-19 $X=4.2 $Y=2.315 $X2=0
+ $Y2=0
cc_387 N_A_526_413#_c_461_n N_A_440_413#_c_909_n 0.0105857f $X=3.03 $Y=2.27
+ $X2=0 $Y2=0
cc_388 N_A_526_413#_c_463_n N_A_440_413#_c_909_n 0.00222725f $X=3.155 $Y=1.19
+ $X2=0 $Y2=0
cc_389 N_A_526_413#_c_462_n N_VGND_M1008_d 0.00981033f $X=3.98 $Y=1.19 $X2=0
+ $Y2=0
cc_390 N_A_526_413#_c_460_n N_VGND_c_948_n 0.00651467f $X=4.325 $Y=1.345 $X2=0
+ $Y2=0
cc_391 N_A_526_413#_c_462_n N_VGND_c_948_n 0.0521967f $X=3.98 $Y=1.19 $X2=0
+ $Y2=0
cc_392 N_A_526_413#_c_463_n N_VGND_c_948_n 0.00295801f $X=3.155 $Y=1.19 $X2=0
+ $Y2=0
cc_393 N_A_526_413#_c_465_n N_VGND_c_948_n 0.00109787f $X=4.325 $Y=1.51 $X2=0
+ $Y2=0
cc_394 N_A_526_413#_c_460_n N_VGND_c_957_n 9.39239e-19 $X=4.325 $Y=1.345 $X2=0
+ $Y2=0
cc_395 N_A_526_413#_c_463_n N_VGND_c_957_n 0.0118065f $X=3.155 $Y=1.19 $X2=0
+ $Y2=0
cc_396 N_A_526_413#_c_462_n A_626_163# 0.00366293f $X=3.98 $Y=1.19 $X2=-0.19
+ $Y2=-0.245
cc_397 N_A_110_70#_M1017_g N_A_1158_93#_M1013_g 0.0409028f $X=5.505 $Y=0.805
+ $X2=0 $Y2=0
cc_398 N_A_110_70#_c_539_n N_A_957_379#_c_744_n 0.00167672f $X=5.43 $Y=0.18
+ $X2=0 $Y2=0
cc_399 N_A_110_70#_M1001_g N_A_957_379#_c_753_n 0.00180094f $X=4.71 $Y=2.315
+ $X2=0 $Y2=0
cc_400 N_A_110_70#_M1001_g N_A_957_379#_c_754_n 0.00918138f $X=4.71 $Y=2.315
+ $X2=0 $Y2=0
cc_401 N_A_110_70#_M1017_g N_A_957_379#_c_747_n 0.003401f $X=5.505 $Y=0.805
+ $X2=0 $Y2=0
cc_402 N_A_110_70#_M1017_g N_A_957_379#_c_748_n 0.00829768f $X=5.505 $Y=0.805
+ $X2=0 $Y2=0
cc_403 N_A_110_70#_c_539_n N_A_957_379#_c_763_n 0.0064181f $X=5.43 $Y=0.18 $X2=0
+ $Y2=0
cc_404 N_A_110_70#_M1001_g N_A_957_379#_c_749_n 3.32162e-19 $X=4.71 $Y=2.315
+ $X2=0 $Y2=0
cc_405 N_A_110_70#_c_545_n N_VPWR_c_824_n 0.0258394f $X=0.69 $Y=2.485 $X2=0
+ $Y2=0
cc_406 N_A_110_70#_M1012_g N_VPWR_c_825_n 0.0162969f $X=1.425 $Y=2.385 $X2=0
+ $Y2=0
cc_407 N_A_110_70#_c_550_n N_VPWR_c_825_n 0.0176692f $X=3.18 $Y=3.15 $X2=0 $Y2=0
cc_408 N_A_110_70#_M1019_g N_VPWR_c_826_n 0.00670905f $X=3.255 $Y=2.275 $X2=0
+ $Y2=0
cc_409 N_A_110_70#_c_553_n N_VPWR_c_826_n 0.0254542f $X=4.635 $Y=3.15 $X2=0
+ $Y2=0
cc_410 N_A_110_70#_M1001_g N_VPWR_c_826_n 0.005747f $X=4.71 $Y=2.315 $X2=0 $Y2=0
cc_411 N_A_110_70#_c_553_n N_VPWR_c_827_n 0.0253881f $X=4.635 $Y=3.15 $X2=0
+ $Y2=0
cc_412 N_A_110_70#_c_551_n N_VPWR_c_830_n 0.00620508f $X=1.5 $Y=3.15 $X2=0 $Y2=0
cc_413 N_A_110_70#_c_545_n N_VPWR_c_830_n 0.00920383f $X=0.69 $Y=2.485 $X2=0
+ $Y2=0
cc_414 N_A_110_70#_c_550_n N_VPWR_c_831_n 0.0524766f $X=3.18 $Y=3.15 $X2=0 $Y2=0
cc_415 N_A_110_70#_c_550_n N_VPWR_c_822_n 0.0408977f $X=3.18 $Y=3.15 $X2=0 $Y2=0
cc_416 N_A_110_70#_c_551_n N_VPWR_c_822_n 0.0113608f $X=1.5 $Y=3.15 $X2=0 $Y2=0
cc_417 N_A_110_70#_c_553_n N_VPWR_c_822_n 0.0537184f $X=4.635 $Y=3.15 $X2=0
+ $Y2=0
cc_418 N_A_110_70#_c_555_n N_VPWR_c_822_n 0.00391025f $X=3.255 $Y=3.15 $X2=0
+ $Y2=0
cc_419 N_A_110_70#_c_545_n N_VPWR_c_822_n 0.00735646f $X=0.69 $Y=2.485 $X2=0
+ $Y2=0
cc_420 N_A_110_70#_M1020_g N_A_440_413#_c_909_n 0.00164914f $X=2.625 $Y=1.025
+ $X2=0 $Y2=0
cc_421 N_A_110_70#_M1011_g N_A_440_413#_c_915_n 7.74111e-19 $X=1.54 $Y=1.025
+ $X2=0 $Y2=0
cc_422 N_A_110_70#_c_536_n N_A_440_413#_c_915_n 0.00410514f $X=2.55 $Y=0.18
+ $X2=0 $Y2=0
cc_423 N_A_110_70#_M1020_g N_A_440_413#_c_915_n 0.00437928f $X=2.625 $Y=1.025
+ $X2=0 $Y2=0
cc_424 N_A_110_70#_M1011_g N_VGND_c_947_n 0.0241986f $X=1.54 $Y=1.025 $X2=0
+ $Y2=0
cc_425 N_A_110_70#_c_536_n N_VGND_c_947_n 0.025695f $X=2.55 $Y=0.18 $X2=0 $Y2=0
cc_426 N_A_110_70#_M1020_g N_VGND_c_947_n 0.0114212f $X=2.625 $Y=1.025 $X2=0
+ $Y2=0
cc_427 N_A_110_70#_c_539_n N_VGND_c_948_n 0.0451286f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_428 N_A_110_70#_c_539_n N_VGND_c_949_n 0.00834065f $X=5.43 $Y=0.18 $X2=0
+ $Y2=0
cc_429 N_A_110_70#_c_537_n N_VGND_c_951_n 0.00950362f $X=1.615 $Y=0.18 $X2=0
+ $Y2=0
cc_430 N_A_110_70#_c_543_n N_VGND_c_951_n 0.00915028f $X=0.69 $Y=0.565 $X2=0
+ $Y2=0
cc_431 N_A_110_70#_c_536_n N_VGND_c_953_n 0.0551589f $X=2.55 $Y=0.18 $X2=0 $Y2=0
cc_432 N_A_110_70#_c_539_n N_VGND_c_954_n 0.0407618f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_433 N_A_110_70#_c_536_n N_VGND_c_957_n 0.023216f $X=2.55 $Y=0.18 $X2=0 $Y2=0
cc_434 N_A_110_70#_c_537_n N_VGND_c_957_n 0.0115931f $X=1.615 $Y=0.18 $X2=0
+ $Y2=0
cc_435 N_A_110_70#_c_539_n N_VGND_c_957_n 0.0862653f $X=5.43 $Y=0.18 $X2=0 $Y2=0
cc_436 N_A_110_70#_c_542_n N_VGND_c_957_n 0.00856335f $X=2.625 $Y=0.18 $X2=0
+ $Y2=0
cc_437 N_A_110_70#_c_543_n N_VGND_c_957_n 0.00923605f $X=0.69 $Y=0.565 $X2=0
+ $Y2=0
cc_438 N_A_1158_93#_M1013_g N_A_957_379#_c_744_n 0.0142464f $X=5.865 $Y=0.805
+ $X2=0 $Y2=0
cc_439 N_A_1158_93#_c_673_n N_A_957_379#_c_744_n 0.00208611f $X=7.685 $Y=1.25
+ $X2=0 $Y2=0
cc_440 N_A_1158_93#_c_676_n N_A_957_379#_c_744_n 0.00199024f $X=6.737 $Y=1.795
+ $X2=0 $Y2=0
cc_441 N_A_1158_93#_M1013_g N_A_957_379#_c_745_n 0.00650191f $X=5.865 $Y=0.805
+ $X2=0 $Y2=0
cc_442 N_A_1158_93#_c_673_n N_A_957_379#_c_745_n 0.0227271f $X=7.685 $Y=1.25
+ $X2=0 $Y2=0
cc_443 N_A_1158_93#_c_675_n N_A_957_379#_c_745_n 5.85455e-19 $X=6.54 $Y=1.71
+ $X2=0 $Y2=0
cc_444 N_A_1158_93#_c_676_n N_A_957_379#_c_745_n 0.0108782f $X=6.737 $Y=1.795
+ $X2=0 $Y2=0
cc_445 N_A_1158_93#_c_677_n N_A_957_379#_c_745_n 0.0205903f $X=5.955 $Y=1.57
+ $X2=0 $Y2=0
cc_446 N_A_1158_93#_M1006_g N_A_957_379#_M1014_g 0.0133316f $X=5.865 $Y=2.105
+ $X2=0 $Y2=0
cc_447 N_A_1158_93#_c_673_n N_A_957_379#_M1014_g 0.0057023f $X=7.685 $Y=1.25
+ $X2=0 $Y2=0
cc_448 N_A_1158_93#_c_675_n N_A_957_379#_M1014_g 0.0154713f $X=6.54 $Y=1.71
+ $X2=0 $Y2=0
cc_449 N_A_1158_93#_c_676_n N_A_957_379#_M1014_g 0.0015192f $X=6.737 $Y=1.795
+ $X2=0 $Y2=0
cc_450 N_A_1158_93#_c_683_n N_A_957_379#_M1014_g 0.00756008f $X=6.625 $Y=2.04
+ $X2=0 $Y2=0
cc_451 N_A_1158_93#_c_684_n N_A_957_379#_M1014_g 9.19115e-19 $X=5.955 $Y=1.57
+ $X2=0 $Y2=0
cc_452 N_A_1158_93#_M1013_g N_A_957_379#_c_748_n 0.0165256f $X=5.865 $Y=0.805
+ $X2=0 $Y2=0
cc_453 N_A_1158_93#_c_675_n N_A_957_379#_c_748_n 0.0102298f $X=6.54 $Y=1.71
+ $X2=0 $Y2=0
cc_454 N_A_1158_93#_c_684_n N_A_957_379#_c_748_n 0.0242145f $X=5.955 $Y=1.57
+ $X2=0 $Y2=0
cc_455 N_A_1158_93#_c_677_n N_A_957_379#_c_748_n 0.00433487f $X=5.955 $Y=1.57
+ $X2=0 $Y2=0
cc_456 N_A_1158_93#_M1013_g N_A_957_379#_c_749_n 0.0021152f $X=5.865 $Y=0.805
+ $X2=0 $Y2=0
cc_457 N_A_1158_93#_c_684_n N_A_957_379#_c_749_n 0.0124098f $X=5.955 $Y=1.57
+ $X2=0 $Y2=0
cc_458 N_A_1158_93#_M1013_g N_A_957_379#_c_751_n 7.41581e-19 $X=5.865 $Y=0.805
+ $X2=0 $Y2=0
cc_459 N_A_1158_93#_c_673_n N_A_957_379#_c_751_n 2.9563e-19 $X=7.685 $Y=1.25
+ $X2=0 $Y2=0
cc_460 N_A_1158_93#_c_675_n N_A_957_379#_c_751_n 0.0148124f $X=6.54 $Y=1.71
+ $X2=0 $Y2=0
cc_461 N_A_1158_93#_c_676_n N_A_957_379#_c_751_n 0.0395863f $X=6.737 $Y=1.795
+ $X2=0 $Y2=0
cc_462 N_A_1158_93#_c_677_n N_A_957_379#_c_751_n 3.56659e-19 $X=5.955 $Y=1.57
+ $X2=0 $Y2=0
cc_463 N_A_1158_93#_M1006_g N_VPWR_c_828_n 0.00410562f $X=5.865 $Y=2.105 $X2=0
+ $Y2=0
cc_464 N_A_1158_93#_c_675_n N_VPWR_c_828_n 0.0170061f $X=6.54 $Y=1.71 $X2=0
+ $Y2=0
cc_465 N_A_1158_93#_c_683_n N_VPWR_c_828_n 0.0293243f $X=6.625 $Y=2.04 $X2=0
+ $Y2=0
cc_466 N_A_1158_93#_c_684_n N_VPWR_c_828_n 0.0112989f $X=5.955 $Y=1.57 $X2=0
+ $Y2=0
cc_467 N_A_1158_93#_c_677_n N_VPWR_c_828_n 8.89017e-19 $X=5.955 $Y=1.57 $X2=0
+ $Y2=0
cc_468 N_A_1158_93#_c_673_n N_VPWR_c_829_n 0.00758183f $X=7.685 $Y=1.25 $X2=0
+ $Y2=0
cc_469 N_A_1158_93#_M1015_g N_VPWR_c_829_n 0.00885086f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_470 N_A_1158_93#_c_683_n N_VPWR_c_829_n 0.045297f $X=6.625 $Y=2.04 $X2=0
+ $Y2=0
cc_471 N_A_1158_93#_c_724_p N_VPWR_c_829_n 0.0253995f $X=6.822 $Y=1.462 $X2=0
+ $Y2=0
cc_472 N_A_1158_93#_c_683_n N_VPWR_c_832_n 0.0089609f $X=6.625 $Y=2.04 $X2=0
+ $Y2=0
cc_473 N_A_1158_93#_M1015_g N_VPWR_c_833_n 0.00585385f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_474 N_A_1158_93#_M1006_g N_VPWR_c_822_n 0.00373935f $X=5.865 $Y=2.105 $X2=0
+ $Y2=0
cc_475 N_A_1158_93#_M1015_g N_VPWR_c_822_n 0.012741f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_476 N_A_1158_93#_c_683_n N_VPWR_c_822_n 0.0124162f $X=6.625 $Y=2.04 $X2=0
+ $Y2=0
cc_477 N_A_1158_93#_M1007_g N_Q_c_932_n 0.030511f $X=7.685 $Y=0.655 $X2=0 $Y2=0
cc_478 N_A_1158_93#_c_676_n N_Q_c_932_n 0.00528143f $X=6.737 $Y=1.795 $X2=0
+ $Y2=0
cc_479 N_A_1158_93#_c_724_p N_Q_c_932_n 0.0318248f $X=6.822 $Y=1.462 $X2=0 $Y2=0
cc_480 N_A_1158_93#_M1013_g N_VGND_c_949_n 0.0056048f $X=5.865 $Y=0.805 $X2=0
+ $Y2=0
cc_481 N_A_1158_93#_c_673_n N_VGND_c_950_n 0.0054111f $X=7.685 $Y=1.25 $X2=0
+ $Y2=0
cc_482 N_A_1158_93#_M1007_g N_VGND_c_950_n 0.00835281f $X=7.685 $Y=0.655 $X2=0
+ $Y2=0
cc_483 N_A_1158_93#_c_676_n N_VGND_c_950_n 0.0367505f $X=6.737 $Y=1.795 $X2=0
+ $Y2=0
cc_484 N_A_1158_93#_c_724_p N_VGND_c_950_n 0.0219327f $X=6.822 $Y=1.462 $X2=0
+ $Y2=0
cc_485 N_A_1158_93#_M1013_g N_VGND_c_954_n 0.00431487f $X=5.865 $Y=0.805 $X2=0
+ $Y2=0
cc_486 N_A_1158_93#_c_676_n N_VGND_c_955_n 0.015356f $X=6.737 $Y=1.795 $X2=0
+ $Y2=0
cc_487 N_A_1158_93#_M1007_g N_VGND_c_956_n 0.00585385f $X=7.685 $Y=0.655 $X2=0
+ $Y2=0
cc_488 N_A_1158_93#_M1013_g N_VGND_c_957_n 0.00477801f $X=5.865 $Y=0.805 $X2=0
+ $Y2=0
cc_489 N_A_1158_93#_M1007_g N_VGND_c_957_n 0.012741f $X=7.685 $Y=0.655 $X2=0
+ $Y2=0
cc_490 N_A_1158_93#_c_676_n N_VGND_c_957_n 0.0162118f $X=6.737 $Y=1.795 $X2=0
+ $Y2=0
cc_491 N_A_957_379#_c_754_n N_VPWR_c_827_n 0.00606476f $X=5.195 $Y=2.04 $X2=0
+ $Y2=0
cc_492 N_A_957_379#_M1014_g N_VPWR_c_828_n 0.0195513f $X=6.41 $Y=2.315 $X2=0
+ $Y2=0
cc_493 N_A_957_379#_c_754_n N_VPWR_c_828_n 0.0149616f $X=5.195 $Y=2.04 $X2=0
+ $Y2=0
cc_494 N_A_957_379#_M1014_g N_VPWR_c_832_n 0.0035863f $X=6.41 $Y=2.315 $X2=0
+ $Y2=0
cc_495 N_A_957_379#_M1014_g N_VPWR_c_822_n 0.00401353f $X=6.41 $Y=2.315 $X2=0
+ $Y2=0
cc_496 N_A_957_379#_c_754_n N_VPWR_c_822_n 0.0083393f $X=5.195 $Y=2.04 $X2=0
+ $Y2=0
cc_497 N_A_957_379#_c_744_n N_VGND_c_949_n 0.0147957f $X=6.37 $Y=1.09 $X2=0
+ $Y2=0
cc_498 N_A_957_379#_c_748_n N_VGND_c_949_n 0.0225599f $X=6.335 $Y=1.21 $X2=0
+ $Y2=0
cc_499 N_A_957_379#_c_763_n N_VGND_c_954_n 0.00712872f $X=5.3 $Y=0.805 $X2=0
+ $Y2=0
cc_500 N_A_957_379#_c_744_n N_VGND_c_955_n 0.00425533f $X=6.37 $Y=1.09 $X2=0
+ $Y2=0
cc_501 N_A_957_379#_c_744_n N_VGND_c_957_n 0.0051163f $X=6.37 $Y=1.09 $X2=0
+ $Y2=0
cc_502 N_A_957_379#_c_763_n N_VGND_c_957_n 0.010251f $X=5.3 $Y=0.805 $X2=0 $Y2=0
cc_503 N_VPWR_c_822_n N_Q_M1015_d 0.0026734f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_504 N_VPWR_c_829_n N_Q_c_932_n 7.36261e-19 $X=7.47 $Y=1.99 $X2=0 $Y2=0
cc_505 N_VPWR_c_833_n N_Q_c_932_n 0.0188755f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_506 N_VPWR_c_822_n N_Q_c_932_n 0.0111968f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_507 N_A_440_413#_c_915_n N_VGND_c_947_n 0.0120979f $X=2.41 $Y=1.025 $X2=0
+ $Y2=0
cc_508 N_A_440_413#_c_915_n N_VGND_c_957_n 0.0108188f $X=2.41 $Y=1.025 $X2=0
+ $Y2=0
cc_509 N_Q_c_932_n N_VGND_c_950_n 0.00153983f $X=7.9 $Y=0.42 $X2=0 $Y2=0
cc_510 N_Q_c_932_n N_VGND_c_956_n 0.0188755f $X=7.9 $Y=0.42 $X2=0 $Y2=0
cc_511 N_Q_M1007_d N_VGND_c_957_n 0.0026734f $X=7.76 $Y=0.235 $X2=0 $Y2=0
cc_512 N_Q_c_932_n N_VGND_c_957_n 0.0111968f $X=7.9 $Y=0.42 $X2=0 $Y2=0
