# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__buf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.390000 1.200000 2.785000 1.540000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.075000 1.855000 1.245000 ;
        RECT 0.095000 1.245000 0.510000 1.775000 ;
        RECT 0.095000 1.775000 1.855000 1.945000 ;
        RECT 0.805000 0.255000 0.995000 1.075000 ;
        RECT 0.805000 1.945000 0.995000 3.075000 ;
        RECT 1.665000 0.255000 1.855000 1.075000 ;
        RECT 1.665000 1.945000 1.855000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.305000  0.085000 0.635000 0.905000 ;
      RECT 0.305000  2.115000 0.635000 3.245000 ;
      RECT 0.700000  1.415000 2.220000 1.605000 ;
      RECT 1.165000  0.085000 1.495000 0.905000 ;
      RECT 1.165000  2.115000 1.495000 3.245000 ;
      RECT 2.025000  0.085000 2.355000 0.690000 ;
      RECT 2.025000  0.860000 2.785000 1.030000 ;
      RECT 2.025000  1.030000 2.220000 1.415000 ;
      RECT 2.025000  1.605000 2.220000 1.755000 ;
      RECT 2.025000  1.755000 2.785000 1.925000 ;
      RECT 2.025000  2.095000 2.355000 3.245000 ;
      RECT 2.525000  0.255000 2.785000 0.860000 ;
      RECT 2.525000  1.925000 2.785000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_lp__buf_4
END LIBRARY
