* File: sky130_fd_sc_lp__and4bb_2.pex.spice
* Created: Wed Sep  2 09:34:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4BB_2%A_N 3 5 7 9 13
c24 7 0 1.1515e-19 $X=0.54 $Y=2.045
r25 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.51 $X2=0.385 $Y2=1.51
r26 9 13 3.98693 $w=4.63e-07 $l=1.55e-07 $layer=LI1_cond $X=0.317 $Y=1.665
+ $X2=0.317 $Y2=1.51
r27 5 12 38.8967 $w=3.59e-07 $l=2.17991e-07 $layer=POLY_cond $X=0.54 $Y=1.675
+ $X2=0.417 $Y2=1.51
r28 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.54 $Y=1.675 $X2=0.54
+ $Y2=2.045
r29 1 12 38.8967 $w=3.59e-07 $l=1.9182e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.417 $Y2=1.51
r30 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.475 $Y=1.345 $X2=0.475
+ $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_2%A_185_23# 1 2 3 12 16 18 22 24 26 28 31 35
+ 38 42 46 47 49 50
c110 38 0 1.2007e-19 $X=3.485 $Y=2.02
c111 35 0 4.80826e-20 $X=1.75 $Y=1.085
r112 49 52 7.18582 $w=4.23e-07 $l=2.65e-07 $layer=LI1_cond $X=2.602 $Y=2.02
+ $X2=2.602 $Y2=2.285
r113 49 50 6.59116 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=2.602 $Y=2.02
+ $X2=2.602 $Y2=1.935
r114 45 47 4.38167 $w=5.03e-07 $l=1.85e-07 $layer=LI1_cond $X=2.29 $Y=0.922
+ $X2=2.475 $Y2=0.922
r115 45 46 9.14837 $w=5.03e-07 $l=1.65e-07 $layer=LI1_cond $X=2.29 $Y=0.922
+ $X2=2.125 $Y2=0.922
r116 40 42 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=3.61 $Y=2.105
+ $X2=3.61 $Y2=2.285
r117 39 49 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=2.815 $Y=2.02
+ $X2=2.602 $Y2=2.02
r118 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.485 $Y=2.02
+ $X2=3.61 $Y2=2.105
r119 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.485 $Y=2.02
+ $X2=2.815 $Y2=2.02
r120 36 47 7.21919 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=2.475 $Y=1.175
+ $X2=2.475 $Y2=0.922
r121 36 50 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.475 $Y=1.175
+ $X2=2.475 $Y2=1.935
r122 35 46 23.1061 $w=1.78e-07 $l=3.75e-07 $layer=LI1_cond $X=1.75 $Y=1.085
+ $X2=2.125 $Y2=1.085
r123 32 54 12.0836 $w=3.59e-07 $l=9e-08 $layer=POLY_cond $X=1.552 $Y=1.45
+ $X2=1.552 $Y2=1.36
r124 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=1.45 $X2=1.585 $Y2=1.45
r125 29 35 7.17723 $w=1.8e-07 $l=1.74284e-07 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.75 $Y2=1.085
r126 29 31 11.7378 $w=2.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.615 $Y=1.175
+ $X2=1.615 $Y2=1.45
r127 24 32 38.8967 $w=3.59e-07 $l=1.9139e-07 $layer=POLY_cond $X=1.495 $Y=1.615
+ $X2=1.552 $Y2=1.45
r128 24 26 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.495 $Y=1.615
+ $X2=1.495 $Y2=2.465
r129 20 54 26.8132 $w=3.59e-07 $l=1.55029e-07 $layer=POLY_cond $X=1.43 $Y=1.285
+ $X2=1.552 $Y2=1.36
r130 20 22 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.43 $Y=1.285
+ $X2=1.43 $Y2=0.665
r131 19 28 5.30422 $w=1.5e-07 $l=1.08e-07 $layer=POLY_cond $X=1.14 $Y=1.36
+ $X2=1.032 $Y2=1.36
r132 18 54 23.2387 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=1.355 $Y=1.36
+ $X2=1.552 $Y2=1.36
r133 18 19 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.355 $Y=1.36
+ $X2=1.14 $Y2=1.36
r134 14 28 20.4101 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.065 $Y=1.435
+ $X2=1.032 $Y2=1.36
r135 14 16 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=1.065 $Y=1.435
+ $X2=1.065 $Y2=2.465
r136 10 28 20.4101 $w=1.5e-07 $l=8.95824e-08 $layer=POLY_cond $X=1 $Y=1.285
+ $X2=1.032 $Y2=1.36
r137 10 12 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1 $Y=1.285 $X2=1
+ $Y2=0.665
r138 3 42 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=2.075 $X2=3.62 $Y2=2.285
r139 2 52 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=2.075 $X2=2.72 $Y2=2.285
r140 1 45 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.625 $X2=2.29 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_2%A_27_133# 1 2 9 13 15 16 19 21 25 26 28 29
+ 32 33 34 37 40
c102 13 0 1.2007e-19 $X=2.505 $Y=2.285
r103 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.51 $X2=2.125 $Y2=1.51
r104 35 37 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=2.09 $Y=1.795
+ $X2=2.09 $Y2=1.51
r105 33 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.96 $Y=1.88
+ $X2=2.09 $Y2=1.795
r106 33 34 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.96 $Y=1.88
+ $X2=1.785 $Y2=1.88
r107 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.7 $Y=1.965
+ $X2=1.785 $Y2=1.88
r108 31 32 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.7 $Y=1.965
+ $X2=1.7 $Y2=2.385
r109 30 40 2.99104 $w=3.17e-07 $l=2.72202e-07 $layer=LI1_cond $X=0.9 $Y=2.47
+ $X2=0.815 $Y2=2.237
r110 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.615 $Y=2.47
+ $X2=1.7 $Y2=2.385
r111 29 30 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.615 $Y=2.47
+ $X2=0.9 $Y2=2.47
r112 28 40 3.66292 $w=1.7e-07 $l=3.17e-07 $layer=LI1_cond $X=0.815 $Y=1.92
+ $X2=0.815 $Y2=2.237
r113 27 28 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.815 $Y=1.245
+ $X2=0.815 $Y2=1.92
r114 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.73 $Y=1.16
+ $X2=0.815 $Y2=1.245
r115 25 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.73 $Y=1.16
+ $X2=0.355 $Y2=1.16
r116 21 40 2.99104 $w=3.17e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.73 $Y=2.152
+ $X2=0.815 $Y2=2.237
r117 21 23 10.4175 $w=4.63e-07 $l=4.05e-07 $layer=LI1_cond $X=0.73 $Y=2.152
+ $X2=0.325 $Y2=2.152
r118 17 26 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=1.075
+ $X2=0.355 $Y2=1.16
r119 17 19 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=0.225 $Y=1.075
+ $X2=0.225 $Y2=0.875
r120 15 38 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.43 $Y=1.51
+ $X2=2.125 $Y2=1.51
r121 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.43 $Y=1.51
+ $X2=2.505 $Y2=1.51
r122 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=1.675
+ $X2=2.505 $Y2=1.51
r123 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.505 $Y=1.675
+ $X2=2.505 $Y2=2.285
r124 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=1.345
+ $X2=2.505 $Y2=1.51
r125 7 9 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.505 $Y=1.345
+ $X2=2.505 $Y2=0.835
r126 2 23 600 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=1.835 $X2=0.325 $Y2=2.085
r127 1 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.665 $X2=0.26 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_2%A_558_99# 1 2 9 12 15 16 17 20 21 23 24 27
+ 31 33
r75 29 33 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.52 $Y=1.765 $X2=4.52
+ $Y2=1.675
r76 29 31 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=4.52 $Y=1.765
+ $X2=4.52 $Y2=2.285
r77 25 33 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.52 $Y=1.585 $X2=4.52
+ $Y2=1.675
r78 25 27 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=4.52 $Y=1.585
+ $X2=4.52 $Y2=0.92
r79 23 33 3.59259 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=1.675
+ $X2=4.52 $Y2=1.675
r80 23 24 76.096 $w=1.78e-07 $l=1.235e-06 $layer=LI1_cond $X=4.355 $Y=1.675
+ $X2=3.12 $Y2=1.675
r81 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.955
+ $Y=1.33 $X2=2.955 $Y2=1.33
r82 18 24 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.955 $Y=1.585
+ $X2=3.12 $Y2=1.675
r83 18 20 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.955 $Y=1.585
+ $X2=2.955 $Y2=1.33
r84 16 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.955 $Y=1.67
+ $X2=2.955 $Y2=1.33
r85 16 17 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.67
+ $X2=2.955 $Y2=1.835
r86 15 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.955 $Y=1.165
+ $X2=2.955 $Y2=1.33
r87 12 17 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.935 $Y=2.285
+ $X2=2.935 $Y2=1.835
r88 9 15 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.865 $Y=0.835
+ $X2=2.865 $Y2=1.165
r89 2 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=2.075 $X2=4.52 $Y2=2.285
r90 1 27 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.625 $X2=4.52 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_2%C 3 6 7 10
r33 10 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=2.855
+ $X2=3.42 $Y2=2.69
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=2.855 $X2=3.42 $Y2=2.855
r35 7 11 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.6 $Y=2.855 $X2=3.42
+ $Y2=2.855
r36 6 12 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.405 $Y=2.285
+ $X2=3.405 $Y2=2.69
r37 3 6 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=3.405 $Y=0.835
+ $X2=3.405 $Y2=2.285
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_2%D 3 6 8 9 13 15
c40 9 0 1.84762e-19 $X=4.08 $Y=1.295
r41 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.32
+ $X2=3.855 $Y2=1.485
r42 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.32
+ $X2=3.855 $Y2=1.155
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.855
+ $Y=1.32 $X2=3.855 $Y2=1.32
r44 9 14 11.034 $w=2.33e-07 $l=2.25e-07 $layer=LI1_cond $X=4.08 $Y=1.297
+ $X2=3.855 $Y2=1.297
r45 8 14 12.5052 $w=2.33e-07 $l=2.55e-07 $layer=LI1_cond $X=3.6 $Y=1.297
+ $X2=3.855 $Y2=1.297
r46 6 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.87 $Y=2.285 $X2=3.87
+ $Y2=1.485
r47 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.765 $Y=0.835
+ $X2=3.765 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_2%B_N 4 7 12 13 14 15 16 20
c44 20 0 2.10206e-19 $X=4.305 $Y=0.35
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.305
+ $Y=0.35 $X2=4.305 $Y2=0.35
r46 16 21 7.43982 $w=3.93e-07 $l=2.55e-07 $layer=LI1_cond $X=4.56 $Y=0.452
+ $X2=4.305 $Y2=0.452
r47 15 21 6.56455 $w=3.93e-07 $l=2.25e-07 $layer=LI1_cond $X=4.08 $Y=0.452
+ $X2=4.305 $Y2=0.452
r48 13 14 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.32 $Y=1.725
+ $X2=4.32 $Y2=1.875
r49 12 13 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.335 $Y=1.305
+ $X2=4.335 $Y2=1.725
r50 11 12 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.32 $Y=1.155
+ $X2=4.32 $Y2=1.305
r51 7 14 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.305 $Y=2.285
+ $X2=4.305 $Y2=1.875
r52 4 11 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.305 $Y=0.835
+ $X2=4.305 $Y2=1.155
r53 1 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=0.515
+ $X2=4.305 $Y2=0.35
r54 1 4 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.305 $Y=0.515
+ $X2=4.305 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_2%VPWR 1 2 3 4 17 21 24 27 32 35 36 37 39 48
+ 54 55 58 61 68
r74 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r75 61 62 6.43606 $w=6.73e-07 $l=1.05e-07 $layer=LI1_cond $X=1.882 $Y=2.83
+ $X2=1.882 $Y2=2.725
r76 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 55 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r79 52 68 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.045 $Y2=3.33
r80 52 54 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 51 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r82 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r83 48 68 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.045 $Y2=3.33
r84 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.6 $Y2=3.33
r85 47 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r86 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 44 46 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.22 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r89 43 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r90 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r91 40 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.85 $Y2=3.33
r92 40 42 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.2 $Y2=3.33
r93 39 44 9.08255 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=1.882 $Y=3.33
+ $X2=2.22 $Y2=3.33
r94 39 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r95 39 61 8.85984 $w=6.73e-07 $l=5e-07 $layer=LI1_cond $X=1.882 $Y=3.33
+ $X2=1.882 $Y2=2.83
r96 39 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r97 37 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r98 37 65 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 35 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.985 $Y=3.33
+ $X2=3.07 $Y2=3.33
r101 34 50 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.6 $Y2=3.33
r102 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.07 $Y2=3.33
r103 29 32 3.76308 $w=2.43e-07 $l=8e-08 $layer=LI1_cond $X=3.07 $Y=2.397
+ $X2=3.15 $Y2=2.397
r104 25 68 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=3.245
+ $X2=4.045 $Y2=3.33
r105 25 27 39.5123 $w=2.78e-07 $l=9.6e-07 $layer=LI1_cond $X=4.045 $Y=3.245
+ $X2=4.045 $Y2=2.285
r106 24 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=3.245
+ $X2=3.07 $Y2=3.33
r107 23 29 2.87745 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=3.07 $Y=2.52
+ $X2=3.07 $Y2=2.397
r108 23 24 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.07 $Y=2.52
+ $X2=3.07 $Y2=3.245
r109 21 62 18.4826 $w=2.63e-07 $l=4.25e-07 $layer=LI1_cond $X=2.087 $Y=2.3
+ $X2=2.087 $Y2=2.725
r110 15 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=3.245
+ $X2=0.85 $Y2=3.33
r111 15 17 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.85 $Y=3.245
+ $X2=0.85 $Y2=2.83
r112 4 27 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=2.075 $X2=4.085 $Y2=2.285
r113 3 32 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=2.075 $X2=3.15 $Y2=2.37
r114 2 61 600 $w=1.7e-07 $l=1.0627e-06 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.835 $X2=1.71 $Y2=2.83
r115 2 21 600 $w=1.7e-07 $l=7.15682e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.835 $X2=2.09 $Y2=2.3
r116 1 17 600 $w=1.7e-07 $l=1.10628e-06 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.835 $X2=0.85 $Y2=2.83
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_2%X 1 2 11 13 14 18
c26 18 0 1.1515e-19 $X=1.215 $Y=0.42
r27 13 14 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.665
r28 13 18 43.8429 $w=2.28e-07 $l=8.75e-07 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=0.42
r29 8 14 13.5287 $w=2.28e-07 $l=2.7e-07 $layer=LI1_cond $X=1.195 $Y=1.935
+ $X2=1.195 $Y2=1.665
r30 7 11 3.49849 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=2.075
+ $X2=1.28 $Y2=2.075
r31 7 8 1.89134 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=1.195 $Y=2.075
+ $X2=1.195 $Y2=1.935
r32 2 11 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.835 $X2=1.28 $Y2=2.1
r33 1 18 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.245 $X2=1.215 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_2%VGND 1 2 3 12 18 21 22 24 26 28 33 38 48 49
+ 52 55 58
c68 24 0 2.54439e-20 $X=3.98 $Y=0.905
r69 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r70 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r71 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r72 49 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r73 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r74 46 58 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.775 $Y=0 $X2=3.605
+ $Y2=0
r75 46 48 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=3.775 $Y=0 $X2=4.56
+ $Y2=0
r76 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r77 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r78 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r79 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r80 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r81 39 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.645
+ $Y2=0
r82 39 41 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=2.16
+ $Y2=0
r83 38 58 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.605
+ $Y2=0
r84 38 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.12
+ $Y2=0
r85 37 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r86 37 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r87 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r88 34 52 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.717
+ $Y2=0
r89 34 36 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.2
+ $Y2=0
r90 33 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=1.645
+ $Y2=0
r91 33 36 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=1.2
+ $Y2=0
r92 31 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r93 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r94 28 52 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.717
+ $Y2=0
r95 28 30 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r96 26 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r97 26 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r98 22 24 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=3.775 $Y=0.915
+ $X2=3.98 $Y2=0.915
r99 21 22 7.55181 $w=1.9e-07 $l=2.1225e-07 $layer=LI1_cond $X=3.605 $Y=0.82
+ $X2=3.775 $Y2=0.915
r100 20 58 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=0.085
+ $X2=3.605 $Y2=0
r101 20 21 24.9131 $w=3.38e-07 $l=7.35e-07 $layer=LI1_cond $X=3.605 $Y=0.085
+ $X2=3.605 $Y2=0.82
r102 16 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0
r103 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.645 $Y=0.085
+ $X2=1.645 $Y2=0.39
r104 12 14 12.8714 $w=3.83e-07 $l=4.3e-07 $layer=LI1_cond $X=0.717 $Y=0.39
+ $X2=0.717 $Y2=0.82
r105 10 52 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.717 $Y=0.085
+ $X2=0.717 $Y2=0
r106 10 12 9.12974 $w=3.83e-07 $l=3.05e-07 $layer=LI1_cond $X=0.717 $Y=0.085
+ $X2=0.717 $Y2=0.39
r107 3 24 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=3.84
+ $Y=0.625 $X2=3.98 $Y2=0.905
r108 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.245 $X2=1.645 $Y2=0.39
r109 1 14 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.665 $X2=0.69 $Y2=0.82
r110 1 12 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.665 $X2=0.785 $Y2=0.39
.ends

