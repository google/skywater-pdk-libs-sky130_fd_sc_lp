* File: sky130_fd_sc_lp__buf_8.pex.spice
* Created: Fri Aug 28 10:10:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUF_8%A 3 7 11 15 19 23 27 30 31 42 44 50 53
c62 27 0 1.64844e-19 $X=1.18 $Y=1.48
r63 44 50 1.0795 $w=3.93e-07 $l=3.7e-08 $layer=LI1_cond $X=0.683 $Y=1.377
+ $X2=0.72 $Y2=1.377
r64 39 53 4.28224 $w=3.93e-07 $l=4e-08 $layer=LI1_cond $X=0.84 $Y=1.377 $X2=0.88
+ $Y2=1.377
r65 38 40 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=0.84 $Y=1.48
+ $X2=0.905 $Y2=1.48
r66 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.48 $X2=0.84 $Y2=1.48
r67 35 38 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=0.475 $Y=1.48
+ $X2=0.84 $Y2=1.48
r68 31 39 2.80087 $w=3.93e-07 $l=9.6e-08 $layer=LI1_cond $X=0.744 $Y=1.377
+ $X2=0.84 $Y2=1.377
r69 31 50 0.700219 $w=3.93e-07 $l=2.4e-08 $layer=LI1_cond $X=0.744 $Y=1.377
+ $X2=0.72 $Y2=1.377
r70 31 44 0.700219 $w=3.93e-07 $l=2.4e-08 $layer=LI1_cond $X=0.659 $Y=1.377
+ $X2=0.683 $Y2=1.377
r71 30 31 12.2246 $w=3.93e-07 $l=4.19e-07 $layer=LI1_cond $X=0.24 $Y=1.377
+ $X2=0.659 $Y2=1.377
r72 28 42 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=1.18 $Y=1.48
+ $X2=1.335 $Y2=1.48
r73 28 40 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=1.18 $Y=1.48
+ $X2=0.905 $Y2=1.48
r74 27 53 17.512 $w=1.88e-07 $l=3e-07 $layer=LI1_cond $X=1.18 $Y=1.48 $X2=0.88
+ $Y2=1.48
r75 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.48 $X2=1.18 $Y2=1.48
r76 21 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.645
+ $X2=1.335 $Y2=1.48
r77 21 23 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.335 $Y=1.645
+ $X2=1.335 $Y2=2.465
r78 17 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.315
+ $X2=1.335 $Y2=1.48
r79 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.335 $Y=1.315
+ $X2=1.335 $Y2=0.655
r80 13 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.645
+ $X2=0.905 $Y2=1.48
r81 13 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.905 $Y=1.645
+ $X2=0.905 $Y2=2.465
r82 9 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.315
+ $X2=0.905 $Y2=1.48
r83 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.905 $Y=1.315
+ $X2=0.905 $Y2=0.655
r84 5 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.645
+ $X2=0.475 $Y2=1.48
r85 5 7 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.475 $Y=1.645
+ $X2=0.475 $Y2=2.465
r86 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.315
+ $X2=0.475 $Y2=1.48
r87 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.475 $Y=1.315
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_8%A_27_47# 1 2 3 4 15 19 23 27 31 35 39 43 47 51
+ 55 59 63 67 71 75 79 83 87 88 89 90 93 97 101 103 106 108 114 117 119 120 131
c192 131 0 1.64844e-19 $X=4.775 $Y=1.48
r193 128 129 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.915 $Y=1.48
+ $X2=4.345 $Y2=1.48
r194 127 128 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.485 $Y=1.48
+ $X2=3.915 $Y2=1.48
r195 126 127 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.055 $Y=1.48
+ $X2=3.485 $Y2=1.48
r196 125 126 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.625 $Y=1.48
+ $X2=3.055 $Y2=1.48
r197 124 125 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.195 $Y=1.48
+ $X2=2.625 $Y2=1.48
r198 117 118 11.0176 $w=2.27e-07 $l=2.05e-07 $layer=LI1_cond $X=1.12 $Y=0.925
+ $X2=1.12 $Y2=1.13
r199 115 131 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=4.575 $Y=1.48
+ $X2=4.775 $Y2=1.48
r200 115 129 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=4.575 $Y=1.48
+ $X2=4.345 $Y2=1.48
r201 114 115 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=4.575
+ $Y=1.48 $X2=4.575 $Y2=1.48
r202 112 124 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.855 $Y=1.48
+ $X2=2.195 $Y2=1.48
r203 112 121 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.855 $Y=1.48
+ $X2=1.765 $Y2=1.48
r204 111 114 167.596 $w=1.78e-07 $l=2.72e-06 $layer=LI1_cond $X=1.855 $Y=1.485
+ $X2=4.575 $Y2=1.485
r205 111 112 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=1.855
+ $Y=1.48 $X2=1.855 $Y2=1.48
r206 109 120 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=1.485
+ $X2=1.61 $Y2=1.485
r207 109 111 9.85859 $w=1.78e-07 $l=1.6e-07 $layer=LI1_cond $X=1.695 $Y=1.485
+ $X2=1.855 $Y2=1.485
r208 107 120 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.61 $Y=1.575
+ $X2=1.61 $Y2=1.485
r209 107 108 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.61 $Y=1.575
+ $X2=1.61 $Y2=1.745
r210 106 120 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.61 $Y=1.395
+ $X2=1.61 $Y2=1.485
r211 105 106 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.61 $Y=1.215
+ $X2=1.61 $Y2=1.395
r212 104 119 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=1.835
+ $X2=1.12 $Y2=1.835
r213 103 108 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.525 $Y=1.835
+ $X2=1.61 $Y2=1.745
r214 103 104 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=1.525 $Y=1.835
+ $X2=1.25 $Y2=1.835
r215 102 118 2.43258 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=1.13
+ $X2=1.12 $Y2=1.13
r216 101 105 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.525 $Y=1.13
+ $X2=1.61 $Y2=1.215
r217 101 102 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.525 $Y=1.13
+ $X2=1.25 $Y2=1.13
r218 97 99 32.8003 $w=2.58e-07 $l=7.4e-07 $layer=LI1_cond $X=1.12 $Y=2.075
+ $X2=1.12 $Y2=2.815
r219 95 119 0.0585112 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=1.12 $Y=1.925
+ $X2=1.12 $Y2=1.835
r220 95 97 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.12 $Y=1.925
+ $X2=1.12 $Y2=2.075
r221 91 117 4.21708 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.84
+ $X2=1.12 $Y2=0.925
r222 91 93 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.12 $Y=0.84
+ $X2=1.12 $Y2=0.47
r223 89 119 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=1.835
+ $X2=1.12 $Y2=1.835
r224 89 90 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=0.99 $Y=1.835
+ $X2=0.39 $Y2=1.835
r225 87 117 2.43258 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=0.925
+ $X2=1.12 $Y2=0.925
r226 87 88 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.99 $Y=0.925
+ $X2=0.39 $Y2=0.925
r227 83 85 28.9087 $w=2.93e-07 $l=7.4e-07 $layer=LI1_cond $X=0.242 $Y=2.075
+ $X2=0.242 $Y2=2.815
r228 81 90 7.34943 $w=1.8e-07 $l=1.87681e-07 $layer=LI1_cond $X=0.242 $Y=1.925
+ $X2=0.39 $Y2=1.835
r229 81 83 5.85988 $w=2.93e-07 $l=1.5e-07 $layer=LI1_cond $X=0.242 $Y=1.925
+ $X2=0.242 $Y2=2.075
r230 77 88 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=0.242 $Y=0.84
+ $X2=0.39 $Y2=0.925
r231 77 79 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=0.84
+ $X2=0.242 $Y2=0.47
r232 73 131 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.775 $Y=1.645
+ $X2=4.775 $Y2=1.48
r233 73 75 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=4.775 $Y=1.645
+ $X2=4.775 $Y2=2.465
r234 69 131 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.775 $Y=1.315
+ $X2=4.775 $Y2=1.48
r235 69 71 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.775 $Y=1.315
+ $X2=4.775 $Y2=0.655
r236 65 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.645
+ $X2=4.345 $Y2=1.48
r237 65 67 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=4.345 $Y=1.645
+ $X2=4.345 $Y2=2.465
r238 61 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.315
+ $X2=4.345 $Y2=1.48
r239 61 63 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.345 $Y=1.315
+ $X2=4.345 $Y2=0.655
r240 57 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.645
+ $X2=3.915 $Y2=1.48
r241 57 59 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.915 $Y=1.645
+ $X2=3.915 $Y2=2.465
r242 53 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.315
+ $X2=3.915 $Y2=1.48
r243 53 55 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.915 $Y=1.315
+ $X2=3.915 $Y2=0.655
r244 49 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.645
+ $X2=3.485 $Y2=1.48
r245 49 51 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.485 $Y=1.645
+ $X2=3.485 $Y2=2.465
r246 45 127 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.315
+ $X2=3.485 $Y2=1.48
r247 45 47 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.485 $Y=1.315
+ $X2=3.485 $Y2=0.655
r248 41 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.645
+ $X2=3.055 $Y2=1.48
r249 41 43 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.055 $Y=1.645
+ $X2=3.055 $Y2=2.465
r250 37 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.315
+ $X2=3.055 $Y2=1.48
r251 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.055 $Y=1.315
+ $X2=3.055 $Y2=0.655
r252 33 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.645
+ $X2=2.625 $Y2=1.48
r253 33 35 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.625 $Y=1.645
+ $X2=2.625 $Y2=2.465
r254 29 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.315
+ $X2=2.625 $Y2=1.48
r255 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.625 $Y=1.315
+ $X2=2.625 $Y2=0.655
r256 25 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.645
+ $X2=2.195 $Y2=1.48
r257 25 27 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.195 $Y=1.645
+ $X2=2.195 $Y2=2.465
r258 21 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.315
+ $X2=2.195 $Y2=1.48
r259 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.195 $Y=1.315
+ $X2=2.195 $Y2=0.655
r260 17 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.645
+ $X2=1.765 $Y2=1.48
r261 17 19 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.765 $Y=1.645
+ $X2=1.765 $Y2=2.465
r262 13 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.315
+ $X2=1.765 $Y2=1.48
r263 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.765 $Y=1.315
+ $X2=1.765 $Y2=0.655
r264 4 99 400 $w=1.7e-07 $l=1.04766e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.815
r265 4 97 400 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.075
r266 3 85 400 $w=1.7e-07 $l=1.04062e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.815
r267 3 83 400 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.075
r268 2 93 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.47
r269 1 79 91 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_8%VPWR 1 2 3 4 5 6 21 27 33 39 43 47 51 53 58 59
+ 61 62 63 64 65 67 82 88 91 95
r84 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 86 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r88 86 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r89 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 83 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.26 $Y=3.33 $X2=4.13
+ $Y2=3.33
r91 83 85 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.26 $Y=3.33 $X2=4.56
+ $Y2=3.33
r92 82 94 3.8143 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=4.86 $Y=3.33 $X2=5.07
+ $Y2=3.33
r93 82 85 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.86 $Y=3.33 $X2=4.56
+ $Y2=3.33
r94 81 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r96 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r97 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 75 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r99 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r100 72 88 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=0.69 $Y2=3.33
r101 72 74 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=3.33
+ $X2=1.2 $Y2=3.33
r102 70 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r104 67 88 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.69 $Y2=3.33
r105 67 69 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r106 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r107 65 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 63 80 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=3.12 $Y2=3.33
r109 63 64 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=3.272 $Y2=3.33
r110 61 77 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.16 $Y2=3.33
r111 61 62 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.275 $Y=3.33
+ $X2=2.405 $Y2=3.33
r112 60 80 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=3.12 $Y2=3.33
r113 60 62 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=2.405 $Y2=3.33
r114 58 74 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.42 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 58 59 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=1.42 $Y=3.33
+ $X2=1.557 $Y2=3.33
r116 57 77 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 57 59 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.557 $Y2=3.33
r118 53 56 33.3473 $w=2.33e-07 $l=6.8e-07 $layer=LI1_cond $X=4.977 $Y=2.26
+ $X2=4.977 $Y2=2.94
r119 51 94 3.23307 $w=2.35e-07 $l=1.28662e-07 $layer=LI1_cond $X=4.977 $Y=3.245
+ $X2=5.07 $Y2=3.33
r120 51 56 14.9572 $w=2.33e-07 $l=3.05e-07 $layer=LI1_cond $X=4.977 $Y=3.245
+ $X2=4.977 $Y2=2.94
r121 47 50 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=4.13 $Y=2.26
+ $X2=4.13 $Y2=2.94
r122 45 91 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=3.33
r123 45 50 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=4.13 $Y=3.245
+ $X2=4.13 $Y2=2.94
r124 44 64 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=3.4 $Y=3.33
+ $X2=3.272 $Y2=3.33
r125 43 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4 $Y=3.33 $X2=4.13
+ $Y2=3.33
r126 43 44 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4 $Y=3.33 $X2=3.4
+ $Y2=3.33
r127 39 42 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=3.272 $Y=2.26
+ $X2=3.272 $Y2=2.94
r128 37 64 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.272 $Y=3.245
+ $X2=3.272 $Y2=3.33
r129 37 42 13.7841 $w=2.53e-07 $l=3.05e-07 $layer=LI1_cond $X=3.272 $Y=3.245
+ $X2=3.272 $Y2=2.94
r130 33 36 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=2.405 $Y=2.26
+ $X2=2.405 $Y2=2.94
r131 31 62 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=3.245
+ $X2=2.405 $Y2=3.33
r132 31 36 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=2.405 $Y=3.245
+ $X2=2.405 $Y2=2.94
r133 27 30 28.4968 $w=2.73e-07 $l=6.8e-07 $layer=LI1_cond $X=1.557 $Y=2.26
+ $X2=1.557 $Y2=2.94
r134 25 59 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.557 $Y=3.245
+ $X2=1.557 $Y2=3.33
r135 25 30 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=1.557 $Y=3.245
+ $X2=1.557 $Y2=2.94
r136 21 24 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.69 $Y=2.26
+ $X2=0.69 $Y2=2.94
r137 19 88 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r138 19 24 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.94
r139 6 56 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=4.85
+ $Y=1.835 $X2=4.99 $Y2=2.94
r140 6 53 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=4.85
+ $Y=1.835 $X2=4.99 $Y2=2.26
r141 5 50 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.835 $X2=4.13 $Y2=2.94
r142 5 47 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.835 $X2=4.13 $Y2=2.26
r143 4 42 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.94
r144 4 39 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.26
r145 3 36 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.94
r146 3 33 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.26
r147 2 30 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.94
r148 2 27 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.26
r149 1 24 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.94
r150 1 21 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_8%X 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 47 49
+ 51 55 59 63 65 69 73 77 79 81 82 83 84 85 86 87 88 93 94 96 100
r111 94 100 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=5.05 $Y=1.745
+ $X2=5.05 $Y2=1.665
r112 93 96 2.88111 $w=2.78e-07 $l=7e-08 $layer=LI1_cond $X=5.05 $Y=1.225
+ $X2=5.05 $Y2=1.295
r113 88 94 2.83462 $w=2.8e-07 $l=9e-08 $layer=LI1_cond $X=5.05 $Y=1.835 $X2=5.05
+ $Y2=1.745
r114 88 100 0.123476 $w=2.78e-07 $l=3e-09 $layer=LI1_cond $X=5.05 $Y=1.662
+ $X2=5.05 $Y2=1.665
r115 87 93 2.83462 $w=2.8e-07 $l=9e-08 $layer=LI1_cond $X=5.05 $Y=1.135 $X2=5.05
+ $Y2=1.225
r116 87 88 14.8171 $w=2.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.05 $Y=1.302
+ $X2=5.05 $Y2=1.662
r117 87 96 0.288111 $w=2.78e-07 $l=7e-09 $layer=LI1_cond $X=5.05 $Y=1.302
+ $X2=5.05 $Y2=1.295
r118 80 86 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=4.69 $Y=1.835
+ $X2=4.56 $Y2=1.835
r119 79 88 4.40942 $w=1.8e-07 $l=1.4e-07 $layer=LI1_cond $X=4.91 $Y=1.835
+ $X2=5.05 $Y2=1.835
r120 79 80 13.5556 $w=1.78e-07 $l=2.2e-07 $layer=LI1_cond $X=4.91 $Y=1.835
+ $X2=4.69 $Y2=1.835
r121 78 85 6.8302 $w=1.8e-07 $l=1.28e-07 $layer=LI1_cond $X=4.685 $Y=1.135
+ $X2=4.557 $Y2=1.135
r122 77 87 4.40942 $w=1.8e-07 $l=1.4e-07 $layer=LI1_cond $X=4.91 $Y=1.135
+ $X2=5.05 $Y2=1.135
r123 77 78 13.8636 $w=1.78e-07 $l=2.25e-07 $layer=LI1_cond $X=4.91 $Y=1.135
+ $X2=4.685 $Y2=1.135
r124 73 75 32.8003 $w=2.58e-07 $l=7.4e-07 $layer=LI1_cond $X=4.56 $Y=2.075
+ $X2=4.56 $Y2=2.815
r125 71 86 0.0585112 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=4.56 $Y=1.925
+ $X2=4.56 $Y2=1.835
r126 71 73 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=4.56 $Y=1.925
+ $X2=4.56 $Y2=2.075
r127 67 85 0.12397 $w=2.55e-07 $l=9e-08 $layer=LI1_cond $X=4.557 $Y=1.045
+ $X2=4.557 $Y2=1.135
r128 67 69 25.9865 $w=2.53e-07 $l=5.75e-07 $layer=LI1_cond $X=4.557 $Y=1.045
+ $X2=4.557 $Y2=0.47
r129 66 84 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=1.835
+ $X2=3.7 $Y2=1.835
r130 65 86 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=4.43 $Y=1.835
+ $X2=4.56 $Y2=1.835
r131 65 66 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=4.43 $Y=1.835
+ $X2=3.83 $Y2=1.835
r132 64 83 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=1.135
+ $X2=3.7 $Y2=1.135
r133 63 85 6.8302 $w=1.8e-07 $l=1.27e-07 $layer=LI1_cond $X=4.43 $Y=1.135
+ $X2=4.557 $Y2=1.135
r134 63 64 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=4.43 $Y=1.135
+ $X2=3.83 $Y2=1.135
r135 59 61 32.8003 $w=2.58e-07 $l=7.4e-07 $layer=LI1_cond $X=3.7 $Y=2.075
+ $X2=3.7 $Y2=2.815
r136 57 84 0.0585112 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=3.7 $Y=1.925 $X2=3.7
+ $Y2=1.835
r137 57 59 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=3.7 $Y=1.925
+ $X2=3.7 $Y2=2.075
r138 53 83 0.0585112 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=3.7 $Y=1.045 $X2=3.7
+ $Y2=1.135
r139 53 55 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=3.7 $Y=1.045
+ $X2=3.7 $Y2=0.47
r140 52 81 7.13466 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=2.975 $Y=1.835
+ $X2=2.84 $Y2=1.835
r141 51 84 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=1.835
+ $X2=3.7 $Y2=1.835
r142 51 52 36.6616 $w=1.78e-07 $l=5.95e-07 $layer=LI1_cond $X=3.57 $Y=1.835
+ $X2=2.975 $Y2=1.835
r143 50 82 6.8302 $w=1.8e-07 $l=1.28e-07 $layer=LI1_cond $X=2.965 $Y=1.135
+ $X2=2.837 $Y2=1.135
r144 49 83 6.93267 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=1.135
+ $X2=3.7 $Y2=1.135
r145 49 50 37.2778 $w=1.78e-07 $l=6.05e-07 $layer=LI1_cond $X=3.57 $Y=1.135
+ $X2=2.965 $Y2=1.135
r146 45 82 0.12397 $w=2.55e-07 $l=9e-08 $layer=LI1_cond $X=2.837 $Y=1.045
+ $X2=2.837 $Y2=1.135
r147 45 47 25.9865 $w=2.53e-07 $l=5.75e-07 $layer=LI1_cond $X=2.837 $Y=1.045
+ $X2=2.837 $Y2=0.47
r148 41 43 31.5855 $w=2.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.84 $Y=2.075
+ $X2=2.84 $Y2=2.815
r149 39 81 0.067832 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=2.84 $Y=1.925
+ $X2=2.84 $Y2=1.835
r150 39 41 6.40246 $w=2.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.84 $Y=1.925
+ $X2=2.84 $Y2=2.075
r151 37 82 6.8302 $w=1.8e-07 $l=1.27e-07 $layer=LI1_cond $X=2.71 $Y=1.135
+ $X2=2.837 $Y2=1.135
r152 37 38 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=2.71 $Y=1.135
+ $X2=2.11 $Y2=1.135
r153 35 81 7.13466 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=2.705 $Y=1.835
+ $X2=2.84 $Y2=1.835
r154 35 36 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=2.705 $Y=1.835
+ $X2=2.105 $Y2=1.835
r155 31 33 35.5337 $w=2.38e-07 $l=7.4e-07 $layer=LI1_cond $X=1.985 $Y=2.075
+ $X2=1.985 $Y2=2.815
r156 29 36 6.999 $w=1.8e-07 $l=1.58745e-07 $layer=LI1_cond $X=1.985 $Y=1.925
+ $X2=2.105 $Y2=1.835
r157 29 31 7.20277 $w=2.38e-07 $l=1.5e-07 $layer=LI1_cond $X=1.985 $Y=1.925
+ $X2=1.985 $Y2=2.075
r158 25 38 7.02594 $w=1.8e-07 $l=1.61861e-07 $layer=LI1_cond $X=1.987 $Y=1.045
+ $X2=2.11 $Y2=1.135
r159 25 27 27.0471 $w=2.43e-07 $l=5.75e-07 $layer=LI1_cond $X=1.987 $Y=1.045
+ $X2=1.987 $Y2=0.47
r160 8 75 400 $w=1.7e-07 $l=1.04766e-06 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.835 $X2=4.56 $Y2=2.815
r161 8 73 400 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.835 $X2=4.56 $Y2=2.075
r162 7 61 400 $w=1.7e-07 $l=1.04766e-06 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.815
r163 7 59 400 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.075
r164 6 43 400 $w=1.7e-07 $l=1.04766e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.815
r165 6 41 400 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.075
r166 5 33 400 $w=1.7e-07 $l=1.04766e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.815
r167 5 31 400 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.075
r168 4 69 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=4.42
+ $Y=0.235 $X2=4.56 $Y2=0.47
r169 3 55 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.47
r170 2 47 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.47
r171 1 27 91 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_8%VGND 1 2 3 4 5 6 21 25 29 33 35 39 41 43 46 47
+ 49 50 51 52 53 55 70 76 79 83
r84 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r85 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r86 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r87 74 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r88 74 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r89 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r90 71 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.26 $Y=0 $X2=4.13
+ $Y2=0
r91 71 73 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.26 $Y=0 $X2=4.56
+ $Y2=0
r92 70 82 4.4394 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=4.855 $Y=0 $X2=5.067
+ $Y2=0
r93 70 73 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=0 $X2=4.56
+ $Y2=0
r94 69 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r95 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r96 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r97 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r98 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r99 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r100 60 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.69
+ $Y2=0
r101 60 62 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=1.2
+ $Y2=0
r102 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r103 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r104 55 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.69
+ $Y2=0
r105 55 57 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r106 53 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r107 53 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r108 51 68 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.12
+ $Y2=0
r109 51 52 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.135 $Y=0
+ $X2=3.267 $Y2=0
r110 49 65 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.16
+ $Y2=0
r111 49 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.41
+ $Y2=0
r112 48 68 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=3.12
+ $Y2=0
r113 48 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.41
+ $Y2=0
r114 46 62 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.2
+ $Y2=0
r115 46 47 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.557
+ $Y2=0
r116 45 65 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.695 $Y=0
+ $X2=2.16 $Y2=0
r117 45 47 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.695 $Y=0
+ $X2=1.557 $Y2=0
r118 41 82 3.07827 $w=3e-07 $l=1.11781e-07 $layer=LI1_cond $X=5.005 $Y=0.085
+ $X2=5.067 $Y2=0
r119 41 43 10.9482 $w=2.98e-07 $l=2.85e-07 $layer=LI1_cond $X=5.005 $Y=0.085
+ $X2=5.005 $Y2=0.37
r120 37 79 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.085
+ $X2=4.13 $Y2=0
r121 37 39 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=4.13 $Y=0.085
+ $X2=4.13 $Y2=0.37
r122 36 52 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.267
+ $Y2=0
r123 35 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4 $Y=0 $X2=4.13
+ $Y2=0
r124 35 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4 $Y=0 $X2=3.4 $Y2=0
r125 31 52 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.267 $Y=0.085
+ $X2=3.267 $Y2=0
r126 31 33 12.3942 $w=2.63e-07 $l=2.85e-07 $layer=LI1_cond $X=3.267 $Y=0.085
+ $X2=3.267 $Y2=0.37
r127 27 50 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0
r128 27 29 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0.37
r129 23 47 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.557 $Y=0.085
+ $X2=1.557 $Y2=0
r130 23 25 11.9435 $w=2.73e-07 $l=2.85e-07 $layer=LI1_cond $X=1.557 $Y=0.085
+ $X2=1.557 $Y2=0.37
r131 19 76 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r132 19 21 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.505
r133 6 43 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=4.85
+ $Y=0.235 $X2=4.99 $Y2=0.37
r134 5 39 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.99
+ $Y=0.235 $X2=4.13 $Y2=0.37
r135 4 33 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.37
r136 3 29 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.37
r137 2 25 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.37
r138 1 21 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.505
.ends

