* File: sky130_fd_sc_lp__lsbufiso0p_lp.pex.spice
* Created: Wed Sep  2 09:59:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%VGND 1 2 3 4 29 45 49 53 57 70 71 75
+ 78 82 91 98
c183 70 0 1.58517e-19 $X=2.87 $Y=3.33
r184 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r185 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r186 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r187 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.32
+ $X2=0.72 $Y2=3.32
r188 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r189 86 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.32 $X2=6.48
+ $Y2=3.32
r190 86 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.32 $X2=5.04
+ $Y2=3.32
r191 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r192 83 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=3.33
+ $X2=5.19 $Y2=3.33
r193 83 85 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.355 $Y=3.33
+ $X2=6 $Y2=3.33
r194 82 97 3.44808 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=6.33 $Y=3.33
+ $X2=6.525 $Y2=3.33
r195 82 85 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.33 $Y=3.33 $X2=6
+ $Y2=3.33
r196 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r197 78 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=3.33
+ $X2=5.19 $Y2=3.33
r198 78 80 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=5.025 $Y=3.33
+ $X2=3.12 $Y2=3.33
r199 76 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.32
+ $X2=3.12 $Y2=3.32
r200 76 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.32
+ $X2=0.72 $Y2=3.32
r201 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r202 73 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r203 73 75 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r204 71 95 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=3.36 $Y=3.32
+ $X2=5.04 $Y2=3.32
r205 71 81 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.32
+ $X2=3.12 $Y2=3.32
r206 69 80 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.04 $Y=3.33 $X2=3.12
+ $Y2=3.33
r207 69 70 3.80956 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.04 $Y=3.33
+ $X2=2.87 $Y2=3.33
r208 64 97 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=6.48 $Y=3.415
+ $X2=6.525 $Y2=3.33
r209 59 97 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=6.48 $Y=3.245
+ $X2=6.525 $Y2=3.33
r210 55 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=3.415
+ $X2=5.19 $Y2=3.33
r211 55 57 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=5.19 $Y=3.415
+ $X2=5.19 $Y2=3.715
r212 51 70 2.88756 $w=3.3e-07 $l=8.74643e-08 $layer=LI1_cond $X=2.875 $Y=3.245
+ $X2=2.87 $Y2=3.33
r213 51 53 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=2.875 $Y=3.245
+ $X2=2.875 $Y2=2.515
r214 47 70 2.88756 $w=3.3e-07 $l=8.74643e-08 $layer=LI1_cond $X=2.865 $Y=3.415
+ $X2=2.87 $Y2=3.33
r215 47 49 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=2.865 $Y=3.415
+ $X2=2.865 $Y2=4.155
r216 43 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=3.33
r217 43 45 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=2.44
r218 42 88 3.44808 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r219 41 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r220 41 42 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.39 $Y2=3.33
r221 36 88 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.24 $Y=3.415
+ $X2=0.195 $Y2=3.33
r222 31 88 3.14896 $w=3e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.195 $Y2=3.33
r223 29 64 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=6.48 $Y=3.855
+ $X2=6.48 $Y2=3.415
r224 29 59 32.8446 $w=2.98e-07 $l=8.55e-07 $layer=LI1_cond $X=6.48 $Y=2.39
+ $X2=6.48 $Y2=3.245
r225 29 36 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=0.24 $Y=3.855
+ $X2=0.24 $Y2=3.415
r226 29 31 32.8446 $w=2.98e-07 $l=8.55e-07 $layer=LI1_cond $X=0.24 $Y=2.39
+ $X2=0.24 $Y2=3.245
r227 4 57 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=3.59 $X2=5.19 $Y2=3.715
r228 3 49 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.74
+ $Y=4.01 $X2=2.865 $Y2=4.155
r229 2 53 91 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=2 $X=2.735
+ $Y=2.23 $X2=2.875 $Y2=2.515
r230 1 45 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=2.23 $X2=0.74 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%VPB 7 9 10 11 12 13 14
r19 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=6.48 $Y=0.925
+ $X2=6.48 $Y2=1.295
r20 12 13 15.3659 $w=2.98e-07 $l=4e-07 $layer=LI1_cond $X=6.48 $Y=0.525 $X2=6.48
+ $Y2=0.925
r21 10 11 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.295
r22 9 10 15.3659 $w=2.98e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=0.525 $X2=0.24
+ $Y2=0.925
r23 7 12 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=6.395 $Y=0.32 $X2=6.48 $Y2=0.525
r24 7 9 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2 $X=0.155
+ $Y=0.32 $X2=0.24 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%DESTVPB 7 9 10 11 12 13 14
c55 7 0 6.60929e-20 $X=-0.025 $Y=4.985
r56 13 14 15.558 $w=2.98e-07 $l=4.05e-07 $layer=LI1_cond $X=6.48 $Y=5.7 $X2=6.48
+ $Y2=6.105
r57 12 13 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.48 $Y=5.365
+ $X2=6.48 $Y2=5.7
r58 10 11 15.558 $w=2.98e-07 $l=4.05e-07 $layer=LI1_cond $X=0.24 $Y=5.7 $X2=0.24
+ $Y2=6.105
r59 9 10 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=5.365
+ $X2=0.24 $Y2=5.7
r60 7 13 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=6.395 $Y=5.495 $X2=6.48 $Y2=5.7
r61 7 10 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=0.155 $Y=5.495 $X2=0.24 $Y2=5.7
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_176_987# 1 2 9 13 15 18 21 24 28 31
+ 35
c75 18 0 1.70849e-20 $X=2.24 $Y=5.355
r76 28 30 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=4.235
+ $X2=2.32 $Y2=4.4
r77 25 35 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.165 $Y=5.1
+ $X2=1.315 $Y2=5.1
r78 25 32 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.165 $Y=5.1
+ $X2=0.955 $Y2=5.1
r79 24 26 16.4603 $w=2.52e-07 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=5.1
+ $X2=1.165 $Y2=5.44
r80 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=5.1 $X2=1.165 $Y2=5.1
r81 19 31 3.70735 $w=2.5e-07 $l=2.38642e-07 $layer=LI1_cond $X=2.32 $Y=5.525
+ $X2=2.155 $Y2=5.355
r82 19 21 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.32 $Y=5.525
+ $X2=2.32 $Y2=5.55
r83 18 31 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=5.355
+ $X2=2.155 $Y2=5.355
r84 18 30 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.24 $Y=5.355
+ $X2=2.24 $Y2=4.4
r85 16 26 3.04159 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.33 $Y=5.44
+ $X2=1.165 $Y2=5.44
r86 15 31 2.76166 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=5.44
+ $X2=2.155 $Y2=5.355
r87 15 16 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.155 $Y=5.44
+ $X2=1.33 $Y2=5.44
r88 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.315 $Y=5.265
+ $X2=1.315 $Y2=5.1
r89 11 13 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.315 $Y=5.265
+ $X2=1.315 $Y2=5.925
r90 7 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=5.265
+ $X2=0.955 $Y2=5.1
r91 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.955 $Y=5.265
+ $X2=0.955 $Y2=5.925
r92 2 21 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.18
+ $Y=5.425 $X2=2.32 $Y2=5.55
r93 1 28 182 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_NDIFF $count=1 $X=2.18
+ $Y=3.59 $X2=2.32 $Y2=4.235
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A 3 5 7 10 12 13 16 21 22 24 27 31 34
+ 43 51
c72 27 0 3.44129e-20 $X=1.16 $Y=2.775
r73 42 43 61.0986 $w=3.4e-07 $l=3.6e-07 $layer=POLY_cond $X=0.955 $Y=1.96
+ $X2=1.315 $Y2=1.96
r74 39 42 34.7923 $w=3.4e-07 $l=2.05e-07 $layer=POLY_cond $X=0.75 $Y=1.96
+ $X2=0.955 $Y2=1.96
r75 34 51 8.5999 $w=6.03e-07 $l=4.35e-07 $layer=LI1_cond $X=0.725 $Y=1.832
+ $X2=1.16 $Y2=1.832
r76 34 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.955 $X2=0.75 $Y2=1.955
r77 32 46 22.0523 $w=3.06e-07 $l=1.4e-07 $layer=POLY_cond $X=1.405 $Y=2.925
+ $X2=1.405 $Y2=3.065
r78 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.405
+ $Y=2.925 $X2=1.405 $Y2=2.925
r79 28 31 9.41162 $w=2.98e-07 $l=2.45e-07 $layer=LI1_cond $X=1.16 $Y=2.925
+ $X2=1.405 $Y2=2.925
r80 27 28 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.16 $Y=2.775 $X2=1.16
+ $Y2=2.925
r81 26 51 8.37032 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=1.16 $Y=2.135
+ $X2=1.16 $Y2=1.832
r82 26 27 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.16 $Y=2.135
+ $X2=1.16 $Y2=2.775
r83 22 46 24.3585 $w=3.06e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.315 $Y=3.14
+ $X2=1.405 $Y2=3.065
r84 22 24 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.315 $Y=3.14
+ $X2=1.315 $Y2=4.01
r85 19 32 38.535 $w=3.06e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.315 $Y=2.76
+ $X2=1.405 $Y2=2.925
r86 19 21 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.315 $Y=2.76
+ $X2=1.315 $Y2=2.44
r87 18 43 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.315 $Y=2.13
+ $X2=1.315 $Y2=1.96
r88 18 21 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.315 $Y=2.13
+ $X2=1.315 $Y2=2.44
r89 14 43 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.315 $Y=1.79
+ $X2=1.315 $Y2=1.96
r90 14 16 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=1.315 $Y=1.79
+ $X2=1.315 $Y2=0.735
r91 12 46 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.24 $Y=3.065
+ $X2=1.405 $Y2=3.065
r92 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.24 $Y=3.065
+ $X2=1.03 $Y2=3.065
r93 8 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.955 $Y=3.14
+ $X2=1.03 $Y2=3.065
r94 8 10 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=0.955 $Y=3.14
+ $X2=0.955 $Y2=4.01
r95 5 42 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.955 $Y=2.13
+ $X2=0.955 $Y2=1.96
r96 5 7 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.955 $Y=2.13
+ $X2=0.955 $Y2=2.44
r97 1 42 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.955 $Y=1.79
+ $X2=0.955 $Y2=1.96
r98 1 3 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=0.955 $Y=1.79
+ $X2=0.955 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_278_47# 1 2 7 9 10 11 13 14 16 17 20
+ 26 28 29 31 33
c71 29 0 3.44129e-20 $X=1.98 $Y=2.925
r72 31 33 41.2959 $w=2.98e-07 $l=1.075e-06 $layer=LI1_cond $X=1.565 $Y=1.36
+ $X2=1.565 $Y2=2.435
r73 29 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=2.925
+ $X2=1.98 $Y2=3.09
r74 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.98
+ $Y=2.925 $X2=1.98 $Y2=2.925
r75 26 33 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.98 $Y=2.52
+ $X2=1.53 $Y2=2.52
r76 26 28 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.98 $Y=2.605
+ $X2=1.98 $Y2=2.925
r77 20 23 23.3781 $w=3.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.54 $Y=0.38
+ $X2=1.54 $Y2=1.09
r78 18 31 6.02978 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=1.54 $Y=1.185
+ $X2=1.54 $Y2=1.36
r79 18 23 3.12806 $w=3.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.54 $Y=1.185
+ $X2=1.54 $Y2=1.09
r80 14 17 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=2.105 $Y=3.515
+ $X2=2.087 $Y2=3.44
r81 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.105 $Y=3.515
+ $X2=2.105 $Y2=4.01
r82 13 17 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=2.07 $Y=3.365
+ $X2=2.087 $Y2=3.44
r83 13 39 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=2.07 $Y=3.365
+ $X2=2.07 $Y2=3.09
r84 10 17 5.30422 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=1.995 $Y=3.44
+ $X2=2.087 $Y2=3.44
r85 10 11 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.995 $Y=3.44
+ $X2=1.82 $Y2=3.44
r86 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.745 $Y=3.515
+ $X2=1.82 $Y2=3.44
r87 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.745 $Y=3.515
+ $X2=1.745 $Y2=4.01
r88 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.39
+ $Y=0.235 $X2=1.53 $Y2=1.09
r89 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.39
+ $Y=0.235 $X2=1.53 $Y2=0.38
r90 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.39
+ $Y=2.23 $X2=1.53 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_123_718# 1 2 7 9 10 12 13 14 17 21
+ 25 29 35 37 40 41 42 44 45 46 48 49 51 54 56 57 61 66 77
c157 77 0 6.8949e-20 $X=5.765 $Y=4.825
c158 49 0 6.60929e-20 $X=4.87 $Y=4.825
c159 14 0 1.8723e-19 $X=2.18 $Y=5.275
c160 7 0 1.70849e-20 $X=1.745 $Y=5.35
r161 66 72 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.58 $Y=5.1
+ $X2=2.58 $Y2=5.275
r162 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=5.1 $X2=2.58 $Y2=5.1
r163 62 67 3.32414 $w=2.9e-07 $l=2e-08 $layer=POLY_cond $X=1.765 $Y=5.142
+ $X2=1.745 $Y2=5.142
r164 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=5.1 $X2=1.765 $Y2=5.1
r165 56 57 5.31505 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.75 $Y=5.57
+ $X2=0.75 $Y2=5.435
r166 52 77 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.495 $Y=4.825
+ $X2=5.765 $Y2=4.825
r167 52 74 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.495 $Y=4.825
+ $X2=5.405 $Y2=4.825
r168 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.495
+ $Y=4.825 $X2=5.495 $Y2=4.825
r169 49 51 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=4.87 $Y=4.825
+ $X2=5.495 $Y2=4.825
r170 47 49 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.785 $Y=4.99
+ $X2=4.87 $Y2=4.825
r171 47 48 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=4.785 $Y=4.99
+ $X2=4.785 $Y2=6.235
r172 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.7 $Y=6.32
+ $X2=4.785 $Y2=6.235
r173 45 46 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.7 $Y=6.32
+ $X2=4.16 $Y2=6.32
r174 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.075 $Y=6.235
+ $X2=4.16 $Y2=6.32
r175 43 44 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=4.075 $Y=5.25
+ $X2=4.075 $Y2=6.235
r176 42 65 8.96033 $w=3.13e-07 $l=1.88348e-07 $layer=LI1_cond $X=2.745 $Y=5.165
+ $X2=2.58 $Y2=5.115
r177 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.99 $Y=5.165
+ $X2=4.075 $Y2=5.25
r178 41 42 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=3.99 $Y=5.165
+ $X2=2.745 $Y2=5.165
r179 40 61 10.1403 $w=1.73e-07 $l=1.6e-07 $layer=LI1_cond $X=1.605 $Y=5.097
+ $X2=1.765 $Y2=5.097
r180 39 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.605 $Y=4.82
+ $X2=1.605 $Y2=5.01
r181 38 54 3.01551 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.855 $Y=4.735
+ $X2=0.715 $Y2=4.735
r182 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.52 $Y=4.735
+ $X2=1.605 $Y2=4.82
r183 37 38 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.52 $Y=4.735
+ $X2=0.855 $Y2=4.735
r184 33 56 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.75 $Y=5.61 $X2=0.75
+ $Y2=5.57
r185 33 35 22.0611 $w=3.48e-07 $l=6.7e-07 $layer=LI1_cond $X=0.75 $Y=5.61
+ $X2=0.75 $Y2=6.28
r186 31 54 3.49088 $w=2.67e-07 $l=9.12688e-08 $layer=LI1_cond $X=0.702 $Y=4.82
+ $X2=0.715 $Y2=4.735
r187 31 57 27.7942 $w=2.53e-07 $l=6.15e-07 $layer=LI1_cond $X=0.702 $Y=4.82
+ $X2=0.702 $Y2=5.435
r188 27 54 3.49088 $w=2.67e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=4.65
+ $X2=0.715 $Y2=4.735
r189 27 29 37.0428 $w=2.78e-07 $l=9e-07 $layer=LI1_cond $X=0.715 $Y=4.65
+ $X2=0.715 $Y2=3.75
r190 23 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.765 $Y=4.99
+ $X2=5.765 $Y2=4.825
r191 23 25 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=5.765 $Y=4.99
+ $X2=5.765 $Y2=5.925
r192 19 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.765 $Y=4.66
+ $X2=5.765 $Y2=4.825
r193 19 21 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=5.765 $Y=4.66
+ $X2=5.765 $Y2=4.01
r194 15 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.405 $Y=4.66
+ $X2=5.405 $Y2=4.825
r195 15 17 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=5.405 $Y=4.66
+ $X2=5.405 $Y2=4.01
r196 13 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=5.275
+ $X2=2.58 $Y2=5.275
r197 13 14 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=2.415 $Y=5.275
+ $X2=2.18 $Y2=5.275
r198 10 14 23.6571 $w=2.9e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.105 $Y=5.35
+ $X2=2.18 $Y2=5.275
r199 10 62 56.5103 $w=2.9e-07 $l=4.31648e-07 $layer=POLY_cond $X=2.105 $Y=5.35
+ $X2=1.765 $Y2=5.142
r200 10 12 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.105 $Y=5.35
+ $X2=2.105 $Y2=5.925
r201 7 67 18.1727 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=1.745 $Y=5.35
+ $X2=1.745 $Y2=5.142
r202 7 9 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.745 $Y=5.35
+ $X2=1.745 $Y2=5.925
r203 2 56 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=5.425 $X2=0.74 $Y2=5.57
r204 2 35 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=5.425 $X2=0.74 $Y2=6.28
r205 1 29 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=0.615
+ $Y=3.59 $X2=0.74 $Y2=3.75
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_517_420# 1 2 7 9 10 11 14 15 16 17
+ 20 24 28
c74 14 0 2.24484e-20 $X=3.702 $Y=4.24
r75 24 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=3.75
+ $X2=3.995 $Y2=3.585
r76 23 26 10.7413 $w=4.6e-07 $l=4.05e-07 $layer=LI1_cond $X=3.785 $Y=3.75
+ $X2=3.785 $Y2=4.155
r77 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.995
+ $Y=3.75 $X2=3.995 $Y2=3.75
r78 18 20 35.4909 $w=1.98e-07 $l=6.4e-07 $layer=LI1_cond $X=4.43 $Y=4.91
+ $X2=4.43 $Y2=5.55
r79 16 18 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.33 $Y=4.825
+ $X2=4.43 $Y2=4.91
r80 16 17 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.33 $Y=4.825
+ $X2=3.815 $Y2=4.825
r81 15 17 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=3.702 $Y=4.74
+ $X2=3.815 $Y2=4.825
r82 14 26 5.44365 $w=4.6e-07 $l=1.19499e-07 $layer=LI1_cond $X=3.702 $Y=4.24
+ $X2=3.785 $Y2=4.155
r83 14 15 25.6098 $w=2.23e-07 $l=5e-07 $layer=LI1_cond $X=3.702 $Y=4.24
+ $X2=3.702 $Y2=4.74
r84 12 28 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.905 $Y=3.295
+ $X2=3.905 $Y2=3.585
r85 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.83 $Y=3.22
+ $X2=3.905 $Y2=3.295
r86 10 11 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=3.83 $Y=3.22
+ $X2=2.735 $Y2=3.22
r87 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.66 $Y=3.145
+ $X2=2.735 $Y2=3.22
r88 7 9 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.66 $Y=3.145 $X2=2.66
+ $Y2=2.65
r89 2 20 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=4.305
+ $Y=5.425 $X2=4.445 $Y2=5.55
r90 1 26 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=4.01 $X2=3.655 $Y2=4.155
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%SLEEP 1 3 4 6 9 11 15 17 20 21 23 24
+ 26 28 30 31 33 35 36 38 39 40 41 42 43 49 51
c115 28 0 2.24484e-20 $X=4.615 $Y=4.505
c116 1 0 1.58517e-19 $X=3.08 $Y=4.505
r117 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.255
+ $Y=4.705 $X2=3.255 $Y2=4.705
r118 43 49 3.84148 $w=4.03e-07 $l=1.35e-07 $layer=LI1_cond $X=3.12 $Y=4.707
+ $X2=3.255 $Y2=4.707
r119 36 38 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.405 $Y=5.35
+ $X2=5.405 $Y2=5.925
r120 33 35 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.975 $Y=4.505
+ $X2=4.975 $Y2=4.01
r121 32 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.69 $Y=4.58
+ $X2=4.615 $Y2=4.58
r122 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.9 $Y=4.58
+ $X2=4.975 $Y2=4.505
r123 31 32 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.9 $Y=4.58
+ $X2=4.69 $Y2=4.58
r124 28 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.615 $Y=4.505
+ $X2=4.615 $Y2=4.58
r125 28 30 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.615 $Y=4.505
+ $X2=4.615 $Y2=4.01
r126 27 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.305 $Y=5.275
+ $X2=4.23 $Y2=5.275
r127 26 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.33 $Y=5.275
+ $X2=5.405 $Y2=5.35
r128 26 27 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=5.33 $Y=5.275
+ $X2=4.305 $Y2=5.275
r129 25 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.305 $Y=4.58
+ $X2=4.23 $Y2=4.58
r130 24 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.54 $Y=4.58
+ $X2=4.615 $Y2=4.58
r131 24 25 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=4.54 $Y=4.58
+ $X2=4.305 $Y2=4.58
r132 21 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.23 $Y=5.35
+ $X2=4.23 $Y2=5.275
r133 21 23 184.767 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=4.23 $Y=5.35
+ $X2=4.23 $Y2=5.925
r134 20 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.23 $Y=5.2
+ $X2=4.23 $Y2=5.275
r135 19 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.23 $Y=4.655
+ $X2=4.23 $Y2=4.58
r136 19 20 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.23 $Y=4.655
+ $X2=4.23 $Y2=5.2
r137 18 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.945 $Y=4.58
+ $X2=3.87 $Y2=4.58
r138 17 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.155 $Y=4.58
+ $X2=4.23 $Y2=4.58
r139 17 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.155 $Y=4.58
+ $X2=3.945 $Y2=4.58
r140 13 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.87 $Y=4.655
+ $X2=3.87 $Y2=4.58
r141 13 15 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=3.87 $Y=4.655
+ $X2=3.87 $Y2=5.925
r142 11 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.795 $Y=4.58
+ $X2=3.87 $Y2=4.58
r143 11 51 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.795 $Y=4.58
+ $X2=3.515 $Y2=4.58
r144 7 9 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=3.44 $Y=4.87
+ $X2=3.44 $Y2=5.925
r145 4 51 32.4387 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=3.44 $Y=4.687
+ $X2=3.515 $Y2=4.687
r146 4 7 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.44 $Y=4.687
+ $X2=3.44 $Y2=4.87
r147 4 48 29.2473 $w=3.65e-07 $l=1.85e-07 $layer=POLY_cond $X=3.44 $Y=4.687
+ $X2=3.255 $Y2=4.687
r148 4 6 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.44 $Y=4.505 $X2=3.44
+ $Y2=4.22
r149 1 48 27.6664 $w=3.65e-07 $l=1.75e-07 $layer=POLY_cond $X=3.08 $Y=4.687
+ $X2=3.255 $Y2=4.687
r150 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.08 $Y=4.505 $X2=3.08
+ $Y2=4.22
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%VPWR 1 6 10 12 22 23 26
r24 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r25 22 23 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r26 20 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r27 19 22 344.471 $w=1.68e-07 $l=5.28e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=6.48
+ $Y2=0
r28 19 20 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r29 17 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.74
+ $Y2=0
r30 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.2
+ $Y2=0
r31 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r32 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 12 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.74
+ $Y2=0
r34 12 14 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.24
+ $Y2=0
r35 10 23 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=6.48
+ $Y2=0
r36 10 20 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=1.2
+ $Y2=0
r37 6 8 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.74 $Y=0.38 $X2=0.74
+ $Y2=1.09
r38 4 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0
r39 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.38
r40 1 8 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.74 $Y2=1.09
r41 1 6 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.74 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_278_1085# 1 2 9 11 12 13 15
r33 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=6.235
+ $X2=3.225 $Y2=6.32
r34 13 15 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.225 $Y=6.235
+ $X2=3.225 $Y2=5.6
r35 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=6.32
+ $X2=3.225 $Y2=6.32
r36 11 12 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=3.06 $Y=6.32
+ $X2=1.695 $Y2=6.32
r37 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.53 $Y=6.235
+ $X2=1.695 $Y2=6.32
r38 7 9 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.53 $Y=6.235
+ $X2=1.53 $Y2=5.78
r39 2 18 400 $w=1.7e-07 $l=9.17701e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=5.425 $X2=3.225 $Y2=6.28
r40 2 15 400 $w=1.7e-07 $l=2.3103e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=5.425 $X2=3.225 $Y2=5.6
r41 1 9 300 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=2 $X=1.39
+ $Y=5.425 $X2=1.53 $Y2=5.78
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%DESTPWR 1 2 9 15 19 21 26 36 37 40 43
c66 15 0 6.8949e-20 $X=5.19 $Y=5.585
r67 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=6.66
+ $X2=5.04 $Y2=6.66
r68 40 41 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=6.66
+ $X2=3.6 $Y2=6.66
r69 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=6.66
+ $X2=6.48 $Y2=6.66
r70 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=6.66
+ $X2=6.48 $Y2=6.66
r71 34 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=6.66
+ $X2=5.04 $Y2=6.66
r72 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=6.66 $X2=6.48
+ $Y2=6.66
r73 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=6.66
+ $X2=5.52 $Y2=6.66
r74 31 43 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=5.355 $Y=6.66
+ $X2=5.197 $Y2=6.66
r75 31 33 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=6.66
+ $X2=5.52 $Y2=6.66
r76 30 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=6.66
+ $X2=5.04 $Y2=6.66
r77 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=6.66
+ $X2=3.6 $Y2=6.66
r78 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=6.66
+ $X2=4.08 $Y2=6.66
r79 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=6.66
+ $X2=3.655 $Y2=6.66
r80 27 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.74 $Y=6.66
+ $X2=4.08 $Y2=6.66
r81 26 43 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=5.04 $Y=6.66
+ $X2=5.197 $Y2=6.66
r82 26 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=6.66 $X2=4.08
+ $Y2=6.66
r83 23 24 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=6.66
+ $X2=0.24 $Y2=6.66
r84 21 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=6.66
+ $X2=3.655 $Y2=6.66
r85 21 23 217.251 $w=1.68e-07 $l=3.33e-06 $layer=LI1_cond $X=3.57 $Y=6.66
+ $X2=0.24 $Y2=6.66
r86 19 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=6.66
+ $X2=3.6 $Y2=6.66
r87 19 24 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=3.36 $Y=6.66
+ $X2=0.24 $Y2=6.66
r88 15 18 26.1586 $w=3.13e-07 $l=7.15e-07 $layer=LI1_cond $X=5.197 $Y=5.585
+ $X2=5.197 $Y2=6.3
r89 13 43 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.197 $Y=6.575
+ $X2=5.197 $Y2=6.66
r90 13 18 10.061 $w=3.13e-07 $l=2.75e-07 $layer=LI1_cond $X=5.197 $Y=6.575
+ $X2=5.197 $Y2=6.3
r91 9 12 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.655 $Y=5.585
+ $X2=3.655 $Y2=6.3
r92 7 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=6.575
+ $X2=3.655 $Y2=6.66
r93 7 12 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.655 $Y=6.575
+ $X2=3.655 $Y2=6.3
r94 2 18 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=5.045
+ $Y=5.425 $X2=5.19 $Y2=6.3
r95 2 15 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=5.045
+ $Y=5.425 $X2=5.19 $Y2=5.585
r96 1 12 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=5.425 $X2=3.655 $Y2=6.3
r97 1 9 400 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=5.425 $X2=3.655 $Y2=5.585
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%X 1 2 3 12 14 15 16 17 18 19 20 21 31
+ 37
r48 29 37 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=5.98 $Y=4.32
+ $X2=5.98 $Y2=4.255
r49 21 50 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=5.98 $Y=5.735
+ $X2=5.98 $Y2=6.28
r50 21 46 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.98 $Y=5.735
+ $X2=5.98 $Y2=5.57
r51 20 46 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.98 $Y=5.365
+ $X2=5.98 $Y2=5.57
r52 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.98 $Y=4.995
+ $X2=5.98 $Y2=5.365
r53 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.98 $Y=4.625
+ $X2=5.98 $Y2=4.995
r54 18 38 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.98 $Y=4.625
+ $X2=5.98 $Y2=4.49
r55 17 29 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=4.405
+ $X2=5.98 $Y2=4.32
r56 17 38 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.98 $Y=4.405
+ $X2=5.98 $Y2=4.49
r57 17 37 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=5.98 $Y=4.245
+ $X2=5.98 $Y2=4.255
r58 16 17 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.98 $Y=3.885
+ $X2=5.98 $Y2=4.245
r59 16 31 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.98 $Y=3.885
+ $X2=5.98 $Y2=3.735
r60 14 17 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=4.405
+ $X2=5.98 $Y2=4.405
r61 14 15 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=5.815 $Y=4.405
+ $X2=4.565 $Y2=4.405
r62 10 15 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.425 $Y=4.32
+ $X2=4.565 $Y2=4.405
r63 10 12 23.2547 $w=2.78e-07 $l=5.65e-07 $layer=LI1_cond $X=4.425 $Y=4.32
+ $X2=4.425 $Y2=3.755
r64 3 50 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=5.84
+ $Y=5.425 $X2=5.98 $Y2=6.28
r65 3 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.84
+ $Y=5.425 $X2=5.98 $Y2=5.57
r66 2 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.84
+ $Y=3.59 $X2=5.98 $Y2=3.735
r67 1 12 91 $w=1.7e-07 $l=2.20624e-07 $layer=licon1_NDIFF $count=2 $X=4.27
+ $Y=3.59 $X2=4.4 $Y2=3.755
.ends

.subckt PM_SKY130_FD_SC_LP__LSBUFISO0P_LP%A_278_718# 1 2 9 13 16 18 19
c38 18 0 1.8723e-19 $X=1.53 $Y=3.75
r39 16 19 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.4 $Y=3.585
+ $X2=2.4 $Y2=3.09
r40 11 19 6.27261 $w=2.13e-07 $l=1.07e-07 $layer=LI1_cond $X=2.422 $Y=2.983
+ $X2=2.422 $Y2=3.09
r41 11 13 26.1578 $w=2.13e-07 $l=4.88e-07 $layer=LI1_cond $X=2.422 $Y=2.983
+ $X2=2.422 $Y2=2.495
r42 10 18 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.645 $Y=3.67
+ $X2=1.505 $Y2=3.67
r43 9 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.315 $Y=3.67
+ $X2=2.4 $Y2=3.585
r44 9 10 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.315 $Y=3.67
+ $X2=1.645 $Y2=3.67
r45 2 13 91 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=2 $X=2.32
+ $Y=2.23 $X2=2.445 $Y2=2.495
r46 1 18 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=1.39
+ $Y=3.59 $X2=1.53 $Y2=3.75
.ends

