* File: sky130_fd_sc_lp__and3_1.pex.spice
* Created: Fri Aug 28 10:05:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3_1%A 3 7 9 12
r29 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.27
+ $X2=0.58 $Y2=1.435
r30 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.27
+ $X2=0.58 $Y2=1.105
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.58
+ $Y=1.27 $X2=0.58 $Y2=1.27
r32 9 13 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.72 $Y=1.27 $X2=0.58
+ $Y2=1.27
r33 7 14 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.67 $Y=0.475
+ $X2=0.67 $Y2=1.105
r34 3 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.645 $Y=2.045
+ $X2=0.645 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_1%B 3 7 9 12
r31 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.27
+ $X2=1.15 $Y2=1.435
r32 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.27
+ $X2=1.15 $Y2=1.105
r33 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.27 $X2=1.15 $Y2=1.27
r34 7 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.095 $Y=2.045
+ $X2=1.095 $Y2=1.435
r35 3 14 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.06 $Y=0.475
+ $X2=1.06 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_1%C 3 7 9 10 11 12 13 22 26 41
c50 26 0 1.86775e-19 $X=1.685 $Y=1.52
r51 41 42 3.31806 $w=2.58e-07 $l=5e-08 $layer=LI1_cond $X=1.645 $Y=2.405
+ $X2=1.645 $Y2=2.355
r52 22 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.38
+ $X2=1.69 $Y2=1.545
r53 22 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.38
+ $X2=1.69 $Y2=1.215
r54 12 33 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=1.645 $Y=2.42
+ $X2=1.645 $Y2=2.485
r55 12 41 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.645 $Y=2.42
+ $X2=1.645 $Y2=2.405
r56 12 13 12.7655 $w=2.58e-07 $l=2.88e-07 $layer=LI1_cond $X=1.645 $Y=2.487
+ $X2=1.645 $Y2=2.775
r57 12 33 0.0886495 $w=2.58e-07 $l=2e-09 $layer=LI1_cond $X=1.645 $Y=2.487
+ $X2=1.645 $Y2=2.485
r58 12 42 1.10909 $w=1.78e-07 $l=1.8e-08 $layer=LI1_cond $X=1.685 $Y=2.337
+ $X2=1.685 $Y2=2.355
r59 11 12 18.6081 $w=1.78e-07 $l=3.02e-07 $layer=LI1_cond $X=1.685 $Y=2.035
+ $X2=1.685 $Y2=2.337
r60 10 11 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=2.035
r61 10 26 8.93434 $w=1.78e-07 $l=1.45e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=1.52
r62 9 26 11.859 $w=2.54e-07 $l=2.45561e-07 $layer=LI1_cond $X=1.642 $Y=1.295
+ $X2=1.685 $Y2=1.52
r63 9 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.38 $X2=1.69 $Y2=1.38
r64 7 25 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.6 $Y=2.045 $X2=1.6
+ $Y2=1.545
r65 3 24 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.6 $Y=0.475 $X2=1.6
+ $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_1%A_61_367# 1 2 3 12 16 19 22 24 26 30 33 35 39
+ 43 49
c83 49 0 1.86775e-19 $X=2.385 $Y=1.47
r84 44 49 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.23 $Y=1.47
+ $X2=2.385 $Y2=1.47
r85 44 46 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.23 $Y=1.47
+ $X2=2.195 $Y2=1.47
r86 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.47 $X2=2.23 $Y2=1.47
r87 40 43 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.035 $Y=1.47
+ $X2=2.23 $Y2=1.47
r88 37 38 7.35235 $w=4.73e-07 $l=8.5e-08 $layer=LI1_cond $X=0.382 $Y=0.85
+ $X2=0.382 $Y2=0.935
r89 35 37 9.44272 $w=4.73e-07 $l=3.75e-07 $layer=LI1_cond $X=0.382 $Y=0.475
+ $X2=0.382 $Y2=0.85
r90 33 40 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=1.305
+ $X2=2.035 $Y2=1.47
r91 32 33 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.035 $Y=0.935
+ $X2=2.035 $Y2=1.305
r92 28 30 12.965 $w=2.38e-07 $l=2.7e-07 $layer=LI1_cond $X=1.305 $Y=1.775
+ $X2=1.305 $Y2=2.045
r93 27 37 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.62 $Y=0.85
+ $X2=0.382 $Y2=0.85
r94 26 32 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.945 $Y=0.85
+ $X2=2.035 $Y2=0.935
r95 26 27 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=1.945 $Y=0.85
+ $X2=0.62 $Y2=0.85
r96 25 39 3.3845 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.565 $Y=1.69
+ $X2=0.355 $Y2=1.69
r97 24 28 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.185 $Y=1.69
+ $X2=1.305 $Y2=1.775
r98 24 25 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.185 $Y=1.69
+ $X2=0.565 $Y2=1.69
r99 20 39 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.355 $Y=1.775
+ $X2=0.355 $Y2=1.69
r100 20 22 7.40856 $w=4.18e-07 $l=2.7e-07 $layer=LI1_cond $X=0.355 $Y=1.775
+ $X2=0.355 $Y2=2.045
r101 19 39 3.19717 $w=2.95e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.23 $Y=1.605
+ $X2=0.355 $Y2=1.69
r102 19 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.23 $Y=1.605
+ $X2=0.23 $Y2=0.935
r103 14 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.635
+ $X2=2.385 $Y2=1.47
r104 14 16 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.385 $Y=1.635
+ $X2=2.385 $Y2=2.465
r105 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.305
+ $X2=2.195 $Y2=1.47
r106 10 12 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.195 $Y=1.305
+ $X2=2.195 $Y2=0.685
r107 3 30 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=1.17
+ $Y=1.835 $X2=1.33 $Y2=2.045
r108 2 22 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.835 $X2=0.43 $Y2=2.045
r109 1 35 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.33
+ $Y=0.265 $X2=0.455 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_1%VPWR 1 2 9 13 18 19 20 26 32 33 36
r28 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 33 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 30 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.135 $Y2=3.33
r32 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 26 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=2.135 $Y2=3.33
r36 26 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 20 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 20 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 18 23 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 18 19 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.875 $Y2=3.33
r42 17 28 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 17 19 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.875 $Y2=3.33
r44 13 16 13.799 $w=3.78e-07 $l=4.55e-07 $layer=LI1_cond $X=2.135 $Y=1.975
+ $X2=2.135 $Y2=2.43
r45 11 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=3.33
r46 11 16 24.7169 $w=3.78e-07 $l=8.15e-07 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=2.43
r47 7 19 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=3.33
r48 7 9 46.7151 $w=2.78e-07 $l=1.135e-06 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=2.11
r49 2 16 300 $w=1.7e-07 $l=8.05326e-07 $layer=licon1_PDIFF $count=2 $X=1.675
+ $Y=1.835 $X2=2.17 $Y2=2.43
r50 2 13 600 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.675
+ $Y=1.835 $X2=2.03 $Y2=1.975
r51 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.835 $X2=0.86 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_1%X 1 2 7 8 9 10 11 12 13 24 45
r19 22 45 1.19608 $w=4.98e-07 $l=5e-08 $layer=LI1_cond $X=2.545 $Y=0.875
+ $X2=2.545 $Y2=0.925
r20 13 42 5.18599 $w=2.98e-07 $l=1.35e-07 $layer=LI1_cond $X=2.645 $Y=2.775
+ $X2=2.645 $Y2=2.91
r21 12 13 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=2.405
+ $X2=2.645 $Y2=2.775
r22 11 12 16.3263 $w=2.98e-07 $l=4.25e-07 $layer=LI1_cond $X=2.645 $Y=1.98
+ $X2=2.645 $Y2=2.405
r23 10 11 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=2.645 $Y=1.665
+ $X2=2.645 $Y2=1.98
r24 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=1.295
+ $X2=2.645 $Y2=1.665
r25 9 47 6.53051 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=2.645 $Y=1.295
+ $X2=2.645 $Y2=1.125
r26 8 47 6.27653 $w=4.98e-07 $l=1.83e-07 $layer=LI1_cond $X=2.545 $Y=0.942
+ $X2=2.545 $Y2=1.125
r27 8 45 0.406667 $w=4.98e-07 $l=1.7e-08 $layer=LI1_cond $X=2.545 $Y=0.942
+ $X2=2.545 $Y2=0.925
r28 8 22 0.430588 $w=4.98e-07 $l=1.8e-08 $layer=LI1_cond $X=2.545 $Y=0.857
+ $X2=2.545 $Y2=0.875
r29 7 8 7.22431 $w=4.98e-07 $l=3.02e-07 $layer=LI1_cond $X=2.545 $Y=0.555
+ $X2=2.545 $Y2=0.857
r30 7 24 3.22941 $w=4.98e-07 $l=1.35e-07 $layer=LI1_cond $X=2.545 $Y=0.555
+ $X2=2.545 $Y2=0.42
r31 2 42 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.835 $X2=2.6 $Y2=2.91
r32 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.835 $X2=2.6 $Y2=1.98
r33 1 24 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.265 $X2=2.41 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_1%VGND 1 6 9 10 11 21 22
r24 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r25 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r26 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r27 14 18 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r28 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 11 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r30 11 15 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.24
+ $Y2=0
r31 9 18 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.68
+ $Y2=0
r32 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.905
+ $Y2=0
r33 8 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.64
+ $Y2=0
r34 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.905
+ $Y2=0
r35 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=0.085
+ $X2=1.905 $Y2=0
r36 4 6 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.905 $Y=0.085
+ $X2=1.905 $Y2=0.455
r37 1 6 182 $w=1.7e-07 $l=3.10805e-07 $layer=licon1_NDIFF $count=1 $X=1.675
+ $Y=0.265 $X2=1.905 $Y2=0.455
.ends

