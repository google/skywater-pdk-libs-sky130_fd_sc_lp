* File: sky130_fd_sc_lp__a221o_lp.pxi.spice
* Created: Wed Sep  2 09:21:29 2020
* 
x_PM_SKY130_FD_SC_LP__A221O_LP%A_96_183# N_A_96_183#_M1011_d N_A_96_183#_M1008_d
+ N_A_96_183#_M1002_d N_A_96_183#_M1003_g N_A_96_183#_M1010_g N_A_96_183#_c_94_n
+ N_A_96_183#_c_95_n N_A_96_183#_c_96_n N_A_96_183#_M1013_g N_A_96_183#_c_97_n
+ N_A_96_183#_c_98_n N_A_96_183#_c_99_n N_A_96_183#_c_100_n N_A_96_183#_c_113_n
+ N_A_96_183#_c_114_n N_A_96_183#_c_101_n N_A_96_183#_c_102_n
+ N_A_96_183#_c_103_n N_A_96_183#_c_104_n N_A_96_183#_c_105_n
+ N_A_96_183#_c_106_n N_A_96_183#_c_107_n N_A_96_183#_c_108_n
+ N_A_96_183#_c_109_n N_A_96_183#_c_116_n N_A_96_183#_c_110_n
+ PM_SKY130_FD_SC_LP__A221O_LP%A_96_183#
x_PM_SKY130_FD_SC_LP__A221O_LP%A2 N_A2_M1005_g N_A2_M1004_g A2 N_A2_c_228_n
+ N_A2_c_229_n PM_SKY130_FD_SC_LP__A221O_LP%A2
x_PM_SKY130_FD_SC_LP__A221O_LP%A1 N_A1_M1012_g N_A1_M1011_g N_A1_c_269_n A1 A1
+ A1 N_A1_c_271_n N_A1_c_272_n PM_SKY130_FD_SC_LP__A221O_LP%A1
x_PM_SKY130_FD_SC_LP__A221O_LP%B1 N_B1_c_313_n N_B1_c_318_n N_B1_c_319_n
+ N_B1_M1000_g N_B1_c_320_n N_B1_M1009_g B1 N_B1_c_316_n
+ PM_SKY130_FD_SC_LP__A221O_LP%B1
x_PM_SKY130_FD_SC_LP__A221O_LP%B2 N_B2_M1001_g N_B2_M1006_g B2 B2 N_B2_c_370_n
+ PM_SKY130_FD_SC_LP__A221O_LP%B2
x_PM_SKY130_FD_SC_LP__A221O_LP%C1 N_C1_c_411_n N_C1_M1007_g N_C1_c_412_n
+ N_C1_c_413_n N_C1_c_414_n N_C1_M1008_g N_C1_c_420_n N_C1_M1002_g N_C1_c_415_n
+ N_C1_c_416_n N_C1_c_417_n C1 C1 N_C1_c_419_n PM_SKY130_FD_SC_LP__A221O_LP%C1
x_PM_SKY130_FD_SC_LP__A221O_LP%X N_X_M1010_s N_X_M1003_s N_X_c_462_n X X X
+ N_X_c_463_n PM_SKY130_FD_SC_LP__A221O_LP%X
x_PM_SKY130_FD_SC_LP__A221O_LP%VPWR N_VPWR_M1003_d N_VPWR_M1012_d N_VPWR_c_489_n
+ N_VPWR_c_490_n N_VPWR_c_491_n VPWR N_VPWR_c_492_n N_VPWR_c_493_n
+ N_VPWR_c_488_n N_VPWR_c_495_n N_VPWR_c_496_n PM_SKY130_FD_SC_LP__A221O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A221O_LP%A_322_419# N_A_322_419#_M1005_d
+ N_A_322_419#_M1009_d N_A_322_419#_c_539_n N_A_322_419#_c_534_n
+ N_A_322_419#_c_535_n N_A_322_419#_c_548_n
+ PM_SKY130_FD_SC_LP__A221O_LP%A_322_419#
x_PM_SKY130_FD_SC_LP__A221O_LP%A_545_400# N_A_545_400#_M1009_s
+ N_A_545_400#_M1006_d N_A_545_400#_c_569_n N_A_545_400#_c_570_n
+ N_A_545_400#_c_571_n N_A_545_400#_c_573_n
+ PM_SKY130_FD_SC_LP__A221O_LP%A_545_400#
x_PM_SKY130_FD_SC_LP__A221O_LP%VGND N_VGND_M1013_d N_VGND_M1001_d N_VGND_c_601_n
+ N_VGND_c_602_n N_VGND_c_603_n N_VGND_c_604_n VGND N_VGND_c_605_n
+ N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n PM_SKY130_FD_SC_LP__A221O_LP%VGND
cc_1 VNB N_A_96_183#_M1003_g 0.00483251f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.595
cc_2 VNB N_A_96_183#_M1010_g 0.0158476f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.54
cc_3 VNB N_A_96_183#_c_94_n 0.0230144f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.18
cc_4 VNB N_A_96_183#_c_95_n 0.0127798f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.18
cc_5 VNB N_A_96_183#_c_96_n 0.0142047f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=0.255
cc_6 VNB N_A_96_183#_c_97_n 0.0287563f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.42
cc_7 VNB N_A_96_183#_c_98_n 0.0151341f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.585
cc_8 VNB N_A_96_183#_c_99_n 0.0310705f $X=-0.19 $Y=-0.245 $X2=1.58 $Y2=1
cc_9 VNB N_A_96_183#_c_100_n 0.00389079f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=1.71
cc_10 VNB N_A_96_183#_c_101_n 0.00357292f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=0.54
cc_11 VNB N_A_96_183#_c_102_n 0.00507726f $X=-0.19 $Y=-0.245 $X2=3.01 $Y2=0.905
cc_12 VNB N_A_96_183#_c_103_n 0.00537921f $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=0.905
cc_13 VNB N_A_96_183#_c_104_n 0.00819525f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=1.71
cc_14 VNB N_A_96_183#_c_105_n 0.00427551f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.08
cc_15 VNB N_A_96_183#_c_106_n 0.0195983f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.08
cc_16 VNB N_A_96_183#_c_107_n 0.00280775f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=0.905
cc_17 VNB N_A_96_183#_c_108_n 0.0177782f $X=-0.19 $Y=-0.245 $X2=4.155 $Y2=0.65
cc_18 VNB N_A_96_183#_c_109_n 0.0475189f $X=-0.19 $Y=-0.245 $X2=4.625 $Y2=0.65
cc_19 VNB N_A_96_183#_c_110_n 0.0324631f $X=-0.19 $Y=-0.245 $X2=4.502 $Y2=2.02
cc_20 VNB N_A2_M1004_g 0.0400805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_c_228_n 0.048675f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.595
cc_22 VNB N_A2_c_229_n 0.0028866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_269_n 0.0471502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB A1 0.00813512f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.585
cc_25 VNB N_A1_c_271_n 0.018028f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.54
cc_26 VNB N_A1_c_272_n 0.0191765f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.18
cc_27 VNB N_B1_c_313_n 0.00687175f $X=-0.19 $Y=-0.245 $X2=4.18 $Y2=0.33
cc_28 VNB N_B1_M1000_g 0.0362774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB B1 0.00424878f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.595
cc_30 VNB N_B1_c_316_n 0.0408453f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.18
cc_31 VNB N_B2_M1001_g 0.0385f $X=-0.19 $Y=-0.245 $X2=4.32 $Y2=2
cc_32 VNB N_B2_M1006_g 0.0079351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB B2 0.00462003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B2_c_370_n 0.0555704f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.18
cc_35 VNB N_C1_c_411_n 0.0152627f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=0.33
cc_36 VNB N_C1_c_412_n 0.0101095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_C1_c_413_n 0.0071232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_C1_c_414_n 0.0182912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_C1_c_415_n 0.00667205f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.915
cc_40 VNB N_C1_c_416_n 0.0168513f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.54
cc_41 VNB N_C1_c_417_n 0.0226263f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=0.18
cc_42 VNB C1 0.00564083f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.18
cc_43 VNB N_C1_c_419_n 0.0175765f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.915
cc_44 VNB N_X_c_462_n 0.0261186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_463_n 0.0439454f $X=-0.19 $Y=-0.245 $X2=3.01 $Y2=1.795
cc_46 VNB N_VPWR_c_488_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1
cc_47 VNB N_VGND_c_601_n 0.00544226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_602_n 0.00545551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_603_n 0.0371607f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.54
cc_50 VNB N_VGND_c_604_n 0.00585462f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.54
cc_51 VNB N_VGND_c_605_n 0.048811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_606_n 0.0354908f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=0.54
cc_53 VNB N_VGND_c_607_n 0.287566f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=0.54
cc_54 VNB N_VGND_c_608_n 0.00585462f $X=-0.19 $Y=-0.245 $X2=2.785 $Y2=0.905
cc_55 VPB N_A_96_183#_M1003_g 0.0521972f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.595
cc_56 VPB N_A_96_183#_c_100_n 5.08562e-19 $X=-0.19 $Y=1.655 $X2=1.665 $Y2=1.71
cc_57 VPB N_A_96_183#_c_113_n 0.0284849f $X=-0.19 $Y=1.655 $X2=3.01 $Y2=1.795
cc_58 VPB N_A_96_183#_c_114_n 6.5944e-19 $X=-0.19 $Y=1.655 $X2=1.75 $Y2=1.795
cc_59 VPB N_A_96_183#_c_104_n 9.89493e-19 $X=-0.19 $Y=1.655 $X2=3.095 $Y2=1.71
cc_60 VPB N_A_96_183#_c_116_n 0.0453272f $X=-0.19 $Y=1.655 $X2=4.46 $Y2=2.185
cc_61 VPB N_A_96_183#_c_110_n 0.0174507f $X=-0.19 $Y=1.655 $X2=4.502 $Y2=2.02
cc_62 VPB N_A2_M1005_g 0.0281814f $X=-0.19 $Y=1.655 $X2=4.32 $Y2=2
cc_63 VPB N_A2_c_228_n 0.0367346f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.595
cc_64 VPB N_A2_c_229_n 0.00325889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A1_M1012_g 0.0423063f $X=-0.19 $Y=1.655 $X2=4.32 $Y2=2
cc_66 VPB N_B1_c_313_n 0.0795019f $X=-0.19 $Y=1.655 $X2=4.18 $Y2=0.33
cc_67 VPB N_B1_c_318_n 0.0381808f $X=-0.19 $Y=1.655 $X2=4.32 $Y2=2
cc_68 VPB N_B1_c_319_n 0.0100618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_B1_c_320_n 0.0198882f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_B2_M1006_g 0.0397126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB B2 0.0029824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_C1_c_420_n 0.013958f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.595
cc_73 VPB N_C1_M1002_g 0.0302692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_C1_c_417_n 0.00134765f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=0.18
cc_75 VPB C1 0.00287287f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.18
cc_76 VPB X 0.0289805f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.595
cc_77 VPB X 0.0377443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_X_c_463_n 0.0132448f $X=-0.19 $Y=1.655 $X2=3.01 $Y2=1.795
cc_79 VPB N_VPWR_c_489_n 0.00562917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_490_n 0.0203665f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.595
cc_81 VPB N_VPWR_c_491_n 0.00823696f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=0.915
cc_82 VPB N_VPWR_c_492_n 0.0279108f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.18
cc_83 VPB N_VPWR_c_493_n 0.0607843f $X=-0.19 $Y=1.655 $X2=1.58 $Y2=1
cc_84 VPB N_VPWR_c_488_n 0.0557165f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1
cc_85 VPB N_VPWR_c_495_n 0.00632158f $X=-0.19 $Y=1.655 $X2=3.01 $Y2=1.795
cc_86 VPB N_VPWR_c_496_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.62 $Y2=0.54
cc_87 VPB N_A_322_419#_c_534_n 0.00789863f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.595
cc_88 VPB N_A_322_419#_c_535_n 0.0024287f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.595
cc_89 VPB N_A_545_400#_c_569_n 0.00377584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_545_400#_c_570_n 0.00410318f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.595
cc_91 VPB N_A_545_400#_c_571_n 0.00344132f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.595
cc_92 N_A_96_183#_M1003_g N_A2_M1005_g 0.0155724f $X=0.685 $Y=2.595 $X2=0 $Y2=0
cc_93 N_A_96_183#_M1010_g N_A2_M1004_g 0.00629906f $X=0.735 $Y=0.54 $X2=0 $Y2=0
cc_94 N_A_96_183#_c_94_n N_A2_M1004_g 0.0150947f $X=1.02 $Y=0.18 $X2=0 $Y2=0
cc_95 N_A_96_183#_c_99_n N_A2_M1004_g 0.0154078f $X=1.58 $Y=1 $X2=0 $Y2=0
cc_96 N_A_96_183#_c_100_n N_A2_M1004_g 0.00901782f $X=1.665 $Y=1.71 $X2=0 $Y2=0
cc_97 N_A_96_183#_c_96_n N_A2_c_228_n 0.00287028f $X=1.095 $Y=0.255 $X2=0 $Y2=0
cc_98 N_A_96_183#_c_97_n N_A2_c_228_n 0.0352391f $X=0.645 $Y=1.42 $X2=0 $Y2=0
cc_99 N_A_96_183#_c_99_n N_A2_c_228_n 0.00729592f $X=1.58 $Y=1 $X2=0 $Y2=0
cc_100 N_A_96_183#_c_100_n N_A2_c_228_n 0.0121273f $X=1.665 $Y=1.71 $X2=0 $Y2=0
cc_101 N_A_96_183#_c_114_n N_A2_c_228_n 0.00653797f $X=1.75 $Y=1.795 $X2=0 $Y2=0
cc_102 N_A_96_183#_c_105_n N_A2_c_228_n 0.00136441f $X=0.645 $Y=1.08 $X2=0 $Y2=0
cc_103 N_A_96_183#_c_97_n N_A2_c_229_n 0.00345003f $X=0.645 $Y=1.42 $X2=0 $Y2=0
cc_104 N_A_96_183#_c_99_n N_A2_c_229_n 0.0250673f $X=1.58 $Y=1 $X2=0 $Y2=0
cc_105 N_A_96_183#_c_100_n N_A2_c_229_n 0.0303225f $X=1.665 $Y=1.71 $X2=0 $Y2=0
cc_106 N_A_96_183#_c_114_n N_A2_c_229_n 0.0129587f $X=1.75 $Y=1.795 $X2=0 $Y2=0
cc_107 N_A_96_183#_c_105_n N_A2_c_229_n 0.0170751f $X=0.645 $Y=1.08 $X2=0 $Y2=0
cc_108 N_A_96_183#_c_113_n N_A1_M1012_g 0.0159895f $X=3.01 $Y=1.795 $X2=0 $Y2=0
cc_109 N_A_96_183#_c_100_n N_A1_c_269_n 0.00633766f $X=1.665 $Y=1.71 $X2=0 $Y2=0
cc_110 N_A_96_183#_c_113_n N_A1_c_269_n 8.25547e-19 $X=3.01 $Y=1.795 $X2=0 $Y2=0
cc_111 N_A_96_183#_M1011_d A1 0.00541429f $X=2.07 $Y=0.33 $X2=0 $Y2=0
cc_112 N_A_96_183#_c_99_n A1 0.013738f $X=1.58 $Y=1 $X2=0 $Y2=0
cc_113 N_A_96_183#_c_100_n A1 0.032071f $X=1.665 $Y=1.71 $X2=0 $Y2=0
cc_114 N_A_96_183#_c_113_n A1 0.0255205f $X=3.01 $Y=1.795 $X2=0 $Y2=0
cc_115 N_A_96_183#_c_101_n A1 0.0294874f $X=2.62 $Y=0.54 $X2=0 $Y2=0
cc_116 N_A_96_183#_c_103_n A1 0.0144844f $X=2.785 $Y=0.905 $X2=0 $Y2=0
cc_117 N_A_96_183#_c_99_n N_A1_c_271_n 0.00113937f $X=1.58 $Y=1 $X2=0 $Y2=0
cc_118 N_A_96_183#_c_103_n N_A1_c_271_n 5.84037e-19 $X=2.785 $Y=0.905 $X2=0
+ $Y2=0
cc_119 N_A_96_183#_c_101_n N_A1_c_272_n 0.00379826f $X=2.62 $Y=0.54 $X2=0 $Y2=0
cc_120 N_A_96_183#_c_113_n N_B1_c_313_n 0.0128416f $X=3.01 $Y=1.795 $X2=0 $Y2=0
cc_121 N_A_96_183#_c_104_n N_B1_c_313_n 0.00306335f $X=3.095 $Y=1.71 $X2=0 $Y2=0
cc_122 N_A_96_183#_c_101_n N_B1_M1000_g 0.0108715f $X=2.62 $Y=0.54 $X2=0 $Y2=0
cc_123 N_A_96_183#_c_102_n N_B1_M1000_g 0.0105137f $X=3.01 $Y=0.905 $X2=0 $Y2=0
cc_124 N_A_96_183#_c_103_n N_B1_M1000_g 0.00334221f $X=2.785 $Y=0.905 $X2=0
+ $Y2=0
cc_125 N_A_96_183#_c_104_n N_B1_M1000_g 0.00643565f $X=3.095 $Y=1.71 $X2=0 $Y2=0
cc_126 N_A_96_183#_c_113_n N_B1_c_320_n 0.00693432f $X=3.01 $Y=1.795 $X2=0 $Y2=0
cc_127 N_A_96_183#_c_113_n B1 0.0213417f $X=3.01 $Y=1.795 $X2=0 $Y2=0
cc_128 N_A_96_183#_c_102_n B1 0.00285671f $X=3.01 $Y=0.905 $X2=0 $Y2=0
cc_129 N_A_96_183#_c_103_n B1 0.0220115f $X=2.785 $Y=0.905 $X2=0 $Y2=0
cc_130 N_A_96_183#_c_104_n B1 0.0237534f $X=3.095 $Y=1.71 $X2=0 $Y2=0
cc_131 N_A_96_183#_c_113_n N_B1_c_316_n 0.0044678f $X=3.01 $Y=1.795 $X2=0 $Y2=0
cc_132 N_A_96_183#_c_103_n N_B1_c_316_n 0.00199686f $X=2.785 $Y=0.905 $X2=0
+ $Y2=0
cc_133 N_A_96_183#_c_101_n N_B2_M1001_g 0.00182338f $X=2.62 $Y=0.54 $X2=0 $Y2=0
cc_134 N_A_96_183#_c_104_n N_B2_M1001_g 0.00949024f $X=3.095 $Y=1.71 $X2=0 $Y2=0
cc_135 N_A_96_183#_c_107_n N_B2_M1001_g 0.00300708f $X=3.095 $Y=0.905 $X2=0
+ $Y2=0
cc_136 N_A_96_183#_c_108_n N_B2_M1001_g 0.0119702f $X=4.155 $Y=0.65 $X2=0 $Y2=0
cc_137 N_A_96_183#_c_113_n N_B2_M1006_g 0.00361944f $X=3.01 $Y=1.795 $X2=0 $Y2=0
cc_138 N_A_96_183#_c_104_n N_B2_M1006_g 7.89164e-19 $X=3.095 $Y=1.71 $X2=0 $Y2=0
cc_139 N_A_96_183#_c_116_n N_B2_M1006_g 3.57329e-19 $X=4.46 $Y=2.185 $X2=0 $Y2=0
cc_140 N_A_96_183#_c_113_n B2 0.00542587f $X=3.01 $Y=1.795 $X2=0 $Y2=0
cc_141 N_A_96_183#_c_104_n B2 0.0339949f $X=3.095 $Y=1.71 $X2=0 $Y2=0
cc_142 N_A_96_183#_c_108_n B2 0.0253375f $X=4.155 $Y=0.65 $X2=0 $Y2=0
cc_143 N_A_96_183#_c_104_n N_B2_c_370_n 0.00869468f $X=3.095 $Y=1.71 $X2=0 $Y2=0
cc_144 N_A_96_183#_c_108_n N_B2_c_370_n 0.00646843f $X=4.155 $Y=0.65 $X2=0 $Y2=0
cc_145 N_A_96_183#_c_108_n N_C1_c_411_n 0.00345935f $X=4.155 $Y=0.65 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_96_183#_c_109_n N_C1_c_411_n 0.00183473f $X=4.625 $Y=0.65 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_96_183#_c_108_n N_C1_c_412_n 0.00628469f $X=4.155 $Y=0.65 $X2=0 $Y2=0
cc_148 N_A_96_183#_c_108_n N_C1_c_413_n 0.00504154f $X=4.155 $Y=0.65 $X2=0 $Y2=0
cc_149 N_A_96_183#_c_108_n N_C1_c_414_n 0.00285973f $X=4.155 $Y=0.65 $X2=0 $Y2=0
cc_150 N_A_96_183#_c_109_n N_C1_c_414_n 0.0120828f $X=4.625 $Y=0.65 $X2=0 $Y2=0
cc_151 N_A_96_183#_c_116_n N_C1_M1002_g 0.0238409f $X=4.46 $Y=2.185 $X2=0 $Y2=0
cc_152 N_A_96_183#_c_110_n N_C1_M1002_g 0.0058018f $X=4.502 $Y=2.02 $X2=0 $Y2=0
cc_153 N_A_96_183#_c_108_n N_C1_c_415_n 0.00175146f $X=4.155 $Y=0.65 $X2=0 $Y2=0
cc_154 N_A_96_183#_c_109_n N_C1_c_415_n 0.00376901f $X=4.625 $Y=0.65 $X2=0 $Y2=0
cc_155 N_A_96_183#_c_108_n N_C1_c_416_n 0.00220795f $X=4.155 $Y=0.65 $X2=0 $Y2=0
cc_156 N_A_96_183#_c_109_n N_C1_c_416_n 6.99906e-19 $X=4.625 $Y=0.65 $X2=0 $Y2=0
cc_157 N_A_96_183#_c_110_n N_C1_c_416_n 0.00502213f $X=4.502 $Y=2.02 $X2=0 $Y2=0
cc_158 N_A_96_183#_c_108_n C1 0.0314368f $X=4.155 $Y=0.65 $X2=0 $Y2=0
cc_159 N_A_96_183#_c_116_n C1 0.00346926f $X=4.46 $Y=2.185 $X2=0 $Y2=0
cc_160 N_A_96_183#_c_110_n C1 0.0488284f $X=4.502 $Y=2.02 $X2=0 $Y2=0
cc_161 N_A_96_183#_c_109_n N_C1_c_419_n 0.00138157f $X=4.625 $Y=0.65 $X2=0 $Y2=0
cc_162 N_A_96_183#_c_110_n N_C1_c_419_n 0.0148853f $X=4.502 $Y=2.02 $X2=0 $Y2=0
cc_163 N_A_96_183#_M1010_g N_X_c_462_n 0.00883276f $X=0.735 $Y=0.54 $X2=0 $Y2=0
cc_164 N_A_96_183#_c_96_n N_X_c_462_n 0.00120799f $X=1.095 $Y=0.255 $X2=0 $Y2=0
cc_165 N_A_96_183#_c_105_n N_X_c_462_n 0.0141589f $X=0.645 $Y=1.08 $X2=0 $Y2=0
cc_166 N_A_96_183#_c_106_n N_X_c_462_n 0.001176f $X=0.645 $Y=1.08 $X2=0 $Y2=0
cc_167 N_A_96_183#_M1003_g X 0.0203465f $X=0.685 $Y=2.595 $X2=0 $Y2=0
cc_168 N_A_96_183#_c_98_n X 5.69591e-19 $X=0.645 $Y=1.585 $X2=0 $Y2=0
cc_169 N_A_96_183#_c_105_n X 0.0164013f $X=0.645 $Y=1.08 $X2=0 $Y2=0
cc_170 N_A_96_183#_M1003_g X 0.0334585f $X=0.685 $Y=2.595 $X2=0 $Y2=0
cc_171 N_A_96_183#_M1003_g N_X_c_463_n 0.0093333f $X=0.685 $Y=2.595 $X2=0 $Y2=0
cc_172 N_A_96_183#_M1010_g N_X_c_463_n 0.00360441f $X=0.735 $Y=0.54 $X2=0 $Y2=0
cc_173 N_A_96_183#_c_97_n N_X_c_463_n 0.0110821f $X=0.645 $Y=1.42 $X2=0 $Y2=0
cc_174 N_A_96_183#_c_105_n N_X_c_463_n 0.0478911f $X=0.645 $Y=1.08 $X2=0 $Y2=0
cc_175 N_A_96_183#_c_106_n N_X_c_463_n 0.00117201f $X=0.645 $Y=1.08 $X2=0 $Y2=0
cc_176 N_A_96_183#_M1003_g N_VPWR_c_489_n 0.00692475f $X=0.685 $Y=2.595 $X2=0
+ $Y2=0
cc_177 N_A_96_183#_M1003_g N_VPWR_c_492_n 0.00599594f $X=0.685 $Y=2.595 $X2=0
+ $Y2=0
cc_178 N_A_96_183#_c_116_n N_VPWR_c_493_n 0.0218588f $X=4.46 $Y=2.185 $X2=0
+ $Y2=0
cc_179 N_A_96_183#_M1003_g N_VPWR_c_488_n 0.00947311f $X=0.685 $Y=2.595 $X2=0
+ $Y2=0
cc_180 N_A_96_183#_c_116_n N_VPWR_c_488_n 0.0154967f $X=4.46 $Y=2.185 $X2=0
+ $Y2=0
cc_181 N_A_96_183#_c_113_n N_A_322_419#_c_534_n 0.0862815f $X=3.01 $Y=1.795
+ $X2=0 $Y2=0
cc_182 N_A_96_183#_c_113_n N_A_322_419#_c_535_n 0.013137f $X=3.01 $Y=1.795 $X2=0
+ $Y2=0
cc_183 N_A_96_183#_c_114_n N_A_322_419#_c_535_n 0.0142469f $X=1.75 $Y=1.795
+ $X2=0 $Y2=0
cc_184 N_A_96_183#_c_116_n N_A_545_400#_c_570_n 0.00890207f $X=4.46 $Y=2.185
+ $X2=0 $Y2=0
cc_185 N_A_96_183#_c_116_n N_A_545_400#_c_573_n 0.0586161f $X=4.46 $Y=2.185
+ $X2=0 $Y2=0
cc_186 N_A_96_183#_c_94_n N_VGND_c_601_n 0.0088238f $X=1.02 $Y=0.18 $X2=0 $Y2=0
cc_187 N_A_96_183#_c_99_n N_VGND_c_601_n 0.0233617f $X=1.58 $Y=1 $X2=0 $Y2=0
cc_188 N_A_96_183#_c_101_n N_VGND_c_602_n 0.0104546f $X=2.62 $Y=0.54 $X2=0 $Y2=0
cc_189 N_A_96_183#_c_108_n N_VGND_c_602_n 0.0226313f $X=4.155 $Y=0.65 $X2=0
+ $Y2=0
cc_190 N_A_96_183#_c_109_n N_VGND_c_602_n 0.0106155f $X=4.625 $Y=0.65 $X2=0
+ $Y2=0
cc_191 N_A_96_183#_c_95_n N_VGND_c_603_n 0.019388f $X=0.81 $Y=0.18 $X2=0 $Y2=0
cc_192 N_A_96_183#_c_101_n N_VGND_c_605_n 0.0173442f $X=2.62 $Y=0.54 $X2=0 $Y2=0
cc_193 N_A_96_183#_c_109_n N_VGND_c_606_n 0.0292523f $X=4.625 $Y=0.65 $X2=0
+ $Y2=0
cc_194 N_A_96_183#_c_94_n N_VGND_c_607_n 0.0237064f $X=1.02 $Y=0.18 $X2=0 $Y2=0
cc_195 N_A_96_183#_c_95_n N_VGND_c_607_n 0.0103891f $X=0.81 $Y=0.18 $X2=0 $Y2=0
cc_196 N_A_96_183#_c_101_n N_VGND_c_607_n 0.0122839f $X=2.62 $Y=0.54 $X2=0 $Y2=0
cc_197 N_A_96_183#_c_102_n N_VGND_c_607_n 0.00698459f $X=3.01 $Y=0.905 $X2=0
+ $Y2=0
cc_198 N_A_96_183#_c_107_n N_VGND_c_607_n 0.00658983f $X=3.095 $Y=0.905 $X2=0
+ $Y2=0
cc_199 N_A_96_183#_c_108_n N_VGND_c_607_n 0.0211591f $X=4.155 $Y=0.65 $X2=0
+ $Y2=0
cc_200 N_A_96_183#_c_109_n N_VGND_c_607_n 0.0208455f $X=4.625 $Y=0.65 $X2=0
+ $Y2=0
cc_201 N_A2_M1005_g N_A1_M1012_g 0.0272808f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_202 N_A2_c_229_n N_A1_M1012_g 3.49069e-19 $X=1.235 $Y=1.43 $X2=0 $Y2=0
cc_203 N_A2_c_228_n N_A1_c_269_n 0.026063f $X=1.235 $Y=1.43 $X2=0 $Y2=0
cc_204 N_A2_M1004_g A1 0.00281503f $X=1.605 $Y=0.54 $X2=0 $Y2=0
cc_205 N_A2_c_228_n N_A1_c_271_n 0.0345034f $X=1.235 $Y=1.43 $X2=0 $Y2=0
cc_206 N_A2_M1004_g N_A1_c_272_n 0.0345034f $X=1.605 $Y=0.54 $X2=0 $Y2=0
cc_207 N_A2_M1005_g X 0.00321251f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_208 N_A2_c_229_n X 9.9346e-19 $X=1.235 $Y=1.43 $X2=0 $Y2=0
cc_209 N_A2_M1005_g N_VPWR_c_489_n 0.00611108f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_210 N_A2_c_228_n N_VPWR_c_489_n 0.00199352f $X=1.235 $Y=1.43 $X2=0 $Y2=0
cc_211 N_A2_c_229_n N_VPWR_c_489_n 0.0210242f $X=1.235 $Y=1.43 $X2=0 $Y2=0
cc_212 N_A2_M1005_g N_VPWR_c_490_n 0.00939541f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_213 N_A2_M1005_g N_VPWR_c_491_n 0.00119667f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_214 N_A2_M1005_g N_VPWR_c_488_n 0.016444f $X=1.485 $Y=2.595 $X2=0 $Y2=0
cc_215 N_A2_M1005_g N_A_322_419#_c_539_n 0.0157038f $X=1.485 $Y=2.595 $X2=0
+ $Y2=0
cc_216 N_A2_M1005_g N_A_322_419#_c_535_n 0.00513626f $X=1.485 $Y=2.595 $X2=0
+ $Y2=0
cc_217 N_A2_c_228_n N_A_322_419#_c_535_n 0.00202318f $X=1.235 $Y=1.43 $X2=0
+ $Y2=0
cc_218 N_A2_M1004_g N_VGND_c_601_n 0.0113532f $X=1.605 $Y=0.54 $X2=0 $Y2=0
cc_219 N_A2_M1004_g N_VGND_c_605_n 0.00411131f $X=1.605 $Y=0.54 $X2=0 $Y2=0
cc_220 N_A2_M1004_g N_VGND_c_607_n 0.00781653f $X=1.605 $Y=0.54 $X2=0 $Y2=0
cc_221 N_A1_c_269_n N_B1_c_313_n 0.0230047f $X=2.09 $Y=1.36 $X2=0 $Y2=0
cc_222 N_A1_M1012_g N_B1_c_319_n 0.0230047f $X=2.015 $Y=2.595 $X2=0 $Y2=0
cc_223 A1 N_B1_M1000_g 0.0044006f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_224 N_A1_c_271_n N_B1_M1000_g 0.00610428f $X=2.095 $Y=1.025 $X2=0 $Y2=0
cc_225 N_A1_c_272_n N_B1_M1000_g 0.00567287f $X=2.09 $Y=0.86 $X2=0 $Y2=0
cc_226 N_A1_c_269_n B1 4.09964e-19 $X=2.09 $Y=1.36 $X2=0 $Y2=0
cc_227 A1 B1 0.0212609f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_228 N_A1_c_269_n N_B1_c_316_n 0.0189232f $X=2.09 $Y=1.36 $X2=0 $Y2=0
cc_229 A1 N_B1_c_316_n 0.00252902f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_230 N_A1_M1012_g N_VPWR_c_490_n 0.00840199f $X=2.015 $Y=2.595 $X2=0 $Y2=0
cc_231 N_A1_M1012_g N_VPWR_c_491_n 0.0169496f $X=2.015 $Y=2.595 $X2=0 $Y2=0
cc_232 N_A1_M1012_g N_VPWR_c_488_n 0.0136033f $X=2.015 $Y=2.595 $X2=0 $Y2=0
cc_233 N_A1_M1012_g N_A_322_419#_c_539_n 0.0183515f $X=2.015 $Y=2.595 $X2=0
+ $Y2=0
cc_234 N_A1_M1012_g N_A_322_419#_c_534_n 0.0182356f $X=2.015 $Y=2.595 $X2=0
+ $Y2=0
cc_235 N_A1_M1012_g N_A_322_419#_c_535_n 0.00116066f $X=2.015 $Y=2.595 $X2=0
+ $Y2=0
cc_236 A1 N_VGND_c_601_n 0.0117597f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_237 N_A1_c_272_n N_VGND_c_601_n 0.00211767f $X=2.09 $Y=0.86 $X2=0 $Y2=0
cc_238 A1 N_VGND_c_605_n 0.00979091f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_239 N_A1_c_272_n N_VGND_c_605_n 0.00339722f $X=2.09 $Y=0.86 $X2=0 $Y2=0
cc_240 A1 N_VGND_c_607_n 0.0112666f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_241 N_A1_c_272_n N_VGND_c_607_n 0.00505909f $X=2.09 $Y=0.86 $X2=0 $Y2=0
cc_242 N_B1_M1000_g N_B2_M1001_g 0.0339362f $X=2.835 $Y=0.54 $X2=0 $Y2=0
cc_243 B1 N_B2_M1001_g 2.85387e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_244 N_B1_c_320_n N_B2_M1006_g 0.0415629f $X=3.135 $Y=3.075 $X2=0 $Y2=0
cc_245 N_B1_c_320_n N_B2_c_370_n 0.00516146f $X=3.135 $Y=3.075 $X2=0 $Y2=0
cc_246 N_B1_c_316_n N_B2_c_370_n 0.0339362f $X=2.835 $Y=1.345 $X2=0 $Y2=0
cc_247 N_B1_c_313_n N_VPWR_c_491_n 0.010615f $X=2.575 $Y=3.075 $X2=0 $Y2=0
cc_248 N_B1_c_319_n N_VPWR_c_493_n 0.020601f $X=2.65 $Y=3.15 $X2=0 $Y2=0
cc_249 N_B1_c_318_n N_VPWR_c_488_n 0.0186572f $X=3.01 $Y=3.15 $X2=0 $Y2=0
cc_250 N_B1_c_319_n N_VPWR_c_488_n 0.0102451f $X=2.65 $Y=3.15 $X2=0 $Y2=0
cc_251 N_B1_c_313_n N_A_322_419#_c_539_n 8.52338e-19 $X=2.575 $Y=3.075 $X2=0
+ $Y2=0
cc_252 N_B1_c_313_n N_A_322_419#_c_534_n 0.0159459f $X=2.575 $Y=3.075 $X2=0
+ $Y2=0
cc_253 N_B1_c_320_n N_A_322_419#_c_534_n 0.0177128f $X=3.135 $Y=3.075 $X2=0
+ $Y2=0
cc_254 N_B1_c_313_n N_A_322_419#_c_548_n 7.78444e-19 $X=2.575 $Y=3.075 $X2=0
+ $Y2=0
cc_255 N_B1_c_320_n N_A_322_419#_c_548_n 0.0109697f $X=3.135 $Y=3.075 $X2=0
+ $Y2=0
cc_256 N_B1_c_313_n N_A_545_400#_c_569_n 0.00483321f $X=2.575 $Y=3.075 $X2=0
+ $Y2=0
cc_257 N_B1_c_320_n N_A_545_400#_c_569_n 0.0104467f $X=3.135 $Y=3.075 $X2=0
+ $Y2=0
cc_258 N_B1_c_320_n N_A_545_400#_c_570_n 0.0136128f $X=3.135 $Y=3.075 $X2=0
+ $Y2=0
cc_259 N_B1_c_313_n N_A_545_400#_c_571_n 9.8192e-19 $X=2.575 $Y=3.075 $X2=0
+ $Y2=0
cc_260 N_B1_c_318_n N_A_545_400#_c_571_n 0.0044168f $X=3.01 $Y=3.15 $X2=0 $Y2=0
cc_261 N_B1_c_320_n N_A_545_400#_c_571_n 0.00314811f $X=3.135 $Y=3.075 $X2=0
+ $Y2=0
cc_262 N_B1_c_320_n N_A_545_400#_c_573_n 0.00120317f $X=3.135 $Y=3.075 $X2=0
+ $Y2=0
cc_263 N_B1_M1000_g N_VGND_c_602_n 0.00162185f $X=2.835 $Y=0.54 $X2=0 $Y2=0
cc_264 N_B1_M1000_g N_VGND_c_605_n 0.0046526f $X=2.835 $Y=0.54 $X2=0 $Y2=0
cc_265 N_B1_M1000_g N_VGND_c_607_n 0.0053614f $X=2.835 $Y=0.54 $X2=0 $Y2=0
cc_266 N_B2_M1001_g N_C1_c_411_n 0.0187636f $X=3.225 $Y=0.54 $X2=-0.19
+ $Y2=-0.245
cc_267 N_B2_c_370_n N_C1_c_413_n 0.00674646f $X=3.665 $Y=1.38 $X2=0 $Y2=0
cc_268 N_B2_M1006_g N_C1_M1002_g 0.0277645f $X=3.665 $Y=2.5 $X2=0 $Y2=0
cc_269 N_B2_M1006_g N_C1_c_417_n 0.0167253f $X=3.665 $Y=2.5 $X2=0 $Y2=0
cc_270 N_B2_M1001_g C1 2.83085e-19 $X=3.225 $Y=0.54 $X2=0 $Y2=0
cc_271 B2 C1 0.0362656f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_272 N_B2_c_370_n C1 0.00564652f $X=3.665 $Y=1.38 $X2=0 $Y2=0
cc_273 B2 N_C1_c_419_n 7.87189e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_274 N_B2_c_370_n N_C1_c_419_n 0.0167253f $X=3.665 $Y=1.38 $X2=0 $Y2=0
cc_275 N_B2_M1006_g N_VPWR_c_493_n 0.00502174f $X=3.665 $Y=2.5 $X2=0 $Y2=0
cc_276 N_B2_M1006_g N_VPWR_c_488_n 0.00675085f $X=3.665 $Y=2.5 $X2=0 $Y2=0
cc_277 N_B2_M1006_g N_A_322_419#_c_534_n 0.00493104f $X=3.665 $Y=2.5 $X2=0 $Y2=0
cc_278 B2 N_A_322_419#_c_534_n 0.00938893f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_279 N_B2_c_370_n N_A_322_419#_c_534_n 0.00404349f $X=3.665 $Y=1.38 $X2=0
+ $Y2=0
cc_280 N_B2_M1006_g N_A_322_419#_c_548_n 0.010058f $X=3.665 $Y=2.5 $X2=0 $Y2=0
cc_281 N_B2_M1006_g N_A_545_400#_c_569_n 8.96863e-19 $X=3.665 $Y=2.5 $X2=0 $Y2=0
cc_282 N_B2_M1006_g N_A_545_400#_c_570_n 0.0175127f $X=3.665 $Y=2.5 $X2=0 $Y2=0
cc_283 N_B2_M1006_g N_A_545_400#_c_573_n 0.019915f $X=3.665 $Y=2.5 $X2=0 $Y2=0
cc_284 N_B2_M1001_g N_VGND_c_602_n 0.0100197f $X=3.225 $Y=0.54 $X2=0 $Y2=0
cc_285 N_B2_M1001_g N_VGND_c_605_n 0.00411131f $X=3.225 $Y=0.54 $X2=0 $Y2=0
cc_286 N_B2_M1001_g N_VGND_c_607_n 0.0040384f $X=3.225 $Y=0.54 $X2=0 $Y2=0
cc_287 N_C1_M1002_g N_VPWR_c_493_n 0.00763034f $X=4.195 $Y=2.5 $X2=0 $Y2=0
cc_288 N_C1_M1002_g N_VPWR_c_488_n 0.0145365f $X=4.195 $Y=2.5 $X2=0 $Y2=0
cc_289 N_C1_M1002_g N_A_322_419#_c_548_n 2.20729e-19 $X=4.195 $Y=2.5 $X2=0 $Y2=0
cc_290 N_C1_M1002_g N_A_545_400#_c_570_n 0.0053574f $X=4.195 $Y=2.5 $X2=0 $Y2=0
cc_291 N_C1_M1002_g N_A_545_400#_c_573_n 0.0189602f $X=4.195 $Y=2.5 $X2=0 $Y2=0
cc_292 C1 N_A_545_400#_c_573_n 0.00841124f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_293 N_C1_c_411_n N_VGND_c_602_n 0.00742492f $X=3.745 $Y=0.825 $X2=0 $Y2=0
cc_294 N_C1_c_411_n N_VGND_c_606_n 0.00495161f $X=3.745 $Y=0.825 $X2=0 $Y2=0
cc_295 N_C1_c_414_n N_VGND_c_606_n 0.0046404f $X=4.105 $Y=0.825 $X2=0 $Y2=0
cc_296 N_C1_c_411_n N_VGND_c_607_n 0.0052607f $X=3.745 $Y=0.825 $X2=0 $Y2=0
cc_297 N_C1_c_414_n N_VGND_c_607_n 0.0054529f $X=4.105 $Y=0.825 $X2=0 $Y2=0
cc_298 X N_VPWR_c_492_n 0.0437825f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_299 N_X_M1003_s N_VPWR_c_488_n 0.0023218f $X=0.275 $Y=2.095 $X2=0 $Y2=0
cc_300 X N_VPWR_c_488_n 0.0261704f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_301 N_X_c_462_n N_VGND_c_601_n 0.00675204f $X=0.21 $Y=0.735 $X2=0 $Y2=0
cc_302 N_X_c_462_n N_VGND_c_603_n 0.0221557f $X=0.21 $Y=0.735 $X2=0 $Y2=0
cc_303 N_X_c_462_n N_VGND_c_607_n 0.0194213f $X=0.21 $Y=0.735 $X2=0 $Y2=0
cc_304 N_VPWR_c_488_n N_A_322_419#_M1005_d 0.00223819f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_305 N_VPWR_c_490_n N_A_322_419#_c_539_n 0.0177952f $X=2.115 $Y=3.33 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_491_n N_A_322_419#_c_539_n 0.0431584f $X=2.28 $Y=2.575 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_488_n N_A_322_419#_c_539_n 0.0123247f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_308 N_VPWR_M1012_d N_A_322_419#_c_534_n 0.00248253f $X=2.14 $Y=2.095 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_491_n N_A_322_419#_c_534_n 0.02102f $X=2.28 $Y=2.575 $X2=0 $Y2=0
cc_310 N_VPWR_c_491_n N_A_545_400#_c_569_n 0.0299607f $X=2.28 $Y=2.575 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_493_n N_A_545_400#_c_570_n 0.0650023f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_488_n N_A_545_400#_c_570_n 0.0377535f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_491_n N_A_545_400#_c_571_n 0.0111564f $X=2.28 $Y=2.575 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_493_n N_A_545_400#_c_571_n 0.0220964f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_488_n N_A_545_400#_c_571_n 0.0113949f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_316 N_A_322_419#_c_534_n N_A_545_400#_M1009_s 0.00477085f $X=3.235 $Y=2.145
+ $X2=-0.19 $Y2=1.655
cc_317 N_A_322_419#_c_534_n N_A_545_400#_c_569_n 0.0209956f $X=3.235 $Y=2.145
+ $X2=0 $Y2=0
cc_318 N_A_322_419#_c_548_n N_A_545_400#_c_569_n 0.0200967f $X=3.4 $Y=2.23 $X2=0
+ $Y2=0
cc_319 N_A_322_419#_M1009_d N_A_545_400#_c_570_n 0.00180746f $X=3.26 $Y=2 $X2=0
+ $Y2=0
cc_320 N_A_322_419#_c_534_n N_A_545_400#_c_570_n 0.00431681f $X=3.235 $Y=2.145
+ $X2=0 $Y2=0
cc_321 N_A_322_419#_c_548_n N_A_545_400#_c_570_n 0.0152642f $X=3.4 $Y=2.23 $X2=0
+ $Y2=0
cc_322 N_A_322_419#_c_534_n N_A_545_400#_c_573_n 0.0119061f $X=3.235 $Y=2.145
+ $X2=0 $Y2=0
cc_323 N_A_322_419#_c_548_n N_A_545_400#_c_573_n 0.031924f $X=3.4 $Y=2.23 $X2=0
+ $Y2=0
