* File: sky130_fd_sc_lp__nand2_lp.pxi.spice
* Created: Fri Aug 28 10:47:41 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2_LP%B N_B_M1000_g N_B_M1003_g N_B_M1002_g B B B B B
+ N_B_c_31_n N_B_c_32_n PM_SKY130_FD_SC_LP__NAND2_LP%B
x_PM_SKY130_FD_SC_LP__NAND2_LP%A N_A_M1004_g N_A_M1001_g N_A_M1005_g N_A_c_60_n
+ N_A_c_61_n A N_A_c_63_n PM_SKY130_FD_SC_LP__NAND2_LP%A
x_PM_SKY130_FD_SC_LP__NAND2_LP%Y N_Y_M1004_d N_Y_M1003_d N_Y_c_87_n N_Y_c_88_n
+ N_Y_c_96_n N_Y_c_89_n Y Y PM_SKY130_FD_SC_LP__NAND2_LP%Y
x_PM_SKY130_FD_SC_LP__NAND2_LP%VPWR N_VPWR_M1002_d N_VPWR_c_123_n VPWR
+ N_VPWR_c_124_n N_VPWR_c_125_n N_VPWR_c_122_n N_VPWR_c_127_n
+ PM_SKY130_FD_SC_LP__NAND2_LP%VPWR
x_PM_SKY130_FD_SC_LP__NAND2_LP%VGND N_VGND_M1000_s N_VGND_c_140_n N_VGND_c_141_n
+ VGND N_VGND_c_142_n N_VGND_c_143_n PM_SKY130_FD_SC_LP__NAND2_LP%VGND
cc_1 VNB N_B_M1000_g 0.0309029f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.495
cc_2 VNB N_B_M1003_g 0.00146606f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.045
cc_3 VNB N_B_c_31_n 0.102851f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_4 VNB N_B_c_32_n 0.00570936f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_5 VNB N_A_M1004_g 0.0289344f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.495
cc_6 VNB N_A_M1001_g 0.00646847f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.045
cc_7 VNB N_A_c_60_n 0.0215617f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_8 VNB N_A_c_61_n 0.0192176f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.69
cc_9 VNB A 0.0319158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_c_63_n 0.0292927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_Y_c_87_n 0.00641568f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.735
cc_12 VNB N_Y_c_88_n 0.00322923f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.735
cc_13 VNB N_Y_c_89_n 0.0223736f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_VPWR_c_122_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_140_n 0.0117944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_141_n 0.0258732f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.045
cc_17 VNB N_VGND_c_142_n 0.0301668f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_VGND_c_143_n 0.118434f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_19 VPB N_B_M1003_g 0.0378647f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.045
cc_20 VPB N_B_c_32_n 0.0537862f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_21 VPB N_A_M1001_g 0.0495993f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.045
cc_22 VPB N_Y_c_87_n 0.00300018f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.735
cc_23 VPB Y 0.0316446f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_123_n 0.00776111f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.045
cc_25 VPB N_VPWR_c_124_n 0.0186227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_VPWR_c_125_n 0.0189497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_122_n 0.0658886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_127_n 0.00619952f $X=-0.19 $Y=1.655 $X2=0.355 $Y2=1.12
cc_29 N_B_M1000_g N_A_M1004_g 0.0233489f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_30 N_B_c_31_n N_A_c_60_n 0.0233489f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_31 N_B_M1003_g N_A_c_61_n 0.0269287f $X=0.53 $Y=2.045 $X2=0 $Y2=0
cc_32 N_B_M1000_g A 6.0997e-19 $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_33 N_B_c_31_n N_A_c_63_n 0.0269287f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_34 N_B_c_32_n A_39_367# 0.0144046f $X=0.27 $Y=1.12 $X2=-0.19 $Y2=-0.245
cc_35 N_B_M1000_g N_Y_c_87_n 0.0106386f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_36 N_B_M1003_g N_Y_c_87_n 0.00968287f $X=0.53 $Y=2.045 $X2=0 $Y2=0
cc_37 N_B_c_31_n N_Y_c_87_n 0.0157347f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_38 N_B_c_32_n N_Y_c_87_n 0.0788471f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_39 N_B_M1000_g N_Y_c_96_n 0.00408602f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_40 N_B_M1000_g N_Y_c_89_n 9.29579e-19 $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_41 N_B_M1003_g N_VPWR_c_123_n 0.0152407f $X=0.53 $Y=2.045 $X2=0 $Y2=0
cc_42 N_B_c_32_n N_VPWR_c_123_n 0.0145454f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_43 N_B_M1003_g N_VPWR_c_124_n 0.00471276f $X=0.53 $Y=2.045 $X2=0 $Y2=0
cc_44 N_B_c_32_n N_VPWR_c_124_n 0.00934611f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_45 N_B_M1003_g N_VPWR_c_122_n 0.0045449f $X=0.53 $Y=2.045 $X2=0 $Y2=0
cc_46 N_B_c_32_n N_VPWR_c_122_n 0.0102088f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_47 N_B_M1000_g N_VGND_c_141_n 0.00543702f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_48 N_B_c_31_n N_VGND_c_141_n 0.0018737f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_49 N_B_c_32_n N_VGND_c_141_n 0.0176025f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_50 N_B_M1000_g N_VGND_c_142_n 0.00509035f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_51 N_B_M1000_g N_VGND_c_143_n 0.0100767f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_52 N_A_M1004_g N_Y_c_87_n 0.00499856f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_53 A N_Y_c_87_n 0.048526f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_54 N_A_c_63_n N_Y_c_87_n 0.00866941f $X=1.055 $Y=1.07 $X2=0 $Y2=0
cc_55 N_A_M1004_g N_Y_c_88_n 0.0108614f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_56 A N_Y_c_88_n 0.00290608f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_57 N_A_M1004_g N_Y_c_89_n 0.00801279f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_58 N_A_c_60_n N_Y_c_89_n 0.00168007f $X=1.032 $Y=1.055 $X2=0 $Y2=0
cc_59 A N_Y_c_89_n 0.0239666f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_60 N_A_M1001_g Y 0.0269842f $X=0.96 $Y=2.045 $X2=0 $Y2=0
cc_61 N_A_c_61_n Y 0.00132428f $X=1.052 $Y=1.575 $X2=0 $Y2=0
cc_62 A Y 0.0252656f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A_M1001_g N_VPWR_c_123_n 0.0277269f $X=0.96 $Y=2.045 $X2=0 $Y2=0
cc_64 N_A_M1001_g N_VPWR_c_125_n 0.00471276f $X=0.96 $Y=2.045 $X2=0 $Y2=0
cc_65 N_A_M1001_g N_VPWR_c_122_n 0.0045449f $X=0.96 $Y=2.045 $X2=0 $Y2=0
cc_66 N_A_M1004_g N_VGND_c_142_n 0.00367856f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_67 N_A_M1004_g N_VGND_c_143_n 0.0058278f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_68 N_Y_c_87_n N_VPWR_c_123_n 0.0125284f $X=0.665 $Y=1.815 $X2=0 $Y2=0
cc_69 Y N_VPWR_c_123_n 0.0113972f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_70 Y A_207_367# 0.00990353f $X=1.115 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_71 N_Y_c_96_n N_VGND_c_141_n 0.00702103f $X=0.75 $Y=0.64 $X2=0 $Y2=0
cc_72 N_Y_c_89_n N_VGND_c_141_n 0.00436551f $X=1.135 $Y=0.495 $X2=0 $Y2=0
cc_73 N_Y_c_88_n N_VGND_c_142_n 0.00396191f $X=0.97 $Y=0.64 $X2=0 $Y2=0
cc_74 N_Y_c_96_n N_VGND_c_142_n 0.00327294f $X=0.75 $Y=0.64 $X2=0 $Y2=0
cc_75 N_Y_c_89_n N_VGND_c_142_n 0.0214013f $X=1.135 $Y=0.495 $X2=0 $Y2=0
cc_76 N_Y_c_88_n N_VGND_c_143_n 0.00605815f $X=0.97 $Y=0.64 $X2=0 $Y2=0
cc_77 N_Y_c_96_n N_VGND_c_143_n 0.00534138f $X=0.75 $Y=0.64 $X2=0 $Y2=0
cc_78 N_Y_c_89_n N_VGND_c_143_n 0.0124501f $X=1.135 $Y=0.495 $X2=0 $Y2=0
cc_79 N_Y_c_88_n A_121_57# 5.83038e-19 $X=0.97 $Y=0.64 $X2=-0.19 $Y2=-0.245
cc_80 N_Y_c_96_n A_121_57# 0.00145152f $X=0.75 $Y=0.64 $X2=-0.19 $Y2=-0.245
