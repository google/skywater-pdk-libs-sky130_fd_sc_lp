* File: sky130_fd_sc_lp__dlrbp_2.pex.spice
* Created: Wed Sep  2 09:46:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRBP_2%A_80_21# 1 2 9 13 17 21 23 28 31 35 39 41
c49 35 0 1.77994e-19 $X=2.02 $Y=0.885
r50 37 41 5.47651 $w=3.07e-07 $l=1.75656e-07 $layer=LI1_cond $X=2.062 $Y=1.63
+ $X2=2.04 $Y2=1.465
r51 37 39 14.355 $w=2.83e-07 $l=3.55e-07 $layer=LI1_cond $X=2.062 $Y=1.63
+ $X2=2.062 $Y2=1.985
r52 33 41 5.47651 $w=3.07e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=1.3
+ $X2=2.04 $Y2=1.465
r53 33 35 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.04 $Y=1.3
+ $X2=2.04 $Y2=0.885
r54 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.465 $X2=1.165 $Y2=1.465
r55 28 41 1.08954 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=1.465
+ $X2=2.04 $Y2=1.465
r56 28 30 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.875 $Y=1.465
+ $X2=1.165 $Y2=1.465
r57 26 27 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.905 $Y=1.465
+ $X2=0.91 $Y2=1.465
r58 24 26 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.465
+ $X2=0.905 $Y2=1.465
r59 23 31 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.985 $Y=1.465
+ $X2=1.165 $Y2=1.465
r60 23 27 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.985 $Y=1.465
+ $X2=0.91 $Y2=1.465
r61 19 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.63
+ $X2=0.91 $Y2=1.465
r62 19 21 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=0.91 $Y=1.63
+ $X2=0.91 $Y2=2.465
r63 15 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.3
+ $X2=0.905 $Y2=1.465
r64 15 17 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.905 $Y=1.3
+ $X2=0.905 $Y2=0.655
r65 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.63
+ $X2=0.475 $Y2=1.465
r66 11 13 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=0.475 $Y=1.63
+ $X2=0.475 $Y2=2.465
r67 7 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.3
+ $X2=0.475 $Y2=1.465
r68 7 9 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.475 $Y=1.3
+ $X2=0.475 $Y2=0.655
r69 2 39 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=1.835 $X2=2.1 $Y2=1.985
r70 1 35 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.675 $X2=2.02 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%A_432_109# 1 2 7 9 12 14 16 19 21 23 26 30
+ 34 39 40 42 43 44 46 48 52 55 63 64 72
c137 63 0 1.79023e-19 $X=4.97 $Y=1.62
c138 55 0 1.9533e-19 $X=3.2 $Y=1.37
c139 14 0 1.77994e-19 $X=2.86 $Y=1.205
r140 69 70 57.3559 $w=4.58e-07 $l=5.45e-07 $layer=POLY_cond $X=2.315 $Y=1.445
+ $X2=2.86 $Y2=1.445
r141 64 73 26.7778 $w=2.52e-07 $l=1.4e-07 $layer=POLY_cond $X=4.97 $Y=1.62
+ $X2=4.83 $Y2=1.62
r142 63 66 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=4.97 $Y=1.62
+ $X2=4.97 $Y2=1.8
r143 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.97
+ $Y=1.62 $X2=4.97 $Y2=1.62
r144 60 61 2.48416 $w=2.21e-07 $l=4.5e-08 $layer=LI1_cond $X=4.055 $Y=1.96
+ $X2=4.055 $Y2=2.005
r145 58 60 8.83258 $w=2.21e-07 $l=1.6e-07 $layer=LI1_cond $X=4.055 $Y=1.8
+ $X2=4.055 $Y2=1.96
r146 56 72 9.47162 $w=4.58e-07 $l=9e-08 $layer=POLY_cond $X=3.2 $Y=1.445
+ $X2=3.29 $Y2=1.445
r147 56 70 35.7817 $w=4.58e-07 $l=3.4e-07 $layer=POLY_cond $X=3.2 $Y=1.445
+ $X2=2.86 $Y2=1.445
r148 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.2
+ $Y=1.37 $X2=3.2 $Y2=1.37
r149 50 52 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.405 $Y=0.835
+ $X2=4.405 $Y2=0.42
r150 49 58 2.27611 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.185 $Y=1.8
+ $X2=4.055 $Y2=1.8
r151 48 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=1.8
+ $X2=4.97 $Y2=1.8
r152 48 49 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.805 $Y=1.8
+ $X2=4.185 $Y2=1.8
r153 44 61 4.29794 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=2.09
+ $X2=4.055 $Y2=2.005
r154 44 46 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=4.055 $Y=2.09
+ $X2=4.055 $Y2=2.91
r155 42 61 2.27611 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.925 $Y=2.005
+ $X2=4.055 $Y2=2.005
r156 42 43 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.925 $Y=2.005
+ $X2=3.335 $Y2=2.005
r157 41 55 3.70735 $w=2.5e-07 $l=2.18403e-07 $layer=LI1_cond $X=3.335 $Y=1.09
+ $X2=3.25 $Y2=1.27
r158 40 50 28.0067 $w=2.21e-07 $l=5.35817e-07 $layer=LI1_cond $X=3.91 $Y=1.09
+ $X2=4.405 $Y2=1.005
r159 40 41 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.91 $Y=1.09
+ $X2=3.335 $Y2=1.09
r160 39 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.25 $Y=1.92
+ $X2=3.335 $Y2=2.005
r161 38 55 2.76166 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.25 $Y=1.535
+ $X2=3.25 $Y2=1.27
r162 38 39 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.25 $Y=1.535
+ $X2=3.25 $Y2=1.92
r163 32 64 55.4683 $w=2.52e-07 $l=3.63249e-07 $layer=POLY_cond $X=5.26 $Y=1.455
+ $X2=4.97 $Y2=1.62
r164 32 34 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=5.26 $Y=1.455
+ $X2=5.26 $Y2=0.805
r165 28 73 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.83 $Y=1.785
+ $X2=4.83 $Y2=1.62
r166 28 30 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.83 $Y=1.785 $X2=4.83
+ $Y2=2.725
r167 24 72 29.2056 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.29 $Y=1.685
+ $X2=3.29 $Y2=1.445
r168 24 26 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.29 $Y=1.685
+ $X2=3.29 $Y2=2.465
r169 21 72 29.2056 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.29 $Y=1.205
+ $X2=3.29 $Y2=1.445
r170 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.29 $Y=1.205
+ $X2=3.29 $Y2=0.675
r171 17 70 29.2056 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.86 $Y=1.685
+ $X2=2.86 $Y2=1.445
r172 17 19 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.86 $Y=1.685
+ $X2=2.86 $Y2=2.465
r173 14 70 29.2056 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.86 $Y=1.205
+ $X2=2.86 $Y2=1.445
r174 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.86 $Y=1.205
+ $X2=2.86 $Y2=0.675
r175 10 69 29.2056 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.315 $Y=1.685
+ $X2=2.315 $Y2=1.445
r176 10 12 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.315 $Y=1.685
+ $X2=2.315 $Y2=2.155
r177 7 69 8.41921 $w=4.58e-07 $l=2.77128e-07 $layer=POLY_cond $X=2.235 $Y=1.205
+ $X2=2.315 $Y2=1.445
r178 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.235 $Y=1.205
+ $X2=2.235 $Y2=0.885
r179 2 60 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.835 $X2=4.09 $Y2=1.96
r180 2 46 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.835 $X2=4.09 $Y2=2.91
r181 1 52 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=4.265
+ $Y=0.255 $X2=4.405 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%RESET_B 3 5 7 8 12
c36 5 0 1.9533e-19 $X=3.875 $Y=1.715
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=1.51 $X2=3.74 $Y2=1.51
r38 8 12 5.58215 $w=3.18e-07 $l=1.55e-07 $layer=LI1_cond $X=3.665 $Y=1.665
+ $X2=3.665 $Y2=1.51
r39 5 11 44.3014 $w=3.48e-07 $l=2.55323e-07 $layer=POLY_cond $X=3.875 $Y=1.715
+ $X2=3.762 $Y2=1.51
r40 5 7 241 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=3.875 $Y=1.715 $X2=3.875
+ $Y2=2.465
r41 1 11 38.7612 $w=3.48e-07 $l=1.96074e-07 $layer=POLY_cond $X=3.83 $Y=1.345
+ $X2=3.762 $Y2=1.51
r42 1 3 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=3.83 $Y=1.345 $X2=3.83
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%A_823_25# 1 2 7 9 12 14 17 20 29 31 33 34 37
c84 37 0 3.79235e-20 $X=4.305 $Y=1.37
c85 33 0 1.66518e-19 $X=5.73 $Y=2.45
r86 33 34 9.98589 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=5.725 $Y=2.45
+ $X2=5.725 $Y2=2.275
r87 26 29 4.57319 $w=3.13e-07 $l=1.25e-07 $layer=LI1_cond $X=5.71 $Y=0.797
+ $X2=5.835 $Y2=0.797
r88 24 37 12.5521 $w=2.88e-07 $l=7.5e-08 $layer=POLY_cond $X=4.38 $Y=1.37
+ $X2=4.305 $Y2=1.37
r89 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.38
+ $Y=1.37 $X2=4.38 $Y2=1.37
r90 20 23 3.90659 $w=2.93e-07 $l=1e-07 $layer=LI1_cond $X=4.397 $Y=1.27
+ $X2=4.397 $Y2=1.37
r91 18 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.71 $Y=1.355
+ $X2=5.71 $Y2=1.27
r92 18 34 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.71 $Y=1.355
+ $X2=5.71 $Y2=2.275
r93 17 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.71 $Y=1.185
+ $X2=5.71 $Y2=1.27
r94 16 26 4.34843 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=5.71 $Y=0.955
+ $X2=5.71 $Y2=0.797
r95 16 17 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.71 $Y=0.955
+ $X2=5.71 $Y2=1.185
r96 15 20 3.96227 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=4.545 $Y=1.27
+ $X2=4.397 $Y2=1.27
r97 14 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=1.27
+ $X2=5.71 $Y2=1.27
r98 14 15 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=5.625 $Y=1.27
+ $X2=4.545 $Y2=1.27
r99 10 37 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.535
+ $X2=4.305 $Y2=1.37
r100 10 12 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=4.305 $Y=1.535
+ $X2=4.305 $Y2=2.465
r101 7 37 19.2465 $w=2.88e-07 $l=2.14942e-07 $layer=POLY_cond $X=4.19 $Y=1.205
+ $X2=4.305 $Y2=1.37
r102 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.19 $Y=1.205
+ $X2=4.19 $Y2=0.675
r103 2 33 600 $w=1.7e-07 $l=2.65518e-07 $layer=licon1_PDIFF $count=1 $X=5.495
+ $Y=2.515 $X2=5.73 $Y2=2.45
r104 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.695
+ $Y=0.595 $X2=5.835 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%A_1023_405# 1 2 9 13 16 19 20 22 24 25 28 30
+ 32 34 35 38 42 45 47 51 54
c137 51 0 1.41099e-19 $X=5.42 $Y=2.19
c138 32 0 1.44644e-19 $X=7.7 $Y=2.64
r139 44 47 7.62646 $w=3.38e-07 $l=2.25e-07 $layer=LI1_cond $X=7.7 $Y=2.81
+ $X2=7.925 $Y2=2.81
r140 44 45 5.76029 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=7.7 $Y=2.81
+ $X2=7.615 $Y2=2.81
r141 39 42 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=7.7 $Y=0.445
+ $X2=7.855 $Y2=0.445
r142 35 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.07 $Y=1.29
+ $X2=6.07 $Y2=1.125
r143 34 37 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=1.29
+ $X2=6.065 $Y2=1.455
r144 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.07
+ $Y=1.29 $X2=6.07 $Y2=1.29
r145 32 44 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.7 $Y=2.64 $X2=7.7
+ $Y2=2.81
r146 31 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.7 $Y=0.61 $X2=7.7
+ $Y2=0.445
r147 31 32 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=7.7 $Y=0.61
+ $X2=7.7 $Y2=2.64
r148 30 45 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.035 $Y=2.895
+ $X2=7.615 $Y2=2.895
r149 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.95 $Y=2.81
+ $X2=7.035 $Y2=2.895
r150 27 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.95 $Y=2.525
+ $X2=6.95 $Y2=2.81
r151 26 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.165 $Y=2.44
+ $X2=6.08 $Y2=2.44
r152 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.865 $Y=2.44
+ $X2=6.95 $Y2=2.525
r153 25 26 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.865 $Y=2.44
+ $X2=6.165 $Y2=2.44
r154 23 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.08 $Y=2.525
+ $X2=6.08 $Y2=2.44
r155 23 24 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.08 $Y=2.525
+ $X2=6.08 $Y2=2.785
r156 22 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.08 $Y=2.355
+ $X2=6.08 $Y2=2.44
r157 22 37 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=6.08 $Y=2.355
+ $X2=6.08 $Y2=1.455
r158 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.995 $Y=2.87
+ $X2=6.08 $Y2=2.785
r159 19 20 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.995 $Y=2.87
+ $X2=5.445 $Y2=2.87
r160 17 51 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.28 $Y=2.19
+ $X2=5.42 $Y2=2.19
r161 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.28
+ $Y=2.19 $X2=5.28 $Y2=2.19
r162 14 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.28 $Y=2.785
+ $X2=5.445 $Y2=2.87
r163 14 16 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=5.28 $Y=2.785
+ $X2=5.28 $Y2=2.19
r164 13 54 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.05 $Y=0.805
+ $X2=6.05 $Y2=1.125
r165 7 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.42 $Y=2.355
+ $X2=5.42 $Y2=2.19
r166 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.42 $Y=2.355
+ $X2=5.42 $Y2=2.725
r167 2 47 600 $w=1.7e-07 $l=4.48163e-07 $layer=licon1_PDIFF $count=1 $X=7.8
+ $Y=2.415 $X2=7.925 $Y2=2.805
r168 1 42 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=7.73
+ $Y=0.235 $X2=7.855 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%A_1246_339# 1 2 9 13 17 20 21 24 28 30 31 36
r76 30 31 9.5763 $w=2.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.32 $Y=2.475
+ $X2=7.32 $Y2=2.3
r77 26 28 4.23118 $w=2.15e-07 $l=1.33918e-07 $layer=LI1_cond $X=7.35 $Y=1.27
+ $X2=7.252 $Y2=1.185
r78 26 31 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=7.35 $Y=1.27
+ $X2=7.35 $Y2=2.3
r79 22 28 4.23118 $w=2.15e-07 $l=1.07912e-07 $layer=LI1_cond $X=7.2 $Y=1.1
+ $X2=7.252 $Y2=1.185
r80 22 24 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=7.2 $Y=1.1 $X2=7.2
+ $Y2=0.805
r81 20 28 2.20034 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.07 $Y=1.185
+ $X2=7.252 $Y2=1.185
r82 20 21 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=7.07 $Y=1.185
+ $X2=6.595 $Y2=1.185
r83 18 36 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.43 $Y=1.86 $X2=6.52
+ $Y2=1.86
r84 18 33 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.43 $Y=1.86
+ $X2=6.305 $Y2=1.86
r85 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.43
+ $Y=1.86 $X2=6.43 $Y2=1.86
r86 15 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.465 $Y=1.27
+ $X2=6.595 $Y2=1.185
r87 15 17 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=6.465 $Y=1.27
+ $X2=6.465 $Y2=1.86
r88 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.52 $Y=1.695
+ $X2=6.52 $Y2=1.86
r89 11 13 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=6.52 $Y=1.695
+ $X2=6.52 $Y2=0.805
r90 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=2.025
+ $X2=6.305 $Y2=1.86
r91 7 9 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.305 $Y=2.025
+ $X2=6.305 $Y2=2.615
r92 2 30 600 $w=1.7e-07 $l=2.47386e-07 $layer=licon1_PDIFF $count=1 $X=7.14
+ $Y=2.295 $X2=7.3 $Y2=2.475
r93 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.025
+ $Y=0.595 $X2=7.165 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%D 3 7 11 12 13 14 18
r48 13 14 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.93 $Y=1.615
+ $X2=6.93 $Y2=2.035
r49 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7 $Y=1.615
+ $X2=7 $Y2=1.615
r50 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7 $Y=1.955 $X2=7
+ $Y2=1.615
r51 11 12 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7 $Y=1.955 $X2=7
+ $Y2=2.12
r52 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7 $Y=1.45 $X2=7
+ $Y2=1.615
r53 7 12 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.065 $Y=2.615
+ $X2=7.065 $Y2=2.12
r54 3 10 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=6.95 $Y=0.805
+ $X2=6.95 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%A_1109_21# 1 2 10 11 12 15 18 19 20 21 23 28
+ 30 33 34 35 36 39 40 42 43 46 49 53 55
c125 15 0 1.66518e-19 $X=5.945 $Y=2.615
r126 51 53 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=8.715 $Y=0.445
+ $X2=8.935 $Y2=0.445
r127 49 55 3.6114 $w=2.57e-07 $l=1.17707e-07 $layer=LI1_cond $X=8.935 $Y=2.3
+ $X2=8.857 $Y2=2.385
r128 48 53 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.935 $Y=0.61
+ $X2=8.935 $Y2=0.445
r129 48 49 104.131 $w=1.78e-07 $l=1.69e-06 $layer=LI1_cond $X=8.935 $Y=0.61
+ $X2=8.935 $Y2=2.3
r130 44 55 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=8.857 $Y=2.47
+ $X2=8.857 $Y2=2.385
r131 44 46 3.09612 $w=3.33e-07 $l=9e-08 $layer=LI1_cond $X=8.857 $Y=2.47
+ $X2=8.857 $Y2=2.56
r132 42 55 2.87242 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=8.69 $Y=2.385
+ $X2=8.857 $Y2=2.385
r133 42 43 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=8.69 $Y=2.385
+ $X2=8.135 $Y2=2.385
r134 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.05
+ $Y=1.75 $X2=8.05 $Y2=1.75
r135 37 43 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=8.045 $Y=2.3
+ $X2=8.135 $Y2=2.385
r136 37 39 33.8889 $w=1.78e-07 $l=5.5e-07 $layer=LI1_cond $X=8.045 $Y=2.3
+ $X2=8.045 $Y2=1.75
r137 34 40 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.05 $Y=2.09
+ $X2=8.05 $Y2=1.75
r138 34 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.05 $Y=2.09
+ $X2=8.05 $Y2=2.255
r139 33 40 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.05 $Y=1.585
+ $X2=8.05 $Y2=1.75
r140 30 31 98.522 $w=1.59e-07 $l=3.25e-07 $layer=POLY_cond $X=5.62 $Y=1.755
+ $X2=5.945 $Y2=1.755
r141 28 35 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.14 $Y=2.735
+ $X2=8.14 $Y2=2.255
r142 24 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.07 $Y=0.915
+ $X2=8.07 $Y2=0.84
r143 24 33 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=8.07 $Y=0.915
+ $X2=8.07 $Y2=1.585
r144 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.07 $Y=0.765
+ $X2=8.07 $Y2=0.84
r145 21 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.07 $Y=0.765
+ $X2=8.07 $Y2=0.445
r146 19 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.995 $Y=0.84
+ $X2=8.07 $Y2=0.84
r147 19 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.995 $Y=0.84
+ $X2=7.655 $Y2=0.84
r148 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.58 $Y=0.765
+ $X2=7.655 $Y2=0.84
r149 17 18 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.58 $Y=0.255
+ $X2=7.58 $Y2=0.765
r150 13 31 4.22461 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.945 $Y=1.845
+ $X2=5.945 $Y2=1.755
r151 13 15 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.945 $Y=1.845
+ $X2=5.945 $Y2=2.615
r152 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.505 $Y=0.18
+ $X2=7.58 $Y2=0.255
r153 11 12 928.106 $w=1.5e-07 $l=1.81e-06 $layer=POLY_cond $X=7.505 $Y=0.18
+ $X2=5.695 $Y2=0.18
r154 8 30 4.22461 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.62 $Y=1.665 $X2=5.62
+ $Y2=1.755
r155 8 10 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.62 $Y=1.665
+ $X2=5.62 $Y2=0.805
r156 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.62 $Y=0.255
+ $X2=5.695 $Y2=0.18
r157 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.62 $Y=0.255
+ $X2=5.62 $Y2=0.805
r158 2 46 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.645
+ $Y=2.415 $X2=8.79 $Y2=2.56
r159 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.575
+ $Y=0.235 $X2=8.715 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%GATE 3 7 11 12 13 14 15 16 22
c35 3 0 1.44644e-19 $X=8.5 $Y=0.445
r36 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.59
+ $Y=1.005 $X2=8.59 $Y2=1.005
r37 15 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.49 $Y=1.665
+ $X2=8.49 $Y2=2.035
r38 14 15 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.49 $Y=1.295
+ $X2=8.49 $Y2=1.665
r39 14 23 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.49 $Y=1.295
+ $X2=8.49 $Y2=1.005
r40 13 23 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=8.49 $Y=0.925 $X2=8.49
+ $Y2=1.005
r41 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.59 $Y=1.345
+ $X2=8.59 $Y2=1.005
r42 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.59 $Y=1.345
+ $X2=8.59 $Y2=1.51
r43 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.59 $Y=0.84
+ $X2=8.59 $Y2=1.005
r44 7 12 628.138 $w=1.5e-07 $l=1.225e-06 $layer=POLY_cond $X=8.57 $Y=2.735
+ $X2=8.57 $Y2=1.51
r45 3 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.5 $Y=0.445 $X2=8.5
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%VPWR 1 2 3 4 5 6 7 22 24 30 36 40 44 50 54
+ 56 58 63 68 73 78 86 96 97 103 106 109 112 115 118
r118 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r119 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r120 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r121 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r124 97 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r125 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r126 94 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.52 $Y=3.33
+ $X2=8.355 $Y2=3.33
r127 94 96 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.52 $Y=3.33
+ $X2=8.88 $Y2=3.33
r128 93 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r129 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r130 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 90 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r132 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r133 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r134 87 115 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.525 $Y2=3.33
r135 87 89 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.96 $Y2=3.33
r136 86 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=8.355 $Y2=3.33
r137 86 92 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=7.92 $Y2=3.33
r138 85 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r139 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r140 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r141 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r142 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r143 79 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.685 $Y=3.33
+ $X2=4.52 $Y2=3.33
r144 79 81 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.685 $Y=3.33
+ $X2=5.04 $Y2=3.33
r145 78 115 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.355 $Y=3.33
+ $X2=6.525 $Y2=3.33
r146 78 84 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.355 $Y=3.33
+ $X2=6 $Y2=3.33
r147 77 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r148 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r149 74 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.58 $Y2=3.33
r150 74 76 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=4.08 $Y2=3.33
r151 73 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.52 $Y2=3.33
r152 73 76 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.08 $Y2=3.33
r153 72 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r154 72 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r155 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r156 69 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=3.33
+ $X2=2.625 $Y2=3.33
r157 69 71 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.79 $Y=3.33
+ $X2=3.12 $Y2=3.33
r158 68 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.58 $Y2=3.33
r159 68 71 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.12 $Y2=3.33
r160 67 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r161 67 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r162 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r163 64 103 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.145 $Y2=3.33
r164 64 66 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=2.16 $Y2=3.33
r165 63 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=3.33
+ $X2=2.625 $Y2=3.33
r166 63 66 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.46 $Y=3.33 $X2=2.16
+ $Y2=3.33
r167 62 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 62 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r169 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r170 59 100 4.40339 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.192 $Y2=3.33
r171 59 61 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.72 $Y2=3.33
r172 58 103 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1 $Y=3.33
+ $X2=1.145 $Y2=3.33
r173 58 61 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r174 56 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r175 56 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r176 56 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r177 52 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=3.245
+ $X2=8.355 $Y2=3.33
r178 52 54 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.355 $Y=3.245
+ $X2=8.355 $Y2=2.765
r179 48 115 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.525 $Y=3.245
+ $X2=6.525 $Y2=3.33
r180 48 50 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=6.525 $Y=3.245
+ $X2=6.525 $Y2=2.81
r181 44 47 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=4.52 $Y=2.14
+ $X2=4.52 $Y2=2.95
r182 42 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.52 $Y2=3.33
r183 42 47 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.52 $Y2=2.95
r184 38 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.58 $Y2=3.33
r185 38 40 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.58 $Y2=2.38
r186 34 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=3.245
+ $X2=2.625 $Y2=3.33
r187 34 36 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=2.625 $Y=3.245
+ $X2=2.625 $Y2=2.79
r188 30 33 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=1.145 $Y=1.98
+ $X2=1.145 $Y2=2.95
r189 28 103 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=3.33
r190 28 33 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.145 $Y=3.245
+ $X2=1.145 $Y2=2.95
r191 24 27 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=0.24 $Y=1.98
+ $X2=0.24 $Y2=2.95
r192 22 100 3.03446 $w=2.9e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.192 $Y2=3.33
r193 22 27 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.95
r194 7 54 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=8.215
+ $Y=2.415 $X2=8.355 $Y2=2.765
r195 6 50 600 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=2.295 $X2=6.53 $Y2=2.81
r196 5 47 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.835 $X2=4.52 $Y2=2.95
r197 5 44 300 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=2 $X=4.38
+ $Y=1.835 $X2=4.52 $Y2=2.14
r198 4 40 300 $w=1.7e-07 $l=6.43584e-07 $layer=licon1_PDIFF $count=2 $X=3.365
+ $Y=1.835 $X2=3.58 $Y2=2.38
r199 3 36 600 $w=1.7e-07 $l=1.06604e-06 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.835 $X2=2.625 $Y2=2.79
r200 2 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.95
r201 2 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=1.98
r202 1 27 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r203 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%Q_N 1 2 7 8 9 14
r18 9 24 39.8117 $w=2.73e-07 $l=9.5e-07 $layer=LI1_cond $X=0.692 $Y=1.96
+ $X2=0.692 $Y2=2.91
r19 8 9 12.3626 $w=2.73e-07 $l=2.95e-07 $layer=LI1_cond $X=0.692 $Y=1.665
+ $X2=0.692 $Y2=1.96
r20 7 8 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.692 $Y=1.295
+ $X2=0.692 $Y2=1.665
r21 7 14 36.6686 $w=2.73e-07 $l=8.75e-07 $layer=LI1_cond $X=0.692 $Y=1.295
+ $X2=0.692 $Y2=0.42
r22 2 24 400 $w=1.7e-07 $l=1.14521e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.695 $Y2=2.91
r23 2 9 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.695 $Y2=1.96
r24 1 14 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%Q 1 2 8 9 10 13 15 16 17 18 25 31 34 38
r55 32 34 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.605 $Y=2.375
+ $X2=2.64 $Y2=2.375
r56 18 31 3.78936 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=3.1 $Y=2.375 $X2=2.96
+ $Y2=2.375
r57 18 38 12.8605 $w=4.48e-07 $l=4.2e-07 $layer=LI1_cond $X=3.1 $Y=2.49 $X2=3.1
+ $Y2=2.91
r58 17 25 4.50329 $w=2e-07 $l=9.88686e-08 $layer=LI1_cond $X=2.52 $Y=2.375
+ $X2=2.435 $Y2=2.405
r59 17 32 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.375 $X2=2.605
+ $Y2=2.375
r60 17 31 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.665 $Y=2.375
+ $X2=2.96 $Y2=2.375
r61 17 34 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.665 $Y=2.375
+ $X2=2.64 $Y2=2.375
r62 16 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.16 $Y=2.405
+ $X2=2.435 $Y2=2.405
r63 15 16 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.405
+ $X2=2.16 $Y2=2.405
r64 11 13 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=3.075 $Y=0.655
+ $X2=3.075 $Y2=0.39
r65 9 11 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.91 $Y=0.745
+ $X2=3.075 $Y2=0.655
r66 9 10 18.7929 $w=1.78e-07 $l=3.05e-07 $layer=LI1_cond $X=2.91 $Y=0.745
+ $X2=2.605 $Y2=0.745
r67 8 17 1.93381 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.52 $Y=2.26 $X2=2.52
+ $Y2=2.375
r68 7 10 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.52 $Y=0.835
+ $X2=2.605 $Y2=0.745
r69 7 8 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=2.52 $Y=0.835
+ $X2=2.52 $Y2=2.26
r70 2 18 600 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.835 $X2=3.075 $Y2=2.385
r71 2 38 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.835 $X2=3.075 $Y2=2.91
r72 1 13 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=2.935
+ $Y=0.255 $X2=3.075 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__DLRBP_2%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 48
+ 51 52 54 55 56 58 63 68 73 92 93 99 102 105 108
r110 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r111 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r112 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r113 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r114 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r115 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r116 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r117 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r118 87 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r119 86 89 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r120 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r121 84 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r122 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r123 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r124 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r125 80 83 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r126 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r127 78 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=0
+ $X2=5.045 $Y2=0
r128 78 80 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.52
+ $Y2=0
r129 74 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=0
+ $X2=3.575 $Y2=0
r130 74 76 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=4.56
+ $Y2=0
r131 73 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.88 $Y=0
+ $X2=5.045 $Y2=0
r132 73 76 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=0 $X2=4.56
+ $Y2=0
r133 72 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r134 72 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=2.64 $Y2=0
r135 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r136 69 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=0
+ $X2=2.565 $Y2=0
r137 69 71 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.73 $Y=0 $X2=3.12
+ $Y2=0
r138 68 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=0
+ $X2=3.575 $Y2=0
r139 68 71 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.41 $Y=0 $X2=3.12
+ $Y2=0
r140 67 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r141 67 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r142 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r143 64 99 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.142 $Y2=0
r144 64 66 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=2.16 $Y2=0
r145 63 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.565
+ $Y2=0
r146 63 66 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r147 62 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r148 62 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r149 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r150 59 96 4.40339 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=0
+ $X2=0.192 $Y2=0
r151 59 61 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=0
+ $X2=0.72 $Y2=0
r152 58 99 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=1 $Y=0 $X2=1.142
+ $Y2=0
r153 58 61 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1 $Y=0 $X2=0.72
+ $Y2=0
r154 56 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r155 56 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r156 56 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r157 54 89 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.15 $Y=0 $X2=7.92
+ $Y2=0
r158 54 55 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.15 $Y=0 $X2=8.282
+ $Y2=0
r159 53 92 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.415 $Y=0
+ $X2=8.88 $Y2=0
r160 53 55 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.415 $Y=0
+ $X2=8.282 $Y2=0
r161 51 83 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.57 $Y=0 $X2=6.48
+ $Y2=0
r162 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.57 $Y=0 $X2=6.735
+ $Y2=0
r163 50 86 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=6.9 $Y=0 $X2=6.96
+ $Y2=0
r164 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.9 $Y=0 $X2=6.735
+ $Y2=0
r165 46 55 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=8.282 $Y=0.085
+ $X2=8.282 $Y2=0
r166 46 48 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=8.282 $Y=0.085
+ $X2=8.282 $Y2=0.445
r167 42 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.735 $Y=0.085
+ $X2=6.735 $Y2=0
r168 42 44 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=6.735 $Y=0.085
+ $X2=6.735 $Y2=0.805
r169 38 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0.085
+ $X2=5.045 $Y2=0
r170 38 40 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=5.045 $Y=0.085
+ $X2=5.045 $Y2=0.805
r171 34 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0
r172 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0.38
r173 30 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=0.085
+ $X2=2.565 $Y2=0
r174 30 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.565 $Y=0.085
+ $X2=2.565 $Y2=0.38
r175 26 99 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.142 $Y=0.085
+ $X2=1.142 $Y2=0
r176 26 28 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=1.142 $Y=0.085
+ $X2=1.142 $Y2=0.38
r177 22 96 3.03446 $w=2.9e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.192 $Y2=0
r178 22 24 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.38
r179 7 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.145
+ $Y=0.235 $X2=8.285 $Y2=0.445
r180 6 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.595
+ $Y=0.595 $X2=6.735 $Y2=0.805
r181 5 40 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=4.92
+ $Y=0.595 $X2=5.045 $Y2=0.805
r182 4 36 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=3.365
+ $Y=0.255 $X2=3.575 $Y2=0.38
r183 3 32 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.675 $X2=2.565 $Y2=0.38
r184 2 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.38
r185 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

