* File: sky130_fd_sc_lp__ha_1.pex.spice
* Created: Wed Sep  2 09:54:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__HA_1%A_80_30# 1 2 9 12 14 18 20 23 24 28 30 34 37
r62 31 34 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.34
+ $X2=1.715 $Y2=2.34
r63 28 38 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.395
+ $X2=0.597 $Y2=1.56
r64 28 37 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.395
+ $X2=0.597 $Y2=1.23
r65 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.395 $X2=0.63 $Y2=1.395
r66 24 27 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=0.665 $Y=1.315
+ $X2=0.665 $Y2=1.395
r67 23 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=2.175
+ $X2=1.63 $Y2=2.34
r68 22 23 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.63 $Y=1.4
+ $X2=1.63 $Y2=2.175
r69 21 30 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.37 $Y=1.315
+ $X2=1.225 $Y2=1.315
r70 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.545 $Y=1.315
+ $X2=1.63 $Y2=1.4
r71 20 21 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.545 $Y=1.315
+ $X2=1.37 $Y2=1.315
r72 16 30 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=1.23
+ $X2=1.225 $Y2=1.315
r73 16 18 28.215 $w=2.88e-07 $l=7.1e-07 $layer=LI1_cond $X=1.225 $Y=1.23
+ $X2=1.225 $Y2=0.52
r74 15 24 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.795 $Y=1.315
+ $X2=0.665 $Y2=1.315
r75 14 30 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.08 $Y=1.315
+ $X2=1.225 $Y2=1.315
r76 14 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.08 $Y=1.315
+ $X2=0.795 $Y2=1.315
r77 12 38 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=0.615 $Y=2.465
+ $X2=0.615 $Y2=1.56
r78 9 37 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.7
+ $X2=0.475 $Y2=1.23
r79 2 34 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=2.14 $X2=1.715 $Y2=2.34
r80 1 18 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.31 $X2=1.245 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__HA_1%A_223_320# 1 2 9 13 17 20 24 27 28 30 31 32 33
+ 39 42 44 47 48 50 51 53 56
c136 53 0 6.14124e-20 $X=1.46 $Y=1.765
r137 53 54 6.14013 $w=3.14e-07 $l=4e-08 $layer=POLY_cond $X=1.46 $Y=1.765
+ $X2=1.5 $Y2=1.765
r138 48 57 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=4.172 $Y=1.425
+ $X2=4.172 $Y2=1.59
r139 48 56 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=4.172 $Y=1.425
+ $X2=4.172 $Y2=1.26
r140 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.14
+ $Y=1.425 $X2=4.14 $Y2=1.425
r141 45 51 0.221902 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=3.68 $Y=1.425
+ $X2=3.56 $Y2=1.425
r142 45 47 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=3.68 $Y=1.425
+ $X2=4.14 $Y2=1.425
r143 44 50 3.70735 $w=2.5e-07 $l=8.9861e-08 $layer=LI1_cond $X=3.56 $Y=1.93
+ $X2=3.55 $Y2=2.015
r144 43 51 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=1.59
+ $X2=3.56 $Y2=1.425
r145 43 44 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=3.56 $Y=1.59
+ $X2=3.56 $Y2=1.93
r146 42 51 7.38875 $w=2.1e-07 $l=1.79374e-07 $layer=LI1_cond $X=3.53 $Y=1.26
+ $X2=3.56 $Y2=1.425
r147 41 42 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=3.53 $Y=1.06 $X2=3.53
+ $Y2=1.26
r148 37 50 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.1 $X2=3.55
+ $Y2=2.015
r149 37 39 10.6379 $w=2.58e-07 $l=2.4e-07 $layer=LI1_cond $X=3.55 $Y=2.1
+ $X2=3.55 $Y2=2.34
r150 33 41 7.42255 $w=3.05e-07 $l=1.92819e-07 $layer=LI1_cond $X=3.44 $Y=0.907
+ $X2=3.53 $Y2=1.06
r151 33 35 13.4137 $w=3.03e-07 $l=3.55e-07 $layer=LI1_cond $X=3.44 $Y=0.907
+ $X2=3.085 $Y2=0.907
r152 31 50 2.76166 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.42 $Y=2.015
+ $X2=3.55 $Y2=2.015
r153 31 32 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.42 $Y=2.015
+ $X2=2.47 $Y2=2.015
r154 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.385 $Y=2.1
+ $X2=2.47 $Y2=2.015
r155 29 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.385 $Y=2.1
+ $X2=2.385 $Y2=2.675
r156 27 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.3 $Y=2.78
+ $X2=2.385 $Y2=2.675
r157 27 28 49.381 $w=2.08e-07 $l=9.35e-07 $layer=LI1_cond $X=2.3 $Y=2.78
+ $X2=1.365 $Y2=2.78
r158 25 53 27.6306 $w=3.14e-07 $l=1.8e-07 $layer=POLY_cond $X=1.28 $Y=1.765
+ $X2=1.46 $Y2=1.765
r159 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.28
+ $Y=1.765 $X2=1.28 $Y2=1.765
r160 22 28 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.28 $Y=2.675
+ $X2=1.365 $Y2=2.78
r161 22 24 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.28 $Y=2.675
+ $X2=1.28 $Y2=1.765
r162 20 57 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.295 $Y=2.465
+ $X2=4.295 $Y2=1.59
r163 17 56 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.215 $Y=0.73
+ $X2=4.215 $Y2=1.26
r164 11 54 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.93 $X2=1.5
+ $Y2=1.765
r165 11 13 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.5 $Y=1.93 $X2=1.5
+ $Y2=2.35
r166 7 53 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.46 $Y=1.6 $X2=1.46
+ $Y2=1.765
r167 7 9 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=1.46 $Y=1.6 $X2=1.46
+ $Y2=0.52
r168 2 39 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=2.14 $X2=3.515 $Y2=2.34
r169 1 35 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.73 $X2=3.085 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_LP__HA_1%B 3 7 9 11 14 18 19 22 25 26 28 33 35
c88 35 0 1.23857e-19 $X=3.3 $Y=1.425
c89 25 0 6.14124e-20 $X=1.98 $Y=1.345
c90 22 0 1.3617e-19 $X=2.96 $Y=1.315
r91 32 35 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.12 $Y=1.425 $X2=3.3
+ $Y2=1.425
r92 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.425 $X2=3.12 $Y2=1.425
r93 28 33 8.92214 $w=3.08e-07 $l=2.4e-07 $layer=LI1_cond $X=3.115 $Y=1.665
+ $X2=3.115 $Y2=1.425
r94 27 33 0.92939 $w=3.08e-07 $l=2.5e-08 $layer=LI1_cond $X=3.115 $Y=1.4
+ $X2=3.115 $Y2=1.425
r95 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.98
+ $Y=1.345 $X2=1.98 $Y2=1.345
r96 23 25 4.21847 $w=1.7e-07 $l=1.41951e-07 $layer=LI1_cond $X=2.145 $Y=1.315
+ $X2=2.015 $Y2=1.29
r97 22 27 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=2.96 $Y=1.315
+ $X2=3.115 $Y2=1.4
r98 22 23 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.96 $Y=1.315
+ $X2=2.145 $Y2=1.315
r99 18 26 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=1.98 $Y=1.735
+ $X2=1.98 $Y2=1.345
r100 18 19 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=1.735
+ $X2=1.98 $Y2=1.9
r101 17 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=1.18
+ $X2=1.98 $Y2=1.345
r102 12 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.59
+ $X2=3.3 $Y2=1.425
r103 12 14 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.3 $Y=1.59 $X2=3.3
+ $Y2=2.35
r104 9 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.26 $X2=3.3
+ $Y2=1.425
r105 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.3 $Y=1.26 $X2=3.3
+ $Y2=0.94
r106 7 19 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.93 $Y=2.35
+ $X2=1.93 $Y2=1.9
r107 3 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.89 $Y=0.52
+ $X2=1.89 $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_LP__HA_1%A 1 3 8 10 11 13 14 15 19 22 28 29 32 34
c91 29 0 1.23857e-19 $X=2.64 $Y=1.665
c92 19 0 2.66955e-19 $X=3.69 $Y=0.94
r93 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.55 $Y=1.665
+ $X2=2.55 $Y2=1.83
r94 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.55 $Y=1.665
+ $X2=2.55 $Y2=1.5
r95 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.55
+ $Y=1.665 $X2=2.55 $Y2=1.665
r96 29 33 5.25359 $w=1.88e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=1.665 $X2=2.55
+ $Y2=1.665
r97 27 28 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=3.71 $Y=1.83
+ $X2=3.71 $Y2=1.98
r98 24 26 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.32 $Y=0.915
+ $X2=2.46 $Y2=0.915
r99 22 28 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.73 $Y=2.35
+ $X2=3.73 $Y2=1.98
r100 19 27 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.69 $Y=0.94
+ $X2=3.69 $Y2=1.83
r101 16 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.69 $Y=0.36
+ $X2=3.69 $Y2=0.94
r102 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.615 $Y=0.285
+ $X2=3.69 $Y2=0.36
r103 14 15 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.615 $Y=0.285
+ $X2=2.885 $Y2=0.285
r104 12 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.81 $Y=0.36
+ $X2=2.885 $Y2=0.285
r105 12 13 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.81 $Y=0.36
+ $X2=2.81 $Y2=0.84
r106 11 26 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.535 $Y=0.915
+ $X2=2.46 $Y2=0.915
r107 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.735 $Y=0.915
+ $X2=2.81 $Y2=0.84
r108 10 11 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.735 $Y=0.915
+ $X2=2.535 $Y2=0.915
r109 8 35 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.46 $Y=2.35
+ $X2=2.46 $Y2=1.83
r110 4 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.46 $Y=0.99
+ $X2=2.46 $Y2=0.915
r111 4 34 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.46 $Y=0.99
+ $X2=2.46 $Y2=1.5
r112 1 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.32 $Y=0.84
+ $X2=2.32 $Y2=0.915
r113 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.32 $Y=0.84 $X2=2.32
+ $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__HA_1%SUM 1 2 7 8 9 10 11 12 13 24 34 37
r16 35 37 0.983793 $w=4.08e-07 $l=3.5e-08 $layer=LI1_cond $X=0.3 $Y=1.945
+ $X2=0.3 $Y2=1.98
r17 34 48 3.20123 $w=2.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.23 $Y=1.665
+ $X2=0.23 $Y2=1.74
r18 13 45 3.79463 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=0.3 $Y=2.775
+ $X2=0.3 $Y2=2.91
r19 12 13 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.3 $Y=2.405 $X2=0.3
+ $Y2=2.775
r20 11 12 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.3 $Y=2.035 $X2=0.3
+ $Y2=2.405
r21 11 37 1.54596 $w=4.08e-07 $l=5.5e-08 $layer=LI1_cond $X=0.3 $Y=2.035 $X2=0.3
+ $Y2=1.98
r22 10 35 5.62167 $w=4.08e-07 $l=2e-07 $layer=LI1_cond $X=0.3 $Y=1.745 $X2=0.3
+ $Y2=1.945
r23 10 48 1.48481 $w=4.08e-07 $l=5e-09 $layer=LI1_cond $X=0.3 $Y=1.745 $X2=0.3
+ $Y2=1.74
r24 10 34 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=0.23 $Y=1.66 $X2=0.23
+ $Y2=1.665
r25 9 10 15.5793 $w=2.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.23 $Y=1.295
+ $X2=0.23 $Y2=1.66
r26 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=0.925 $X2=0.23
+ $Y2=1.295
r27 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=0.555 $X2=0.23
+ $Y2=0.925
r28 7 24 5.5488 $w=2.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.23 $Y=0.555 $X2=0.23
+ $Y2=0.425
r29 2 45 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.835 $X2=0.4 $Y2=2.91
r30 2 37 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.835 $X2=0.4 $Y2=1.98
r31 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.28 $X2=0.26 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_LP__HA_1%VPWR 1 2 3 12 20 24 31 32 33 39 43 50 51 54 59
c59 24 0 1.30785e-19 $X=4.08 $Y=1.98
r60 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 55 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 54 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r64 51 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r66 48 59 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.037 $Y2=3.33
r67 48 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.56 $Y2=3.33
r68 47 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r69 47 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r71 44 54 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=3.25 $Y=3.33
+ $X2=2.945 $Y2=3.33
r72 44 46 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=3.33 $X2=3.6
+ $Y2=3.33
r73 43 59 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=3.85 $Y=3.33
+ $X2=4.037 $Y2=3.33
r74 43 46 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.85 $Y=3.33 $X2=3.6
+ $Y2=3.33
r75 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r76 39 54 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=2.945 $Y2=3.33
r77 39 41 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r78 37 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r79 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 33 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 33 42 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r82 31 36 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r83 31 32 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.875 $Y2=3.33
r84 30 41 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.2 $Y2=3.33
r85 30 32 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.875 $Y2=3.33
r86 27 29 15.9805 $w=3.73e-07 $l=5.2e-07 $layer=LI1_cond $X=4.037 $Y=2.43
+ $X2=4.037 $Y2=2.95
r87 24 27 13.8293 $w=3.73e-07 $l=4.5e-07 $layer=LI1_cond $X=4.037 $Y=1.98
+ $X2=4.037 $Y2=2.43
r88 22 59 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.037 $Y=3.245
+ $X2=4.037 $Y2=3.33
r89 22 29 9.06588 $w=3.73e-07 $l=2.95e-07 $layer=LI1_cond $X=4.037 $Y=3.245
+ $X2=4.037 $Y2=2.95
r90 18 54 2.55884 $w=6.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=3.245
+ $X2=2.945 $Y2=3.33
r91 18 20 15.8824 $w=6.08e-07 $l=8.1e-07 $layer=LI1_cond $X=2.945 $Y=3.245
+ $X2=2.945 $Y2=2.435
r92 15 17 18.247 $w=2.98e-07 $l=4.75e-07 $layer=LI1_cond $X=0.875 $Y=2.475
+ $X2=0.875 $Y2=2.95
r93 12 15 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=0.875 $Y=1.98
+ $X2=0.875 $Y2=2.475
r94 10 32 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=3.33
r95 10 17 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=2.95
r96 3 29 600 $w=1.7e-07 $l=9.3747e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=2.14 $X2=4.08 $Y2=2.95
r97 3 27 600 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=2.14 $X2=3.945 $Y2=2.43
r98 3 24 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=2.14 $X2=4.08 $Y2=1.98
r99 2 20 300 $w=1.7e-07 $l=6.81726e-07 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=2.14 $X2=3.085 $Y2=2.435
r100 1 17 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.835 $X2=0.83 $Y2=2.95
r101 1 15 600 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.835 $X2=0.83 $Y2=2.475
r102 1 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.835 $X2=0.83 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__HA_1%COUT 1 2 7 8 9 10 11 12 13 24 45
r16 22 45 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=4.52 $Y=0.895
+ $X2=4.52 $Y2=0.925
r17 13 42 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=4.555 $Y=2.775
+ $X2=4.555 $Y2=2.91
r18 12 13 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=4.555 $Y=2.405
+ $X2=4.555 $Y2=2.775
r19 11 12 15.3059 $w=3.18e-07 $l=4.25e-07 $layer=LI1_cond $X=4.555 $Y=1.98
+ $X2=4.555 $Y2=2.405
r20 10 11 11.3444 $w=3.18e-07 $l=3.15e-07 $layer=LI1_cond $X=4.555 $Y=1.665
+ $X2=4.555 $Y2=1.98
r21 9 10 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=4.555 $Y=1.295
+ $X2=4.555 $Y2=1.665
r22 9 47 7.38284 $w=3.18e-07 $l=2.05e-07 $layer=LI1_cond $X=4.555 $Y=1.295
+ $X2=4.555 $Y2=1.09
r23 8 47 4.48322 $w=3.88e-07 $l=1.38e-07 $layer=LI1_cond $X=4.52 $Y=0.952
+ $X2=4.52 $Y2=1.09
r24 8 45 0.797845 $w=3.88e-07 $l=2.7e-08 $layer=LI1_cond $X=4.52 $Y=0.952
+ $X2=4.52 $Y2=0.925
r25 8 22 0.827395 $w=3.88e-07 $l=2.8e-08 $layer=LI1_cond $X=4.52 $Y=0.867
+ $X2=4.52 $Y2=0.895
r26 7 8 9.21954 $w=3.88e-07 $l=3.12e-07 $layer=LI1_cond $X=4.52 $Y=0.555
+ $X2=4.52 $Y2=0.867
r27 7 24 2.95498 $w=3.88e-07 $l=1e-07 $layer=LI1_cond $X=4.52 $Y=0.555 $X2=4.52
+ $Y2=0.455
r28 2 42 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.835 $X2=4.51 $Y2=2.91
r29 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.37
+ $Y=1.835 $X2=4.51 $Y2=1.98
r30 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.29
+ $Y=0.31 $X2=4.43 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__HA_1%VGND 1 2 3 12 16 20 25 26 27 29 34 47 48 51 54
r55 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r56 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r57 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r58 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r59 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r60 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r61 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r62 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r63 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.105
+ $Y2=0
r64 39 41 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.64
+ $Y2=0
r65 38 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r66 38 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r67 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r68 35 51 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.695
+ $Y2=0
r69 35 37 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.68
+ $Y2=0
r70 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.105
+ $Y2=0
r71 34 37 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.68
+ $Y2=0
r72 32 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r73 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r74 29 51 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.695
+ $Y2=0
r75 29 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r76 27 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r77 27 55 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r78 25 44 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.79 $Y=0 $X2=3.6
+ $Y2=0
r79 25 26 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.79 $Y=0 $X2=3.972
+ $Y2=0
r80 24 47 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.155 $Y=0 $X2=4.56
+ $Y2=0
r81 24 26 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=4.155 $Y=0 $X2=3.972
+ $Y2=0
r82 20 22 14.8397 $w=3.63e-07 $l=4.7e-07 $layer=LI1_cond $X=3.972 $Y=0.455
+ $X2=3.972 $Y2=0.925
r83 18 26 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.972 $Y=0.085
+ $X2=3.972 $Y2=0
r84 18 20 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.972 $Y=0.085
+ $X2=3.972 $Y2=0.455
r85 14 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r86 14 16 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.52
r87 10 51 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0
r88 10 12 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0.425
r89 3 22 182 $w=1.7e-07 $l=2.73998e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.73 $X2=3.955 $Y2=0.925
r90 3 20 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.73 $X2=4 $Y2=0.455
r91 2 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.31 $X2=2.105 $Y2=0.52
r92 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.28 $X2=0.69 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_LP__HA_1%A_307_62# 1 2 9 11 12 15
r27 13 15 14.1839 $w=2.58e-07 $l=3.2e-07 $layer=LI1_cond $X=2.57 $Y=0.84
+ $X2=2.57 $Y2=0.52
r28 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.44 $Y=0.925
+ $X2=2.57 $Y2=0.84
r29 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.44 $Y=0.925
+ $X2=1.77 $Y2=0.925
r30 7 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.655 $Y=0.84
+ $X2=1.77 $Y2=0.925
r31 7 9 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.655 $Y=0.84 $X2=1.655
+ $Y2=0.52
r32 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.31 $X2=2.535 $Y2=0.52
r33 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.31 $X2=1.675 $Y2=0.52
.ends

