* File: sky130_fd_sc_lp__clkbuflp_16.spice
* Created: Wed Sep  2 09:38:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkbuflp_16.pex.spice"
.subckt sky130_fd_sc_lp__clkbuflp_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1018 A_110_47# N_A_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75010.8 A=0.0825 P=1.4 MULT=1
MM1002 N_A_130_417#_M1002_d N_A_M1002_g A_110_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.5
+ SB=75010.5 A=0.0825 P=1.4 MULT=1
MM1007 N_A_130_417#_M1002_d N_A_M1007_g A_584_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001
+ SB=75010 A=0.0825 P=1.4 MULT=1
MM1009 A_584_47# N_A_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75001.3 SB=75009.7
+ A=0.0825 P=1.4 MULT=1
MM1021 A_268_47# N_A_M1021_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75001.8 SB=75009.3
+ A=0.0825 P=1.4 MULT=1
MM1033 N_A_130_417#_M1033_d N_A_M1033_g A_268_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75002.1
+ SB=75008.9 A=0.0825 P=1.4 MULT=1
MM1038 N_A_130_417#_M1033_d N_A_M1038_g A_426_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75002.6
+ SB=75008.5 A=0.0825 P=1.4 MULT=1
MM1035 A_426_47# N_A_M1035_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.55 AD=0.05775
+ AS=0.0825 PD=0.76 PS=0.85 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75002.9 SB=75008.1
+ A=0.0825 P=1.4 MULT=1
MM1010 A_1378_47# N_A_130_417#_M1010_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.0825 PD=0.76 PS=0.85 NRD=10.908 NRS=4.356 M=1 R=3.66667
+ SA=75003.4 SB=75007.7 A=0.0825 P=1.4 MULT=1
MM1000 N_X_M1000_d N_A_130_417#_M1000_g A_1378_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75003.7
+ SB=75007.3 A=0.0825 P=1.4 MULT=1
MM1001 N_X_M1000_d N_A_130_417#_M1001_g A_2010_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75004.2
+ SB=75006.9 A=0.0825 P=1.4 MULT=1
MM1008 A_2010_47# N_A_130_417#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75004.5
+ SB=75006.5 A=0.0825 P=1.4 MULT=1
MM1040 A_1852_47# N_A_130_417#_M1040_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75004.9
+ SB=75006.1 A=0.0825 P=1.4 MULT=1
MM1003 N_X_M1003_d N_A_130_417#_M1003_g A_1852_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75005.3
+ SB=75005.7 A=0.0825 P=1.4 MULT=1
MM1049 N_X_M1003_d N_A_130_417#_M1049_g A_746_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75005.7
+ SB=75005.3 A=0.0825 P=1.4 MULT=1
MM1011 A_746_47# N_A_130_417#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75006.1
+ SB=75004.9 A=0.0825 P=1.4 MULT=1
MM1019 A_904_47# N_A_130_417#_M1019_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75006.5
+ SB=75004.5 A=0.0825 P=1.4 MULT=1
MM1014 N_X_M1014_d N_A_130_417#_M1014_g A_904_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75006.9
+ SB=75004.1 A=0.0825 P=1.4 MULT=1
MM1030 N_X_M1014_d N_A_130_417#_M1030_g A_1536_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75007.3
+ SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1015 A_1536_47# N_A_130_417#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75007.7
+ SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1020 A_2168_47# N_A_130_417#_M1020_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75008.1
+ SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1032 N_X_M1032_d N_A_130_417#_M1032_g A_2168_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75008.5
+ SB=75002.6 A=0.0825 P=1.4 MULT=1
MM1027 N_X_M1032_d N_A_130_417#_M1027_g A_1062_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75008.9
+ SB=75002.1 A=0.0825 P=1.4 MULT=1
MM1024 A_1062_47# N_A_130_417#_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75009.3
+ SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1031 A_1220_47# N_A_130_417#_M1031_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75009.7
+ SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1028 N_X_M1028_d N_A_130_417#_M1028_g A_1220_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75010
+ SB=75001 A=0.0825 P=1.4 MULT=1
MM1036 N_X_M1028_d N_A_130_417#_M1036_g A_1694_47# VNB NSHORT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75010.5
+ SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1034 A_1694_47# N_A_130_417#_M1034_g N_VGND_M1034_s VNB NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75010.8 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_130_417#_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125011
+ A=0.25 P=2.5 MULT=1
MM1016 N_VPWR_M1016_d N_A_M1016_g N_A_130_417#_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125011 A=0.25
+ P=2.5 MULT=1
MM1025 N_VPWR_M1016_d N_A_M1025_g N_A_130_417#_M1025_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125010 A=0.25
+ P=2.5 MULT=1
MM1029 N_VPWR_M1029_d N_A_M1029_g N_A_130_417#_M1025_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125010 A=0.25
+ P=2.5 MULT=1
MM1046 N_VPWR_M1029_d N_A_M1046_g N_A_130_417#_M1046_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125009 A=0.25
+ P=2.5 MULT=1
MM1047 N_VPWR_M1047_d N_A_M1047_g N_A_130_417#_M1046_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125009 A=0.25
+ P=2.5 MULT=1
MM1004 N_VPWR_M1047_d N_A_130_417#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125008 A=0.25
+ P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_A_130_417#_M1006_g N_X_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125008 A=0.25
+ P=2.5 MULT=1
MM1012 N_VPWR_M1006_d N_A_130_417#_M1012_g N_X_M1012_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125004 SB=125007 A=0.25
+ P=2.5 MULT=1
MM1013 N_VPWR_M1013_d N_A_130_417#_M1013_g N_X_M1012_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125005 SB=125006 A=0.25
+ P=2.5 MULT=1
MM1017 N_VPWR_M1013_d N_A_130_417#_M1017_g N_X_M1017_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125005 SB=125006 A=0.25
+ P=2.5 MULT=1
MM1022 N_VPWR_M1022_d N_A_130_417#_M1022_g N_X_M1017_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125006 SB=125005 A=0.25
+ P=2.5 MULT=1
MM1023 N_VPWR_M1022_d N_A_130_417#_M1023_g N_X_M1023_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125006 SB=125005 A=0.25
+ P=2.5 MULT=1
MM1026 N_VPWR_M1026_d N_A_130_417#_M1026_g N_X_M1023_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125007 SB=125004 A=0.25
+ P=2.5 MULT=1
MM1037 N_VPWR_M1026_d N_A_130_417#_M1037_g N_X_M1037_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125008 SB=125004 A=0.25
+ P=2.5 MULT=1
MM1039 N_VPWR_M1039_d N_A_130_417#_M1039_g N_X_M1037_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125008 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1041 N_VPWR_M1039_d N_A_130_417#_M1041_g N_X_M1041_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125009 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1042 N_VPWR_M1042_d N_A_130_417#_M1042_g N_X_M1041_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125009 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1043 N_VPWR_M1042_d N_A_130_417#_M1043_g N_X_M1043_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125010 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1044 N_VPWR_M1044_d N_A_130_417#_M1044_g N_X_M1043_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125010 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1045 N_VPWR_M1044_d N_A_130_417#_M1045_g N_X_M1045_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125011 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1048 N_VPWR_M1048_d N_A_130_417#_M1048_g N_X_M1045_s VPB PHIGHVT L=0.25 W=1
+ AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125011 SB=125000
+ A=0.25 P=2.5 MULT=1
DX50_noxref VNB VPB NWDIODE A=23.9839 P=29.45
*
.include "sky130_fd_sc_lp__clkbuflp_16.pxi.spice"
*
.ends
*
*
