* File: sky130_fd_sc_lp__invlp_8.pxi.spice
* Created: Fri Aug 28 10:40:11 2020
* 
x_PM_SKY130_FD_SC_LP__INVLP_8%A N_A_M1001_g N_A_M1003_g N_A_M1004_g N_A_M1006_g
+ N_A_M1011_g N_A_M1010_g N_A_M1013_g N_A_M1017_g N_A_M1015_g N_A_M1020_g
+ N_A_M1016_g N_A_M1021_g N_A_M1022_g N_A_M1028_g N_A_M1000_g N_A_M1005_g
+ N_A_M1002_g N_A_M1008_g N_A_M1007_g N_A_M1012_g N_A_M1009_g N_A_M1018_g
+ N_A_M1014_g N_A_M1019_g N_A_M1025_g N_A_M1024_g N_A_M1026_g N_A_M1030_g
+ N_A_M1027_g N_A_M1031_g N_A_M1023_g N_A_M1029_g N_A_c_112_n N_A_c_113_n A A A
+ A N_A_c_133_n N_A_c_114_n N_A_c_135_n PM_SKY130_FD_SC_LP__INVLP_8%A
x_PM_SKY130_FD_SC_LP__INVLP_8%VPWR N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_M1017_d
+ N_VPWR_M1021_d N_VPWR_M1029_d N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n
+ N_VPWR_c_412_n N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n
+ N_VPWR_c_417_n N_VPWR_c_418_n N_VPWR_c_419_n VPWR N_VPWR_c_420_n
+ N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_408_n PM_SKY130_FD_SC_LP__INVLP_8%VPWR
x_PM_SKY130_FD_SC_LP__INVLP_8%A_114_367# N_A_114_367#_M1003_s
+ N_A_114_367#_M1010_s N_A_114_367#_M1020_s N_A_114_367#_M1028_s
+ N_A_114_367#_M1008_s N_A_114_367#_M1018_s N_A_114_367#_M1024_s
+ N_A_114_367#_M1031_s N_A_114_367#_c_518_n N_A_114_367#_c_520_n
+ N_A_114_367#_c_521_n N_A_114_367#_c_523_n N_A_114_367#_c_525_n
+ N_A_114_367#_c_527_n N_A_114_367#_c_529_n N_A_114_367#_c_533_n
+ N_A_114_367#_c_535_n N_A_114_367#_c_537_n N_A_114_367#_c_541_n
+ N_A_114_367#_c_543_n N_A_114_367#_c_547_n N_A_114_367#_c_549_n
+ N_A_114_367#_c_553_n N_A_114_367#_c_594_n N_A_114_367#_c_555_n
+ N_A_114_367#_c_557_n N_A_114_367#_c_596_n N_A_114_367#_c_558_n
+ N_A_114_367#_c_562_n N_A_114_367#_c_564_n N_A_114_367#_c_566_n
+ PM_SKY130_FD_SC_LP__INVLP_8%A_114_367#
x_PM_SKY130_FD_SC_LP__INVLP_8%Y N_Y_M1000_d N_Y_M1007_d N_Y_M1014_d N_Y_M1026_d
+ N_Y_M1005_d N_Y_M1012_d N_Y_M1019_d N_Y_M1030_d N_Y_c_632_n N_Y_c_640_n
+ N_Y_c_633_n N_Y_c_660_n N_Y_c_662_n N_Y_c_672_n N_Y_c_673_n N_Y_c_758_n
+ N_Y_c_634_n N_Y_c_679_n N_Y_c_683_n N_Y_c_635_n N_Y_c_689_n N_Y_c_693_n
+ N_Y_c_636_n N_Y_c_703_n N_Y_c_707_n N_Y_c_641_n N_Y_c_642_n N_Y_c_637_n
+ N_Y_c_718_n N_Y_c_638_n N_Y_c_723_n N_Y_c_639_n N_Y_c_729_n N_Y_c_731_n Y
+ PM_SKY130_FD_SC_LP__INVLP_8%Y
x_PM_SKY130_FD_SC_LP__INVLP_8%VGND N_VGND_M1001_s N_VGND_M1004_s N_VGND_M1013_s
+ N_VGND_M1016_s N_VGND_M1023_s N_VGND_c_807_n N_VGND_c_808_n N_VGND_c_809_n
+ N_VGND_c_810_n N_VGND_c_811_n N_VGND_c_812_n N_VGND_c_813_n N_VGND_c_814_n
+ N_VGND_c_815_n N_VGND_c_816_n N_VGND_c_817_n VGND N_VGND_c_818_n
+ N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n PM_SKY130_FD_SC_LP__INVLP_8%VGND
x_PM_SKY130_FD_SC_LP__INVLP_8%A_114_53# N_A_114_53#_M1001_d N_A_114_53#_M1011_d
+ N_A_114_53#_M1015_d N_A_114_53#_M1022_d N_A_114_53#_M1002_s
+ N_A_114_53#_M1009_s N_A_114_53#_M1025_s N_A_114_53#_M1027_s
+ N_A_114_53#_c_922_n N_A_114_53#_c_923_n N_A_114_53#_c_939_n
+ N_A_114_53#_c_924_n N_A_114_53#_c_944_n N_A_114_53#_c_925_n
+ N_A_114_53#_c_948_n N_A_114_53#_c_926_n N_A_114_53#_c_927_n
+ N_A_114_53#_c_953_n N_A_114_53#_c_928_n N_A_114_53#_c_993_n
+ N_A_114_53#_c_929_n N_A_114_53#_c_930_n N_A_114_53#_c_963_n
+ N_A_114_53#_c_1001_n N_A_114_53#_c_1002_n N_A_114_53#_c_931_n
+ N_A_114_53#_c_932_n N_A_114_53#_c_933_n N_A_114_53#_c_934_n
+ PM_SKY130_FD_SC_LP__INVLP_8%A_114_53#
cc_1 VNB N_A_M1001_g 0.0316821f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.685
cc_2 VNB N_A_M1004_g 0.021659f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.685
cc_3 VNB N_A_M1011_g 0.0220136f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.685
cc_4 VNB N_A_M1013_g 0.0220539f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.685
cc_5 VNB N_A_M1015_g 0.0220752f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.685
cc_6 VNB N_A_M1016_g 0.0220752f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.685
cc_7 VNB N_A_M1022_g 0.022076f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=0.685
cc_8 VNB N_A_M1000_g 0.0222364f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=0.685
cc_9 VNB N_A_M1002_g 0.0222372f $X=-0.19 $Y=-0.245 $X2=3.935 $Y2=0.685
cc_10 VNB N_A_M1007_g 0.0222372f $X=-0.19 $Y=-0.245 $X2=4.365 $Y2=0.685
cc_11 VNB N_A_M1009_g 0.0222372f $X=-0.19 $Y=-0.245 $X2=4.795 $Y2=0.685
cc_12 VNB N_A_M1014_g 0.0222372f $X=-0.19 $Y=-0.245 $X2=5.225 $Y2=0.685
cc_13 VNB N_A_M1025_g 0.0232397f $X=-0.19 $Y=-0.245 $X2=5.655 $Y2=0.685
cc_14 VNB N_A_M1026_g 0.0242421f $X=-0.19 $Y=-0.245 $X2=6.155 $Y2=0.685
cc_15 VNB N_A_M1027_g 0.0245555f $X=-0.19 $Y=-0.245 $X2=6.655 $Y2=0.685
cc_16 VNB N_A_M1023_g 0.0327026f $X=-0.19 $Y=-0.245 $X2=7.155 $Y2=0.685
cc_17 VNB N_A_c_112_n 0.0125848f $X=-0.19 $Y=-0.245 $X2=7.25 $Y2=1.51
cc_18 VNB N_A_c_113_n 0.306282f $X=-0.19 $Y=-0.245 $X2=7.25 $Y2=1.51
cc_19 VNB N_A_c_114_n 0.00139588f $X=-0.19 $Y=-0.245 $X2=2 $Y2=1.562
cc_20 VNB N_VPWR_c_408_n 0.322901f $X=-0.19 $Y=-0.245 $X2=4.365 $Y2=0.685
cc_21 VNB N_Y_c_632_n 0.00159633f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.685
cc_22 VNB N_Y_c_633_n 0.0148755f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.675
cc_23 VNB N_Y_c_634_n 0.00324651f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.345
cc_24 VNB N_Y_c_635_n 0.00225436f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=0.685
cc_25 VNB N_Y_c_636_n 0.00537496f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.675
cc_26 VNB N_Y_c_637_n 0.00177357f $X=-0.19 $Y=-0.245 $X2=4.365 $Y2=1.345
cc_27 VNB N_Y_c_638_n 0.00177357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_639_n 0.00229801f $X=-0.19 $Y=-0.245 $X2=4.505 $Y2=2.465
cc_29 VNB N_VGND_c_807_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_808_n 0.0479102f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.685
cc_31 VNB N_VGND_c_809_n 8.31601e-19 $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=2.465
cc_32 VNB N_VGND_c_810_n 7.97178e-19 $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.685
cc_33 VNB N_VGND_c_811_n 0.00102933f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=2.465
cc_34 VNB N_VGND_c_812_n 0.011635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_813_n 0.0441817f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.685
cc_36 VNB N_VGND_c_814_n 0.011999f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.675
cc_37 VNB N_VGND_c_815_n 0.00472949f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=2.465
cc_38 VNB N_VGND_c_816_n 0.011999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_817_n 0.00472949f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.345
cc_40 VNB N_VGND_c_818_n 0.0152756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_819_n 0.0960093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_820_n 0.00472949f $X=-0.19 $Y=-0.245 $X2=3.935 $Y2=0.685
cc_43 VNB N_VGND_c_821_n 0.400508f $X=-0.19 $Y=-0.245 $X2=4.075 $Y2=2.465
cc_44 VNB N_A_114_53#_c_922_n 0.00170023f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.685
cc_45 VNB N_A_114_53#_c_923_n 0.00366139f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=2.465
cc_46 VNB N_A_114_53#_c_924_n 0.0013877f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.675
cc_47 VNB N_A_114_53#_c_925_n 0.0013877f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.685
cc_48 VNB N_A_114_53#_c_926_n 0.00237811f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=0.685
cc_49 VNB N_A_114_53#_c_927_n 0.00130493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_114_53#_c_928_n 0.00237811f $X=-0.19 $Y=-0.245 $X2=3.505 $Y2=1.345
cc_51 VNB N_A_114_53#_c_929_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=2.465
cc_52 VNB N_A_114_53#_c_930_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=3.935 $Y2=0.685
cc_53 VNB N_A_114_53#_c_931_n 0.00203277f $X=-0.19 $Y=-0.245 $X2=4.365 $Y2=0.685
cc_54 VNB N_A_114_53#_c_932_n 0.00121966f $X=-0.19 $Y=-0.245 $X2=4.365 $Y2=0.685
cc_55 VNB N_A_114_53#_c_933_n 0.00220701f $X=-0.19 $Y=-0.245 $X2=4.505 $Y2=1.675
cc_56 VNB N_A_114_53#_c_934_n 0.0049581f $X=-0.19 $Y=-0.245 $X2=4.505 $Y2=2.465
cc_57 VPB N_A_M1003_g 0.0255339f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_58 VPB N_A_M1006_g 0.0174225f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_59 VPB N_A_M1010_g 0.0184795f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=2.465
cc_60 VPB N_A_M1017_g 0.0176783f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=2.465
cc_61 VPB N_A_M1020_g 0.017887f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=2.465
cc_62 VPB N_A_M1021_g 0.0193454f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.465
cc_63 VPB N_A_M1028_g 0.019776f $X=-0.19 $Y=1.655 $X2=3.215 $Y2=2.465
cc_64 VPB N_A_M1005_g 0.0187367f $X=-0.19 $Y=1.655 $X2=3.645 $Y2=2.465
cc_65 VPB N_A_M1008_g 0.0187483f $X=-0.19 $Y=1.655 $X2=4.075 $Y2=2.465
cc_66 VPB N_A_M1012_g 0.0187483f $X=-0.19 $Y=1.655 $X2=4.505 $Y2=2.465
cc_67 VPB N_A_M1018_g 0.0187483f $X=-0.19 $Y=1.655 $X2=4.935 $Y2=2.465
cc_68 VPB N_A_M1019_g 0.0187483f $X=-0.19 $Y=1.655 $X2=5.365 $Y2=2.465
cc_69 VPB N_A_M1024_g 0.0187483f $X=-0.19 $Y=1.655 $X2=5.795 $Y2=2.465
cc_70 VPB N_A_M1030_g 0.0195411f $X=-0.19 $Y=1.655 $X2=6.225 $Y2=2.465
cc_71 VPB N_A_M1031_g 0.0195411f $X=-0.19 $Y=1.655 $X2=6.725 $Y2=2.465
cc_72 VPB N_A_M1029_g 0.0252388f $X=-0.19 $Y=1.655 $X2=7.155 $Y2=2.465
cc_73 VPB N_A_c_112_n 7.73822e-19 $X=-0.19 $Y=1.655 $X2=7.25 $Y2=1.51
cc_74 VPB N_A_c_113_n 0.067013f $X=-0.19 $Y=1.655 $X2=7.25 $Y2=1.51
cc_75 VPB N_A_c_133_n 0.00668504f $X=-0.19 $Y=1.655 $X2=3.018 $Y2=1.562
cc_76 VPB N_A_c_114_n 0.00404148f $X=-0.19 $Y=1.655 $X2=2 $Y2=1.562
cc_77 VPB N_A_c_135_n 0.00113907f $X=-0.19 $Y=1.655 $X2=3.235 $Y2=1.562
cc_78 VPB N_VPWR_c_409_n 0.0106521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_410_n 0.0618081f $X=-0.19 $Y=1.655 $X2=1.355 $Y2=0.685
cc_80 VPB N_VPWR_c_411_n 3.22457e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_412_n 0.00229788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_413_n 0.00552394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_414_n 0.0119347f $X=-0.19 $Y=1.655 $X2=2.215 $Y2=0.685
cc_84 VPB N_VPWR_c_415_n 0.0508336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_416_n 0.0131279f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=1.345
cc_86 VPB N_VPWR_c_417_n 0.00356964f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=0.685
cc_87 VPB N_VPWR_c_418_n 0.0182639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_419_n 0.00631455f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=1.675
cc_89 VPB N_VPWR_c_420_n 0.0158404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_421_n 0.0930962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_422_n 0.00436868f $X=-0.19 $Y=1.655 $X2=4.075 $Y2=2.465
cc_92 VPB N_VPWR_c_408_n 0.0470032f $X=-0.19 $Y=1.655 $X2=4.365 $Y2=0.685
cc_93 VPB N_Y_c_640_n 5.1007e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_Y_c_641_n 0.00363384f $X=-0.19 $Y=1.655 $X2=4.075 $Y2=2.465
cc_95 VPB N_Y_c_642_n 8.75554e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 N_A_M1003_g N_VPWR_c_410_n 0.0073203f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A_M1003_g N_VPWR_c_411_n 6.19298e-19 $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_M1006_g N_VPWR_c_411_n 0.0100242f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_M1010_g N_VPWR_c_411_n 0.0098444f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_M1017_g N_VPWR_c_411_n 5.82718e-19 $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A_M1010_g N_VPWR_c_412_n 5.77413e-19 $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_M1017_g N_VPWR_c_412_n 0.00925199f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A_M1020_g N_VPWR_c_412_n 0.00313805f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A_M1021_g N_VPWR_c_413_n 0.00598313f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A_M1028_g N_VPWR_c_413_n 0.00598313f $X=3.215 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A_M1031_g N_VPWR_c_415_n 0.00109254f $X=6.725 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_M1029_g N_VPWR_c_415_n 0.0225088f $X=7.155 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_c_112_n N_VPWR_c_415_n 0.0145929f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A_c_113_n N_VPWR_c_415_n 0.00413601f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_110 N_A_M1010_g N_VPWR_c_416_n 0.00486043f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_M1017_g N_VPWR_c_416_n 0.00486043f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_M1020_g N_VPWR_c_418_n 0.0054895f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_M1021_g N_VPWR_c_418_n 0.0054895f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A_M1003_g N_VPWR_c_420_n 0.0054895f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_M1006_g N_VPWR_c_420_n 0.00486043f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_M1028_g N_VPWR_c_421_n 0.00547432f $X=3.215 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_M1005_g N_VPWR_c_421_n 0.00357842f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_M1008_g N_VPWR_c_421_n 0.00357842f $X=4.075 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_M1012_g N_VPWR_c_421_n 0.00357842f $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A_M1018_g N_VPWR_c_421_n 0.00357842f $X=4.935 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_M1019_g N_VPWR_c_421_n 0.00357842f $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_M1024_g N_VPWR_c_421_n 0.00357842f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_M1030_g N_VPWR_c_421_n 0.00357842f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_M1031_g N_VPWR_c_421_n 0.00357877f $X=6.725 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_M1029_g N_VPWR_c_421_n 0.00486043f $X=7.155 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_M1003_g N_VPWR_c_408_n 0.010744f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_M1006_g N_VPWR_c_408_n 0.00824727f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_M1010_g N_VPWR_c_408_n 0.00824727f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A_M1017_g N_VPWR_c_408_n 0.00824727f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A_M1020_g N_VPWR_c_408_n 0.00990036f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A_M1021_g N_VPWR_c_408_n 0.0102184f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A_M1028_g N_VPWR_c_408_n 0.0101814f $X=3.215 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A_M1005_g N_VPWR_c_408_n 0.00535118f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A_M1008_g N_VPWR_c_408_n 0.00535118f $X=4.075 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_M1012_g N_VPWR_c_408_n 0.00535118f $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_M1018_g N_VPWR_c_408_n 0.00535118f $X=4.935 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_M1019_g N_VPWR_c_408_n 0.00535118f $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A_M1024_g N_VPWR_c_408_n 0.00535118f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_M1030_g N_VPWR_c_408_n 0.00553547f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A_M1031_g N_VPWR_c_408_n 0.00553549f $X=6.725 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_M1029_g N_VPWR_c_408_n 0.00824727f $X=7.155 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_M1003_g N_A_114_367#_c_518_n 0.00489293f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_c_113_n N_A_114_367#_c_518_n 6.09546e-19 $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A_M1003_g N_A_114_367#_c_520_n 0.00698794f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_M1006_g N_A_114_367#_c_521_n 0.0135977f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_M1010_g N_A_114_367#_c_521_n 0.0122595f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_M1017_g N_A_114_367#_c_523_n 0.0122595f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_M1020_g N_A_114_367#_c_523_n 0.01115f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_M1021_g N_A_114_367#_c_525_n 0.0118691f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_M1028_g N_A_114_367#_c_525_n 0.0118691f $X=3.215 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_M1028_g N_A_114_367#_c_527_n 7.32094e-19 $X=3.215 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_M1005_g N_A_114_367#_c_527_n 0.0021125f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_M1021_g N_A_114_367#_c_529_n 5.85908e-19 $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_154 N_A_M1028_g N_A_114_367#_c_529_n 0.00704975f $X=3.215 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_M1005_g N_A_114_367#_c_529_n 0.00656286f $X=3.645 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_M1008_g N_A_114_367#_c_529_n 5.16617e-19 $X=4.075 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_M1005_g N_A_114_367#_c_533_n 0.0105205f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_M1008_g N_A_114_367#_c_533_n 0.0105205f $X=4.075 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A_M1028_g N_A_114_367#_c_535_n 0.00196648f $X=3.215 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_M1005_g N_A_114_367#_c_535_n 5.89773e-19 $X=3.645 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_M1005_g N_A_114_367#_c_537_n 5.9898e-19 $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A_M1008_g N_A_114_367#_c_537_n 0.0110126f $X=4.075 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_M1012_g N_A_114_367#_c_537_n 0.0110126f $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A_M1018_g N_A_114_367#_c_537_n 5.9898e-19 $X=4.935 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_M1012_g N_A_114_367#_c_541_n 0.0105205f $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A_M1018_g N_A_114_367#_c_541_n 0.0105205f $X=4.935 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A_M1012_g N_A_114_367#_c_543_n 5.9898e-19 $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A_M1018_g N_A_114_367#_c_543_n 0.0110126f $X=4.935 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A_M1019_g N_A_114_367#_c_543_n 0.0110126f $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_M1024_g N_A_114_367#_c_543_n 5.9898e-19 $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A_M1019_g N_A_114_367#_c_547_n 0.0105205f $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A_M1024_g N_A_114_367#_c_547_n 0.0105205f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A_M1019_g N_A_114_367#_c_549_n 5.9898e-19 $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_M1024_g N_A_114_367#_c_549_n 0.0119757f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A_M1030_g N_A_114_367#_c_549_n 0.0122249f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_M1031_g N_A_114_367#_c_549_n 9.39294e-19 $X=6.725 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_M1030_g N_A_114_367#_c_553_n 0.0109138f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_M1031_g N_A_114_367#_c_553_n 0.0118963f $X=6.725 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A_c_112_n N_A_114_367#_c_555_n 0.0137839f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A_c_113_n N_A_114_367#_c_555_n 0.00232957f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_181 N_A_M1003_g N_A_114_367#_c_557_n 0.00192234f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_M1017_g N_A_114_367#_c_558_n 6.73728e-19 $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_M1020_g N_A_114_367#_c_558_n 0.00947025f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_184 N_A_M1021_g N_A_114_367#_c_558_n 0.0097425f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_M1028_g N_A_114_367#_c_558_n 6.19919e-19 $X=3.215 $Y=2.465 $X2=0
+ $Y2=0
cc_186 N_A_M1008_g N_A_114_367#_c_562_n 5.89773e-19 $X=4.075 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_M1012_g N_A_114_367#_c_562_n 5.89773e-19 $X=4.505 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_M1018_g N_A_114_367#_c_564_n 5.89773e-19 $X=4.935 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_A_M1019_g N_A_114_367#_c_564_n 5.89773e-19 $X=5.365 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A_M1024_g N_A_114_367#_c_566_n 5.89773e-19 $X=5.795 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A_M1030_g N_A_114_367#_c_566_n 5.89773e-19 $X=6.225 $Y=2.465 $X2=0
+ $Y2=0
cc_192 N_A_M1001_g N_Y_c_632_n 8.44792e-19 $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_193 N_A_M1004_g N_Y_c_632_n 0.00419028f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_194 N_A_M1011_g N_Y_c_632_n 0.00360365f $X=1.355 $Y=0.685 $X2=0 $Y2=0
cc_195 N_A_c_113_n N_Y_c_632_n 0.0155104f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A_c_114_n N_Y_c_632_n 0.0155819f $X=2 $Y=1.562 $X2=0 $Y2=0
cc_197 N_A_M1003_g N_Y_c_640_n 5.2502e-19 $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A_M1006_g N_Y_c_640_n 0.00437719f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A_M1010_g N_Y_c_640_n 0.00358934f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A_M1011_g N_Y_c_633_n 0.0112067f $X=1.355 $Y=0.685 $X2=0 $Y2=0
cc_201 N_A_M1013_g N_Y_c_633_n 0.0104864f $X=1.785 $Y=0.685 $X2=0 $Y2=0
cc_202 N_A_M1015_g N_Y_c_633_n 0.0104926f $X=2.215 $Y=0.685 $X2=0 $Y2=0
cc_203 N_A_M1016_g N_Y_c_633_n 0.0104926f $X=2.645 $Y=0.685 $X2=0 $Y2=0
cc_204 N_A_M1022_g N_Y_c_633_n 0.0104926f $X=3.075 $Y=0.685 $X2=0 $Y2=0
cc_205 N_A_M1000_g N_Y_c_633_n 0.00899033f $X=3.505 $Y=0.685 $X2=0 $Y2=0
cc_206 N_A_c_113_n N_Y_c_633_n 0.0113474f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_207 N_A_c_133_n N_Y_c_633_n 0.116577f $X=3.018 $Y=1.562 $X2=0 $Y2=0
cc_208 N_A_c_114_n N_Y_c_633_n 0.0521718f $X=2 $Y=1.562 $X2=0 $Y2=0
cc_209 N_A_M1001_g N_Y_c_660_n 2.89663e-19 $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_210 N_A_M1004_g N_Y_c_660_n 0.00487892f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_211 N_A_M1010_g N_Y_c_662_n 0.011757f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A_M1017_g N_Y_c_662_n 0.0104864f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A_M1020_g N_Y_c_662_n 0.0104915f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A_M1021_g N_Y_c_662_n 0.0112106f $X=2.645 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A_M1028_g N_Y_c_662_n 0.0114042f $X=3.215 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A_M1005_g N_Y_c_662_n 0.0128314f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_c_112_n N_Y_c_662_n 0.0227098f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_218 N_A_c_113_n N_Y_c_662_n 0.00724546f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_219 N_A_c_133_n N_Y_c_662_n 0.0853812f $X=3.018 $Y=1.562 $X2=0 $Y2=0
cc_220 N_A_c_114_n N_Y_c_662_n 0.0412355f $X=2 $Y=1.562 $X2=0 $Y2=0
cc_221 N_A_M1006_g N_Y_c_672_n 0.0043809f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A_M1022_g N_Y_c_673_n 9.24842e-19 $X=3.075 $Y=0.685 $X2=0 $Y2=0
cc_223 N_A_M1000_g N_Y_c_673_n 0.00644131f $X=3.505 $Y=0.685 $X2=0 $Y2=0
cc_224 N_A_M1002_g N_Y_c_634_n 0.0115018f $X=3.935 $Y=0.685 $X2=0 $Y2=0
cc_225 N_A_M1007_g N_Y_c_634_n 0.0115018f $X=4.365 $Y=0.685 $X2=0 $Y2=0
cc_226 N_A_c_112_n N_Y_c_634_n 0.0506643f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_227 N_A_c_113_n N_Y_c_634_n 0.00263605f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A_M1008_g N_Y_c_679_n 0.0122595f $X=4.075 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A_M1012_g N_Y_c_679_n 0.0122306f $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A_c_112_n N_Y_c_679_n 0.0420181f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_231 N_A_c_113_n N_Y_c_679_n 0.00263605f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_232 N_A_M1009_g N_Y_c_683_n 0.00640964f $X=4.795 $Y=0.685 $X2=0 $Y2=0
cc_233 N_A_M1014_g N_Y_c_683_n 5.72721e-19 $X=5.225 $Y=0.685 $X2=0 $Y2=0
cc_234 N_A_M1009_g N_Y_c_635_n 0.00899033f $X=4.795 $Y=0.685 $X2=0 $Y2=0
cc_235 N_A_M1014_g N_Y_c_635_n 0.00899033f $X=5.225 $Y=0.685 $X2=0 $Y2=0
cc_236 N_A_c_112_n N_Y_c_635_n 0.0388321f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_237 N_A_c_113_n N_Y_c_635_n 0.00263605f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_238 N_A_M1018_g N_Y_c_689_n 0.0122595f $X=4.935 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A_M1019_g N_Y_c_689_n 0.0122595f $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_c_112_n N_Y_c_689_n 0.0420181f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_241 N_A_c_113_n N_Y_c_689_n 0.00263605f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_242 N_A_M1009_g N_Y_c_693_n 5.71288e-19 $X=4.795 $Y=0.685 $X2=0 $Y2=0
cc_243 N_A_M1014_g N_Y_c_693_n 0.00661193f $X=5.225 $Y=0.685 $X2=0 $Y2=0
cc_244 N_A_M1025_g N_Y_c_693_n 0.00701103f $X=5.655 $Y=0.685 $X2=0 $Y2=0
cc_245 N_A_M1026_g N_Y_c_693_n 2.75259e-19 $X=6.155 $Y=0.685 $X2=0 $Y2=0
cc_246 N_A_M1025_g N_Y_c_636_n 0.00938357f $X=5.655 $Y=0.685 $X2=0 $Y2=0
cc_247 N_A_M1026_g N_Y_c_636_n 0.012905f $X=6.155 $Y=0.685 $X2=0 $Y2=0
cc_248 N_A_M1027_g N_Y_c_636_n 0.00492244f $X=6.655 $Y=0.685 $X2=0 $Y2=0
cc_249 N_A_M1023_g N_Y_c_636_n 2.71338e-19 $X=7.155 $Y=0.685 $X2=0 $Y2=0
cc_250 N_A_c_112_n N_Y_c_636_n 0.0766181f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_251 N_A_c_113_n N_Y_c_636_n 0.00857451f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_252 N_A_M1024_g N_Y_c_703_n 0.0122595f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_253 N_A_M1030_g N_Y_c_703_n 0.014733f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_254 N_A_c_112_n N_Y_c_703_n 0.0416768f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_255 N_A_c_113_n N_Y_c_703_n 0.00251785f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_256 N_A_M1027_g N_Y_c_707_n 0.00488246f $X=6.655 $Y=0.685 $X2=0 $Y2=0
cc_257 N_A_M1003_g N_Y_c_641_n 0.00317194f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A_M1006_g N_Y_c_641_n 0.00497313f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A_c_113_n N_Y_c_641_n 0.0228188f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_260 N_A_M1006_g N_Y_c_642_n 0.00107549f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A_M1010_g N_Y_c_642_n 0.00107962f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A_c_113_n N_Y_c_642_n 0.00476357f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_263 N_A_c_114_n N_Y_c_642_n 0.0154195f $X=2 $Y=1.562 $X2=0 $Y2=0
cc_264 N_A_M1000_g N_Y_c_637_n 0.0021743f $X=3.505 $Y=0.685 $X2=0 $Y2=0
cc_265 N_A_c_112_n N_Y_c_637_n 0.020702f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_266 N_A_c_113_n N_Y_c_637_n 0.00270932f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_267 N_A_c_112_n N_Y_c_718_n 0.0138593f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_268 N_A_c_113_n N_Y_c_718_n 0.00272398f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_269 N_A_M1009_g N_Y_c_638_n 0.0021743f $X=4.795 $Y=0.685 $X2=0 $Y2=0
cc_270 N_A_c_112_n N_Y_c_638_n 0.020702f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_271 N_A_c_113_n N_Y_c_638_n 0.00270932f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_272 N_A_c_112_n N_Y_c_723_n 0.0138593f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_273 N_A_c_113_n N_Y_c_723_n 0.00272398f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_274 N_A_M1014_g N_Y_c_639_n 0.0021743f $X=5.225 $Y=0.685 $X2=0 $Y2=0
cc_275 N_A_M1025_g N_Y_c_639_n 0.0021743f $X=5.655 $Y=0.685 $X2=0 $Y2=0
cc_276 N_A_c_112_n N_Y_c_639_n 0.0272511f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_277 N_A_c_113_n N_Y_c_639_n 0.00270932f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_278 N_A_c_112_n N_Y_c_729_n 0.0138593f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_279 N_A_c_113_n N_Y_c_729_n 0.00272398f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_280 N_A_M1031_g N_Y_c_731_n 0.011928f $X=6.725 $Y=2.465 $X2=0 $Y2=0
cc_281 N_A_c_112_n N_Y_c_731_n 0.024044f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_282 N_A_c_113_n N_Y_c_731_n 0.00423635f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_283 N_A_M1001_g N_VGND_c_808_n 0.0066302f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_284 N_A_M1001_g N_VGND_c_809_n 4.89794e-19 $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_285 N_A_M1004_g N_VGND_c_809_n 0.00656226f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_286 N_A_M1011_g N_VGND_c_809_n 0.00641832f $X=1.355 $Y=0.685 $X2=0 $Y2=0
cc_287 N_A_M1013_g N_VGND_c_809_n 4.59873e-19 $X=1.785 $Y=0.685 $X2=0 $Y2=0
cc_288 N_A_M1011_g N_VGND_c_810_n 4.59873e-19 $X=1.355 $Y=0.685 $X2=0 $Y2=0
cc_289 N_A_M1013_g N_VGND_c_810_n 0.00641832f $X=1.785 $Y=0.685 $X2=0 $Y2=0
cc_290 N_A_M1015_g N_VGND_c_810_n 0.00641832f $X=2.215 $Y=0.685 $X2=0 $Y2=0
cc_291 N_A_M1016_g N_VGND_c_810_n 4.59873e-19 $X=2.645 $Y=0.685 $X2=0 $Y2=0
cc_292 N_A_M1015_g N_VGND_c_811_n 4.59873e-19 $X=2.215 $Y=0.685 $X2=0 $Y2=0
cc_293 N_A_M1016_g N_VGND_c_811_n 0.00641832f $X=2.645 $Y=0.685 $X2=0 $Y2=0
cc_294 N_A_M1022_g N_VGND_c_811_n 0.00733695f $X=3.075 $Y=0.685 $X2=0 $Y2=0
cc_295 N_A_M1000_g N_VGND_c_811_n 9.92089e-19 $X=3.505 $Y=0.685 $X2=0 $Y2=0
cc_296 N_A_M1023_g N_VGND_c_813_n 0.00787605f $X=7.155 $Y=0.685 $X2=0 $Y2=0
cc_297 N_A_c_112_n N_VGND_c_813_n 0.00897005f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_298 N_A_c_113_n N_VGND_c_813_n 0.00292725f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_299 N_A_M1011_g N_VGND_c_814_n 0.00336564f $X=1.355 $Y=0.685 $X2=0 $Y2=0
cc_300 N_A_M1013_g N_VGND_c_814_n 0.00336564f $X=1.785 $Y=0.685 $X2=0 $Y2=0
cc_301 N_A_M1015_g N_VGND_c_816_n 0.00336564f $X=2.215 $Y=0.685 $X2=0 $Y2=0
cc_302 N_A_M1016_g N_VGND_c_816_n 0.00336564f $X=2.645 $Y=0.685 $X2=0 $Y2=0
cc_303 N_A_M1001_g N_VGND_c_818_n 0.00520505f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_304 N_A_M1004_g N_VGND_c_818_n 0.00336564f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_305 N_A_M1022_g N_VGND_c_819_n 0.00336564f $X=3.075 $Y=0.685 $X2=0 $Y2=0
cc_306 N_A_M1000_g N_VGND_c_819_n 0.00338313f $X=3.505 $Y=0.685 $X2=0 $Y2=0
cc_307 N_A_M1002_g N_VGND_c_819_n 0.0033828f $X=3.935 $Y=0.685 $X2=0 $Y2=0
cc_308 N_A_M1007_g N_VGND_c_819_n 0.0033828f $X=4.365 $Y=0.685 $X2=0 $Y2=0
cc_309 N_A_M1009_g N_VGND_c_819_n 0.00338313f $X=4.795 $Y=0.685 $X2=0 $Y2=0
cc_310 N_A_M1014_g N_VGND_c_819_n 0.00338313f $X=5.225 $Y=0.685 $X2=0 $Y2=0
cc_311 N_A_M1025_g N_VGND_c_819_n 0.00338313f $X=5.655 $Y=0.685 $X2=0 $Y2=0
cc_312 N_A_M1026_g N_VGND_c_819_n 0.0033828f $X=6.155 $Y=0.685 $X2=0 $Y2=0
cc_313 N_A_M1027_g N_VGND_c_819_n 0.00338313f $X=6.655 $Y=0.685 $X2=0 $Y2=0
cc_314 N_A_M1023_g N_VGND_c_819_n 0.00519058f $X=7.155 $Y=0.685 $X2=0 $Y2=0
cc_315 N_A_M1001_g N_VGND_c_821_n 0.0104451f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_316 N_A_M1004_g N_VGND_c_821_n 0.00409996f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_317 N_A_M1011_g N_VGND_c_821_n 0.00409996f $X=1.355 $Y=0.685 $X2=0 $Y2=0
cc_318 N_A_M1013_g N_VGND_c_821_n 0.00409996f $X=1.785 $Y=0.685 $X2=0 $Y2=0
cc_319 N_A_M1015_g N_VGND_c_821_n 0.00409996f $X=2.215 $Y=0.685 $X2=0 $Y2=0
cc_320 N_A_M1016_g N_VGND_c_821_n 0.00409996f $X=2.645 $Y=0.685 $X2=0 $Y2=0
cc_321 N_A_M1022_g N_VGND_c_821_n 0.00409996f $X=3.075 $Y=0.685 $X2=0 $Y2=0
cc_322 N_A_M1000_g N_VGND_c_821_n 0.00509124f $X=3.505 $Y=0.685 $X2=0 $Y2=0
cc_323 N_A_M1002_g N_VGND_c_821_n 0.00509122f $X=3.935 $Y=0.685 $X2=0 $Y2=0
cc_324 N_A_M1007_g N_VGND_c_821_n 0.00509122f $X=4.365 $Y=0.685 $X2=0 $Y2=0
cc_325 N_A_M1009_g N_VGND_c_821_n 0.00509124f $X=4.795 $Y=0.685 $X2=0 $Y2=0
cc_326 N_A_M1014_g N_VGND_c_821_n 0.00509124f $X=5.225 $Y=0.685 $X2=0 $Y2=0
cc_327 N_A_M1025_g N_VGND_c_821_n 0.00523603f $X=5.655 $Y=0.685 $X2=0 $Y2=0
cc_328 N_A_M1026_g N_VGND_c_821_n 0.00538081f $X=6.155 $Y=0.685 $X2=0 $Y2=0
cc_329 N_A_M1027_g N_VGND_c_821_n 0.00538083f $X=6.655 $Y=0.685 $X2=0 $Y2=0
cc_330 N_A_M1023_g N_VGND_c_821_n 0.0105745f $X=7.155 $Y=0.685 $X2=0 $Y2=0
cc_331 N_A_M1001_g N_A_114_53#_c_922_n 0.00518192f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_332 N_A_M1004_g N_A_114_53#_c_922_n 2.81313e-19 $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_333 N_A_M1001_g N_A_114_53#_c_923_n 0.0045732f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_334 N_A_c_113_n N_A_114_53#_c_923_n 0.00254615f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_335 N_A_M1004_g N_A_114_53#_c_939_n 0.0143358f $X=0.925 $Y=0.685 $X2=0 $Y2=0
cc_336 N_A_M1011_g N_A_114_53#_c_939_n 0.0107718f $X=1.355 $Y=0.685 $X2=0 $Y2=0
cc_337 N_A_c_113_n N_A_114_53#_c_939_n 2.2967e-19 $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_338 N_A_M1011_g N_A_114_53#_c_924_n 4.26168e-19 $X=1.355 $Y=0.685 $X2=0 $Y2=0
cc_339 N_A_M1013_g N_A_114_53#_c_924_n 4.26168e-19 $X=1.785 $Y=0.685 $X2=0 $Y2=0
cc_340 N_A_M1013_g N_A_114_53#_c_944_n 0.0107855f $X=1.785 $Y=0.685 $X2=0 $Y2=0
cc_341 N_A_M1015_g N_A_114_53#_c_944_n 0.0107855f $X=2.215 $Y=0.685 $X2=0 $Y2=0
cc_342 N_A_M1015_g N_A_114_53#_c_925_n 4.26168e-19 $X=2.215 $Y=0.685 $X2=0 $Y2=0
cc_343 N_A_M1016_g N_A_114_53#_c_925_n 4.26168e-19 $X=2.645 $Y=0.685 $X2=0 $Y2=0
cc_344 N_A_M1016_g N_A_114_53#_c_948_n 0.0107389f $X=2.645 $Y=0.685 $X2=0 $Y2=0
cc_345 N_A_M1022_g N_A_114_53#_c_948_n 0.0105157f $X=3.075 $Y=0.685 $X2=0 $Y2=0
cc_346 N_A_M1000_g N_A_114_53#_c_926_n 0.0100634f $X=3.505 $Y=0.685 $X2=0 $Y2=0
cc_347 N_A_M1002_g N_A_114_53#_c_926_n 0.00822656f $X=3.935 $Y=0.685 $X2=0 $Y2=0
cc_348 N_A_M1022_g N_A_114_53#_c_927_n 4.37262e-19 $X=3.075 $Y=0.685 $X2=0 $Y2=0
cc_349 N_A_M1000_g N_A_114_53#_c_953_n 6.19364e-19 $X=3.505 $Y=0.685 $X2=0 $Y2=0
cc_350 N_A_M1002_g N_A_114_53#_c_953_n 0.00712923f $X=3.935 $Y=0.685 $X2=0 $Y2=0
cc_351 N_A_M1007_g N_A_114_53#_c_953_n 0.00712923f $X=4.365 $Y=0.685 $X2=0 $Y2=0
cc_352 N_A_M1009_g N_A_114_53#_c_953_n 6.19364e-19 $X=4.795 $Y=0.685 $X2=0 $Y2=0
cc_353 N_A_M1007_g N_A_114_53#_c_928_n 0.00827312f $X=4.365 $Y=0.685 $X2=0 $Y2=0
cc_354 N_A_M1009_g N_A_114_53#_c_928_n 0.0103332f $X=4.795 $Y=0.685 $X2=0 $Y2=0
cc_355 N_A_M1014_g N_A_114_53#_c_929_n 0.0103332f $X=5.225 $Y=0.685 $X2=0 $Y2=0
cc_356 N_A_M1025_g N_A_114_53#_c_929_n 0.0116441f $X=5.655 $Y=0.685 $X2=0 $Y2=0
cc_357 N_A_M1026_g N_A_114_53#_c_930_n 0.00866637f $X=6.155 $Y=0.685 $X2=0 $Y2=0
cc_358 N_A_M1027_g N_A_114_53#_c_930_n 0.0142587f $X=6.655 $Y=0.685 $X2=0 $Y2=0
cc_359 N_A_M1001_g N_A_114_53#_c_963_n 0.00306596f $X=0.495 $Y=0.685 $X2=0 $Y2=0
cc_360 N_A_M1002_g N_A_114_53#_c_931_n 0.00171638f $X=3.935 $Y=0.685 $X2=0 $Y2=0
cc_361 N_A_M1007_g N_A_114_53#_c_931_n 0.00171638f $X=4.365 $Y=0.685 $X2=0 $Y2=0
cc_362 N_A_M1026_g N_A_114_53#_c_933_n 0.00686149f $X=6.155 $Y=0.685 $X2=0 $Y2=0
cc_363 N_A_M1027_g N_A_114_53#_c_933_n 6.03526e-19 $X=6.655 $Y=0.685 $X2=0 $Y2=0
cc_364 N_A_M1027_g N_A_114_53#_c_934_n 0.00371159f $X=6.655 $Y=0.685 $X2=0 $Y2=0
cc_365 N_A_M1023_g N_A_114_53#_c_934_n 0.0122586f $X=7.155 $Y=0.685 $X2=0 $Y2=0
cc_366 N_A_c_112_n N_A_114_53#_c_934_n 0.022699f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_367 N_A_c_113_n N_A_114_53#_c_934_n 0.00411924f $X=7.25 $Y=1.51 $X2=0 $Y2=0
cc_368 N_VPWR_c_408_n N_A_114_367#_M1003_s 0.0041489f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_369 N_VPWR_c_408_n N_A_114_367#_M1010_s 0.00606222f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_408_n N_A_114_367#_M1020_s 0.00223559f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_408_n N_A_114_367#_M1028_s 0.00223559f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_372 N_VPWR_c_408_n N_A_114_367#_M1008_s 0.00223559f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_408_n N_A_114_367#_M1018_s 0.00223559f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_408_n N_A_114_367#_M1024_s 0.00223559f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_408_n N_A_114_367#_M1031_s 0.00411415f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_420_n N_A_114_367#_c_520_n 0.0153332f $X=0.975 $Y=3.33 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_408_n N_A_114_367#_c_520_n 0.00945339f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_378 N_VPWR_M1006_d N_A_114_367#_c_521_n 0.0034343f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_379 N_VPWR_c_411_n N_A_114_367#_c_521_n 0.0171619f $X=1.14 $Y=2.87 $X2=0
+ $Y2=0
cc_380 N_VPWR_M1017_d N_A_114_367#_c_523_n 0.00344593f $X=1.86 $Y=1.835 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_412_n N_A_114_367#_c_523_n 0.0153337f $X=2 $Y=2.87 $X2=0 $Y2=0
cc_382 N_VPWR_M1021_d N_A_114_367#_c_525_n 0.00686131f $X=2.72 $Y=1.835 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_413_n N_A_114_367#_c_525_n 0.0248957f $X=2.93 $Y=2.87 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_421_n N_A_114_367#_c_533_n 0.0298674f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_408_n N_A_114_367#_c_533_n 0.0187823f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_421_n N_A_114_367#_c_535_n 0.01906f $X=7.205 $Y=3.33 $X2=0 $Y2=0
cc_387 N_VPWR_c_408_n N_A_114_367#_c_535_n 0.0124545f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_421_n N_A_114_367#_c_541_n 0.0298674f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_408_n N_A_114_367#_c_541_n 0.0187823f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_421_n N_A_114_367#_c_547_n 0.0298674f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_408_n N_A_114_367#_c_547_n 0.0187823f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_421_n N_A_114_367#_c_553_n 0.037782f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_408_n N_A_114_367#_c_553_n 0.024237f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_394 N_VPWR_c_421_n N_A_114_367#_c_594_n 0.0118138f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_408_n N_A_114_367#_c_594_n 0.00658808f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_416_n N_A_114_367#_c_596_n 0.0117428f $X=1.835 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_408_n N_A_114_367#_c_596_n 0.00652089f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_418_n N_A_114_367#_c_558_n 0.0189236f $X=2.765 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_408_n N_A_114_367#_c_558_n 0.0123859f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_421_n N_A_114_367#_c_562_n 0.01906f $X=7.205 $Y=3.33 $X2=0 $Y2=0
cc_401 N_VPWR_c_408_n N_A_114_367#_c_562_n 0.0124545f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_421_n N_A_114_367#_c_564_n 0.01906f $X=7.205 $Y=3.33 $X2=0 $Y2=0
cc_403 N_VPWR_c_408_n N_A_114_367#_c_564_n 0.0124545f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_421_n N_A_114_367#_c_566_n 0.01906f $X=7.205 $Y=3.33 $X2=0 $Y2=0
cc_405 N_VPWR_c_408_n N_A_114_367#_c_566_n 0.0124545f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_408_n N_Y_M1005_d 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_407 N_VPWR_c_408_n N_Y_M1012_d 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_408 N_VPWR_c_408_n N_Y_M1019_d 0.00225186f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_409 N_VPWR_c_408_n N_Y_M1030_d 0.00281482f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_410 N_VPWR_M1006_d N_Y_c_640_n 0.00130164f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_411 N_VPWR_c_410_n N_Y_c_640_n 0.00190934f $X=0.28 $Y=1.98 $X2=0 $Y2=0
cc_412 N_VPWR_M1006_d N_Y_c_662_n 0.00286567f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_413 N_VPWR_M1017_d N_Y_c_662_n 0.00334119f $X=1.86 $Y=1.835 $X2=0 $Y2=0
cc_414 N_VPWR_M1021_d N_Y_c_662_n 0.00661192f $X=2.72 $Y=1.835 $X2=0 $Y2=0
cc_415 N_VPWR_M1006_d N_Y_c_672_n 8.54197e-19 $X=1 $Y=1.835 $X2=0 $Y2=0
cc_416 N_A_114_367#_c_533_n N_Y_M1005_d 0.00332344f $X=4.125 $Y=2.99 $X2=0.495
+ $Y2=1.675
cc_417 N_A_114_367#_c_541_n N_Y_M1012_d 0.00332344f $X=4.985 $Y=2.99 $X2=0.495
+ $Y2=2.465
cc_418 N_A_114_367#_c_547_n N_Y_M1019_d 0.00332344f $X=5.845 $Y=2.99 $X2=0.495
+ $Y2=2.465
cc_419 N_A_114_367#_c_553_n N_Y_M1030_d 0.00472489f $X=6.855 $Y=2.99 $X2=0 $Y2=0
cc_420 N_A_114_367#_M1010_s N_Y_c_662_n 0.00350572f $X=1.43 $Y=1.835 $X2=1.785
+ $Y2=2.465
cc_421 N_A_114_367#_M1020_s N_Y_c_662_n 0.00333871f $X=2.29 $Y=1.835 $X2=1.785
+ $Y2=2.465
cc_422 N_A_114_367#_M1028_s N_Y_c_662_n 0.00369844f $X=3.29 $Y=1.835 $X2=1.785
+ $Y2=2.465
cc_423 N_A_114_367#_c_521_n N_Y_c_662_n 0.0164886f $X=1.485 $Y=2.375 $X2=1.785
+ $Y2=2.465
cc_424 N_A_114_367#_c_523_n N_Y_c_662_n 0.0306289f $X=2.265 $Y=2.375 $X2=1.785
+ $Y2=2.465
cc_425 N_A_114_367#_c_525_n N_Y_c_662_n 0.0391031f $X=3.265 $Y=2.375 $X2=1.785
+ $Y2=2.465
cc_426 N_A_114_367#_c_527_n N_Y_c_662_n 0.01723f $X=3.43 $Y=2.46 $X2=1.785
+ $Y2=2.465
cc_427 N_A_114_367#_c_596_n N_Y_c_662_n 0.0135055f $X=1.57 $Y=2.455 $X2=1.785
+ $Y2=2.465
cc_428 N_A_114_367#_c_558_n N_Y_c_662_n 0.01723f $X=2.43 $Y=2.455 $X2=1.785
+ $Y2=2.465
cc_429 N_A_114_367#_c_521_n N_Y_c_672_n 0.0089251f $X=1.485 $Y=2.375 $X2=0 $Y2=0
cc_430 N_A_114_367#_c_533_n N_Y_c_758_n 0.0126348f $X=4.125 $Y=2.99 $X2=2.215
+ $Y2=2.465
cc_431 N_A_114_367#_M1008_s N_Y_c_679_n 0.00330483f $X=4.15 $Y=1.835 $X2=2.645
+ $Y2=0.685
cc_432 N_A_114_367#_c_537_n N_Y_c_679_n 0.0170777f $X=4.29 $Y=2.35 $X2=2.645
+ $Y2=0.685
cc_433 N_A_114_367#_M1018_s N_Y_c_689_n 0.00330483f $X=5.01 $Y=1.835 $X2=3.215
+ $Y2=1.675
cc_434 N_A_114_367#_c_543_n N_Y_c_689_n 0.0170777f $X=5.15 $Y=2.35 $X2=3.215
+ $Y2=1.675
cc_435 N_A_114_367#_M1024_s N_Y_c_703_n 0.00330483f $X=5.87 $Y=1.835 $X2=3.645
+ $Y2=2.465
cc_436 N_A_114_367#_c_549_n N_Y_c_703_n 0.0170777f $X=6.01 $Y=2.27 $X2=3.645
+ $Y2=2.465
cc_437 N_A_114_367#_c_518_n N_Y_c_641_n 0.0149317f $X=0.71 $Y=2.115 $X2=4.075
+ $Y2=2.465
cc_438 N_A_114_367#_c_521_n N_Y_c_641_n 0.0042396f $X=1.485 $Y=2.375 $X2=4.075
+ $Y2=2.465
cc_439 N_A_114_367#_c_541_n N_Y_c_723_n 0.0126348f $X=4.985 $Y=2.99 $X2=4.505
+ $Y2=2.465
cc_440 N_A_114_367#_c_547_n N_Y_c_729_n 0.0126348f $X=5.845 $Y=2.99 $X2=4.795
+ $Y2=1.345
cc_441 N_A_114_367#_c_553_n N_Y_c_731_n 0.0196355f $X=6.855 $Y=2.99 $X2=4.795
+ $Y2=0.685
cc_442 N_Y_c_633_n N_VGND_M1004_s 9.27081e-19 $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_443 N_Y_c_660_n N_VGND_M1004_s 8.65291e-19 $X=1.135 $Y=1.09 $X2=0 $Y2=0
cc_444 N_Y_c_633_n N_VGND_M1013_s 0.00176891f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_445 N_Y_c_633_n N_VGND_M1016_s 0.00176891f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_446 N_Y_c_633_n N_A_114_53#_M1011_d 0.00176461f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_447 N_Y_c_633_n N_A_114_53#_M1015_d 0.00176461f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_448 N_Y_c_633_n N_A_114_53#_M1022_d 0.00176461f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_449 N_Y_c_634_n N_A_114_53#_M1002_s 0.00176461f $X=4.495 $Y=1.09 $X2=0 $Y2=0
cc_450 N_Y_c_635_n N_A_114_53#_M1009_s 0.00176461f $X=5.275 $Y=1.09 $X2=0 $Y2=0
cc_451 N_Y_c_636_n N_A_114_53#_M1025_s 0.00250873f $X=6.275 $Y=1.09 $X2=0 $Y2=0
cc_452 N_Y_c_660_n N_A_114_53#_c_923_n 0.00581604f $X=1.135 $Y=1.09 $X2=0 $Y2=0
cc_453 N_Y_c_641_n N_A_114_53#_c_923_n 0.00786795f $X=0.965 $Y=1.665 $X2=0 $Y2=0
cc_454 N_Y_c_633_n N_A_114_53#_c_939_n 0.0165225f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_455 N_Y_c_660_n N_A_114_53#_c_939_n 0.0090121f $X=1.135 $Y=1.09 $X2=0 $Y2=0
cc_456 N_Y_c_633_n N_A_114_53#_c_944_n 0.0323912f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_457 N_Y_c_633_n N_A_114_53#_c_948_n 0.045723f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_458 N_Y_M1000_d N_A_114_53#_c_926_n 0.00176461f $X=3.58 $Y=0.265 $X2=0 $Y2=0
cc_459 N_Y_c_633_n N_A_114_53#_c_926_n 0.00305513f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_460 N_Y_c_673_n N_A_114_53#_c_926_n 0.01417f $X=3.72 $Y=0.86 $X2=0 $Y2=0
cc_461 N_Y_c_634_n N_A_114_53#_c_926_n 0.00305513f $X=4.495 $Y=1.09 $X2=0 $Y2=0
cc_462 N_Y_c_634_n N_A_114_53#_c_953_n 0.0169399f $X=4.495 $Y=1.09 $X2=0 $Y2=0
cc_463 N_Y_M1007_d N_A_114_53#_c_928_n 0.00176461f $X=4.44 $Y=0.265 $X2=0 $Y2=0
cc_464 N_Y_c_634_n N_A_114_53#_c_928_n 0.00305513f $X=4.495 $Y=1.09 $X2=0 $Y2=0
cc_465 N_Y_c_683_n N_A_114_53#_c_928_n 0.01417f $X=4.58 $Y=0.86 $X2=0 $Y2=0
cc_466 N_Y_c_635_n N_A_114_53#_c_928_n 0.00305513f $X=5.275 $Y=1.09 $X2=0 $Y2=0
cc_467 N_Y_c_635_n N_A_114_53#_c_993_n 0.0133318f $X=5.275 $Y=1.09 $X2=0 $Y2=0
cc_468 N_Y_M1014_d N_A_114_53#_c_929_n 0.00176461f $X=5.3 $Y=0.265 $X2=0 $Y2=0
cc_469 N_Y_c_635_n N_A_114_53#_c_929_n 0.00305513f $X=5.275 $Y=1.09 $X2=0 $Y2=0
cc_470 N_Y_c_693_n N_A_114_53#_c_929_n 0.0158587f $X=5.44 $Y=0.86 $X2=0 $Y2=0
cc_471 N_Y_c_636_n N_A_114_53#_c_929_n 0.00306745f $X=6.275 $Y=1.09 $X2=0 $Y2=0
cc_472 N_Y_M1026_d N_A_114_53#_c_930_n 0.00250873f $X=6.23 $Y=0.265 $X2=0 $Y2=0
cc_473 N_Y_c_636_n N_A_114_53#_c_930_n 0.00306745f $X=6.275 $Y=1.09 $X2=0 $Y2=0
cc_474 N_Y_c_707_n N_A_114_53#_c_930_n 0.0194333f $X=6.44 $Y=0.82 $X2=0 $Y2=0
cc_475 N_Y_c_633_n N_A_114_53#_c_1001_n 0.0133318f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_476 N_Y_c_633_n N_A_114_53#_c_1002_n 0.0133318f $X=3.555 $Y=1.09 $X2=0 $Y2=0
cc_477 N_Y_c_636_n N_A_114_53#_c_933_n 0.0207166f $X=6.275 $Y=1.09 $X2=0 $Y2=0
cc_478 N_Y_c_636_n N_A_114_53#_c_934_n 0.00584871f $X=6.275 $Y=1.09 $X2=0 $Y2=0
cc_479 N_VGND_c_808_n N_A_114_53#_c_922_n 0.0143933f $X=0.28 $Y=0.41 $X2=0 $Y2=0
cc_480 N_VGND_c_809_n N_A_114_53#_c_922_n 0.00894674f $X=1.14 $Y=0.41 $X2=0
+ $Y2=0
cc_481 N_VGND_c_818_n N_A_114_53#_c_922_n 0.017694f $X=0.975 $Y=0 $X2=0 $Y2=0
cc_482 N_VGND_c_821_n N_A_114_53#_c_922_n 0.00953185f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_483 N_VGND_c_808_n N_A_114_53#_c_923_n 0.0106547f $X=0.28 $Y=0.41 $X2=0 $Y2=0
cc_484 N_VGND_M1004_s N_A_114_53#_c_939_n 0.00334726f $X=1 $Y=0.265 $X2=0 $Y2=0
cc_485 N_VGND_c_809_n N_A_114_53#_c_939_n 0.0161464f $X=1.14 $Y=0.41 $X2=0 $Y2=0
cc_486 N_VGND_c_814_n N_A_114_53#_c_939_n 0.00238814f $X=1.835 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_c_818_n N_A_114_53#_c_939_n 0.00239434f $X=0.975 $Y=0 $X2=0 $Y2=0
cc_488 N_VGND_c_821_n N_A_114_53#_c_939_n 0.0102174f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_489 N_VGND_c_809_n N_A_114_53#_c_924_n 0.00892713f $X=1.14 $Y=0.41 $X2=0
+ $Y2=0
cc_490 N_VGND_c_810_n N_A_114_53#_c_924_n 0.00892713f $X=2 $Y=0.41 $X2=0 $Y2=0
cc_491 N_VGND_c_814_n N_A_114_53#_c_924_n 0.0118996f $X=1.835 $Y=0 $X2=0 $Y2=0
cc_492 N_VGND_c_821_n N_A_114_53#_c_924_n 0.00650442f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_493 N_VGND_M1013_s N_A_114_53#_c_944_n 0.00335857f $X=1.86 $Y=0.265 $X2=0
+ $Y2=0
cc_494 N_VGND_c_810_n N_A_114_53#_c_944_n 0.0161464f $X=2 $Y=0.41 $X2=0 $Y2=0
cc_495 N_VGND_c_814_n N_A_114_53#_c_944_n 0.00238814f $X=1.835 $Y=0 $X2=0 $Y2=0
cc_496 N_VGND_c_816_n N_A_114_53#_c_944_n 0.00238814f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_497 N_VGND_c_821_n N_A_114_53#_c_944_n 0.0102073f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_498 N_VGND_c_810_n N_A_114_53#_c_925_n 0.00892713f $X=2 $Y=0.41 $X2=0 $Y2=0
cc_499 N_VGND_c_811_n N_A_114_53#_c_925_n 0.00892713f $X=2.86 $Y=0.41 $X2=0
+ $Y2=0
cc_500 N_VGND_c_816_n N_A_114_53#_c_925_n 0.0118996f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_501 N_VGND_c_821_n N_A_114_53#_c_925_n 0.00650442f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_502 N_VGND_M1016_s N_A_114_53#_c_948_n 0.00335857f $X=2.72 $Y=0.265 $X2=0
+ $Y2=0
cc_503 N_VGND_c_811_n N_A_114_53#_c_948_n 0.0161464f $X=2.86 $Y=0.41 $X2=0 $Y2=0
cc_504 N_VGND_c_816_n N_A_114_53#_c_948_n 0.00238814f $X=2.695 $Y=0 $X2=0 $Y2=0
cc_505 N_VGND_c_819_n N_A_114_53#_c_948_n 0.00238814f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_506 N_VGND_c_821_n N_A_114_53#_c_948_n 0.0102073f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_507 N_VGND_c_819_n N_A_114_53#_c_926_n 0.0384393f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_508 N_VGND_c_821_n N_A_114_53#_c_926_n 0.0216758f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_509 N_VGND_c_811_n N_A_114_53#_c_927_n 0.00652315f $X=2.86 $Y=0.41 $X2=0
+ $Y2=0
cc_510 N_VGND_c_819_n N_A_114_53#_c_927_n 0.0120413f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_511 N_VGND_c_821_n N_A_114_53#_c_927_n 0.00658185f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_512 N_VGND_c_819_n N_A_114_53#_c_928_n 0.0384393f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_c_821_n N_A_114_53#_c_928_n 0.0216758f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_819_n N_A_114_53#_c_929_n 0.0428729f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_515 N_VGND_c_821_n N_A_114_53#_c_929_n 0.0241933f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_516 N_VGND_c_819_n N_A_114_53#_c_930_n 0.0423044f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_821_n N_A_114_53#_c_930_n 0.0239316f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_819_n N_A_114_53#_c_931_n 0.0232038f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_821_n N_A_114_53#_c_931_n 0.0125481f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_819_n N_A_114_53#_c_932_n 0.012043f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_821_n N_A_114_53#_c_932_n 0.00658217f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_819_n N_A_114_53#_c_933_n 0.0232899f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_523 N_VGND_c_821_n N_A_114_53#_c_933_n 0.0126625f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_524 N_VGND_c_813_n N_A_114_53#_c_934_n 0.0329656f $X=7.37 $Y=0.41 $X2=0 $Y2=0
cc_525 N_VGND_c_819_n N_A_114_53#_c_934_n 0.0235688f $X=7.285 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_821_n N_A_114_53#_c_934_n 0.0127152f $X=7.44 $Y=0 $X2=0 $Y2=0
