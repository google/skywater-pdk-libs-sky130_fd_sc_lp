* File: sky130_fd_sc_lp__dlxbn_1.spice
* Created: Wed Sep  2 09:47:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxbn_1.pex.spice"
.subckt sky130_fd_sc_lp__dlxbn_1  VNB VPB D GATE_N VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_D_M1015_g N_A_34_407#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_219_135#_M1008_d N_GATE_N_M1008_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_219_135#_M1010_g N_A_363_483#_M1010_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1019 A_554_47# N_A_34_407#_M1019_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_626_47#_M1011_d N_A_219_135#_M1011_g A_554_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=17.136 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1002 A_734_47# N_A_363_483#_M1002_g N_A_626_47#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=14.28 M=1 R=2.8
+ SA=75001.5 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_806_385#_M1007_g A_734_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.0819 PD=0.81 PS=0.81 NRD=15.708 NRS=39.996 M=1 R=2.8 SA=75002.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_806_385#_M1017_d N_A_626_47#_M1017_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=2.856 M=1 R=5.6
+ SA=75001.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_806_385#_M1004_g N_A_1069_161#_M1004_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.2121 AS=0.1113 PD=1.16 PS=1.37 NRD=128.568 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1018 N_Q_N_M1018_d N_A_1069_161#_M1018_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.4242 PD=2.21 PS=2.32 NRD=0 NRS=49.992 M=1 R=5.6
+ SA=75000.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_Q_M1003_d N_A_806_385#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_D_M1012_g N_A_34_407#_M1012_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1152 AS=0.1696 PD=1 PS=1.81 NRD=24.6053 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1005 N_A_219_135#_M1005_d N_GATE_N_M1005_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.3459 AS=0.1152 PD=2.7 PS=1 NRD=149.424 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1014 N_VPWR_M1014_d N_A_219_135#_M1014_g N_A_363_483#_M1014_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1728 AS=0.1696 PD=1.18 PS=1.81 NRD=44.6205 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1021 A_584_483# N_A_34_407#_M1021_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1728 PD=0.85 PS=1.18 NRD=15.3857 NRS=35.3812 M=1 R=4.26667
+ SA=75000.9 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1000 N_A_626_47#_M1000_d N_A_363_483#_M1000_g A_584_483# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.134098 AS=0.0672 PD=1.24377 PS=0.85 NRD=16.9223 NRS=15.3857 M=1
+ R=4.26667 SA=75001.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1006 A_764_483# N_A_219_135#_M1006_g N_A_626_47#_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0880019 PD=0.63 PS=0.816226 NRD=23.443 NRS=26.9693 M=1
+ R=2.8 SA=75001.8 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_806_385#_M1009_g A_764_483# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1239 AS=0.0441 PD=0.94 PS=0.63 NRD=112.566 NRS=23.443 M=1 R=2.8
+ SA=75002.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1020 N_A_806_385#_M1020_d N_A_626_47#_M1020_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3717 PD=3.05 PS=2.82 NRD=0 NRS=2.3443 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_A_806_385#_M1016_g N_A_1069_161#_M1016_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.12864 AS=0.1696 PD=1.07789 PS=1.81 NRD=13.8491 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1001 N_Q_N_M1001_d N_A_1069_161#_M1001_g N_VPWR_M1016_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.25326 PD=3.05 PS=2.12211 NRD=0 NRS=1.8124 M=1 R=8.4
+ SA=75000.4 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1013 N_Q_M1013_d N_A_806_385#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX22_noxref VNB VPB NWDIODE A=16.1256 P=21.03
*
.include "sky130_fd_sc_lp__dlxbn_1.pxi.spice"
*
.ends
*
*
