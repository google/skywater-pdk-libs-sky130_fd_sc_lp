* File: sky130_fd_sc_lp__a2111oi_2.pex.spice
* Created: Fri Aug 28 09:46:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111OI_2%C1 3 7 11 15 17 20 25 29 32 33
c73 32 0 1.20436e-19 $X=1.81 $Y=1.46
c74 20 0 7.76129e-20 $X=0.29 $Y=1.46
c75 7 0 1.16478e-19 $X=0.5 $Y=2.465
r76 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.46
+ $X2=1.81 $Y2=1.625
r77 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.81 $Y=1.46
+ $X2=1.81 $Y2=1.295
r78 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.46 $X2=1.81 $Y2=1.46
r79 25 40 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.69
r80 25 33 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.46
r81 21 29 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.29 $Y=1.46 $X2=0.5
+ $Y2=1.46
r82 20 23 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.29 $Y=1.46
+ $X2=0.29 $Y2=1.69
r83 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.46 $X2=0.29 $Y2=1.46
r84 18 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=1.69
+ $X2=0.29 $Y2=1.69
r85 17 40 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=1.525 $Y=1.69
+ $X2=1.71 $Y2=1.69
r86 17 18 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=1.525 $Y=1.69
+ $X2=0.455 $Y2=1.69
r87 15 34 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.9 $Y=0.655 $X2=1.9
+ $Y2=1.295
r88 11 35 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.79 $Y=2.465
+ $X2=1.79 $Y2=1.625
r89 5 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.625 $X2=0.5
+ $Y2=1.46
r90 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.5 $Y=1.625 $X2=0.5
+ $Y2=2.465
r91 1 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.295 $X2=0.5
+ $Y2=1.46
r92 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.5 $Y=1.295 $X2=0.5
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%D1 1 3 6 8 10 13 15 16 24
c51 16 0 1.20436e-19 $X=1.2 $Y=1.295
c52 6 0 7.76129e-20 $X=0.93 $Y=2.465
r53 22 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.02 $Y=1.35
+ $X2=1.36 $Y2=1.35
r54 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.02
+ $Y=1.35 $X2=1.02 $Y2=1.35
r55 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.93 $Y=1.35 $X2=1.02
+ $Y2=1.35
r56 16 23 9.21954 $w=2.23e-07 $l=1.8e-07 $layer=LI1_cond $X=1.2 $Y=1.322
+ $X2=1.02 $Y2=1.322
r57 15 23 15.3659 $w=2.23e-07 $l=3e-07 $layer=LI1_cond $X=0.72 $Y=1.322 $X2=1.02
+ $Y2=1.322
r58 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.515
+ $X2=1.36 $Y2=1.35
r59 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.36 $Y=1.515
+ $X2=1.36 $Y2=2.465
r60 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.36 $Y2=1.35
r61 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.36 $Y2=0.655
r62 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.515
+ $X2=0.93 $Y2=1.35
r63 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.93 $Y=1.515 $X2=0.93
+ $Y2=2.465
r64 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=1.35
r65 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.93 $Y=1.185 $X2=0.93
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%B1 3 7 11 15 17 18 26 27
c48 26 0 1.74471e-19 $X=2.69 $Y=1.51
c49 7 0 1.47259e-19 $X=2.375 $Y=0.655
r50 25 27 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=2.69 $Y=1.51
+ $X2=2.915 $Y2=1.51
r51 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.69
+ $Y=1.51 $X2=2.69 $Y2=1.51
r52 23 25 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=2.375 $Y=1.51
+ $X2=2.69 $Y2=1.51
r53 21 23 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=2.26 $Y=1.51
+ $X2=2.375 $Y2=1.51
r54 18 26 1.64635 $w=3.48e-07 $l=5e-08 $layer=LI1_cond $X=2.64 $Y=1.6 $X2=2.69
+ $Y2=1.6
r55 17 18 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.6 $X2=2.64
+ $Y2=1.6
r56 13 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.345
+ $X2=2.915 $Y2=1.51
r57 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.915 $Y=1.345
+ $X2=2.915 $Y2=0.655
r58 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.675
+ $X2=2.69 $Y2=1.51
r59 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.69 $Y=1.675
+ $X2=2.69 $Y2=2.465
r60 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.345
+ $X2=2.375 $Y2=1.51
r61 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.375 $Y=1.345
+ $X2=2.375 $Y2=0.655
r62 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.675
+ $X2=2.26 $Y2=1.51
r63 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.26 $Y=1.675 $X2=2.26
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%A1 3 7 11 15 17 20 21 25 26 34 39 46
c77 34 0 1.74471e-19 $X=3.64 $Y=1.51
r78 32 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.55 $Y=1.51 $X2=3.64
+ $Y2=1.51
r79 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.51 $X2=3.55 $Y2=1.51
r80 29 32 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.345 $Y=1.51
+ $X2=3.55 $Y2=1.51
r81 26 46 7.2638 $w=4.38e-07 $l=1.05e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.185 $Y2=1.565
r82 26 39 3.01207 $w=4.38e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.965 $Y2=1.565
r83 25 39 9.56004 $w=4.38e-07 $l=3.65e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.965 $Y2=1.565
r84 25 33 1.30959 $w=4.38e-07 $l=5e-08 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.55
+ $Y2=1.565
r85 21 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.06 $Y=1.51
+ $X2=5.06 $Y2=1.675
r86 21 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.06 $Y=1.51
+ $X2=5.06 $Y2=1.345
r87 20 23 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=5.025 $Y=1.51
+ $X2=5.025 $Y2=1.7
r88 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.06
+ $Y=1.51 $X2=5.06 $Y2=1.51
r89 17 23 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.895 $Y=1.7
+ $X2=5.025 $Y2=1.7
r90 17 46 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.895 $Y=1.7
+ $X2=4.185 $Y2=1.7
r91 15 38 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.97 $Y=2.465
+ $X2=4.97 $Y2=1.675
r92 11 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.97 $Y=0.655
+ $X2=4.97 $Y2=1.345
r93 5 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.64 $Y=1.675
+ $X2=3.64 $Y2=1.51
r94 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.64 $Y=1.675 $X2=3.64
+ $Y2=2.465
r95 1 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.345
+ $X2=3.345 $Y2=1.51
r96 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.345 $Y=1.345
+ $X2=3.345 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%A2 1 3 6 8 12 16 17 18 20 21
r59 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=1.35
+ $X2=4.52 $Y2=1.515
r60 20 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.52 $Y=1.26 $X2=4.52
+ $Y2=1.35
r61 20 21 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.52 $Y=1.26 $X2=4.52
+ $Y2=1.185
r62 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.52
+ $Y=1.35 $X2=4.52 $Y2=1.35
r63 16 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.54 $Y=0.655
+ $X2=4.54 $Y2=1.185
r64 12 25 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.5 $Y=2.465 $X2=4.5
+ $Y2=1.515
r65 9 17 5.30422 $w=1.5e-07 $l=8.8e-08 $layer=POLY_cond $X=4.145 $Y=1.26
+ $X2=4.057 $Y2=1.26
r66 8 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.26
+ $X2=4.52 $Y2=1.26
r67 8 9 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.355 $Y=1.26
+ $X2=4.145 $Y2=1.26
r68 4 17 20.4101 $w=1.5e-07 $l=8.12404e-08 $layer=POLY_cond $X=4.07 $Y=1.335
+ $X2=4.057 $Y2=1.26
r69 4 6 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=4.07 $Y=1.335
+ $X2=4.07 $Y2=2.465
r70 1 17 20.4101 $w=1.5e-07 $l=8.07775e-08 $layer=POLY_cond $X=4.045 $Y=1.185
+ $X2=4.057 $Y2=1.26
r71 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.045 $Y=1.185
+ $X2=4.045 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%A_32_367# 1 2 3 10 12 14 18 22 27
c36 3 0 4.98153e-20 $X=2.765 $Y=1.835
r37 20 27 6.21488 $w=2.35e-07 $l=1.48e-07 $layer=LI1_cond $X=2.165 $Y=2.945
+ $X2=2.017 $Y2=2.945
r38 20 22 32.8003 $w=2.58e-07 $l=7.4e-07 $layer=LI1_cond $X=2.165 $Y=2.945
+ $X2=2.905 $Y2=2.945
r39 16 27 0.538047 $w=2.95e-07 $l=1.3e-07 $layer=LI1_cond $X=2.017 $Y=2.815
+ $X2=2.017 $Y2=2.945
r40 16 18 13.8684 $w=2.93e-07 $l=3.55e-07 $layer=LI1_cond $X=2.017 $Y=2.815
+ $X2=2.017 $Y2=2.46
r41 15 25 3.99943 $w=2.1e-07 $l=1.4e-07 $layer=LI1_cond $X=0.4 $Y=2.97 $X2=0.26
+ $Y2=2.97
r42 14 27 6.21488 $w=2.35e-07 $l=1.59009e-07 $layer=LI1_cond $X=1.87 $Y=2.97
+ $X2=2.017 $Y2=2.945
r43 14 15 77.6364 $w=2.08e-07 $l=1.47e-06 $layer=LI1_cond $X=1.87 $Y=2.97
+ $X2=0.4 $Y2=2.97
r44 10 25 2.99957 $w=2.8e-07 $l=1.05e-07 $layer=LI1_cond $X=0.26 $Y=2.865
+ $X2=0.26 $Y2=2.97
r45 10 12 30.6632 $w=2.78e-07 $l=7.45e-07 $layer=LI1_cond $X=0.26 $Y=2.865
+ $X2=0.26 $Y2=2.12
r46 3 22 600 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.835 $X2=2.905 $Y2=2.93
r47 2 27 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.835 $X2=2.005 $Y2=2.91
r48 2 18 600 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.835 $X2=2.005 $Y2=2.46
r49 1 25 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=2.91
r50 1 12 400 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%A_115_367# 1 2 9 11 12 14
r17 14 16 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=1.575 $Y=2.46
+ $X2=1.575 $Y2=2.61
r18 11 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.45 $Y=2.61
+ $X2=1.575 $Y2=2.61
r19 11 12 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.45 $Y=2.61
+ $X2=0.83 $Y2=2.61
r20 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.7 $Y=2.525
+ $X2=0.83 $Y2=2.61
r21 7 9 17.9515 $w=2.58e-07 $l=4.05e-07 $layer=LI1_cond $X=0.7 $Y=2.525 $X2=0.7
+ $Y2=2.12
r22 2 14 600 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=1 $X=1.435
+ $Y=1.835 $X2=1.575 $Y2=2.46
r23 1 9 300 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=1.835 $X2=0.715 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%Y 1 2 3 4 5 6 21 23 24 27 29 31 35 37 41
+ 43 46 47 52 53 56 59 60 61 69
c130 61 0 4.98153e-20 $X=3.12 $Y=2.035
c131 53 0 1.47259e-19 $X=2.13 $Y=0.955
c132 47 0 1.16478e-19 $X=1.132 $Y=2.035
r133 66 69 1.70732 $w=2.68e-07 $l=4e-08 $layer=LI1_cond $X=3.16 $Y=1.255
+ $X2=3.16 $Y2=1.295
r134 61 67 0.161356 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=3.16 $Y=2.035
+ $X2=3.16 $Y2=1.945
r135 60 67 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.16 $Y=1.665
+ $X2=3.16 $Y2=1.945
r136 59 66 3.14896 $w=3e-07 $l=9.88686e-08 $layer=LI1_cond $X=3.13 $Y=1.17
+ $X2=3.16 $Y2=1.255
r137 59 60 14.8537 $w=2.68e-07 $l=3.48e-07 $layer=LI1_cond $X=3.16 $Y=1.317
+ $X2=3.16 $Y2=1.665
r138 59 69 0.939028 $w=2.68e-07 $l=2.2e-08 $layer=LI1_cond $X=3.16 $Y=1.317
+ $X2=3.16 $Y2=1.295
r139 56 58 15.3188 $w=6.38e-07 $l=6.75e-07 $layer=LI1_cond $X=5.34 $Y=0.42
+ $X2=5.34 $Y2=1.095
r140 53 54 9.57299 $w=2.74e-07 $l=2.15e-07 $layer=LI1_cond $X=2.13 $Y=0.955
+ $X2=2.13 $Y2=1.17
r141 47 50 6.7407 $w=2.63e-07 $l=1.55e-07 $layer=LI1_cond $X=1.132 $Y=2.035
+ $X2=1.132 $Y2=2.19
r142 46 58 29.5851 $w=3.33e-07 $l=8.6e-07 $layer=LI1_cond $X=5.492 $Y=1.955
+ $X2=5.492 $Y2=1.095
r143 44 61 7.28786 $w=1.75e-07 $l=1.37477e-07 $layer=LI1_cond $X=3.295 $Y=2.04
+ $X2=3.16 $Y2=2.035
r144 43 46 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=5.325 $Y=2.04
+ $X2=5.492 $Y2=1.955
r145 43 44 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=5.325 $Y=2.04
+ $X2=3.295 $Y2=2.04
r146 39 59 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=1.085 $X2=3.13
+ $Y2=1.17
r147 39 41 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.13 $Y=1.085
+ $X2=3.13 $Y2=0.375
r148 38 54 3.52985 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=1.17
+ $X2=2.13 $Y2=1.17
r149 37 59 3.44808 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=1.17
+ $X2=3.13 $Y2=1.17
r150 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.965 $Y=1.17
+ $X2=2.295 $Y2=1.17
r151 33 53 3.52979 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=0.87
+ $X2=2.13 $Y2=0.955
r152 33 35 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.13 $Y=0.87
+ $X2=2.13 $Y2=0.42
r153 32 52 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.295 $Y=0.955
+ $X2=1.172 $Y2=0.955
r154 31 53 3.52985 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=0.955
+ $X2=2.13 $Y2=0.955
r155 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.965 $Y=0.955
+ $X2=1.295 $Y2=0.955
r156 30 47 3.00163 $w=1.8e-07 $l=1.33e-07 $layer=LI1_cond $X=1.265 $Y=2.035
+ $X2=1.132 $Y2=2.035
r157 29 61 7.28786 $w=1.75e-07 $l=1.35e-07 $layer=LI1_cond $X=3.025 $Y=2.035
+ $X2=3.16 $Y2=2.035
r158 29 30 108.444 $w=1.78e-07 $l=1.76e-06 $layer=LI1_cond $X=3.025 $Y=2.035
+ $X2=1.265 $Y2=2.035
r159 25 52 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.172 $Y=0.87
+ $X2=1.172 $Y2=0.955
r160 25 27 20.6969 $w=2.43e-07 $l=4.4e-07 $layer=LI1_cond $X=1.172 $Y=0.87
+ $X2=1.172 $Y2=0.43
r161 23 52 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=1.05 $Y=0.955
+ $X2=1.172 $Y2=0.955
r162 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.05 $Y=0.955
+ $X2=0.38 $Y2=0.955
r163 19 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.25 $Y=0.87
+ $X2=0.38 $Y2=0.955
r164 19 21 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=0.25 $Y=0.87
+ $X2=0.25 $Y2=0.43
r165 6 50 600 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.005
+ $Y=1.835 $X2=1.145 $Y2=2.19
r166 5 56 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.045
+ $Y=0.235 $X2=5.185 $Y2=0.42
r167 4 41 91 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=2 $X=2.99
+ $Y=0.235 $X2=3.13 $Y2=0.375
r168 3 35 91 $w=1.7e-07 $l=2.56271e-07 $layer=licon1_NDIFF $count=2 $X=1.975
+ $Y=0.235 $X2=2.145 $Y2=0.42
r169 2 27 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.235 $X2=1.145 $Y2=0.43
r170 1 21 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%A_467_367# 1 2 3 4 13 19 21 25 27 29 31 34
+ 36
r44 29 38 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.21 $Y=2.465
+ $X2=5.21 $Y2=2.38
r45 29 31 18.3156 $w=2.78e-07 $l=4.45e-07 $layer=LI1_cond $X=5.21 $Y=2.465
+ $X2=5.21 $Y2=2.91
r46 28 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.4 $Y=2.38
+ $X2=4.295 $Y2=2.38
r47 27 38 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.07 $Y=2.38 $X2=5.21
+ $Y2=2.38
r48 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.07 $Y=2.38 $X2=4.4
+ $Y2=2.38
r49 23 36 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=2.465
+ $X2=4.295 $Y2=2.38
r50 23 25 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=4.295 $Y=2.465
+ $X2=4.295 $Y2=2.91
r51 22 34 5.16603 $w=2.6e-07 $l=1.69115e-07 $layer=LI1_cond $X=3.52 $Y=2.38
+ $X2=3.39 $Y2=2.47
r52 21 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.19 $Y=2.38
+ $X2=4.295 $Y2=2.38
r53 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.19 $Y=2.38
+ $X2=3.52 $Y2=2.38
r54 17 34 1.34256 $w=2.6e-07 $l=1.75e-07 $layer=LI1_cond $X=3.39 $Y=2.645
+ $X2=3.39 $Y2=2.47
r55 17 19 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=3.39 $Y=2.645
+ $X2=3.39 $Y2=2.91
r56 13 34 5.16603 $w=2.6e-07 $l=1.3e-07 $layer=LI1_cond $X=3.26 $Y=2.47 $X2=3.39
+ $Y2=2.47
r57 13 15 25.8477 $w=3.48e-07 $l=7.85e-07 $layer=LI1_cond $X=3.26 $Y=2.47
+ $X2=2.475 $Y2=2.47
r58 4 38 600 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=1 $X=5.045
+ $Y=1.835 $X2=5.185 $Y2=2.38
r59 4 31 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.045
+ $Y=1.835 $X2=5.185 $Y2=2.91
r60 3 36 600 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=1 $X=4.145
+ $Y=1.835 $X2=4.285 $Y2=2.38
r61 3 25 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.145
+ $Y=1.835 $X2=4.285 $Y2=2.91
r62 2 34 600 $w=1.7e-07 $l=6.04276e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.835 $X2=3.425 $Y2=2.38
r63 2 19 600 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.835 $X2=3.425 $Y2=2.91
r64 1 15 600 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=1 $X=2.335
+ $Y=1.835 $X2=2.475 $Y2=2.48
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%VPWR 1 2 9 13 16 17 19 20 21 34 35
r67 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r68 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r69 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r70 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r71 28 29 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r72 24 28 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=3.6 $Y2=3.33
r73 24 25 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 21 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r75 21 25 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 19 31 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=4.57 $Y=3.33 $X2=4.56
+ $Y2=3.33
r77 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.57 $Y=3.33
+ $X2=4.735 $Y2=3.33
r78 18 34 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.9 $Y=3.33 $X2=5.52
+ $Y2=3.33
r79 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=3.33
+ $X2=4.735 $Y2=3.33
r80 16 28 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.69 $Y=3.33 $X2=3.6
+ $Y2=3.33
r81 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.69 $Y=3.33
+ $X2=3.855 $Y2=3.33
r82 15 31 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=4.56 $Y2=3.33
r83 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=3.855 $Y2=3.33
r84 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.735 $Y=3.245
+ $X2=4.735 $Y2=3.33
r85 11 13 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=4.735 $Y=3.245
+ $X2=4.735 $Y2=2.76
r86 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=3.245
+ $X2=3.855 $Y2=3.33
r87 7 9 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.855 $Y=3.245
+ $X2=3.855 $Y2=2.76
r88 2 13 600 $w=1.7e-07 $l=1.00181e-06 $layer=licon1_PDIFF $count=1 $X=4.575
+ $Y=1.835 $X2=4.735 $Y2=2.76
r89 1 9 600 $w=1.7e-07 $l=9.92535e-07 $layer=licon1_PDIFF $count=1 $X=3.715
+ $Y=1.835 $X2=3.855 $Y2=2.76
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39 44
+ 60 61 64 67 70
r71 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r72 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r73 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r74 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r75 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r76 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r77 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r78 55 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r79 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r80 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r81 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r82 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r83 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.63
+ $Y2=0
r84 49 51 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.12
+ $Y2=0
r85 48 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r86 48 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r87 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r88 45 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=1.63
+ $Y2=0
r89 45 47 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0 $X2=2.16
+ $Y2=0
r90 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.63
+ $Y2=0
r91 44 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.16
+ $Y2=0
r92 43 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r93 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r94 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r95 40 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.715
+ $Y2=0
r96 40 42 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.2
+ $Y2=0
r97 39 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.63
+ $Y2=0
r98 39 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.2
+ $Y2=0
r99 37 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r100 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r101 34 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.715
+ $Y2=0
r102 34 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r103 32 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r104 32 71 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r105 30 54 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.125 $Y=0 $X2=4.08
+ $Y2=0
r106 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.125 $Y=0 $X2=4.29
+ $Y2=0
r107 29 57 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.455 $Y=0
+ $X2=4.56 $Y2=0
r108 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=0 $X2=4.29
+ $Y2=0
r109 25 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=0.085
+ $X2=4.29 $Y2=0
r110 25 27 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.29 $Y=0.085
+ $X2=4.29 $Y2=0.575
r111 21 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0
r112 21 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.38
r113 17 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0
r114 17 19 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0.575
r115 13 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r116 13 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.575
r117 4 27 182 $w=1.7e-07 $l=4.16413e-07 $layer=licon1_NDIFF $count=1 $X=4.12
+ $Y=0.235 $X2=4.29 $Y2=0.575
r118 3 23 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=2.45
+ $Y=0.235 $X2=2.63 $Y2=0.38
r119 2 19 182 $w=1.7e-07 $l=4.26497e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.235 $X2=1.63 $Y2=0.575
r120 1 15 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__A2111OI_2%A_684_47# 1 2 9 11 12 15
r22 13 15 23.0489 $w=2.23e-07 $l=4.5e-07 $layer=LI1_cond $X=4.737 $Y=0.87
+ $X2=4.737 $Y2=0.42
r23 11 13 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=4.625 $Y=0.955
+ $X2=4.737 $Y2=0.87
r24 11 12 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.625 $Y=0.955
+ $X2=3.86 $Y2=0.955
r25 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.695 $Y=0.87
+ $X2=3.86 $Y2=0.955
r26 7 9 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.695 $Y=0.87
+ $X2=3.695 $Y2=0.375
r27 2 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.615
+ $Y=0.235 $X2=4.755 $Y2=0.42
r28 1 9 91 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.235 $X2=3.695 $Y2=0.375
.ends

