* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21ba_lp A1 A2 B1_N VGND VNB VPB VPWR X
X0 VPWR B1_N a_317_29# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_708_75# a_253_389# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_317_29# B1_N a_550_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_550_75# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_253_389# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VPWR A1 a_155_389# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VGND A2 a_34_55# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_34_55# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_34_55# a_317_29# a_253_389# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_155_389# A2 a_253_389# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VGND a_253_389# a_708_75# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_253_389# a_317_29# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
