* File: sky130_fd_sc_lp__a31o_2.pex.spice
* Created: Fri Aug 28 09:59:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31O_2%A_85_23# 1 2 9 13 15 17 20 23 26 27 28 29 32
+ 36 41 42 43
c100 41 0 5.77941e-20 $X=1.07 $Y=1.36
r101 45 46 48.406 $w=2.34e-07 $l=2.35e-07 $layer=POLY_cond $X=0.695 $Y=1.375
+ $X2=0.93 $Y2=1.375
r102 42 48 11.3291 $w=2.34e-07 $l=5.5e-08 $layer=POLY_cond $X=1.07 $Y=1.375
+ $X2=1.125 $Y2=1.375
r103 42 46 28.8376 $w=2.34e-07 $l=1.4e-07 $layer=POLY_cond $X=1.07 $Y=1.375
+ $X2=0.93 $Y2=1.375
r104 41 43 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=1.36
+ $X2=1.165 $Y2=1.195
r105 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.36 $X2=1.07 $Y2=1.36
r106 36 38 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=3.39 $Y=1.98
+ $X2=3.39 $Y2=2.91
r107 34 36 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=3.39 $Y=1.875
+ $X2=3.39 $Y2=1.98
r108 30 32 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.855 $Y=0.855
+ $X2=2.855 $Y2=0.395
r109 28 34 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.26 $Y=1.79
+ $X2=3.39 $Y2=1.875
r110 28 29 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=3.26 $Y=1.79
+ $X2=1.345 $Y2=1.79
r111 26 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.69 $Y=0.94
+ $X2=2.855 $Y2=0.855
r112 26 27 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=2.69 $Y=0.94
+ $X2=1.345 $Y2=0.94
r113 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.26 $Y=1.025
+ $X2=1.345 $Y2=0.94
r114 24 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.26 $Y=1.025
+ $X2=1.26 $Y2=1.195
r115 23 29 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=1.165 $Y=1.705
+ $X2=1.345 $Y2=1.79
r116 22 41 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.165 $Y=1.375
+ $X2=1.165 $Y2=1.36
r117 22 23 10.5641 $w=3.58e-07 $l=3.3e-07 $layer=LI1_cond $X=1.165 $Y=1.375
+ $X2=1.165 $Y2=1.705
r118 18 48 13.1928 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.125 $Y=1.525
+ $X2=1.125 $Y2=1.375
r119 18 20 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.125 $Y=1.525
+ $X2=1.125 $Y2=2.465
r120 15 46 13.1928 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.93 $Y=1.195
+ $X2=0.93 $Y2=1.375
r121 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.93 $Y=1.195
+ $X2=0.93 $Y2=0.665
r122 11 45 13.1928 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.695 $Y=1.525
+ $X2=0.695 $Y2=1.375
r123 11 13 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=0.695 $Y=1.525
+ $X2=0.695 $Y2=2.465
r124 7 45 40.1667 $w=2.34e-07 $l=1.95e-07 $layer=POLY_cond $X=0.5 $Y=1.375
+ $X2=0.695 $Y2=1.375
r125 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.5 $Y=1.375 $X2=0.5
+ $Y2=0.665
r126 2 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.835 $X2=3.355 $Y2=2.91
r127 2 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.835 $X2=3.355 $Y2=1.98
r128 1 32 91 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_NDIFF $count=2 $X=2.675
+ $Y=0.245 $X2=2.855 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_2%A3 3 7 8 11 13
r31 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.36
+ $X2=1.61 $Y2=1.525
r32 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.36
+ $X2=1.61 $Y2=1.195
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.36 $X2=1.61 $Y2=1.36
r34 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.7 $Y=0.665 $X2=1.7
+ $Y2=1.195
r35 3 14 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.635 $Y=2.465 $X2=1.635
+ $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_2%A2 3 6 8 11 13
c33 8 0 5.77941e-20 $X=2.16 $Y=1.295
r34 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.36
+ $X2=2.15 $Y2=1.525
r35 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.36
+ $X2=2.15 $Y2=1.195
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.36 $X2=2.15 $Y2=1.36
r37 6 14 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.065 $Y=2.465 $X2=2.065
+ $Y2=1.525
r38 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.06 $Y=0.665
+ $X2=2.06 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_2%A1 3 6 8 9 13 15
r34 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.36
+ $X2=2.69 $Y2=1.525
r35 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.36
+ $X2=2.69 $Y2=1.195
r36 8 9 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.32 $X2=3.12
+ $Y2=1.32
r37 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.36 $X2=2.69 $Y2=1.36
r38 6 16 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.71 $Y=2.465 $X2=2.71
+ $Y2=1.525
r39 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.6 $Y=0.665 $X2=2.6
+ $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_2%B1 1 3 6 8 13
r23 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.47
+ $Y=1.36 $X2=3.47 $Y2=1.36
r24 10 13 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.14 $Y=1.36
+ $X2=3.47 $Y2=1.36
r25 8 14 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.6 $Y=1.36 $X2=3.47
+ $Y2=1.36
r26 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.14 $Y=1.525
+ $X2=3.14 $Y2=1.36
r27 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.14 $Y=1.525 $X2=3.14
+ $Y2=2.465
r28 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.14 $Y=1.195
+ $X2=3.14 $Y2=1.36
r29 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.14 $Y=1.195 $X2=3.14
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_2%VPWR 1 2 3 10 12 18 24 27 28 30 31 32 45 46
r51 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r53 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 42 45 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 40 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 37 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 34 49 3.99156 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r61 34 36 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=1.2 $Y2=3.33
r62 32 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 32 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 30 39 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=3.33
+ $X2=2.39 $Y2=3.33
r66 29 42 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.39 $Y2=3.33
r68 27 36 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.22 $Y=3.33 $X2=1.2
+ $Y2=3.33
r69 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=3.33
+ $X2=1.385 $Y2=3.33
r70 26 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=3.33
+ $X2=1.385 $Y2=3.33
r72 22 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=3.245
+ $X2=2.39 $Y2=3.33
r73 22 24 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.39 $Y=3.245
+ $X2=2.39 $Y2=2.57
r74 18 21 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=1.385 $Y=2.13
+ $X2=1.385 $Y2=2.95
r75 16 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.385 $Y=3.245
+ $X2=1.385 $Y2=3.33
r76 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=3.245
+ $X2=1.385 $Y2=2.95
r77 12 15 42.5517 $w=2.58e-07 $l=9.6e-07 $layer=LI1_cond $X=0.335 $Y=1.99
+ $X2=0.335 $Y2=2.95
r78 10 49 3.22066 $w=2.6e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.335 $Y=3.245
+ $X2=0.232 $Y2=3.33
r79 10 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=3.245
+ $X2=0.335 $Y2=2.95
r80 3 24 300 $w=1.7e-07 $l=8.50867e-07 $layer=licon1_PDIFF $count=2 $X=2.14
+ $Y=1.835 $X2=2.39 $Y2=2.57
r81 2 21 400 $w=1.7e-07 $l=1.20395e-06 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=1.835 $X2=1.385 $Y2=2.95
r82 2 18 400 $w=1.7e-07 $l=3.76298e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=1.835 $X2=1.385 $Y2=2.13
r83 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.95
r84 1 12 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_2%X 1 2 9 10 11 12 13 14 15 16 26 39
r25 40 51 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=0.842 $Y=2.252
+ $X2=0.842 $Y2=2.21
r26 39 49 0.633766 $w=1.73e-07 $l=1e-08 $layer=LI1_cond $X=0.722 $Y=2.035
+ $X2=0.722 $Y2=2.045
r27 16 46 3.47121 $w=4.13e-07 $l=1.25e-07 $layer=LI1_cond $X=0.842 $Y=2.775
+ $X2=0.842 $Y2=2.9
r28 15 16 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.842 $Y=2.405
+ $X2=0.842 $Y2=2.775
r29 15 40 4.24877 $w=4.13e-07 $l=1.53e-07 $layer=LI1_cond $X=0.842 $Y=2.405
+ $X2=0.842 $Y2=2.252
r30 14 51 3.55452 $w=4.13e-07 $l=1.28e-07 $layer=LI1_cond $X=0.842 $Y=2.082
+ $X2=0.842 $Y2=2.21
r31 14 49 4.97156 $w=4.13e-07 $l=3.7e-08 $layer=LI1_cond $X=0.842 $Y=2.082
+ $X2=0.842 $Y2=2.045
r32 14 39 2.40831 $w=1.73e-07 $l=3.8e-08 $layer=LI1_cond $X=0.722 $Y=1.997
+ $X2=0.722 $Y2=2.035
r33 13 14 21.041 $w=1.73e-07 $l=3.32e-07 $layer=LI1_cond $X=0.722 $Y=1.665
+ $X2=0.722 $Y2=1.997
r34 12 13 23.4494 $w=1.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=1.295
+ $X2=0.722 $Y2=1.665
r35 10 11 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.555
+ $X2=0.715 $Y2=0.925
r36 10 26 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=0.715 $Y=0.555
+ $X2=0.715 $Y2=0.42
r37 9 12 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=0.722 $Y=1.125
+ $X2=0.722 $Y2=1.295
r38 7 11 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=0.715 $Y=1.03
+ $X2=0.715 $Y2=0.925
r39 7 9 5.63364 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.715 $Y=1.03
+ $X2=0.715 $Y2=1.125
r40 2 51 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=0.77
+ $Y=1.835 $X2=0.91 $Y2=2.21
r41 2 46 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=0.77
+ $Y=1.835 $X2=0.91 $Y2=2.9
r42 1 26 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.245 $X2=0.715 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_2%A_342_367# 1 2 7 9 11 13 15
r25 13 20 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.925 $Y=2.225
+ $X2=2.925 $Y2=2.135
r26 13 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.925 $Y=2.225
+ $X2=2.925 $Y2=2.935
r27 12 18 4.57023 $w=1.8e-07 $l=1.48e-07 $layer=LI1_cond $X=2.015 $Y=2.135
+ $X2=1.867 $Y2=2.135
r28 11 20 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=2.135
+ $X2=2.925 $Y2=2.135
r29 11 12 45.904 $w=1.78e-07 $l=7.45e-07 $layer=LI1_cond $X=2.76 $Y=2.135
+ $X2=2.015 $Y2=2.135
r30 7 18 2.7792 $w=2.95e-07 $l=9e-08 $layer=LI1_cond $X=1.867 $Y=2.225 $X2=1.867
+ $Y2=2.135
r31 7 9 26.7601 $w=2.93e-07 $l=6.85e-07 $layer=LI1_cond $X=1.867 $Y=2.225
+ $X2=1.867 $Y2=2.91
r32 2 20 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.835 $X2=2.925 $Y2=2.13
r33 2 15 400 $w=1.7e-07 $l=1.1679e-06 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.835 $X2=2.925 $Y2=2.935
r34 1 18 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.835 $X2=1.85 $Y2=2.21
r35 1 9 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.835 $X2=1.85 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_2%VGND 1 2 3 10 12 16 19 20 21 23 36 37 44
r51 44 47 9.90781 $w=6.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.315 $Y=0
+ $X2=1.315 $Y2=0.555
r52 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r54 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 34 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r56 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r58 30 33 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r59 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 28 44 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.315
+ $Y2=0
r61 28 30 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.68
+ $Y2=0
r62 27 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r63 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r64 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 24 40 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.225
+ $Y2=0
r66 24 26 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.72
+ $Y2=0
r67 23 44 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.315
+ $Y2=0
r68 23 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.72
+ $Y2=0
r69 21 34 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r70 21 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r71 19 33 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.12
+ $Y2=0
r72 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.355
+ $Y2=0
r73 18 36 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.52 $Y=0 $X2=3.6
+ $Y2=0
r74 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.52 $Y=0 $X2=3.355
+ $Y2=0
r75 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.355 $Y2=0
r76 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.355 $Y=0.085
+ $X2=3.355 $Y2=0.39
r77 10 40 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=0.085
+ $X2=0.225 $Y2=0
r78 10 12 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.285 $Y=0.085
+ $X2=0.285 $Y2=0.39
r79 3 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.215
+ $Y=0.245 $X2=3.355 $Y2=0.39
r80 2 47 91 $w=1.7e-07 $l=6.15792e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.245 $X2=1.485 $Y2=0.555
r81 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.245 $X2=0.285 $Y2=0.39
.ends

