* File: sky130_fd_sc_lp__sdfxtp_lp.pxi.spice
* Created: Fri Aug 28 11:31:09 2020
* 
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_27_409# N_A_27_409#_M1032_s
+ N_A_27_409#_M1005_s N_A_27_409#_M1011_g N_A_27_409#_M1025_g
+ N_A_27_409#_c_228_n N_A_27_409#_c_229_n N_A_27_409#_c_238_n
+ N_A_27_409#_c_230_n N_A_27_409#_c_231_n N_A_27_409#_c_232_n
+ N_A_27_409#_c_233_n N_A_27_409#_c_234_n N_A_27_409#_c_235_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_27_409#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%D N_D_M1003_g N_D_M1000_g N_D_c_295_n
+ N_D_c_300_n D N_D_c_296_n N_D_c_297_n PM_SKY130_FD_SC_LP__SDFXTP_LP%D
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%SCE N_SCE_M1005_g N_SCE_M1032_g N_SCE_c_335_n
+ N_SCE_M1015_g N_SCE_c_337_n N_SCE_c_338_n N_SCE_M1034_g N_SCE_c_340_n
+ N_SCE_M1030_g SCE N_SCE_c_343_n PM_SKY130_FD_SC_LP__SDFXTP_LP%SCE
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%SCD N_SCD_M1019_g N_SCD_c_414_n N_SCD_M1014_g
+ N_SCD_c_419_n SCD SCD N_SCD_c_416_n PM_SKY130_FD_SC_LP__SDFXTP_LP%SCD
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%CLK N_CLK_M1018_g N_CLK_M1029_g N_CLK_M1020_g
+ CLK N_CLK_c_458_n PM_SKY130_FD_SC_LP__SDFXTP_LP%CLK
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1576_99# N_A_1576_99#_M1016_d
+ N_A_1576_99#_M1010_d N_A_1576_99#_M1036_d N_A_1576_99#_M1037_g
+ N_A_1576_99#_M1022_g N_A_1576_99#_c_497_n N_A_1576_99#_c_498_n
+ N_A_1576_99#_c_507_n N_A_1576_99#_c_508_n N_A_1576_99#_c_499_n
+ N_A_1576_99#_c_500_n N_A_1576_99#_c_501_n N_A_1576_99#_c_502_n
+ N_A_1576_99#_c_503_n N_A_1576_99#_c_504_n N_A_1576_99#_c_505_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1576_99#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1263_155# N_A_1263_155#_M1023_d
+ N_A_1263_155#_M1021_d N_A_1263_155#_M1028_g N_A_1263_155#_M1016_g
+ N_A_1263_155#_M1036_g N_A_1263_155#_c_594_n N_A_1263_155#_c_595_n
+ N_A_1263_155#_c_596_n N_A_1263_155#_c_601_n N_A_1263_155#_c_602_n
+ N_A_1263_155#_c_597_n N_A_1263_155#_c_598_n N_A_1263_155#_c_599_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1263_155#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_733_66# N_A_733_66#_M1018_s
+ N_A_733_66#_M1029_s N_A_733_66#_c_676_n N_A_733_66#_M1004_g
+ N_A_733_66#_M1012_g N_A_733_66#_M1027_g N_A_733_66#_c_679_n
+ N_A_733_66#_c_680_n N_A_733_66#_M1009_g N_A_733_66#_c_682_n
+ N_A_733_66#_M1007_g N_A_733_66#_c_684_n N_A_733_66#_c_685_n
+ N_A_733_66#_M1017_g N_A_733_66#_c_687_n N_A_733_66#_M1008_g
+ N_A_733_66#_c_688_n N_A_733_66#_c_689_n N_A_733_66#_c_690_n
+ N_A_733_66#_c_691_n N_A_733_66#_c_692_n N_A_733_66#_c_693_n
+ N_A_733_66#_c_694_n N_A_733_66#_c_695_n N_A_733_66#_c_703_n
+ N_A_733_66#_c_696_n N_A_733_66#_c_697_n N_A_733_66#_c_698_n
+ N_A_733_66#_c_699_n PM_SKY130_FD_SC_LP__SDFXTP_LP%A_733_66#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_998_347# N_A_998_347#_M1027_d
+ N_A_998_347#_M1012_d N_A_998_347#_c_849_n N_A_998_347#_c_842_n
+ N_A_998_347#_c_843_n N_A_998_347#_c_850_n N_A_998_347#_c_851_n
+ N_A_998_347#_c_844_n N_A_998_347#_M1023_g N_A_998_347#_M1021_g
+ N_A_998_347#_c_853_n N_A_998_347#_M1033_g N_A_998_347#_c_855_n
+ N_A_998_347#_M1010_g N_A_998_347#_c_857_n N_A_998_347#_c_858_n
+ N_A_998_347#_c_846_n N_A_998_347#_c_847_n N_A_998_347#_c_848_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_998_347#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_2148_185# N_A_2148_185#_M1013_d
+ N_A_2148_185#_M1031_d N_A_2148_185#_M1026_g N_A_2148_185#_M1001_g
+ N_A_2148_185#_c_947_n N_A_2148_185#_c_948_n N_A_2148_185#_M1002_g
+ N_A_2148_185#_M1006_g N_A_2148_185#_M1035_g N_A_2148_185#_c_952_n
+ N_A_2148_185#_c_953_n N_A_2148_185#_c_954_n N_A_2148_185#_c_955_n
+ N_A_2148_185#_c_956_n N_A_2148_185#_c_963_n N_A_2148_185#_c_957_n
+ N_A_2148_185#_c_958_n N_A_2148_185#_c_959_n N_A_2148_185#_c_960_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_2148_185#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1957_347# N_A_1957_347#_M1008_d
+ N_A_1957_347#_M1017_d N_A_1957_347#_c_1047_n N_A_1957_347#_M1031_g
+ N_A_1957_347#_M1024_g N_A_1957_347#_c_1049_n N_A_1957_347#_M1013_g
+ N_A_1957_347#_c_1057_n N_A_1957_347#_c_1051_n N_A_1957_347#_c_1052_n
+ N_A_1957_347#_c_1053_n N_A_1957_347#_c_1054_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1957_347#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%VPWR N_VPWR_M1005_d N_VPWR_M1030_d
+ N_VPWR_M1029_d N_VPWR_M1022_d N_VPWR_M1026_d N_VPWR_M1006_d N_VPWR_c_1130_n
+ N_VPWR_c_1131_n N_VPWR_c_1132_n N_VPWR_c_1133_n N_VPWR_c_1134_n
+ N_VPWR_c_1135_n N_VPWR_c_1136_n N_VPWR_c_1137_n N_VPWR_c_1138_n VPWR
+ N_VPWR_c_1139_n N_VPWR_c_1140_n N_VPWR_c_1141_n N_VPWR_c_1142_n
+ N_VPWR_c_1143_n N_VPWR_c_1144_n N_VPWR_c_1145_n N_VPWR_c_1146_n
+ N_VPWR_c_1129_n PM_SKY130_FD_SC_LP__SDFXTP_LP%VPWR
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_244_417# N_A_244_417#_M1011_s
+ N_A_244_417#_M1014_d N_A_244_417#_c_1237_n N_A_244_417#_c_1238_n
+ N_A_244_417#_c_1239_n N_A_244_417#_c_1240_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_244_417#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_351_417# N_A_351_417#_M1003_d
+ N_A_351_417#_M1009_d N_A_351_417#_M1011_d N_A_351_417#_M1021_s
+ N_A_351_417#_c_1284_n N_A_351_417#_c_1278_n N_A_351_417#_c_1279_n
+ N_A_351_417#_c_1280_n N_A_351_417#_c_1281_n N_A_351_417#_c_1287_n
+ N_A_351_417#_c_1282_n N_A_351_417#_c_1283_n N_A_351_417#_c_1307_n
+ N_A_351_417#_c_1288_n N_A_351_417#_c_1289_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_351_417#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%Q N_Q_M1002_s N_Q_M1006_s N_Q_c_1383_n Q Q Q
+ N_Q_c_1384_n PM_SKY130_FD_SC_LP__SDFXTP_LP%Q
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%VGND N_VGND_M1015_d N_VGND_M1019_d
+ N_VGND_M1020_d N_VGND_M1037_d N_VGND_M1001_d N_VGND_M1035_d N_VGND_c_1413_n
+ N_VGND_c_1414_n N_VGND_c_1415_n N_VGND_c_1416_n N_VGND_c_1417_n
+ N_VGND_c_1418_n N_VGND_c_1419_n N_VGND_c_1420_n N_VGND_c_1421_n VGND
+ N_VGND_c_1422_n N_VGND_c_1423_n N_VGND_c_1424_n N_VGND_c_1425_n
+ N_VGND_c_1426_n N_VGND_c_1427_n N_VGND_c_1428_n N_VGND_c_1429_n
+ N_VGND_c_1430_n N_VGND_c_1431_n PM_SKY130_FD_SC_LP__SDFXTP_LP%VGND
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1160_155# N_A_1160_155#_M1023_s
+ N_A_1160_155#_M1037_s N_A_1160_155#_c_1545_n N_A_1160_155#_c_1546_n
+ N_A_1160_155#_c_1547_n N_A_1160_155#_c_1548_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1160_155#
x_PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1910_155# N_A_1910_155#_M1008_s
+ N_A_1910_155#_M1001_s N_A_1910_155#_c_1581_n N_A_1910_155#_c_1582_n
+ N_A_1910_155#_c_1583_n N_A_1910_155#_c_1584_n
+ PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1910_155#
cc_1 VNB N_A_27_409#_c_228_n 0.0169966f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.165
cc_2 VNB N_A_27_409#_c_229_n 0.0224156f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.67
cc_3 VNB N_A_27_409#_c_230_n 0.034521f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.835
cc_4 VNB N_A_27_409#_c_231_n 0.0172128f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.19
cc_5 VNB N_A_27_409#_c_232_n 0.0234774f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.25
cc_6 VNB N_A_27_409#_c_233_n 0.0134272f $X=-0.19 $Y=-0.245 $X2=0.392 $Y2=1.25
cc_7 VNB N_A_27_409#_c_234_n 0.00668666f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.33
cc_8 VNB N_A_27_409#_c_235_n 0.0145799f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.33
cc_9 VNB N_D_M1003_g 0.0193139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_D_c_295_n 0.0186885f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.165
cc_11 VNB N_D_c_296_n 0.016334f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.67
cc_12 VNB N_D_c_297_n 0.00431482f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.835
cc_13 VNB N_SCE_M1032_g 0.0411412f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.835
cc_14 VNB N_SCE_c_335_n 0.00847643f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=2.585
cc_15 VNB N_SCE_M1015_g 0.0504344f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.33
cc_16 VNB N_SCE_c_337_n 0.112697f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.165
cc_17 VNB N_SCE_c_338_n 0.0126405f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.67
cc_18 VNB N_SCE_M1034_g 0.0327782f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.835
cc_19 VNB N_SCE_c_340_n 0.0127735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_SCE_M1030_g 0.0217626f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.19
cc_21 VNB SCE 9.34446e-19 $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.9
cc_22 VNB N_SCE_c_343_n 0.0163969f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.33
cc_23 VNB N_SCD_M1019_g 0.0286291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_SCD_c_414_n 0.0184588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB SCD 0.017832f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.835
cc_26 VNB N_SCD_c_416_n 0.0202686f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.835
cc_27 VNB N_CLK_M1018_g 0.0394111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_CLK_M1029_g 0.00329302f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.835
cc_29 VNB N_CLK_M1020_g 0.0295534f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.165
cc_30 VNB CLK 0.00284951f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.835
cc_31 VNB N_CLK_c_458_n 0.0434819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1576_99#_M1022_g 0.00451939f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.165
cc_33 VNB N_A_1576_99#_c_497_n 0.00659583f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.835
cc_34 VNB N_A_1576_99#_c_498_n 0.00480125f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.335
cc_35 VNB N_A_1576_99#_c_499_n 0.00463592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1576_99#_c_500_n 0.0240402f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.25
cc_37 VNB N_A_1576_99#_c_501_n 0.00913979f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.33
cc_38 VNB N_A_1576_99#_c_502_n 0.0267893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1576_99#_c_503_n 0.00350992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1576_99#_c_504_n 0.0108983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1576_99#_c_505_n 0.0172307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1263_155#_M1028_g 0.0197366f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=2.585
cc_43 VNB N_A_1263_155#_M1016_g 0.0186694f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.835
cc_44 VNB N_A_1263_155#_c_594_n 0.00240272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1263_155#_c_595_n 0.00427122f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.19
cc_46 VNB N_A_1263_155#_c_596_n 0.00534608f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.19
cc_47 VNB N_A_1263_155#_c_597_n 2.86565e-19 $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.33
cc_48 VNB N_A_1263_155#_c_598_n 0.00605958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1263_155#_c_599_n 0.0369929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_733_66#_c_676_n 0.0155006f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.835
cc_51 VNB N_A_733_66#_M1012_g 0.0017237f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.835
cc_52 VNB N_A_733_66#_M1027_g 0.0108826f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.835
cc_53 VNB N_A_733_66#_c_679_n 0.116644f $X=-0.19 $Y=-0.245 $X2=0.392 $Y2=1.165
cc_54 VNB N_A_733_66#_c_680_n 0.0113293f $X=-0.19 $Y=-0.245 $X2=0.392 $Y2=0.835
cc_55 VNB N_A_733_66#_M1009_g 0.0450639f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.335
cc_56 VNB N_A_733_66#_c_682_n 0.021289f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.19
cc_57 VNB N_A_733_66#_M1007_g 0.0203087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_733_66#_c_684_n 0.140572f $X=-0.19 $Y=-0.245 $X2=0.392 $Y2=1.25
cc_59 VNB N_A_733_66#_c_685_n 0.0656694f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.33
cc_60 VNB N_A_733_66#_M1017_g 0.0102111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_733_66#_c_687_n 0.013679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_733_66#_c_688_n 0.0268974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_733_66#_c_689_n 0.0141414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_733_66#_c_690_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_733_66#_c_691_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_733_66#_c_692_n 0.0502545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_733_66#_c_693_n 0.0141929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_733_66#_c_694_n 0.0337938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_733_66#_c_695_n 0.00777936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_733_66#_c_696_n 0.0201252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_733_66#_c_697_n 0.0125017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_733_66#_c_698_n 4.51335e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_733_66#_c_699_n 0.0253007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_998_347#_c_842_n 0.0446627f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=2.585
cc_75 VNB N_A_998_347#_c_843_n 0.0174909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_998_347#_c_844_n 0.0178618f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.835
cc_77 VNB N_A_998_347#_M1010_g 0.0319335f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.25
cc_78 VNB N_A_998_347#_c_846_n 0.0159125f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.33
cc_79 VNB N_A_998_347#_c_847_n 0.0121388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_998_347#_c_848_n 0.00564795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_2148_185#_M1026_g 0.021524f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=2.585
cc_82 VNB N_A_2148_185#_M1001_g 0.0252722f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.835
cc_83 VNB N_A_2148_185#_c_947_n 0.0175844f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.165
cc_84 VNB N_A_2148_185#_c_948_n 0.0221224f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.67
cc_85 VNB N_A_2148_185#_M1002_g 0.0259061f $X=-0.19 $Y=-0.245 $X2=0.392
+ $Y2=0.835
cc_86 VNB N_A_2148_185#_M1006_g 0.0545527f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.19
cc_87 VNB N_A_2148_185#_M1035_g 0.0274426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_2148_185#_c_952_n 0.0252184f $X=-0.19 $Y=-0.245 $X2=0.392 $Y2=1.25
cc_89 VNB N_A_2148_185#_c_953_n 0.0114002f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.33
cc_90 VNB N_A_2148_185#_c_954_n 0.00280285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2148_185#_c_955_n 0.0010781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2148_185#_c_956_n 0.0580959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2148_185#_c_957_n 0.00559263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2148_185#_c_958_n 0.024562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2148_185#_c_959_n 0.0533226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2148_185#_c_960_n 0.00766569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1957_347#_c_1047_n 0.0446278f $X=-0.19 $Y=-0.245 $X2=1.63
+ $Y2=1.835
cc_98 VNB N_A_1957_347#_M1024_g 0.0290511f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0.835
cc_99 VNB N_A_1957_347#_c_1049_n 0.0232461f $X=-0.19 $Y=-0.245 $X2=1.59
+ $Y2=1.165
cc_100 VNB N_A_1957_347#_M1013_g 0.0335999f $X=-0.19 $Y=-0.245 $X2=0.392
+ $Y2=0.835
cc_101 VNB N_A_1957_347#_c_1051_n 5.37725e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1957_347#_c_1052_n 0.0146304f $X=-0.19 $Y=-0.245 $X2=1.59
+ $Y2=1.25
cc_103 VNB N_A_1957_347#_c_1053_n 0.00181106f $X=-0.19 $Y=-0.245 $X2=1.59
+ $Y2=1.33
cc_104 VNB N_A_1957_347#_c_1054_n 0.00276933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VPWR_c_1129_n 0.581632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_351_417#_c_1278_n 0.00455364f $X=-0.19 $Y=-0.245 $X2=0.392
+ $Y2=1.165
cc_107 VNB N_A_351_417#_c_1279_n 0.00483827f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.335
cc_108 VNB N_A_351_417#_c_1280_n 0.0082733f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.19
cc_109 VNB N_A_351_417#_c_1281_n 0.00133203f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.19
cc_110 VNB N_A_351_417#_c_1282_n 0.00381761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_351_417#_c_1283_n 0.00323792f $X=-0.19 $Y=-0.245 $X2=1.59
+ $Y2=1.33
cc_112 VNB N_Q_c_1383_n 0.00888668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_Q_c_1384_n 0.013384f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.25
cc_114 VNB N_VGND_c_1413_n 0.0116153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1414_n 0.0216405f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.9
cc_116 VNB N_VGND_c_1415_n 0.00293489f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.25
cc_117 VNB N_VGND_c_1416_n 0.00879115f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=1.25
cc_118 VNB N_VGND_c_1417_n 0.0054388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1418_n 0.0118377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1419_n 0.0377882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1420_n 0.072687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1421_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1422_n 0.035397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1423_n 0.0477062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1424_n 0.0290432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1425_n 0.0823484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1426_n 0.0508558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1427_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1428_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1429_n 0.00555411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1430_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1431_n 0.725468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_1160_155#_c_1545_n 0.0167725f $X=-0.19 $Y=-0.245 $X2=1.63
+ $Y2=2.585
cc_134 VNB N_A_1160_155#_c_1546_n 0.0306959f $X=-0.19 $Y=-0.245 $X2=1.68
+ $Y2=1.165
cc_135 VNB N_A_1160_155#_c_1547_n 0.0044524f $X=-0.19 $Y=-0.245 $X2=1.68
+ $Y2=0.835
cc_136 VNB N_A_1160_155#_c_1548_n 0.00694917f $X=-0.19 $Y=-0.245 $X2=1.59
+ $Y2=1.165
cc_137 VNB N_A_1910_155#_c_1581_n 0.00823906f $X=-0.19 $Y=-0.245 $X2=1.63
+ $Y2=2.585
cc_138 VNB N_A_1910_155#_c_1582_n 0.0159726f $X=-0.19 $Y=-0.245 $X2=1.68
+ $Y2=1.165
cc_139 VNB N_A_1910_155#_c_1583_n 0.00379749f $X=-0.19 $Y=-0.245 $X2=1.68
+ $Y2=0.835
cc_140 VNB N_A_1910_155#_c_1584_n 0.0101557f $X=-0.19 $Y=-0.245 $X2=1.59
+ $Y2=1.165
cc_141 VPB N_A_27_409#_M1011_g 0.0402816f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.585
cc_142 VPB N_A_27_409#_c_229_n 9.02489e-19 $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.67
cc_143 VPB N_A_27_409#_c_238_n 0.0154498f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.835
cc_144 VPB N_A_27_409#_c_231_n 0.0601925f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=2.19
cc_145 VPB N_A_27_409#_c_234_n 8.2657e-19 $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.33
cc_146 VPB N_D_M1000_g 0.0274235f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=1.835
cc_147 VPB N_D_c_295_n 0.00436519f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.165
cc_148 VPB N_D_c_300_n 0.0134868f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=0.835
cc_149 VPB N_D_c_297_n 7.46703e-19 $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.835
cc_150 VPB N_SCE_M1005_g 0.0391252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_SCE_c_335_n 0.0147784f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.585
cc_152 VPB N_SCE_M1030_g 0.0384005f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.19
cc_153 VPB SCE 0.00192552f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=2.9
cc_154 VPB N_SCE_c_343_n 0.0247123f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.33
cc_155 VPB N_SCD_c_414_n 0.00625759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_SCD_M1014_g 0.0330381f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.585
cc_157 VPB N_SCD_c_419_n 0.0188891f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.165
cc_158 VPB SCD 0.00839715f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=0.835
cc_159 VPB N_CLK_M1029_g 0.030195f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=1.835
cc_160 VPB N_A_1576_99#_M1022_g 0.0252751f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.165
cc_161 VPB N_A_1576_99#_c_507_n 0.00394496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_1576_99#_c_508_n 0.00325268f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.25
cc_163 VPB N_A_1576_99#_c_504_n 0.00366358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_1263_155#_M1036_g 0.0279231f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.835
cc_165 VPB N_A_1263_155#_c_601_n 0.00264581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_1263_155#_c_602_n 0.0131922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_1263_155#_c_597_n 0.0016987f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.33
cc_168 VPB N_A_1263_155#_c_598_n 0.00186343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_1263_155#_c_599_n 0.0141725f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_733_66#_M1012_g 0.0295748f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=0.835
cc_171 VPB N_A_733_66#_M1007_g 0.0230911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_733_66#_M1017_g 0.0278438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_733_66#_c_703_n 0.00650044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_733_66#_c_698_n 0.00289943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_998_347#_c_849_n 0.0950106f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.585
cc_176 VPB N_A_998_347#_c_850_n 0.0873395f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.165
cc_177 VPB N_A_998_347#_c_851_n 0.012806f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=0.835
cc_178 VPB N_A_998_347#_M1021_g 0.0525443f $X=-0.19 $Y=1.655 $X2=0.392 $Y2=1.165
cc_179 VPB N_A_998_347#_c_853_n 0.253774f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.835
cc_180 VPB N_A_998_347#_M1033_g 0.0256516f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.9
cc_181 VPB N_A_998_347#_c_855_n 0.0128819f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=2.9
cc_182 VPB N_A_998_347#_M1010_g 0.0031546f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.25
cc_183 VPB N_A_998_347#_c_857_n 0.0189649f $X=-0.19 $Y=1.655 $X2=0.392 $Y2=1.25
cc_184 VPB N_A_998_347#_c_858_n 0.0124845f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.25
cc_185 VPB N_A_998_347#_c_847_n 0.0187143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_998_347#_c_848_n 0.0212566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_2148_185#_M1026_g 0.0271335f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.585
cc_188 VPB N_A_2148_185#_M1006_g 0.0477578f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.19
cc_189 VPB N_A_2148_185#_c_963_n 0.0282475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_2148_185#_c_957_n 0.00954435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_1957_347#_c_1047_n 0.00722543f $X=-0.19 $Y=1.655 $X2=1.63
+ $Y2=1.835
cc_192 VPB N_A_1957_347#_M1031_g 0.0311752f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.585
cc_193 VPB N_A_1957_347#_c_1057_n 0.00686499f $X=-0.19 $Y=1.655 $X2=0.24
+ $Y2=2.19
cc_194 VPB N_A_1957_347#_c_1052_n 0.0144188f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.25
cc_195 VPB N_A_1957_347#_c_1053_n 0.00365521f $X=-0.19 $Y=1.655 $X2=1.59
+ $Y2=1.33
cc_196 VPB N_A_1957_347#_c_1054_n 7.45669e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1130_n 0.0163446f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.19
cc_198 VPB N_VPWR_c_1131_n 7.46595e-19 $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.25
cc_199 VPB N_VPWR_c_1132_n 0.0229058f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.25
cc_200 VPB N_VPWR_c_1133_n 0.018503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1134_n 0.0159517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1135_n 0.012153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1136_n 0.0626402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1137_n 0.0466449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1138_n 0.0044842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1139_n 0.0388222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1140_n 0.101885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1141_n 0.0758525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1142_n 0.0616554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1143_n 0.0251504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1144_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1145_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1146_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1129_n 0.180934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_244_417#_c_1237_n 0.0136392f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.585
cc_216 VPB N_A_244_417#_c_1238_n 0.00317291f $X=-0.19 $Y=1.655 $X2=1.68
+ $Y2=0.835
cc_217 VPB N_A_244_417#_c_1239_n 0.0107853f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.835
cc_218 VPB N_A_244_417#_c_1240_n 0.00506195f $X=-0.19 $Y=1.655 $X2=0.392
+ $Y2=0.835
cc_219 VPB N_A_351_417#_c_1284_n 0.014634f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=0.835
cc_220 VPB N_A_351_417#_c_1278_n 0.00315441f $X=-0.19 $Y=1.655 $X2=0.392
+ $Y2=1.165
cc_221 VPB N_A_351_417#_c_1279_n 0.00553385f $X=-0.19 $Y=1.655 $X2=0.24
+ $Y2=1.335
cc_222 VPB N_A_351_417#_c_1287_n 0.019273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_351_417#_c_1288_n 0.0681701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_351_417#_c_1289_n 0.0376134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB Q 0.0253344f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=0.835
cc_226 VPB Q 0.0297894f $X=-0.19 $Y=1.655 $X2=1.59 $Y2=1.33
cc_227 VPB N_Q_c_1384_n 0.01163f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=1.25
cc_228 N_A_27_409#_c_228_n N_D_M1003_g 0.0380232f $X=1.59 $Y=1.165 $X2=0 $Y2=0
cc_229 N_A_27_409#_c_234_n N_D_M1003_g 3.1836e-19 $X=1.59 $Y=1.33 $X2=0 $Y2=0
cc_230 N_A_27_409#_M1011_g N_D_M1000_g 0.0495982f $X=1.63 $Y=2.585 $X2=0 $Y2=0
cc_231 N_A_27_409#_c_229_n N_D_c_295_n 0.013728f $X=1.59 $Y=1.67 $X2=0 $Y2=0
cc_232 N_A_27_409#_c_238_n N_D_c_300_n 0.013728f $X=1.59 $Y=1.835 $X2=0 $Y2=0
cc_233 N_A_27_409#_c_234_n N_D_c_296_n 0.00215095f $X=1.59 $Y=1.33 $X2=0 $Y2=0
cc_234 N_A_27_409#_c_235_n N_D_c_296_n 0.013728f $X=1.59 $Y=1.33 $X2=0 $Y2=0
cc_235 N_A_27_409#_c_229_n N_D_c_297_n 0.0020827f $X=1.59 $Y=1.67 $X2=0 $Y2=0
cc_236 N_A_27_409#_c_234_n N_D_c_297_n 0.0396062f $X=1.59 $Y=1.33 $X2=0 $Y2=0
cc_237 N_A_27_409#_c_230_n N_SCE_M1032_g 0.0138875f $X=0.505 $Y=0.835 $X2=0
+ $Y2=0
cc_238 N_A_27_409#_c_231_n N_SCE_M1032_g 0.00570404f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_239 N_A_27_409#_c_232_n N_SCE_M1032_g 0.0107693f $X=1.425 $Y=1.25 $X2=0 $Y2=0
cc_240 N_A_27_409#_c_233_n N_SCE_M1032_g 0.00464376f $X=0.392 $Y=1.25 $X2=0
+ $Y2=0
cc_241 N_A_27_409#_c_229_n N_SCE_c_335_n 0.0140381f $X=1.59 $Y=1.67 $X2=0 $Y2=0
cc_242 N_A_27_409#_c_232_n N_SCE_c_335_n 0.00203214f $X=1.425 $Y=1.25 $X2=0
+ $Y2=0
cc_243 N_A_27_409#_c_228_n N_SCE_M1015_g 0.0126314f $X=1.59 $Y=1.165 $X2=0 $Y2=0
cc_244 N_A_27_409#_c_230_n N_SCE_M1015_g 0.00195403f $X=0.505 $Y=0.835 $X2=0
+ $Y2=0
cc_245 N_A_27_409#_c_232_n N_SCE_M1015_g 0.0177902f $X=1.425 $Y=1.25 $X2=0 $Y2=0
cc_246 N_A_27_409#_c_234_n N_SCE_M1015_g 0.00190179f $X=1.59 $Y=1.33 $X2=0 $Y2=0
cc_247 N_A_27_409#_c_235_n N_SCE_M1015_g 0.0140381f $X=1.59 $Y=1.33 $X2=0 $Y2=0
cc_248 N_A_27_409#_c_228_n N_SCE_c_337_n 0.00907339f $X=1.59 $Y=1.165 $X2=0
+ $Y2=0
cc_249 N_A_27_409#_c_229_n SCE 0.00106622f $X=1.59 $Y=1.67 $X2=0 $Y2=0
cc_250 N_A_27_409#_c_231_n SCE 0.0244713f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_251 N_A_27_409#_c_232_n SCE 0.0142514f $X=1.425 $Y=1.25 $X2=0 $Y2=0
cc_252 N_A_27_409#_c_233_n SCE 0.00994925f $X=0.392 $Y=1.25 $X2=0 $Y2=0
cc_253 N_A_27_409#_c_234_n SCE 0.0091394f $X=1.59 $Y=1.33 $X2=0 $Y2=0
cc_254 N_A_27_409#_M1011_g N_SCE_c_343_n 2.12182e-19 $X=1.63 $Y=2.585 $X2=0
+ $Y2=0
cc_255 N_A_27_409#_c_229_n N_SCE_c_343_n 0.00329978f $X=1.59 $Y=1.67 $X2=0 $Y2=0
cc_256 N_A_27_409#_c_231_n N_SCE_c_343_n 0.0183672f $X=0.28 $Y=2.19 $X2=0 $Y2=0
cc_257 N_A_27_409#_c_233_n N_SCE_c_343_n 0.00679978f $X=0.392 $Y=1.25 $X2=0
+ $Y2=0
cc_258 N_A_27_409#_c_234_n N_SCE_c_343_n 7.6928e-19 $X=1.59 $Y=1.33 $X2=0 $Y2=0
cc_259 N_A_27_409#_M1011_g N_VPWR_c_1130_n 0.00575148f $X=1.63 $Y=2.585 $X2=0
+ $Y2=0
cc_260 N_A_27_409#_c_231_n N_VPWR_c_1130_n 0.0272606f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_261 N_A_27_409#_M1011_g N_VPWR_c_1137_n 0.00689754f $X=1.63 $Y=2.585 $X2=0
+ $Y2=0
cc_262 N_A_27_409#_c_231_n N_VPWR_c_1143_n 0.0167213f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_263 N_A_27_409#_M1011_g N_VPWR_c_1129_n 0.0101052f $X=1.63 $Y=2.585 $X2=0
+ $Y2=0
cc_264 N_A_27_409#_c_231_n N_VPWR_c_1129_n 0.0095959f $X=0.28 $Y=2.19 $X2=0
+ $Y2=0
cc_265 N_A_27_409#_M1011_g N_A_244_417#_c_1237_n 0.0103575f $X=1.63 $Y=2.585
+ $X2=0 $Y2=0
cc_266 N_A_27_409#_c_238_n N_A_244_417#_c_1237_n 5.96864e-19 $X=1.59 $Y=1.835
+ $X2=0 $Y2=0
cc_267 N_A_27_409#_c_234_n N_A_244_417#_c_1237_n 0.00719112f $X=1.59 $Y=1.33
+ $X2=0 $Y2=0
cc_268 N_A_27_409#_M1011_g N_A_244_417#_c_1238_n 0.0168096f $X=1.63 $Y=2.585
+ $X2=0 $Y2=0
cc_269 N_A_27_409#_c_234_n N_A_244_417#_c_1238_n 0.00480834f $X=1.59 $Y=1.33
+ $X2=0 $Y2=0
cc_270 N_A_27_409#_M1011_g N_A_244_417#_c_1240_n 0.0125111f $X=1.63 $Y=2.585
+ $X2=0 $Y2=0
cc_271 N_A_27_409#_M1011_g N_A_351_417#_c_1284_n 0.00560657f $X=1.63 $Y=2.585
+ $X2=0 $Y2=0
cc_272 N_A_27_409#_c_234_n N_A_351_417#_c_1284_n 0.00147549f $X=1.59 $Y=1.33
+ $X2=0 $Y2=0
cc_273 N_A_27_409#_c_228_n N_VGND_c_1413_n 0.013096f $X=1.59 $Y=1.165 $X2=0
+ $Y2=0
cc_274 N_A_27_409#_c_230_n N_VGND_c_1413_n 0.0125366f $X=0.505 $Y=0.835 $X2=0
+ $Y2=0
cc_275 N_A_27_409#_c_232_n N_VGND_c_1413_n 0.0182523f $X=1.425 $Y=1.25 $X2=0
+ $Y2=0
cc_276 N_A_27_409#_c_234_n N_VGND_c_1413_n 0.00534387f $X=1.59 $Y=1.33 $X2=0
+ $Y2=0
cc_277 N_A_27_409#_c_235_n N_VGND_c_1413_n 4.97464e-19 $X=1.59 $Y=1.33 $X2=0
+ $Y2=0
cc_278 N_A_27_409#_c_230_n N_VGND_c_1422_n 0.0118767f $X=0.505 $Y=0.835 $X2=0
+ $Y2=0
cc_279 N_A_27_409#_c_228_n N_VGND_c_1431_n 9.49986e-19 $X=1.59 $Y=1.165 $X2=0
+ $Y2=0
cc_280 N_A_27_409#_c_230_n N_VGND_c_1431_n 0.017127f $X=0.505 $Y=0.835 $X2=0
+ $Y2=0
cc_281 N_D_M1003_g N_SCE_c_337_n 0.00907339f $X=2.07 $Y=0.835 $X2=0 $Y2=0
cc_282 N_D_M1003_g N_SCE_M1034_g 0.0156566f $X=2.07 $Y=0.835 $X2=0 $Y2=0
cc_283 N_D_c_296_n N_SCE_c_340_n 0.0208967f $X=2.13 $Y=1.38 $X2=0 $Y2=0
cc_284 N_D_c_297_n N_SCE_c_340_n 7.93125e-19 $X=2.13 $Y=1.38 $X2=0 $Y2=0
cc_285 N_D_M1000_g N_SCE_M1030_g 0.0846943f $X=2.16 $Y=2.585 $X2=0 $Y2=0
cc_286 N_D_c_295_n N_SCE_M1030_g 0.0208967f $X=2.13 $Y=1.72 $X2=0 $Y2=0
cc_287 N_D_M1000_g N_VPWR_c_1131_n 0.00189839f $X=2.16 $Y=2.585 $X2=0 $Y2=0
cc_288 N_D_M1000_g N_VPWR_c_1137_n 0.00699368f $X=2.16 $Y=2.585 $X2=0 $Y2=0
cc_289 N_D_M1000_g N_VPWR_c_1129_n 0.00878302f $X=2.16 $Y=2.585 $X2=0 $Y2=0
cc_290 N_D_M1000_g N_A_244_417#_c_1237_n 6.31982e-19 $X=2.16 $Y=2.585 $X2=0
+ $Y2=0
cc_291 N_D_M1000_g N_A_244_417#_c_1238_n 0.0168827f $X=2.16 $Y=2.585 $X2=0 $Y2=0
cc_292 N_D_M1000_g N_A_244_417#_c_1240_n 0.00167569f $X=2.16 $Y=2.585 $X2=0
+ $Y2=0
cc_293 N_D_M1000_g N_A_351_417#_c_1284_n 0.0158567f $X=2.16 $Y=2.585 $X2=0 $Y2=0
cc_294 N_D_c_300_n N_A_351_417#_c_1284_n 5.5436e-19 $X=2.13 $Y=1.885 $X2=0 $Y2=0
cc_295 N_D_c_297_n N_A_351_417#_c_1284_n 0.0248611f $X=2.13 $Y=1.38 $X2=0 $Y2=0
cc_296 N_D_M1003_g N_A_351_417#_c_1278_n 0.00302497f $X=2.07 $Y=0.835 $X2=0
+ $Y2=0
cc_297 N_D_M1000_g N_A_351_417#_c_1278_n 0.00355667f $X=2.16 $Y=2.585 $X2=0
+ $Y2=0
cc_298 N_D_c_296_n N_A_351_417#_c_1278_n 0.00353574f $X=2.13 $Y=1.38 $X2=0 $Y2=0
cc_299 N_D_c_297_n N_A_351_417#_c_1278_n 0.0481605f $X=2.13 $Y=1.38 $X2=0 $Y2=0
cc_300 N_D_M1003_g N_A_351_417#_c_1283_n 0.00268596f $X=2.07 $Y=0.835 $X2=0
+ $Y2=0
cc_301 N_D_c_296_n N_A_351_417#_c_1283_n 6.90803e-19 $X=2.13 $Y=1.38 $X2=0 $Y2=0
cc_302 N_D_c_297_n N_A_351_417#_c_1283_n 0.00746632f $X=2.13 $Y=1.38 $X2=0 $Y2=0
cc_303 N_D_M1003_g N_VGND_c_1431_n 9.49986e-19 $X=2.07 $Y=0.835 $X2=0 $Y2=0
cc_304 N_SCE_M1034_g N_SCD_M1019_g 0.0227131f $X=2.58 $Y=0.835 $X2=0 $Y2=0
cc_305 N_SCE_c_340_n N_SCD_M1019_g 0.0246635f $X=2.63 $Y=1.245 $X2=0 $Y2=0
cc_306 N_SCE_M1030_g N_SCD_c_414_n 0.0246635f $X=2.63 $Y=2.585 $X2=0 $Y2=0
cc_307 N_SCE_M1030_g N_SCD_M1014_g 0.0464731f $X=2.63 $Y=2.585 $X2=0 $Y2=0
cc_308 N_SCE_M1030_g SCD 0.00223867f $X=2.63 $Y=2.585 $X2=0 $Y2=0
cc_309 N_SCE_M1005_g N_VPWR_c_1130_n 0.0231779f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_310 N_SCE_c_335_n N_VPWR_c_1130_n 0.0035377f $X=1.035 $Y=1.59 $X2=0 $Y2=0
cc_311 SCE N_VPWR_c_1130_n 0.0183937f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_312 N_SCE_c_343_n N_VPWR_c_1130_n 0.00158396f $X=0.875 $Y=1.68 $X2=0 $Y2=0
cc_313 N_SCE_M1030_g N_VPWR_c_1131_n 0.00974128f $X=2.63 $Y=2.585 $X2=0 $Y2=0
cc_314 N_SCE_M1030_g N_VPWR_c_1137_n 0.00628722f $X=2.63 $Y=2.585 $X2=0 $Y2=0
cc_315 N_SCE_M1005_g N_VPWR_c_1143_n 0.00802402f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_316 N_SCE_M1005_g N_VPWR_c_1129_n 0.0149742f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_317 N_SCE_M1030_g N_VPWR_c_1129_n 0.00697167f $X=2.63 $Y=2.585 $X2=0 $Y2=0
cc_318 N_SCE_M1030_g N_A_244_417#_c_1238_n 0.0166126f $X=2.63 $Y=2.585 $X2=0
+ $Y2=0
cc_319 N_SCE_M1030_g N_A_244_417#_c_1239_n 5.47451e-19 $X=2.63 $Y=2.585 $X2=0
+ $Y2=0
cc_320 N_SCE_M1005_g N_A_244_417#_c_1240_n 7.10786e-19 $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_321 N_SCE_M1034_g N_A_351_417#_c_1278_n 0.00304023f $X=2.58 $Y=0.835 $X2=0
+ $Y2=0
cc_322 N_SCE_c_340_n N_A_351_417#_c_1278_n 0.00394799f $X=2.63 $Y=1.245 $X2=0
+ $Y2=0
cc_323 N_SCE_M1030_g N_A_351_417#_c_1278_n 0.0223309f $X=2.63 $Y=2.585 $X2=0
+ $Y2=0
cc_324 N_SCE_c_337_n N_A_351_417#_c_1283_n 0.00412283f $X=2.505 $Y=0.18 $X2=0
+ $Y2=0
cc_325 N_SCE_M1034_g N_A_351_417#_c_1283_n 0.0140781f $X=2.58 $Y=0.835 $X2=0
+ $Y2=0
cc_326 N_SCE_M1030_g N_A_351_417#_c_1307_n 0.00950797f $X=2.63 $Y=2.585 $X2=0
+ $Y2=0
cc_327 N_SCE_M1030_g N_A_351_417#_c_1288_n 0.0100578f $X=2.63 $Y=2.585 $X2=0
+ $Y2=0
cc_328 N_SCE_M1032_g N_VGND_c_1413_n 0.00162086f $X=0.72 $Y=0.835 $X2=0 $Y2=0
cc_329 N_SCE_M1015_g N_VGND_c_1413_n 0.0255268f $X=1.11 $Y=0.835 $X2=0 $Y2=0
cc_330 N_SCE_c_337_n N_VGND_c_1413_n 0.0187754f $X=2.505 $Y=0.18 $X2=0 $Y2=0
cc_331 N_SCE_c_338_n N_VGND_c_1413_n 0.00388727f $X=1.185 $Y=0.18 $X2=0 $Y2=0
cc_332 N_SCE_c_337_n N_VGND_c_1414_n 0.00978633f $X=2.505 $Y=0.18 $X2=0 $Y2=0
cc_333 N_SCE_M1034_g N_VGND_c_1414_n 0.00185483f $X=2.58 $Y=0.835 $X2=0 $Y2=0
cc_334 N_SCE_M1032_g N_VGND_c_1422_n 0.00399929f $X=0.72 $Y=0.835 $X2=0 $Y2=0
cc_335 N_SCE_c_338_n N_VGND_c_1422_n 0.00486043f $X=1.185 $Y=0.18 $X2=0 $Y2=0
cc_336 N_SCE_c_337_n N_VGND_c_1423_n 0.0370899f $X=2.505 $Y=0.18 $X2=0 $Y2=0
cc_337 N_SCE_M1032_g N_VGND_c_1431_n 0.00469432f $X=0.72 $Y=0.835 $X2=0 $Y2=0
cc_338 N_SCE_c_337_n N_VGND_c_1431_n 0.0470752f $X=2.505 $Y=0.18 $X2=0 $Y2=0
cc_339 N_SCE_c_338_n N_VGND_c_1431_n 0.00983503f $X=1.185 $Y=0.18 $X2=0 $Y2=0
cc_340 SCD N_CLK_M1029_g 0.00671113f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_341 SCD CLK 0.0175443f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_342 N_SCD_c_416_n CLK 2.01561e-19 $X=3.17 $Y=1.41 $X2=0 $Y2=0
cc_343 SCD N_CLK_c_458_n 0.0029648f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_344 N_SCD_c_416_n N_CLK_c_458_n 0.00350019f $X=3.17 $Y=1.41 $X2=0 $Y2=0
cc_345 N_SCD_M1019_g N_A_733_66#_c_695_n 8.92906e-19 $X=3.04 $Y=0.835 $X2=0
+ $Y2=0
cc_346 N_SCD_c_414_n N_A_733_66#_c_703_n 7.20184e-19 $X=3.15 $Y=1.73 $X2=0 $Y2=0
cc_347 N_SCD_M1014_g N_A_733_66#_c_703_n 0.00158703f $X=3.16 $Y=2.585 $X2=0
+ $Y2=0
cc_348 SCD N_A_733_66#_c_703_n 0.0171954f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_349 SCD N_A_733_66#_c_697_n 0.00505442f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_350 N_SCD_M1014_g N_VPWR_c_1131_n 0.0098582f $X=3.16 $Y=2.585 $X2=0 $Y2=0
cc_351 N_SCD_M1014_g N_VPWR_c_1139_n 0.00619108f $X=3.16 $Y=2.585 $X2=0 $Y2=0
cc_352 N_SCD_M1014_g N_VPWR_c_1129_n 0.00830296f $X=3.16 $Y=2.585 $X2=0 $Y2=0
cc_353 N_SCD_M1014_g N_A_244_417#_c_1238_n 0.0161244f $X=3.16 $Y=2.585 $X2=0
+ $Y2=0
cc_354 N_SCD_M1014_g N_A_244_417#_c_1239_n 0.00908033f $X=3.16 $Y=2.585 $X2=0
+ $Y2=0
cc_355 N_SCD_M1019_g N_A_351_417#_c_1278_n 0.00316203f $X=3.04 $Y=0.835 $X2=0
+ $Y2=0
cc_356 N_SCD_M1014_g N_A_351_417#_c_1278_n 7.95258e-19 $X=3.16 $Y=2.585 $X2=0
+ $Y2=0
cc_357 SCD N_A_351_417#_c_1278_n 0.0278453f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_358 N_SCD_M1019_g N_A_351_417#_c_1283_n 0.00154665f $X=3.04 $Y=0.835 $X2=0
+ $Y2=0
cc_359 N_SCD_M1014_g N_A_351_417#_c_1307_n 4.72088e-19 $X=3.16 $Y=2.585 $X2=0
+ $Y2=0
cc_360 N_SCD_M1014_g N_A_351_417#_c_1288_n 0.0176685f $X=3.16 $Y=2.585 $X2=0
+ $Y2=0
cc_361 N_SCD_c_419_n N_A_351_417#_c_1288_n 0.00177823f $X=3.15 $Y=1.915 $X2=0
+ $Y2=0
cc_362 SCD N_A_351_417#_c_1288_n 0.0414625f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_363 N_SCD_M1019_g N_VGND_c_1414_n 0.0140026f $X=3.04 $Y=0.835 $X2=0 $Y2=0
cc_364 SCD N_VGND_c_1414_n 0.0281216f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_365 N_SCD_c_416_n N_VGND_c_1414_n 0.0059387f $X=3.17 $Y=1.41 $X2=0 $Y2=0
cc_366 N_SCD_M1019_g N_VGND_c_1423_n 0.00345209f $X=3.04 $Y=0.835 $X2=0 $Y2=0
cc_367 N_SCD_M1019_g N_VGND_c_1431_n 0.00394323f $X=3.04 $Y=0.835 $X2=0 $Y2=0
cc_368 N_CLK_M1020_g N_A_733_66#_c_676_n 0.0150576f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_369 N_CLK_M1029_g N_A_733_66#_M1012_g 0.0451631f $X=4.335 $Y=2.235 $X2=0
+ $Y2=0
cc_370 N_CLK_M1020_g N_A_733_66#_c_688_n 0.0108173f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_371 N_CLK_M1029_g N_A_733_66#_c_689_n 0.0108173f $X=4.335 $Y=2.235 $X2=0
+ $Y2=0
cc_372 N_CLK_M1018_g N_A_733_66#_c_695_n 0.0113373f $X=4.025 $Y=0.54 $X2=0 $Y2=0
cc_373 N_CLK_M1020_g N_A_733_66#_c_695_n 0.0018251f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_374 N_CLK_M1029_g N_A_733_66#_c_703_n 0.0214107f $X=4.335 $Y=2.235 $X2=0
+ $Y2=0
cc_375 CLK N_A_733_66#_c_703_n 0.0219514f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_376 N_CLK_c_458_n N_A_733_66#_c_703_n 0.00179859f $X=4.385 $Y=1.345 $X2=0
+ $Y2=0
cc_377 N_CLK_M1018_g N_A_733_66#_c_696_n 0.00808961f $X=4.025 $Y=0.54 $X2=0
+ $Y2=0
cc_378 N_CLK_M1020_g N_A_733_66#_c_696_n 0.0230306f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_379 CLK N_A_733_66#_c_696_n 0.0476895f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_380 N_CLK_c_458_n N_A_733_66#_c_696_n 2.07958e-19 $X=4.385 $Y=1.345 $X2=0
+ $Y2=0
cc_381 N_CLK_M1018_g N_A_733_66#_c_697_n 0.00417744f $X=4.025 $Y=0.54 $X2=0
+ $Y2=0
cc_382 CLK N_A_733_66#_c_697_n 0.00184056f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_383 N_CLK_c_458_n N_A_733_66#_c_698_n 0.00729993f $X=4.385 $Y=1.345 $X2=0
+ $Y2=0
cc_384 CLK N_A_733_66#_c_699_n 2.15138e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_385 N_CLK_c_458_n N_A_733_66#_c_699_n 0.0108173f $X=4.385 $Y=1.345 $X2=0
+ $Y2=0
cc_386 N_CLK_M1029_g N_VPWR_c_1132_n 0.0184641f $X=4.335 $Y=2.235 $X2=0 $Y2=0
cc_387 N_CLK_M1029_g N_VPWR_c_1139_n 0.00646289f $X=4.335 $Y=2.235 $X2=0 $Y2=0
cc_388 N_CLK_M1029_g N_VPWR_c_1129_n 0.00719887f $X=4.335 $Y=2.235 $X2=0 $Y2=0
cc_389 N_CLK_M1029_g N_A_244_417#_c_1238_n 0.00460716f $X=4.335 $Y=2.235 $X2=0
+ $Y2=0
cc_390 N_CLK_M1029_g N_A_244_417#_c_1239_n 0.0046584f $X=4.335 $Y=2.235 $X2=0
+ $Y2=0
cc_391 N_CLK_M1029_g N_A_351_417#_c_1288_n 0.0234019f $X=4.335 $Y=2.235 $X2=0
+ $Y2=0
cc_392 N_CLK_M1018_g N_VGND_c_1414_n 0.00583836f $X=4.025 $Y=0.54 $X2=0 $Y2=0
cc_393 N_CLK_M1018_g N_VGND_c_1415_n 0.00163126f $X=4.025 $Y=0.54 $X2=0 $Y2=0
cc_394 N_CLK_M1020_g N_VGND_c_1415_n 0.00983975f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_395 N_CLK_M1018_g N_VGND_c_1424_n 0.0046526f $X=4.025 $Y=0.54 $X2=0 $Y2=0
cc_396 N_CLK_M1020_g N_VGND_c_1424_n 0.00411131f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_397 N_CLK_M1018_g N_VGND_c_1431_n 0.00553875f $X=4.025 $Y=0.54 $X2=0 $Y2=0
cc_398 N_CLK_M1020_g N_VGND_c_1431_n 0.00401821f $X=4.385 $Y=0.54 $X2=0 $Y2=0
cc_399 N_A_1576_99#_c_497_n N_A_1263_155#_M1028_g 0.0114317f $X=8.945 $Y=0.98
+ $X2=0 $Y2=0
cc_400 N_A_1576_99#_c_498_n N_A_1263_155#_M1028_g 0.00152347f $X=9.11 $Y=0.835
+ $X2=0 $Y2=0
cc_401 N_A_1576_99#_c_501_n N_A_1263_155#_M1028_g 0.00340622f $X=8.045 $Y=0.98
+ $X2=0 $Y2=0
cc_402 N_A_1576_99#_c_502_n N_A_1263_155#_M1028_g 0.0170772f $X=8.045 $Y=1.32
+ $X2=0 $Y2=0
cc_403 N_A_1576_99#_c_505_n N_A_1263_155#_M1028_g 0.0147763f $X=8.045 $Y=1.155
+ $X2=0 $Y2=0
cc_404 N_A_1576_99#_c_497_n N_A_1263_155#_M1016_g 0.011364f $X=8.945 $Y=0.98
+ $X2=0 $Y2=0
cc_405 N_A_1576_99#_c_498_n N_A_1263_155#_M1016_g 0.00883554f $X=9.11 $Y=0.835
+ $X2=0 $Y2=0
cc_406 N_A_1576_99#_c_503_n N_A_1263_155#_M1016_g 0.00205768f $X=9.11 $Y=0.98
+ $X2=0 $Y2=0
cc_407 N_A_1576_99#_c_504_n N_A_1263_155#_M1016_g 0.00401245f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_408 N_A_1576_99#_M1022_g N_A_1263_155#_M1036_g 0.0115593f $X=8.005 $Y=2.235
+ $X2=0 $Y2=0
cc_409 N_A_1576_99#_c_507_n N_A_1263_155#_M1036_g 0.00325853f $X=9.27 $Y=1.88
+ $X2=0 $Y2=0
cc_410 N_A_1576_99#_M1022_g N_A_1263_155#_c_602_n 0.0229662f $X=8.005 $Y=2.235
+ $X2=0 $Y2=0
cc_411 N_A_1576_99#_c_497_n N_A_1263_155#_c_602_n 0.00780235f $X=8.945 $Y=0.98
+ $X2=0 $Y2=0
cc_412 N_A_1576_99#_c_501_n N_A_1263_155#_c_602_n 0.0234901f $X=8.045 $Y=0.98
+ $X2=0 $Y2=0
cc_413 N_A_1576_99#_c_502_n N_A_1263_155#_c_602_n 5.56982e-19 $X=8.045 $Y=1.32
+ $X2=0 $Y2=0
cc_414 N_A_1576_99#_c_504_n N_A_1263_155#_c_602_n 0.00380683f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_415 N_A_1576_99#_M1022_g N_A_1263_155#_c_597_n 0.00263657f $X=8.005 $Y=2.235
+ $X2=0 $Y2=0
cc_416 N_A_1576_99#_c_497_n N_A_1263_155#_c_597_n 0.0242553f $X=8.945 $Y=0.98
+ $X2=0 $Y2=0
cc_417 N_A_1576_99#_c_501_n N_A_1263_155#_c_597_n 0.0132832f $X=8.045 $Y=0.98
+ $X2=0 $Y2=0
cc_418 N_A_1576_99#_c_502_n N_A_1263_155#_c_597_n 3.07663e-19 $X=8.045 $Y=1.32
+ $X2=0 $Y2=0
cc_419 N_A_1576_99#_c_504_n N_A_1263_155#_c_597_n 0.0202502f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_420 N_A_1576_99#_M1022_g N_A_1263_155#_c_598_n 0.00481573f $X=8.005 $Y=2.235
+ $X2=0 $Y2=0
cc_421 N_A_1576_99#_c_501_n N_A_1263_155#_c_598_n 0.00398664f $X=8.045 $Y=0.98
+ $X2=0 $Y2=0
cc_422 N_A_1576_99#_M1022_g N_A_1263_155#_c_599_n 0.00393945f $X=8.005 $Y=2.235
+ $X2=0 $Y2=0
cc_423 N_A_1576_99#_c_497_n N_A_1263_155#_c_599_n 2.08868e-19 $X=8.945 $Y=0.98
+ $X2=0 $Y2=0
cc_424 N_A_1576_99#_c_503_n N_A_1263_155#_c_599_n 0.00550457f $X=9.11 $Y=0.98
+ $X2=0 $Y2=0
cc_425 N_A_1576_99#_c_504_n N_A_1263_155#_c_599_n 0.00325853f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_426 N_A_1576_99#_c_502_n N_A_733_66#_M1007_g 0.0481599f $X=8.045 $Y=1.32
+ $X2=0 $Y2=0
cc_427 N_A_1576_99#_c_497_n N_A_733_66#_c_684_n 0.0046157f $X=8.945 $Y=0.98
+ $X2=0 $Y2=0
cc_428 N_A_1576_99#_c_499_n N_A_733_66#_c_684_n 0.00674097f $X=9.275 $Y=0.35
+ $X2=0 $Y2=0
cc_429 N_A_1576_99#_c_501_n N_A_733_66#_c_684_n 4.00292e-19 $X=8.045 $Y=0.98
+ $X2=0 $Y2=0
cc_430 N_A_1576_99#_c_505_n N_A_733_66#_c_684_n 0.00907339f $X=8.045 $Y=1.155
+ $X2=0 $Y2=0
cc_431 N_A_1576_99#_c_498_n N_A_733_66#_c_685_n 0.00867788f $X=9.11 $Y=0.835
+ $X2=0 $Y2=0
cc_432 N_A_1576_99#_c_500_n N_A_733_66#_c_685_n 0.0179839f $X=10.52 $Y=0.35
+ $X2=0 $Y2=0
cc_433 N_A_1576_99#_c_503_n N_A_733_66#_c_685_n 0.00184673f $X=9.11 $Y=0.98
+ $X2=0 $Y2=0
cc_434 N_A_1576_99#_c_504_n N_A_733_66#_c_685_n 0.00422154f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_435 N_A_1576_99#_c_507_n N_A_733_66#_M1017_g 0.013319f $X=9.27 $Y=1.88 $X2=0
+ $Y2=0
cc_436 N_A_1576_99#_c_504_n N_A_733_66#_M1017_g 0.00300278f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_437 N_A_1576_99#_c_500_n N_A_733_66#_c_687_n 9.5131e-19 $X=10.52 $Y=0.35
+ $X2=0 $Y2=0
cc_438 N_A_1576_99#_c_505_n N_A_733_66#_c_692_n 0.0116667f $X=8.045 $Y=1.155
+ $X2=0 $Y2=0
cc_439 N_A_1576_99#_c_501_n N_A_733_66#_c_693_n 0.00183507f $X=8.045 $Y=0.98
+ $X2=0 $Y2=0
cc_440 N_A_1576_99#_c_505_n N_A_733_66#_c_693_n 0.0481599f $X=8.045 $Y=1.155
+ $X2=0 $Y2=0
cc_441 N_A_1576_99#_c_507_n N_A_733_66#_c_694_n 0.00461428f $X=9.27 $Y=1.88
+ $X2=0 $Y2=0
cc_442 N_A_1576_99#_M1022_g N_A_998_347#_c_853_n 0.0172549f $X=8.005 $Y=2.235
+ $X2=0 $Y2=0
cc_443 N_A_1576_99#_c_508_n N_A_998_347#_c_853_n 0.00666278f $X=9.27 $Y=2.59
+ $X2=0 $Y2=0
cc_444 N_A_1576_99#_c_500_n N_A_998_347#_M1010_g 9.5131e-19 $X=10.52 $Y=0.35
+ $X2=0 $Y2=0
cc_445 N_A_1576_99#_c_500_n N_A_2148_185#_M1001_g 0.00121906f $X=10.52 $Y=0.35
+ $X2=0 $Y2=0
cc_446 N_A_1576_99#_c_507_n N_A_1957_347#_c_1057_n 0.0228766f $X=9.27 $Y=1.88
+ $X2=0 $Y2=0
cc_447 N_A_1576_99#_c_504_n N_A_1957_347#_c_1057_n 0.00235193f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_448 N_A_1576_99#_c_504_n N_A_1957_347#_c_1051_n 0.00700601f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_449 N_A_1576_99#_c_504_n N_A_1957_347#_c_1053_n 0.00615404f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_450 N_A_1576_99#_M1022_g N_VPWR_c_1133_n 0.0198184f $X=8.005 $Y=2.235 $X2=0
+ $Y2=0
cc_451 N_A_1576_99#_c_508_n N_VPWR_c_1133_n 0.0108646f $X=9.27 $Y=2.59 $X2=0
+ $Y2=0
cc_452 N_A_1576_99#_c_508_n N_VPWR_c_1141_n 0.00755126f $X=9.27 $Y=2.59 $X2=0
+ $Y2=0
cc_453 N_A_1576_99#_M1022_g N_VPWR_c_1129_n 0.00141512f $X=8.005 $Y=2.235 $X2=0
+ $Y2=0
cc_454 N_A_1576_99#_c_508_n N_VPWR_c_1129_n 0.00910022f $X=9.27 $Y=2.59 $X2=0
+ $Y2=0
cc_455 N_A_1576_99#_c_501_n N_A_351_417#_c_1282_n 9.39913e-19 $X=8.045 $Y=0.98
+ $X2=0 $Y2=0
cc_456 N_A_1576_99#_c_497_n N_VGND_M1037_d 0.00222975f $X=8.945 $Y=0.98 $X2=0
+ $Y2=0
cc_457 N_A_1576_99#_c_501_n N_VGND_M1037_d 0.00182503f $X=8.045 $Y=0.98 $X2=0
+ $Y2=0
cc_458 N_A_1576_99#_c_497_n N_VGND_c_1416_n 0.0150101f $X=8.945 $Y=0.98 $X2=0
+ $Y2=0
cc_459 N_A_1576_99#_c_498_n N_VGND_c_1416_n 0.00786051f $X=9.11 $Y=0.835 $X2=0
+ $Y2=0
cc_460 N_A_1576_99#_c_499_n N_VGND_c_1416_n 0.00677668f $X=9.275 $Y=0.35 $X2=0
+ $Y2=0
cc_461 N_A_1576_99#_c_501_n N_VGND_c_1416_n 0.0105123f $X=8.045 $Y=0.98 $X2=0
+ $Y2=0
cc_462 N_A_1576_99#_c_502_n N_VGND_c_1416_n 5.63174e-19 $X=8.045 $Y=1.32 $X2=0
+ $Y2=0
cc_463 N_A_1576_99#_c_505_n N_VGND_c_1416_n 0.00195644f $X=8.045 $Y=1.155 $X2=0
+ $Y2=0
cc_464 N_A_1576_99#_c_500_n N_VGND_c_1417_n 0.00178819f $X=10.52 $Y=0.35 $X2=0
+ $Y2=0
cc_465 N_A_1576_99#_c_499_n N_VGND_c_1420_n 0.0222419f $X=9.275 $Y=0.35 $X2=0
+ $Y2=0
cc_466 N_A_1576_99#_c_500_n N_VGND_c_1420_n 0.0847403f $X=10.52 $Y=0.35 $X2=0
+ $Y2=0
cc_467 N_A_1576_99#_M1010_d N_VGND_c_1431_n 0.00272517f $X=10.375 $Y=0.205 $X2=0
+ $Y2=0
cc_468 N_A_1576_99#_c_499_n N_VGND_c_1431_n 0.0114525f $X=9.275 $Y=0.35 $X2=0
+ $Y2=0
cc_469 N_A_1576_99#_c_500_n N_VGND_c_1431_n 0.0517766f $X=10.52 $Y=0.35 $X2=0
+ $Y2=0
cc_470 N_A_1576_99#_c_505_n N_VGND_c_1431_n 9.49986e-19 $X=8.045 $Y=1.155 $X2=0
+ $Y2=0
cc_471 N_A_1576_99#_c_505_n N_A_1160_155#_c_1548_n 0.00124446f $X=8.045 $Y=1.155
+ $X2=0 $Y2=0
cc_472 N_A_1576_99#_c_497_n A_1722_125# 0.00166171f $X=8.945 $Y=0.98 $X2=-0.19
+ $Y2=-0.245
cc_473 N_A_1576_99#_c_498_n N_A_1910_155#_c_1581_n 0.00667074f $X=9.11 $Y=0.835
+ $X2=0 $Y2=0
cc_474 N_A_1576_99#_c_503_n N_A_1910_155#_c_1581_n 0.0110511f $X=9.11 $Y=0.98
+ $X2=0 $Y2=0
cc_475 N_A_1576_99#_c_504_n N_A_1910_155#_c_1581_n 0.00870173f $X=9.27 $Y=1.715
+ $X2=0 $Y2=0
cc_476 N_A_1576_99#_M1010_d N_A_1910_155#_c_1582_n 0.0109989f $X=10.375 $Y=0.205
+ $X2=0 $Y2=0
cc_477 N_A_1576_99#_c_500_n N_A_1910_155#_c_1582_n 0.0613851f $X=10.52 $Y=0.35
+ $X2=0 $Y2=0
cc_478 N_A_1576_99#_c_498_n N_A_1910_155#_c_1583_n 0.0113026f $X=9.11 $Y=0.835
+ $X2=0 $Y2=0
cc_479 N_A_1576_99#_c_500_n N_A_1910_155#_c_1583_n 0.0179592f $X=10.52 $Y=0.35
+ $X2=0 $Y2=0
cc_480 N_A_1576_99#_c_500_n N_A_1910_155#_c_1584_n 0.00776387f $X=10.52 $Y=0.35
+ $X2=0 $Y2=0
cc_481 N_A_1263_155#_c_594_n N_A_733_66#_M1009_g 0.00753045f $X=6.725 $Y=1.05
+ $X2=0 $Y2=0
cc_482 N_A_1263_155#_c_595_n N_A_733_66#_M1009_g 0.00178743f $X=7.085 $Y=1.45
+ $X2=0 $Y2=0
cc_483 N_A_1263_155#_c_594_n N_A_733_66#_M1007_g 0.00136496f $X=6.725 $Y=1.05
+ $X2=0 $Y2=0
cc_484 N_A_1263_155#_c_595_n N_A_733_66#_M1007_g 5.70967e-19 $X=7.085 $Y=1.45
+ $X2=0 $Y2=0
cc_485 N_A_1263_155#_c_601_n N_A_733_66#_M1007_g 0.0186025f $X=7.25 $Y=1.88
+ $X2=0 $Y2=0
cc_486 N_A_1263_155#_c_602_n N_A_733_66#_M1007_g 0.0254285f $X=8.46 $Y=1.75
+ $X2=0 $Y2=0
cc_487 N_A_1263_155#_c_598_n N_A_733_66#_M1007_g 0.0142842f $X=7.25 $Y=1.45
+ $X2=0 $Y2=0
cc_488 N_A_1263_155#_M1028_g N_A_733_66#_c_684_n 0.00868355f $X=8.535 $Y=0.835
+ $X2=0 $Y2=0
cc_489 N_A_1263_155#_M1016_g N_A_733_66#_c_684_n 0.00847339f $X=8.895 $Y=0.835
+ $X2=0 $Y2=0
cc_490 N_A_1263_155#_M1016_g N_A_733_66#_c_685_n 0.0144468f $X=8.895 $Y=0.835
+ $X2=0 $Y2=0
cc_491 N_A_1263_155#_c_599_n N_A_733_66#_c_685_n 0.00926782f $X=8.96 $Y=1.41
+ $X2=0 $Y2=0
cc_492 N_A_1263_155#_c_599_n N_A_733_66#_M1017_g 0.0198561f $X=8.96 $Y=1.41
+ $X2=0 $Y2=0
cc_493 N_A_1263_155#_c_594_n N_A_733_66#_c_693_n 4.83474e-19 $X=6.725 $Y=1.05
+ $X2=0 $Y2=0
cc_494 N_A_1263_155#_c_598_n N_A_733_66#_c_693_n 0.00104994f $X=7.25 $Y=1.45
+ $X2=0 $Y2=0
cc_495 N_A_1263_155#_c_596_n N_A_998_347#_c_842_n 5.76687e-19 $X=6.89 $Y=1.45
+ $X2=0 $Y2=0
cc_496 N_A_1263_155#_c_594_n N_A_998_347#_c_844_n 0.0015522f $X=6.725 $Y=1.05
+ $X2=0 $Y2=0
cc_497 N_A_1263_155#_c_595_n N_A_998_347#_M1021_g 0.00636688f $X=7.085 $Y=1.45
+ $X2=0 $Y2=0
cc_498 N_A_1263_155#_c_596_n N_A_998_347#_M1021_g 5.03796e-19 $X=6.89 $Y=1.45
+ $X2=0 $Y2=0
cc_499 N_A_1263_155#_c_601_n N_A_998_347#_M1021_g 0.0167798f $X=7.25 $Y=1.88
+ $X2=0 $Y2=0
cc_500 N_A_1263_155#_c_598_n N_A_998_347#_M1021_g 0.00901252f $X=7.25 $Y=1.45
+ $X2=0 $Y2=0
cc_501 N_A_1263_155#_M1036_g N_A_998_347#_c_853_n 0.0173606f $X=8.96 $Y=2.235
+ $X2=0 $Y2=0
cc_502 N_A_1263_155#_c_601_n N_A_998_347#_c_853_n 0.00392786f $X=7.25 $Y=1.88
+ $X2=0 $Y2=0
cc_503 N_A_1263_155#_c_602_n N_VPWR_M1022_d 0.0197619f $X=8.46 $Y=1.75 $X2=0
+ $Y2=0
cc_504 N_A_1263_155#_M1036_g N_VPWR_c_1133_n 0.010454f $X=8.96 $Y=2.235 $X2=0
+ $Y2=0
cc_505 N_A_1263_155#_c_602_n N_VPWR_c_1133_n 0.0209601f $X=8.46 $Y=1.75 $X2=0
+ $Y2=0
cc_506 N_A_1263_155#_c_601_n N_VPWR_c_1140_n 0.0074415f $X=7.25 $Y=1.88 $X2=0
+ $Y2=0
cc_507 N_A_1263_155#_M1036_g N_VPWR_c_1129_n 0.0015654f $X=8.96 $Y=2.235 $X2=0
+ $Y2=0
cc_508 N_A_1263_155#_c_601_n N_VPWR_c_1129_n 0.00902447f $X=7.25 $Y=1.88 $X2=0
+ $Y2=0
cc_509 N_A_1263_155#_M1023_d N_A_351_417#_c_1279_n 0.00493789f $X=6.315 $Y=0.775
+ $X2=0 $Y2=0
cc_510 N_A_1263_155#_c_594_n N_A_351_417#_c_1279_n 0.0297498f $X=6.725 $Y=1.05
+ $X2=0 $Y2=0
cc_511 N_A_1263_155#_c_596_n N_A_351_417#_c_1279_n 0.0134997f $X=6.89 $Y=1.45
+ $X2=0 $Y2=0
cc_512 N_A_1263_155#_M1023_d N_A_351_417#_c_1280_n 0.00965206f $X=6.315 $Y=0.775
+ $X2=0 $Y2=0
cc_513 N_A_1263_155#_c_594_n N_A_351_417#_c_1280_n 0.0206612f $X=6.725 $Y=1.05
+ $X2=0 $Y2=0
cc_514 N_A_1263_155#_c_595_n N_A_351_417#_c_1280_n 0.00437128f $X=7.085 $Y=1.45
+ $X2=0 $Y2=0
cc_515 N_A_1263_155#_c_601_n N_A_351_417#_c_1287_n 0.028333f $X=7.25 $Y=1.88
+ $X2=0 $Y2=0
cc_516 N_A_1263_155#_c_595_n N_A_351_417#_c_1282_n 0.00105288f $X=7.085 $Y=1.45
+ $X2=0 $Y2=0
cc_517 N_A_1263_155#_c_598_n N_A_351_417#_c_1282_n 0.0203227f $X=7.25 $Y=1.45
+ $X2=0 $Y2=0
cc_518 N_A_1263_155#_c_596_n N_A_351_417#_c_1289_n 0.0283831f $X=6.89 $Y=1.45
+ $X2=0 $Y2=0
cc_519 N_A_1263_155#_c_598_n N_A_351_417#_c_1289_n 0.0425307f $X=7.25 $Y=1.45
+ $X2=0 $Y2=0
cc_520 N_A_1263_155#_c_602_n A_1528_347# 0.0048076f $X=8.46 $Y=1.75 $X2=-0.19
+ $Y2=-0.245
cc_521 N_A_1263_155#_M1028_g N_VGND_c_1416_n 0.002478f $X=8.535 $Y=0.835 $X2=0
+ $Y2=0
cc_522 N_A_1263_155#_M1028_g N_VGND_c_1431_n 9.49986e-19 $X=8.535 $Y=0.835 $X2=0
+ $Y2=0
cc_523 N_A_1263_155#_M1016_g N_VGND_c_1431_n 7.94319e-19 $X=8.895 $Y=0.835 $X2=0
+ $Y2=0
cc_524 N_A_733_66#_M1012_g N_A_998_347#_c_849_n 0.0172245f $X=4.865 $Y=2.235
+ $X2=0 $Y2=0
cc_525 N_A_733_66#_c_699_n N_A_998_347#_c_843_n 0.00248017f $X=4.88 $Y=1.025
+ $X2=0 $Y2=0
cc_526 N_A_733_66#_c_679_n N_A_998_347#_c_844_n 0.00377117f $X=6.865 $Y=0.18
+ $X2=0 $Y2=0
cc_527 N_A_733_66#_M1009_g N_A_998_347#_c_844_n 0.00822585f $X=6.94 $Y=0.985
+ $X2=0 $Y2=0
cc_528 N_A_733_66#_M1009_g N_A_998_347#_M1021_g 0.00667669f $X=6.94 $Y=0.985
+ $X2=0 $Y2=0
cc_529 N_A_733_66#_M1007_g N_A_998_347#_M1021_g 0.0128253f $X=7.515 $Y=2.235
+ $X2=0 $Y2=0
cc_530 N_A_733_66#_M1007_g N_A_998_347#_c_853_n 0.0172445f $X=7.515 $Y=2.235
+ $X2=0 $Y2=0
cc_531 N_A_733_66#_M1017_g N_A_998_347#_c_853_n 0.0173606f $X=9.66 $Y=2.235
+ $X2=0 $Y2=0
cc_532 N_A_733_66#_M1017_g N_A_998_347#_c_855_n 0.0233693f $X=9.66 $Y=2.235
+ $X2=0 $Y2=0
cc_533 N_A_733_66#_M1017_g N_A_998_347#_M1010_g 0.00502515f $X=9.66 $Y=2.235
+ $X2=0 $Y2=0
cc_534 N_A_733_66#_c_687_n N_A_998_347#_M1010_g 0.0197043f $X=9.89 $Y=1.27 $X2=0
+ $Y2=0
cc_535 N_A_733_66#_c_676_n N_A_998_347#_c_846_n 0.00185108f $X=4.815 $Y=0.86
+ $X2=0 $Y2=0
cc_536 N_A_733_66#_M1027_g N_A_998_347#_c_846_n 0.0123097f $X=5.175 $Y=0.54
+ $X2=0 $Y2=0
cc_537 N_A_733_66#_c_679_n N_A_998_347#_c_846_n 0.00516985f $X=6.865 $Y=0.18
+ $X2=0 $Y2=0
cc_538 N_A_733_66#_c_688_n N_A_998_347#_c_846_n 0.00614714f $X=5.175 $Y=0.935
+ $X2=0 $Y2=0
cc_539 N_A_733_66#_c_696_n N_A_998_347#_c_846_n 0.0368438f $X=4.46 $Y=0.915
+ $X2=0 $Y2=0
cc_540 N_A_733_66#_c_699_n N_A_998_347#_c_846_n 0.00665921f $X=4.88 $Y=1.025
+ $X2=0 $Y2=0
cc_541 N_A_733_66#_M1012_g N_A_998_347#_c_847_n 0.00766477f $X=4.865 $Y=2.235
+ $X2=0 $Y2=0
cc_542 N_A_733_66#_c_689_n N_A_998_347#_c_847_n 3.82421e-19 $X=4.88 $Y=1.53
+ $X2=0 $Y2=0
cc_543 N_A_733_66#_c_703_n N_A_998_347#_c_847_n 0.0134797f $X=4.46 $Y=1.845
+ $X2=0 $Y2=0
cc_544 N_A_733_66#_c_696_n N_A_998_347#_c_847_n 0.0247267f $X=4.46 $Y=0.915
+ $X2=0 $Y2=0
cc_545 N_A_733_66#_c_698_n N_A_998_347#_c_847_n 0.00634447f $X=4.545 $Y=1.715
+ $X2=0 $Y2=0
cc_546 N_A_733_66#_c_699_n N_A_998_347#_c_847_n 0.00199386f $X=4.88 $Y=1.025
+ $X2=0 $Y2=0
cc_547 N_A_733_66#_M1012_g N_A_998_347#_c_848_n 0.00604777f $X=4.865 $Y=2.235
+ $X2=0 $Y2=0
cc_548 N_A_733_66#_c_689_n N_A_998_347#_c_848_n 0.00248017f $X=4.88 $Y=1.53
+ $X2=0 $Y2=0
cc_549 N_A_733_66#_M1017_g N_A_1957_347#_c_1057_n 0.0106972f $X=9.66 $Y=2.235
+ $X2=0 $Y2=0
cc_550 N_A_733_66#_c_685_n N_A_1957_347#_c_1051_n 2.29661e-19 $X=9.4 $Y=1.27
+ $X2=0 $Y2=0
cc_551 N_A_733_66#_M1017_g N_A_1957_347#_c_1051_n 7.77819e-19 $X=9.66 $Y=2.235
+ $X2=0 $Y2=0
cc_552 N_A_733_66#_c_687_n N_A_1957_347#_c_1051_n 0.00482451f $X=9.89 $Y=1.27
+ $X2=0 $Y2=0
cc_553 N_A_733_66#_c_694_n N_A_1957_347#_c_1051_n 0.00673731f $X=9.89 $Y=1.345
+ $X2=0 $Y2=0
cc_554 N_A_733_66#_M1017_g N_A_1957_347#_c_1053_n 0.00306756f $X=9.66 $Y=2.235
+ $X2=0 $Y2=0
cc_555 N_A_733_66#_c_694_n N_A_1957_347#_c_1053_n 0.00548523f $X=9.89 $Y=1.345
+ $X2=0 $Y2=0
cc_556 N_A_733_66#_c_703_n N_VPWR_M1029_d 0.00399987f $X=4.46 $Y=1.845 $X2=0
+ $Y2=0
cc_557 N_A_733_66#_M1012_g N_VPWR_c_1132_n 0.0184641f $X=4.865 $Y=2.235 $X2=0
+ $Y2=0
cc_558 N_A_733_66#_M1007_g N_VPWR_c_1133_n 0.0036745f $X=7.515 $Y=2.235 $X2=0
+ $Y2=0
cc_559 N_A_733_66#_M1012_g N_VPWR_c_1140_n 0.00646289f $X=4.865 $Y=2.235 $X2=0
+ $Y2=0
cc_560 N_A_733_66#_M1012_g N_VPWR_c_1129_n 0.00719887f $X=4.865 $Y=2.235 $X2=0
+ $Y2=0
cc_561 N_A_733_66#_M1007_g N_VPWR_c_1129_n 0.0015654f $X=7.515 $Y=2.235 $X2=0
+ $Y2=0
cc_562 N_A_733_66#_M1017_g N_VPWR_c_1129_n 0.0015654f $X=9.66 $Y=2.235 $X2=0
+ $Y2=0
cc_563 N_A_733_66#_M1009_g N_A_351_417#_c_1279_n 0.00302119f $X=6.94 $Y=0.985
+ $X2=0 $Y2=0
cc_564 N_A_733_66#_M1009_g N_A_351_417#_c_1280_n 0.0130136f $X=6.94 $Y=0.985
+ $X2=0 $Y2=0
cc_565 N_A_733_66#_c_692_n N_A_351_417#_c_1280_n 0.00184673f $X=7.505 $Y=1.12
+ $X2=0 $Y2=0
cc_566 N_A_733_66#_c_692_n N_A_351_417#_c_1282_n 0.00711127f $X=7.505 $Y=1.12
+ $X2=0 $Y2=0
cc_567 N_A_733_66#_M1029_s N_A_351_417#_c_1288_n 0.011995f $X=3.925 $Y=1.735
+ $X2=0 $Y2=0
cc_568 N_A_733_66#_M1012_g N_A_351_417#_c_1288_n 0.0258518f $X=4.865 $Y=2.235
+ $X2=0 $Y2=0
cc_569 N_A_733_66#_c_703_n N_A_351_417#_c_1288_n 0.043359f $X=4.46 $Y=1.845
+ $X2=0 $Y2=0
cc_570 N_A_733_66#_c_696_n N_A_351_417#_c_1288_n 0.00849888f $X=4.46 $Y=0.915
+ $X2=0 $Y2=0
cc_571 N_A_733_66#_c_695_n N_VGND_c_1414_n 0.0355608f $X=3.81 $Y=0.54 $X2=0
+ $Y2=0
cc_572 N_A_733_66#_c_697_n N_VGND_c_1414_n 0.0123489f $X=3.975 $Y=0.915 $X2=0
+ $Y2=0
cc_573 N_A_733_66#_c_676_n N_VGND_c_1415_n 0.00983875f $X=4.815 $Y=0.86 $X2=0
+ $Y2=0
cc_574 N_A_733_66#_c_680_n N_VGND_c_1415_n 0.0038616f $X=5.25 $Y=0.18 $X2=0
+ $Y2=0
cc_575 N_A_733_66#_c_695_n N_VGND_c_1415_n 0.0113755f $X=3.81 $Y=0.54 $X2=0
+ $Y2=0
cc_576 N_A_733_66#_c_696_n N_VGND_c_1415_n 0.0224996f $X=4.46 $Y=0.915 $X2=0
+ $Y2=0
cc_577 N_A_733_66#_c_684_n N_VGND_c_1416_n 0.0255216f $X=9.325 $Y=0.18 $X2=0
+ $Y2=0
cc_578 N_A_733_66#_c_692_n N_VGND_c_1416_n 0.001031f $X=7.505 $Y=1.12 $X2=0
+ $Y2=0
cc_579 N_A_733_66#_c_684_n N_VGND_c_1420_n 0.0304792f $X=9.325 $Y=0.18 $X2=0
+ $Y2=0
cc_580 N_A_733_66#_c_695_n N_VGND_c_1424_n 0.0173629f $X=3.81 $Y=0.54 $X2=0
+ $Y2=0
cc_581 N_A_733_66#_c_676_n N_VGND_c_1425_n 0.00411131f $X=4.815 $Y=0.86 $X2=0
+ $Y2=0
cc_582 N_A_733_66#_c_680_n N_VGND_c_1425_n 0.0729479f $X=5.25 $Y=0.18 $X2=0
+ $Y2=0
cc_583 N_A_733_66#_c_676_n N_VGND_c_1431_n 0.00401612f $X=4.815 $Y=0.86 $X2=0
+ $Y2=0
cc_584 N_A_733_66#_c_679_n N_VGND_c_1431_n 0.0449542f $X=6.865 $Y=0.18 $X2=0
+ $Y2=0
cc_585 N_A_733_66#_c_680_n N_VGND_c_1431_n 0.0101746f $X=5.25 $Y=0.18 $X2=0
+ $Y2=0
cc_586 N_A_733_66#_c_682_n N_VGND_c_1431_n 0.00848224f $X=7.37 $Y=0.18 $X2=0
+ $Y2=0
cc_587 N_A_733_66#_c_684_n N_VGND_c_1431_n 0.055636f $X=9.325 $Y=0.18 $X2=0
+ $Y2=0
cc_588 N_A_733_66#_c_690_n N_VGND_c_1431_n 0.00371014f $X=6.94 $Y=0.18 $X2=0
+ $Y2=0
cc_589 N_A_733_66#_c_691_n N_VGND_c_1431_n 0.00371014f $X=7.445 $Y=0.18 $X2=0
+ $Y2=0
cc_590 N_A_733_66#_c_695_n N_VGND_c_1431_n 0.0122896f $X=3.81 $Y=0.54 $X2=0
+ $Y2=0
cc_591 N_A_733_66#_c_696_n N_VGND_c_1431_n 0.0256668f $X=4.46 $Y=0.915 $X2=0
+ $Y2=0
cc_592 N_A_733_66#_M1027_g N_A_1160_155#_c_1545_n 0.00151807f $X=5.175 $Y=0.54
+ $X2=0 $Y2=0
cc_593 N_A_733_66#_c_679_n N_A_1160_155#_c_1546_n 0.0152969f $X=6.865 $Y=0.18
+ $X2=0 $Y2=0
cc_594 N_A_733_66#_M1009_g N_A_1160_155#_c_1546_n 0.0123198f $X=6.94 $Y=0.985
+ $X2=0 $Y2=0
cc_595 N_A_733_66#_c_682_n N_A_1160_155#_c_1546_n 0.00408708f $X=7.37 $Y=0.18
+ $X2=0 $Y2=0
cc_596 N_A_733_66#_c_684_n N_A_1160_155#_c_1546_n 0.00529313f $X=9.325 $Y=0.18
+ $X2=0 $Y2=0
cc_597 N_A_733_66#_c_692_n N_A_1160_155#_c_1546_n 0.0161867f $X=7.505 $Y=1.12
+ $X2=0 $Y2=0
cc_598 N_A_733_66#_c_693_n N_A_1160_155#_c_1546_n 0.00133371f $X=7.505 $Y=1.27
+ $X2=0 $Y2=0
cc_599 N_A_733_66#_M1027_g N_A_1160_155#_c_1547_n 0.00160285f $X=5.175 $Y=0.54
+ $X2=0 $Y2=0
cc_600 N_A_733_66#_c_679_n N_A_1160_155#_c_1547_n 0.00615835f $X=6.865 $Y=0.18
+ $X2=0 $Y2=0
cc_601 N_A_733_66#_c_692_n N_A_1160_155#_c_1548_n 0.00907827f $X=7.505 $Y=1.12
+ $X2=0 $Y2=0
cc_602 N_A_733_66#_c_693_n N_A_1160_155#_c_1548_n 0.00317658f $X=7.505 $Y=1.27
+ $X2=0 $Y2=0
cc_603 N_A_733_66#_c_685_n N_A_1910_155#_c_1581_n 0.00399925f $X=9.4 $Y=1.27
+ $X2=0 $Y2=0
cc_604 N_A_733_66#_c_687_n N_A_1910_155#_c_1581_n 2.61813e-19 $X=9.89 $Y=1.27
+ $X2=0 $Y2=0
cc_605 N_A_733_66#_c_694_n N_A_1910_155#_c_1581_n 0.00859761f $X=9.89 $Y=1.345
+ $X2=0 $Y2=0
cc_606 N_A_733_66#_c_687_n N_A_1910_155#_c_1582_n 0.0130709f $X=9.89 $Y=1.27
+ $X2=0 $Y2=0
cc_607 N_A_733_66#_c_685_n N_A_1910_155#_c_1583_n 0.0022214f $X=9.4 $Y=1.27
+ $X2=0 $Y2=0
cc_608 N_A_998_347#_c_855_n N_A_2148_185#_M1026_g 0.0646095f $X=10.32 $Y=1.65
+ $X2=0 $Y2=0
cc_609 N_A_998_347#_M1010_g N_A_2148_185#_c_955_n 0.00116492f $X=10.32 $Y=0.985
+ $X2=0 $Y2=0
cc_610 N_A_998_347#_M1010_g N_A_2148_185#_c_956_n 0.0258395f $X=10.32 $Y=0.985
+ $X2=0 $Y2=0
cc_611 N_A_998_347#_c_853_n N_A_1957_347#_c_1057_n 0.00629123f $X=10.225 $Y=3.15
+ $X2=0 $Y2=0
cc_612 N_A_998_347#_c_855_n N_A_1957_347#_c_1057_n 0.0113727f $X=10.32 $Y=1.65
+ $X2=0 $Y2=0
cc_613 N_A_998_347#_M1010_g N_A_1957_347#_c_1057_n 8.44101e-19 $X=10.32 $Y=0.985
+ $X2=0 $Y2=0
cc_614 N_A_998_347#_M1010_g N_A_1957_347#_c_1051_n 0.0128976f $X=10.32 $Y=0.985
+ $X2=0 $Y2=0
cc_615 N_A_998_347#_c_855_n N_A_1957_347#_c_1052_n 0.00397798f $X=10.32 $Y=1.65
+ $X2=0 $Y2=0
cc_616 N_A_998_347#_M1010_g N_A_1957_347#_c_1052_n 0.0152449f $X=10.32 $Y=0.985
+ $X2=0 $Y2=0
cc_617 N_A_998_347#_c_855_n N_A_1957_347#_c_1053_n 0.00112041f $X=10.32 $Y=1.65
+ $X2=0 $Y2=0
cc_618 N_A_998_347#_M1010_g N_A_1957_347#_c_1053_n 0.00426042f $X=10.32 $Y=0.985
+ $X2=0 $Y2=0
cc_619 N_A_998_347#_c_853_n N_VPWR_c_1133_n 0.025796f $X=10.225 $Y=3.15 $X2=0
+ $Y2=0
cc_620 N_A_998_347#_M1033_g N_VPWR_c_1134_n 0.0114903f $X=10.35 $Y=2.305 $X2=0
+ $Y2=0
cc_621 N_A_998_347#_c_851_n N_VPWR_c_1140_n 0.0809525f $X=5.82 $Y=3.15 $X2=0
+ $Y2=0
cc_622 N_A_998_347#_c_853_n N_VPWR_c_1141_n 0.0655751f $X=10.225 $Y=3.15 $X2=0
+ $Y2=0
cc_623 N_A_998_347#_c_850_n N_VPWR_c_1129_n 0.0487619f $X=6.86 $Y=3.15 $X2=0
+ $Y2=0
cc_624 N_A_998_347#_c_851_n N_VPWR_c_1129_n 0.0116041f $X=5.82 $Y=3.15 $X2=0
+ $Y2=0
cc_625 N_A_998_347#_c_853_n N_VPWR_c_1129_n 0.121235f $X=10.225 $Y=3.15 $X2=0
+ $Y2=0
cc_626 N_A_998_347#_c_858_n N_VPWR_c_1129_n 0.0138136f $X=6.985 $Y=3.15 $X2=0
+ $Y2=0
cc_627 N_A_998_347#_c_842_n N_A_351_417#_c_1279_n 0.00892391f $X=6.165 $Y=1.38
+ $X2=0 $Y2=0
cc_628 N_A_998_347#_c_844_n N_A_351_417#_c_1279_n 0.0155972f $X=6.24 $Y=1.305
+ $X2=0 $Y2=0
cc_629 N_A_998_347#_M1021_g N_A_351_417#_c_1279_n 0.00288505f $X=6.985 $Y=2.235
+ $X2=0 $Y2=0
cc_630 N_A_998_347#_c_846_n N_A_351_417#_c_1279_n 0.00487387f $X=5.39 $Y=0.54
+ $X2=0 $Y2=0
cc_631 N_A_998_347#_c_847_n N_A_351_417#_c_1279_n 0.016764f $X=5.39 $Y=1.64
+ $X2=0 $Y2=0
cc_632 N_A_998_347#_c_848_n N_A_351_417#_c_1279_n 9.97538e-19 $X=5.655 $Y=1.47
+ $X2=0 $Y2=0
cc_633 N_A_998_347#_c_844_n N_A_351_417#_c_1281_n 0.00552634f $X=6.24 $Y=1.305
+ $X2=0 $Y2=0
cc_634 N_A_998_347#_c_850_n N_A_351_417#_c_1287_n 0.00420701f $X=6.86 $Y=3.15
+ $X2=0 $Y2=0
cc_635 N_A_998_347#_M1021_g N_A_351_417#_c_1287_n 0.00816224f $X=6.985 $Y=2.235
+ $X2=0 $Y2=0
cc_636 N_A_998_347#_M1012_d N_A_351_417#_c_1288_n 0.0121584f $X=4.99 $Y=1.735
+ $X2=0 $Y2=0
cc_637 N_A_998_347#_c_849_n N_A_351_417#_c_1288_n 0.0185931f $X=5.745 $Y=3.075
+ $X2=0 $Y2=0
cc_638 N_A_998_347#_c_857_n N_A_351_417#_c_1288_n 0.00123832f $X=5.655 $Y=1.975
+ $X2=0 $Y2=0
cc_639 N_A_998_347#_c_847_n N_A_351_417#_c_1288_n 0.0605008f $X=5.39 $Y=1.64
+ $X2=0 $Y2=0
cc_640 N_A_998_347#_c_849_n N_A_351_417#_c_1289_n 0.0057967f $X=5.745 $Y=3.075
+ $X2=0 $Y2=0
cc_641 N_A_998_347#_c_842_n N_A_351_417#_c_1289_n 3.83008e-19 $X=6.165 $Y=1.38
+ $X2=0 $Y2=0
cc_642 N_A_998_347#_M1021_g N_A_351_417#_c_1289_n 0.0111913f $X=6.985 $Y=2.235
+ $X2=0 $Y2=0
cc_643 N_A_998_347#_c_847_n N_A_351_417#_c_1289_n 0.0123583f $X=5.39 $Y=1.64
+ $X2=0 $Y2=0
cc_644 N_A_998_347#_c_848_n N_A_351_417#_c_1289_n 0.00181484f $X=5.655 $Y=1.47
+ $X2=0 $Y2=0
cc_645 N_A_998_347#_c_846_n N_VGND_c_1415_n 0.0113755f $X=5.39 $Y=0.54 $X2=0
+ $Y2=0
cc_646 N_A_998_347#_c_846_n N_VGND_c_1425_n 0.0173367f $X=5.39 $Y=0.54 $X2=0
+ $Y2=0
cc_647 N_A_998_347#_c_846_n N_VGND_c_1431_n 0.0110393f $X=5.39 $Y=0.54 $X2=0
+ $Y2=0
cc_648 N_A_998_347#_c_842_n N_A_1160_155#_c_1545_n 0.00848258f $X=6.165 $Y=1.38
+ $X2=0 $Y2=0
cc_649 N_A_998_347#_c_843_n N_A_1160_155#_c_1545_n 3.02817e-19 $X=5.82 $Y=1.38
+ $X2=0 $Y2=0
cc_650 N_A_998_347#_c_844_n N_A_1160_155#_c_1545_n 0.00972362f $X=6.24 $Y=1.305
+ $X2=0 $Y2=0
cc_651 N_A_998_347#_c_846_n N_A_1160_155#_c_1545_n 0.0462272f $X=5.39 $Y=0.54
+ $X2=0 $Y2=0
cc_652 N_A_998_347#_c_847_n N_A_1160_155#_c_1545_n 0.0032901f $X=5.39 $Y=1.64
+ $X2=0 $Y2=0
cc_653 N_A_998_347#_c_844_n N_A_1160_155#_c_1546_n 0.00134976f $X=6.24 $Y=1.305
+ $X2=0 $Y2=0
cc_654 N_A_998_347#_c_846_n N_A_1160_155#_c_1547_n 0.00908019f $X=5.39 $Y=0.54
+ $X2=0 $Y2=0
cc_655 N_A_998_347#_M1010_g N_A_1910_155#_c_1582_n 0.0150172f $X=10.32 $Y=0.985
+ $X2=0 $Y2=0
cc_656 N_A_2148_185#_M1026_g N_A_1957_347#_c_1047_n 0.0415414f $X=10.865
+ $Y=2.305 $X2=0 $Y2=0
cc_657 N_A_2148_185#_c_953_n N_A_1957_347#_c_1047_n 0.0019863f $X=11.855 $Y=1.05
+ $X2=0 $Y2=0
cc_658 N_A_2148_185#_c_956_n N_A_1957_347#_c_1047_n 0.00111824f $X=10.94 $Y=1.13
+ $X2=0 $Y2=0
cc_659 N_A_2148_185#_c_963_n N_A_1957_347#_c_1047_n 0.00623112f $X=11.735
+ $Y=1.99 $X2=0 $Y2=0
cc_660 N_A_2148_185#_c_957_n N_A_1957_347#_c_1047_n 0.00441692f $X=11.797
+ $Y=1.825 $X2=0 $Y2=0
cc_661 N_A_2148_185#_c_959_n N_A_1957_347#_c_1047_n 0.00431422f $X=12.56 $Y=1.13
+ $X2=0 $Y2=0
cc_662 N_A_2148_185#_c_963_n N_A_1957_347#_M1031_g 0.0222436f $X=11.735 $Y=1.99
+ $X2=0 $Y2=0
cc_663 N_A_2148_185#_c_957_n N_A_1957_347#_M1031_g 0.00555926f $X=11.797
+ $Y=1.825 $X2=0 $Y2=0
cc_664 N_A_2148_185#_M1001_g N_A_1957_347#_M1024_g 0.0224671f $X=11.29 $Y=0.555
+ $X2=0 $Y2=0
cc_665 N_A_2148_185#_c_953_n N_A_1957_347#_M1024_g 0.017639f $X=11.855 $Y=1.05
+ $X2=0 $Y2=0
cc_666 N_A_2148_185#_c_955_n N_A_1957_347#_M1024_g 0.00103348f $X=10.94 $Y=1.05
+ $X2=0 $Y2=0
cc_667 N_A_2148_185#_c_956_n N_A_1957_347#_M1024_g 0.00516117f $X=10.94 $Y=1.13
+ $X2=0 $Y2=0
cc_668 N_A_2148_185#_c_957_n N_A_1957_347#_M1024_g 6.79797e-19 $X=11.797
+ $Y=1.825 $X2=0 $Y2=0
cc_669 N_A_2148_185#_c_960_n N_A_1957_347#_M1024_g 0.0021612f $X=12.295 $Y=0.555
+ $X2=0 $Y2=0
cc_670 N_A_2148_185#_c_963_n N_A_1957_347#_c_1049_n 0.00201617f $X=11.735
+ $Y=1.99 $X2=0 $Y2=0
cc_671 N_A_2148_185#_c_957_n N_A_1957_347#_c_1049_n 0.014676f $X=11.797 $Y=1.825
+ $X2=0 $Y2=0
cc_672 N_A_2148_185#_c_958_n N_A_1957_347#_c_1049_n 3.55305e-19 $X=12.56 $Y=1.13
+ $X2=0 $Y2=0
cc_673 N_A_2148_185#_c_959_n N_A_1957_347#_c_1049_n 0.00953691f $X=12.56 $Y=1.13
+ $X2=0 $Y2=0
cc_674 N_A_2148_185#_c_948_n N_A_1957_347#_M1013_g 0.00953691f $X=12.725 $Y=1.04
+ $X2=0 $Y2=0
cc_675 N_A_2148_185#_c_954_n N_A_1957_347#_M1013_g 0.00614242f $X=12.215
+ $Y=0.965 $X2=0 $Y2=0
cc_676 N_A_2148_185#_c_957_n N_A_1957_347#_M1013_g 6.32775e-19 $X=11.797
+ $Y=1.825 $X2=0 $Y2=0
cc_677 N_A_2148_185#_c_958_n N_A_1957_347#_M1013_g 0.0171482f $X=12.56 $Y=1.13
+ $X2=0 $Y2=0
cc_678 N_A_2148_185#_c_960_n N_A_1957_347#_M1013_g 0.00896472f $X=12.295
+ $Y=0.555 $X2=0 $Y2=0
cc_679 N_A_2148_185#_c_955_n N_A_1957_347#_c_1051_n 0.010184f $X=10.94 $Y=1.05
+ $X2=0 $Y2=0
cc_680 N_A_2148_185#_c_956_n N_A_1957_347#_c_1051_n 0.002094f $X=10.94 $Y=1.13
+ $X2=0 $Y2=0
cc_681 N_A_2148_185#_M1026_g N_A_1957_347#_c_1052_n 0.0235291f $X=10.865
+ $Y=2.305 $X2=0 $Y2=0
cc_682 N_A_2148_185#_c_953_n N_A_1957_347#_c_1052_n 0.0111857f $X=11.855 $Y=1.05
+ $X2=0 $Y2=0
cc_683 N_A_2148_185#_c_955_n N_A_1957_347#_c_1052_n 0.022915f $X=10.94 $Y=1.05
+ $X2=0 $Y2=0
cc_684 N_A_2148_185#_c_956_n N_A_1957_347#_c_1052_n 0.00209257f $X=10.94 $Y=1.13
+ $X2=0 $Y2=0
cc_685 N_A_2148_185#_M1026_g N_A_1957_347#_c_1054_n 0.00111993f $X=10.865
+ $Y=2.305 $X2=0 $Y2=0
cc_686 N_A_2148_185#_c_953_n N_A_1957_347#_c_1054_n 0.0236129f $X=11.855 $Y=1.05
+ $X2=0 $Y2=0
cc_687 N_A_2148_185#_c_963_n N_A_1957_347#_c_1054_n 0.00560763f $X=11.735
+ $Y=1.99 $X2=0 $Y2=0
cc_688 N_A_2148_185#_c_957_n N_A_1957_347#_c_1054_n 0.0237523f $X=11.797
+ $Y=1.825 $X2=0 $Y2=0
cc_689 N_A_2148_185#_M1026_g N_VPWR_c_1134_n 0.0281129f $X=10.865 $Y=2.305 $X2=0
+ $Y2=0
cc_690 N_A_2148_185#_c_963_n N_VPWR_c_1134_n 0.0273743f $X=11.735 $Y=1.99 $X2=0
+ $Y2=0
cc_691 N_A_2148_185#_M1006_g N_VPWR_c_1136_n 0.0278522f $X=13.375 $Y=2.44 $X2=0
+ $Y2=0
cc_692 N_A_2148_185#_M1026_g N_VPWR_c_1141_n 0.00707094f $X=10.865 $Y=2.305
+ $X2=0 $Y2=0
cc_693 N_A_2148_185#_M1006_g N_VPWR_c_1142_n 0.00817829f $X=13.375 $Y=2.44 $X2=0
+ $Y2=0
cc_694 N_A_2148_185#_c_963_n N_VPWR_c_1142_n 0.0123069f $X=11.735 $Y=1.99 $X2=0
+ $Y2=0
cc_695 N_A_2148_185#_M1026_g N_VPWR_c_1129_n 0.0075026f $X=10.865 $Y=2.305 $X2=0
+ $Y2=0
cc_696 N_A_2148_185#_M1006_g N_VPWR_c_1129_n 0.00812777f $X=13.375 $Y=2.44 $X2=0
+ $Y2=0
cc_697 N_A_2148_185#_c_963_n N_VPWR_c_1129_n 0.0150765f $X=11.735 $Y=1.99 $X2=0
+ $Y2=0
cc_698 N_A_2148_185#_c_948_n N_Q_c_1383_n 0.00855454f $X=12.725 $Y=1.04 $X2=0
+ $Y2=0
cc_699 N_A_2148_185#_M1002_g N_Q_c_1383_n 0.0108661f $X=13.065 $Y=0.555 $X2=0
+ $Y2=0
cc_700 N_A_2148_185#_M1035_g N_Q_c_1383_n 0.00239934f $X=13.425 $Y=0.555 $X2=0
+ $Y2=0
cc_701 N_A_2148_185#_c_958_n N_Q_c_1383_n 0.00291485f $X=12.56 $Y=1.13 $X2=0
+ $Y2=0
cc_702 N_A_2148_185#_c_960_n N_Q_c_1383_n 0.0318905f $X=12.295 $Y=0.555 $X2=0
+ $Y2=0
cc_703 N_A_2148_185#_M1006_g Q 0.0077196f $X=13.375 $Y=2.44 $X2=0 $Y2=0
cc_704 N_A_2148_185#_c_963_n Q 0.0173569f $X=11.735 $Y=1.99 $X2=0 $Y2=0
cc_705 N_A_2148_185#_c_958_n Q 0.00698704f $X=12.56 $Y=1.13 $X2=0 $Y2=0
cc_706 N_A_2148_185#_c_959_n Q 8.69545e-19 $X=12.56 $Y=1.13 $X2=0 $Y2=0
cc_707 N_A_2148_185#_M1006_g Q 0.0133579f $X=13.375 $Y=2.44 $X2=0 $Y2=0
cc_708 N_A_2148_185#_c_963_n Q 0.0173569f $X=11.735 $Y=1.99 $X2=0 $Y2=0
cc_709 N_A_2148_185#_c_947_n N_Q_c_1384_n 0.00721701f $X=12.99 $Y=1.04 $X2=0
+ $Y2=0
cc_710 N_A_2148_185#_M1002_g N_Q_c_1384_n 0.00706462f $X=13.065 $Y=0.555 $X2=0
+ $Y2=0
cc_711 N_A_2148_185#_M1006_g N_Q_c_1384_n 0.0228825f $X=13.375 $Y=2.44 $X2=0
+ $Y2=0
cc_712 N_A_2148_185#_c_952_n N_Q_c_1384_n 0.00947522f $X=13.425 $Y=1.04 $X2=0
+ $Y2=0
cc_713 N_A_2148_185#_c_954_n N_Q_c_1384_n 0.00404804f $X=12.215 $Y=0.965 $X2=0
+ $Y2=0
cc_714 N_A_2148_185#_c_958_n N_Q_c_1384_n 0.0482464f $X=12.56 $Y=1.13 $X2=0
+ $Y2=0
cc_715 N_A_2148_185#_c_959_n N_Q_c_1384_n 0.00458652f $X=12.56 $Y=1.13 $X2=0
+ $Y2=0
cc_716 N_A_2148_185#_M1001_g N_VGND_c_1417_n 0.0108146f $X=11.29 $Y=0.555 $X2=0
+ $Y2=0
cc_717 N_A_2148_185#_c_953_n N_VGND_c_1417_n 0.0262009f $X=11.855 $Y=1.05 $X2=0
+ $Y2=0
cc_718 N_A_2148_185#_c_960_n N_VGND_c_1417_n 0.0153904f $X=12.295 $Y=0.555 $X2=0
+ $Y2=0
cc_719 N_A_2148_185#_M1002_g N_VGND_c_1419_n 0.00186275f $X=13.065 $Y=0.555
+ $X2=0 $Y2=0
cc_720 N_A_2148_185#_M1035_g N_VGND_c_1419_n 0.0142291f $X=13.425 $Y=0.555 $X2=0
+ $Y2=0
cc_721 N_A_2148_185#_M1001_g N_VGND_c_1420_n 0.00400407f $X=11.29 $Y=0.555 $X2=0
+ $Y2=0
cc_722 N_A_2148_185#_M1002_g N_VGND_c_1426_n 0.00381277f $X=13.065 $Y=0.555
+ $X2=0 $Y2=0
cc_723 N_A_2148_185#_M1035_g N_VGND_c_1426_n 0.00400407f $X=13.425 $Y=0.555
+ $X2=0 $Y2=0
cc_724 N_A_2148_185#_c_960_n N_VGND_c_1426_n 0.015931f $X=12.295 $Y=0.555 $X2=0
+ $Y2=0
cc_725 N_A_2148_185#_M1001_g N_VGND_c_1431_n 0.00804497f $X=11.29 $Y=0.555 $X2=0
+ $Y2=0
cc_726 N_A_2148_185#_M1002_g N_VGND_c_1431_n 0.00670522f $X=13.065 $Y=0.555
+ $X2=0 $Y2=0
cc_727 N_A_2148_185#_M1035_g N_VGND_c_1431_n 0.00769986f $X=13.425 $Y=0.555
+ $X2=0 $Y2=0
cc_728 N_A_2148_185#_c_960_n N_VGND_c_1431_n 0.0120937f $X=12.295 $Y=0.555 $X2=0
+ $Y2=0
cc_729 N_A_2148_185#_M1001_g N_A_1910_155#_c_1582_n 7.48457e-19 $X=11.29
+ $Y=0.555 $X2=0 $Y2=0
cc_730 N_A_2148_185#_c_953_n N_A_1910_155#_c_1582_n 0.00411296f $X=11.855
+ $Y=1.05 $X2=0 $Y2=0
cc_731 N_A_2148_185#_c_955_n N_A_1910_155#_c_1582_n 0.0249021f $X=10.94 $Y=1.05
+ $X2=0 $Y2=0
cc_732 N_A_2148_185#_c_956_n N_A_1910_155#_c_1582_n 0.0114306f $X=10.94 $Y=1.13
+ $X2=0 $Y2=0
cc_733 N_A_2148_185#_M1001_g N_A_1910_155#_c_1584_n 7.31217e-19 $X=11.29
+ $Y=0.555 $X2=0 $Y2=0
cc_734 N_A_1957_347#_M1031_g N_VPWR_c_1134_n 0.00914188f $X=11.47 $Y=2.305 $X2=0
+ $Y2=0
cc_735 N_A_1957_347#_c_1052_n N_VPWR_c_1134_n 0.0231064f $X=11.345 $Y=1.56 $X2=0
+ $Y2=0
cc_736 N_A_1957_347#_c_1057_n N_VPWR_c_1141_n 0.00894219f $X=10.005 $Y=1.88
+ $X2=0 $Y2=0
cc_737 N_A_1957_347#_M1031_g N_VPWR_c_1142_n 0.00767722f $X=11.47 $Y=2.305 $X2=0
+ $Y2=0
cc_738 N_A_1957_347#_M1031_g N_VPWR_c_1129_n 0.00829933f $X=11.47 $Y=2.305 $X2=0
+ $Y2=0
cc_739 N_A_1957_347#_c_1057_n N_VPWR_c_1129_n 0.00962586f $X=10.005 $Y=1.88
+ $X2=0 $Y2=0
cc_740 N_A_1957_347#_M1013_g N_Q_c_1383_n 9.74305e-19 $X=12.08 $Y=0.555 $X2=0
+ $Y2=0
cc_741 N_A_1957_347#_M1024_g N_VGND_c_1417_n 0.0123079f $X=11.72 $Y=0.555 $X2=0
+ $Y2=0
cc_742 N_A_1957_347#_M1013_g N_VGND_c_1417_n 0.00190651f $X=12.08 $Y=0.555 $X2=0
+ $Y2=0
cc_743 N_A_1957_347#_M1024_g N_VGND_c_1426_n 0.00400407f $X=11.72 $Y=0.555 $X2=0
+ $Y2=0
cc_744 N_A_1957_347#_M1013_g N_VGND_c_1426_n 0.00453398f $X=12.08 $Y=0.555 $X2=0
+ $Y2=0
cc_745 N_A_1957_347#_M1024_g N_VGND_c_1431_n 0.00769986f $X=11.72 $Y=0.555 $X2=0
+ $Y2=0
cc_746 N_A_1957_347#_M1013_g N_VGND_c_1431_n 0.00891576f $X=12.08 $Y=0.555 $X2=0
+ $Y2=0
cc_747 N_A_1957_347#_c_1051_n N_A_1910_155#_c_1581_n 0.0101339f $X=10.105
+ $Y=1.05 $X2=0 $Y2=0
cc_748 N_A_1957_347#_M1008_d N_A_1910_155#_c_1582_n 0.00180746f $X=9.965
+ $Y=0.775 $X2=0 $Y2=0
cc_749 N_A_1957_347#_c_1051_n N_A_1910_155#_c_1582_n 0.0163515f $X=10.105
+ $Y=1.05 $X2=0 $Y2=0
cc_750 N_VPWR_c_1129_n N_A_244_417#_M1011_s 0.0022865f $X=13.68 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_751 N_VPWR_c_1129_n N_A_244_417#_M1014_d 0.00229455f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_752 N_VPWR_c_1130_n N_A_244_417#_c_1237_n 0.0300845f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_753 N_VPWR_M1030_d N_A_244_417#_c_1238_n 0.00354096f $X=2.755 $Y=2.085 $X2=0
+ $Y2=0
cc_754 N_VPWR_c_1131_n N_A_244_417#_c_1238_n 0.0152929f $X=2.895 $Y=2.94 $X2=0
+ $Y2=0
cc_755 N_VPWR_c_1137_n N_A_244_417#_c_1238_n 0.0175598f $X=2.73 $Y=3.33 $X2=0
+ $Y2=0
cc_756 N_VPWR_c_1139_n N_A_244_417#_c_1238_n 0.00310358f $X=4.435 $Y=3.33 $X2=0
+ $Y2=0
cc_757 N_VPWR_c_1129_n N_A_244_417#_c_1238_n 0.0363669f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_758 N_VPWR_c_1131_n N_A_244_417#_c_1239_n 0.013837f $X=2.895 $Y=2.94 $X2=0
+ $Y2=0
cc_759 N_VPWR_c_1139_n N_A_244_417#_c_1239_n 0.0195379f $X=4.435 $Y=3.33 $X2=0
+ $Y2=0
cc_760 N_VPWR_c_1129_n N_A_244_417#_c_1239_n 0.0125146f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_761 N_VPWR_c_1130_n N_A_244_417#_c_1240_n 0.0390108f $X=0.81 $Y=2.19 $X2=0
+ $Y2=0
cc_762 N_VPWR_c_1137_n N_A_244_417#_c_1240_n 0.019758f $X=2.73 $Y=3.33 $X2=0
+ $Y2=0
cc_763 N_VPWR_c_1129_n N_A_244_417#_c_1240_n 0.012508f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_764 N_VPWR_c_1129_n N_A_351_417#_M1011_d 0.00333718f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_765 N_VPWR_c_1140_n N_A_351_417#_c_1287_n 0.00725013f $X=8.105 $Y=3.33 $X2=0
+ $Y2=0
cc_766 N_VPWR_c_1129_n N_A_351_417#_c_1287_n 0.00884694f $X=13.68 $Y=3.33 $X2=0
+ $Y2=0
cc_767 N_VPWR_M1030_d N_A_351_417#_c_1288_n 0.00780837f $X=2.755 $Y=2.085 $X2=0
+ $Y2=0
cc_768 N_VPWR_M1029_d N_A_351_417#_c_1288_n 0.00411515f $X=4.46 $Y=1.735 $X2=0
+ $Y2=0
cc_769 N_VPWR_c_1132_n N_A_351_417#_c_1288_n 0.0163515f $X=4.6 $Y=2.59 $X2=0
+ $Y2=0
cc_770 N_VPWR_c_1129_n A_457_417# 0.00262207f $X=13.68 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_771 N_VPWR_c_1136_n Q 0.0724063f $X=13.64 $Y=2.085 $X2=0 $Y2=0
cc_772 N_VPWR_c_1142_n Q 0.0275196f $X=13.475 $Y=3.33 $X2=0 $Y2=0
cc_773 N_VPWR_c_1129_n Q 0.0243516f $X=13.68 $Y=3.33 $X2=0 $Y2=0
cc_774 N_A_244_417#_c_1238_n N_A_351_417#_M1011_d 0.00475803f $X=3.26 $Y=2.59
+ $X2=0 $Y2=0
cc_775 N_A_244_417#_c_1237_n N_A_351_417#_c_1284_n 0.0180693f $X=1.365 $Y=2.23
+ $X2=0 $Y2=0
cc_776 N_A_244_417#_c_1238_n N_A_351_417#_c_1284_n 0.0378599f $X=3.26 $Y=2.59
+ $X2=0 $Y2=0
cc_777 N_A_244_417#_c_1238_n N_A_351_417#_c_1307_n 0.0101437f $X=3.26 $Y=2.59
+ $X2=0 $Y2=0
cc_778 N_A_244_417#_M1014_d N_A_351_417#_c_1288_n 0.00628932f $X=3.285 $Y=2.085
+ $X2=0 $Y2=0
cc_779 N_A_244_417#_c_1238_n N_A_351_417#_c_1288_n 0.0540631f $X=3.26 $Y=2.59
+ $X2=0 $Y2=0
cc_780 N_A_244_417#_c_1238_n A_457_417# 0.00304514f $X=3.26 $Y=2.59 $X2=-0.19
+ $Y2=1.655
cc_781 N_A_351_417#_c_1284_n A_457_417# 0.00117218f $X=2.475 $Y=2.195 $X2=-0.19
+ $Y2=-0.245
cc_782 N_A_351_417#_c_1278_n N_VGND_c_1414_n 9.82691e-19 $X=2.56 $Y=2.065 $X2=0
+ $Y2=0
cc_783 N_A_351_417#_c_1283_n N_VGND_c_1414_n 0.0151116f $X=2.56 $Y=0.82 $X2=0
+ $Y2=0
cc_784 N_A_351_417#_c_1283_n N_VGND_c_1423_n 0.00893874f $X=2.56 $Y=0.82 $X2=0
+ $Y2=0
cc_785 N_A_351_417#_c_1283_n N_VGND_c_1431_n 0.0115756f $X=2.56 $Y=0.82 $X2=0
+ $Y2=0
cc_786 N_A_351_417#_c_1279_n N_A_1160_155#_c_1545_n 0.0235109f $X=6.295 $Y=1.715
+ $X2=0 $Y2=0
cc_787 N_A_351_417#_c_1281_n N_A_1160_155#_c_1545_n 0.0135022f $X=6.38 $Y=0.7
+ $X2=0 $Y2=0
cc_788 N_A_351_417#_c_1280_n N_A_1160_155#_c_1546_n 0.0642913f $X=7.07 $Y=0.7
+ $X2=0 $Y2=0
cc_789 N_A_351_417#_c_1281_n N_A_1160_155#_c_1546_n 0.0128424f $X=6.38 $Y=0.7
+ $X2=0 $Y2=0
cc_790 N_A_351_417#_c_1280_n N_A_1160_155#_c_1548_n 0.0110827f $X=7.07 $Y=0.7
+ $X2=0 $Y2=0
cc_791 N_A_351_417#_c_1282_n N_A_1160_155#_c_1548_n 0.011388f $X=7.155 $Y=0.97
+ $X2=0 $Y2=0
cc_792 N_Q_c_1383_n N_VGND_c_1419_n 0.0175456f $X=12.85 $Y=0.555 $X2=0 $Y2=0
cc_793 N_Q_c_1383_n N_VGND_c_1426_n 0.0186721f $X=12.85 $Y=0.555 $X2=0 $Y2=0
cc_794 N_Q_c_1383_n N_VGND_c_1431_n 0.0140413f $X=12.85 $Y=0.555 $X2=0 $Y2=0
cc_795 N_VGND_c_1416_n N_A_1160_155#_c_1546_n 0.011323f $X=8.245 $Y=0.55 $X2=0
+ $Y2=0
cc_796 N_VGND_c_1425_n N_A_1160_155#_c_1546_n 0.10965f $X=8.08 $Y=0 $X2=0 $Y2=0
cc_797 N_VGND_c_1431_n N_A_1160_155#_c_1546_n 0.0599641f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_798 N_VGND_c_1425_n N_A_1160_155#_c_1547_n 0.0168491f $X=8.08 $Y=0 $X2=0
+ $Y2=0
cc_799 N_VGND_c_1431_n N_A_1160_155#_c_1547_n 0.00867615f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_800 N_VGND_c_1416_n N_A_1160_155#_c_1548_n 0.0115783f $X=8.245 $Y=0.55 $X2=0
+ $Y2=0
cc_801 N_VGND_c_1417_n N_A_1910_155#_c_1582_n 0.0069708f $X=11.505 $Y=0.555
+ $X2=0 $Y2=0
cc_802 N_VGND_c_1420_n N_A_1910_155#_c_1582_n 0.00427436f $X=11.34 $Y=0 $X2=0
+ $Y2=0
cc_803 N_VGND_c_1431_n N_A_1910_155#_c_1582_n 0.00848415f $X=13.68 $Y=0 $X2=0
+ $Y2=0
cc_804 N_VGND_c_1417_n N_A_1910_155#_c_1584_n 0.011122f $X=11.505 $Y=0.555 $X2=0
+ $Y2=0
cc_805 N_VGND_c_1420_n N_A_1910_155#_c_1584_n 0.0119522f $X=11.34 $Y=0 $X2=0
+ $Y2=0
cc_806 N_VGND_c_1431_n N_A_1910_155#_c_1584_n 0.00918135f $X=13.68 $Y=0 $X2=0
+ $Y2=0
