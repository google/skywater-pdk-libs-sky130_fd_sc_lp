* NGSPICE file created from sky130_fd_sc_lp__a22oi_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a22oi_m A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 a_39_496# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=3.822e+11p pd=4.34e+06u as=1.176e+11p ps=1.4e+06u
M1001 VPWR A1 a_39_496# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_314_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.659e+11p ps=1.63e+06u
M1003 Y B1 a_133_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 VGND A2 a_314_47# VNB nshort w=420000u l=150000u
+  ad=2.52e+11p pd=2.88e+06u as=0p ps=0u
M1005 Y B2 a_39_496# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1006 a_39_496# B1 Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_133_47# B2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

