# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nor4bb_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nor4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.195000 1.185000 6.635000 1.515000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.185000 4.715000 1.515000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.580000 0.885000 2.250000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 1.580000 1.420000 2.500000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.293600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.705000 1.675000 4.230000 1.845000 ;
        RECT 2.705000 1.845000 3.035000 2.735000 ;
        RECT 2.775000 0.255000 2.965000 0.995000 ;
        RECT 2.775000 0.995000 5.165000 1.015000 ;
        RECT 2.775000 1.015000 4.230000 1.165000 ;
        RECT 3.635000 0.255000 3.825000 0.840000 ;
        RECT 3.635000 0.840000 5.165000 0.995000 ;
        RECT 3.995000 1.165000 4.230000 1.675000 ;
        RECT 4.885000 1.015000 5.165000 1.065000 ;
        RECT 4.885000 1.065000 6.025000 1.235000 ;
        RECT 4.975000 0.255000 5.165000 0.840000 ;
        RECT 5.835000 0.255000 6.025000 1.065000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.720000 0.085000 ;
        RECT 0.615000  0.085000 0.955000 1.070000 ;
        RECT 2.275000  0.085000 2.605000 0.490000 ;
        RECT 3.135000  0.085000 3.465000 0.825000 ;
        RECT 3.995000  0.085000 4.805000 0.670000 ;
        RECT 5.335000  0.085000 5.665000 0.885000 ;
        RECT 6.195000  0.085000 6.525000 1.015000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.720000 3.415000 ;
        RECT 0.635000 2.670000 1.305000 3.245000 ;
        RECT 5.845000 2.025000 6.175000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.185000 0.865000 0.435000 1.240000 ;
      RECT 0.185000 1.240000 1.295000 1.410000 ;
      RECT 0.185000 1.410000 0.435000 2.605000 ;
      RECT 0.185000 2.605000 0.465000 2.935000 ;
      RECT 1.125000 0.660000 2.555000 0.830000 ;
      RECT 1.125000 0.830000 1.295000 1.240000 ;
      RECT 1.475000 1.000000 2.205000 1.260000 ;
      RECT 1.475000 2.670000 1.975000 3.000000 ;
      RECT 1.805000 1.260000 2.205000 1.600000 ;
      RECT 1.805000 1.600000 1.975000 2.670000 ;
      RECT 2.275000 1.755000 2.535000 2.905000 ;
      RECT 2.275000 2.905000 3.415000 3.075000 ;
      RECT 2.385000 0.830000 2.555000 1.335000 ;
      RECT 2.385000 1.335000 3.825000 1.505000 ;
      RECT 3.205000 2.015000 4.365000 2.185000 ;
      RECT 3.205000 2.185000 3.415000 2.905000 ;
      RECT 3.585000 2.355000 3.915000 2.905000 ;
      RECT 3.585000 2.905000 5.315000 3.075000 ;
      RECT 4.085000 2.185000 4.365000 2.735000 ;
      RECT 4.555000 1.685000 6.605000 1.855000 ;
      RECT 4.555000 1.855000 4.815000 2.735000 ;
      RECT 4.985000 2.025000 5.315000 2.905000 ;
      RECT 5.485000 1.855000 5.675000 3.075000 ;
      RECT 6.345000 1.855000 6.605000 3.075000 ;
  END
END sky130_fd_sc_lp__nor4bb_2
