* File: sky130_fd_sc_lp__o31a_lp.pex.spice
* Created: Wed Sep  2 10:24:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31A_LP%B1 3 7 11 12 13 14 18 19
c38 12 0 1.55458e-19 $X=0.605 $Y=1.795
r39 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.29 $X2=0.605 $Y2=1.29
r40 13 14 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.622 $Y=1.295
+ $X2=0.622 $Y2=1.665
r41 13 19 0.157869 $w=3.63e-07 $l=5e-09 $layer=LI1_cond $X=0.622 $Y=1.295
+ $X2=0.622 $Y2=1.29
r42 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.605 $Y=1.63
+ $X2=0.605 $Y2=1.29
r43 11 12 31.2043 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.63
+ $X2=0.605 $Y2=1.795
r44 10 18 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.125
+ $X2=0.605 $Y2=1.29
r45 7 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.625 $Y=0.495
+ $X2=0.625 $Y2=1.125
r46 3 12 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.625 $Y=2.55
+ $X2=0.625 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_LP%A3 3 7 11 12 13 14 18
c47 12 0 1.9714e-19 $X=1.145 $Y=1.795
r48 13 14 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.15 $Y=1.29
+ $X2=1.15 $Y2=1.665
r49 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.145
+ $Y=1.29 $X2=1.145 $Y2=1.29
r50 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.145 $Y=1.63
+ $X2=1.145 $Y2=1.29
r51 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.63
+ $X2=1.145 $Y2=1.795
r52 10 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.125
+ $X2=1.145 $Y2=1.29
r53 7 12 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.155 $Y=2.55
+ $X2=1.155 $Y2=1.795
r54 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.085 $Y=0.495
+ $X2=1.085 $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_LP%A2 3 7 11 12 13 14 18
c44 3 0 1.92213e-19 $X=1.675 $Y=2.55
r45 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.295
+ $X2=1.685 $Y2=1.665
r46 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.685
+ $Y=1.335 $X2=1.685 $Y2=1.335
r47 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.685 $Y=1.675
+ $X2=1.685 $Y2=1.335
r48 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.685 $Y=1.675
+ $X2=1.685 $Y2=1.84
r49 10 18 40.0117 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.685 $Y=1.17
+ $X2=1.685 $Y2=1.335
r50 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.645 $Y=0.495
+ $X2=1.645 $Y2=1.17
r51 3 12 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.675 $Y=2.55
+ $X2=1.675 $Y2=1.84
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_LP%A1 3 8 10 11 13 14 15 16 17 21
r49 16 17 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.217 $Y=1.295
+ $X2=2.217 $Y2=1.665
r50 16 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.225
+ $Y=1.335 $X2=2.225 $Y2=1.335
r51 14 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.225 $Y=1.675
+ $X2=2.225 $Y2=1.335
r52 14 15 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.675
+ $X2=2.225 $Y2=1.84
r53 13 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.17
+ $X2=2.225 $Y2=1.335
r54 11 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.135 $Y=0.93
+ $X2=2.135 $Y2=1.17
r55 10 11 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=2.105 $Y=0.78
+ $X2=2.105 $Y2=0.93
r56 8 15 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.215 $Y=2.55
+ $X2=2.215 $Y2=1.84
r57 3 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.075 $Y=0.495
+ $X2=2.075 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_LP%A_37_57# 1 2 7 9 12 16 19 21 23 24 25 28 32
+ 36 37 40 44 46 47
c93 46 0 3.47671e-19 $X=0.89 $Y=2.082
c94 32 0 1.9714e-19 $X=2.575 $Y=2.105
r95 41 44 4.03026 $w=4.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.175 $Y=0.495
+ $X2=0.33 $Y2=0.495
r96 40 47 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.66 $Y=2.02
+ $X2=2.66 $Y2=1.6
r97 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.765
+ $Y=1.095 $X2=2.765 $Y2=1.095
r98 34 47 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=2.747 $Y=1.428
+ $X2=2.747 $Y2=1.6
r99 34 36 11.1236 $w=3.43e-07 $l=3.33e-07 $layer=LI1_cond $X=2.747 $Y=1.428
+ $X2=2.747 $Y2=1.095
r100 33 46 8.61065 $w=1.7e-07 $l=1.76125e-07 $layer=LI1_cond $X=1.055 $Y=2.105
+ $X2=0.89 $Y2=2.082
r101 32 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=2.105
+ $X2=2.66 $Y2=2.02
r102 32 33 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=2.575 $Y=2.105
+ $X2=1.055 $Y2=2.105
r103 28 30 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.89 $Y=2.195
+ $X2=0.89 $Y2=2.9
r104 26 46 0.89609 $w=3.3e-07 $l=1.08e-07 $layer=LI1_cond $X=0.89 $Y=2.19
+ $X2=0.89 $Y2=2.082
r105 26 28 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.89 $Y=2.19
+ $X2=0.89 $Y2=2.195
r106 24 46 8.61065 $w=1.7e-07 $l=1.75656e-07 $layer=LI1_cond $X=0.725 $Y=2.06
+ $X2=0.89 $Y2=2.082
r107 24 25 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.725 $Y=2.06
+ $X2=0.26 $Y2=2.06
r108 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.175 $Y=1.975
+ $X2=0.26 $Y2=2.06
r109 22 41 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.175 $Y=0.725
+ $X2=0.175 $Y2=0.495
r110 22 23 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=0.175 $Y=0.725
+ $X2=0.175 $Y2=1.975
r111 20 37 56.8556 $w=3.4e-07 $l=3.35e-07 $layer=POLY_cond $X=2.77 $Y=1.43
+ $X2=2.77 $Y2=1.095
r112 20 21 31.7294 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=2.77 $Y=1.43
+ $X2=2.77 $Y2=1.6
r113 19 37 28.0035 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=0.93
+ $X2=2.77 $Y2=1.095
r114 12 21 236.031 $w=2.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.745 $Y=2.55
+ $X2=2.745 $Y2=1.6
r115 7 19 26.4004 $w=3.4e-07 $l=1.5e-07 $layer=POLY_cond $X=2.685 $Y=0.78
+ $X2=2.685 $Y2=0.93
r116 7 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.865 $Y=0.78
+ $X2=2.865 $Y2=0.495
r117 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.505 $Y=0.78
+ $X2=2.505 $Y2=0.495
r118 2 30 400 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=0.75
+ $Y=2.05 $X2=0.89 $Y2=2.9
r119 2 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.75
+ $Y=2.05 $X2=0.89 $Y2=2.195
r120 1 44 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.285 $X2=0.33 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_LP%VPWR 1 2 7 9 13 16 17 18 28 29
r35 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 26 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 23 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 20 32 4.57961 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.262 $Y2=3.33
r43 20 22 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 18 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 18 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 16 25 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.48 $Y2=3.33
r48 15 28 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.48 $Y2=3.33
r50 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=3.245
+ $X2=2.48 $Y2=3.33
r51 11 13 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.48 $Y=3.245
+ $X2=2.48 $Y2=2.535
r52 7 32 3.18657 $w=3.3e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.262 $Y2=3.33
r53 7 9 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.36 $Y=3.245
+ $X2=0.36 $Y2=2.49
r54 2 13 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=2.34
+ $Y=2.05 $X2=2.48 $Y2=2.535
r55 1 9 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=0.215
+ $Y=2.05 $X2=0.36 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_LP%X 1 2 10 13 14 15 32 34
r19 20 34 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=3.097 $Y=2.092
+ $X2=3.097 $Y2=2.035
r20 15 29 4.17552 $w=3.43e-07 $l=1.25e-07 $layer=LI1_cond $X=3.097 $Y=2.775
+ $X2=3.097 $Y2=2.9
r21 14 15 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.097 $Y=2.405
+ $X2=3.097 $Y2=2.775
r22 14 23 7.01487 $w=3.43e-07 $l=2.1e-07 $layer=LI1_cond $X=3.097 $Y=2.405
+ $X2=3.097 $Y2=2.195
r23 13 34 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=3.097 $Y=2.021
+ $X2=3.097 $Y2=2.035
r24 13 32 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=3.097 $Y=2.021
+ $X2=3.097 $Y2=1.92
r25 13 23 2.97297 $w=3.43e-07 $l=8.9e-08 $layer=LI1_cond $X=3.097 $Y=2.106
+ $X2=3.097 $Y2=2.195
r26 13 20 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=3.097 $Y=2.106
+ $X2=3.097 $Y2=2.092
r27 12 32 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=3.185 $Y=0.725
+ $X2=3.185 $Y2=1.92
r28 10 12 10.6092 $w=3.53e-07 $l=2.3e-07 $layer=LI1_cond $X=3.092 $Y=0.495
+ $X2=3.092 $Y2=0.725
r29 2 29 400 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=2.05 $X2=3.01 $Y2=2.9
r30 2 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.87
+ $Y=2.05 $X2=3.01 $Y2=2.195
r31 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.285 $X2=3.08 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_LP%A_140_57# 1 2 9 11 12 15
r35 13 15 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.82 $Y=0.775
+ $X2=1.82 $Y2=0.495
r36 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.695 $Y=0.86
+ $X2=1.82 $Y2=0.775
r37 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.695 $Y=0.86
+ $X2=1.005 $Y2=0.86
r38 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.84 $Y=0.775
+ $X2=1.005 $Y2=0.86
r39 7 9 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.84 $Y=0.775 $X2=0.84
+ $Y2=0.495
r40 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.285 $X2=1.86 $Y2=0.495
r41 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.7
+ $Y=0.285 $X2=0.84 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_LP%VGND 1 2 9 11 15 17 19 26 27 30 33
r42 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r43 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 27 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r45 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.29
+ $Y2=0
r47 24 26 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=3.12
+ $Y2=0
r48 22 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r49 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.35
+ $Y2=0
r51 19 21 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=0.24
+ $Y2=0
r52 17 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r53 17 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0
r55 13 15 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0.495
r56 12 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.35
+ $Y2=0
r57 11 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.29
+ $Y2=0
r58 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=1.515
+ $Y2=0
r59 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=0.085 $X2=1.35
+ $Y2=0
r60 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0.43
r61 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.15
+ $Y=0.285 $X2=2.29 $Y2=0.495
r62 1 9 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.285 $X2=1.35 $Y2=0.43
.ends

