* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 Y a_223_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND A_N a_223_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y a_223_49# a_357_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_614_47# a_27_373# a_357_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR A_N a_223_49# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR a_27_373# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_357_47# a_223_49# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_27_373# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_357_47# a_27_373# a_614_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_27_373# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 VPWR a_223_49# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Y a_27_373# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_821_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VGND D a_821_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_821_47# C a_614_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_614_47# C a_821_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
