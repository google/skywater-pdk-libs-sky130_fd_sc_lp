* File: sky130_fd_sc_lp__a41o_lp.pex.spice
* Created: Wed Sep  2 09:29:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41O_LP%A4 3 7 11 12 13 16 17
r35 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=0.99 $X2=0.27 $Y2=0.99
r36 13 17 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=0.99
r37 12 16 32.6516 $w=4.65e-07 $l=2.73e-07 $layer=POLY_cond $X=0.337 $Y=1.263
+ $X2=0.337 $Y2=0.99
r38 11 16 1.79404 $w=4.65e-07 $l=1.5e-08 $layer=POLY_cond $X=0.337 $Y=0.975
+ $X2=0.337 $Y2=0.99
r39 10 11 45.5629 $w=4.65e-07 $l=1.5e-07 $layer=POLY_cond $X=0.372 $Y=0.825
+ $X2=0.372 $Y2=0.975
r40 7 10 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.565 $Y=0.445
+ $X2=0.565 $Y2=0.825
r41 1 12 44.235 $w=3.89e-07 $l=4.49116e-07 $layer=POLY_cond $X=0.545 $Y=1.62
+ $X2=0.337 $Y2=1.263
r42 1 3 229.82 $w=2.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.545 $Y=1.62
+ $X2=0.545 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_LP%A3 3 6 9 10 11 12 13 14 19
c47 19 0 2.64121e-20 $X=1.045 $Y=0.93
c48 11 0 6.7672e-20 $X=1.045 $Y=1.435
c49 6 0 7.16571e-20 $X=1.075 $Y=2.545
r50 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.045
+ $Y=0.93 $X2=1.045 $Y2=0.93
r51 14 20 7.33729 $w=5.93e-07 $l=3.65e-07 $layer=LI1_cond $X=0.912 $Y=1.295
+ $X2=0.912 $Y2=0.93
r52 13 20 0.100511 $w=5.93e-07 $l=5e-09 $layer=LI1_cond $X=0.912 $Y=0.925
+ $X2=0.912 $Y2=0.93
r53 12 13 7.4378 $w=5.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.912 $Y=0.555
+ $X2=0.912 $Y2=0.925
r54 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.045 $Y=1.27
+ $X2=1.045 $Y2=0.93
r55 10 11 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=1.27
+ $X2=1.045 $Y2=1.435
r56 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=0.765
+ $X2=1.045 $Y2=0.93
r57 6 11 275.784 $w=2.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.075 $Y=2.545
+ $X2=1.075 $Y2=1.435
r58 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.955 $Y=0.445
+ $X2=0.955 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_LP%A2 3 6 9 10 11 12 13 14 19
c46 11 0 1.08738e-19 $X=1.585 $Y=1.435
c47 6 0 1.01004e-19 $X=1.605 $Y=2.545
r48 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.585
+ $Y=0.93 $X2=1.585 $Y2=0.93
r49 14 20 11.2171 $w=3.73e-07 $l=3.65e-07 $layer=LI1_cond $X=1.607 $Y=1.295
+ $X2=1.607 $Y2=0.93
r50 13 20 0.153659 $w=3.73e-07 $l=5e-09 $layer=LI1_cond $X=1.607 $Y=0.925
+ $X2=1.607 $Y2=0.93
r51 12 13 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.607 $Y=0.555
+ $X2=1.607 $Y2=0.925
r52 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.585 $Y=1.27
+ $X2=1.585 $Y2=0.93
r53 10 11 31.2043 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.27
+ $X2=1.585 $Y2=1.435
r54 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=0.765
+ $X2=1.585 $Y2=0.93
r55 6 11 275.784 $w=2.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.605 $Y=2.545
+ $X2=1.605 $Y2=1.435
r56 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.495 $Y=0.445
+ $X2=1.495 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_LP%A1 3 5 7 11 12 15
c43 12 0 1.76692e-19 $X=2.16 $Y=1.295
c44 7 0 8.40218e-20 $X=2.155 $Y=2.545
c45 5 0 1.88811e-19 $X=2.155 $Y=1.745
r46 12 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.155
+ $Y=1.24 $X2=2.155 $Y2=1.24
r47 11 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.155 $Y=1.58
+ $X2=2.155 $Y2=1.24
r48 10 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.075
+ $X2=2.155 $Y2=1.24
r49 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.745
+ $X2=2.155 $Y2=1.58
r50 5 7 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=2.155 $Y=1.745 $X2=2.155
+ $Y2=2.545
r51 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.065 $Y=0.445
+ $X2=2.065 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_LP%B1 3 7 11 15 16 17 20 21
c51 15 0 1.89903e-19 $X=2.815 $Y=1.225
r52 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.825
+ $Y=1.24 $X2=2.825 $Y2=1.24
r53 17 21 3.3026 $w=6.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.64 $Y=1.41
+ $X2=2.825 $Y2=1.41
r54 16 20 40.6942 $w=4.1e-07 $l=3e-07 $layer=POLY_cond $X=2.865 $Y=1.54
+ $X2=2.865 $Y2=1.24
r55 15 20 2.03471 $w=4.1e-07 $l=1.5e-08 $layer=POLY_cond $X=2.865 $Y=1.225
+ $X2=2.865 $Y2=1.24
r56 5 16 45.5759 $w=3.49e-07 $l=4.10244e-07 $layer=POLY_cond $X=2.685 $Y=1.87
+ $X2=2.865 $Y2=1.54
r57 5 7 167.706 $w=2.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.685 $Y=1.87
+ $X2=2.685 $Y2=2.545
r58 1 15 24.4548 $w=4.1e-07 $l=1.5e-07 $layer=POLY_cond $X=2.815 $Y=1.075
+ $X2=2.815 $Y2=1.225
r59 1 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.995 $Y=1.075
+ $X2=2.995 $Y2=0.445
r60 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.635 $Y=1.075
+ $X2=2.635 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_LP%A_428_47# 1 2 7 9 12 14 16 19 21 22 25 29 30
+ 34 35
c74 35 0 1.72253e-19 $X=3.49 $Y=0.93
c75 30 0 8.40218e-20 $X=3.115 $Y=2.01
r76 35 37 64.3909 $w=5.75e-07 $l=5.05e-07 $layer=POLY_cond $X=3.612 $Y=0.93
+ $X2=3.612 $Y2=1.435
r77 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.49
+ $Y=0.93 $X2=3.49 $Y2=0.93
r78 32 34 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=3.49 $Y=1.925
+ $X2=3.49 $Y2=0.93
r79 31 34 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=3.49 $Y=0.895
+ $X2=3.49 $Y2=0.93
r80 29 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.325 $Y=2.01
+ $X2=3.49 $Y2=1.925
r81 29 30 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.325 $Y=2.01
+ $X2=3.115 $Y2=2.01
r82 25 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.95 $Y=2.19 $X2=2.95
+ $Y2=2.9
r83 23 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.95 $Y=2.095
+ $X2=3.115 $Y2=2.01
r84 23 25 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.95 $Y=2.095
+ $X2=2.95 $Y2=2.19
r85 21 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.325 $Y=0.81
+ $X2=3.49 $Y2=0.895
r86 21 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.325 $Y=0.81
+ $X2=2.585 $Y2=0.81
r87 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.42 $Y=0.725
+ $X2=2.585 $Y2=0.81
r88 17 19 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.42 $Y=0.725
+ $X2=2.42 $Y2=0.47
r89 14 35 30.1985 $w=2.87e-07 $l=2.41814e-07 $layer=POLY_cond $X=3.785 $Y=0.765
+ $X2=3.612 $Y2=0.93
r90 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.785 $Y=0.765
+ $X2=3.785 $Y2=0.445
r91 12 37 275.784 $w=2.5e-07 $l=1.11e-06 $layer=POLY_cond $X=3.775 $Y=2.545
+ $X2=3.775 $Y2=1.435
r92 7 35 30.1985 $w=2.87e-07 $l=2.56562e-07 $layer=POLY_cond $X=3.425 $Y=0.765
+ $X2=3.612 $Y2=0.93
r93 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.425 $Y=0.765
+ $X2=3.425 $Y2=0.445
r94 2 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.045 $X2=2.95 $Y2=2.9
r95 2 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.81
+ $Y=2.045 $X2=2.95 $Y2=2.19
r96 1 19 182 $w=1.7e-07 $l=3.79737e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.235 $X2=2.42 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_LP%A_27_409# 1 2 3 12 16 17 20 24 28 32
c52 32 0 2.56483e-19 $X=1.34 $Y=1.76
c53 24 0 1.93606e-19 $X=2.255 $Y=2.01
c54 16 0 1.01004e-19 $X=1.175 $Y=1.76
r55 32 34 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.34 $Y=1.76
+ $X2=1.34 $Y2=2.01
r56 28 30 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.42 $Y=2.19 $X2=2.42
+ $Y2=2.9
r57 26 28 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.42 $Y=2.095
+ $X2=2.42 $Y2=2.19
r58 25 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=2.01
+ $X2=1.34 $Y2=2.01
r59 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.255 $Y=2.01
+ $X2=2.42 $Y2=2.095
r60 24 25 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.255 $Y=2.01
+ $X2=1.505 $Y2=2.01
r61 20 22 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.34 $Y=2.19 $X2=1.34
+ $Y2=2.9
r62 18 34 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.34 $Y=2.095
+ $X2=1.34 $Y2=2.01
r63 18 20 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.34 $Y=2.095
+ $X2=1.34 $Y2=2.19
r64 16 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=1.76
+ $X2=1.34 $Y2=1.76
r65 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.175 $Y=1.76
+ $X2=0.445 $Y2=1.76
r66 12 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.19 $X2=0.28
+ $Y2=2.9
r67 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.845
+ $X2=0.445 $Y2=1.76
r68 10 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.28 $Y=1.845
+ $X2=0.28 $Y2=2.19
r69 3 30 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=2.045 $X2=2.42 $Y2=2.9
r70 3 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=2.045 $X2=2.42 $Y2=2.19
r71 2 22 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.045 $X2=1.34 $Y2=2.9
r72 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.2
+ $Y=2.045 $X2=1.34 $Y2=2.19
r73 1 14 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r74 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_LP%VPWR 1 2 3 14 20 24 27 28 30 31 32 45 46 49
r53 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r58 37 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r61 34 36 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 32 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 32 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 32 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r65 30 42 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.51 $Y2=3.33
r67 29 45 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=4.08 $Y2=3.33
r68 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=3.51 $Y2=3.33
r69 27 36 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.87 $Y2=3.33
r71 26 39 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.87 $Y2=3.33
r73 22 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.51 $Y=3.245
+ $X2=3.51 $Y2=3.33
r74 22 24 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=3.51 $Y=3.245
+ $X2=3.51 $Y2=2.44
r75 18 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=3.33
r76 18 20 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=2.44
r77 14 17 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.19 $X2=0.81
+ $Y2=2.9
r78 12 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r79 12 17 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.9
r80 3 24 300 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=2 $X=3.365
+ $Y=2.045 $X2=3.51 $Y2=2.44
r81 2 20 300 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=2 $X=1.73
+ $Y=2.045 $X2=1.87 $Y2=2.44
r82 1 17 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.9
r83 1 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_LP%X 1 2 7 8 9 10 11 12 13
r19 13 37 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=4.04 $Y=2.775
+ $X2=4.04 $Y2=2.9
r20 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.04 $Y=2.405
+ $X2=4.04 $Y2=2.775
r21 12 31 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.04 $Y=2.405
+ $X2=4.04 $Y2=2.19
r22 11 31 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.04 $Y=2.035
+ $X2=4.04 $Y2=2.19
r23 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=2.035
r24 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.04 $Y=1.295
+ $X2=4.04 $Y2=1.665
r25 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.04 $Y=0.925 $X2=4.04
+ $Y2=1.295
r26 8 43 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=4.04 $Y=0.925
+ $X2=4.04 $Y2=0.675
r27 7 43 6.54674 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.02 $Y=0.47
+ $X2=4.02 $Y2=0.675
r28 2 37 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=2.045 $X2=4.04 $Y2=2.9
r29 2 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=2.045 $X2=4.04 $Y2=2.19
r30 1 7 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.86
+ $Y=0.235 $X2=4 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A41O_LP%VGND 1 2 7 9 13 15 17 24 25 31
c55 25 0 2.64121e-20 $X=4.08 $Y=0
c56 24 0 1.72253e-19 $X=4.08 $Y=0
r57 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r58 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r59 25 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r60 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r61 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.21
+ $Y2=0
r62 22 24 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=4.08
+ $Y2=0
r63 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r64 20 21 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 18 28 3.93235 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r66 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.72
+ $Y2=0
r67 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.21
+ $Y2=0
r68 17 20 151.684 $w=1.68e-07 $l=2.325e-06 $layer=LI1_cond $X=3.045 $Y=0
+ $X2=0.72 $Y2=0
r69 15 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r70 15 21 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=0.72
+ $Y2=0
r71 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0
r72 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.21 $Y=0.085
+ $X2=3.21 $Y2=0.38
r73 7 28 3.21082 $w=2.5e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.217 $Y2=0
r74 7 9 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.31 $Y2=0.43
r75 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.235 $X2=3.21 $Y2=0.38
r76 1 9 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.235 $X2=0.35 $Y2=0.43
.ends

