* File: sky130_fd_sc_lp__or4_2.pxi.spice
* Created: Wed Sep  2 10:31:56 2020
* 
x_PM_SKY130_FD_SC_LP__OR4_2%D N_D_c_79_n N_D_c_80_n N_D_c_81_n N_D_c_82_n
+ N_D_M1010_g N_D_M1008_g D D D N_D_c_86_n PM_SKY130_FD_SC_LP__OR4_2%D
x_PM_SKY130_FD_SC_LP__OR4_2%C N_C_M1005_g N_C_M1002_g N_C_c_116_n N_C_c_117_n C
+ C C C C N_C_c_118_n N_C_c_119_n PM_SKY130_FD_SC_LP__OR4_2%C
x_PM_SKY130_FD_SC_LP__OR4_2%B N_B_M1001_g N_B_M1000_g N_B_c_159_n N_B_c_160_n B
+ B B B B N_B_c_161_n N_B_c_162_n PM_SKY130_FD_SC_LP__OR4_2%B
x_PM_SKY130_FD_SC_LP__OR4_2%A N_A_M1006_g N_A_M1007_g A A A A N_A_c_205_n
+ N_A_c_206_n A PM_SKY130_FD_SC_LP__OR4_2%A
x_PM_SKY130_FD_SC_LP__OR4_2%A_72_367# N_A_72_367#_M1010_d N_A_72_367#_M1000_d
+ N_A_72_367#_M1008_s N_A_72_367#_c_254_n N_A_72_367#_M1004_g
+ N_A_72_367#_M1003_g N_A_72_367#_c_257_n N_A_72_367#_M1011_g
+ N_A_72_367#_M1009_g N_A_72_367#_c_260_n N_A_72_367#_c_261_n
+ N_A_72_367#_c_290_n N_A_72_367#_c_262_n N_A_72_367#_c_263_n
+ N_A_72_367#_c_297_n N_A_72_367#_c_264_n N_A_72_367#_c_265_n
+ N_A_72_367#_c_266_n N_A_72_367#_c_267_n N_A_72_367#_c_272_n
+ N_A_72_367#_c_268_n PM_SKY130_FD_SC_LP__OR4_2%A_72_367#
x_PM_SKY130_FD_SC_LP__OR4_2%VPWR N_VPWR_M1007_d N_VPWR_M1009_s N_VPWR_c_384_n
+ N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_398_n VPWR N_VPWR_c_387_n
+ N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_383_n PM_SKY130_FD_SC_LP__OR4_2%VPWR
x_PM_SKY130_FD_SC_LP__OR4_2%X N_X_M1003_s N_X_M1004_d X X X X X X X N_X_c_417_n
+ X PM_SKY130_FD_SC_LP__OR4_2%X
x_PM_SKY130_FD_SC_LP__OR4_2%VGND N_VGND_M1010_s N_VGND_M1002_d N_VGND_M1006_d
+ N_VGND_M1011_d N_VGND_c_438_n N_VGND_c_439_n N_VGND_c_440_n N_VGND_c_441_n
+ N_VGND_c_442_n N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n VGND
+ N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n N_VGND_c_449_n
+ PM_SKY130_FD_SC_LP__OR4_2%VGND
cc_1 VNB N_D_c_79_n 0.0192249f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.915
cc_2 VNB N_D_c_80_n 0.0189035f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.915
cc_3 VNB N_D_c_81_n 0.0194222f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.435
cc_4 VNB N_D_c_82_n 0.0191156f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.435
cc_5 VNB N_D_M1010_g 0.0242448f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.455
cc_6 VNB N_D_M1008_g 0.00875446f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.045
cc_7 VNB D 0.0379652f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_8 VNB N_D_c_86_n 0.0285789f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_9 VNB N_C_M1002_g 0.0297324f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.455
cc_10 VNB N_C_c_116_n 0.0228454f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.045
cc_11 VNB N_C_c_117_n 0.00896639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C_c_118_n 0.0170727f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=0.925
cc_13 VNB N_C_c_119_n 0.00390733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_M1000_g 0.0296024f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.455
cc_15 VNB N_B_c_159_n 0.0209044f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.045
cc_16 VNB N_B_c_160_n 0.00895555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_c_161_n 0.0152775f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=0.925
cc_18 VNB N_B_c_162_n 0.00584667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_M1006_g 0.0473827f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.435
cc_20 VNB N_A_c_205_n 0.0219669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_206_n 0.00445194f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_22 VNB N_A_72_367#_c_254_n 0.0331201f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.045
cc_23 VNB N_A_72_367#_M1004_g 0.00224613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_72_367#_M1003_g 0.0238474f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_25 VNB N_A_72_367#_c_257_n 0.0102961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_72_367#_M1011_g 0.0287405f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_27 VNB N_A_72_367#_M1009_g 0.0175949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_72_367#_c_260_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_72_367#_c_261_n 0.00719691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_72_367#_c_262_n 0.00810487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_72_367#_c_263_n 0.0132623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_72_367#_c_264_n 0.00717429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_72_367#_c_265_n 0.00486896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_72_367#_c_266_n 0.00688826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_72_367#_c_267_n 0.00200012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_72_367#_c_268_n 0.00896796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_383_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB X 0.00189758f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.51
cc_39 VNB N_X_c_417_n 3.86013e-19 $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=0.925
cc_40 VNB X 0.00481904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_438_n 0.0158051f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_42 VNB N_VGND_c_439_n 0.00463806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_440_n 0.0116069f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_44 VNB N_VGND_c_441_n 0.0498891f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_45 VNB N_VGND_c_442_n 0.0109511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_443_n 0.00529368f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=1.295
cc_47 VNB N_VGND_c_444_n 0.0148029f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=1.665
cc_48 VNB N_VGND_c_445_n 0.00630897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_446_n 0.0140401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_447_n 0.0149435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_448_n 0.0137896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_449_n 0.210677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_D_M1008_g 0.029498f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.045
cc_54 VPB D 0.0146328f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_55 VPB N_C_M1005_g 0.018465f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.435
cc_56 VPB N_C_c_117_n 0.00636408f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_C_c_119_n 0.0378018f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_B_M1001_g 0.0187723f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.435
cc_59 VPB N_B_c_160_n 0.0069088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_B_c_162_n 0.0219286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_M1007_g 0.0202303f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.455
cc_62 VPB A 0.00488318f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.51
cc_63 VPB A 0.0153998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_c_205_n 0.00788628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_c_206_n 5.0252e-19 $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_66 VPB A 0.00407259f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_72_367#_M1004_g 0.0236089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_72_367#_M1009_g 0.0272796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_72_367#_c_261_n 0.00379278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_72_367#_c_272_n 0.0131138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_384_n 0.0150635f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.045
cc_72 VPB N_VPWR_c_385_n 0.011581f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.045
cc_73 VPB N_VPWR_c_386_n 0.0653514f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.99
cc_74 VPB N_VPWR_c_387_n 0.0747893f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_75 VPB N_VPWR_c_388_n 0.0149952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_389_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_383_n 0.112287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB X 0.00478821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 N_D_M1010_g N_C_M1002_g 0.0229713f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_80 N_D_c_81_n N_C_c_116_n 0.0295647f $X=0.625 $Y=1.435 $X2=0 $Y2=0
cc_81 N_D_M1008_g N_C_c_117_n 0.0295647f $X=0.7 $Y=2.045 $X2=0 $Y2=0
cc_82 N_D_c_86_n N_C_c_118_n 0.00280064f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_83 N_D_c_81_n N_C_c_119_n 0.00403263f $X=0.625 $Y=1.435 $X2=0 $Y2=0
cc_84 N_D_c_79_n N_A_72_367#_c_261_n 0.00612458f $X=0.625 $Y=0.915 $X2=0 $Y2=0
cc_85 N_D_c_81_n N_A_72_367#_c_261_n 0.0100781f $X=0.625 $Y=1.435 $X2=0 $Y2=0
cc_86 N_D_M1008_g N_A_72_367#_c_261_n 0.0125178f $X=0.7 $Y=2.045 $X2=0 $Y2=0
cc_87 D N_A_72_367#_c_261_n 0.0627012f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_88 N_D_c_86_n N_A_72_367#_c_261_n 0.00202077f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_89 N_D_c_79_n N_A_72_367#_c_263_n 0.0054837f $X=0.625 $Y=0.915 $X2=0 $Y2=0
cc_90 N_D_c_81_n N_A_72_367#_c_263_n 4.31636e-19 $X=0.625 $Y=1.435 $X2=0 $Y2=0
cc_91 N_D_M1010_g N_A_72_367#_c_263_n 0.010317f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_92 D N_A_72_367#_c_263_n 0.0119075f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_93 N_D_c_81_n N_A_72_367#_c_272_n 2.41657e-19 $X=0.625 $Y=1.435 $X2=0 $Y2=0
cc_94 N_D_c_82_n N_A_72_367#_c_272_n 0.00542222f $X=0.435 $Y=1.435 $X2=0 $Y2=0
cc_95 N_D_M1008_g N_A_72_367#_c_272_n 0.00810816f $X=0.7 $Y=2.045 $X2=0 $Y2=0
cc_96 D N_A_72_367#_c_272_n 0.00385066f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_97 N_D_c_79_n N_VGND_c_438_n 4.07435e-19 $X=0.625 $Y=0.915 $X2=0 $Y2=0
cc_98 N_D_c_80_n N_VGND_c_438_n 0.0070146f $X=0.435 $Y=0.915 $X2=0 $Y2=0
cc_99 N_D_M1010_g N_VGND_c_438_n 0.00722672f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_100 D N_VGND_c_438_n 0.00504474f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_101 D N_VGND_c_442_n 0.00340198f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_102 N_D_M1010_g N_VGND_c_444_n 0.00415294f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_103 N_D_M1010_g N_VGND_c_449_n 0.00496559f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_104 D N_VGND_c_449_n 0.00623922f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_105 N_C_M1005_g N_B_M1001_g 0.0203646f $X=1.06 $Y=2.045 $X2=0 $Y2=0
cc_106 N_C_M1002_g N_B_M1000_g 0.0225376f $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_107 N_C_c_116_n N_B_c_159_n 0.0144008f $X=1.15 $Y=1.51 $X2=0 $Y2=0
cc_108 N_C_c_117_n N_B_c_160_n 0.0144008f $X=1.15 $Y=1.675 $X2=0 $Y2=0
cc_109 N_C_c_118_n N_B_c_161_n 0.0144008f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_110 N_C_c_119_n N_B_c_161_n 0.00473631f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_111 N_C_M1005_g N_B_c_162_n 9.4204e-19 $X=1.06 $Y=2.045 $X2=0 $Y2=0
cc_112 N_C_c_118_n N_B_c_162_n 0.0033482f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_113 N_C_c_119_n N_B_c_162_n 0.139491f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_114 N_C_M1002_g N_A_72_367#_c_261_n 8.72084e-19 $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_115 N_C_c_116_n N_A_72_367#_c_261_n 0.00165706f $X=1.15 $Y=1.51 $X2=0 $Y2=0
cc_116 N_C_c_118_n N_A_72_367#_c_261_n 0.00594168f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_117 N_C_c_119_n N_A_72_367#_c_261_n 0.0418294f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_118 N_C_M1002_g N_A_72_367#_c_290_n 0.00674994f $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_119 N_C_M1002_g N_A_72_367#_c_262_n 0.00907497f $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_120 N_C_c_118_n N_A_72_367#_c_262_n 0.00292201f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_121 N_C_c_119_n N_A_72_367#_c_262_n 0.0151653f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_122 N_C_M1002_g N_A_72_367#_c_263_n 0.00522893f $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_123 N_C_c_118_n N_A_72_367#_c_263_n 0.00197525f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_124 N_C_c_119_n N_A_72_367#_c_263_n 0.00667886f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_125 N_C_M1002_g N_A_72_367#_c_297_n 5.77015e-19 $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_126 N_C_M1005_g N_A_72_367#_c_272_n 7.85707e-19 $X=1.06 $Y=2.045 $X2=0 $Y2=0
cc_127 N_C_c_119_n N_A_72_367#_c_272_n 0.0148391f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_128 N_C_c_119_n A_227_367# 0.00426898f $X=1.15 $Y=1.17 $X2=-0.19 $Y2=-0.245
cc_129 N_C_c_119_n N_VPWR_c_387_n 0.0149923f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_130 N_C_c_119_n N_VPWR_c_383_n 0.0132441f $X=1.15 $Y=1.17 $X2=0 $Y2=0
cc_131 N_C_M1002_g N_VGND_c_438_n 4.46421e-19 $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_132 N_C_M1002_g N_VGND_c_439_n 0.00314256f $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_133 N_C_M1002_g N_VGND_c_444_n 0.00405108f $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_134 N_C_M1002_g N_VGND_c_449_n 0.0060424f $X=1.13 $Y=0.455 $X2=0 $Y2=0
cc_135 N_B_M1000_g N_A_M1006_g 0.0231594f $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_136 N_B_c_161_n N_A_M1006_g 0.0210108f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_137 N_B_c_162_n N_A_M1006_g 0.00128313f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_138 N_B_M1001_g N_A_M1007_g 0.0203617f $X=1.6 $Y=2.045 $X2=0 $Y2=0
cc_139 N_B_c_162_n N_A_M1007_g 0.00233528f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_140 N_B_M1001_g A 0.00177964f $X=1.6 $Y=2.045 $X2=0 $Y2=0
cc_141 N_B_c_162_n A 0.104217f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_142 N_B_c_159_n N_A_c_205_n 0.0210108f $X=1.69 $Y=1.51 $X2=0 $Y2=0
cc_143 N_B_c_162_n N_A_c_205_n 3.39391e-19 $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_144 N_B_c_159_n N_A_c_206_n 0.00189478f $X=1.69 $Y=1.51 $X2=0 $Y2=0
cc_145 N_B_c_162_n N_A_c_206_n 0.0255055f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_146 N_B_M1000_g N_A_72_367#_c_290_n 5.86431e-19 $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_147 N_B_M1000_g N_A_72_367#_c_262_n 0.00929679f $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_148 N_B_c_161_n N_A_72_367#_c_262_n 7.55836e-19 $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_149 N_B_c_162_n N_A_72_367#_c_262_n 0.0233692f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_150 N_B_M1000_g N_A_72_367#_c_297_n 0.00648647f $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_151 N_B_M1000_g N_A_72_367#_c_264_n 0.00284619f $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_152 N_B_c_161_n N_A_72_367#_c_264_n 0.00119119f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_153 N_B_M1000_g N_A_72_367#_c_265_n 0.00386056f $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_154 N_B_c_162_n N_A_72_367#_c_265_n 7.37894e-19 $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_155 N_B_c_161_n N_A_72_367#_c_267_n 0.00108182f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_156 N_B_c_162_n N_A_72_367#_c_267_n 0.0142533f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_157 N_B_c_162_n A_335_367# 0.00366165f $X=1.69 $Y=1.17 $X2=-0.19 $Y2=-0.245
cc_158 N_B_c_162_n N_VPWR_c_387_n 0.0129272f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_159 N_B_c_162_n N_VPWR_c_383_n 0.0114198f $X=1.69 $Y=1.17 $X2=0 $Y2=0
cc_160 N_B_M1000_g N_VGND_c_439_n 0.00317866f $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_161 N_B_M1000_g N_VGND_c_446_n 0.00408645f $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_162 N_B_M1000_g N_VGND_c_448_n 4.90419e-19 $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_163 N_B_M1000_g N_VGND_c_449_n 0.00607192f $X=1.71 $Y=0.455 $X2=0 $Y2=0
cc_164 N_A_M1006_g N_A_72_367#_c_254_n 0.00160957f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_165 N_A_c_205_n N_A_72_367#_c_254_n 0.0175254f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_166 N_A_c_206_n N_A_72_367#_c_254_n 3.03886e-19 $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_167 N_A_M1007_g N_A_72_367#_M1004_g 0.00846661f $X=2.14 $Y=2.045 $X2=0 $Y2=0
cc_168 A N_A_72_367#_M1004_g 0.0028849f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A_c_205_n N_A_72_367#_M1004_g 0.00140339f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A_c_206_n N_A_72_367#_M1004_g 2.25808e-19 $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_171 A N_A_72_367#_M1004_g 0.00115795f $X=2.16 $Y=2.405 $X2=0 $Y2=0
cc_172 N_A_M1006_g N_A_72_367#_M1003_g 0.00777245f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_173 N_A_M1006_g N_A_72_367#_c_264_n 0.00991177f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_174 N_A_M1006_g N_A_72_367#_c_265_n 0.00611924f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_175 N_A_c_205_n N_A_72_367#_c_266_n 0.00249308f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_176 N_A_c_206_n N_A_72_367#_c_266_n 0.00821009f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A_M1006_g N_A_72_367#_c_267_n 0.00823792f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_178 N_A_c_205_n N_A_72_367#_c_267_n 0.00161905f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A_c_206_n N_A_72_367#_c_267_n 0.0220067f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A_M1006_g N_A_72_367#_c_268_n 0.00303091f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_181 N_A_c_205_n N_A_72_367#_c_268_n 0.00108451f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A_c_206_n N_A_72_367#_c_268_n 0.0198058f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_183 A A_335_367# 0.00377917f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_184 N_A_M1007_g N_VPWR_c_384_n 8.49077e-19 $X=2.14 $Y=2.045 $X2=0 $Y2=0
cc_185 A N_VPWR_c_384_n 0.00731158f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_186 A N_VPWR_c_384_n 0.0513971f $X=2.16 $Y=2.405 $X2=0 $Y2=0
cc_187 N_A_M1007_g N_VPWR_c_398_n 0.00140651f $X=2.14 $Y=2.045 $X2=0 $Y2=0
cc_188 A N_VPWR_c_387_n 0.0143401f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_189 A N_VPWR_c_383_n 0.0126828f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_190 N_A_c_206_n X 0.00168656f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A_M1006_g N_VGND_c_446_n 0.00348975f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_192 N_A_M1006_g N_VGND_c_448_n 0.00976192f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_193 N_A_M1006_g N_VGND_c_449_n 0.00417764f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_194 N_A_72_367#_M1004_g N_VPWR_c_384_n 0.0177296f $X=2.905 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_72_367#_M1009_g N_VPWR_c_386_n 0.00763511f $X=3.34 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A_72_367#_c_254_n N_VPWR_c_398_n 0.00151275f $X=2.905 $Y=1.615 $X2=0
+ $Y2=0
cc_197 N_A_72_367#_M1004_g N_VPWR_c_398_n 0.00956649f $X=2.905 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A_72_367#_M1009_g N_VPWR_c_398_n 8.07815e-19 $X=3.34 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A_72_367#_c_266_n N_VPWR_c_398_n 0.00469563f $X=2.575 $Y=1.1 $X2=0
+ $Y2=0
cc_200 N_A_72_367#_c_268_n N_VPWR_c_398_n 0.0168248f $X=2.715 $Y=1.1 $X2=0 $Y2=0
cc_201 N_A_72_367#_M1004_g N_VPWR_c_388_n 0.00486043f $X=2.905 $Y=2.465 $X2=0
+ $Y2=0
cc_202 N_A_72_367#_M1009_g N_VPWR_c_388_n 0.00585385f $X=3.34 $Y=2.465 $X2=0
+ $Y2=0
cc_203 N_A_72_367#_M1004_g N_VPWR_c_383_n 0.00826027f $X=2.905 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_A_72_367#_M1009_g N_VPWR_c_383_n 0.0115045f $X=3.34 $Y=2.465 $X2=0
+ $Y2=0
cc_205 N_A_72_367#_M1003_g X 0.00163925f $X=2.91 $Y=0.665 $X2=0 $Y2=0
cc_206 N_A_72_367#_c_268_n X 0.0103037f $X=2.715 $Y=1.1 $X2=0 $Y2=0
cc_207 N_A_72_367#_M1003_g N_X_c_417_n 7.31235e-19 $X=2.91 $Y=0.665 $X2=0 $Y2=0
cc_208 N_A_72_367#_M1011_g N_X_c_417_n 0.00560396f $X=3.34 $Y=0.665 $X2=0 $Y2=0
cc_209 N_A_72_367#_c_268_n N_X_c_417_n 0.00328831f $X=2.715 $Y=1.1 $X2=0 $Y2=0
cc_210 N_A_72_367#_c_254_n X 0.00709794f $X=2.905 $Y=1.615 $X2=0 $Y2=0
cc_211 N_A_72_367#_c_257_n X 0.0162666f $X=3.265 $Y=1.36 $X2=0 $Y2=0
cc_212 N_A_72_367#_M1009_g X 0.0111747f $X=3.34 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A_72_367#_c_268_n X 0.0246569f $X=2.715 $Y=1.1 $X2=0 $Y2=0
cc_214 N_A_72_367#_c_262_n N_VGND_M1002_d 0.00327539f $X=1.76 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A_72_367#_c_264_n N_VGND_M1006_d 2.23166e-19 $X=2.145 $Y=0.825 $X2=0
+ $Y2=0
cc_216 N_A_72_367#_c_266_n N_VGND_M1006_d 0.00171947f $X=2.575 $Y=1.1 $X2=0
+ $Y2=0
cc_217 N_A_72_367#_c_268_n N_VGND_M1006_d 0.0032193f $X=2.715 $Y=1.1 $X2=0 $Y2=0
cc_218 N_A_72_367#_c_263_n N_VGND_c_438_n 0.00567631f $X=1.09 $Y=0.74 $X2=0
+ $Y2=0
cc_219 N_A_72_367#_c_262_n N_VGND_c_439_n 0.0242399f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_72_367#_M1011_g N_VGND_c_441_n 0.00698674f $X=3.34 $Y=0.665 $X2=0
+ $Y2=0
cc_221 N_A_72_367#_c_290_n N_VGND_c_444_n 0.0170002f $X=0.915 $Y=0.42 $X2=0
+ $Y2=0
cc_222 N_A_72_367#_c_262_n N_VGND_c_444_n 0.00228867f $X=1.76 $Y=0.74 $X2=0
+ $Y2=0
cc_223 N_A_72_367#_c_263_n N_VGND_c_444_n 0.00236596f $X=1.09 $Y=0.74 $X2=0
+ $Y2=0
cc_224 N_A_72_367#_c_262_n N_VGND_c_446_n 0.00473472f $X=1.76 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_72_367#_c_297_n N_VGND_c_446_n 0.0151921f $X=1.925 $Y=0.42 $X2=0
+ $Y2=0
cc_226 N_A_72_367#_M1003_g N_VGND_c_447_n 0.00477554f $X=2.91 $Y=0.665 $X2=0
+ $Y2=0
cc_227 N_A_72_367#_M1011_g N_VGND_c_447_n 0.00575161f $X=3.34 $Y=0.665 $X2=0
+ $Y2=0
cc_228 N_A_72_367#_c_254_n N_VGND_c_448_n 9.84837e-19 $X=2.905 $Y=1.615 $X2=0
+ $Y2=0
cc_229 N_A_72_367#_M1003_g N_VGND_c_448_n 0.011673f $X=2.91 $Y=0.665 $X2=0 $Y2=0
cc_230 N_A_72_367#_M1011_g N_VGND_c_448_n 6.29286e-19 $X=3.34 $Y=0.665 $X2=0
+ $Y2=0
cc_231 N_A_72_367#_c_264_n N_VGND_c_448_n 0.017619f $X=2.145 $Y=0.825 $X2=0
+ $Y2=0
cc_232 N_A_72_367#_c_265_n N_VGND_c_448_n 0.00164685f $X=2.145 $Y=1.015 $X2=0
+ $Y2=0
cc_233 N_A_72_367#_c_266_n N_VGND_c_448_n 0.015811f $X=2.575 $Y=1.1 $X2=0 $Y2=0
cc_234 N_A_72_367#_c_268_n N_VGND_c_448_n 0.0182116f $X=2.715 $Y=1.1 $X2=0 $Y2=0
cc_235 N_A_72_367#_M1010_d N_VGND_c_449_n 0.00234862f $X=0.775 $Y=0.245 $X2=0
+ $Y2=0
cc_236 N_A_72_367#_M1000_d N_VGND_c_449_n 0.00241004f $X=1.785 $Y=0.245 $X2=0
+ $Y2=0
cc_237 N_A_72_367#_M1003_g N_VGND_c_449_n 0.00820931f $X=2.91 $Y=0.665 $X2=0
+ $Y2=0
cc_238 N_A_72_367#_M1011_g N_VGND_c_449_n 0.0115045f $X=3.34 $Y=0.665 $X2=0
+ $Y2=0
cc_239 N_A_72_367#_c_290_n N_VGND_c_449_n 0.0109407f $X=0.915 $Y=0.42 $X2=0
+ $Y2=0
cc_240 N_A_72_367#_c_262_n N_VGND_c_449_n 0.013933f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A_72_367#_c_263_n N_VGND_c_449_n 0.00429042f $X=1.09 $Y=0.74 $X2=0
+ $Y2=0
cc_242 N_A_72_367#_c_297_n N_VGND_c_449_n 0.00971501f $X=1.925 $Y=0.42 $X2=0
+ $Y2=0
cc_243 N_A_72_367#_c_264_n N_VGND_c_449_n 4.01127e-19 $X=2.145 $Y=0.825 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_383_n N_X_M1004_d 0.00401517f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_c_386_n X 0.00152603f $X=3.555 $Y=1.98 $X2=0 $Y2=0
cc_246 N_VPWR_c_388_n X 0.0142233f $X=3.43 $Y=3.33 $X2=0 $Y2=0
cc_247 N_VPWR_c_383_n X 0.0090585f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_248 N_X_c_417_n N_VGND_c_441_n 0.0014842f $X=3.125 $Y=0.42 $X2=0 $Y2=0
cc_249 N_X_c_417_n N_VGND_c_447_n 0.0138717f $X=3.125 $Y=0.42 $X2=0 $Y2=0
cc_250 N_X_M1003_s N_VGND_c_449_n 0.00397496f $X=2.985 $Y=0.245 $X2=0 $Y2=0
cc_251 N_X_c_417_n N_VGND_c_449_n 0.00886411f $X=3.125 $Y=0.42 $X2=0 $Y2=0
