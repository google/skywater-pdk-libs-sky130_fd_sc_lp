* File: sky130_fd_sc_lp__a211o_m.spice
* Created: Fri Aug 28 09:48:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a211o_m.pex.spice"
.subckt sky130_fd_sc_lp__a211o_m  VNB VPB A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_82_483#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.18165 AS=0.1113 PD=1.285 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1001 A_322_145# N_A2_M1001_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.18165 PD=0.63 PS=1.285 NRD=14.28 NRS=167.136 M=1 R=2.8 SA=75001.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1009 N_A_82_483#_M1009_d N_A1_M1009_g A_322_145# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_B1_M1000_g N_A_82_483#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_82_483#_M1004_d N_C1_M1004_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0756 PD=1.37 PS=0.78 NRD=0 NRS=0 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_82_483#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A2_M1002_g N_A_225_389#_M1002_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1008 N_A_225_389#_M1008_d N_A1_M1008_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_480_389# N_B1_M1003_g N_A_225_389#_M1008_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_82_483#_M1005_d N_C1_M1005_g A_480_389# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_62 VPB 0 1.41162e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a211o_m.pxi.spice"
*
.ends
*
*
