* File: sky130_fd_sc_lp__ha_2.spice
* Created: Fri Aug 28 10:36:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ha_2.pex.spice"
.subckt sky130_fd_sc_lp__ha_2  VNB VPB B A VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_M1010_g N_A_45_121#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_45_121#_M1009_d N_B_M1009_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1011 N_A_227_397#_M1011_d N_A_270_95#_M1011_g N_A_45_121#_M1009_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_492_131# N_B_M1004_g N_A_270_95#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g A_492_131# VNB NSHORT L=0.15 W=0.42 AD=0.098
+ AS=0.0441 PD=0.85 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1001_d N_A_270_95#_M1005_g N_COUT_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.196 AS=0.1176 PD=1.7 PS=1.12 NRD=11.064 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_A_270_95#_M1015_g N_COUT_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1827 AS=0.1176 PD=1.275 PS=1.12 NRD=12.132 NRS=0 M=1 R=5.6
+ SA=75001.1 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1015_d N_A_227_397#_M1000_g N_SUM_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1827 AS=0.1176 PD=1.275 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6
+ SA=75001.7 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A_227_397#_M1012_g N_SUM_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 A_155_397# N_A_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.1696 PD=0.85 PS=1.81 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75004.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_227_397#_M1006_d N_B_M1006_g A_155_397# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75003.8 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A_270_95#_M1003_g N_A_227_397#_M1006_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2 AS=0.1248 PD=1.265 PS=1.03 NRD=23.0687 NRS=33.8446 M=1
+ R=4.26667 SA=75001.1 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1014 N_A_270_95#_M1014_d N_B_M1014_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.2 PD=0.92 PS=1.265 NRD=0 NRS=83.0946 M=1 R=4.26667 SA=75001.9
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_270_95#_M1014_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.136185 AS=0.0896 PD=1.10147 PS=0.92 NRD=48.5605 NRS=0 M=1 R=4.26667
+ SA=75002.3 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1007_d N_A_270_95#_M1008_g N_COUT_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.268115 AS=0.1764 PD=2.16853 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_A_270_95#_M1016_g N_COUT_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1002 N_SUM_M1002_d N_A_227_397#_M1002_g N_VPWR_M1016_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1017 N_SUM_M1002_d N_A_227_397#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.4284 PD=1.54 PS=3.2 NRD=0 NRS=10.1455 M=1 R=8.4
+ SA=75002.8 SB=75000.3 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=10.5559 P=15.05
c_101 VPB 0 1.74012e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__ha_2.pxi.spice"
*
.ends
*
*
