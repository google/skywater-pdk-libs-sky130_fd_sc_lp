* File: sky130_fd_sc_lp__clkinvlp_4.pex.spice
* Created: Fri Aug 28 10:18:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKINVLP_4%A 3 7 11 15 19 23 27 31 33 34 46
r69 41 42 45.142 $w=3.31e-07 $l=3.1e-07 $layer=POLY_cond $X=0.525 $Y=1.407
+ $X2=0.835 $Y2=1.407
r70 40 41 7.28097 $w=3.31e-07 $l=5e-08 $layer=POLY_cond $X=0.475 $Y=1.407
+ $X2=0.525 $Y2=1.407
r71 38 40 22.571 $w=3.31e-07 $l=1.55e-07 $layer=POLY_cond $X=0.32 $Y=1.407
+ $X2=0.475 $Y2=1.407
r72 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.415 $X2=0.32 $Y2=1.415
r73 34 39 8.1158 $w=3.53e-07 $l=2.5e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.415
r74 33 39 3.89558 $w=3.53e-07 $l=1.2e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.415
r75 29 46 71.3535 $w=3.31e-07 $l=4.9e-07 $layer=POLY_cond $X=2.115 $Y=1.407
+ $X2=1.625 $Y2=1.407
r76 29 31 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=2.115 $Y=1.565
+ $X2=2.115 $Y2=2.48
r77 25 46 21.295 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=1.407
r78 25 27 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=0.61
r79 21 46 5.82477 $w=3.31e-07 $l=4e-08 $layer=POLY_cond $X=1.585 $Y=1.407
+ $X2=1.625 $Y2=1.407
r80 21 44 46.5982 $w=3.31e-07 $l=3.2e-07 $layer=POLY_cond $X=1.585 $Y=1.407
+ $X2=1.265 $Y2=1.407
r81 21 23 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=1.585 $Y=1.565
+ $X2=1.585 $Y2=2.48
r82 17 44 21.295 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=1.265 $Y=1.235
+ $X2=1.265 $Y2=1.407
r83 17 19 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.265 $Y=1.235
+ $X2=1.265 $Y2=0.61
r84 13 44 30.5801 $w=3.31e-07 $l=2.1e-07 $layer=POLY_cond $X=1.055 $Y=1.407
+ $X2=1.265 $Y2=1.407
r85 13 42 32.0363 $w=3.31e-07 $l=2.2e-07 $layer=POLY_cond $X=1.055 $Y=1.407
+ $X2=0.835 $Y2=1.407
r86 13 15 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=1.055 $Y=1.565
+ $X2=1.055 $Y2=2.48
r87 9 42 21.295 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=1.407
r88 9 11 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=0.61
r89 5 41 9.41475 $w=2.5e-07 $l=1.73e-07 $layer=POLY_cond $X=0.525 $Y=1.58
+ $X2=0.525 $Y2=1.407
r90 5 7 223.608 $w=2.5e-07 $l=9e-07 $layer=POLY_cond $X=0.525 $Y=1.58 $X2=0.525
+ $Y2=2.48
r91 1 40 21.295 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=1.407
r92 1 3 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_4%VPWR 1 2 3 10 12 16 20 26 31 32 33 40 41
+ 47
r39 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 38 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 35 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.32 $Y2=3.33
r46 35 37 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 33 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 33 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 31 37 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.38 $Y2=3.33
r51 30 40 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 30 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.38 $Y2=3.33
r53 26 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.38 $Y=2.125
+ $X2=2.38 $Y2=2.835
r54 24 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=3.33
r55 24 29 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=2.835
r56 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.32 $Y=2.125
+ $X2=1.32 $Y2=2.835
r57 18 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=3.245
+ $X2=1.32 $Y2=3.33
r58 18 23 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.32 $Y=3.245
+ $X2=1.32 $Y2=2.835
r59 17 44 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r60 16 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.32 $Y2=3.33
r61 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=0.425 $Y2=3.33
r62 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.26 $Y=2.125
+ $X2=0.26 $Y2=2.835
r63 10 44 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r64 10 15 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.835
r65 3 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.98 $X2=2.38 $Y2=2.835
r66 3 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.98 $X2=2.38 $Y2=2.125
r67 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.98 $X2=1.32 $Y2=2.835
r68 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.98 $X2=1.32 $Y2=2.125
r69 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.98 $X2=0.26 $Y2=2.835
r70 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.98 $X2=0.26 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_4%Y 1 2 3 10 14 22 24 25 26 27 28 29
r41 28 29 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.79 $Y=2.405
+ $X2=0.79 $Y2=2.775
r42 28 47 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.79 $Y=2.405
+ $X2=0.79 $Y2=2.125
r43 27 47 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.79 $Y=2.035 $X2=0.79
+ $Y2=2.125
r44 26 27 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.79 $Y=1.665
+ $X2=0.79 $Y2=2.035
r45 26 41 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.79 $Y=1.665 $X2=0.79
+ $Y2=1.565
r46 25 37 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=1.4 $X2=0.79
+ $Y2=1.235
r47 25 41 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=1.4 $X2=0.79
+ $Y2=1.565
r48 25 37 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=0.79 $Y=1.222
+ $X2=0.79 $Y2=1.235
r49 24 25 10.372 $w=3.28e-07 $l=2.97e-07 $layer=LI1_cond $X=0.79 $Y=0.925
+ $X2=0.79 $Y2=1.222
r50 19 24 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.79 $Y=0.78
+ $X2=0.79 $Y2=0.925
r51 18 22 6.68775 $w=4.63e-07 $l=2.6e-07 $layer=LI1_cond $X=0.79 $Y=0.547
+ $X2=1.05 $Y2=0.547
r52 18 19 2.74626 $w=3.3e-07 $l=2.33e-07 $layer=LI1_cond $X=0.79 $Y=0.547
+ $X2=0.79 $Y2=0.78
r53 14 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.85 $Y=2.125
+ $X2=1.85 $Y2=2.835
r54 12 14 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.85 $Y=1.565
+ $X2=1.85 $Y2=2.125
r55 11 25 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=1.4
+ $X2=0.79 $Y2=1.4
r56 10 12 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=1.685 $Y=1.4
+ $X2=1.85 $Y2=1.565
r57 10 11 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=1.685 $Y=1.4
+ $X2=0.955 $Y2=1.4
r58 3 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.98 $X2=1.85 $Y2=2.835
r59 3 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.98 $X2=1.85 $Y2=2.125
r60 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.98 $X2=0.79 $Y2=2.835
r61 2 47 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.98 $X2=0.79 $Y2=2.125
r62 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.335 $X2=1.05 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_4%VGND 1 2 7 9 13 15 17 24 25 31
r27 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r28 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 25 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r30 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r31 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.84
+ $Y2=0
r32 22 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.64
+ $Y2=0
r33 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r34 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r35 18 28 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r36 18 20 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r37 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.84
+ $Y2=0
r38 17 20 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=0.72
+ $Y2=0
r39 15 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r40 15 21 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r41 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0
r42 11 13 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0.61
r43 7 28 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r44 7 9 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.61
r45 2 13 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.335 $X2=1.84 $Y2=0.61
r46 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.335 $X2=0.26 $Y2=0.61
.ends

