* File: sky130_fd_sc_lp__o41a_4.pex.spice
* Created: Wed Sep  2 10:27:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41A_4%A_83_23# 1 2 3 12 16 20 24 28 32 36 40 42 51
+ 52 54 58 59 60 64 71 81
c128 58 0 6.65354e-20 $X=2.79 $Y=0.95
r129 78 79 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.92 $Y=1.49
+ $X2=1.35 $Y2=1.49
r130 71 73 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.955 $Y=0.735
+ $X2=2.955 $Y2=0.95
r131 68 69 14.2011 $w=1.89e-07 $l=2.2e-07 $layer=LI1_cond $X=2.42 $Y=1.49
+ $X2=2.42 $Y2=1.71
r132 64 66 42.0287 $w=1.88e-07 $l=7.2e-07 $layer=LI1_cond $X=3.815 $Y=1.85
+ $X2=3.815 $Y2=2.57
r133 62 64 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=3.815 $Y=1.815
+ $X2=3.815 $Y2=1.85
r134 61 69 0.0633028 $w=2.1e-07 $l=1e-07 $layer=LI1_cond $X=2.52 $Y=1.71
+ $X2=2.42 $Y2=1.71
r135 60 62 6.83868 $w=2.1e-07 $l=1.44914e-07 $layer=LI1_cond $X=3.72 $Y=1.71
+ $X2=3.815 $Y2=1.815
r136 60 61 63.3766 $w=2.08e-07 $l=1.2e-06 $layer=LI1_cond $X=3.72 $Y=1.71
+ $X2=2.52 $Y2=1.71
r137 58 73 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0.95
+ $X2=2.955 $Y2=0.95
r138 58 59 17.2525 $w=1.78e-07 $l=2.8e-07 $layer=LI1_cond $X=2.79 $Y=0.95
+ $X2=2.51 $Y2=0.95
r139 54 56 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.425 $Y=1.98
+ $X2=2.425 $Y2=2.91
r140 52 69 6.74211 $w=1.9e-07 $l=1.07471e-07 $layer=LI1_cond $X=2.425 $Y=1.815
+ $X2=2.42 $Y2=1.71
r141 52 54 9.63158 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=1.815
+ $X2=2.425 $Y2=1.98
r142 51 68 6.1 $w=1.9e-07 $l=9.74679e-08 $layer=LI1_cond $X=2.415 $Y=1.395
+ $X2=2.42 $Y2=1.49
r143 50 59 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=2.415 $Y=1.04
+ $X2=2.51 $Y2=0.95
r144 50 51 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=2.415 $Y=1.04
+ $X2=2.415 $Y2=1.395
r145 49 81 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.69 $Y=1.49 $X2=1.78
+ $Y2=1.49
r146 49 79 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.69 $Y=1.49
+ $X2=1.35 $Y2=1.49
r147 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.49 $X2=1.69 $Y2=1.49
r148 45 78 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.67 $Y=1.49
+ $X2=0.92 $Y2=1.49
r149 45 75 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.67 $Y=1.49
+ $X2=0.49 $Y2=1.49
r150 44 48 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=0.67 $Y=1.49
+ $X2=1.69 $Y2=1.49
r151 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.67
+ $Y=1.49 $X2=0.67 $Y2=1.49
r152 42 68 0.684278 $w=1.9e-07 $l=1e-07 $layer=LI1_cond $X=2.32 $Y=1.49 $X2=2.42
+ $Y2=1.49
r153 42 48 36.7751 $w=1.88e-07 $l=6.3e-07 $layer=LI1_cond $X=2.32 $Y=1.49
+ $X2=1.69 $Y2=1.49
r154 38 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.655
+ $X2=1.78 $Y2=1.49
r155 38 40 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.78 $Y=1.655
+ $X2=1.78 $Y2=2.465
r156 34 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=1.49
r157 34 36 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.78 $Y=1.325
+ $X2=1.78 $Y2=0.665
r158 30 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.655
+ $X2=1.35 $Y2=1.49
r159 30 32 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.35 $Y=1.655
+ $X2=1.35 $Y2=2.465
r160 26 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=1.49
r161 26 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.35 $Y=1.325
+ $X2=1.35 $Y2=0.665
r162 22 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.655
+ $X2=0.92 $Y2=1.49
r163 22 24 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.92 $Y=1.655
+ $X2=0.92 $Y2=2.465
r164 18 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.325
+ $X2=0.92 $Y2=1.49
r165 18 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.92 $Y=1.325
+ $X2=0.92 $Y2=0.665
r166 14 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.655
+ $X2=0.49 $Y2=1.49
r167 14 16 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.49 $Y=1.655
+ $X2=0.49 $Y2=2.465
r168 10 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=1.49
r169 10 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.49 $Y=1.325
+ $X2=0.49 $Y2=0.665
r170 3 66 400 $w=1.7e-07 $l=9.12318e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.725 $X2=3.815 $Y2=2.57
r171 3 64 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.675
+ $Y=1.725 $X2=3.815 $Y2=1.85
r172 2 56 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.835 $X2=2.425 $Y2=2.91
r173 2 54 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.285
+ $Y=1.835 $X2=2.425 $Y2=1.98
r174 1 71 182 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.235 $X2=2.955 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%B1 3 7 9 11 12 14 15 24
c54 12 0 6.65354e-20 $X=3.17 $Y=1.185
r55 22 24 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=3.17 $Y2=1.35
r56 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.855
+ $Y=1.35 $X2=2.855 $Y2=1.35
r57 20 22 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=2.74 $Y=1.35
+ $X2=2.855 $Y2=1.35
r58 19 20 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.64 $Y=1.35 $X2=2.74
+ $Y2=1.35
r59 17 19 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.21 $Y=1.35
+ $X2=2.64 $Y2=1.35
r60 15 23 13.5732 $w=2.23e-07 $l=2.65e-07 $layer=LI1_cond $X=3.12 $Y=1.322
+ $X2=2.855 $Y2=1.322
r61 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.185
+ $X2=3.17 $Y2=1.35
r62 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.17 $Y=1.185
+ $X2=3.17 $Y2=0.655
r63 9 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.185
+ $X2=2.74 $Y2=1.35
r64 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.74 $Y=1.185
+ $X2=2.74 $Y2=0.655
r65 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=1.515
+ $X2=2.64 $Y2=1.35
r66 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.64 $Y=1.515 $X2=2.64
+ $Y2=2.465
r67 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.515
+ $X2=2.21 $Y2=1.35
r68 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.21 $Y=1.515 $X2=2.21
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%A4 1 3 6 8 10 13 15 22
c46 15 0 1.07548e-19 $X=3.6 $Y=1.295
c47 6 0 1.00671e-19 $X=3.6 $Y=2.355
r48 20 22 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=3.65 $Y=1.35
+ $X2=4.03 $Y2=1.35
r49 17 20 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=3.6 $Y=1.35 $X2=3.65
+ $Y2=1.35
r50 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.65
+ $Y=1.35 $X2=3.65 $Y2=1.35
r51 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.03 $Y=1.515
+ $X2=4.03 $Y2=1.35
r52 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.03 $Y=1.515
+ $X2=4.03 $Y2=2.355
r53 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.03 $Y=1.185
+ $X2=4.03 $Y2=1.35
r54 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.03 $Y=1.185
+ $X2=4.03 $Y2=0.655
r55 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=1.515 $X2=3.6
+ $Y2=1.35
r56 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.6 $Y=1.515 $X2=3.6
+ $Y2=2.355
r57 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=1.185 $X2=3.6
+ $Y2=1.35
r58 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.6 $Y=1.185 $X2=3.6
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%A3 1 3 6 8 10 13 15 16 17 26
c52 26 0 2.86603e-19 $X=4.89 $Y=1.35
c53 13 0 8.70115e-20 $X=4.89 $Y=2.355
r54 24 26 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.87 $Y=1.35 $X2=4.89
+ $Y2=1.35
r55 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.87
+ $Y=1.35 $X2=4.87 $Y2=1.35
r56 21 24 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=4.46 $Y=1.35
+ $X2=4.87 $Y2=1.35
r57 17 25 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=5.04 $Y=1.322
+ $X2=4.87 $Y2=1.322
r58 16 25 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=4.56 $Y=1.322
+ $X2=4.87 $Y2=1.322
r59 15 16 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.322
+ $X2=4.56 $Y2=1.322
r60 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.515
+ $X2=4.89 $Y2=1.35
r61 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.89 $Y=1.515
+ $X2=4.89 $Y2=2.355
r62 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.89 $Y=1.185
+ $X2=4.89 $Y2=1.35
r63 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.89 $Y=1.185
+ $X2=4.89 $Y2=0.655
r64 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.46 $Y=1.515
+ $X2=4.46 $Y2=1.35
r65 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.46 $Y=1.515 $X2=4.46
+ $Y2=2.355
r66 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.46 $Y=1.185
+ $X2=4.46 $Y2=1.35
r67 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.46 $Y=1.185 $X2=4.46
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%A2 1 3 4 5 8 10 12 15 17 18 26
c49 18 0 3.29205e-19 $X=6 $Y=1.295
r50 25 26 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.24 $Y=1.35 $X2=6.31
+ $Y2=1.35
r51 23 25 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=6.06 $Y=1.35 $X2=6.24
+ $Y2=1.35
r52 21 23 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.88 $Y=1.35 $X2=6.06
+ $Y2=1.35
r53 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.06
+ $Y=1.35 $X2=6.06 $Y2=1.35
r54 17 18 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.322 $X2=6
+ $Y2=1.322
r55 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.31 $Y=1.515
+ $X2=6.31 $Y2=1.35
r56 13 15 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.31 $Y=1.515
+ $X2=6.31 $Y2=2.465
r57 10 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.24 $Y=1.185
+ $X2=6.24 $Y2=1.35
r58 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.24 $Y=1.185
+ $X2=6.24 $Y2=0.655
r59 6 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.88 $Y=1.515
+ $X2=5.88 $Y2=1.35
r60 6 8 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.88 $Y=1.515 $X2=5.88
+ $Y2=2.465
r61 4 21 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.805 $Y=1.35
+ $X2=5.88 $Y2=1.35
r62 4 5 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=5.805 $Y=1.35
+ $X2=5.395 $Y2=1.35
r63 1 5 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.32 $Y=1.185
+ $X2=5.395 $Y2=1.35
r64 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.32 $Y=1.185 $X2=5.32
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%A1 1 3 6 8 10 13 15 16 17 24
c37 24 0 1.5015e-19 $X=7.1 $Y=1.35
r38 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.1 $Y=1.35
+ $X2=7.1 $Y2=1.35
r39 22 24 52.1081 $w=3.33e-07 $l=3.6e-07 $layer=POLY_cond $X=6.74 $Y=1.355
+ $X2=7.1 $Y2=1.355
r40 21 22 10.1321 $w=3.33e-07 $l=7e-08 $layer=POLY_cond $X=6.67 $Y=1.355
+ $X2=6.74 $Y2=1.355
r41 17 25 17.4147 $w=2.23e-07 $l=3.4e-07 $layer=LI1_cond $X=7.44 $Y=1.322
+ $X2=7.1 $Y2=1.322
r42 16 25 7.17076 $w=2.23e-07 $l=1.4e-07 $layer=LI1_cond $X=6.96 $Y=1.322
+ $X2=7.1 $Y2=1.322
r43 15 16 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.322
+ $X2=6.96 $Y2=1.322
r44 11 24 10.1321 $w=3.33e-07 $l=7e-08 $layer=POLY_cond $X=7.17 $Y=1.355 $X2=7.1
+ $Y2=1.355
r45 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.17 $Y=1.515
+ $X2=7.17 $Y2=2.465
r46 8 24 21.4384 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.1 $Y=1.185 $X2=7.1
+ $Y2=1.355
r47 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.1 $Y=1.185 $X2=7.1
+ $Y2=0.655
r48 4 22 21.4384 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.74 $Y=1.525
+ $X2=6.74 $Y2=1.355
r49 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=6.74 $Y=1.525 $X2=6.74
+ $Y2=2.465
r50 1 21 21.4384 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.67 $Y=1.185
+ $X2=6.67 $Y2=1.355
r51 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.67 $Y=1.185 $X2=6.67
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%VPWR 1 2 3 4 5 16 18 24 30 36 42 47 48 50 51
+ 52 54 66 75 76 82 85
r102 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r103 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r104 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 76 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r106 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r107 73 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.12 $Y=3.33
+ $X2=6.955 $Y2=3.33
r108 73 75 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.12 $Y=3.33
+ $X2=7.44 $Y2=3.33
r109 72 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r110 71 72 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r111 68 71 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 68 69 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r113 66 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.79 $Y=3.33
+ $X2=6.955 $Y2=3.33
r114 66 71 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.79 $Y=3.33
+ $X2=6.48 $Y2=3.33
r115 65 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r116 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 62 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 59 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.135 $Y2=3.33
r121 59 61 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.68 $Y2=3.33
r122 58 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 58 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r124 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 55 79 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r126 55 57 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 54 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.135 $Y2=3.33
r128 54 57 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 52 72 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=6.48 $Y2=3.33
r130 52 69 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.12 $Y2=3.33
r131 50 64 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=3.33 $X2=2.64
+ $Y2=3.33
r132 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=2.855 $Y2=3.33
r133 49 68 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.02 $Y=3.33 $X2=3.12
+ $Y2=3.33
r134 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=2.855 $Y2=3.33
r135 47 61 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=1.68 $Y2=3.33
r136 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=1.995 $Y2=3.33
r137 46 64 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=1.995 $Y2=3.33
r139 42 45 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=6.955 $Y=2.19
+ $X2=6.955 $Y2=2.95
r140 40 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.955 $Y=3.245
+ $X2=6.955 $Y2=3.33
r141 40 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.955 $Y=3.245
+ $X2=6.955 $Y2=2.95
r142 36 39 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=2.855 $Y=2.07
+ $X2=2.855 $Y2=2.95
r143 34 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=3.245
+ $X2=2.855 $Y2=3.33
r144 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.855 $Y=3.245
+ $X2=2.855 $Y2=2.95
r145 30 33 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=1.995 $Y=1.98
+ $X2=1.995 $Y2=2.95
r146 28 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=3.245
+ $X2=1.995 $Y2=3.33
r147 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.995 $Y=3.245
+ $X2=1.995 $Y2=2.95
r148 24 27 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.135 $Y=2.19
+ $X2=1.135 $Y2=2.95
r149 22 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=3.33
r150 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=2.95
r151 18 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.275 $Y=2.18
+ $X2=0.275 $Y2=2.95
r152 16 79 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r153 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.95
r154 5 45 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.815
+ $Y=1.835 $X2=6.955 $Y2=2.95
r155 5 42 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=6.815
+ $Y=1.835 $X2=6.955 $Y2=2.19
r156 4 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=1.835 $X2=2.855 $Y2=2.95
r157 4 36 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=1.835 $X2=2.855 $Y2=2.07
r158 3 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=1.995 $Y2=2.95
r159 3 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=1.995 $Y2=1.98
r160 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.95
r161 2 24 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.835 $X2=1.135 $Y2=2.19
r162 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.95
r163 1 18 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%X 1 2 3 4 13 15 16 19 23 27 29 33 37 42 43 44
+ 45 49 51
r58 49 51 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=0.21 $Y=1.225 $X2=0.21
+ $Y2=1.295
r59 44 49 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.21 $Y=1.14 $X2=0.21
+ $Y2=1.225
r60 44 45 16.7335 $w=2.48e-07 $l=3.63e-07 $layer=LI1_cond $X=0.21 $Y=1.302
+ $X2=0.21 $Y2=1.665
r61 44 51 0.322684 $w=2.48e-07 $l=7e-09 $layer=LI1_cond $X=0.21 $Y=1.302
+ $X2=0.21 $Y2=1.295
r62 41 45 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.21 $Y=1.755 $X2=0.21
+ $Y2=1.665
r63 37 39 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.565 $Y=1.98
+ $X2=1.565 $Y2=2.91
r64 35 37 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.565 $Y=1.925
+ $X2=1.565 $Y2=1.98
r65 31 33 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=1.565 $Y=1.055
+ $X2=1.565 $Y2=0.42
r66 30 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.8 $Y=1.84 $X2=0.705
+ $Y2=1.84
r67 29 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.47 $Y=1.84
+ $X2=1.565 $Y2=1.925
r68 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.47 $Y=1.84 $X2=0.8
+ $Y2=1.84
r69 28 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.8 $Y=1.14 $X2=0.705
+ $Y2=1.14
r70 27 31 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.47 $Y=1.14
+ $X2=1.565 $Y2=1.055
r71 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.47 $Y=1.14 $X2=0.8
+ $Y2=1.14
r72 23 25 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.705 $Y=1.98
+ $X2=0.705 $Y2=2.91
r73 21 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.925
+ $X2=0.705 $Y2=1.84
r74 21 23 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=0.705 $Y=1.925
+ $X2=0.705 $Y2=1.98
r75 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.055
+ $X2=0.705 $Y2=1.14
r76 17 19 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=0.705 $Y=1.055
+ $X2=0.705 $Y2=0.42
r77 16 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.335 $Y=1.84
+ $X2=0.21 $Y2=1.755
r78 15 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.61 $Y=1.84
+ $X2=0.705 $Y2=1.84
r79 15 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.61 $Y=1.84
+ $X2=0.335 $Y2=1.84
r80 14 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.335 $Y=1.14
+ $X2=0.21 $Y2=1.14
r81 13 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.61 $Y=1.14
+ $X2=0.705 $Y2=1.14
r82 13 14 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.61 $Y=1.14
+ $X2=0.335 $Y2=1.14
r83 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=2.91
r84 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.425
+ $Y=1.835 $X2=1.565 $Y2=1.98
r85 3 25 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.91
r86 3 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=1.98
r87 2 33 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.425
+ $Y=0.245 $X2=1.565 $Y2=0.42
r88 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.245 $X2=0.705 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%A_652_345# 1 2 3 12 16 17 21 24 25 28
c50 25 0 1.00671e-19 $X=4.41 $Y=1.69
c51 16 0 8.70115e-20 $X=4.08 $Y=2.99
r52 28 30 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=5.105 $Y=1.87
+ $X2=5.105 $Y2=2.64
r53 26 28 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.105 $Y=1.775
+ $X2=5.105 $Y2=1.87
r54 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.94 $Y=1.69
+ $X2=5.105 $Y2=1.775
r55 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.94 $Y=1.69
+ $X2=4.41 $Y2=1.69
r56 21 23 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=4.245 $Y=1.87
+ $X2=4.245 $Y2=2.84
r57 19 23 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=4.245 $Y=2.905
+ $X2=4.245 $Y2=2.84
r58 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.245 $Y=1.775
+ $X2=4.41 $Y2=1.69
r59 18 21 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.245 $Y=1.775
+ $X2=4.245 $Y2=1.87
r60 16 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.08 $Y=2.99
+ $X2=4.245 $Y2=2.905
r61 16 17 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.08 $Y=2.99
+ $X2=3.55 $Y2=2.99
r62 12 15 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.385 $Y=2.07
+ $X2=3.385 $Y2=2.84
r63 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.385 $Y=2.905
+ $X2=3.55 $Y2=2.99
r64 10 15 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=3.385 $Y=2.905
+ $X2=3.385 $Y2=2.84
r65 3 30 400 $w=1.7e-07 $l=9.8251e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.725 $X2=5.105 $Y2=2.64
r66 3 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=1.725 $X2=5.105 $Y2=1.87
r67 2 23 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.725 $X2=4.245 $Y2=2.84
r68 2 21 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=1.725 $X2=4.245 $Y2=1.87
r69 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.725 $X2=3.385 $Y2=2.84
r70 1 12 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.725 $X2=3.385 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%A_907_345# 1 2 9 13 14 15 17
r25 15 20 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.095 $Y=2.895
+ $X2=6.095 $Y2=2.985
r26 15 17 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=6.095 $Y=2.895
+ $X2=6.095 $Y2=2.14
r27 13 20 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.93 $Y=2.985
+ $X2=6.095 $Y2=2.985
r28 13 14 71.4747 $w=1.78e-07 $l=1.16e-06 $layer=LI1_cond $X=5.93 $Y=2.985
+ $X2=4.77 $Y2=2.985
r29 9 12 42.6124 $w=1.88e-07 $l=7.3e-07 $layer=LI1_cond $X=4.675 $Y=2.11
+ $X2=4.675 $Y2=2.84
r30 7 14 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=4.675 $Y=2.895
+ $X2=4.77 $Y2=2.985
r31 7 12 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=4.675 $Y=2.895
+ $X2=4.675 $Y2=2.84
r32 2 20 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=5.955
+ $Y=1.835 $X2=6.095 $Y2=2.9
r33 2 17 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=5.955
+ $Y=1.835 $X2=6.095 $Y2=2.14
r34 1 12 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.535
+ $Y=1.725 $X2=4.675 $Y2=2.84
r35 1 9 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=4.535
+ $Y=1.725 $X2=4.675 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%A_1108_367# 1 2 3 12 14 15 18 22 26 30
r39 26 28 51.5727 $w=1.98e-07 $l=9.3e-07 $layer=LI1_cond $X=7.39 $Y=1.98
+ $X2=7.39 $Y2=2.91
r40 24 26 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=7.39 $Y=1.875
+ $X2=7.39 $Y2=1.98
r41 23 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.62 $Y=1.79
+ $X2=6.525 $Y2=1.79
r42 22 24 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=7.29 $Y=1.79
+ $X2=7.39 $Y2=1.875
r43 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.29 $Y=1.79
+ $X2=6.62 $Y2=1.79
r44 18 20 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=6.525 $Y=1.96
+ $X2=6.525 $Y2=2.91
r45 16 30 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.525 $Y=1.875
+ $X2=6.525 $Y2=1.79
r46 16 18 4.96172 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=6.525 $Y=1.875
+ $X2=6.525 $Y2=1.96
r47 14 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.43 $Y=1.79
+ $X2=6.525 $Y2=1.79
r48 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.43 $Y=1.79
+ $X2=5.76 $Y2=1.79
r49 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.63 $Y=1.875
+ $X2=5.76 $Y2=1.79
r50 10 12 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=5.63 $Y=1.875
+ $X2=5.63 $Y2=1.98
r51 3 28 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.835 $X2=7.385 $Y2=2.91
r52 3 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.835 $X2=7.385 $Y2=1.98
r53 2 20 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.385
+ $Y=1.835 $X2=6.525 $Y2=2.91
r54 2 18 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=6.385
+ $Y=1.835 $X2=6.525 $Y2=1.96
r55 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.54
+ $Y=1.835 $X2=5.665 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 38 42 46 49
+ 50 51 52 54 55 56 58 83 84 90 93 98 104
r114 103 104 10.732 $w=7.83e-07 $l=1.25e-07 $layer=LI1_cond $X=6.025 $Y=0.307
+ $X2=6.15 $Y2=0.307
r115 100 103 0.380917 $w=7.83e-07 $l=2.5e-08 $layer=LI1_cond $X=6 $Y=0.307
+ $X2=6.025 $Y2=0.307
r116 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r117 97 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r118 96 100 7.3136 $w=7.83e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=0.307 $X2=6
+ $Y2=0.307
r119 96 98 10.5797 $w=7.83e-07 $l=1.15e-07 $layer=LI1_cond $X=5.52 $Y=0.307
+ $X2=5.405 $Y2=0.307
r120 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r121 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r122 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r123 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r124 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r125 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r126 81 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r127 80 104 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=6.15
+ $Y2=0
r128 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r129 77 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r130 77 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r131 76 98 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.04 $Y=0
+ $X2=5.405 $Y2=0
r132 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r133 74 93 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=4.672
+ $Y2=0
r134 74 76 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r135 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r136 69 72 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r137 68 71 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r138 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r139 66 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r140 66 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r141 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r142 63 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.135
+ $Y2=0
r143 63 65 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.68
+ $Y2=0
r144 62 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r145 62 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r146 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r147 59 87 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r148 59 61 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.72
+ $Y2=0
r149 58 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.135
+ $Y2=0
r150 58 61 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.72
+ $Y2=0
r151 56 94 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=4.56
+ $Y2=0
r152 56 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r153 54 80 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.48 $Y2=0
r154 54 55 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.885
+ $Y2=0
r155 53 83 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.015 $Y=0
+ $X2=7.44 $Y2=0
r156 53 55 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.015 $Y=0 $X2=6.885
+ $Y2=0
r157 51 71 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.6
+ $Y2=0
r158 51 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.815
+ $Y2=0
r159 49 65 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.68
+ $Y2=0
r160 49 50 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.99
+ $Y2=0
r161 48 68 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.16
+ $Y2=0
r162 48 50 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=1.99
+ $Y2=0
r163 44 55 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.885 $Y=0.085
+ $X2=6.885 $Y2=0
r164 44 46 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=6.885 $Y=0.085
+ $X2=6.885 $Y2=0.535
r165 40 93 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.672 $Y=0.085
+ $X2=4.672 $Y2=0
r166 40 42 20.3372 $w=2.53e-07 $l=4.5e-07 $layer=LI1_cond $X=4.672 $Y=0.085
+ $X2=4.672 $Y2=0.535
r167 39 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.945 $Y=0 $X2=3.815
+ $Y2=0
r168 38 93 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.545 $Y=0
+ $X2=4.672 $Y2=0
r169 38 39 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.545 $Y=0 $X2=3.945
+ $Y2=0
r170 34 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0
r171 34 36 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0.535
r172 30 50 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0
r173 30 32 10.9842 $w=3.18e-07 $l=3.05e-07 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0.39
r174 26 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0
r175 26 28 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0.37
r176 22 87 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r177 22 24 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.39
r178 7 46 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=6.745
+ $Y=0.235 $X2=6.885 $Y2=0.535
r179 6 103 91 $w=1.7e-07 $l=7.65441e-07 $layer=licon1_NDIFF $count=2 $X=5.395
+ $Y=0.235 $X2=6.025 $Y2=0.535
r180 5 42 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=4.535
+ $Y=0.235 $X2=4.675 $Y2=0.535
r181 4 36 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=3.675
+ $Y=0.235 $X2=3.815 $Y2=0.535
r182 3 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.855
+ $Y=0.245 $X2=1.995 $Y2=0.39
r183 2 28 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.995
+ $Y=0.245 $X2=1.135 $Y2=0.37
r184 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.245 $X2=0.275 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_4%A_480_47# 1 2 3 4 5 6 19 25 26 29 31 35 37 41
+ 43 47 49 54 55 56
r72 49 52 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=2.49 $Y=0.34
+ $X2=2.49 $Y2=0.525
r73 45 47 16.0976 $w=3.13e-07 $l=4.4e-07 $layer=LI1_cond $X=7.342 $Y=0.87
+ $X2=7.342 $Y2=0.43
r74 44 56 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=6.585 $Y=0.955
+ $X2=6.452 $Y2=0.955
r75 43 45 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=7.185 $Y=0.955
+ $X2=7.342 $Y2=0.87
r76 43 44 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.185 $Y=0.955
+ $X2=6.585 $Y2=0.955
r77 39 56 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=6.452 $Y=0.87
+ $X2=6.452 $Y2=0.955
r78 39 41 19.5698 $w=2.63e-07 $l=4.5e-07 $layer=LI1_cond $X=6.452 $Y=0.87
+ $X2=6.452 $Y2=0.42
r79 38 55 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.235 $Y=0.955
+ $X2=5.102 $Y2=0.955
r80 37 56 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=6.32 $Y=0.955
+ $X2=6.452 $Y2=0.955
r81 37 38 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=6.32 $Y=0.955
+ $X2=5.235 $Y2=0.955
r82 33 55 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.102 $Y=0.87
+ $X2=5.102 $Y2=0.955
r83 33 35 19.5698 $w=2.63e-07 $l=4.5e-07 $layer=LI1_cond $X=5.102 $Y=0.87
+ $X2=5.102 $Y2=0.42
r84 32 54 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.375 $Y=0.955
+ $X2=4.245 $Y2=0.955
r85 31 55 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.97 $Y=0.955
+ $X2=5.102 $Y2=0.955
r86 31 32 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.97 $Y=0.955
+ $X2=4.375 $Y2=0.955
r87 27 54 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.245 $Y=0.87
+ $X2=4.245 $Y2=0.955
r88 27 29 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=4.245 $Y=0.87
+ $X2=4.245 $Y2=0.42
r89 25 54 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.115 $Y=0.955
+ $X2=4.245 $Y2=0.955
r90 25 26 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.115 $Y=0.955
+ $X2=3.515 $Y2=0.955
r91 22 26 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=3.402 $Y=0.87
+ $X2=3.515 $Y2=0.955
r92 22 24 22.5367 $w=2.23e-07 $l=4.4e-07 $layer=LI1_cond $X=3.402 $Y=0.87
+ $X2=3.402 $Y2=0.43
r93 21 24 0.256098 $w=2.23e-07 $l=5e-09 $layer=LI1_cond $X=3.402 $Y=0.425
+ $X2=3.402 $Y2=0.43
r94 20 49 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.62 $Y=0.34 $X2=2.49
+ $Y2=0.34
r95 19 21 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.29 $Y=0.34
+ $X2=3.402 $Y2=0.425
r96 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.29 $Y=0.34
+ $X2=2.62 $Y2=0.34
r97 6 47 91 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=2 $X=7.175
+ $Y=0.235 $X2=7.335 $Y2=0.43
r98 5 41 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.315
+ $Y=0.235 $X2=6.455 $Y2=0.42
r99 4 35 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.965
+ $Y=0.235 $X2=5.105 $Y2=0.42
r100 3 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.105
+ $Y=0.235 $X2=4.245 $Y2=0.42
r101 2 24 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=3.245
+ $Y=0.235 $X2=3.385 $Y2=0.43
r102 1 52 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.235 $X2=2.525 $Y2=0.525
.ends

