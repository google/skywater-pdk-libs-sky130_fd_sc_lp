* File: sky130_fd_sc_lp__a311o_m.spice
* Created: Wed Sep  2 09:25:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311o_m.pex.spice"
.subckt sky130_fd_sc_lp__a311o_m  VNB VPB A3 A2 A1 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_54_154#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1006 A_220_48# N_A3_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0672 PD=0.63 PS=0.74 NRD=14.28 NRS=11.424 M=1 R=2.8 SA=75000.7 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1008 A_292_48# N_A2_M1008_g A_220_48# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_54_154#_M1009_d N_A1_M1009_g A_292_48# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_B1_M1000_g N_A_54_154#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0588 PD=0.81 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_54_154#_M1005_d N_C1_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=25.704 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_54_154#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1011 N_A_196_403#_M1011_d N_A3_M1011_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_196_403#_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.100375 AS=0.0588 PD=0.915 PS=0.7 NRD=39.8531 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_196_403#_M1010_d N_A1_M1010_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.100375 PD=0.7 PS=0.915 NRD=0 NRS=39.8531 M=1 R=2.8
+ SA=75001.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1004 A_486_403# N_B1_M1004_g N_A_196_403#_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_54_154#_M1007_d N_C1_M1007_g A_486_403# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_42 VNB 0 6.36774e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__a311o_m.pxi.spice"
*
.ends
*
*
