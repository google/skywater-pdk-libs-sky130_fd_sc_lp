* File: sky130_fd_sc_lp__dfstp_1.pex.spice
* Created: Fri Aug 28 10:23:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFSTP_1%CLK 2 3 5 6 8 11 13 14 22
c45 22 0 1.29179e-19 $X=0.545 $Y=1.075
r46 20 22 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.525 $Y=1.075
+ $X2=0.545 $Y2=1.075
r47 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.075 $X2=0.525 $Y2=1.075
r48 17 20 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=0.22 $Y=1.075
+ $X2=0.525 $Y2=1.075
r49 14 21 5.82845 $w=4.33e-07 $l=2.2e-07 $layer=LI1_cond $X=0.657 $Y=1.295
+ $X2=0.657 $Y2=1.075
r50 13 21 3.97394 $w=4.33e-07 $l=1.5e-07 $layer=LI1_cond $X=0.657 $Y=0.925
+ $X2=0.657 $Y2=1.075
r51 9 11 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.22 $Y=2.125
+ $X2=0.505 $Y2=2.125
r52 6 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=0.91
+ $X2=0.545 $Y2=1.075
r53 6 8 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.545 $Y=0.91 $X2=0.545
+ $Y2=0.58
r54 3 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.505 $Y=2.2
+ $X2=0.505 $Y2=2.125
r55 3 5 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.505 $Y=2.2 $X2=0.505
+ $Y2=2.635
r56 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.22 $Y=2.05 $X2=0.22
+ $Y2=2.125
r57 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.22 $Y=1.24
+ $X2=0.22 $Y2=1.075
r58 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.22 $Y=1.24 $X2=0.22
+ $Y2=2.05
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%D 1 3 4 6 10 15 17 20
c48 20 0 1.01515e-19 $X=1.6 $Y=1.99
r49 17 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.99 $X2=1.6 $Y2=1.99
r50 13 20 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=1.6 $Y=2.055 $X2=1.6
+ $Y2=1.99
r51 13 15 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.6 $Y=2.13
+ $X2=1.975 $Y2=2.13
r52 8 20 125.026 $w=3.3e-07 $l=7.15e-07 $layer=POLY_cond $X=1.6 $Y=1.275 $X2=1.6
+ $Y2=1.99
r53 8 10 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.6 $Y=1.2 $X2=1.925
+ $Y2=1.2
r54 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.975 $Y=2.205
+ $X2=1.975 $Y2=2.13
r55 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.975 $Y=2.205
+ $X2=1.975 $Y2=2.525
r56 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=1.125
+ $X2=1.925 $Y2=1.2
r57 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.925 $Y=1.125
+ $X2=1.925 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_202_463# 1 2 9 11 15 19 23 25 26 27 28 31
+ 33 36 37 43 44 50 51 60
c170 51 0 1.47832e-19 $X=5.52 $Y=1.295
c171 50 0 9.3441e-20 $X=5.52 $Y=1.295
c172 27 0 4.26559e-20 $X=5.725 $Y=1.51
r173 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.54
+ $Y=1.51 $X2=5.54 $Y2=1.51
r174 51 57 8.65677 $w=3.03e-07 $l=2.15e-07 $layer=LI1_cond $X=5.54 $Y=1.295
+ $X2=5.54 $Y2=1.51
r175 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r176 47 60 26.7664 $w=3.08e-07 $l=7.2e-07 $layer=LI1_cond $X=1.2 $Y=1.295
+ $X2=1.2 $Y2=0.575
r177 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.295
+ $X2=1.2 $Y2=1.295
r178 44 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.295
+ $X2=1.2 $Y2=1.295
r179 43 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=5.52 $Y2=1.295
r180 43 44 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=1.345 $Y2=1.295
r181 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.68 $X2=2.14 $Y2=1.68
r182 37 40 4.0085 $w=2.28e-07 $l=8e-08 $layer=LI1_cond $X=2.12 $Y=1.6 $X2=2.12
+ $Y2=1.68
r183 35 47 8.17863 $w=3.08e-07 $l=2.2e-07 $layer=LI1_cond $X=1.2 $Y=1.515
+ $X2=1.2 $Y2=1.295
r184 35 36 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.515 $X2=1.2
+ $Y2=1.6
r185 34 36 2.90867 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.355 $Y=1.6
+ $X2=1.2 $Y2=1.6
r186 33 37 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.005 $Y=1.6
+ $X2=2.12 $Y2=1.6
r187 33 34 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.005 $Y=1.6
+ $X2=1.355 $Y2=1.6
r188 29 36 3.58051 $w=2.6e-07 $l=1.07121e-07 $layer=LI1_cond $X=1.15 $Y=1.685
+ $X2=1.2 $Y2=1.6
r189 29 31 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=1.15 $Y=1.685
+ $X2=1.15 $Y2=2.46
r190 27 56 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=5.725 $Y=1.51
+ $X2=5.54 $Y2=1.51
r191 27 28 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.725 $Y=1.51
+ $X2=5.725 $Y2=1.345
r192 25 41 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.33 $Y=1.68
+ $X2=2.14 $Y2=1.68
r193 25 26 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=2.33 $Y=1.68
+ $X2=2.405 $Y2=1.68
r194 21 28 37.0704 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=5.835 $Y=1.345
+ $X2=5.725 $Y2=1.345
r195 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.835 $Y=1.345
+ $X2=5.835 $Y2=0.555
r196 17 28 37.0704 $w=1.5e-07 $l=3.65582e-07 $layer=POLY_cond $X=5.8 $Y=1.675
+ $X2=5.725 $Y2=1.345
r197 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.8 $Y=1.675
+ $X2=5.8 $Y2=2.295
r198 13 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.785 $Y=1.515
+ $X2=2.785 $Y2=0.805
r199 12 26 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.48 $Y=1.59
+ $X2=2.405 $Y2=1.68
r200 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.71 $Y=1.59
+ $X2=2.785 $Y2=1.515
r201 11 12 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.71 $Y=1.59
+ $X2=2.48 $Y2=1.59
r202 7 26 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.845
+ $X2=2.405 $Y2=1.68
r203 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.405 $Y=1.845
+ $X2=2.405 $Y2=2.525
r204 2 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=2.315 $X2=1.15 $Y2=2.46
r205 1 60 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.37 $X2=1.19 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_614_93# 1 2 9 14 16 19 21 24 27 29 33 38
+ 41 44
r86 42 44 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.195 $Y=1.455
+ $X2=3.195 $Y2=1.825
r87 35 38 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.835 $Y=2.525
+ $X2=3.95 $Y2=2.525
r88 33 42 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.252 $Y=1.29
+ $X2=3.252 $Y2=1.455
r89 33 41 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.252 $Y=1.29
+ $X2=3.252 $Y2=1.125
r90 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.29 $X2=3.27 $Y2=1.29
r91 29 32 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.27 $Y=1.02
+ $X2=3.27 $Y2=1.29
r92 25 27 20.9147 $w=2.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.945 $Y=0.935
+ $X2=3.945 $Y2=0.445
r93 24 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.835 $Y=2.36
+ $X2=3.835 $Y2=2.525
r94 23 24 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.835 $Y=2.155
+ $X2=3.835 $Y2=2.36
r95 22 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=1.02
+ $X2=3.27 $Y2=1.02
r96 21 25 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.81 $Y=1.02
+ $X2=3.945 $Y2=0.935
r97 21 22 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.81 $Y=1.02
+ $X2=3.435 $Y2=1.02
r98 19 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.99
+ $X2=3.285 $Y2=2.155
r99 19 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.99
+ $X2=3.285 $Y2=1.825
r100 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.285
+ $Y=1.99 $X2=3.285 $Y2=1.99
r101 16 23 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.75 $Y=2.025
+ $X2=3.835 $Y2=2.155
r102 16 18 20.611 $w=2.58e-07 $l=4.65e-07 $layer=LI1_cond $X=3.75 $Y=2.025
+ $X2=3.285 $Y2=2.025
r103 14 45 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.195 $Y=2.525
+ $X2=3.195 $Y2=2.155
r104 9 41 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.145 $Y=0.805
+ $X2=3.145 $Y2=1.125
r105 2 38 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=2.315 $X2=3.95 $Y2=2.525
r106 1 27 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.85
+ $Y=0.235 $X2=3.975 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%SET_B 3 7 10 14 17 18 20 21 24 27 29 30 31
+ 32 42 46 59 61 62
c129 32 0 2.99331e-19 $X=7.44 $Y=1.665
c130 10 0 1.61779e-19 $X=7.08 $Y=0.665
r131 61 62 0.953396 $w=6.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6 $Y=1.59
+ $X2=6.055 $Y2=1.59
r132 46 48 36.572 $w=5.14e-07 $l=3.9e-07 $layer=POLY_cond $X=7.44 $Y=1.58
+ $X2=7.83 $Y2=1.58
r133 32 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.44
+ $Y=1.41 $X2=7.44 $Y2=1.41
r134 31 32 8.56892 $w=6.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.58
+ $X2=7.44 $Y2=1.58
r135 30 31 8.56892 $w=6.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.58
+ $X2=6.96 $Y2=1.58
r136 29 61 0.260017 $w=6.88e-07 $l=1.5e-08 $layer=LI1_cond $X=5.985 $Y=1.59
+ $X2=6 $Y2=1.59
r137 29 59 9.6141 $w=6.88e-07 $l=1e-07 $layer=LI1_cond $X=5.985 $Y=1.59
+ $X2=5.885 $Y2=1.59
r138 29 30 7.31929 $w=6.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.07 $Y=1.58
+ $X2=6.48 $Y2=1.58
r139 29 62 0.267779 $w=6.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.07 $Y=1.58
+ $X2=6.055 $Y2=1.58
r140 27 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.185 $Y=1.99
+ $X2=4.185 $Y2=2.155
r141 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.185
+ $Y=1.99 $X2=4.185 $Y2=1.99
r142 24 59 94.2727 $w=1.68e-07 $l=1.445e-06 $layer=LI1_cond $X=4.44 $Y=1.85
+ $X2=5.885 $Y2=1.85
r143 21 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.64 $Y=0.93
+ $X2=4.64 $Y2=0.765
r144 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.64
+ $Y=0.93 $X2=4.64 $Y2=0.93
r145 18 20 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=4.44 $Y=0.97 $X2=4.64
+ $Y2=0.97
r146 17 24 5.7456 $w=3.02e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.355 $Y=1.765
+ $X2=4.44 $Y2=1.85
r147 17 26 6.86755 $w=3.02e-07 $l=2.66786e-07 $layer=LI1_cond $X=4.355 $Y=1.765
+ $X2=4.185 $Y2=1.96
r148 16 18 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.355 $Y=1.095
+ $X2=4.44 $Y2=0.97
r149 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=1.095
+ $X2=4.355 $Y2=1.765
r150 12 48 32.1071 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.83 $Y=1.915
+ $X2=7.83 $Y2=1.58
r151 12 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.83 $Y=1.915
+ $X2=7.83 $Y2=2.525
r152 8 46 33.7588 $w=5.14e-07 $l=5.002e-07 $layer=POLY_cond $X=7.08 $Y=1.245
+ $X2=7.44 $Y2=1.58
r153 8 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.08 $Y=1.245
+ $X2=7.08 $Y2=0.665
r154 7 42 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.55 $Y=0.445
+ $X2=4.55 $Y2=0.765
r155 3 40 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.165 $Y=2.525
+ $X2=4.165 $Y2=2.155
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_486_119# 1 2 9 13 15 16 19 22 23 24 25 27
+ 29 31 36 38 39 44 46 48
c149 29 0 9.3441e-20 $X=5.09 $Y=1.41
r150 49 55 65.1593 $w=2.7e-07 $l=3.65e-07 $layer=POLY_cond $X=3.825 $Y=1.45
+ $X2=4.19 $Y2=1.45
r151 49 53 16.0667 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=3.825 $Y=1.45
+ $X2=3.735 $Y2=1.45
r152 48 51 8.4217 $w=2.58e-07 $l=1.9e-07 $layer=LI1_cond $X=3.79 $Y=1.45
+ $X2=3.79 $Y2=1.64
r153 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.45 $X2=3.825 $Y2=1.45
r154 42 44 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.62 $Y=2.52
+ $X2=2.84 $Y2=2.52
r155 40 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=1.64
+ $X2=2.84 $Y2=1.64
r156 39 51 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.66 $Y=1.64
+ $X2=3.79 $Y2=1.64
r157 39 40 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.66 $Y=1.64
+ $X2=2.925 $Y2=1.64
r158 38 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=2.355
+ $X2=2.84 $Y2=2.52
r159 37 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=1.725
+ $X2=2.84 $Y2=1.64
r160 37 38 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.84 $Y=1.725
+ $X2=2.84 $Y2=2.355
r161 36 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=1.555
+ $X2=2.84 $Y2=1.64
r162 35 36 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.84 $Y=0.975
+ $X2=2.84 $Y2=1.555
r163 31 35 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.755 $Y=0.81
+ $X2=2.84 $Y2=0.975
r164 31 33 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.755 $Y=0.81
+ $X2=2.57 $Y2=0.81
r165 28 29 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.85 $Y=1.41
+ $X2=5.09 $Y2=1.41
r166 25 27 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.475 $Y=0.985
+ $X2=5.475 $Y2=0.555
r167 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.4 $Y=1.06
+ $X2=5.475 $Y2=0.985
r168 23 24 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.4 $Y=1.06
+ $X2=5.165 $Y2=1.06
r169 22 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.09 $Y=1.335
+ $X2=5.09 $Y2=1.41
r170 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.09 $Y=1.135
+ $X2=5.165 $Y2=1.06
r171 21 22 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.09 $Y=1.135
+ $X2=5.09 $Y2=1.335
r172 17 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.85 $Y=1.485
+ $X2=4.85 $Y2=1.41
r173 17 19 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.85 $Y=1.485
+ $X2=4.85 $Y2=2.315
r174 16 55 22.8359 $w=2.7e-07 $l=9.28709e-08 $layer=POLY_cond $X=4.265 $Y=1.41
+ $X2=4.19 $Y2=1.45
r175 15 28 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.85 $Y2=1.41
r176 15 16 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.265 $Y2=1.41
r177 11 55 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=1.285
+ $X2=4.19 $Y2=1.45
r178 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.19 $Y=1.285
+ $X2=4.19 $Y2=0.445
r179 7 53 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.735 $Y=1.615
+ $X2=3.735 $Y2=1.45
r180 7 9 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3.735 $Y=1.615
+ $X2=3.735 $Y2=2.525
r181 2 42 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=2.315 $X2=2.62 $Y2=2.52
r182 1 33 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.595 $X2=2.57 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_33_463# 1 2 10 14 15 16 17 18 21 25 27 32
+ 35 37 39 41 44 48 54 56 58
c137 48 0 1.01515e-19 $X=0.7 $Y=1.645
c138 35 0 1.47832e-19 $X=6.36 $Y=0.665
r139 58 59 6.10127 $w=3.16e-07 $l=4e-08 $layer=POLY_cond $X=0.935 $Y=1.645
+ $X2=0.975 $Y2=1.645
r140 51 54 6.3796 $w=2.78e-07 $l=1.55e-07 $layer=LI1_cond $X=0.175 $Y=0.53
+ $X2=0.33 $Y2=0.53
r141 49 58 35.8449 $w=3.16e-07 $l=2.35e-07 $layer=POLY_cond $X=0.7 $Y=1.645
+ $X2=0.935 $Y2=1.645
r142 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.7
+ $Y=1.645 $X2=0.7 $Y2=1.645
r143 46 56 1.15852 $w=2.5e-07 $l=1.53e-07 $layer=LI1_cond $X=0.395 $Y=1.685
+ $X2=0.242 $Y2=1.685
r144 46 48 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.395 $Y=1.685
+ $X2=0.7 $Y2=1.685
r145 42 56 5.39018 $w=2.37e-07 $l=1.25e-07 $layer=LI1_cond $X=0.242 $Y=1.81
+ $X2=0.242 $Y2=1.685
r146 42 44 24.5603 $w=3.03e-07 $l=6.5e-07 $layer=LI1_cond $X=0.242 $Y=1.81
+ $X2=0.242 $Y2=2.46
r147 41 56 5.39018 $w=2.37e-07 $l=1.54919e-07 $layer=LI1_cond $X=0.175 $Y=1.56
+ $X2=0.242 $Y2=1.685
r148 40 51 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.175 $Y=0.67
+ $X2=0.175 $Y2=0.53
r149 40 41 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=0.175 $Y=0.67
+ $X2=0.175 $Y2=1.56
r150 38 39 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=6.342 $Y=1.825
+ $X2=6.342 $Y2=1.975
r151 35 38 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=6.36 $Y=0.665
+ $X2=6.36 $Y2=1.825
r152 32 39 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.325 $Y=2.505
+ $X2=6.325 $Y2=1.975
r153 30 32 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=6.325 $Y=3.075
+ $X2=6.325 $Y2=2.505
r154 28 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.91 $Y=3.15
+ $X2=2.835 $Y2=3.15
r155 27 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.25 $Y=3.15
+ $X2=6.325 $Y2=3.075
r156 27 28 1712.64 $w=1.5e-07 $l=3.34e-06 $layer=POLY_cond $X=6.25 $Y=3.15
+ $X2=2.91 $Y2=3.15
r157 23 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.835 $Y=3.075
+ $X2=2.835 $Y2=3.15
r158 23 25 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.835 $Y=3.075
+ $X2=2.835 $Y2=2.525
r159 19 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.355 $Y=0.255
+ $X2=2.355 $Y2=0.805
r160 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.28 $Y=0.18
+ $X2=2.355 $Y2=0.255
r161 17 18 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=2.28 $Y=0.18
+ $X2=1.05 $Y2=0.18
r162 15 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.76 $Y=3.15
+ $X2=2.835 $Y2=3.15
r163 15 16 897.34 $w=1.5e-07 $l=1.75e-06 $layer=POLY_cond $X=2.76 $Y=3.15
+ $X2=1.01 $Y2=3.15
r164 12 59 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.48
+ $X2=0.975 $Y2=1.645
r165 12 14 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=0.975 $Y=1.48
+ $X2=0.975 $Y2=0.58
r166 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.975 $Y=0.255
+ $X2=1.05 $Y2=0.18
r167 11 14 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.975 $Y=0.255
+ $X2=0.975 $Y2=0.58
r168 8 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.935 $Y=3.075
+ $X2=1.01 $Y2=3.15
r169 8 10 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.935 $Y=3.075
+ $X2=0.935 $Y2=2.635
r170 7 58 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.81
+ $X2=0.935 $Y2=1.645
r171 7 10 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=0.935 $Y=1.81
+ $X2=0.935 $Y2=2.635
r172 2 44 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.315 $X2=0.29 $Y2=2.46
r173 1 54 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.37 $X2=0.33 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_1329_65# 1 2 9 12 13 14 17 19 23 25 27 31
+ 34 36
c89 36 0 1.61779e-19 $X=7.825 $Y=0.4
c90 27 0 1.01861e-19 $X=8.65 $Y=0.4
c91 17 0 1.60057e-19 $X=7.4 $Y=2.525
r92 36 39 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=7.825 $Y=0.4
+ $X2=7.825 $Y2=0.63
r93 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.745
+ $Y=2.56 $X2=8.745 $Y2=2.56
r94 31 33 33.3385 $w=2.78e-07 $l=8.1e-07 $layer=LI1_cond $X=8.79 $Y=1.75
+ $X2=8.79 $Y2=2.56
r95 29 31 52.0657 $w=2.78e-07 $l=1.265e-06 $layer=LI1_cond $X=8.79 $Y=0.485
+ $X2=8.79 $Y2=1.75
r96 28 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.99 $Y=0.4
+ $X2=7.825 $Y2=0.4
r97 27 29 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=8.65 $Y=0.4
+ $X2=8.79 $Y2=0.485
r98 27 28 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.65 $Y=0.4 $X2=7.99
+ $Y2=0.4
r99 26 34 90.0536 $w=3.3e-07 $l=5.15e-07 $layer=POLY_cond $X=8.745 $Y=3.075
+ $X2=8.745 $Y2=2.56
r100 21 23 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.72 $Y=1.935
+ $X2=6.91 $Y2=1.935
r101 20 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.475 $Y=3.15
+ $X2=7.4 $Y2=3.15
r102 19 26 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.58 $Y=3.15
+ $X2=8.745 $Y2=3.075
r103 19 20 566.606 $w=1.5e-07 $l=1.105e-06 $layer=POLY_cond $X=8.58 $Y=3.15
+ $X2=7.475 $Y2=3.15
r104 15 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.4 $Y=3.075
+ $X2=7.4 $Y2=3.15
r105 15 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.4 $Y=3.075
+ $X2=7.4 $Y2=2.525
r106 13 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.325 $Y=3.15
+ $X2=7.4 $Y2=3.15
r107 13 14 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.325 $Y=3.15
+ $X2=6.985 $Y2=3.15
r108 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.91 $Y=3.075
+ $X2=6.985 $Y2=3.15
r109 11 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.91 $Y=2.01
+ $X2=6.91 $Y2=1.935
r110 11 12 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=6.91 $Y=2.01
+ $X2=6.91 $Y2=3.075
r111 7 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.72 $Y=1.86
+ $X2=6.72 $Y2=1.935
r112 7 9 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=6.72 $Y=1.86
+ $X2=6.72 $Y2=0.665
r113 2 31 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.625
+ $Y=1.605 $X2=8.765 $Y2=1.75
r114 1 39 182 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_NDIFF $count=1 $X=7.665
+ $Y=0.455 $X2=7.825 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_1175_417# 1 2 3 10 12 13 14 17 19 21 23 26
+ 30 31 34 40 41 42 45 48 50 51 52 55 56
c117 30 0 4.15052e-20 $X=8.385 $Y=1.26
c118 10 0 1.99629e-19 $X=7.59 $Y=0.345
r119 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.31
+ $Y=0.83 $X2=8.31 $Y2=0.83
r120 52 54 9.02528 $w=5.38e-07 $l=3.98e-07 $layer=LI1_cond $X=7.912 $Y=1
+ $X2=8.31 $Y2=1
r121 50 51 9.53052 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=6.235 $Y=2.21
+ $X2=6.405 $Y2=2.21
r122 46 56 3.49088 $w=2.67e-07 $l=1.08305e-07 $layer=LI1_cond $X=8.01 $Y=2.265
+ $X2=7.957 $Y2=2.18
r123 46 48 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=8.01 $Y=2.265
+ $X2=8.01 $Y2=2.525
r124 45 56 3.49088 $w=2.67e-07 $l=1.05119e-07 $layer=LI1_cond $X=7.912 $Y=2.095
+ $X2=7.957 $Y2=2.18
r125 44 52 4.68134 $w=2.75e-07 $l=3.35e-07 $layer=LI1_cond $X=7.912 $Y=1.335
+ $X2=7.912 $Y2=1
r126 44 45 31.8493 $w=2.73e-07 $l=7.6e-07 $layer=LI1_cond $X=7.912 $Y=1.335
+ $X2=7.912 $Y2=2.095
r127 42 56 3.01551 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.775 $Y=2.18
+ $X2=7.957 $Y2=2.18
r128 42 51 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=7.775 $Y=2.18
+ $X2=6.405 $Y2=2.18
r129 40 52 9.31536 $w=5.38e-07 $l=1.41912e-07 $layer=LI1_cond $X=7.775 $Y=0.99
+ $X2=7.912 $Y2=1
r130 40 41 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=7.775 $Y=0.99
+ $X2=6.305 $Y2=0.99
r131 38 50 7.85757 $w=2.18e-07 $l=1.5e-07 $layer=LI1_cond $X=6.085 $Y=2.215
+ $X2=6.235 $Y2=2.215
r132 32 41 8.54503 $w=1.7e-07 $l=2.48898e-07 $layer=LI1_cond $X=6.095 $Y=0.905
+ $X2=6.305 $Y2=0.99
r133 32 34 14.1311 $w=4.18e-07 $l=5.15e-07 $layer=LI1_cond $X=6.095 $Y=0.905
+ $X2=6.095 $Y2=0.39
r134 29 55 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=8.31 $Y=1.185
+ $X2=8.31 $Y2=0.83
r135 29 30 13.5877 $w=2.4e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.31 $Y=1.185
+ $X2=8.385 $Y2=1.26
r136 28 55 84.8077 $w=3.3e-07 $l=4.85e-07 $layer=POLY_cond $X=8.31 $Y=0.345
+ $X2=8.31 $Y2=0.83
r137 24 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.5 $Y=1.335
+ $X2=9.5 $Y2=1.26
r138 24 26 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=9.5 $Y=1.335
+ $X2=9.5 $Y2=2.155
r139 21 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.5 $Y=1.185
+ $X2=9.5 $Y2=1.26
r140 21 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.5 $Y=1.185
+ $X2=9.5 $Y2=0.865
r141 20 30 12.1617 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.625 $Y=1.26
+ $X2=8.385 $Y2=1.26
r142 19 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.425 $Y=1.26
+ $X2=9.5 $Y2=1.26
r143 19 20 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=9.425 $Y=1.26
+ $X2=8.625 $Y2=1.26
r144 15 30 13.5877 $w=2.4e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.55 $Y=1.335
+ $X2=8.385 $Y2=1.26
r145 15 17 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.55 $Y=1.335
+ $X2=8.55 $Y2=1.815
r146 13 28 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.145 $Y=0.27
+ $X2=8.31 $Y2=0.345
r147 13 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.145 $Y=0.27
+ $X2=7.665 $Y2=0.27
r148 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.59 $Y=0.345
+ $X2=7.665 $Y2=0.27
r149 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.59 $Y=0.345
+ $X2=7.59 $Y2=0.665
r150 3 48 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.905
+ $Y=2.315 $X2=8.045 $Y2=2.525
r151 2 38 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.875
+ $Y=2.085 $X2=6.085 $Y2=2.23
r152 1 34 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=5.91
+ $Y=0.235 $X2=6.05 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_1832_131# 1 2 9 13 17 21 25 26 28
c42 21 0 1.94585e-19 $X=9.285 $Y=1.98
r43 26 31 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.972 $Y=1.48
+ $X2=9.972 $Y2=1.645
r44 26 30 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.972 $Y=1.48
+ $X2=9.972 $Y2=1.315
r45 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.95
+ $Y=1.48 $X2=9.95 $Y2=1.48
r46 23 28 0.630948 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=9.39 $Y=1.48
+ $X2=9.255 $Y2=1.48
r47 23 25 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=9.39 $Y=1.48
+ $X2=9.95 $Y2=1.48
r48 19 28 6.08426 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.255 $Y=1.645
+ $X2=9.255 $Y2=1.48
r49 19 21 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.255 $Y=1.645
+ $X2=9.255 $Y2=1.98
r50 15 28 6.08426 $w=2.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.255 $Y=1.315
+ $X2=9.255 $Y2=1.48
r51 15 17 19.2074 $w=2.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.255 $Y=1.315
+ $X2=9.255 $Y2=0.865
r52 13 31 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=10.085 $Y=2.465
+ $X2=10.085 $Y2=1.645
r53 9 30 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.01 $Y=0.655
+ $X2=10.01 $Y2=1.315
r54 2 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=9.16
+ $Y=1.835 $X2=9.285 $Y2=1.98
r55 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.16
+ $Y=0.655 $X2=9.285 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%VPWR 1 2 3 4 5 6 7 24 28 32 34 35 38 41 44
+ 49 50 54 55 57 60 62 67 79 90 94 101 102 105 108 111 114 117
r135 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r136 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r137 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r139 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 102 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r141 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r142 99 117 10.9443 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=10.035 $Y=3.33
+ $X2=9.797 $Y2=3.33
r143 99 101 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.035 $Y=3.33
+ $X2=10.32 $Y2=3.33
r144 98 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r145 98 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.4 $Y2=3.33
r146 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r147 95 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.48 $Y=3.33
+ $X2=8.395 $Y2=3.33
r148 95 97 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=8.48 $Y=3.33
+ $X2=9.36 $Y2=3.33
r149 94 117 10.9443 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=9.56 $Y=3.33
+ $X2=9.797 $Y2=3.33
r150 94 97 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.56 $Y=3.33 $X2=9.36
+ $Y2=3.33
r151 93 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r152 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r153 90 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.31 $Y=3.33
+ $X2=8.395 $Y2=3.33
r154 90 92 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.31 $Y=3.33
+ $X2=7.92 $Y2=3.33
r155 89 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r156 88 89 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r157 86 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 85 88 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r159 85 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r160 83 111 10.508 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=4.507 $Y2=3.33
r161 83 85 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=5.04 $Y2=3.33
r162 82 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r163 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r164 79 111 10.508 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.507 $Y2=3.33
r165 79 81 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.08 $Y2=3.33
r166 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r167 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r168 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r169 75 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r170 74 77 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r171 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r172 72 108 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=1.745 $Y2=3.33
r173 72 74 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.895 $Y=3.33
+ $X2=2.16 $Y2=3.33
r174 71 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r175 71 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r176 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r177 68 105 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.72 $Y2=3.33
r178 68 70 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=1.2 $Y2=3.33
r179 67 108 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.745 $Y2=3.33
r180 67 70 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.2 $Y2=3.33
r181 65 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r182 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r183 62 105 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.72 $Y2=3.33
r184 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r185 60 89 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=7.44 $Y2=3.33
r186 60 86 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r187 57 59 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.355 $Y=1.76
+ $X2=8.355 $Y2=1.925
r188 54 88 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.53 $Y=3.33 $X2=7.44
+ $Y2=3.33
r189 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.53 $Y=3.33
+ $X2=7.615 $Y2=3.33
r190 53 92 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.7 $Y=3.33
+ $X2=7.92 $Y2=3.33
r191 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.7 $Y=3.33
+ $X2=7.615 $Y2=3.33
r192 49 77 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.12 $Y2=3.33
r193 49 50 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.437 $Y2=3.33
r194 48 81 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.58 $Y=3.33 $X2=4.08
+ $Y2=3.33
r195 48 50 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.58 $Y=3.33
+ $X2=3.437 $Y2=3.33
r196 44 47 11.709 $w=4.73e-07 $l=4.65e-07 $layer=LI1_cond $X=9.797 $Y=2.02
+ $X2=9.797 $Y2=2.485
r197 42 117 1.94084 $w=4.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.797 $Y=3.245
+ $X2=9.797 $Y2=3.33
r198 42 47 19.1373 $w=4.73e-07 $l=7.6e-07 $layer=LI1_cond $X=9.797 $Y=3.245
+ $X2=9.797 $Y2=2.485
r199 41 114 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.395 $Y=3.245
+ $X2=8.395 $Y2=3.33
r200 41 59 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=8.395 $Y=3.245
+ $X2=8.395 $Y2=1.925
r201 36 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.615 $Y=3.245
+ $X2=7.615 $Y2=3.33
r202 36 38 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=7.615 $Y=3.245
+ $X2=7.615 $Y2=2.6
r203 35 111 1.76584 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.507 $Y=3.245
+ $X2=4.507 $Y2=3.33
r204 34 52 9.04117 $w=4.45e-07 $l=3.07e-07 $layer=LI1_cond $X=4.507 $Y=2.577
+ $X2=4.507 $Y2=2.27
r205 34 35 17.2996 $w=4.43e-07 $l=6.68e-07 $layer=LI1_cond $X=4.507 $Y=2.577
+ $X2=4.507 $Y2=3.245
r206 30 50 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.437 $Y=3.245
+ $X2=3.437 $Y2=3.33
r207 30 32 29.1143 $w=2.83e-07 $l=7.2e-07 $layer=LI1_cond $X=3.437 $Y=3.245
+ $X2=3.437 $Y2=2.525
r208 26 108 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=3.245
+ $X2=1.745 $Y2=3.33
r209 26 28 27.6586 $w=2.98e-07 $l=7.2e-07 $layer=LI1_cond $X=1.745 $Y=3.245
+ $X2=1.745 $Y2=2.525
r210 22 105 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r211 22 24 28.8111 $w=3.08e-07 $l=7.75e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.47
r212 7 47 300 $w=1.7e-07 $l=7.83741e-07 $layer=licon1_PDIFF $count=2 $X=9.575
+ $Y=1.835 $X2=9.87 $Y2=2.485
r213 7 44 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=9.575
+ $Y=1.835 $X2=9.775 $Y2=2.02
r214 6 57 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.605 $X2=8.335 $Y2=1.76
r215 5 38 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=7.475
+ $Y=2.315 $X2=7.615 $Y2=2.6
r216 4 52 300 $w=1.7e-07 $l=4.16893e-07 $layer=licon1_PDIFF $count=2 $X=4.24
+ $Y=2.315 $X2=4.635 $Y2=2.27
r217 3 32 600 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=2.315 $X2=3.46 $Y2=2.525
r218 2 28 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.635
+ $Y=2.315 $X2=1.76 $Y2=2.525
r219 1 24 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=2.315 $X2=0.72 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_400_119# 1 2 9 13 16 19 23
r51 16 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=2.015
+ $X2=2.49 $Y2=2.1
r52 15 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=1.345
+ $X2=2.49 $Y2=1.26
r53 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.49 $Y=1.345
+ $X2=2.49 $Y2=2.015
r54 11 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.175 $Y=2.1
+ $X2=2.49 $Y2=2.1
r55 11 13 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=2.175 $Y=2.185
+ $X2=2.175 $Y2=2.525
r56 7 19 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.125 $Y=1.26
+ $X2=2.49 $Y2=1.26
r57 7 9 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.125 $Y=1.175
+ $X2=2.125 $Y2=0.805
r58 2 13 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=2.315 $X2=2.19 $Y2=2.525
r59 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.595
+ $X2=2.14 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_985_379# 1 2 9 11 13
r26 11 13 67.4659 $w=2.38e-07 $l=1.405e-06 $layer=LI1_cond $X=5.23 $Y=2.955
+ $X2=6.635 $Y2=2.955
r27 7 11 7.03987 $w=2.4e-07 $l=2.16852e-07 $layer=LI1_cond $X=5.065 $Y=2.835
+ $X2=5.23 $Y2=2.955
r28 7 9 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=5.065 $Y=2.835
+ $X2=5.065 $Y2=2.22
r29 2 13 600 $w=1.7e-07 $l=9.55301e-07 $layer=licon1_PDIFF $count=1 $X=6.4
+ $Y=2.085 $X2=6.635 $Y2=2.93
r30 1 9 300 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_PDIFF $count=2 $X=4.925
+ $Y=1.895 $X2=5.065 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%A_1092_417# 1 2 9 12 14 15
r26 14 15 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.185 $Y=2.55
+ $X2=7.02 $Y2=2.55
r27 12 15 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=5.75 $Y=2.58
+ $X2=7.02 $Y2=2.58
r28 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.585 $Y=2.495
+ $X2=5.75 $Y2=2.58
r29 7 9 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.585 $Y=2.495
+ $X2=5.585 $Y2=2.29
r30 2 14 600 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_PDIFF $count=1 $X=7.06
+ $Y=2.315 $X2=7.185 $Y2=2.56
r31 1 9 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=2.085 $X2=5.585 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%Q 1 2 9 12 13 14 15 16 17
r17 17 35 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=10.34 $Y=2.775
+ $X2=10.34 $Y2=2.91
r18 16 17 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.34 $Y=2.405
+ $X2=10.34 $Y2=2.775
r19 15 16 16.6464 $w=2.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.34 $Y=2.015
+ $X2=10.34 $Y2=2.405
r20 14 15 14.9391 $w=2.68e-07 $l=3.5e-07 $layer=LI1_cond $X=10.34 $Y=1.665
+ $X2=10.34 $Y2=2.015
r21 13 14 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.34 $Y=1.295
+ $X2=10.34 $Y2=1.665
r22 12 13 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=10.34 $Y=1.095
+ $X2=10.34 $Y2=1.295
r23 7 12 6.74395 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=10.285 $Y=0.905
+ $X2=10.285 $Y2=1.095
r24 7 9 14.7088 $w=3.78e-07 $l=4.85e-07 $layer=LI1_cond $X=10.285 $Y=0.905
+ $X2=10.285 $Y2=0.42
r25 2 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.835 $X2=10.3 $Y2=2.91
r26 2 15 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.835 $X2=10.3 $Y2=2.015
r27 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=10.085
+ $Y=0.235 $X2=10.225 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_1%VGND 1 2 3 4 5 6 23 27 31 35 39 43 45 50 58
+ 63 71 78 79 82 85 88 94 98 101
c123 94 0 4.26559e-20 $X=5.26 $Y=0.38
c124 23 0 1.29179e-19 $X=0.76 $Y=0.505
r125 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r126 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r127 94 96 1.1443 $w=6.93e-07 $l=6.5e-08 $layer=LI1_cond $X=5.012 $Y=0.38
+ $X2=5.012 $Y2=0.445
r128 91 94 6.68975 $w=6.93e-07 $l=3.8e-07 $layer=LI1_cond $X=5.012 $Y=0
+ $X2=5.012 $Y2=0.38
r129 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r130 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r131 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r132 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r133 79 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r134 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r135 76 101 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=9.925 $Y=0
+ $X2=9.747 $Y2=0
r136 76 78 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.925 $Y=0
+ $X2=10.32 $Y2=0
r137 75 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r138 75 99 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=7.44 $Y2=0
r139 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r140 72 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.46 $Y=0 $X2=7.295
+ $Y2=0
r141 72 74 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=7.46 $Y=0 $X2=9.36
+ $Y2=0
r142 71 101 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=9.57 $Y=0
+ $X2=9.747 $Y2=0
r143 71 74 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.57 $Y=0 $X2=9.36
+ $Y2=0
r144 70 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r145 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r146 67 70 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.96 $Y2=0
r147 66 69 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=6.96
+ $Y2=0
r148 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r149 64 91 9.25536 $w=1.7e-07 $l=4.13e-07 $layer=LI1_cond $X=5.425 $Y=0
+ $X2=5.012 $Y2=0
r150 64 66 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.425 $Y=0 $X2=5.52
+ $Y2=0
r151 63 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.13 $Y=0 $X2=7.295
+ $Y2=0
r152 63 69 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.13 $Y=0 $X2=6.96
+ $Y2=0
r153 62 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r154 62 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r155 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r156 59 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.455
+ $Y2=0
r157 59 61 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=4.56
+ $Y2=0
r158 58 91 9.25536 $w=1.7e-07 $l=4.12e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=5.012
+ $Y2=0
r159 58 61 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.56
+ $Y2=0
r160 57 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r161 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r162 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r163 54 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r164 53 56 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r165 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r166 51 85 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=1.695
+ $Y2=0
r167 51 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.845 $Y=0
+ $X2=2.16 $Y2=0
r168 50 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=0 $X2=3.455
+ $Y2=0
r169 50 56 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.29 $Y=0 $X2=3.12
+ $Y2=0
r170 49 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r171 49 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r172 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r173 46 82 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.765
+ $Y2=0
r174 46 48 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r175 45 85 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.695
+ $Y2=0
r176 45 48 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.2
+ $Y2=0
r177 43 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.52 $Y2=0
r178 43 92 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.04 $Y2=0
r179 39 41 17.6924 $w=3.53e-07 $l=5.45e-07 $layer=LI1_cond $X=9.747 $Y=0.385
+ $X2=9.747 $Y2=0.93
r180 37 101 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=9.747 $Y=0.085
+ $X2=9.747 $Y2=0
r181 37 39 9.73895 $w=3.53e-07 $l=3e-07 $layer=LI1_cond $X=9.747 $Y=0.085
+ $X2=9.747 $Y2=0.385
r182 33 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0
r183 33 35 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=7.295 $Y=0.085
+ $X2=7.295 $Y2=0.625
r184 29 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0
r185 29 31 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0.67
r186 25 85 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0
r187 25 27 27.6586 $w=2.98e-07 $l=7.2e-07 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0.805
r188 21 82 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0
r189 21 23 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0.505
r190 6 41 182 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_NDIFF $count=1 $X=9.575
+ $Y=0.655 $X2=9.735 $Y2=0.93
r191 6 39 182 $w=1.7e-07 $l=3.63731e-07 $layer=licon1_NDIFF $count=1 $X=9.575
+ $Y=0.655 $X2=9.795 $Y2=0.385
r192 5 35 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=7.155
+ $Y=0.455 $X2=7.295 $Y2=0.625
r193 4 96 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.235 $X2=4.765 $Y2=0.445
r194 4 94 91 $w=1.7e-07 $l=7.03776e-07 $layer=licon1_NDIFF $count=2 $X=4.625
+ $Y=0.235 $X2=5.26 $Y2=0.38
r195 3 31 182 $w=1.7e-07 $l=2.69907e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.595 $X2=3.455 $Y2=0.67
r196 2 27 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.595 $X2=1.71 $Y2=0.805
r197 1 23 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.37 $X2=0.76 $Y2=0.505
.ends

