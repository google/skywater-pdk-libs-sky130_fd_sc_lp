* NGSPICE file created from sky130_fd_sc_lp__o41ai_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o41ai_lp A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_153_57# A3 VGND VNB nshort w=420000u l=150000u
+  ad=3.549e+11p pd=4.21e+06u as=3.906e+11p ps=3.54e+06u
M1001 a_359_419# A3 a_259_419# VPB phighvt w=1e+06u l=250000u
+  ad=3.2e+11p pd=2.64e+06u as=2.5e+11p ps=2.5e+06u
M1002 Y B1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.8e+11p pd=2.56e+06u as=5.7e+11p ps=5.14e+06u
M1003 VGND A4 a_153_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A2 a_153_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_153_57# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A1 a_473_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1007 a_153_57# B1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.533e+11p ps=1.57e+06u
M1008 a_473_419# A2 a_359_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_259_419# A4 Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

