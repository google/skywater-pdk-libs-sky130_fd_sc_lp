* File: sky130_fd_sc_lp__a2111oi_2.pxi.spice
* Created: Fri Aug 28 09:46:49 2020
* 
x_PM_SKY130_FD_SC_LP__A2111OI_2%C1 N_C1_M1012_g N_C1_M1005_g N_C1_M1008_g
+ N_C1_M1017_g N_C1_c_104_n N_C1_c_105_n C1 N_C1_c_106_n N_C1_c_107_n
+ N_C1_c_108_n PM_SKY130_FD_SC_LP__A2111OI_2%C1
x_PM_SKY130_FD_SC_LP__A2111OI_2%D1 N_D1_c_173_n N_D1_M1007_g N_D1_M1009_g
+ N_D1_c_175_n N_D1_M1015_g N_D1_M1016_g D1 D1 N_D1_c_178_n
+ PM_SKY130_FD_SC_LP__A2111OI_2%D1
x_PM_SKY130_FD_SC_LP__A2111OI_2%B1 N_B1_M1001_g N_B1_M1003_g N_B1_M1010_g
+ N_B1_M1011_g B1 B1 N_B1_c_226_n N_B1_c_227_n PM_SKY130_FD_SC_LP__A2111OI_2%B1
x_PM_SKY130_FD_SC_LP__A2111OI_2%A1 N_A1_M1000_g N_A1_M1002_g N_A1_M1013_g
+ N_A1_M1014_g N_A1_c_274_n N_A1_c_275_n N_A1_c_276_n A1 A1 N_A1_c_277_n
+ N_A1_c_278_n N_A1_c_279_n PM_SKY130_FD_SC_LP__A2111OI_2%A1
x_PM_SKY130_FD_SC_LP__A2111OI_2%A2 N_A2_c_349_n N_A2_M1004_g N_A2_M1006_g
+ N_A2_c_351_n N_A2_M1018_g N_A2_M1019_g N_A2_c_353_n A2 N_A2_c_355_n
+ N_A2_c_356_n PM_SKY130_FD_SC_LP__A2111OI_2%A2
x_PM_SKY130_FD_SC_LP__A2111OI_2%A_32_367# N_A_32_367#_M1005_d
+ N_A_32_367#_M1008_d N_A_32_367#_M1010_s N_A_32_367#_c_408_n
+ N_A_32_367#_c_409_n N_A_32_367#_c_413_n N_A_32_367#_c_427_p
+ N_A_32_367#_c_410_n N_A_32_367#_c_436_p
+ PM_SKY130_FD_SC_LP__A2111OI_2%A_32_367#
x_PM_SKY130_FD_SC_LP__A2111OI_2%A_115_367# N_A_115_367#_M1005_s
+ N_A_115_367#_M1016_d N_A_115_367#_c_444_n N_A_115_367#_c_447_n
+ N_A_115_367#_c_446_n N_A_115_367#_c_453_n
+ PM_SKY130_FD_SC_LP__A2111OI_2%A_115_367#
x_PM_SKY130_FD_SC_LP__A2111OI_2%Y N_Y_M1012_d N_Y_M1007_s N_Y_M1017_d
+ N_Y_M1011_s N_Y_M1013_s N_Y_M1009_s N_Y_c_461_n N_Y_c_473_n N_Y_c_462_n
+ N_Y_c_478_n N_Y_c_479_n N_Y_c_483_n N_Y_c_487_n N_Y_c_463_n N_Y_c_509_n
+ N_Y_c_469_n N_Y_c_464_n N_Y_c_488_n N_Y_c_498_n N_Y_c_465_n N_Y_c_466_n Y Y Y
+ Y PM_SKY130_FD_SC_LP__A2111OI_2%Y
x_PM_SKY130_FD_SC_LP__A2111OI_2%A_467_367# N_A_467_367#_M1001_d
+ N_A_467_367#_M1002_s N_A_467_367#_M1006_d N_A_467_367#_M1014_s
+ N_A_467_367#_c_591_n N_A_467_367#_c_592_n N_A_467_367#_c_598_n
+ N_A_467_367#_c_625_p N_A_467_367#_c_599_n N_A_467_367#_c_593_n
+ N_A_467_367#_c_594_n N_A_467_367#_c_595_n N_A_467_367#_c_618_n
+ PM_SKY130_FD_SC_LP__A2111OI_2%A_467_367#
x_PM_SKY130_FD_SC_LP__A2111OI_2%VPWR N_VPWR_M1002_d N_VPWR_M1018_s
+ N_VPWR_c_636_n N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_640_n
+ N_VPWR_c_641_n VPWR N_VPWR_c_642_n N_VPWR_c_635_n
+ PM_SKY130_FD_SC_LP__A2111OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A2111OI_2%VGND N_VGND_M1012_s N_VGND_M1015_d
+ N_VGND_M1003_d N_VGND_M1004_s N_VGND_c_702_n N_VGND_c_703_n N_VGND_c_704_n
+ N_VGND_c_705_n N_VGND_c_706_n N_VGND_c_707_n VGND N_VGND_c_708_n
+ N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n N_VGND_c_712_n N_VGND_c_713_n
+ N_VGND_c_714_n N_VGND_c_715_n PM_SKY130_FD_SC_LP__A2111OI_2%VGND
x_PM_SKY130_FD_SC_LP__A2111OI_2%A_684_47# N_A_684_47#_M1000_d
+ N_A_684_47#_M1019_d N_A_684_47#_c_773_n N_A_684_47#_c_774_n
+ N_A_684_47#_c_776_n N_A_684_47#_c_793_n
+ PM_SKY130_FD_SC_LP__A2111OI_2%A_684_47#
cc_1 VNB N_C1_M1012_g 0.0310872f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_2 VNB N_C1_M1005_g 0.00167964f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_3 VNB N_C1_M1008_g 0.00128182f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.465
cc_4 VNB N_C1_M1017_g 0.0245225f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.655
cc_5 VNB N_C1_c_104_n 0.00660143f $X=-0.19 $Y=-0.245 $X2=1.525 $Y2=1.69
cc_6 VNB N_C1_c_105_n 0.00436011f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_7 VNB N_C1_c_106_n 0.0565962f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.46
cc_8 VNB N_C1_c_107_n 0.030946f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.46
cc_9 VNB N_C1_c_108_n 0.00609175f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.46
cc_10 VNB N_D1_c_173_n 0.016201f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.295
cc_11 VNB N_D1_M1009_g 0.00680537f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_12 VNB N_D1_c_175_n 0.0173798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D1_M1016_g 0.00648617f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=1.295
cc_14 VNB D1 0.00628515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_D1_c_178_n 0.0364545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_M1003_g 0.0254101f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_17 VNB N_B1_M1011_g 0.0246525f $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.655
cc_18 VNB N_B1_c_226_n 0.00248748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_227_n 0.0446055f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_20 VNB N_A1_M1000_g 0.0271945f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.655
cc_21 VNB N_A1_M1013_g 0.0288494f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=2.465
cc_22 VNB N_A1_c_274_n 0.00660959f $X=-0.19 $Y=-0.245 $X2=1.525 $Y2=1.69
cc_23 VNB N_A1_c_275_n 0.00117023f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_24 VNB N_A1_c_276_n 0.0285696f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_25 VNB N_A1_c_277_n 0.0337245f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.295
cc_26 VNB N_A1_c_278_n 0.00291389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_c_279_n 0.00319211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_c_349_n 0.0190805f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.295
cc_29 VNB N_A2_M1006_g 0.0131658f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_30 VNB N_A2_c_351_n 0.011605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_M1018_g 0.00707205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_c_353_n 0.00777799f $X=-0.19 $Y=-0.245 $X2=1.525 $Y2=1.69
cc_33 VNB A2 0.00257775f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.69
cc_34 VNB N_A2_c_355_n 0.0246865f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_35 VNB N_A2_c_356_n 0.0170526f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_36 VNB N_Y_c_461_n 0.0233935f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_37 VNB N_Y_c_462_n 0.00766836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_463_n 0.00819344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_464_n 0.0321296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_465_n 0.00385023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_466_n 0.053114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB Y 0.00142546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB Y 0.00340489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VPWR_c_635_n 0.243291f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.625
cc_45 VNB N_VGND_c_702_n 4.08532e-19 $X=-0.19 $Y=-0.245 $X2=1.9 $Y2=0.655
cc_46 VNB N_VGND_c_703_n 0.00437091f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_47 VNB N_VGND_c_704_n 0.00504266f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.69
cc_48 VNB N_VGND_c_705_n 0.00561423f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_49 VNB N_VGND_c_706_n 0.0358113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_707_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.46
cc_51 VNB N_VGND_c_708_n 0.0161714f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.295
cc_52 VNB N_VGND_c_709_n 0.0152636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_710_n 0.0180522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_711_n 0.0354435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_712_n 0.292458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_713_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_714_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_715_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_C1_M1005_g 0.0252493f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_60 VPB N_C1_M1008_g 0.0195885f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=2.465
cc_61 VPB N_C1_c_104_n 0.00688527f $X=-0.19 $Y=1.655 $X2=1.525 $Y2=1.69
cc_62 VPB N_C1_c_105_n 0.00808067f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_63 VPB N_C1_c_108_n 0.00302903f $X=-0.19 $Y=1.655 $X2=1.81 $Y2=1.46
cc_64 VPB N_D1_M1009_g 0.0189866f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_65 VPB N_D1_M1016_g 0.0189866f $X=-0.19 $Y=1.655 $X2=1.9 $Y2=1.295
cc_66 VPB N_B1_M1001_g 0.0185357f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.655
cc_67 VPB N_B1_M1010_g 0.0224575f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=2.465
cc_68 VPB N_B1_c_226_n 0.00622855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_B1_c_227_n 0.0115954f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_70 VPB N_A1_M1002_g 0.0223792f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_71 VPB N_A1_M1014_g 0.0228363f $X=-0.19 $Y=1.655 $X2=1.9 $Y2=0.655
cc_72 VPB N_A1_c_274_n 0.00509854f $X=-0.19 $Y=1.655 $X2=1.525 $Y2=1.69
cc_73 VPB N_A1_c_275_n 0.00203394f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_74 VPB N_A1_c_276_n 0.00642776f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_75 VPB N_A1_c_277_n 0.00971062f $X=-0.19 $Y=1.655 $X2=1.81 $Y2=1.295
cc_76 VPB N_A1_c_278_n 0.00412729f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A1_c_279_n 6.53693e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A2_M1006_g 0.0186439f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_79 VPB N_A2_M1018_g 0.0191203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_32_367#_c_408_n 0.00915464f $X=-0.19 $Y=1.655 $X2=1.79 $Y2=2.465
cc_81 VPB N_A_32_367#_c_409_n 0.0349476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_32_367#_c_410_n 0.00299093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_Y_c_469_n 0.0225609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_Y_c_464_n 0.0175309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB Y 0.00437508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB Y 0.00513515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_467_367#_c_591_n 0.0080356f $X=-0.19 $Y=1.655 $X2=1.9 $Y2=1.295
cc_88 VPB N_A_467_367#_c_592_n 0.00511077f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_89 VPB N_A_467_367#_c_593_n 0.00754096f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.46
cc_90 VPB N_A_467_367#_c_594_n 0.0234065f $X=-0.19 $Y=1.655 $X2=1.81 $Y2=1.46
cc_91 VPB N_A_467_367#_c_595_n 8.35298e-19 $X=-0.19 $Y=1.655 $X2=1.81 $Y2=1.295
cc_92 VPB N_VPWR_c_636_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=1.79 $Y2=1.625
cc_93 VPB N_VPWR_c_637_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=1.9 $Y2=1.295
cc_94 VPB N_VPWR_c_638_n 0.0867886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_639_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.525 $Y2=1.69
cc_96 VPB N_VPWR_c_640_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_97 VPB N_VPWR_c_641_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_98 VPB N_VPWR_c_642_n 0.0258481f $X=-0.19 $Y=1.655 $X2=1.81 $Y2=1.295
cc_99 VPB N_VPWR_c_635_n 0.0624103f $X=-0.19 $Y=1.655 $X2=1.81 $Y2=1.625
cc_100 N_C1_M1012_g N_D1_c_173_n 0.0302991f $X=0.5 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_101 N_C1_M1005_g N_D1_M1009_g 0.0302991f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_102 N_C1_c_104_n N_D1_M1009_g 0.0148037f $X=1.525 $Y=1.69 $X2=0 $Y2=0
cc_103 N_C1_M1017_g N_D1_c_175_n 0.0239381f $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_104 N_C1_M1008_g N_D1_M1016_g 0.0563404f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_105 N_C1_c_104_n N_D1_M1016_g 0.0104497f $X=1.525 $Y=1.69 $X2=0 $Y2=0
cc_106 N_C1_c_108_n N_D1_M1016_g 2.47149e-19 $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_107 N_C1_M1012_g D1 0.00397349f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_108 N_C1_M1017_g D1 4.1474e-19 $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_109 N_C1_c_104_n D1 0.0533828f $X=1.525 $Y=1.69 $X2=0 $Y2=0
cc_110 N_C1_c_105_n D1 0.0117206f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_111 N_C1_c_108_n D1 0.0117644f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_112 N_C1_c_104_n N_D1_c_178_n 0.00246472f $X=1.525 $Y=1.69 $X2=0 $Y2=0
cc_113 N_C1_c_105_n N_D1_c_178_n 0.00100972f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_114 N_C1_c_106_n N_D1_c_178_n 0.0302991f $X=0.5 $Y=1.46 $X2=0 $Y2=0
cc_115 N_C1_c_107_n N_D1_c_178_n 0.0207278f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_116 N_C1_c_108_n N_D1_c_178_n 0.00549537f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_117 N_C1_M1017_g N_B1_M1003_g 0.0191151f $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_118 N_C1_c_108_n N_B1_M1003_g 2.56577e-19 $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_119 N_C1_M1008_g N_B1_c_226_n 5.73065e-19 $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_120 N_C1_c_107_n N_B1_c_226_n 0.00143544f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_121 N_C1_c_108_n N_B1_c_226_n 0.030199f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_122 N_C1_M1008_g N_B1_c_227_n 0.0338122f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_123 N_C1_c_107_n N_B1_c_227_n 0.018237f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_124 N_C1_c_108_n N_B1_c_227_n 0.00110112f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_125 N_C1_c_105_n N_A_32_367#_c_409_n 0.022163f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_126 N_C1_c_106_n N_A_32_367#_c_409_n 0.00143676f $X=0.5 $Y=1.46 $X2=0 $Y2=0
cc_127 N_C1_M1005_g N_A_32_367#_c_413_n 0.01317f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_128 N_C1_M1008_g N_A_32_367#_c_413_n 0.0133817f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_129 N_C1_M1005_g N_A_115_367#_c_444_n 0.00546781f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_130 N_C1_c_104_n N_A_115_367#_c_444_n 0.016611f $X=1.525 $Y=1.69 $X2=0 $Y2=0
cc_131 N_C1_M1005_g N_A_115_367#_c_446_n 0.00158305f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_132 N_C1_M1012_g N_Y_c_473_n 0.0138217f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_133 N_C1_c_104_n N_Y_c_473_n 0.00384587f $X=1.525 $Y=1.69 $X2=0 $Y2=0
cc_134 N_C1_c_105_n N_Y_c_473_n 0.00282338f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_135 N_C1_c_105_n N_Y_c_462_n 0.015481f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_136 N_C1_c_106_n N_Y_c_462_n 0.00186882f $X=0.5 $Y=1.46 $X2=0 $Y2=0
cc_137 N_C1_M1017_g N_Y_c_478_n 4.45014e-19 $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_138 N_C1_M1008_g N_Y_c_479_n 0.0156368f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_139 N_C1_c_104_n N_Y_c_479_n 0.0155623f $X=1.525 $Y=1.69 $X2=0 $Y2=0
cc_140 N_C1_c_107_n N_Y_c_479_n 0.0027101f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_141 N_C1_c_108_n N_Y_c_479_n 0.025653f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_142 N_C1_M1017_g N_Y_c_483_n 0.0150098f $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_143 N_C1_c_104_n N_Y_c_483_n 0.00398103f $X=1.525 $Y=1.69 $X2=0 $Y2=0
cc_144 N_C1_c_107_n N_Y_c_483_n 0.00100408f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_145 N_C1_c_108_n N_Y_c_483_n 0.0193845f $X=1.81 $Y=1.46 $X2=0 $Y2=0
cc_146 N_C1_M1017_g N_Y_c_487_n 0.00883979f $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_147 N_C1_c_104_n N_Y_c_488_n 0.0169962f $X=1.525 $Y=1.69 $X2=0 $Y2=0
cc_148 N_C1_M1017_g N_Y_c_465_n 0.00679627f $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_149 N_C1_M1005_g N_VPWR_c_638_n 0.00357877f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_150 N_C1_M1008_g N_VPWR_c_638_n 0.00357877f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_151 N_C1_M1005_g N_VPWR_c_635_n 0.00633391f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_152 N_C1_M1008_g N_VPWR_c_635_n 0.00549753f $X=1.79 $Y=2.465 $X2=0 $Y2=0
cc_153 N_C1_M1012_g N_VGND_c_702_n 0.0121813f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_154 N_C1_M1017_g N_VGND_c_703_n 0.00268356f $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_155 N_C1_M1012_g N_VGND_c_708_n 0.00486043f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_156 N_C1_M1017_g N_VGND_c_710_n 0.00571722f $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_157 N_C1_M1012_g N_VGND_c_712_n 0.00920269f $X=0.5 $Y=0.655 $X2=0 $Y2=0
cc_158 N_C1_M1017_g N_VGND_c_712_n 0.0108063f $X=1.9 $Y=0.655 $X2=0 $Y2=0
cc_159 N_D1_M1009_g N_A_32_367#_c_413_n 0.0111577f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_160 N_D1_M1016_g N_A_32_367#_c_413_n 0.011213f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_161 N_D1_M1009_g N_A_115_367#_c_447_n 0.0127458f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_162 N_D1_M1016_g N_A_115_367#_c_447_n 0.0097886f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_163 N_D1_c_173_n N_Y_c_473_n 0.0122129f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_164 D1 N_Y_c_473_n 0.0270141f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_165 N_D1_c_175_n N_Y_c_478_n 0.00784816f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_166 N_D1_M1016_g N_Y_c_479_n 0.0100803f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_167 N_D1_c_175_n N_Y_c_483_n 0.0137966f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_168 D1 N_Y_c_483_n 0.00412248f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_169 N_D1_c_175_n N_Y_c_487_n 4.45507e-19 $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_170 N_D1_M1009_g N_Y_c_488_n 0.00413383f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_171 N_D1_c_175_n N_Y_c_498_n 2.74535e-19 $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_172 D1 N_Y_c_498_n 0.0165392f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_173 N_D1_c_178_n N_Y_c_498_n 0.00240082f $X=1.36 $Y=1.35 $X2=0 $Y2=0
cc_174 N_D1_M1009_g N_VPWR_c_638_n 0.00357877f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_175 N_D1_M1016_g N_VPWR_c_638_n 0.00357877f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_176 N_D1_M1009_g N_VPWR_c_635_n 0.00544922f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_177 N_D1_M1016_g N_VPWR_c_635_n 0.00544922f $X=1.36 $Y=2.465 $X2=0 $Y2=0
cc_178 N_D1_c_173_n N_VGND_c_702_n 0.0107016f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_179 N_D1_c_175_n N_VGND_c_702_n 6.28665e-19 $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_180 N_D1_c_175_n N_VGND_c_703_n 0.00257225f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_181 N_D1_c_173_n N_VGND_c_709_n 0.00486043f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_182 N_D1_c_175_n N_VGND_c_709_n 0.00571847f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_183 N_D1_c_173_n N_VGND_c_712_n 0.00824727f $X=0.93 $Y=1.185 $X2=0 $Y2=0
cc_184 N_D1_c_175_n N_VGND_c_712_n 0.0106761f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_185 N_B1_M1011_g N_A1_M1000_g 0.0202198f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_186 N_B1_c_227_n N_A1_c_277_n 0.0202198f $X=2.915 $Y=1.51 $X2=0 $Y2=0
cc_187 N_B1_M1001_g N_A_32_367#_c_410_n 0.0149068f $X=2.26 $Y=2.465 $X2=0 $Y2=0
cc_188 N_B1_M1010_g N_A_32_367#_c_410_n 0.0100622f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_189 N_B1_M1001_g N_Y_c_479_n 0.0156923f $X=2.26 $Y=2.465 $X2=0 $Y2=0
cc_190 N_B1_M1010_g N_Y_c_479_n 0.0130331f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_191 N_B1_c_226_n N_Y_c_479_n 0.0517958f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_192 N_B1_c_227_n N_Y_c_479_n 0.00598493f $X=2.915 $Y=1.51 $X2=0 $Y2=0
cc_193 N_B1_M1003_g N_Y_c_463_n 0.0153809f $X=2.375 $Y=0.655 $X2=0 $Y2=0
cc_194 N_B1_M1011_g N_Y_c_463_n 0.0147291f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_195 N_B1_c_226_n N_Y_c_463_n 0.0416237f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_196 N_B1_c_227_n N_Y_c_463_n 0.00622066f $X=2.915 $Y=1.51 $X2=0 $Y2=0
cc_197 N_B1_M1003_g N_Y_c_509_n 4.0821e-19 $X=2.375 $Y=0.655 $X2=0 $Y2=0
cc_198 N_B1_M1011_g N_Y_c_509_n 0.012425f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_199 N_B1_c_226_n N_Y_c_465_n 0.0199734f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_200 N_B1_c_227_n N_Y_c_465_n 0.00329766f $X=2.915 $Y=1.51 $X2=0 $Y2=0
cc_201 N_B1_M1011_g Y 0.00358694f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_202 N_B1_M1010_g Y 0.00617651f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B1_M1011_g Y 0.00706032f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_204 N_B1_c_226_n Y 0.0292136f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_205 N_B1_M1010_g N_A_467_367#_c_591_n 0.0174574f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_206 N_B1_M1010_g N_A_467_367#_c_592_n 0.00339302f $X=2.69 $Y=2.465 $X2=0
+ $Y2=0
cc_207 N_B1_M1001_g N_VPWR_c_638_n 0.00357877f $X=2.26 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B1_M1010_g N_VPWR_c_638_n 0.00357877f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_209 N_B1_M1001_g N_VPWR_c_635_n 0.00547024f $X=2.26 $Y=2.465 $X2=0 $Y2=0
cc_210 N_B1_M1010_g N_VPWR_c_635_n 0.00665089f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_211 N_B1_M1003_g N_VGND_c_704_n 0.00227546f $X=2.375 $Y=0.655 $X2=0 $Y2=0
cc_212 N_B1_M1011_g N_VGND_c_704_n 0.00700237f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_213 N_B1_M1011_g N_VGND_c_706_n 0.0054895f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_214 N_B1_M1003_g N_VGND_c_710_n 0.00585385f $X=2.375 $Y=0.655 $X2=0 $Y2=0
cc_215 N_B1_M1003_g N_VGND_c_712_n 0.0109254f $X=2.375 $Y=0.655 $X2=0 $Y2=0
cc_216 N_B1_M1011_g N_VGND_c_712_n 0.0101773f $X=2.915 $Y=0.655 $X2=0 $Y2=0
cc_217 N_A1_M1000_g N_A2_c_349_n 0.0205299f $X=3.345 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_218 N_A1_M1000_g N_A2_M1006_g 2.36326e-19 $X=3.345 $Y=0.655 $X2=0 $Y2=0
cc_219 N_A1_c_277_n N_A2_M1006_g 0.0687862f $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_220 N_A1_c_279_n N_A2_M1006_g 0.0192401f $X=4.185 $Y=1.565 $X2=0 $Y2=0
cc_221 N_A1_c_274_n N_A2_c_351_n 0.00357572f $X=4.895 $Y=1.7 $X2=0 $Y2=0
cc_222 N_A1_c_279_n N_A2_c_351_n 0.00137879f $X=4.185 $Y=1.565 $X2=0 $Y2=0
cc_223 N_A1_c_274_n N_A2_M1018_g 0.0107263f $X=4.895 $Y=1.7 $X2=0 $Y2=0
cc_224 N_A1_c_275_n N_A2_M1018_g 7.23036e-19 $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_225 N_A1_c_276_n N_A2_M1018_g 0.0525548f $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_226 N_A1_c_279_n N_A2_M1018_g 0.00253358f $X=4.185 $Y=1.565 $X2=0 $Y2=0
cc_227 N_A1_c_279_n N_A2_c_353_n 8.79738e-19 $X=4.185 $Y=1.565 $X2=0 $Y2=0
cc_228 N_A1_M1013_g A2 0.00191376f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_229 N_A1_c_274_n A2 0.0254515f $X=4.895 $Y=1.7 $X2=0 $Y2=0
cc_230 N_A1_c_275_n A2 0.00706677f $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_231 N_A1_c_279_n A2 0.00760075f $X=4.185 $Y=1.565 $X2=0 $Y2=0
cc_232 N_A1_M1013_g N_A2_c_355_n 0.0208275f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_233 N_A1_c_274_n N_A2_c_355_n 0.00479299f $X=4.895 $Y=1.7 $X2=0 $Y2=0
cc_234 N_A1_c_275_n N_A2_c_355_n 6.77015e-19 $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_235 N_A1_c_279_n N_A2_c_355_n 0.00272805f $X=4.185 $Y=1.565 $X2=0 $Y2=0
cc_236 N_A1_M1013_g N_A2_c_356_n 0.0144943f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_237 N_A1_M1000_g N_Y_c_509_n 0.0126487f $X=3.345 $Y=0.655 $X2=0 $Y2=0
cc_238 N_A1_M1002_g N_Y_c_469_n 0.0124865f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A1_M1014_g N_Y_c_469_n 0.0125146f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A1_c_275_n N_Y_c_469_n 0.0176075f $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_241 N_A1_c_276_n N_Y_c_469_n 0.00285046f $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_242 N_A1_c_277_n N_Y_c_469_n 0.00653136f $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_243 N_A1_c_278_n N_Y_c_469_n 0.0924642f $X=3.965 $Y=1.565 $X2=0 $Y2=0
cc_244 N_A1_M1013_g N_Y_c_464_n 0.00664016f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_245 N_A1_M1014_g N_Y_c_464_n 0.00622183f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A1_c_275_n N_Y_c_464_n 0.0347076f $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_247 N_A1_c_276_n N_Y_c_464_n 0.00817785f $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_248 N_A1_M1013_g N_Y_c_466_n 0.0128725f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_249 N_A1_c_275_n N_Y_c_466_n 0.00849342f $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_250 N_A1_c_276_n N_Y_c_466_n 0.00371886f $X=5.06 $Y=1.51 $X2=0 $Y2=0
cc_251 N_A1_M1000_g Y 0.00610921f $X=3.345 $Y=0.655 $X2=0 $Y2=0
cc_252 N_A1_M1002_g Y 3.69313e-19 $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_253 N_A1_M1000_g Y 0.00294631f $X=3.345 $Y=0.655 $X2=0 $Y2=0
cc_254 N_A1_M1002_g Y 0.00583628f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_255 N_A1_c_277_n Y 0.00897059f $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_256 N_A1_c_278_n Y 0.0354909f $X=3.965 $Y=1.565 $X2=0 $Y2=0
cc_257 N_A1_M1002_g N_A_467_367#_c_598_n 0.0122129f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A1_M1014_g N_A_467_367#_c_599_n 0.0129814f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A1_c_277_n N_A_467_367#_c_595_n 3.23119e-19 $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_260 N_A1_M1002_g N_VPWR_c_636_n 0.0120604f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A1_M1014_g N_VPWR_c_637_n 0.010819f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A1_M1002_g N_VPWR_c_638_n 0.00486043f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A1_M1014_g N_VPWR_c_642_n 0.00564095f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A1_M1002_g N_VPWR_c_635_n 0.00954696f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A1_M1014_g N_VPWR_c_635_n 0.0106077f $X=4.97 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A1_M1000_g N_VGND_c_706_n 0.0054895f $X=3.345 $Y=0.655 $X2=0 $Y2=0
cc_267 N_A1_M1013_g N_VGND_c_711_n 0.0054895f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_268 N_A1_M1000_g N_VGND_c_712_n 0.0106313f $X=3.345 $Y=0.655 $X2=0 $Y2=0
cc_269 N_A1_M1013_g N_VGND_c_712_n 0.0110629f $X=4.97 $Y=0.655 $X2=0 $Y2=0
cc_270 N_A1_M1000_g N_A_684_47#_c_773_n 0.00646387f $X=3.345 $Y=0.655 $X2=0
+ $Y2=0
cc_271 N_A1_c_274_n N_A_684_47#_c_774_n 0.00931302f $X=4.895 $Y=1.7 $X2=0 $Y2=0
cc_272 N_A1_c_278_n N_A_684_47#_c_774_n 0.0133285f $X=3.965 $Y=1.565 $X2=0 $Y2=0
cc_273 N_A1_M1000_g N_A_684_47#_c_776_n 0.00191791f $X=3.345 $Y=0.655 $X2=0
+ $Y2=0
cc_274 N_A1_c_277_n N_A_684_47#_c_776_n 0.00449783f $X=3.64 $Y=1.51 $X2=0 $Y2=0
cc_275 N_A1_c_278_n N_A_684_47#_c_776_n 0.0183892f $X=3.965 $Y=1.565 $X2=0 $Y2=0
cc_276 N_A2_c_349_n N_Y_c_509_n 4.25868e-19 $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A2_M1006_g N_Y_c_469_n 0.010446f $X=4.07 $Y=2.465 $X2=0 $Y2=0
cc_278 N_A2_M1018_g N_Y_c_469_n 0.0106163f $X=4.5 $Y=2.465 $X2=0 $Y2=0
cc_279 A2 N_Y_c_464_n 0.00467638f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_280 N_A2_c_356_n N_Y_c_466_n 2.01187e-19 $X=4.52 $Y=1.185 $X2=0 $Y2=0
cc_281 N_A2_c_349_n Y 7.89594e-19 $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_282 N_A2_c_353_n Y 4.24706e-19 $X=4.057 $Y=1.26 $X2=0 $Y2=0
cc_283 N_A2_M1006_g N_A_467_367#_c_598_n 0.0122129f $X=4.07 $Y=2.465 $X2=0 $Y2=0
cc_284 N_A2_M1018_g N_A_467_367#_c_599_n 0.0129951f $X=4.5 $Y=2.465 $X2=0 $Y2=0
cc_285 N_A2_M1006_g N_VPWR_c_636_n 0.0104312f $X=4.07 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A2_M1018_g N_VPWR_c_636_n 5.82565e-19 $X=4.5 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A2_M1006_g N_VPWR_c_637_n 5.54009e-19 $X=4.07 $Y=2.465 $X2=0 $Y2=0
cc_288 N_A2_M1018_g N_VPWR_c_637_n 0.00920327f $X=4.5 $Y=2.465 $X2=0 $Y2=0
cc_289 N_A2_M1006_g N_VPWR_c_640_n 0.00486043f $X=4.07 $Y=2.465 $X2=0 $Y2=0
cc_290 N_A2_M1018_g N_VPWR_c_640_n 0.00564095f $X=4.5 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A2_M1006_g N_VPWR_c_635_n 0.00824727f $X=4.07 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A2_M1018_g N_VPWR_c_635_n 0.00948291f $X=4.5 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A2_c_349_n N_VGND_c_705_n 0.00411639f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_294 N_A2_c_356_n N_VGND_c_705_n 0.00407566f $X=4.52 $Y=1.185 $X2=0 $Y2=0
cc_295 N_A2_c_349_n N_VGND_c_706_n 0.00585385f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_296 N_A2_c_356_n N_VGND_c_711_n 0.00585385f $X=4.52 $Y=1.185 $X2=0 $Y2=0
cc_297 N_A2_c_349_n N_VGND_c_712_n 0.0114812f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_298 N_A2_c_356_n N_VGND_c_712_n 0.010827f $X=4.52 $Y=1.185 $X2=0 $Y2=0
cc_299 N_A2_c_349_n N_A_684_47#_c_773_n 0.00964758f $X=4.045 $Y=1.185 $X2=0
+ $Y2=0
cc_300 N_A2_c_349_n N_A_684_47#_c_774_n 0.0169846f $X=4.045 $Y=1.185 $X2=0 $Y2=0
cc_301 N_A2_c_351_n N_A_684_47#_c_774_n 0.00392667f $X=4.355 $Y=1.26 $X2=0 $Y2=0
cc_302 A2 N_A_684_47#_c_774_n 0.022584f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_303 N_A2_c_355_n N_A_684_47#_c_774_n 0.00128968f $X=4.52 $Y=1.26 $X2=0 $Y2=0
cc_304 N_A2_c_356_n N_A_684_47#_c_774_n 0.0133548f $X=4.52 $Y=1.185 $X2=0 $Y2=0
cc_305 N_A_32_367#_c_413_n N_A_115_367#_M1005_s 0.00334517f $X=1.87 $Y=2.97
+ $X2=-0.19 $Y2=1.655
cc_306 N_A_32_367#_c_413_n N_A_115_367#_M1016_d 0.00334517f $X=1.87 $Y=2.97
+ $X2=0 $Y2=0
cc_307 N_A_32_367#_c_413_n N_A_115_367#_c_447_n 0.0312112f $X=1.87 $Y=2.97 $X2=0
+ $Y2=0
cc_308 N_A_32_367#_c_413_n N_A_115_367#_c_446_n 0.0132625f $X=1.87 $Y=2.97 $X2=0
+ $Y2=0
cc_309 N_A_32_367#_c_413_n N_A_115_367#_c_453_n 0.0124294f $X=1.87 $Y=2.97 $X2=0
+ $Y2=0
cc_310 N_A_32_367#_c_413_n N_Y_M1009_s 0.0033495f $X=1.87 $Y=2.97 $X2=0 $Y2=0
cc_311 N_A_32_367#_M1008_d N_Y_c_479_n 0.00702272f $X=1.865 $Y=1.835 $X2=0 $Y2=0
cc_312 N_A_32_367#_M1010_s N_Y_c_479_n 0.00623139f $X=2.765 $Y=1.835 $X2=0 $Y2=0
cc_313 N_A_32_367#_c_427_p N_Y_c_479_n 0.0168246f $X=2.005 $Y=2.46 $X2=0 $Y2=0
cc_314 N_A_32_367#_M1010_s Y 0.00145169f $X=2.765 $Y=1.835 $X2=0 $Y2=0
cc_315 N_A_32_367#_c_410_n N_A_467_367#_M1001_d 0.0033716f $X=2.905 $Y=2.93
+ $X2=-0.19 $Y2=1.655
cc_316 N_A_32_367#_M1010_s N_A_467_367#_c_591_n 0.00585539f $X=2.765 $Y=1.835
+ $X2=0 $Y2=0
cc_317 N_A_32_367#_c_410_n N_A_467_367#_c_591_n 0.0419588f $X=2.905 $Y=2.93
+ $X2=0 $Y2=0
cc_318 N_A_32_367#_c_410_n N_A_467_367#_c_592_n 0.0207418f $X=2.905 $Y=2.93
+ $X2=0 $Y2=0
cc_319 N_A_32_367#_c_408_n N_VPWR_c_638_n 0.0186279f $X=0.26 $Y=2.865 $X2=0
+ $Y2=0
cc_320 N_A_32_367#_c_413_n N_VPWR_c_638_n 0.0824808f $X=1.87 $Y=2.97 $X2=0 $Y2=0
cc_321 N_A_32_367#_c_410_n N_VPWR_c_638_n 0.0527154f $X=2.905 $Y=2.93 $X2=0
+ $Y2=0
cc_322 N_A_32_367#_c_436_p N_VPWR_c_638_n 0.0176422f $X=2.005 $Y=2.91 $X2=0
+ $Y2=0
cc_323 N_A_32_367#_M1005_d N_VPWR_c_635_n 0.0021516f $X=0.16 $Y=1.835 $X2=0
+ $Y2=0
cc_324 N_A_32_367#_M1008_d N_VPWR_c_635_n 0.0025251f $X=1.865 $Y=1.835 $X2=0
+ $Y2=0
cc_325 N_A_32_367#_M1010_s N_VPWR_c_635_n 0.00215176f $X=2.765 $Y=1.835 $X2=0
+ $Y2=0
cc_326 N_A_32_367#_c_408_n N_VPWR_c_635_n 0.0108858f $X=0.26 $Y=2.865 $X2=0
+ $Y2=0
cc_327 N_A_32_367#_c_413_n N_VPWR_c_635_n 0.0526325f $X=1.87 $Y=2.97 $X2=0 $Y2=0
cc_328 N_A_32_367#_c_410_n N_VPWR_c_635_n 0.0328282f $X=2.905 $Y=2.93 $X2=0
+ $Y2=0
cc_329 N_A_32_367#_c_436_p N_VPWR_c_635_n 0.0114689f $X=2.005 $Y=2.91 $X2=0
+ $Y2=0
cc_330 N_A_115_367#_c_447_n N_Y_M1009_s 0.00346461f $X=1.45 $Y=2.61 $X2=0.5
+ $Y2=2.465
cc_331 N_A_115_367#_M1016_d N_Y_c_479_n 0.00350245f $X=1.435 $Y=1.835 $X2=0.5
+ $Y2=1.46
cc_332 N_A_115_367#_c_447_n N_Y_c_479_n 0.00509093f $X=1.45 $Y=2.61 $X2=0.5
+ $Y2=1.46
cc_333 N_A_115_367#_c_453_n N_Y_c_479_n 0.0129938f $X=1.575 $Y=2.46 $X2=0.5
+ $Y2=1.46
cc_334 N_A_115_367#_c_447_n N_Y_c_488_n 0.0132201f $X=1.45 $Y=2.61 $X2=0 $Y2=0
cc_335 N_A_115_367#_M1005_s N_VPWR_c_635_n 0.00225186f $X=0.575 $Y=1.835
+ $X2=1.81 $Y2=1.625
cc_336 N_A_115_367#_M1016_d N_VPWR_c_635_n 0.00224381f $X=1.435 $Y=1.835
+ $X2=1.81 $Y2=1.625
cc_337 N_Y_c_479_n N_A_467_367#_M1001_d 0.00334717f $X=3.025 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_338 N_Y_c_469_n N_A_467_367#_M1002_s 0.00546176f $X=5.325 $Y=2.04 $X2=0 $Y2=0
cc_339 N_Y_c_469_n N_A_467_367#_M1006_d 0.00337418f $X=5.325 $Y=2.04 $X2=0 $Y2=0
cc_340 N_Y_c_469_n N_A_467_367#_M1014_s 0.00759464f $X=5.325 $Y=2.04 $X2=0 $Y2=0
cc_341 N_Y_c_479_n N_A_467_367#_c_591_n 0.0391788f $X=3.025 $Y=2.035 $X2=0 $Y2=0
cc_342 Y N_A_467_367#_c_591_n 0.0207726f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_343 N_Y_c_469_n N_A_467_367#_c_598_n 0.0323235f $X=5.325 $Y=2.04 $X2=0 $Y2=0
cc_344 N_Y_c_469_n N_A_467_367#_c_599_n 0.035161f $X=5.325 $Y=2.04 $X2=0 $Y2=0
cc_345 N_Y_c_469_n N_A_467_367#_c_593_n 0.0204473f $X=5.325 $Y=2.04 $X2=0 $Y2=0
cc_346 N_Y_c_469_n N_A_467_367#_c_595_n 0.0173071f $X=5.325 $Y=2.04 $X2=0 $Y2=0
cc_347 Y N_A_467_367#_c_595_n 0.00327941f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_348 N_Y_c_469_n N_A_467_367#_c_618_n 0.0135055f $X=5.325 $Y=2.04 $X2=0 $Y2=0
cc_349 N_Y_c_469_n N_VPWR_M1002_d 0.00353783f $X=5.325 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_350 N_Y_c_469_n N_VPWR_M1018_s 0.0043175f $X=5.325 $Y=2.04 $X2=0 $Y2=0
cc_351 N_Y_M1009_s N_VPWR_c_635_n 0.00225186f $X=1.005 $Y=1.835 $X2=0 $Y2=0
cc_352 N_Y_c_473_n N_VGND_M1012_s 0.00353353f $X=1.05 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_353 N_Y_c_483_n N_VGND_M1015_d 0.0066154f $X=1.965 $Y=0.955 $X2=0 $Y2=0
cc_354 N_Y_c_473_n N_VGND_c_702_n 0.0170777f $X=1.05 $Y=0.955 $X2=0 $Y2=0
cc_355 N_Y_c_483_n N_VGND_c_703_n 0.022455f $X=1.965 $Y=0.955 $X2=0 $Y2=0
cc_356 N_Y_c_463_n N_VGND_c_704_n 0.0247883f $X=2.965 $Y=1.17 $X2=0 $Y2=0
cc_357 N_Y_c_509_n N_VGND_c_706_n 0.0189236f $X=3.13 $Y=0.375 $X2=0 $Y2=0
cc_358 N_Y_c_461_n N_VGND_c_708_n 0.0178111f $X=0.285 $Y=0.43 $X2=0 $Y2=0
cc_359 N_Y_c_478_n N_VGND_c_709_n 0.01379f $X=1.145 $Y=0.43 $X2=0 $Y2=0
cc_360 N_Y_c_487_n N_VGND_c_710_n 0.0192488f $X=2.145 $Y=0.42 $X2=0 $Y2=0
cc_361 N_Y_c_466_n N_VGND_c_711_n 0.0432696f $X=5.185 $Y=0.42 $X2=0 $Y2=0
cc_362 N_Y_M1012_d N_VGND_c_712_n 0.00371702f $X=0.16 $Y=0.235 $X2=0 $Y2=0
cc_363 N_Y_M1007_s N_VGND_c_712_n 0.00380321f $X=1.005 $Y=0.235 $X2=0 $Y2=0
cc_364 N_Y_M1017_d N_VGND_c_712_n 0.0027714f $X=1.975 $Y=0.235 $X2=0 $Y2=0
cc_365 N_Y_M1011_s N_VGND_c_712_n 0.00223559f $X=2.99 $Y=0.235 $X2=0 $Y2=0
cc_366 N_Y_M1013_s N_VGND_c_712_n 0.00215158f $X=5.045 $Y=0.235 $X2=0 $Y2=0
cc_367 N_Y_c_461_n N_VGND_c_712_n 0.0100304f $X=0.285 $Y=0.43 $X2=0 $Y2=0
cc_368 N_Y_c_478_n N_VGND_c_712_n 0.0092882f $X=1.145 $Y=0.43 $X2=0 $Y2=0
cc_369 N_Y_c_487_n N_VGND_c_712_n 0.0126375f $X=2.145 $Y=0.42 $X2=0 $Y2=0
cc_370 N_Y_c_509_n N_VGND_c_712_n 0.0123859f $X=3.13 $Y=0.375 $X2=0 $Y2=0
cc_371 N_Y_c_466_n N_VGND_c_712_n 0.024621f $X=5.185 $Y=0.42 $X2=0 $Y2=0
cc_372 N_Y_c_509_n N_A_684_47#_c_773_n 0.037202f $X=3.13 $Y=0.375 $X2=0 $Y2=0
cc_373 N_Y_c_509_n N_A_684_47#_c_776_n 0.0109407f $X=3.13 $Y=0.375 $X2=0 $Y2=0
cc_374 N_A_467_367#_c_598_n N_VPWR_M1002_d 0.00353353f $X=4.19 $Y=2.38 $X2=-0.19
+ $Y2=1.655
cc_375 N_A_467_367#_c_599_n N_VPWR_M1018_s 0.00438498f $X=5.07 $Y=2.38 $X2=0
+ $Y2=0
cc_376 N_A_467_367#_c_598_n N_VPWR_c_636_n 0.0170777f $X=4.19 $Y=2.38 $X2=0
+ $Y2=0
cc_377 N_A_467_367#_c_599_n N_VPWR_c_637_n 0.017251f $X=5.07 $Y=2.38 $X2=0 $Y2=0
cc_378 N_A_467_367#_c_591_n N_VPWR_c_638_n 0.00328876f $X=3.26 $Y=2.47 $X2=0
+ $Y2=0
cc_379 N_A_467_367#_c_592_n N_VPWR_c_638_n 0.0178111f $X=3.425 $Y=2.91 $X2=0
+ $Y2=0
cc_380 N_A_467_367#_c_625_p N_VPWR_c_640_n 0.0131621f $X=4.285 $Y=2.91 $X2=0
+ $Y2=0
cc_381 N_A_467_367#_c_594_n N_VPWR_c_642_n 0.0185207f $X=5.185 $Y=2.91 $X2=0
+ $Y2=0
cc_382 N_A_467_367#_M1001_d N_VPWR_c_635_n 0.00225186f $X=2.335 $Y=1.835 $X2=0
+ $Y2=0
cc_383 N_A_467_367#_M1002_s N_VPWR_c_635_n 0.00371702f $X=3.3 $Y=1.835 $X2=0
+ $Y2=0
cc_384 N_A_467_367#_M1006_d N_VPWR_c_635_n 0.00467071f $X=4.145 $Y=1.835 $X2=0
+ $Y2=0
cc_385 N_A_467_367#_M1014_s N_VPWR_c_635_n 0.00302127f $X=5.045 $Y=1.835 $X2=0
+ $Y2=0
cc_386 N_A_467_367#_c_591_n N_VPWR_c_635_n 0.00684347f $X=3.26 $Y=2.47 $X2=0
+ $Y2=0
cc_387 N_A_467_367#_c_592_n N_VPWR_c_635_n 0.0100304f $X=3.425 $Y=2.91 $X2=0
+ $Y2=0
cc_388 N_A_467_367#_c_625_p N_VPWR_c_635_n 0.00808656f $X=4.285 $Y=2.91 $X2=0
+ $Y2=0
cc_389 N_A_467_367#_c_594_n N_VPWR_c_635_n 0.010808f $X=5.185 $Y=2.91 $X2=0
+ $Y2=0
cc_390 N_VGND_c_712_n N_A_684_47#_M1000_d 0.0122096f $X=5.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_391 N_VGND_c_712_n N_A_684_47#_M1019_d 0.0041489f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_706_n N_A_684_47#_c_773_n 0.0230625f $X=4.125 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_712_n N_A_684_47#_c_773_n 0.0127519f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_394 N_VGND_M1004_s N_A_684_47#_c_774_n 0.00557461f $X=4.12 $Y=0.235 $X2=0
+ $Y2=0
cc_395 N_VGND_c_705_n N_A_684_47#_c_774_n 0.0187938f $X=4.29 $Y=0.575 $X2=0
+ $Y2=0
cc_396 N_VGND_c_711_n N_A_684_47#_c_793_n 0.0136943f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_c_712_n N_A_684_47#_c_793_n 0.00866972f $X=5.52 $Y=0 $X2=0 $Y2=0
