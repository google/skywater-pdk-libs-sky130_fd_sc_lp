# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.150000 1.295000 1.395000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.145000 1.845000 10.475000 3.075000 ;
        RECT 10.155000 0.255000 10.475000 1.090000 ;
        RECT 10.205000 1.090000 10.475000 1.845000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.565000 0.680000 2.120000 ;
        RECT 2.555000 1.565000 3.375000 1.750000 ;
        RECT 6.855000 1.580000 7.295000 1.835000 ;
        RECT 7.045000 1.835000 7.295000 2.250000 ;
      LAYER mcon ;
        RECT 0.155000 1.580000 0.325000 1.750000 ;
        RECT 2.555000 1.580000 2.725000 1.750000 ;
        RECT 6.875000 1.580000 7.045000 1.750000 ;
      LAYER met1 ;
        RECT 0.095000 1.550000 0.385000 1.595000 ;
        RECT 0.095000 1.595000 7.105000 1.735000 ;
        RECT 0.095000 1.735000 0.385000 1.780000 ;
        RECT 2.495000 1.550000 2.785000 1.595000 ;
        RECT 2.495000 1.735000 2.785000 1.780000 ;
        RECT 6.815000 1.550000 7.105000 1.595000 ;
        RECT 6.815000 1.735000 7.105000 1.780000 ;
    END
  END RESET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.570000 8.505000 2.215000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.560000 0.085000 ;
        RECT 0.255000  0.085000  0.585000 0.980000 ;
        RECT 3.250000  0.085000  3.580000 0.540000 ;
        RECT 4.470000  0.085000  4.800000 0.415000 ;
        RECT 6.790000  0.085000  7.120000 0.710000 ;
        RECT 8.760000  0.085000  8.930000 0.890000 ;
        RECT 8.760000  0.890000  9.215000 1.060000 ;
        RECT 9.015000  1.060000  9.215000 1.320000 ;
        RECT 9.725000  0.085000  9.985000 1.090000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 10.560000 3.415000 ;
        RECT 0.640000 2.630000  0.970000 3.245000 ;
        RECT 2.830000 2.610000  3.160000 3.245000 ;
        RECT 4.525000 2.965000  4.855000 3.245000 ;
        RECT 6.720000 2.785000  6.920000 3.245000 ;
        RECT 8.145000 2.745000  8.335000 3.245000 ;
        RECT 9.605000 1.845000  9.975000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.100000 2.290000  1.565000 2.460000 ;
      RECT 0.100000 2.460000  0.470000 2.735000 ;
      RECT 1.150000 0.650000  1.635000 0.980000 ;
      RECT 1.160000 1.565000  1.635000 1.820000 ;
      RECT 1.160000 1.820000  1.565000 2.290000 ;
      RECT 1.160000 2.460000  1.565000 2.735000 ;
      RECT 1.465000 0.980000  1.635000 1.565000 ;
      RECT 1.470000 0.255000  2.335000 0.480000 ;
      RECT 1.735000 2.085000  1.985000 2.270000 ;
      RECT 1.735000 2.270000  4.845000 2.440000 ;
      RECT 1.735000 2.440000  2.040000 2.735000 ;
      RECT 1.805000 0.675000  1.985000 2.085000 ;
      RECT 2.155000 0.480000  2.335000 0.710000 ;
      RECT 2.155000 0.710000  5.140000 0.765000 ;
      RECT 2.155000 0.765000  4.165000 0.880000 ;
      RECT 2.155000 0.880000  2.335000 1.920000 ;
      RECT 2.155000 1.920000  4.275000 2.100000 ;
      RECT 2.505000 1.050000  5.480000 1.105000 ;
      RECT 2.505000 1.105000  4.505000 1.220000 ;
      RECT 2.505000 1.220000  2.835000 1.395000 ;
      RECT 3.330000 2.440000  3.645000 2.735000 ;
      RECT 3.915000 0.550000  4.245000 0.585000 ;
      RECT 3.915000 0.585000  5.140000 0.710000 ;
      RECT 4.025000 2.625000  5.370000 2.765000 ;
      RECT 4.025000 2.765000  6.245000 2.795000 ;
      RECT 4.025000 2.795000  4.355000 3.065000 ;
      RECT 4.335000 0.935000  5.480000 1.050000 ;
      RECT 4.675000 1.275000  4.845000 2.270000 ;
      RECT 4.970000 0.255000  6.375000 0.425000 ;
      RECT 4.970000 0.425000  5.140000 0.585000 ;
      RECT 5.025000 1.105000  5.480000 1.205000 ;
      RECT 5.025000 1.205000  5.205000 2.245000 ;
      RECT 5.025000 2.245000  5.370000 2.455000 ;
      RECT 5.200000 2.795000  6.245000 2.935000 ;
      RECT 5.310000 0.595000  5.480000 0.935000 ;
      RECT 5.385000 1.480000  5.830000 1.735000 ;
      RECT 5.385000 1.735000  5.555000 1.810000 ;
      RECT 5.540000 1.980000  6.170000 2.075000 ;
      RECT 5.540000 2.075000  5.830000 2.100000 ;
      RECT 5.540000 2.100000  5.800000 2.115000 ;
      RECT 5.540000 2.115000  5.770000 2.155000 ;
      RECT 5.540000 2.155000  5.720000 2.585000 ;
      RECT 5.610000 1.975000  6.170000 1.980000 ;
      RECT 5.625000 1.965000  6.170000 1.975000 ;
      RECT 5.640000 1.960000  6.170000 1.965000 ;
      RECT 5.655000 1.950000  6.170000 1.960000 ;
      RECT 5.660000 0.425000  6.375000 0.435000 ;
      RECT 5.660000 0.435000  5.830000 1.480000 ;
      RECT 5.680000 1.935000  6.170000 1.950000 ;
      RECT 5.700000 1.905000  6.170000 1.935000 ;
      RECT 5.920000 2.245000  6.250000 2.430000 ;
      RECT 5.920000 2.430000  7.260000 2.600000 ;
      RECT 5.920000 2.600000  6.245000 2.765000 ;
      RECT 6.000000 0.605000  6.225000 0.880000 ;
      RECT 6.000000 0.880000  7.490000 1.060000 ;
      RECT 6.000000 1.060000  6.170000 1.905000 ;
      RECT 6.515000 1.230000  7.990000 1.400000 ;
      RECT 6.515000 1.400000  6.685000 2.050000 ;
      RECT 7.090000 2.600000  7.260000 2.895000 ;
      RECT 7.090000 2.895000  7.975000 3.065000 ;
      RECT 7.310000 0.265000  8.360000 0.490000 ;
      RECT 7.310000 0.490000  7.490000 0.880000 ;
      RECT 7.465000 1.400000  7.635000 2.725000 ;
      RECT 7.660000 0.660000  7.990000 1.230000 ;
      RECT 7.805000 2.405000  8.845000 2.575000 ;
      RECT 7.805000 2.575000  7.975000 2.895000 ;
      RECT 8.215000 0.940000  8.475000 1.230000 ;
      RECT 8.215000 1.230000  8.845000 1.400000 ;
      RECT 8.505000 2.575000  8.845000 3.075000 ;
      RECT 8.675000 1.400000  8.845000 2.405000 ;
      RECT 9.120000 1.505000 10.035000 1.675000 ;
      RECT 9.120000 1.675000  9.435000 2.495000 ;
      RECT 9.180000 0.280000  9.555000 0.610000 ;
      RECT 9.385000 0.610000  9.555000 1.345000 ;
      RECT 9.385000 1.345000 10.035000 1.505000 ;
  END
END sky130_fd_sc_lp__dfrtn_1
