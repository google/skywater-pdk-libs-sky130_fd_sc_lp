* File: sky130_fd_sc_lp__o41a_0.pex.spice
* Created: Fri Aug 28 11:19:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41A_0%A_80_21# 1 2 9 11 14 16 20 21 22 23 24 25 28
+ 31 35 38
r73 32 35 8.93541 $w=6.78e-07 $l=5.08e-07 $layer=LI1_cond $X=1.317 $Y=2.735
+ $X2=1.825 $Y2=2.735
r74 31 32 7.62417 $w=2.15e-07 $l=3.4e-07 $layer=LI1_cond $X=1.317 $Y=2.395
+ $X2=1.317 $Y2=2.735
r75 30 31 9.64836 $w=2.13e-07 $l=1.8e-07 $layer=LI1_cond $X=1.317 $Y=2.215
+ $X2=1.317 $Y2=2.395
r76 26 28 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=1.29 $Y=0.74
+ $X2=1.29 $Y2=0.465
r77 24 30 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=1.21 $Y=2.13
+ $X2=1.317 $Y2=2.215
r78 24 25 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.21 $Y=2.13
+ $X2=0.775 $Y2=2.13
r79 22 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.14 $Y=0.825
+ $X2=1.29 $Y2=0.74
r80 22 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.14 $Y=0.825
+ $X2=0.775 $Y2=0.825
r81 21 38 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=0.93
+ $X2=0.587 $Y2=0.765
r82 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=0.93 $X2=0.61 $Y2=0.93
r83 18 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.65 $Y=2.045
+ $X2=0.775 $Y2=2.13
r84 18 20 51.399 $w=2.48e-07 $l=1.115e-06 $layer=LI1_cond $X=0.65 $Y=2.045
+ $X2=0.65 $Y2=0.93
r85 17 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.65 $Y=0.91
+ $X2=0.775 $Y2=0.825
r86 17 20 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=0.65 $Y=0.91 $X2=0.65
+ $Y2=0.93
r87 14 16 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=0.66 $Y=2.735
+ $X2=0.66 $Y2=1.435
r88 11 16 43.0937 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.587 $Y=1.248
+ $X2=0.587 $Y2=1.435
r89 10 21 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.587 $Y=0.952
+ $X2=0.587 $Y2=0.93
r90 10 11 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.587 $Y=0.952
+ $X2=0.587 $Y2=1.248
r91 9 38 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.765
r92 2 35 150 $w=1.7e-07 $l=7.28903e-07 $layer=licon1_PDIFF $count=4 $X=1.165
+ $Y=2.415 $X2=1.825 $Y2=2.56
r93 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.18
+ $Y=0.255 $X2=1.305 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_0%B1 3 7 12 15 16 17 21
r47 16 17 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.18 $Y=1.245
+ $X2=1.18 $Y2=1.665
r48 16 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.18
+ $Y=1.245 $X2=1.18 $Y2=1.245
r49 14 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.18 $Y=1.585
+ $X2=1.18 $Y2=1.245
r50 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.585
+ $X2=1.18 $Y2=1.75
r51 10 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.18 $Y=1.23
+ $X2=1.18 $Y2=1.245
r52 10 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.18 $Y=1.155
+ $X2=1.52 $Y2=1.155
r53 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.52 $Y=1.08 $X2=1.52
+ $Y2=1.155
r54 5 7 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.52 $Y=1.08 $X2=1.52
+ $Y2=0.465
r55 3 15 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=1.09 $Y=2.735
+ $X2=1.09 $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_0%A4 1 3 7 10 11 12 13 14
c50 12 0 3.31551e-20 $X=1.68 $Y=1.295
c51 3 0 1.26066e-19 $X=1.95 $Y=0.465
r52 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.95
+ $Y=1.635 $X2=1.95 $Y2=1.635
r53 13 14 6.91483 $w=6.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.915 $Y=1.665
+ $X2=1.915 $Y2=2.035
r54 13 20 0.560662 $w=6.38e-07 $l=3e-08 $layer=LI1_cond $X=1.915 $Y=1.665
+ $X2=1.915 $Y2=1.635
r55 12 20 6.35417 $w=6.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.915 $Y=1.295
+ $X2=1.915 $Y2=1.635
r56 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.95 $Y=1.975
+ $X2=1.95 $Y2=1.635
r57 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.95 $Y=1.975
+ $X2=1.95 $Y2=2.14
r58 7 11 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=2.04 $Y=2.735
+ $X2=2.04 $Y2=2.14
r59 1 19 87.7993 $w=2.69e-07 $l=4.9e-07 $layer=POLY_cond $X=1.95 $Y=1.145
+ $X2=1.95 $Y2=1.635
r60 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.95 $Y=1.145 $X2=1.95
+ $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_0%A3 3 5 7 11 12 13 14 15 16 24 41
c54 24 0 2.95765e-20 $X=2.49 $Y=1.7
c55 12 0 1.26066e-19 $X=2.64 $Y=1.295
c56 7 0 3.31551e-20 $X=2.49 $Y=2.735
r57 26 41 0.467207 $w=3.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.59 $Y=2.02
+ $X2=2.59 $Y2=2.035
r58 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.49 $Y=1.7
+ $X2=2.49 $Y2=1.7
r59 15 16 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.405
+ $X2=2.62 $Y2=2.775
r60 15 43 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=2.62 $Y=2.405 $X2=2.62
+ $Y2=2.205
r61 14 43 4.54172 $w=3.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.59 $Y=2.07
+ $X2=2.59 $Y2=2.205
r62 14 41 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.59 $Y=2.07
+ $X2=2.59 $Y2=2.035
r63 14 26 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.59 $Y=1.985
+ $X2=2.59 $Y2=2.02
r64 14 25 8.87693 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.59 $Y=1.985
+ $X2=2.59 $Y2=1.7
r65 13 25 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.59 $Y=1.665
+ $X2=2.59 $Y2=1.7
r66 12 13 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.59 $Y=1.295
+ $X2=2.59 $Y2=1.665
r67 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.49 $Y=2.04
+ $X2=2.49 $Y2=1.7
r68 10 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=1.535
+ $X2=2.49 $Y2=1.7
r69 5 11 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.49 $Y=2.205
+ $X2=2.49 $Y2=2.04
r70 5 7 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.49 $Y=2.205 $X2=2.49
+ $Y2=2.735
r71 3 10 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.4 $Y=0.465 $X2=2.4
+ $Y2=1.535
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_0%A2 1 3 8 12 15 16 17 18 19 20 21 22 29
r56 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.03
+ $Y=1.41 $X2=3.03 $Y2=1.41
r57 21 22 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.075 $Y=2.405
+ $X2=3.075 $Y2=2.775
r58 20 21 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=3.075 $Y2=2.405
r59 19 20 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.075 $Y=1.665
+ $X2=3.075 $Y2=2.035
r60 19 30 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=3.075 $Y=1.665
+ $X2=3.075 $Y2=1.41
r61 18 30 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=3.075 $Y=1.295
+ $X2=3.075 $Y2=1.41
r62 16 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.03 $Y=1.75
+ $X2=3.03 $Y2=1.41
r63 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.03 $Y=1.75
+ $X2=3.03 $Y2=1.915
r64 15 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.03 $Y=1.245
+ $X2=3.03 $Y2=1.41
r65 10 12 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=2.83 $Y=0.86
+ $X2=2.94 $Y2=0.86
r66 8 17 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.94 $Y=2.735
+ $X2=2.94 $Y2=1.915
r67 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.94 $Y=0.935
+ $X2=2.94 $Y2=0.86
r68 4 15 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=2.94 $Y=0.935
+ $X2=2.94 $Y2=1.245
r69 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.83 $Y=0.785
+ $X2=2.83 $Y2=0.86
r70 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.83 $Y=0.785 $X2=2.83
+ $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_0%A1 3 5 7 9 13 17 20 21 22 23 28 29
r38 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.12 $X2=3.57 $Y2=1.12
r39 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=2.035
r40 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.295
+ $X2=3.57 $Y2=1.665
r41 21 29 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=3.57 $Y=1.295
+ $X2=3.57 $Y2=1.12
r42 19 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.57 $Y=1.46
+ $X2=3.57 $Y2=1.12
r43 19 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.57 $Y=1.46
+ $X2=3.57 $Y2=1.625
r44 15 17 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.3 $Y=2.23 $X2=3.48
+ $Y2=2.23
r45 13 28 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.57 $Y=1.005
+ $X2=3.57 $Y2=1.12
r46 10 13 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.3 $Y=0.93 $X2=3.57
+ $Y2=0.93
r47 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.48 $Y=2.155
+ $X2=3.48 $Y2=2.23
r48 9 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.48 $Y=2.155
+ $X2=3.48 $Y2=1.625
r49 5 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.3 $Y=2.305 $X2=3.3
+ $Y2=2.23
r50 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.3 $Y=2.305 $X2=3.3
+ $Y2=2.735
r51 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.3 $Y=0.855 $X2=3.3
+ $Y2=0.93
r52 1 3 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.3 $Y=0.855 $X2=3.3
+ $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_0%X 1 2 7 8 9 10 11 12 13 24 38
r16 38 39 2.22423 $w=4.53e-07 $l=1e-08 $layer=LI1_cond $X=0.312 $Y=2.405
+ $X2=0.312 $Y2=2.395
r17 13 42 5.6518 $w=4.53e-07 $l=2.15e-07 $layer=LI1_cond $X=0.312 $Y=2.775
+ $X2=0.312 $Y2=2.56
r18 12 42 3.10192 $w=4.53e-07 $l=1.18e-07 $layer=LI1_cond $X=0.312 $Y=2.442
+ $X2=0.312 $Y2=2.56
r19 12 38 0.972635 $w=4.53e-07 $l=3.7e-08 $layer=LI1_cond $X=0.312 $Y=2.442
+ $X2=0.312 $Y2=2.405
r20 12 39 1.62196 $w=2.68e-07 $l=3.8e-08 $layer=LI1_cond $X=0.22 $Y=2.357
+ $X2=0.22 $Y2=2.395
r21 11 12 13.7439 $w=2.68e-07 $l=3.22e-07 $layer=LI1_cond $X=0.22 $Y=2.035
+ $X2=0.22 $Y2=2.357
r22 10 11 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=2.035
r23 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.665
r24 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.925 $X2=0.22
+ $Y2=1.295
r25 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.555 $X2=0.22
+ $Y2=0.925
r26 7 24 4.90855 $w=2.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.22 $Y=0.555
+ $X2=0.22 $Y2=0.44
r27 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.32
+ $Y=2.415 $X2=0.445 $Y2=2.56
r28 1 24 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_0%VPWR 1 2 11 13 15 17 19 28 32
r37 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r38 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r40 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 20 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=0.875 $Y2=3.33
r45 20 22 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.04 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 19 31 4.52193 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.607 $Y2=3.33
r47 19 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 17 26 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 17 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 13 31 3.11857 $w=3.15e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.532 $Y=3.245
+ $X2=3.607 $Y2=3.33
r51 13 15 25.0611 $w=3.13e-07 $l=6.85e-07 $layer=LI1_cond $X=3.532 $Y=3.245
+ $X2=3.532 $Y2=2.56
r52 9 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=3.33
r53 9 11 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=2.56
r54 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.375
+ $Y=2.415 $X2=3.515 $Y2=2.56
r55 1 11 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.735
+ $Y=2.415 $X2=0.875 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_0%VGND 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
r56 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r58 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r59 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r60 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r61 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=0 $X2=3.065
+ $Y2=0
r62 39 41 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.23 $Y=0 $X2=3.6
+ $Y2=0
r63 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r64 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r65 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r66 35 48 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.175
+ $Y2=0
r67 35 37 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.64
+ $Y2=0
r68 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=3.065
+ $Y2=0
r69 34 37 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=0 $X2=2.64
+ $Y2=0
r70 33 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r71 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r72 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r73 30 32 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.68
+ $Y2=0
r74 29 48 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.175
+ $Y2=0
r75 29 32 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.68
+ $Y2=0
r76 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r77 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r78 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r79 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r80 22 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r81 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r82 18 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.065 $Y2=0
r83 18 20 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.065 $Y=0.085
+ $X2=3.065 $Y2=0.415
r84 14 48 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0
r85 14 16 15.6403 $w=2.78e-07 $l=3.8e-07 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0.465
r86 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r87 10 12 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.445
r88 3 20 182 $w=1.7e-07 $l=2.26274e-07 $layer=licon1_NDIFF $count=1 $X=2.905
+ $Y=0.255 $X2=3.065 $Y2=0.415
r89 2 16 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.255 $X2=2.18 $Y2=0.465
r90 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_0%A_319_51# 1 2 3 12 14 15 18 20 24 26
c48 14 0 2.95765e-20 $X=2.485 $Y=0.885
r49 22 24 8.69055 $w=3.03e-07 $l=2.3e-07 $layer=LI1_cond $X=3.552 $Y=0.695
+ $X2=3.552 $Y2=0.465
r50 21 26 6.92067 $w=1.7e-07 $l=2.84341e-07 $layer=LI1_cond $X=2.73 $Y=0.78
+ $X2=2.485 $Y2=0.695
r51 20 22 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=3.4 $Y=0.78
+ $X2=3.552 $Y2=0.695
r52 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.4 $Y=0.78 $X2=2.73
+ $Y2=0.78
r53 16 26 0.066131 $w=2.45e-07 $l=1.22e-07 $layer=LI1_cond $X=2.607 $Y=0.695
+ $X2=2.485 $Y2=0.695
r54 16 18 10.8189 $w=2.43e-07 $l=2.3e-07 $layer=LI1_cond $X=2.607 $Y=0.695
+ $X2=2.607 $Y2=0.465
r55 14 26 6.92067 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.485 $Y=0.885
+ $X2=2.485 $Y2=0.695
r56 14 15 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.485 $Y=0.885
+ $X2=1.865 $Y2=0.885
r57 10 15 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=1.737 $Y=0.8
+ $X2=1.865 $Y2=0.885
r58 10 12 15.1399 $w=2.53e-07 $l=3.35e-07 $layer=LI1_cond $X=1.737 $Y=0.8
+ $X2=1.737 $Y2=0.465
r59 3 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.255 $X2=3.515 $Y2=0.465
r60 2 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.255 $X2=2.615 $Y2=0.465
r61 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.255 $X2=1.735 $Y2=0.465
.ends

