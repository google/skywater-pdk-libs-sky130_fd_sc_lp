* File: sky130_fd_sc_lp__dlrtn_1.spice
* Created: Wed Sep  2 09:46:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrtn_1.pex.spice"
.subckt sky130_fd_sc_lp__dlrtn_1  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_D_M1018_g N_A_47_47#_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.1113 PD=0.98 PS=1.37 NRD=79.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1002 N_A_270_465#_M1002_d N_GATE_N_M1002_g N_VGND_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1176 PD=1.37 PS=0.98 NRD=0 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_270_465#_M1009_g N_A_387_385#_M1009_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1012 A_598_125# N_A_47_47#_M1012_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=31.428 M=1 R=2.8 SA=75000.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1015 N_A_670_125#_M1015_d N_A_270_465#_M1015_g A_598_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 A_756_125# N_A_387_385#_M1006_g N_A_670_125#_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_820_99#_M1019_g A_756_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1013 A_1040_47# N_A_670_125#_M1013_g N_A_820_99#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_RESET_B_M1005_g A_1040_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.0882 PD=1.23 PS=1.05 NRD=7.848 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1010 N_Q_M1010_d N_A_820_99#_M1010_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1638 PD=2.25 PS=1.23 NRD=2.856 NRS=7.848 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_D_M1008_g N_A_47_47#_M1008_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.176 AS=0.1696 PD=1.19 PS=1.81 NRD=6.1464 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.9 A=0.096 P=1.58 MULT=1
MM1011 N_A_270_465#_M1011_d N_GATE_N_M1011_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.176 PD=1.81 PS=1.19 NRD=0 NRS=76.9482 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A_270_465#_M1001_g N_A_387_385#_M1001_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1136 AS=0.3459 PD=0.995 PS=2.7 NRD=12.2928 NRS=149.424 M=1
+ R=4.26667 SA=75000.3 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1004 A_598_447# N_A_47_47#_M1004_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1136 PD=0.85 PS=0.995 NRD=15.3857 NRS=10.7562 M=1 R=4.26667
+ SA=75000.8 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1003 N_A_670_125#_M1003_d N_A_387_385#_M1003_g A_598_447# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.137419 AS=0.0672 PD=1.24377 PS=0.85 NRD=4.6098 NRS=15.3857 M=1
+ R=4.26667 SA=75001.2 SB=75002 A=0.096 P=1.58 MULT=1
MM1016 A_778_447# N_A_270_465#_M1016_g N_A_670_125#_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0901811 PD=0.63 PS=0.816226 NRD=23.443 NRS=45.7237 M=1
+ R=2.8 SA=75001.7 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_820_99#_M1014_g A_778_447# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.13755 AS=0.0441 PD=0.995 PS=0.63 NRD=201.689 NRS=23.443 M=1 R=2.8
+ SA=75002.1 SB=75002 A=0.063 P=1.14 MULT=1
MM1000 N_A_820_99#_M1000_d N_A_670_125#_M1000_g N_VPWR_M1014_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.41265 PD=1.54 PS=2.985 NRD=0 NRS=3.9006 M=1 R=8.4
+ SA=75001.1 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_RESET_B_M1007_g N_A_820_99#_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.1764 PD=1.65 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75001.6 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1017 N_Q_M1017_d N_A_820_99#_M1017_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=10.9335 M=1 R=8.4 SA=75002.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=13.2415 P=17.93
c_72 VNB 0 1.91944e-19 $X=0 $Y=0
c_128 VPB 0 1.73265e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlrtn_1.pxi.spice"
*
.ends
*
*
