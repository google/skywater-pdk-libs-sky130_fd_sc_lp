* File: sky130_fd_sc_lp__xnor3_1.pex.spice
* Created: Wed Sep  2 10:40:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XNOR3_1%A_81_259# 1 2 9 13 18 19 20 22 23 25 28 29
+ 30 34 36
c90 19 0 2.53008e-20 $X=2.245 $Y=0.62
r91 36 39 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.41 $Y=0.62
+ $X2=2.41 $Y2=0.765
r92 32 34 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.695 $Y=2.035
+ $X2=1.035 $Y2=2.035
r93 29 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.46
+ $X2=0.57 $Y2=1.625
r94 29 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.46
+ $X2=0.57 $Y2=1.295
r95 28 31 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=1.46
+ $X2=0.61 $Y2=1.625
r96 28 30 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=1.46
+ $X2=0.61 $Y2=1.295
r97 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.57
+ $Y=1.46 $X2=0.57 $Y2=1.46
r98 23 25 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=1.12 $Y=2.95
+ $X2=2.34 $Y2=2.95
r99 22 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.035 $Y=2.865
+ $X2=1.12 $Y2=2.95
r100 21 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.035 $Y=2.12
+ $X2=1.035 $Y2=2.035
r101 21 22 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.035 $Y=2.12
+ $X2=1.035 $Y2=2.865
r102 19 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0.62
+ $X2=2.41 $Y2=0.62
r103 19 20 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=2.245 $Y=0.62
+ $X2=0.78 $Y2=0.62
r104 18 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=1.95
+ $X2=0.695 $Y2=2.035
r105 18 31 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.695 $Y=1.95
+ $X2=0.695 $Y2=1.625
r106 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.695 $Y=0.705
+ $X2=0.78 $Y2=0.62
r107 15 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.695 $Y=0.705
+ $X2=0.695 $Y2=1.295
r108 13 42 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.49 $Y=0.685
+ $X2=0.49 $Y2=1.295
r109 9 43 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.48 $Y=2.465
+ $X2=0.48 $Y2=1.625
r110 2 25 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=2.255 $X2=2.34 $Y2=2.95
r111 1 39 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=2.2
+ $Y=0.545 $X2=2.41 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%C 3 7 9 13 17 19 20 22 26
c70 7 0 1.71647e-19 $X=1.16 $Y=2.155
c71 3 0 1.62474e-19 $X=1.145 $Y=0.895
r72 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.51
+ $X2=1.19 $Y2=1.675
r73 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=1.51 $X2=1.19 $Y2=1.51
r74 22 25 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.19 $Y=1.42 $X2=1.19
+ $Y2=1.51
r75 22 23 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.19 $Y=1.42 $X2=1.19
+ $Y2=1.345
r76 20 26 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.51
r77 15 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.125 $Y=1.495
+ $X2=2.125 $Y2=1.42
r78 15 17 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=2.125 $Y=1.495
+ $X2=2.125 $Y2=2.675
r79 11 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.125 $Y=1.345
+ $X2=2.125 $Y2=1.42
r80 11 13 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.125 $Y=1.345
+ $X2=2.125 $Y2=0.865
r81 10 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.42
+ $X2=1.19 $Y2=1.42
r82 9 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.05 $Y=1.42
+ $X2=2.125 $Y2=1.42
r83 9 10 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.05 $Y=1.42
+ $X2=1.355 $Y2=1.42
r84 7 27 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.16 $Y=2.155
+ $X2=1.16 $Y2=1.675
r85 3 23 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.145 $Y=0.895
+ $X2=1.145 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%A_244_137# 1 2 9 13 15 20 21 23 24
c66 9 0 2.53008e-20 $X=2.625 $Y=0.865
r67 24 31 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.577 $Y=1.72
+ $X2=2.577 $Y2=1.885
r68 24 30 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.577 $Y=1.72
+ $X2=2.577 $Y2=1.555
r69 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.575
+ $Y=1.72 $X2=2.575 $Y2=1.72
r70 21 28 21.5548 $w=2.83e-07 $l=5.8438e-07 $layer=LI1_cond $X=1.655 $Y=1.72
+ $X2=1.472 $Y2=2.22
r71 21 23 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=1.655 $Y=1.72
+ $X2=2.575 $Y2=1.72
r72 20 21 9.04317 $w=2.83e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.57 $Y=1.555
+ $X2=1.655 $Y2=1.72
r73 19 20 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.57 $Y=1.125
+ $X2=1.57 $Y2=1.555
r74 15 19 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.485 $Y=1
+ $X2=1.57 $Y2=1.125
r75 15 17 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.485 $Y=1 $X2=1.36
+ $Y2=1
r76 13 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.67 $Y=2.465
+ $X2=2.67 $Y2=1.885
r77 9 30 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.625 $Y=0.865
+ $X2=2.625 $Y2=1.555
r78 2 28 600 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.835 $X2=1.375 $Y2=2.22
r79 1 17 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.22
+ $Y=0.685 $X2=1.36 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%A_754_367# 1 2 9 14 15 16 19 24 27 30 31 34
+ 39 41 45 50
c115 50 0 1.30013e-19 $X=4.83 $Y=1.54
c116 45 0 1.11774e-19 $X=4.655 $Y=1.54
c117 39 0 8.84612e-20 $X=4.185 $Y=2.075
c118 27 0 2.6204e-19 $X=5.95 $Y=1.415
c119 14 0 1.01023e-19 $X=4.905 $Y=0.945
r120 50 51 11.9702 $w=3.02e-07 $l=7.5e-08 $layer=POLY_cond $X=4.83 $Y=1.54
+ $X2=4.905 $Y2=1.54
r121 46 50 27.9305 $w=3.02e-07 $l=1.75e-07 $layer=POLY_cond $X=4.655 $Y=1.54
+ $X2=4.83 $Y2=1.54
r122 45 48 8.49766 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=4.637 $Y=1.54
+ $X2=4.637 $Y2=1.705
r123 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.655
+ $Y=1.54 $X2=4.655 $Y2=1.54
r124 38 39 5.10546 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=2.075
+ $X2=4.185 $Y2=2.075
r125 36 38 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=3.91 $Y=2.075
+ $X2=4.1 $Y2=2.075
r126 34 48 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.575 $Y=2.03
+ $X2=4.575 $Y2=1.705
r127 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=2.115
+ $X2=4.575 $Y2=2.03
r128 31 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.49 $Y=2.115
+ $X2=4.185 $Y2=2.115
r129 30 38 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.1 $Y=1.95 $X2=4.1
+ $Y2=2.075
r130 29 41 0.716491 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.1 $Y=1.125
+ $X2=4.015 $Y2=1.04
r131 29 30 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.1 $Y=1.125
+ $X2=4.1 $Y2=1.95
r132 25 27 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=5.805 $Y=1.415
+ $X2=5.95 $Y2=1.415
r133 22 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.95 $Y=1.34
+ $X2=5.95 $Y2=1.415
r134 22 24 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.95 $Y=1.34
+ $X2=5.95 $Y2=0.79
r135 21 24 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.95 $Y=0.255
+ $X2=5.95 $Y2=0.79
r136 17 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.805 $Y=1.49
+ $X2=5.805 $Y2=1.415
r137 17 19 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.805 $Y=1.49
+ $X2=5.805 $Y2=2.185
r138 15 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.875 $Y=0.18
+ $X2=5.95 $Y2=0.255
r139 15 16 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=5.875 $Y=0.18
+ $X2=4.98 $Y2=0.18
r140 12 51 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.905 $Y=1.375
+ $X2=4.905 $Y2=1.54
r141 12 14 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.905 $Y=1.375
+ $X2=4.905 $Y2=0.945
r142 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.905 $Y=0.255
+ $X2=4.98 $Y2=0.18
r143 11 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.905 $Y=0.255
+ $X2=4.905 $Y2=0.945
r144 7 50 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.83 $Y=1.705
+ $X2=4.83 $Y2=1.54
r145 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.83 $Y=1.705
+ $X2=4.83 $Y2=2.285
r146 2 36 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=3.77
+ $Y=1.835 $X2=3.91 $Y2=2.035
r147 1 41 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.875
+ $Y=0.345 $X2=4.015 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%B 3 7 9 12 13 14 18 21 23 28 31 34 35 38 40
+ 43 44
c130 38 0 1.66518e-19 $X=6.54 $Y=1.63
c131 31 0 7.27944e-20 $X=6.54 $Y=0.68
c132 21 0 1.29867e-19 $X=5.405 $Y=0.945
c133 9 0 8.84612e-20 $X=4.13 $Y=1.6
r134 43 46 14.4261 $w=3.6e-07 $l=9e-08 $layer=POLY_cond $X=3.695 $Y=1.51
+ $X2=3.695 $Y2=1.6
r135 43 45 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=1.51
+ $X2=3.695 $Y2=1.345
r136 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.68
+ $Y=1.51 $X2=3.68 $Y2=1.51
r137 40 44 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.68 $Y=1.665
+ $X2=3.68 $Y2=1.51
r138 36 38 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.45 $Y=1.63 $X2=6.54
+ $Y2=1.63
r139 33 34 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.39 $Y=1.605
+ $X2=5.39 $Y2=1.755
r140 29 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.54 $Y=1.555
+ $X2=6.54 $Y2=1.63
r141 29 31 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=6.54 $Y=1.555
+ $X2=6.54 $Y2=0.68
r142 26 28 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.45 $Y=3.075
+ $X2=6.45 $Y2=2.285
r143 25 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.45 $Y=1.705
+ $X2=6.45 $Y2=1.63
r144 25 28 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.45 $Y=1.705
+ $X2=6.45 $Y2=2.285
r145 24 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.45 $Y=3.15
+ $X2=5.375 $Y2=3.15
r146 23 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.375 $Y=3.15
+ $X2=6.45 $Y2=3.075
r147 23 24 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=6.375 $Y=3.15
+ $X2=5.45 $Y2=3.15
r148 21 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.405 $Y=0.945
+ $X2=5.405 $Y2=1.605
r149 18 34 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.375 $Y=2.185
+ $X2=5.375 $Y2=1.755
r150 16 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.375 $Y=3.075
+ $X2=5.375 $Y2=3.15
r151 16 18 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=5.375 $Y=3.075
+ $X2=5.375 $Y2=2.185
r152 13 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.3 $Y=3.15
+ $X2=5.375 $Y2=3.15
r153 13 14 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=5.3 $Y=3.15
+ $X2=4.28 $Y2=3.15
r154 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.205 $Y=3.075
+ $X2=4.28 $Y2=3.15
r155 11 12 717.872 $w=1.5e-07 $l=1.4e-06 $layer=POLY_cond $X=4.205 $Y=1.675
+ $X2=4.205 $Y2=3.075
r156 10 46 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.875 $Y=1.6
+ $X2=3.695 $Y2=1.6
r157 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.13 $Y=1.6
+ $X2=4.205 $Y2=1.675
r158 9 10 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=4.13 $Y=1.6
+ $X2=3.875 $Y2=1.6
r159 7 45 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.8 $Y=0.765 $X2=3.8
+ $Y2=1.345
r160 1 46 32.1566 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=3.695 $Y=1.675
+ $X2=3.695 $Y2=1.6
r161 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.695 $Y=1.675
+ $X2=3.695 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%A 3 7 9 12
c50 12 0 1.19914e-19 $X=7.02 $Y=1.345
c51 7 0 1.89142e-19 $X=7.11 $Y=2.415
c52 3 0 1.50571e-20 $X=6.995 $Y=0.68
r53 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.02 $Y=1.345
+ $X2=7.02 $Y2=1.51
r54 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.02 $Y=1.345
+ $X2=7.02 $Y2=1.18
r55 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.02
+ $Y=1.345 $X2=7.02 $Y2=1.345
r56 7 15 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=7.11 $Y=2.415
+ $X2=7.11 $Y2=1.51
r57 3 14 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.995 $Y=0.68 $X2=6.995
+ $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%A_871_373# 1 2 3 4 15 19 21 23 28 29 32 35
+ 36 37 42 44 51 55 56 57
c122 56 0 1.66176e-19 $X=7.56 $Y=1.355
r123 56 61 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.575 $Y=1.355
+ $X2=7.575 $Y2=1.52
r124 56 60 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.575 $Y=1.355
+ $X2=7.575 $Y2=1.19
r125 55 58 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.5 $Y=1.355
+ $X2=7.5 $Y2=1.52
r126 55 57 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.5 $Y=1.355
+ $X2=7.5 $Y2=1.19
r127 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.56
+ $Y=1.355 $X2=7.56 $Y2=1.355
r128 49 51 9.77977 $w=1.88e-07 $l=1.65e-07 $layer=LI1_cond $X=4.575 $Y=0.35
+ $X2=4.74 $Y2=0.35
r129 44 46 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.5 $Y=2.795
+ $X2=4.5 $Y2=2.98
r130 42 58 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.44 $Y=1.845
+ $X2=7.44 $Y2=1.52
r131 39 57 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.44 $Y=0.945
+ $X2=7.44 $Y2=1.19
r132 38 53 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.945 $Y=2.01
+ $X2=6.78 $Y2=2.01
r133 37 42 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.355 $Y=2.01
+ $X2=7.44 $Y2=1.845
r134 37 38 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.355 $Y=2.01
+ $X2=6.945 $Y2=2.01
r135 35 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.355 $Y=0.86
+ $X2=7.44 $Y2=0.945
r136 35 36 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=7.355 $Y=0.86
+ $X2=6.945 $Y2=0.86
r137 32 34 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.78 $Y=2.43
+ $X2=6.78 $Y2=2.77
r138 30 34 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=6.78 $Y=2.895
+ $X2=6.78 $Y2=2.77
r139 29 53 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=2.175
+ $X2=6.78 $Y2=2.01
r140 29 32 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.78 $Y=2.175
+ $X2=6.78 $Y2=2.43
r141 26 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.78 $Y=0.775
+ $X2=6.945 $Y2=0.86
r142 26 28 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.78 $Y=0.775
+ $X2=6.78 $Y2=0.505
r143 25 28 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.78 $Y=0.425 $X2=6.78
+ $Y2=0.505
r144 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.615 $Y=0.34
+ $X2=6.78 $Y2=0.425
r145 23 51 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=6.615 $Y=0.34
+ $X2=4.74 $Y2=0.34
r146 22 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=2.98
+ $X2=4.5 $Y2=2.98
r147 21 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.615 $Y=2.98
+ $X2=6.78 $Y2=2.895
r148 21 22 127.219 $w=1.68e-07 $l=1.95e-06 $layer=LI1_cond $X=6.615 $Y=2.98
+ $X2=4.665 $Y2=2.98
r149 19 61 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=7.645 $Y=2.415
+ $X2=7.645 $Y2=1.52
r150 15 60 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.645 $Y=0.68
+ $X2=7.645 $Y2=1.19
r151 4 53 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.865 $X2=6.78 $Y2=2.01
r152 4 34 600 $w=1.7e-07 $l=1.0246e-06 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.865 $X2=6.78 $Y2=2.77
r153 4 32 600 $w=1.7e-07 $l=6.80661e-07 $layer=licon1_PDIFF $count=1 $X=6.525
+ $Y=1.865 $X2=6.78 $Y2=2.43
r154 3 44 600 $w=1.7e-07 $l=9.99875e-07 $layer=licon1_PDIFF $count=1 $X=4.355
+ $Y=1.865 $X2=4.5 $Y2=2.795
r155 2 28 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=6.615
+ $Y=0.36 $X2=6.78 $Y2=0.505
r156 1 49 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.215 $X2=4.575 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%X 1 2 9 11 15 16 17 23 29
c22 23 0 1.62474e-19 $X=0.275 $Y=0.42
r23 21 29 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=0.27 $Y=0.955 $X2=0.27
+ $Y2=0.925
r24 17 31 7.72622 $w=3.38e-07 $l=1.43e-07 $layer=LI1_cond $X=0.27 $Y=0.982
+ $X2=0.27 $Y2=1.125
r25 17 21 0.915175 $w=3.38e-07 $l=2.7e-08 $layer=LI1_cond $X=0.27 $Y=0.982
+ $X2=0.27 $Y2=0.955
r26 17 29 0.949071 $w=3.38e-07 $l=2.8e-08 $layer=LI1_cond $X=0.27 $Y=0.897
+ $X2=0.27 $Y2=0.925
r27 16 17 11.5922 $w=3.38e-07 $l=3.42e-07 $layer=LI1_cond $X=0.27 $Y=0.555
+ $X2=0.27 $Y2=0.897
r28 16 23 4.57588 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=0.27 $Y=0.555
+ $X2=0.27 $Y2=0.42
r29 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.185 $Y=1.815
+ $X2=0.185 $Y2=1.125
r30 11 13 42.8709 $w=2.48e-07 $l=9.3e-07 $layer=LI1_cond $X=0.225 $Y=1.98
+ $X2=0.225 $Y2=2.91
r31 9 15 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.225 $Y=1.94
+ $X2=0.225 $Y2=1.815
r32 9 11 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=0.225 $Y=1.94 $X2=0.225
+ $Y2=1.98
r33 2 13 400 $w=1.7e-07 $l=1.13815e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.265 $Y2=2.91
r34 2 11 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.265 $Y2=1.98
r35 1 23 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.265 $X2=0.275 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%VPWR 1 2 3 12 16 20 23 24 25 27 32 42 43 46
+ 49
c78 32 0 1.71647e-19 $X=3.315 $Y=3.33
r79 49 50 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r80 46 47 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r82 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r83 39 40 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r84 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=3.48 $Y2=3.33
r85 37 39 216.273 $w=1.68e-07 $l=3.315e-06 $layer=LI1_cond $X=3.645 $Y=3.33
+ $X2=6.96 $Y2=3.33
r86 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r87 36 47 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=0.72 $Y2=3.33
r88 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r89 33 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.78 $Y=3.33
+ $X2=0.655 $Y2=3.33
r90 33 35 152.663 $w=1.68e-07 $l=2.34e-06 $layer=LI1_cond $X=0.78 $Y=3.33
+ $X2=3.12 $Y2=3.33
r91 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.48 $Y2=3.33
r92 32 35 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.12 $Y2=3.33
r93 30 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r94 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r95 27 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.655 $Y2=3.33
r96 27 29 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.24 $Y2=3.33
r97 25 40 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6.96 $Y2=3.33
r98 25 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r99 23 39 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.16 $Y=3.33 $X2=6.96
+ $Y2=3.33
r100 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.16 $Y=3.33
+ $X2=7.325 $Y2=3.33
r101 22 42 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.49 $Y=3.33
+ $X2=7.92 $Y2=3.33
r102 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.49 $Y=3.33
+ $X2=7.325 $Y2=3.33
r103 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.325 $Y=3.245
+ $X2=7.325 $Y2=3.33
r104 18 20 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=7.325 $Y=3.245
+ $X2=7.325 $Y2=2.43
r105 14 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=3.245
+ $X2=3.48 $Y2=3.33
r106 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.48 $Y=3.245
+ $X2=3.48 $Y2=2.95
r107 10 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.655 $Y=3.245
+ $X2=0.655 $Y2=3.33
r108 10 12 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.655 $Y=3.245
+ $X2=0.655 $Y2=2.455
r109 3 20 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=7.185
+ $Y=1.915 $X2=7.325 $Y2=2.43
r110 2 16 600 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=3.335
+ $Y=1.835 $X2=3.48 $Y2=2.95
r111 1 12 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.835 $X2=0.695 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%A_355_451# 1 2 3 4 15 17 18 20 22 23 25 27
+ 29 34 39 40 41
c136 41 0 1.66518e-19 $X=6.28 $Y=0.68
c137 29 0 1.51199e-19 $X=6.115 $Y=0.68
c138 27 0 1.30013e-19 $X=5.045 $Y=2.04
r139 41 44 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.28 $Y=0.68
+ $X2=6.28 $Y2=0.765
r140 39 40 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=4.91 $Y=0.69
+ $X2=5.08 $Y2=0.69
r141 34 35 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.26 $Y=2.455
+ $X2=3.26 $Y2=2.61
r142 32 33 9.61712 $w=4.44e-07 $l=3.5e-07 $layer=LI1_cond $X=2.91 $Y=0.767
+ $X2=3.26 $Y2=0.767
r143 29 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=0.68
+ $X2=6.28 $Y2=0.68
r144 29 40 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=6.115 $Y=0.68
+ $X2=5.08 $Y2=0.68
r145 25 38 3.16731 $w=3.3e-07 $l=1.77e-07 $layer=LI1_cond $X=5.045 $Y=2.37
+ $X2=5.045 $Y2=2.547
r146 25 27 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.045 $Y=2.37
+ $X2=5.045 $Y2=2.04
r147 24 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=2.455
+ $X2=3.26 $Y2=2.455
r148 23 38 4.59886 $w=1.7e-07 $l=2.05925e-07 $layer=LI1_cond $X=4.88 $Y=2.455
+ $X2=5.045 $Y2=2.547
r149 23 24 100.144 $w=1.68e-07 $l=1.535e-06 $layer=LI1_cond $X=4.88 $Y=2.455
+ $X2=3.345 $Y2=2.455
r150 22 33 7.17697 $w=4.44e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.345 $Y=0.7
+ $X2=3.26 $Y2=0.767
r151 22 39 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=3.345 $Y=0.7
+ $X2=4.91 $Y2=0.7
r152 20 34 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=2.37
+ $X2=3.26 $Y2=2.455
r153 19 33 6.41743 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=3.26 $Y=1.01
+ $X2=3.26 $Y2=0.767
r154 19 20 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.26 $Y=1.01
+ $X2=3.26 $Y2=2.37
r155 17 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.175 $Y=2.61
+ $X2=3.26 $Y2=2.61
r156 17 18 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=3.175 $Y=2.61
+ $X2=2.075 $Y2=2.61
r157 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.95 $Y=2.525
+ $X2=2.075 $Y2=2.61
r158 13 15 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=1.95 $Y=2.525
+ $X2=1.95 $Y2=2.465
r159 4 38 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=1.865 $X2=5.045 $Y2=2.56
r160 4 27 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=1.865 $X2=5.045 $Y2=2.04
r161 3 15 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=1.775
+ $Y=2.255 $X2=1.91 $Y2=2.465
r162 2 44 182 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_NDIFF $count=1 $X=6.025
+ $Y=0.58 $X2=6.28 $Y2=0.765
r163 1 32 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.545 $X2=2.91 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%A_354_109# 1 2 3 4 15 19 21 22 25 27 28 31
+ 35 36 42 43
r104 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.295
r105 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.295
r106 36 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.295
+ $X2=2.64 $Y2=1.295
r107 35 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=5.04 $Y2=1.295
r108 35 36 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=2.785 $Y2=1.295
r109 34 43 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.12 $Y=1.455
+ $X2=5.12 $Y2=1.295
r110 33 43 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.12 $Y=1.205
+ $X2=5.12 $Y2=1.295
r111 31 33 5.38305 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.105 $Y=1.04
+ $X2=5.105 $Y2=1.205
r112 28 39 10.5499 $w=2.03e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=1.282
+ $X2=2.64 $Y2=1.282
r113 27 39 30.5676 $w=2.03e-07 $l=5.65e-07 $layer=LI1_cond $X=2.075 $Y=1.282
+ $X2=2.64 $Y2=1.282
r114 23 25 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=6.02 $Y=1.625
+ $X2=6.02 $Y2=2.095
r115 22 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.285 $Y=1.54
+ $X2=5.12 $Y2=1.455
r116 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.935 $Y=1.54
+ $X2=6.02 $Y2=1.625
r117 21 22 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.935 $Y=1.54
+ $X2=5.285 $Y2=1.54
r118 17 28 6.89401 $w=2.05e-07 $l=1.39155e-07 $layer=LI1_cond $X=2.92 $Y=1.385
+ $X2=2.835 $Y2=1.282
r119 17 19 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=2.92 $Y=1.385
+ $X2=2.92 $Y2=2.19
r120 13 27 6.90357 $w=2.05e-07 $l=1.68449e-07 $layer=LI1_cond $X=1.95 $Y=1.18
+ $X2=2.075 $Y2=1.282
r121 13 15 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=1.95 $Y=1.18
+ $X2=1.95 $Y2=1.04
r122 4 25 600 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_PDIFF $count=1 $X=5.88
+ $Y=1.865 $X2=6.02 $Y2=2.095
r123 3 19 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=2.045 $X2=2.92 $Y2=2.19
r124 2 31 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=4.98
+ $Y=0.625 $X2=5.12 $Y2=1.04
r125 1 15 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.545 $X2=1.91 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%A_1090_373# 1 2 3 4 13 14 15 18 20 23 29 33
+ 34 37 38 39 40 46 47 50
c108 37 0 1.89142e-19 $X=7.86 $Y=2.06
c109 34 0 1.50571e-20 $X=7.885 $Y=1.02
c110 33 0 1.36914e-19 $X=6.42 $Y=1.675
c111 29 0 1.73817e-19 $X=5.62 $Y=1.11
c112 18 0 1.1084e-19 $X=6.42 $Y=1.53
c113 15 0 1.38007e-19 $X=6.275 $Y=1.2
r114 47 55 11.0695 $w=3.78e-07 $l=3.65e-07 $layer=LI1_cond $X=7.885 $Y=2.405
+ $X2=7.885 $Y2=2.77
r115 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.405
+ $X2=7.92 $Y2=2.405
r116 43 50 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=5.59 $Y=2.405
+ $X2=5.59 $Y2=2.01
r117 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.405
+ $X2=5.52 $Y2=2.405
r118 40 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.405
+ $X2=5.52 $Y2=2.405
r119 39 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.405
+ $X2=7.92 $Y2=2.405
r120 39 40 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=7.775 $Y=2.405
+ $X2=5.665 $Y2=2.405
r121 37 38 6.56115 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=7.885 $Y=2.06
+ $X2=7.885 $Y2=1.895
r122 35 47 9.70478 $w=3.78e-07 $l=3.2e-07 $layer=LI1_cond $X=7.885 $Y=2.085
+ $X2=7.885 $Y2=2.405
r123 35 37 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=7.885 $Y=2.085
+ $X2=7.885 $Y2=2.06
r124 34 38 42.0162 $w=2.38e-07 $l=8.75e-07 $layer=LI1_cond $X=7.955 $Y=1.02
+ $X2=7.955 $Y2=1.895
r125 29 31 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.62 $Y=1.11 $X2=5.62
+ $Y2=1.2
r126 27 43 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=5.59 $Y=2.515
+ $X2=5.59 $Y2=2.405
r127 21 34 7.31933 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=7.885 $Y=0.83
+ $X2=7.885 $Y2=1.02
r128 21 23 9.85642 $w=3.78e-07 $l=3.25e-07 $layer=LI1_cond $X=7.885 $Y=0.83
+ $X2=7.885 $Y2=0.505
r129 20 33 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.36 $Y=2.515
+ $X2=6.36 $Y2=1.675
r130 18 33 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=6.42 $Y=1.53
+ $X2=6.42 $Y2=1.675
r131 17 18 9.73616 $w=2.88e-07 $l=2.45e-07 $layer=LI1_cond $X=6.42 $Y=1.285
+ $X2=6.42 $Y2=1.53
r132 16 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=1.2
+ $X2=5.62 $Y2=1.2
r133 15 17 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=6.275 $Y=1.2
+ $X2=6.42 $Y2=1.285
r134 15 16 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=6.275 $Y=1.2
+ $X2=5.785 $Y2=1.2
r135 14 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.755 $Y=2.6
+ $X2=5.59 $Y2=2.515
r136 13 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.275 $Y=2.6
+ $X2=6.36 $Y2=2.515
r137 13 14 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.275 $Y=2.6
+ $X2=5.755 $Y2=2.6
r138 4 55 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=7.72
+ $Y=1.915 $X2=7.86 $Y2=2.77
r139 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.72
+ $Y=1.915 $X2=7.86 $Y2=2.06
r140 3 50 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=5.45
+ $Y=1.865 $X2=5.59 $Y2=2.01
r141 2 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.72
+ $Y=0.36 $X2=7.86 $Y2=0.505
r142 1 29 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.625 $X2=5.62 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LP__XNOR3_1%VGND 1 2 3 14 18 21 22 23 25 38 39 43 49
c65 18 0 1.66176e-19 $X=7.28 $Y=0.505
r66 49 50 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r67 43 46 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.815
+ $Y2=0.28
r68 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r70 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r71 35 36 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r72 33 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=0 $X2=3.47
+ $Y2=0
r73 33 35 216.925 $w=1.68e-07 $l=3.325e-06 $layer=LI1_cond $X=3.635 $Y=0
+ $X2=6.96 $Y2=0
r74 32 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r75 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r76 29 32 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r77 29 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r78 28 31 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r79 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r80 26 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r81 26 28 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r82 25 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.47
+ $Y2=0
r83 25 31 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.12
+ $Y2=0
r84 23 36 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6.96
+ $Y2=0
r85 23 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r86 21 35 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.115 $Y=0 $X2=6.96
+ $Y2=0
r87 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.115 $Y=0 $X2=7.28
+ $Y2=0
r88 20 38 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=7.445 $Y=0 $X2=7.92
+ $Y2=0
r89 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.445 $Y=0 $X2=7.28
+ $Y2=0
r90 16 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.28 $Y=0.085
+ $X2=7.28 $Y2=0
r91 16 18 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=7.28 $Y=0.085
+ $X2=7.28 $Y2=0.505
r92 12 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=0.085
+ $X2=3.47 $Y2=0
r93 12 14 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.47 $Y=0.085
+ $X2=3.47 $Y2=0.36
r94 3 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.07
+ $Y=0.36 $X2=7.28 $Y2=0.505
r95 2 14 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.215 $X2=3.47 $Y2=0.36
r96 1 46 182 $w=1.7e-07 $l=2.57391e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.265 $X2=0.815 $Y2=0.28
.ends

