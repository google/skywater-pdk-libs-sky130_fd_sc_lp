* NGSPICE file created from sky130_fd_sc_lp__a41oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_103_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.079e+12p pd=1.842e+07u as=2.5641e+12p ps=1.415e+07u
M1001 a_103_367# B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1002 a_318_69# A2 a_577_69# VNB nshort w=840000u l=150000u
+  ad=7.56e+11p pd=6.84e+06u as=4.704e+11p ps=4.48e+06u
M1003 VPWR A4 a_103_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_318_69# A1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.48e+06u
M1005 a_788_69# A3 a_577_69# VNB nshort w=840000u l=150000u
+  ad=7.392e+11p pd=6.8e+06u as=0p ps=0u
M1006 VPWR A3 a_103_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_103_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_103_367# A3 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A4 a_788_69# VNB nshort w=840000u l=150000u
+  ad=6.804e+11p pd=6.66e+06u as=0p ps=0u
M1010 VPWR A2 a_103_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_103_367# A4 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_577_69# A2 a_318_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A1 a_103_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A1 a_318_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_577_69# A3 a_788_69# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_103_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_788_69# A4 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

