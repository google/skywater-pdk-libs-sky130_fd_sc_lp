* File: sky130_fd_sc_lp__nand4b_4.spice
* Created: Fri Aug 28 10:51:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4b_4.pex.spice"
.subckt sky130_fd_sc_lp__nand4b_4  VNB VPB A_N B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1027 N_VGND_M1027_d N_A_N_M1027_g N_A_27_51#_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_217_51#_M1001_d N_A_27_51#_M1001_g N_Y_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1005 N_A_217_51#_M1005_d N_A_27_51#_M1005_g N_Y_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1018 N_A_217_51#_M1005_d N_A_27_51#_M1018_g N_Y_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1020 N_A_217_51#_M1020_d N_A_27_51#_M1020_g N_Y_M1018_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1002 N_A_644_51#_M1002_d N_B_M1002_g N_A_217_51#_M1020_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=11.424 NRS=0 M=1 R=5.6
+ SA=75001.9 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1011 N_A_644_51#_M1002_d N_B_M1011_g N_A_217_51#_M1011_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1512 AS=0.1176 PD=1.2 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1013 N_A_644_51#_M1013_d N_B_M1013_g N_A_217_51#_M1011_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1023 N_A_644_51#_M1013_d N_B_M1023_g N_A_217_51#_M1023_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_A_1025_65#_M1003_d N_C_M1003_g N_A_644_51#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1014 N_A_1025_65#_M1014_d N_C_M1014_g N_A_644_51#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1025 N_A_1025_65#_M1014_d N_C_M1025_g N_A_644_51#_M1025_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6
+ SA=75001.1 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1028 N_A_1025_65#_M1028_d N_C_M1028_g N_A_644_51#_M1025_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_D_M1012_g N_A_1025_65#_M1028_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1012_d N_D_M1015_g N_A_1025_65#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1024_d N_D_M1024_g N_A_1025_65#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1032 N_VGND_M1024_d N_D_M1032_g N_A_1025_65#_M1032_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_27_51#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1827 AS=0.3339 PD=1.55 PS=3.05 NRD=1.5563 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75007.9 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1000_d N_A_27_51#_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1827 AS=0.1764 PD=1.55 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75007.4 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A_27_51#_M1008_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75007 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1008_d N_A_27_51#_M1021_g N_Y_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75006.5 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1026_d N_A_27_51#_M1026_g N_Y_M1021_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.189 AS=0.1764 PD=1.56 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75006.1
+ A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1026_d N_B_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.26 AD=0.189
+ AS=0.1764 PD=1.56 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75002.4 SB=75005.6
+ A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_B_M1017_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75005.2 A=0.189 P=2.82 MULT=1
MM1029 N_VPWR_M1017_d N_B_M1029_g N_Y_M1029_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.3
+ SB=75004.8 A=0.189 P=2.82 MULT=1
MM1033 N_VPWR_M1033_d N_B_M1033_g N_Y_M1029_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.1764 PD=1.88 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1033_d N_C_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.1764 PD=1.88 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_C_M1010_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.9
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1010_d N_C_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.4
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1031 N_VPWR_M1031_d N_C_M1031_g N_Y_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4095 AS=0.1764 PD=1.91 PS=1.54 NRD=4.6886 NRS=0 M=1 R=8.4 SA=75005.8
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1031_d N_D_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4095 AS=0.1764 PD=1.91 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_D_M1016_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007 SB=75001.1
+ A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1016_d N_D_M1022_g N_Y_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1030 N_VPWR_M1030_d N_D_M1030_g N_Y_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75007.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=17.7175 P=22.73
*
.include "sky130_fd_sc_lp__nand4b_4.pxi.spice"
*
.ends
*
*
