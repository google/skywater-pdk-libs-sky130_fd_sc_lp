* NGSPICE file created from sky130_fd_sc_lp__a32o_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a32o_lp A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_30_419# B1 a_137_419# VPB phighvt w=1e+06u l=250000u
+  ad=8.45e+11p pd=7.69e+06u as=2.8e+11p ps=2.56e+06u
M1001 a_137_141# B2 VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.192e+11p ps=3.2e+06u
M1002 X a_137_419# a_682_141# VNB nshort w=420000u l=150000u
+  ad=1.575e+11p pd=1.59e+06u as=1.008e+11p ps=1.32e+06u
M1003 VPWR A3 a_30_419# VPB phighvt w=1e+06u l=250000u
+  ad=1.125e+12p pd=6.25e+06u as=0p ps=0u
M1004 X a_137_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1005 a_682_141# a_137_419# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_137_419# B2 a_30_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_30_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_329_141# A1 a_137_419# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=1.764e+11p ps=1.68e+06u
M1009 VGND A3 a_443_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
M1010 a_137_419# B1 a_137_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_443_141# A2 a_329_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_30_419# A2 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

