* File: sky130_fd_sc_lp__or4bb_2.pxi.spice
* Created: Wed Sep  2 10:33:12 2020
* 
x_PM_SKY130_FD_SC_LP__OR4BB_2%C_N N_C_N_M1003_g N_C_N_c_105_n N_C_N_c_106_n
+ N_C_N_c_112_n N_C_N_c_113_n N_C_N_M1007_g N_C_N_c_107_n C_N C_N C_N
+ N_C_N_c_109_n N_C_N_c_110_n PM_SKY130_FD_SC_LP__OR4BB_2%C_N
x_PM_SKY130_FD_SC_LP__OR4BB_2%A N_A_M1000_g N_A_M1002_g N_A_c_152_n N_A_c_153_n
+ N_A_c_154_n A A N_A_c_156_n PM_SKY130_FD_SC_LP__OR4BB_2%A
x_PM_SKY130_FD_SC_LP__OR4BB_2%B N_B_M1004_g N_B_M1006_g B N_B_c_192_n
+ N_B_c_193_n PM_SKY130_FD_SC_LP__OR4BB_2%B
x_PM_SKY130_FD_SC_LP__OR4BB_2%A_40_47# N_A_40_47#_M1003_s N_A_40_47#_M1007_s
+ N_A_40_47#_M1012_g N_A_40_47#_M1010_g N_A_40_47#_c_229_n N_A_40_47#_c_230_n
+ N_A_40_47#_c_236_n N_A_40_47#_c_231_n N_A_40_47#_c_232_n N_A_40_47#_c_233_n
+ N_A_40_47#_c_234_n PM_SKY130_FD_SC_LP__OR4BB_2%A_40_47#
x_PM_SKY130_FD_SC_LP__OR4BB_2%A_462_351# N_A_462_351#_M1009_d
+ N_A_462_351#_M1011_d N_A_462_351#_c_308_n N_A_462_351#_M1015_g
+ N_A_462_351#_c_309_n N_A_462_351#_c_310_n N_A_462_351#_c_301_n
+ N_A_462_351#_M1001_g N_A_462_351#_c_312_n N_A_462_351#_c_303_n
+ N_A_462_351#_c_313_n N_A_462_351#_c_314_n N_A_462_351#_c_315_n
+ N_A_462_351#_c_316_n N_A_462_351#_c_304_n N_A_462_351#_c_318_n
+ N_A_462_351#_c_305_n N_A_462_351#_c_306_n N_A_462_351#_c_319_n
+ N_A_462_351#_c_307_n N_A_462_351#_c_343_p N_A_462_351#_c_320_n
+ PM_SKY130_FD_SC_LP__OR4BB_2%A_462_351#
x_PM_SKY130_FD_SC_LP__OR4BB_2%A_276_47# N_A_276_47#_M1000_d N_A_276_47#_M1010_d
+ N_A_276_47#_M1015_d N_A_276_47#_c_410_n N_A_276_47#_M1008_g
+ N_A_276_47#_c_411_n N_A_276_47#_M1005_g N_A_276_47#_c_412_n
+ N_A_276_47#_c_413_n N_A_276_47#_M1014_g N_A_276_47#_M1013_g
+ N_A_276_47#_c_415_n N_A_276_47#_c_516_p N_A_276_47#_c_416_n
+ N_A_276_47#_c_417_n N_A_276_47#_c_418_n N_A_276_47#_c_419_n
+ N_A_276_47#_c_420_n N_A_276_47#_c_421_n N_A_276_47#_c_426_n
+ N_A_276_47#_c_422_n PM_SKY130_FD_SC_LP__OR4BB_2%A_276_47#
x_PM_SKY130_FD_SC_LP__OR4BB_2%D_N N_D_N_M1009_g N_D_N_M1011_g D_N N_D_N_c_531_n
+ PM_SKY130_FD_SC_LP__OR4BB_2%D_N
x_PM_SKY130_FD_SC_LP__OR4BB_2%VPWR N_VPWR_M1007_d N_VPWR_M1005_s N_VPWR_M1013_s
+ N_VPWR_c_556_n N_VPWR_c_557_n N_VPWR_c_558_n VPWR N_VPWR_c_559_n
+ N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_555_n N_VPWR_c_564_n
+ N_VPWR_c_565_n N_VPWR_c_566_n PM_SKY130_FD_SC_LP__OR4BB_2%VPWR
x_PM_SKY130_FD_SC_LP__OR4BB_2%X N_X_M1008_s N_X_M1005_d X X X X X N_X_c_606_n
+ PM_SKY130_FD_SC_LP__OR4BB_2%X
x_PM_SKY130_FD_SC_LP__OR4BB_2%VGND N_VGND_M1003_d N_VGND_M1006_d N_VGND_M1001_d
+ N_VGND_M1014_d N_VGND_c_627_n N_VGND_c_628_n N_VGND_c_629_n N_VGND_c_630_n
+ N_VGND_c_631_n N_VGND_c_632_n N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n
+ VGND N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n
+ PM_SKY130_FD_SC_LP__OR4BB_2%VGND
cc_1 VNB N_C_N_c_105_n 0.0234648f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.248
cc_2 VNB N_C_N_c_106_n 0.0108435f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.685
cc_3 VNB N_C_N_c_107_n 0.0177249f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.435
cc_4 VNB C_N 0.00259293f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB N_C_N_c_109_n 0.0216353f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.93
cc_6 VNB N_C_N_c_110_n 0.0211191f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=0.765
cc_7 VNB N_A_M1002_g 0.0146457f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.435
cc_8 VNB N_A_c_152_n 0.0192983f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.76
cc_9 VNB N_A_c_153_n 0.0208705f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.835
cc_10 VNB N_A_c_154_n 0.0155102f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.225
cc_11 VNB A 0.00811283f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.225
cc_12 VNB N_A_c_156_n 0.0155836f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_B_M1004_g 0.0205989f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.445
cc_14 VNB N_B_M1006_g 0.0226959f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.685
cc_15 VNB N_B_c_192_n 0.030449f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.225
cc_16 VNB N_B_c_193_n 0.00842937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_40_47#_M1012_g 0.00609692f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.76
cc_18 VNB N_A_40_47#_M1010_g 0.0236226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_40_47#_c_229_n 0.0522528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_40_47#_c_230_n 0.0641837f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=0.765
cc_21 VNB N_A_40_47#_c_231_n 0.0161005f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.295
cc_22 VNB N_A_40_47#_c_232_n 0.00504292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_40_47#_c_233_n 0.00127237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_40_47#_c_234_n 0.01582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_462_351#_c_301_n 0.0323401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_462_351#_M1001_g 0.0182119f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_27 VNB N_A_462_351#_c_303_n 0.0122341f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=0.93
cc_28 VNB N_A_462_351#_c_304_n 0.00315987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_462_351#_c_305_n 0.0158322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_462_351#_c_306_n 6.42811e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_462_351#_c_307_n 0.0146462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_276_47#_c_410_n 0.0171341f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.835
cc_33 VNB N_A_276_47#_c_411_n 0.0470709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_276_47#_c_412_n 0.0111523f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_35 VNB N_A_276_47#_c_413_n 0.0188722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_276_47#_M1013_g 0.0158543f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.93
cc_37 VNB N_A_276_47#_c_415_n 0.00706701f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=0.555
cc_38 VNB N_A_276_47#_c_416_n 0.00584181f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.295
cc_39 VNB N_A_276_47#_c_417_n 0.00299166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_276_47#_c_418_n 0.00322341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_276_47#_c_419_n 9.88026e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_276_47#_c_420_n 0.00902339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_276_47#_c_421_n 0.00701766f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_276_47#_c_422_n 0.00205633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_D_N_M1009_g 0.0346493f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.445
cc_46 VNB D_N 0.012763f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.76
cc_47 VNB N_D_N_c_531_n 0.0323258f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=2.225
cc_48 VNB N_VPWR_c_555_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_X_c_606_n 0.00640576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_627_n 0.00243645f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_51 VNB N_VGND_c_628_n 0.00476851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_629_n 0.016849f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=0.555
cc_53 VNB N_VGND_c_630_n 0.0298283f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=0.925
cc_54 VNB N_VGND_c_631_n 0.00382155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_632_n 0.0109617f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.295
cc_56 VNB N_VGND_c_633_n 0.0154337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_634_n 0.0151002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_635_n 0.00528623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_636_n 0.0204163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_637_n 0.021863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_638_n 0.261548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_639_n 0.00455727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VPB N_C_N_c_106_n 0.00128929f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.685
cc_64 VPB N_C_N_c_112_n 0.018789f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.76
cc_65 VPB N_C_N_c_113_n 0.0127874f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.76
cc_66 VPB N_C_N_M1007_g 0.0262793f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=2.225
cc_67 VPB N_A_M1002_g 0.0285338f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.435
cc_68 VPB N_B_M1004_g 0.0276925f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.445
cc_69 VPB N_A_40_47#_M1012_g 0.0288233f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.76
cc_70 VPB N_A_40_47#_c_236_n 0.0242331f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=0.925
cc_71 VPB N_A_40_47#_c_231_n 0.0266129f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.295
cc_72 VPB N_A_40_47#_c_232_n 0.0167816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_462_351#_c_308_n 0.0180899f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.685
cc_74 VPB N_A_462_351#_c_309_n 0.0160742f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.835
cc_75 VPB N_A_462_351#_c_310_n 0.00619204f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=2.225
cc_76 VPB N_A_462_351#_c_301_n 0.00617721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_A_462_351#_c_312_n 0.0445699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_462_351#_c_313_n 0.0124904f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.93
cc_79 VPB N_A_462_351#_c_314_n 0.0059257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_462_351#_c_315_n 0.0115379f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.295
cc_81 VPB N_A_462_351#_c_316_n 0.00680667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_462_351#_c_304_n 0.00139567f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A_462_351#_c_318_n 0.00344177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_462_351#_c_319_n 0.0270485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A_462_351#_c_320_n 0.0661353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_276_47#_c_411_n 0.0245941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_276_47#_M1013_g 0.0213807f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.93
cc_88 VPB N_A_276_47#_c_419_n 0.00206588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_276_47#_c_426_n 0.00510431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_D_N_M1011_g 0.0305895f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.685
cc_91 VPB D_N 0.00833411f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.76
cc_92 VPB N_D_N_c_531_n 0.00699532f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=2.225
cc_93 VPB N_VPWR_c_556_n 0.0499917f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=2.225
cc_94 VPB N_VPWR_c_557_n 0.00550494f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_95 VPB N_VPWR_c_558_n 0.0148774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_559_n 0.0326924f $X=-0.19 $Y=1.655 $X2=0.652 $Y2=0.765
cc_97 VPB N_VPWR_c_560_n 0.05097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_561_n 0.0127083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_562_n 0.021922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_555_n 0.135208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_564_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_565_n 0.00510584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_566_n 0.00510584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_X_c_606_n 0.00426245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 N_C_N_c_106_n N_A_M1002_g 0.0017234f $X=0.54 $Y=1.685 $X2=0 $Y2=0
cc_106 N_C_N_c_112_n N_A_M1002_g 0.0217489f $X=0.8 $Y=1.76 $X2=0 $Y2=0
cc_107 C_N N_A_c_152_n 0.00149009f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_108 N_C_N_c_109_n N_A_c_152_n 3.32112e-19 $X=0.675 $Y=0.93 $X2=0 $Y2=0
cc_109 N_C_N_c_110_n N_A_c_152_n 0.00630672f $X=0.652 $Y=0.765 $X2=0 $Y2=0
cc_110 N_C_N_c_105_n N_A_c_153_n 0.0138947f $X=0.652 $Y=1.248 $X2=0 $Y2=0
cc_111 N_C_N_c_107_n N_A_c_154_n 0.0138947f $X=0.652 $Y=1.435 $X2=0 $Y2=0
cc_112 C_N A 0.0413757f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_113 N_C_N_c_109_n A 0.00393613f $X=0.675 $Y=0.93 $X2=0 $Y2=0
cc_114 C_N N_A_c_156_n 7.79501e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_115 N_C_N_c_109_n N_A_c_156_n 0.0138947f $X=0.675 $Y=0.93 $X2=0 $Y2=0
cc_116 C_N N_A_40_47#_c_230_n 0.0653428f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_117 N_C_N_c_110_n N_A_40_47#_c_230_n 0.0290706f $X=0.652 $Y=0.765 $X2=0 $Y2=0
cc_118 N_C_N_c_112_n N_A_40_47#_c_236_n 0.00580557f $X=0.8 $Y=1.76 $X2=0 $Y2=0
cc_119 N_C_N_c_113_n N_A_40_47#_c_236_n 0.00512954f $X=0.615 $Y=1.76 $X2=0 $Y2=0
cc_120 N_C_N_M1007_g N_A_40_47#_c_236_n 0.00810347f $X=0.875 $Y=2.225 $X2=0
+ $Y2=0
cc_121 N_C_N_c_112_n N_A_40_47#_c_231_n 0.0117242f $X=0.8 $Y=1.76 $X2=0 $Y2=0
cc_122 N_C_N_c_107_n N_A_40_47#_c_231_n 5.47305e-19 $X=0.652 $Y=1.435 $X2=0
+ $Y2=0
cc_123 N_C_N_c_106_n N_A_40_47#_c_232_n 0.00761331f $X=0.54 $Y=1.685 $X2=0 $Y2=0
cc_124 N_C_N_c_112_n N_A_40_47#_c_232_n 0.00305241f $X=0.8 $Y=1.76 $X2=0 $Y2=0
cc_125 N_C_N_c_113_n N_A_40_47#_c_232_n 0.00526373f $X=0.615 $Y=1.76 $X2=0 $Y2=0
cc_126 N_C_N_c_107_n N_A_40_47#_c_232_n 6.16582e-19 $X=0.652 $Y=1.435 $X2=0
+ $Y2=0
cc_127 C_N N_A_40_47#_c_232_n 0.016948f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_128 C_N N_A_276_47#_c_417_n 0.00475323f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_129 N_C_N_M1007_g N_VPWR_c_556_n 0.00369603f $X=0.875 $Y=2.225 $X2=0 $Y2=0
cc_130 N_C_N_M1007_g N_VPWR_c_559_n 0.00297774f $X=0.875 $Y=2.225 $X2=0 $Y2=0
cc_131 N_C_N_M1007_g N_VPWR_c_555_n 0.00400849f $X=0.875 $Y=2.225 $X2=0 $Y2=0
cc_132 C_N N_VGND_M1003_d 0.00428381f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_133 C_N N_VGND_c_627_n 0.0103712f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_134 N_C_N_c_110_n N_VGND_c_627_n 0.00470553f $X=0.652 $Y=0.765 $X2=0 $Y2=0
cc_135 C_N N_VGND_c_630_n 0.00592215f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_136 N_C_N_c_109_n N_VGND_c_630_n 0.00104552f $X=0.675 $Y=0.93 $X2=0 $Y2=0
cc_137 N_C_N_c_110_n N_VGND_c_630_n 0.00543046f $X=0.652 $Y=0.765 $X2=0 $Y2=0
cc_138 C_N N_VGND_c_638_n 0.00778885f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_139 N_C_N_c_109_n N_VGND_c_638_n 6.86715e-19 $X=0.675 $Y=0.93 $X2=0 $Y2=0
cc_140 N_C_N_c_110_n N_VGND_c_638_n 0.0115225f $X=0.652 $Y=0.765 $X2=0 $Y2=0
cc_141 N_A_c_154_n N_B_M1004_g 0.053995f $X=1.215 $Y=1.445 $X2=0 $Y2=0
cc_142 N_A_c_152_n N_B_M1006_g 0.0165991f $X=1.215 $Y=0.775 $X2=0 $Y2=0
cc_143 A N_B_M1006_g 4.32331e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_144 A N_B_c_192_n 9.19075e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_145 N_A_c_156_n N_B_c_192_n 0.053995f $X=1.215 $Y=0.94 $X2=0 $Y2=0
cc_146 A N_B_c_193_n 0.0380392f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_147 N_A_c_156_n N_B_c_193_n 0.00373464f $X=1.215 $Y=0.94 $X2=0 $Y2=0
cc_148 A N_A_40_47#_c_230_n 3.21901e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_149 N_A_M1002_g N_A_40_47#_c_231_n 0.0167972f $X=1.305 $Y=2.225 $X2=0 $Y2=0
cc_150 N_A_c_154_n N_A_40_47#_c_231_n 0.00123832f $X=1.215 $Y=1.445 $X2=0 $Y2=0
cc_151 A N_A_40_47#_c_231_n 0.02063f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_152 N_A_c_152_n N_A_276_47#_c_417_n 0.00223261f $X=1.215 $Y=0.775 $X2=0 $Y2=0
cc_153 N_A_M1002_g N_VPWR_c_556_n 0.0113489f $X=1.305 $Y=2.225 $X2=0 $Y2=0
cc_154 N_A_M1002_g N_VPWR_c_560_n 0.00247589f $X=1.305 $Y=2.225 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_VPWR_c_555_n 0.00336713f $X=1.305 $Y=2.225 $X2=0 $Y2=0
cc_156 N_A_c_152_n N_VGND_c_627_n 0.00804053f $X=1.215 $Y=0.775 $X2=0 $Y2=0
cc_157 A N_VGND_c_627_n 0.0150424f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_158 N_A_c_156_n N_VGND_c_627_n 0.00123287f $X=1.215 $Y=0.94 $X2=0 $Y2=0
cc_159 N_A_c_152_n N_VGND_c_633_n 0.00525069f $X=1.215 $Y=0.775 $X2=0 $Y2=0
cc_160 N_A_c_152_n N_VGND_c_638_n 0.00689178f $X=1.215 $Y=0.775 $X2=0 $Y2=0
cc_161 A N_VGND_c_638_n 0.00296617f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_162 N_B_M1006_g N_A_40_47#_M1010_g 0.0157474f $X=1.735 $Y=0.445 $X2=0 $Y2=0
cc_163 N_B_c_192_n N_A_40_47#_M1010_g 7.81606e-19 $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_164 N_B_M1004_g N_A_40_47#_c_229_n 0.0808844f $X=1.665 $Y=2.225 $X2=0 $Y2=0
cc_165 N_B_c_193_n N_A_40_47#_c_229_n 0.00220573f $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_166 N_B_M1004_g N_A_40_47#_c_231_n 0.0140641f $X=1.665 $Y=2.225 $X2=0 $Y2=0
cc_167 N_B_c_192_n N_A_40_47#_c_231_n 6.86847e-19 $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_168 N_B_c_193_n N_A_40_47#_c_231_n 0.0333665f $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_169 N_B_M1004_g N_A_40_47#_c_233_n 6.56108e-19 $X=1.665 $Y=2.225 $X2=0 $Y2=0
cc_170 N_B_c_192_n N_A_40_47#_c_233_n 9.0492e-19 $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_171 N_B_c_193_n N_A_40_47#_c_233_n 0.0353262f $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_172 N_B_c_192_n N_A_40_47#_c_234_n 0.0195294f $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_173 N_B_c_193_n N_A_40_47#_c_234_n 9.01708e-19 $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_174 N_B_M1006_g N_A_276_47#_c_416_n 0.0115956f $X=1.735 $Y=0.445 $X2=0 $Y2=0
cc_175 N_B_c_192_n N_A_276_47#_c_416_n 0.00297706f $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_176 N_B_c_193_n N_A_276_47#_c_416_n 0.020476f $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_177 N_B_c_192_n N_A_276_47#_c_417_n 0.00175861f $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_178 N_B_c_193_n N_A_276_47#_c_417_n 0.0131068f $X=1.755 $Y=1.02 $X2=0 $Y2=0
cc_179 N_B_M1006_g N_A_276_47#_c_421_n 8.52336e-19 $X=1.735 $Y=0.445 $X2=0 $Y2=0
cc_180 N_B_M1004_g N_VPWR_c_556_n 0.00261274f $X=1.665 $Y=2.225 $X2=0 $Y2=0
cc_181 N_B_M1004_g N_VPWR_c_560_n 0.00297774f $X=1.665 $Y=2.225 $X2=0 $Y2=0
cc_182 N_B_M1004_g N_VPWR_c_555_n 0.00400849f $X=1.665 $Y=2.225 $X2=0 $Y2=0
cc_183 N_B_M1006_g N_VGND_c_627_n 5.65736e-19 $X=1.735 $Y=0.445 $X2=0 $Y2=0
cc_184 N_B_M1006_g N_VGND_c_632_n 0.00302501f $X=1.735 $Y=0.445 $X2=0 $Y2=0
cc_185 N_B_M1006_g N_VGND_c_633_n 0.00417536f $X=1.735 $Y=0.445 $X2=0 $Y2=0
cc_186 N_B_M1006_g N_VGND_c_638_n 0.00623895f $X=1.735 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A_40_47#_M1012_g N_A_462_351#_c_310_n 0.0518652f $X=2.025 $Y=2.225
+ $X2=0 $Y2=0
cc_188 N_A_40_47#_c_229_n N_A_462_351#_c_310_n 0.00982047f $X=2.295 $Y=1.395
+ $X2=0 $Y2=0
cc_189 N_A_40_47#_c_231_n N_A_462_351#_c_310_n 0.00978967f $X=2.13 $Y=1.71 $X2=0
+ $Y2=0
cc_190 N_A_40_47#_M1012_g N_A_462_351#_c_301_n 0.00300247f $X=2.025 $Y=2.225
+ $X2=0 $Y2=0
cc_191 N_A_40_47#_c_229_n N_A_462_351#_c_301_n 0.0233415f $X=2.295 $Y=1.395
+ $X2=0 $Y2=0
cc_192 N_A_40_47#_c_231_n N_A_462_351#_c_301_n 5.84432e-19 $X=2.13 $Y=1.71 $X2=0
+ $Y2=0
cc_193 N_A_40_47#_c_233_n N_A_462_351#_c_301_n 3.19283e-19 $X=2.295 $Y=1.04
+ $X2=0 $Y2=0
cc_194 N_A_40_47#_M1010_g N_A_462_351#_M1001_g 0.0140423f $X=2.385 $Y=0.445
+ $X2=0 $Y2=0
cc_195 N_A_40_47#_M1010_g N_A_462_351#_c_303_n 0.0233415f $X=2.385 $Y=0.445
+ $X2=0 $Y2=0
cc_196 N_A_40_47#_c_233_n N_A_462_351#_c_303_n 7.4128e-19 $X=2.295 $Y=1.04 $X2=0
+ $Y2=0
cc_197 N_A_40_47#_M1010_g N_A_276_47#_c_416_n 0.00980019f $X=2.385 $Y=0.445
+ $X2=0 $Y2=0
cc_198 N_A_40_47#_c_229_n N_A_276_47#_c_416_n 0.00446188f $X=2.295 $Y=1.395
+ $X2=0 $Y2=0
cc_199 N_A_40_47#_c_233_n N_A_276_47#_c_416_n 0.023826f $X=2.295 $Y=1.04 $X2=0
+ $Y2=0
cc_200 N_A_40_47#_c_234_n N_A_276_47#_c_416_n 0.00496807f $X=2.295 $Y=1.04 $X2=0
+ $Y2=0
cc_201 N_A_40_47#_M1010_g N_A_276_47#_c_418_n 0.00474928f $X=2.385 $Y=0.445
+ $X2=0 $Y2=0
cc_202 N_A_40_47#_c_233_n N_A_276_47#_c_418_n 0.018645f $X=2.295 $Y=1.04 $X2=0
+ $Y2=0
cc_203 N_A_40_47#_M1012_g N_A_276_47#_c_419_n 7.29736e-19 $X=2.025 $Y=2.225
+ $X2=0 $Y2=0
cc_204 N_A_40_47#_c_231_n N_A_276_47#_c_419_n 0.0134511f $X=2.13 $Y=1.71 $X2=0
+ $Y2=0
cc_205 N_A_40_47#_c_233_n N_A_276_47#_c_419_n 0.00817468f $X=2.295 $Y=1.04 $X2=0
+ $Y2=0
cc_206 N_A_40_47#_M1010_g N_A_276_47#_c_421_n 0.0081622f $X=2.385 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_40_47#_c_233_n N_A_276_47#_c_421_n 0.00189525f $X=2.295 $Y=1.04 $X2=0
+ $Y2=0
cc_208 N_A_40_47#_M1012_g N_A_276_47#_c_426_n 0.00139428f $X=2.025 $Y=2.225
+ $X2=0 $Y2=0
cc_209 N_A_40_47#_c_231_n N_A_276_47#_c_426_n 0.00173035f $X=2.13 $Y=1.71 $X2=0
+ $Y2=0
cc_210 N_A_40_47#_c_229_n N_A_276_47#_c_422_n 0.00204519f $X=2.295 $Y=1.395
+ $X2=0 $Y2=0
cc_211 N_A_40_47#_c_233_n N_A_276_47#_c_422_n 0.0264882f $X=2.295 $Y=1.04 $X2=0
+ $Y2=0
cc_212 N_A_40_47#_c_231_n N_VPWR_c_556_n 0.0146725f $X=2.13 $Y=1.71 $X2=0 $Y2=0
cc_213 N_A_40_47#_M1012_g N_VPWR_c_560_n 0.00297774f $X=2.025 $Y=2.225 $X2=0
+ $Y2=0
cc_214 N_A_40_47#_M1012_g N_VPWR_c_555_n 0.00400849f $X=2.025 $Y=2.225 $X2=0
+ $Y2=0
cc_215 N_A_40_47#_c_230_n N_VGND_c_630_n 0.0150394f $X=0.325 $Y=0.445 $X2=0
+ $Y2=0
cc_216 N_A_40_47#_M1010_g N_VGND_c_632_n 0.00530547f $X=2.385 $Y=0.445 $X2=0
+ $Y2=0
cc_217 N_A_40_47#_M1010_g N_VGND_c_636_n 0.00409905f $X=2.385 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_A_40_47#_M1003_s N_VGND_c_638_n 0.00411505f $X=0.2 $Y=0.235 $X2=0 $Y2=0
cc_219 N_A_40_47#_M1010_g N_VGND_c_638_n 0.00634624f $X=2.385 $Y=0.445 $X2=0
+ $Y2=0
cc_220 N_A_40_47#_c_230_n N_VGND_c_638_n 0.00951889f $X=0.325 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_462_351#_c_301_n N_A_276_47#_c_410_n 0.00432275f $X=2.745 $Y=1.755
+ $X2=0 $Y2=0
cc_222 N_A_462_351#_M1001_g N_A_276_47#_c_410_n 0.0143626f $X=2.815 $Y=0.445
+ $X2=0 $Y2=0
cc_223 N_A_462_351#_c_301_n N_A_276_47#_c_411_n 0.0270348f $X=2.745 $Y=1.755
+ $X2=0 $Y2=0
cc_224 N_A_462_351#_c_313_n N_A_276_47#_c_411_n 0.0419806f $X=2.875 $Y=1.83
+ $X2=0 $Y2=0
cc_225 N_A_462_351#_c_314_n N_A_276_47#_c_411_n 5.72737e-19 $X=2.64 $Y=2.94
+ $X2=0 $Y2=0
cc_226 N_A_462_351#_c_315_n N_A_276_47#_c_411_n 0.0167618f $X=3.865 $Y=2.53
+ $X2=0 $Y2=0
cc_227 N_A_462_351#_c_318_n N_A_276_47#_c_411_n 7.37073e-19 $X=4.035 $Y=2.445
+ $X2=0 $Y2=0
cc_228 N_A_462_351#_c_306_n N_A_276_47#_c_413_n 0.00112337f $X=4.035 $Y=1.15
+ $X2=0 $Y2=0
cc_229 N_A_462_351#_c_307_n N_A_276_47#_c_413_n 5.05935e-19 $X=4.5 $Y=0.865
+ $X2=0 $Y2=0
cc_230 N_A_462_351#_c_315_n N_A_276_47#_M1013_g 0.0176208f $X=3.865 $Y=2.53
+ $X2=0 $Y2=0
cc_231 N_A_462_351#_c_304_n N_A_276_47#_M1013_g 0.0107949f $X=3.95 $Y=1.93 $X2=0
+ $Y2=0
cc_232 N_A_462_351#_c_318_n N_A_276_47#_M1013_g 0.00580816f $X=4.035 $Y=2.445
+ $X2=0 $Y2=0
cc_233 N_A_462_351#_c_343_p N_A_276_47#_M1013_g 0.00775485f $X=4.035 $Y=2.095
+ $X2=0 $Y2=0
cc_234 N_A_462_351#_c_304_n N_A_276_47#_c_415_n 0.00229108f $X=3.95 $Y=1.93
+ $X2=0 $Y2=0
cc_235 N_A_462_351#_c_306_n N_A_276_47#_c_415_n 0.00151582f $X=4.035 $Y=1.15
+ $X2=0 $Y2=0
cc_236 N_A_462_351#_c_301_n N_A_276_47#_c_418_n 0.00639506f $X=2.745 $Y=1.755
+ $X2=0 $Y2=0
cc_237 N_A_462_351#_M1001_g N_A_276_47#_c_418_n 7.3836e-19 $X=2.815 $Y=0.445
+ $X2=0 $Y2=0
cc_238 N_A_462_351#_c_303_n N_A_276_47#_c_418_n 0.00489486f $X=2.78 $Y=0.945
+ $X2=0 $Y2=0
cc_239 N_A_462_351#_c_308_n N_A_276_47#_c_419_n 0.0030315f $X=2.385 $Y=1.905
+ $X2=0 $Y2=0
cc_240 N_A_462_351#_c_309_n N_A_276_47#_c_419_n 0.00399575f $X=2.67 $Y=1.83
+ $X2=0 $Y2=0
cc_241 N_A_462_351#_c_301_n N_A_276_47#_c_419_n 0.0085136f $X=2.745 $Y=1.755
+ $X2=0 $Y2=0
cc_242 N_A_462_351#_c_312_n N_A_276_47#_c_419_n 0.00166753f $X=2.875 $Y=2.775
+ $X2=0 $Y2=0
cc_243 N_A_462_351#_c_313_n N_A_276_47#_c_419_n 0.00526037f $X=2.875 $Y=1.83
+ $X2=0 $Y2=0
cc_244 N_A_462_351#_c_301_n N_A_276_47#_c_420_n 0.00407557f $X=2.745 $Y=1.755
+ $X2=0 $Y2=0
cc_245 N_A_462_351#_c_303_n N_A_276_47#_c_420_n 0.00288063f $X=2.78 $Y=0.945
+ $X2=0 $Y2=0
cc_246 N_A_462_351#_c_313_n N_A_276_47#_c_420_n 0.00534975f $X=2.875 $Y=1.83
+ $X2=0 $Y2=0
cc_247 N_A_462_351#_M1001_g N_A_276_47#_c_421_n 0.00830045f $X=2.815 $Y=0.445
+ $X2=0 $Y2=0
cc_248 N_A_462_351#_c_308_n N_A_276_47#_c_426_n 0.00650489f $X=2.385 $Y=1.905
+ $X2=0 $Y2=0
cc_249 N_A_462_351#_c_309_n N_A_276_47#_c_426_n 0.00407568f $X=2.67 $Y=1.83
+ $X2=0 $Y2=0
cc_250 N_A_462_351#_c_312_n N_A_276_47#_c_426_n 0.00915797f $X=2.875 $Y=2.775
+ $X2=0 $Y2=0
cc_251 N_A_462_351#_c_315_n N_A_276_47#_c_426_n 2.8192e-19 $X=3.865 $Y=2.53
+ $X2=0 $Y2=0
cc_252 N_A_462_351#_c_316_n N_A_276_47#_c_426_n 0.0266162f $X=2.805 $Y=2.53
+ $X2=0 $Y2=0
cc_253 N_A_462_351#_c_320_n N_A_276_47#_c_426_n 0.00111493f $X=2.875 $Y=2.94
+ $X2=0 $Y2=0
cc_254 N_A_462_351#_c_301_n N_A_276_47#_c_422_n 0.00505914f $X=2.745 $Y=1.755
+ $X2=0 $Y2=0
cc_255 N_A_462_351#_c_304_n N_D_N_M1009_g 0.00552905f $X=3.95 $Y=1.93 $X2=0
+ $Y2=0
cc_256 N_A_462_351#_c_305_n N_D_N_M1009_g 0.0154196f $X=4.335 $Y=1.15 $X2=0
+ $Y2=0
cc_257 N_A_462_351#_c_307_n N_D_N_M1009_g 0.0058872f $X=4.5 $Y=0.865 $X2=0 $Y2=0
cc_258 N_A_462_351#_c_304_n N_D_N_M1011_g 0.00377566f $X=3.95 $Y=1.93 $X2=0
+ $Y2=0
cc_259 N_A_462_351#_c_318_n N_D_N_M1011_g 0.00360439f $X=4.035 $Y=2.445 $X2=0
+ $Y2=0
cc_260 N_A_462_351#_c_319_n N_D_N_M1011_g 0.0177558f $X=4.535 $Y=2.055 $X2=0
+ $Y2=0
cc_261 N_A_462_351#_c_304_n D_N 0.0267291f $X=3.95 $Y=1.93 $X2=0 $Y2=0
cc_262 N_A_462_351#_c_305_n D_N 0.0364039f $X=4.335 $Y=1.15 $X2=0 $Y2=0
cc_263 N_A_462_351#_c_319_n D_N 0.0353923f $X=4.535 $Y=2.055 $X2=0 $Y2=0
cc_264 N_A_462_351#_c_305_n N_D_N_c_531_n 0.00474042f $X=4.335 $Y=1.15 $X2=0
+ $Y2=0
cc_265 N_A_462_351#_c_319_n N_D_N_c_531_n 7.69561e-19 $X=4.535 $Y=2.055 $X2=0
+ $Y2=0
cc_266 N_A_462_351#_c_315_n N_VPWR_M1005_s 0.0100895f $X=3.865 $Y=2.53 $X2=0
+ $Y2=0
cc_267 N_A_462_351#_c_315_n N_VPWR_M1013_s 0.00303057f $X=3.865 $Y=2.53 $X2=0
+ $Y2=0
cc_268 N_A_462_351#_c_304_n N_VPWR_M1013_s 0.00112177f $X=3.95 $Y=1.93 $X2=0
+ $Y2=0
cc_269 N_A_462_351#_c_343_p N_VPWR_M1013_s 0.00718195f $X=4.035 $Y=2.095 $X2=0
+ $Y2=0
cc_270 N_A_462_351#_c_314_n N_VPWR_c_557_n 0.0219818f $X=2.64 $Y=2.94 $X2=0
+ $Y2=0
cc_271 N_A_462_351#_c_315_n N_VPWR_c_557_n 0.0210984f $X=3.865 $Y=2.53 $X2=0
+ $Y2=0
cc_272 N_A_462_351#_c_320_n N_VPWR_c_557_n 0.003772f $X=2.875 $Y=2.94 $X2=0
+ $Y2=0
cc_273 N_A_462_351#_c_315_n N_VPWR_c_558_n 0.0230659f $X=3.865 $Y=2.53 $X2=0
+ $Y2=0
cc_274 N_A_462_351#_c_308_n N_VPWR_c_560_n 0.00297774f $X=2.385 $Y=1.905 $X2=0
+ $Y2=0
cc_275 N_A_462_351#_c_314_n N_VPWR_c_560_n 0.0222366f $X=2.64 $Y=2.94 $X2=0
+ $Y2=0
cc_276 N_A_462_351#_c_315_n N_VPWR_c_560_n 0.00250852f $X=3.865 $Y=2.53 $X2=0
+ $Y2=0
cc_277 N_A_462_351#_c_320_n N_VPWR_c_560_n 0.0091353f $X=2.875 $Y=2.94 $X2=0
+ $Y2=0
cc_278 N_A_462_351#_c_315_n N_VPWR_c_561_n 0.0067515f $X=3.865 $Y=2.53 $X2=0
+ $Y2=0
cc_279 N_A_462_351#_c_315_n N_VPWR_c_562_n 5.11315e-19 $X=3.865 $Y=2.53 $X2=0
+ $Y2=0
cc_280 N_A_462_351#_c_308_n N_VPWR_c_555_n 0.00400849f $X=2.385 $Y=1.905 $X2=0
+ $Y2=0
cc_281 N_A_462_351#_c_314_n N_VPWR_c_555_n 0.0112257f $X=2.64 $Y=2.94 $X2=0
+ $Y2=0
cc_282 N_A_462_351#_c_315_n N_VPWR_c_555_n 0.0207904f $X=3.865 $Y=2.53 $X2=0
+ $Y2=0
cc_283 N_A_462_351#_c_320_n N_VPWR_c_555_n 0.0120503f $X=2.875 $Y=2.94 $X2=0
+ $Y2=0
cc_284 N_A_462_351#_c_315_n N_X_M1005_d 0.00491577f $X=3.865 $Y=2.53 $X2=0 $Y2=0
cc_285 N_A_462_351#_c_315_n N_X_c_606_n 0.0135055f $X=3.865 $Y=2.53 $X2=0 $Y2=0
cc_286 N_A_462_351#_c_304_n N_X_c_606_n 0.0468819f $X=3.95 $Y=1.93 $X2=0 $Y2=0
cc_287 N_A_462_351#_c_306_n N_X_c_606_n 0.0132748f $X=4.035 $Y=1.15 $X2=0 $Y2=0
cc_288 N_A_462_351#_c_307_n N_X_c_606_n 0.00412477f $X=4.5 $Y=0.865 $X2=0 $Y2=0
cc_289 N_A_462_351#_c_305_n N_VGND_M1014_d 0.00162909f $X=4.335 $Y=1.15 $X2=0
+ $Y2=0
cc_290 N_A_462_351#_c_306_n N_VGND_M1014_d 0.00158247f $X=4.035 $Y=1.15 $X2=0
+ $Y2=0
cc_291 N_A_462_351#_c_301_n N_VGND_c_628_n 5.22849e-19 $X=2.745 $Y=1.755 $X2=0
+ $Y2=0
cc_292 N_A_462_351#_M1001_g N_VGND_c_628_n 0.00916688f $X=2.815 $Y=0.445 $X2=0
+ $Y2=0
cc_293 N_A_462_351#_c_305_n N_VGND_c_629_n 0.00842481f $X=4.335 $Y=1.15 $X2=0
+ $Y2=0
cc_294 N_A_462_351#_c_306_n N_VGND_c_629_n 0.0128931f $X=4.035 $Y=1.15 $X2=0
+ $Y2=0
cc_295 N_A_462_351#_c_307_n N_VGND_c_629_n 0.013429f $X=4.5 $Y=0.865 $X2=0 $Y2=0
cc_296 N_A_462_351#_M1001_g N_VGND_c_636_n 0.00483021f $X=2.815 $Y=0.445 $X2=0
+ $Y2=0
cc_297 N_A_462_351#_c_307_n N_VGND_c_637_n 0.00495237f $X=4.5 $Y=0.865 $X2=0
+ $Y2=0
cc_298 N_A_462_351#_M1001_g N_VGND_c_638_n 0.00866235f $X=2.815 $Y=0.445 $X2=0
+ $Y2=0
cc_299 N_A_462_351#_c_307_n N_VGND_c_638_n 0.00933518f $X=4.5 $Y=0.865 $X2=0
+ $Y2=0
cc_300 N_A_276_47#_c_413_n N_D_N_M1009_g 0.0118302f $X=3.76 $Y=1.185 $X2=0 $Y2=0
cc_301 N_A_276_47#_c_415_n N_D_N_M1009_g 0.00802494f $X=3.777 $Y=1.26 $X2=0
+ $Y2=0
cc_302 N_A_276_47#_M1013_g N_D_N_M1011_g 0.0205588f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_276_47#_M1013_g D_N 5.02724e-19 $X=3.795 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A_276_47#_M1013_g N_D_N_c_531_n 0.00802494f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_A_276_47#_c_411_n N_VPWR_c_557_n 0.0104937f $X=3.365 $Y=1.725 $X2=0
+ $Y2=0
cc_306 N_A_276_47#_M1013_g N_VPWR_c_557_n 0.00133982f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_276_47#_c_411_n N_VPWR_c_558_n 0.00133982f $X=3.365 $Y=1.725 $X2=0
+ $Y2=0
cc_308 N_A_276_47#_M1013_g N_VPWR_c_558_n 0.0106038f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_276_47#_c_411_n N_VPWR_c_561_n 0.00362954f $X=3.365 $Y=1.725 $X2=0
+ $Y2=0
cc_310 N_A_276_47#_M1013_g N_VPWR_c_561_n 0.00362954f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A_276_47#_c_411_n N_VPWR_c_555_n 0.00435695f $X=3.365 $Y=1.725 $X2=0
+ $Y2=0
cc_312 N_A_276_47#_M1013_g N_VPWR_c_555_n 0.00435695f $X=3.795 $Y=2.465 $X2=0
+ $Y2=0
cc_313 N_A_276_47#_c_410_n N_X_c_606_n 0.00201477f $X=3.33 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A_276_47#_c_411_n N_X_c_606_n 0.00670408f $X=3.365 $Y=1.725 $X2=0 $Y2=0
cc_315 N_A_276_47#_c_412_n N_X_c_606_n 0.0109951f $X=3.685 $Y=1.26 $X2=0 $Y2=0
cc_316 N_A_276_47#_c_413_n N_X_c_606_n 0.0124653f $X=3.76 $Y=1.185 $X2=0 $Y2=0
cc_317 N_A_276_47#_M1013_g N_X_c_606_n 0.00431806f $X=3.795 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A_276_47#_c_415_n N_X_c_606_n 0.00210532f $X=3.777 $Y=1.26 $X2=0 $Y2=0
cc_319 N_A_276_47#_c_418_n N_X_c_606_n 0.00358746f $X=2.725 $Y=1.185 $X2=0 $Y2=0
cc_320 N_A_276_47#_c_419_n N_X_c_606_n 0.0103003f $X=2.725 $Y=1.995 $X2=0 $Y2=0
cc_321 N_A_276_47#_c_420_n N_X_c_606_n 0.0262053f $X=3.195 $Y=1.35 $X2=0 $Y2=0
cc_322 N_A_276_47#_c_416_n N_VGND_M1006_d 0.00479128f $X=2.435 $Y=0.67 $X2=0
+ $Y2=0
cc_323 N_A_276_47#_c_417_n N_VGND_c_627_n 6.3314e-19 $X=1.65 $Y=0.67 $X2=0 $Y2=0
cc_324 N_A_276_47#_c_410_n N_VGND_c_628_n 0.0130558f $X=3.33 $Y=1.185 $X2=0
+ $Y2=0
cc_325 N_A_276_47#_c_411_n N_VGND_c_628_n 0.00506784f $X=3.365 $Y=1.725 $X2=0
+ $Y2=0
cc_326 N_A_276_47#_c_413_n N_VGND_c_628_n 7.39791e-19 $X=3.76 $Y=1.185 $X2=0
+ $Y2=0
cc_327 N_A_276_47#_c_420_n N_VGND_c_628_n 0.0221599f $X=3.195 $Y=1.35 $X2=0
+ $Y2=0
cc_328 N_A_276_47#_c_421_n N_VGND_c_628_n 0.0564761f $X=2.6 $Y=0.445 $X2=0 $Y2=0
cc_329 N_A_276_47#_c_413_n N_VGND_c_629_n 0.00327135f $X=3.76 $Y=1.185 $X2=0
+ $Y2=0
cc_330 N_A_276_47#_c_416_n N_VGND_c_632_n 0.024516f $X=2.435 $Y=0.67 $X2=0 $Y2=0
cc_331 N_A_276_47#_c_421_n N_VGND_c_632_n 0.00811879f $X=2.6 $Y=0.445 $X2=0
+ $Y2=0
cc_332 N_A_276_47#_c_516_p N_VGND_c_633_n 0.012879f $X=1.52 $Y=0.43 $X2=0 $Y2=0
cc_333 N_A_276_47#_c_416_n N_VGND_c_633_n 0.00347982f $X=2.435 $Y=0.67 $X2=0
+ $Y2=0
cc_334 N_A_276_47#_c_410_n N_VGND_c_634_n 0.00486043f $X=3.33 $Y=1.185 $X2=0
+ $Y2=0
cc_335 N_A_276_47#_c_413_n N_VGND_c_634_n 0.00571722f $X=3.76 $Y=1.185 $X2=0
+ $Y2=0
cc_336 N_A_276_47#_c_416_n N_VGND_c_636_n 0.00407273f $X=2.435 $Y=0.67 $X2=0
+ $Y2=0
cc_337 N_A_276_47#_c_421_n N_VGND_c_636_n 0.0187435f $X=2.6 $Y=0.445 $X2=0 $Y2=0
cc_338 N_A_276_47#_M1000_d N_VGND_c_638_n 0.00347322f $X=1.38 $Y=0.235 $X2=0
+ $Y2=0
cc_339 N_A_276_47#_M1010_d N_VGND_c_638_n 0.00226149f $X=2.46 $Y=0.235 $X2=0
+ $Y2=0
cc_340 N_A_276_47#_c_410_n N_VGND_c_638_n 0.00824727f $X=3.33 $Y=1.185 $X2=0
+ $Y2=0
cc_341 N_A_276_47#_c_413_n N_VGND_c_638_n 0.0115803f $X=3.76 $Y=1.185 $X2=0
+ $Y2=0
cc_342 N_A_276_47#_c_516_p N_VGND_c_638_n 0.0089129f $X=1.52 $Y=0.43 $X2=0 $Y2=0
cc_343 N_A_276_47#_c_416_n N_VGND_c_638_n 0.0137342f $X=2.435 $Y=0.67 $X2=0
+ $Y2=0
cc_344 N_A_276_47#_c_421_n N_VGND_c_638_n 0.0137942f $X=2.6 $Y=0.445 $X2=0 $Y2=0
cc_345 N_D_N_M1009_g N_X_c_606_n 7.31097e-19 $X=4.285 $Y=0.865 $X2=0 $Y2=0
cc_346 N_D_N_M1009_g N_VGND_c_629_n 0.00638834f $X=4.285 $Y=0.865 $X2=0 $Y2=0
cc_347 N_D_N_M1009_g N_VGND_c_637_n 0.00385987f $X=4.285 $Y=0.865 $X2=0 $Y2=0
cc_348 N_D_N_M1009_g N_VGND_c_638_n 0.0046122f $X=4.285 $Y=0.865 $X2=0 $Y2=0
cc_349 N_VPWR_c_555_n N_X_M1005_d 0.00358487f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_350 N_X_c_606_n N_VGND_c_634_n 0.0146655f $X=3.545 $Y=0.42 $X2=0 $Y2=0
cc_351 N_X_M1008_s N_VGND_c_638_n 0.00380103f $X=3.405 $Y=0.235 $X2=0 $Y2=0
cc_352 N_X_c_606_n N_VGND_c_638_n 0.00933292f $X=3.545 $Y=0.42 $X2=0 $Y2=0
