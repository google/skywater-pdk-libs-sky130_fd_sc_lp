* File: sky130_fd_sc_lp__a32o_0.pex.spice
* Created: Wed Sep  2 09:27:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32O_0%A_80_21# 1 2 9 15 17 18 21 22 24 25 26 27 32
+ 40 41
c99 21 0 6.57343e-20 $X=0.59 $Y=1.45
c100 18 0 1.44493e-19 $X=0.657 $Y=1.995
r101 40 41 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.037 $Y=1.785
+ $X2=3.037 $Y2=1.955
r102 34 40 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=3.17 $Y=0.61
+ $X2=3.17 $Y2=1.785
r103 32 41 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.985 $Y=2.27
+ $X2=2.985 $Y2=1.955
r104 27 29 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.85 $Y=0.445
+ $X2=2.465 $Y2=0.445
r105 26 34 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.085 $Y=0.445
+ $X2=3.17 $Y2=0.61
r106 26 29 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=3.085 $Y=0.445
+ $X2=2.465 $Y2=0.445
r107 24 27 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=1.722 $Y=0.76
+ $X2=1.722 $Y2=0.445
r108 24 25 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.595 $Y=0.76
+ $X2=0.755 $Y2=0.76
r109 22 43 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.45
+ $X2=0.577 $Y2=1.285
r110 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.45 $X2=0.59 $Y2=1.45
r111 19 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.63 $Y=0.845
+ $X2=0.755 $Y2=0.76
r112 19 21 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=0.63 $Y=0.845
+ $X2=0.63 $Y2=1.45
r113 17 18 44.0658 $w=3.55e-07 $l=1.5e-07 $layer=POLY_cond $X=0.657 $Y=1.845
+ $X2=0.657 $Y2=1.995
r114 15 18 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.84 $Y=2.465 $X2=0.84
+ $Y2=1.995
r115 11 22 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.577 $Y=1.462
+ $X2=0.577 $Y2=1.45
r116 11 17 62.2555 $w=3.55e-07 $l=3.83e-07 $layer=POLY_cond $X=0.577 $Y=1.462
+ $X2=0.577 $Y2=1.845
r117 9 43 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=1.285
r118 2 32 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.845
+ $Y=2.145 $X2=2.985 $Y2=2.27
r119 1 29 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.235 $X2=2.465 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_0%A3 2 5 9 11 12 13 17 18
c51 18 0 2.80382e-20 $X=1.13 $Y=1.1
c52 13 0 1.44493e-19 $X=1.2 $Y=1.665
c53 11 0 6.57343e-20 $X=1.17 $Y=1.605
r54 17 19 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.1
+ $X2=1.17 $Y2=0.935
r55 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.13 $Y=1.1
+ $X2=1.13 $Y2=1.1
r56 13 20 3.54909 $w=3.85e-07 $l=1.12e-07 $layer=LI1_cond $X=1.157 $Y=1.665
+ $X2=1.157 $Y2=1.553
r57 12 20 7.72286 $w=3.83e-07 $l=2.58e-07 $layer=LI1_cond $X=1.157 $Y=1.295
+ $X2=1.157 $Y2=1.553
r58 12 18 5.83705 $w=3.83e-07 $l=1.95e-07 $layer=LI1_cond $X=1.157 $Y=1.295
+ $X2=1.157 $Y2=1.1
r59 9 19 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.3 $Y=0.445 $X2=1.3
+ $Y2=0.935
r60 5 11 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.27 $Y=2.465
+ $X2=1.27 $Y2=1.605
r61 2 11 46.9225 $w=4.1e-07 $l=2.05e-07 $layer=POLY_cond $X=1.17 $Y=1.4 $X2=1.17
+ $Y2=1.605
r62 1 17 5.42589 $w=4.1e-07 $l=4e-08 $layer=POLY_cond $X=1.17 $Y=1.14 $X2=1.17
+ $Y2=1.1
r63 1 2 35.2683 $w=4.1e-07 $l=2.6e-07 $layer=POLY_cond $X=1.17 $Y=1.14 $X2=1.17
+ $Y2=1.4
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_0%A2 3 7 11 12 13 16 17
c52 7 0 1.38141e-20 $X=1.795 $Y=2.465
r53 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.75
+ $Y=1.18 $X2=1.75 $Y2=1.18
r54 13 17 1.24963 $w=6.68e-07 $l=7e-08 $layer=LI1_cond $X=1.68 $Y=1.35 $X2=1.75
+ $Y2=1.35
r55 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.75 $Y=1.52
+ $X2=1.75 $Y2=1.18
r56 11 12 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.52
+ $X2=1.75 $Y2=1.685
r57 10 16 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.015
+ $X2=1.75 $Y2=1.18
r58 7 12 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.795 $Y=2.465
+ $X2=1.795 $Y2=1.685
r59 3 10 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.74 $Y=0.445
+ $X2=1.74 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_0%A1 3 7 11 12 13 14 18
c41 13 0 2.01831e-19 $X=2.16 $Y=0.925
c42 3 0 1.83092e-19 $X=2.2 $Y=0.445
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.005 $X2=2.29 $Y2=1.005
r44 14 19 9.41432 $w=3.53e-07 $l=2.9e-07 $layer=LI1_cond $X=2.197 $Y=1.295
+ $X2=2.197 $Y2=1.005
r45 13 19 2.59705 $w=3.53e-07 $l=8e-08 $layer=LI1_cond $X=2.197 $Y=0.925
+ $X2=2.197 $Y2=1.005
r46 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.29 $Y=1.345
+ $X2=2.29 $Y2=1.005
r47 11 12 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.345
+ $X2=2.29 $Y2=1.51
r48 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=0.84
+ $X2=2.29 $Y2=1.005
r49 7 12 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=2.32 $Y=2.465
+ $X2=2.32 $Y2=1.51
r50 3 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.2 $Y=0.445 $X2=2.2
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_0%B1 3 7 11 12 13 14 18
c40 13 0 1.83092e-19 $X=2.64 $Y=0.925
c41 7 0 3.11233e-20 $X=2.77 $Y=2.465
c42 3 0 1.73793e-19 $X=2.74 $Y=0.445
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.83
+ $Y=1.005 $X2=2.83 $Y2=1.005
r44 14 19 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.73 $Y=1.295
+ $X2=2.73 $Y2=1.005
r45 13 19 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=2.73 $Y=0.925 $X2=2.73
+ $Y2=1.005
r46 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.83 $Y=1.345
+ $X2=2.83 $Y2=1.005
r47 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.345
+ $X2=2.83 $Y2=1.51
r48 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=0.84
+ $X2=2.83 $Y2=1.005
r49 7 12 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=2.77 $Y=2.465
+ $X2=2.77 $Y2=1.51
r50 3 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.74 $Y=0.445
+ $X2=2.74 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_0%B2 1 3 7 15 17 18 19 24
c35 17 0 3.11233e-20 $X=3.6 $Y=0.925
r36 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.12 $X2=3.57 $Y2=1.12
r37 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.59 $Y=1.295
+ $X2=3.59 $Y2=1.665
r38 18 25 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=3.59 $Y=1.295
+ $X2=3.59 $Y2=1.12
r39 17 25 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.59 $Y=0.925
+ $X2=3.59 $Y2=1.12
r40 15 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.57 $Y=1.105
+ $X2=3.57 $Y2=1.12
r41 12 15 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.28 $Y=1.03
+ $X2=3.57 $Y2=1.03
r42 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.57 $Y=1.46
+ $X2=3.57 $Y2=1.12
r43 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.28 $Y=0.955
+ $X2=3.28 $Y2=1.03
r44 5 7 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.28 $Y=0.955 $X2=3.28
+ $Y2=0.445
r45 1 11 79.2622 $w=2.25e-07 $l=5.96992e-07 $layer=POLY_cond $X=3.2 $Y=1.9
+ $X2=3.57 $Y2=1.46
r46 1 3 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.2 $Y=1.9 $X2=3.2
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_0%X 1 2 7 8 9 10 11 12 13 34 38 41
r17 41 42 7.86913 $w=6.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.42 $Y=2.29
+ $X2=0.42 $Y2=2.125
r18 38 39 1.36218 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=0.555 $X2=0.22
+ $Y2=0.585
r19 12 13 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.42 $Y=2.405
+ $X2=0.42 $Y2=2.775
r20 12 41 2.05297 $w=6.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.42 $Y=2.405
+ $X2=0.42 $Y2=2.29
r21 11 42 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.21 $Y=2.035 $X2=0.21
+ $Y2=2.125
r22 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=2.035
r23 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.295
+ $X2=0.21 $Y2=1.665
r24 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=0.925 $X2=0.21
+ $Y2=1.295
r25 7 38 1.19513 $w=2.68e-07 $l=2.8e-08 $layer=LI1_cond $X=0.22 $Y=0.527
+ $X2=0.22 $Y2=0.555
r26 7 34 4.56709 $w=2.68e-07 $l=1.07e-07 $layer=LI1_cond $X=0.22 $Y=0.527
+ $X2=0.22 $Y2=0.42
r27 7 8 14.4286 $w=2.48e-07 $l=3.13e-07 $layer=LI1_cond $X=0.21 $Y=0.612
+ $X2=0.21 $Y2=0.925
r28 7 39 1.24464 $w=2.48e-07 $l=2.7e-08 $layer=LI1_cond $X=0.21 $Y=0.612
+ $X2=0.21 $Y2=0.585
r29 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.5
+ $Y=2.145 $X2=0.625 $Y2=2.29
r30 1 34 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_0%VPWR 1 2 9 13 16 17 18 24 30 31 34
r41 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 31 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.03 $Y2=3.33
r45 28 30 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=3.6 $Y2=3.33
r46 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=2.03 $Y2=3.33
r48 24 26 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 18 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 16 21 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 16 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.065 $Y2=3.33
r55 15 26 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 15 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=1.065 $Y2=3.33
r57 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=3.33
r58 11 13 33.351 $w=3.28e-07 $l=9.55e-07 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=2.29
r59 7 17 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=3.245
+ $X2=1.065 $Y2=3.33
r60 7 9 39.3065 $w=2.78e-07 $l=9.55e-07 $layer=LI1_cond $X=1.065 $Y=3.245
+ $X2=1.065 $Y2=2.29
r61 2 13 300 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=2 $X=1.87
+ $Y=2.145 $X2=2.03 $Y2=2.29
r62 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=2.145 $X2=1.055 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_0%A_269_429# 1 2 3 12 14 15 19 20 21 24
c44 21 0 1.38141e-20 $X=2.65 $Y=2.98
r45 22 24 24.901 $w=2.78e-07 $l=6.05e-07 $layer=LI1_cond $X=3.46 $Y=2.895
+ $X2=3.46 $Y2=2.29
r46 20 22 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.32 $Y=2.98
+ $X2=3.46 $Y2=2.895
r47 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.32 $Y=2.98
+ $X2=2.65 $Y2=2.98
r48 17 21 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=2.507 $Y=2.895
+ $X2=2.65 $Y2=2.98
r49 17 19 24.4641 $w=2.83e-07 $l=6.05e-07 $layer=LI1_cond $X=2.507 $Y=2.895
+ $X2=2.507 $Y2=2.29
r50 16 19 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=2.507 $Y=2.035
+ $X2=2.507 $Y2=2.29
r51 14 16 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=2.365 $Y=1.95
+ $X2=2.507 $Y2=2.035
r52 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.365 $Y=1.95
+ $X2=1.695 $Y2=1.95
r53 10 15 20.7559 $w=9e-08 $l=1.9799e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.695 $Y2=1.95
r54 10 12 9.18353 $w=3.18e-07 $l=2.55e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.535 $Y2=2.29
r55 3 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.275
+ $Y=2.145 $X2=3.415 $Y2=2.29
r56 2 19 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.395
+ $Y=2.145 $X2=2.535 $Y2=2.29
r57 1 12 300 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=2 $X=1.345
+ $Y=2.145 $X2=1.54 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_0%VGND 1 2 7 9 11 18 26 32 35
r44 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 30 32 7.75958 $w=5.88e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=0.21 $X2=1.25
+ $Y2=0.21
r46 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r47 28 30 2.33134 $w=5.88e-07 $l=1.15e-07 $layer=LI1_cond $X=1.085 $Y=0.21
+ $X2=1.2 $Y2=0.21
r48 25 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r49 24 28 7.39947 $w=5.88e-07 $l=3.65e-07 $layer=LI1_cond $X=0.72 $Y=0.21
+ $X2=1.085 $Y2=0.21
r50 24 26 10.6991 $w=5.88e-07 $l=1.95e-07 $layer=LI1_cond $X=0.72 $Y=0.21
+ $X2=0.525 $Y2=0.21
r51 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 22 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r53 21 32 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=1.25
+ $Y2=0
r54 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r55 18 34 3.95357 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.632
+ $Y2=0
r56 18 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=0 $X2=3.12
+ $Y2=0
r57 16 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r58 15 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.525
+ $Y2=0
r59 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r60 11 22 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r61 11 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r62 7 34 3.18959 $w=2.5e-07 $l=1.19143e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.632 $Y2=0
r63 7 9 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=3.55 $Y=0.085 $X2=3.55
+ $Y2=0.445
r64 2 9 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=3.355
+ $Y=0.235 $X2=3.51 $Y2=0.445
r65 1 28 91 $w=1.7e-07 $l=6.07577e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=1.085 $Y2=0.39
.ends

