* File: sky130_fd_sc_lp__dlygate4s18_1.pex.spice
* Created: Wed Sep  2 09:50:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLYGATE4S18_1%A 3 7 11 12 13 14 18
r37 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.565
+ $Y=1.355 $X2=0.565 $Y2=1.355
r38 14 19 5.88547 $w=6.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.415 $Y=1.665
+ $X2=0.415 $Y2=1.355
r39 13 19 1.13912 $w=6.28e-07 $l=6e-08 $layer=LI1_cond $X=0.415 $Y=1.295
+ $X2=0.415 $Y2=1.355
r40 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.565 $Y=1.695
+ $X2=0.565 $Y2=1.355
r41 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.695
+ $X2=0.565 $Y2=1.86
r42 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.19
+ $X2=0.565 $Y2=1.355
r43 7 12 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.475 $Y=2.545
+ $X2=0.475 $Y2=1.86
r44 3 10 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.475 $Y=0.47
+ $X2=0.475 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_LP__DLYGATE4S18_1%A_27_52# 1 2 8 11 15 19 23 25 26 27 28
+ 32 33 36
r60 36 40 40.7881 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.765
+ $X2=1.19 $Y2=1.93
r61 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.765 $X2=1.14 $Y2=1.765
r62 33 38 40.7881 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.19 $Y=1.085
+ $X2=1.19 $Y2=0.92
r63 32 35 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.14 $Y=1.085
+ $X2=1.14 $Y2=1.765
r64 32 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.085 $X2=1.14 $Y2=1.085
r65 30 35 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.14 $Y=2.03
+ $X2=1.14 $Y2=1.765
r66 29 32 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.14 $Y=1.02
+ $X2=1.14 $Y2=1.085
r67 27 29 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=0.975 $Y=0.92
+ $X2=1.14 $Y2=1.02
r68 27 28 31.3318 $w=1.98e-07 $l=5.65e-07 $layer=LI1_cond $X=0.975 $Y=0.92
+ $X2=0.41 $Y2=0.92
r69 25 30 7.68689 $w=1.75e-07 $l=2.03912e-07 $layer=LI1_cond $X=0.975 $Y=2.117
+ $X2=1.14 $Y2=2.03
r70 25 26 36.4416 $w=1.73e-07 $l=5.75e-07 $layer=LI1_cond $X=0.975 $Y=2.117
+ $X2=0.4 $Y2=2.117
r71 21 26 7.48781 $w=1.75e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.247 $Y=2.205
+ $X2=0.4 $Y2=2.117
r72 21 23 13.4137 $w=3.03e-07 $l=3.55e-07 $layer=LI1_cond $X=0.247 $Y=2.205
+ $X2=0.247 $Y2=2.56
r73 17 28 7.26812 $w=2e-07 $l=2.01901e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.41 $Y2=0.92
r74 17 19 12.8049 $w=3.13e-07 $l=3.5e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.252 $Y2=0.47
r75 15 40 239.056 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=1.35 $Y=2.545
+ $X2=1.35 $Y2=1.93
r76 11 38 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=1.35 $Y=0.47
+ $X2=1.35 $Y2=0.92
r77 8 36 9.0955 $w=5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.19 $Y=1.68 $X2=1.19
+ $Y2=1.765
r78 7 33 9.0955 $w=5e-07 $l=8.5e-08 $layer=POLY_cond $X=1.19 $Y=1.17 $X2=1.19
+ $Y2=1.085
r79 7 8 54.573 $w=5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.19 $Y=1.17 $X2=1.19
+ $Y2=1.68
r80 2 23 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.335 $X2=0.26 $Y2=2.56
r81 1 19 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.26 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLYGATE4S18_1%A_288_52# 1 2 9 13 16 21 22 25 29 30
+ 32
c57 21 0 2.41794e-20 $X=2.575 $Y=1.51
r58 29 30 6.71392 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.567 $Y=2.56
+ $X2=1.567 $Y2=2.395
r59 25 27 6.71392 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.567 $Y=0.47
+ $X2=1.567 $Y2=0.635
r60 22 33 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.575 $Y=1.51
+ $X2=2.38 $Y2=1.51
r61 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.575
+ $Y=1.51 $X2=2.575 $Y2=1.51
r62 19 32 0.995122 $w=2.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.72 $Y=1.52
+ $X2=1.597 $Y2=1.52
r63 19 21 36.494 $w=2.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.72 $Y=1.52
+ $X2=2.575 $Y2=1.52
r64 17 32 5.59678 $w=2.45e-07 $l=1.35e-07 $layer=LI1_cond $X=1.597 $Y=1.655
+ $X2=1.597 $Y2=1.52
r65 17 30 34.8085 $w=2.43e-07 $l=7.4e-07 $layer=LI1_cond $X=1.597 $Y=1.655
+ $X2=1.597 $Y2=2.395
r66 16 32 5.59678 $w=2.45e-07 $l=1.35e-07 $layer=LI1_cond $X=1.597 $Y=1.385
+ $X2=1.597 $Y2=1.52
r67 16 27 35.2789 $w=2.43e-07 $l=7.5e-07 $layer=LI1_cond $X=1.597 $Y=1.385
+ $X2=1.597 $Y2=0.635
r68 11 33 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.675
+ $X2=2.38 $Y2=1.51
r69 11 13 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.38 $Y=1.675
+ $X2=2.38 $Y2=2.045
r70 7 33 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.345
+ $X2=2.38 $Y2=1.51
r71 7 9 176.863 $w=1.8e-07 $l=4.55e-07 $layer=POLY_cond $X=2.38 $Y=1.345
+ $X2=2.38 $Y2=0.89
r72 2 29 600 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=1 $X=1.44
+ $Y=2.335 $X2=1.58 $Y2=2.56
r73 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.26 $X2=1.58 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLYGATE4S18_1%A_405_136# 1 2 9 13 15 17 19 20 22 26
+ 34
c64 20 0 1.65637e-19 $X=3.032 $Y=1.825
c65 13 0 2.41794e-20 $X=3.205 $Y=2.465
r66 34 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.46
+ $X2=3.165 $Y2=1.625
r67 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.46
+ $X2=3.165 $Y2=1.295
r68 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.165
+ $Y=1.46 $X2=3.165 $Y2=1.46
r69 31 33 12.7405 $w=3.16e-07 $l=3.3e-07 $layer=LI1_cond $X=3.095 $Y=1.13
+ $X2=3.095 $Y2=1.46
r70 26 29 3.68142 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=2.165 $Y=1.91
+ $X2=2.165 $Y2=2.025
r71 22 24 8.16314 $w=3.58e-07 $l=2.55e-07 $layer=LI1_cond $X=2.165 $Y=0.875
+ $X2=2.165 $Y2=1.13
r72 19 33 7.01833 $w=3.16e-07 $l=1.93959e-07 $layer=LI1_cond $X=3.032 $Y=1.625
+ $X2=3.095 $Y2=1.46
r73 19 20 9.4077 $w=2.43e-07 $l=2e-07 $layer=LI1_cond $X=3.032 $Y=1.625
+ $X2=3.032 $Y2=1.825
r74 18 26 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.345 $Y=1.91
+ $X2=2.165 $Y2=1.91
r75 17 20 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.91 $Y=1.91
+ $X2=3.032 $Y2=1.825
r76 17 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.91 $Y=1.91
+ $X2=2.345 $Y2=1.91
r77 16 24 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.345 $Y=1.13
+ $X2=2.165 $Y2=1.13
r78 15 31 4.36715 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.91 $Y=1.13
+ $X2=3.095 $Y2=1.13
r79 15 16 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.91 $Y=1.13
+ $X2=2.345 $Y2=1.13
r80 13 37 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.205 $Y=2.465
+ $X2=3.205 $Y2=1.625
r81 9 36 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.205 $Y=0.68
+ $X2=3.205 $Y2=1.295
r82 2 29 600 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_PDIFF $count=1 $X=2.025
+ $Y=1.835 $X2=2.15 $Y2=2.025
r83 1 22 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.68 $X2=2.15 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__DLYGATE4S18_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
r32 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r34 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r35 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 29 32 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r39 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=0.735 $Y2=3.33
r40 27 29 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=1.2
+ $Y2=3.33
r41 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.735 $Y2=3.33
r44 22 24 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 20 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 20 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 18 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.99 $Y2=3.33
r49 17 35 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.6 $Y2=3.33
r50 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=2.99 $Y2=3.33
r51 13 16 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.99 $Y=2.27
+ $X2=2.99 $Y2=2.95
r52 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=3.245
+ $X2=2.99 $Y2=3.33
r53 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.99 $Y=3.245
+ $X2=2.99 $Y2=2.95
r54 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r55 7 9 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.735 $Y=3.245 $X2=0.735
+ $Y2=2.545
r56 2 16 400 $w=1.7e-07 $l=1.35019e-06 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.835 $X2=2.99 $Y2=2.95
r57 2 13 400 $w=1.7e-07 $l=7.04699e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=1.835 $X2=2.99 $Y2=2.27
r58 1 9 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.335 $X2=0.735 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__DLYGATE4S18_1%X 1 2 7 8 9 10 11 12 13 25 38 48 52
r22 52 53 5.64022 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.532 $Y=1.98
+ $X2=3.532 $Y2=1.815
r23 36 38 0.361006 $w=4.13e-07 $l=1.3e-08 $layer=LI1_cond $X=3.532 $Y=2.022
+ $X2=3.532 $Y2=2.035
r24 23 48 0.333237 $w=4.13e-07 $l=1.2e-08 $layer=LI1_cond $X=3.532 $Y=0.913
+ $X2=3.532 $Y2=0.925
r25 13 45 3.74891 $w=4.13e-07 $l=1.35e-07 $layer=LI1_cond $X=3.532 $Y=2.775
+ $X2=3.532 $Y2=2.91
r26 12 13 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.532 $Y=2.405
+ $X2=3.532 $Y2=2.775
r27 11 36 0.99971 $w=4.13e-07 $l=3.6e-08 $layer=LI1_cond $X=3.532 $Y=1.986
+ $X2=3.532 $Y2=2.022
r28 11 52 0.166618 $w=4.13e-07 $l=6e-09 $layer=LI1_cond $X=3.532 $Y=1.986
+ $X2=3.532 $Y2=1.98
r29 11 12 9.27508 $w=4.13e-07 $l=3.34e-07 $layer=LI1_cond $X=3.532 $Y=2.071
+ $X2=3.532 $Y2=2.405
r30 11 38 0.99971 $w=4.13e-07 $l=3.6e-08 $layer=LI1_cond $X=3.532 $Y=2.071
+ $X2=3.532 $Y2=2.035
r31 10 53 5.96091 $w=2.88e-07 $l=1.5e-07 $layer=LI1_cond $X=3.595 $Y=1.665
+ $X2=3.595 $Y2=1.815
r32 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.595 $Y=1.295
+ $X2=3.595 $Y2=1.665
r33 9 50 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=3.595 $Y=1.295
+ $X2=3.595 $Y2=1.12
r34 8 50 5.4736 $w=4.13e-07 $l=1.59e-07 $layer=LI1_cond $X=3.532 $Y=0.961
+ $X2=3.532 $Y2=1.12
r35 8 48 0.99971 $w=4.13e-07 $l=3.6e-08 $layer=LI1_cond $X=3.532 $Y=0.961
+ $X2=3.532 $Y2=0.925
r36 8 23 1.02748 $w=4.13e-07 $l=3.7e-08 $layer=LI1_cond $X=3.532 $Y=0.876
+ $X2=3.532 $Y2=0.913
r37 7 8 8.91408 $w=4.13e-07 $l=3.21e-07 $layer=LI1_cond $X=3.532 $Y=0.555
+ $X2=3.532 $Y2=0.876
r38 7 25 3.74891 $w=4.13e-07 $l=1.35e-07 $layer=LI1_cond $X=3.532 $Y=0.555
+ $X2=3.532 $Y2=0.42
r39 2 52 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.835 $X2=3.42 $Y2=1.98
r40 2 45 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.835 $X2=3.42 $Y2=2.91
r41 1 25 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=3.28
+ $Y=0.26 $X2=3.42 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLYGATE4S18_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r38 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r40 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r41 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r44 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.745
+ $Y2=0
r46 25 27 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.2
+ $Y2=0
r47 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r48 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r49 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.745
+ $Y2=0
r50 20 22 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.24
+ $Y2=0
r51 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r52 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r53 16 30 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.64
+ $Y2=0
r54 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.99
+ $Y2=0
r55 15 33 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=3.6
+ $Y2=0
r56 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=2.99
+ $Y2=0
r57 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=2.99 $Y2=0
r58 11 13 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=2.99 $Y2=0.415
r59 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r60 7 9 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.47
r61 2 13 91 $w=1.7e-07 $l=6.38905e-07 $layer=licon1_NDIFF $count=2 $X=2.47
+ $Y=0.68 $X2=2.99 $Y2=0.415
r62 1 9 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.26 $X2=0.745 $Y2=0.47
.ends

