* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_2 A0 A1 S VGND VNB VPB VPWR X
M1000 a_350_449# a_284_279# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.05375e+12p ps=8.59e+06u
M1001 a_319_48# a_284_279# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=7.269e+11p ps=6.53e+06u
M1002 VPWR S a_508_449# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.048e+11p ps=1.92e+06u
M1003 VGND S a_499_48# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 a_508_449# A0 a_86_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1005 a_499_48# A1 a_86_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.638e+11p ps=1.62e+06u
M1006 X a_86_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1007 X a_86_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1008 VGND a_86_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_284_279# S VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1010 a_86_21# A1 a_350_449# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_86_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_284_279# S VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1013 a_86_21# A0 a_319_48# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
