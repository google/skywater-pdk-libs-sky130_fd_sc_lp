* File: sky130_fd_sc_lp__sdfxtp_2.spice
* Created: Wed Sep  2 10:36:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfxtp_2.pex.spice"
.subckt sky130_fd_sc_lp__sdfxtp_2  VNB VPB D SCE SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* SCE	SCE
* D	D
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_SCE_M1008_g N_A_55_119#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.1197 PD=0.84 PS=1.41 NRD=2.856 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1007 A_256_119# N_A_55_119#_M1007_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0882 PD=0.63 PS=0.84 NRD=14.28 NRS=37.14 M=1 R=2.8 SA=75000.8
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1004 N_A_328_119#_M1004_d N_D_M1004_g A_256_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=0.95 PS=0.63 NRD=68.568 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1017 A_464_119# N_SCE_M1017_g N_A_328_119#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=0.95 NRD=14.28 NRS=2.856 M=1 R=2.8 SA=75001.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_SCD_M1009_g A_464_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.0441 PD=0.79 PS=0.63 NRD=11.424 NRS=14.28 M=1 R=2.8 SA=75002.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1023 N_A_610_487#_M1023_d N_CLK_M1023_g N_VGND_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0777 PD=1.37 PS=0.79 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75002.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 N_A_831_47#_M1032_d N_A_610_487#_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1428 AS=0.1134 PD=1.52 PS=1.38 NRD=0 NRS=1.428 M=1 R=2.8
+ SA=75000.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1012 N_A_1047_125#_M1012_d N_A_610_487#_M1012_g N_A_328_119#_M1012_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0756 AS=0.1197 PD=0.78 PS=1.41 NRD=0 NRS=5.712 M=1
+ R=2.8 SA=75000.2 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1027 A_1149_125# N_A_831_47#_M1027_g N_A_1047_125#_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=22.848 M=1 R=2.8
+ SA=75000.7 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1178_399#_M1020_g A_1149_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.195855 AS=0.0504 PD=1.19264 PS=0.66 NRD=117.516 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1015 N_A_1178_399#_M1015_d N_A_1047_125#_M1015_g N_VGND_M1020_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.130294 AS=0.298445 PD=1.22566 PS=1.81736 NRD=0 NRS=73.116
+ M=1 R=4.26667 SA=75001.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1033 N_A_1517_63#_M1033_d N_A_831_47#_M1033_g N_A_1178_399#_M1015_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.12915 AS=0.0855057 PD=1.035 PS=0.80434 NRD=39.996
+ NRS=42.444 M=1 R=2.8 SA=75001.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1026 A_1670_63# N_A_610_487#_M1026_g N_A_1517_63#_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.12915 PD=0.63 PS=1.035 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_A_1665_381#_M1028_g A_1670_63# VNB NSHORT L=0.15 W=0.42
+ AD=0.0855057 AS=0.0441 PD=0.80434 PS=0.63 NRD=28.56 NRS=14.28 M=1 R=2.8
+ SA=75002.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1025 N_A_1665_381#_M1025_d N_A_1517_63#_M1025_g N_VGND_M1028_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.130294 PD=1.81 PS=1.22566 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_Q_M1003_d N_A_1665_381#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_Q_M1003_d N_A_1665_381#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1029 N_VPWR_M1029_d N_SCE_M1029_g N_A_55_119#_M1029_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1152 AS=0.1824 PD=1 PS=1.85 NRD=10.7562 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1030 A_256_487# N_SCE_M1030_g N_VPWR_M1029_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1152 PD=0.85 PS=1 NRD=15.3857 NRS=13.8491 M=1 R=4.26667
+ SA=75000.7 SB=75002 A=0.096 P=1.58 MULT=1
MM1018 N_A_328_119#_M1018_d N_D_M1018_g A_256_487# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.1
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1005 A_414_487# N_A_55_119#_M1005_g N_A_328_119#_M1018_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=32.308 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_SCD_M1001_g A_414_487# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1152 AS=0.1024 PD=1 PS=0.96 NRD=18.4589 NRS=32.308 M=1 R=4.26667 SA=75002
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1031 N_A_610_487#_M1031_d N_CLK_M1031_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1152 PD=1.81 PS=1 NRD=0 NRS=6.1464 M=1 R=4.26667
+ SA=75002.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_831_47#_M1006_d N_A_610_487#_M1006_g N_VPWR_M1006_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.3424 PD=1.81 PS=2.35 NRD=0 NRS=80.0214 M=1
+ R=4.26667 SA=75000.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1021 N_A_1047_125#_M1021_d N_A_831_47#_M1021_g N_A_328_119#_M1021_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1011 A_1136_451# N_A_610_487#_M1011_g N_A_1047_125#_M1021_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_1178_399#_M1002_g A_1136_451# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1855 AS=0.0441 PD=1.02667 PS=0.63 NRD=39.8531 NRS=23.443 M=1 R=2.8
+ SA=75001 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_1178_399#_M1014_d N_A_1047_125#_M1014_g N_VPWR_M1002_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.231 AS=0.371 PD=1.39 PS=2.05333 NRD=0 NRS=79.7259 M=1 R=5.6
+ SA=75001.2 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1019 N_A_1517_63#_M1019_d N_A_610_487#_M1019_g N_A_1178_399#_M1014_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1792 AS=0.231 PD=1.62 PS=1.39 NRD=0 NRS=63.3158 M=1
+ R=5.6 SA=75001.9 SB=75001 A=0.126 P=1.98 MULT=1
MM1016 A_1623_493# N_A_831_47#_M1016_g N_A_1517_63#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0896 PD=0.63 PS=0.81 NRD=23.443 NRS=46.886 M=1 R=2.8
+ SA=75002.4 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1022_d N_A_1665_381#_M1022_g A_1623_493# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1274 AS=0.0441 PD=0.976667 PS=0.63 NRD=164.16 NRS=23.443 M=1 R=2.8
+ SA=75002.8 SB=75001 A=0.063 P=1.14 MULT=1
MM1000 N_A_1665_381#_M1000_d N_A_1517_63#_M1000_g N_VPWR_M1022_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.2548 PD=2.21 PS=1.95333 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_Q_M1013_d N_A_1665_381#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1024 N_Q_M1013_d N_A_1665_381#_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=21.2983 P=26.57
c_116 VNB 0 9.65774e-20 $X=0 $Y=0
c_1577 A_414_487# 0 1.20926e-19 $X=2.07 $Y=2.435
*
.include "sky130_fd_sc_lp__sdfxtp_2.pxi.spice"
*
.ends
*
*
