* File: sky130_fd_sc_lp__invkapwr_8.pex.spice
* Created: Fri Aug 28 10:39:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INVKAPWR_8%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55
+ 59 63 67 71 75 79 81 82 83 84 85 86 87 88 89 90 119
r179 117 119 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.1 $Y=1.375
+ $X2=5.275 $Y2=1.375
r180 115 117 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=4.845 $Y=1.375
+ $X2=5.1 $Y2=1.375
r181 114 115 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.415 $Y=1.375
+ $X2=4.845 $Y2=1.375
r182 113 114 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.985 $Y=1.375
+ $X2=4.415 $Y2=1.375
r183 112 113 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.555 $Y=1.375
+ $X2=3.985 $Y2=1.375
r184 111 112 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.125 $Y=1.375
+ $X2=3.555 $Y2=1.375
r185 110 111 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.695 $Y=1.375
+ $X2=3.125 $Y2=1.375
r186 109 110 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.265 $Y=1.375
+ $X2=2.695 $Y2=1.375
r187 108 109 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.835 $Y=1.375
+ $X2=2.265 $Y2=1.375
r188 107 108 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.405 $Y=1.375
+ $X2=1.835 $Y2=1.375
r189 106 107 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.975 $Y=1.375
+ $X2=1.405 $Y2=1.375
r190 104 106 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=0.68 $Y=1.375
+ $X2=0.975 $Y2=1.375
r191 101 104 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=0.545 $Y=1.375
+ $X2=0.68 $Y2=1.375
r192 90 117 20.7543 $w=1.7e-07 $l=1.19e-06 $layer=licon1_POLY $count=7 $X=5.1
+ $Y=1.375 $X2=5.1 $Y2=1.375
r193 89 90 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.375
+ $X2=5.04 $Y2=1.375
r194 88 89 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.375
+ $X2=4.56 $Y2=1.375
r195 87 88 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.375
+ $X2=4.08 $Y2=1.375
r196 86 87 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.375
+ $X2=3.6 $Y2=1.375
r197 85 86 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.375
+ $X2=3.12 $Y2=1.375
r198 84 85 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.375
+ $X2=2.64 $Y2=1.375
r199 83 84 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.375
+ $X2=2.16 $Y2=1.375
r200 82 83 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.375
+ $X2=1.68 $Y2=1.375
r201 81 82 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=0.68 $Y=1.375
+ $X2=1.2 $Y2=1.375
r202 81 104 20.7543 $w=1.7e-07 $l=1.19e-06 $layer=licon1_POLY $count=7 $X=0.68
+ $Y=1.375 $X2=0.68 $Y2=1.375
r203 77 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.275 $Y=1.54
+ $X2=5.275 $Y2=1.375
r204 77 79 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=5.275 $Y=1.54
+ $X2=5.275 $Y2=2.465
r205 73 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.845 $Y=1.54
+ $X2=4.845 $Y2=1.375
r206 73 75 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=4.845 $Y=1.54
+ $X2=4.845 $Y2=2.465
r207 69 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.54
+ $X2=4.415 $Y2=1.375
r208 69 71 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=4.415 $Y=1.54
+ $X2=4.415 $Y2=2.465
r209 65 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.21
+ $X2=4.415 $Y2=1.375
r210 65 67 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=4.415 $Y=1.21
+ $X2=4.415 $Y2=0.56
r211 61 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.54
+ $X2=3.985 $Y2=1.375
r212 61 63 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.985 $Y=1.54
+ $X2=3.985 $Y2=2.465
r213 57 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.21
+ $X2=3.985 $Y2=1.375
r214 57 59 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.985 $Y=1.21
+ $X2=3.985 $Y2=0.56
r215 53 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.555 $Y=1.54
+ $X2=3.555 $Y2=1.375
r216 53 55 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.555 $Y=1.54
+ $X2=3.555 $Y2=2.465
r217 49 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.555 $Y=1.21
+ $X2=3.555 $Y2=1.375
r218 49 51 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.555 $Y=1.21
+ $X2=3.555 $Y2=0.56
r219 45 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.54
+ $X2=3.125 $Y2=1.375
r220 45 47 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.125 $Y=1.54
+ $X2=3.125 $Y2=2.465
r221 41 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.21
+ $X2=3.125 $Y2=1.375
r222 41 43 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.125 $Y=1.21
+ $X2=3.125 $Y2=0.56
r223 37 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.54
+ $X2=2.695 $Y2=1.375
r224 37 39 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.695 $Y=1.54
+ $X2=2.695 $Y2=2.465
r225 33 110 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.21
+ $X2=2.695 $Y2=1.375
r226 33 35 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.695 $Y=1.21
+ $X2=2.695 $Y2=0.56
r227 29 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.54
+ $X2=2.265 $Y2=1.375
r228 29 31 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.265 $Y=1.54
+ $X2=2.265 $Y2=2.465
r229 25 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.21
+ $X2=2.265 $Y2=1.375
r230 25 27 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.265 $Y=1.21
+ $X2=2.265 $Y2=0.56
r231 21 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.54
+ $X2=1.835 $Y2=1.375
r232 21 23 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.835 $Y=1.54
+ $X2=1.835 $Y2=2.465
r233 17 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.21
+ $X2=1.835 $Y2=1.375
r234 17 19 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.835 $Y=1.21
+ $X2=1.835 $Y2=0.56
r235 13 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.54
+ $X2=1.405 $Y2=1.375
r236 13 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.405 $Y=1.54
+ $X2=1.405 $Y2=2.465
r237 9 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.21
+ $X2=1.405 $Y2=1.375
r238 9 11 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.405 $Y=1.21
+ $X2=1.405 $Y2=0.56
r239 5 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.54
+ $X2=0.975 $Y2=1.375
r240 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.975 $Y=1.54
+ $X2=0.975 $Y2=2.465
r241 1 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.54
+ $X2=0.545 $Y2=1.375
r242 1 3 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.545 $Y=1.54
+ $X2=0.545 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_8%KAPWR 1 2 3 4 5 6 7 22 25 33 41 49 57 65
+ 73 77
r77 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.495 $Y=2.81
+ $X2=5.495 $Y2=2.81
r78 73 76 26.6644 $w=2.53e-07 $l=5.9e-07 $layer=LI1_cond $X=5.487 $Y=2.22
+ $X2=5.487 $Y2=2.81
r79 69 77 0.497684 $w=2.55e-07 $l=8.6e-07 $layer=MET1_cond $X=4.635 $Y=2.817
+ $X2=5.495 $Y2=2.817
r80 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.635 $Y=2.81
+ $X2=4.635 $Y2=2.81
r81 65 68 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=4.63 $Y=2.22
+ $X2=4.63 $Y2=2.81
r82 61 69 0.497684 $w=2.55e-07 $l=8.6e-07 $layer=MET1_cond $X=3.775 $Y=2.817
+ $X2=4.635 $Y2=2.817
r83 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.775 $Y=2.81
+ $X2=3.775 $Y2=2.81
r84 57 60 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=3.77 $Y=2.22
+ $X2=3.77 $Y2=2.81
r85 49 52 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=2.91 $Y=2.22
+ $X2=2.91 $Y2=2.81
r86 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.055 $Y=2.81
+ $X2=2.055 $Y2=2.81
r87 41 44 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=2.05 $Y=2.22
+ $X2=2.05 $Y2=2.81
r88 37 45 0.503471 $w=2.55e-07 $l=8.7e-07 $layer=MET1_cond $X=1.185 $Y=2.817
+ $X2=2.055 $Y2=2.817
r89 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.185 $Y=2.81
+ $X2=1.185 $Y2=2.81
r90 33 36 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=1.19 $Y=2.22
+ $X2=1.19 $Y2=2.81
r91 29 37 0.49479 $w=2.55e-07 $l=8.55e-07 $layer=MET1_cond $X=0.33 $Y=2.817
+ $X2=1.185 $Y2=2.817
r92 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.33 $Y=2.81
+ $X2=0.33 $Y2=2.81
r93 25 28 26.1516 $w=2.58e-07 $l=5.9e-07 $layer=LI1_cond $X=0.33 $Y=2.22
+ $X2=0.33 $Y2=2.81
r94 22 61 0.517938 $w=2.55e-07 $l=8.95e-07 $layer=MET1_cond $X=2.88 $Y=2.817
+ $X2=3.775 $Y2=2.817
r95 22 45 0.477429 $w=2.55e-07 $l=8.25e-07 $layer=MET1_cond $X=2.88 $Y=2.817
+ $X2=2.055 $Y2=2.817
r96 22 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.91 $Y=2.81
+ $X2=2.91 $Y2=2.81
r97 7 76 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.835 $X2=5.49 $Y2=2.91
r98 7 73 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.835 $X2=5.49 $Y2=2.22
r99 6 68 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.49
+ $Y=1.835 $X2=4.63 $Y2=2.91
r100 6 65 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=4.49
+ $Y=1.835 $X2=4.63 $Y2=2.22
r101 5 60 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.63
+ $Y=1.835 $X2=3.77 $Y2=2.91
r102 5 57 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=3.63
+ $Y=1.835 $X2=3.77 $Y2=2.22
r103 4 52 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.835 $X2=2.91 $Y2=2.91
r104 4 49 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.835 $X2=2.91 $Y2=2.22
r105 3 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=2.91
r106 3 41 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=2.22
r107 2 36 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.91
r108 2 33 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.22
r109 1 28 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.91
r110 1 25 400 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_8%Y 1 2 3 4 5 6 7 8 9 10 32 33 34 35 36 39
+ 43 47 51 55 57 61 65 69 71 75 79 83 85 89 93 97 101 105 107 108 109 110 111
+ 112 113 115 116 117 119 120 124
r197 120 124 15.2875 $w=1.83e-07 $l=2.55e-07 $layer=LI1_cond $X=5.527 $Y=1.295
+ $X2=5.527 $Y2=1.04
r198 119 124 3.55727 $w=1.85e-07 $l=1e-07 $layer=LI1_cond $X=5.527 $Y=0.94
+ $X2=5.527 $Y2=1.04
r199 118 120 24.8796 $w=1.83e-07 $l=4.15e-07 $layer=LI1_cond $X=5.527 $Y=1.71
+ $X2=5.527 $Y2=1.295
r200 114 119 35.7429 $w=3.68e-07 $l=1.105e-06 $layer=LI1_cond $X=4.33 $Y=0.94
+ $X2=5.435 $Y2=0.94
r201 114 115 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=4.33 $Y=0.94 $X2=4.2
+ $Y2=0.94
r202 106 117 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=5.19 $Y=1.797
+ $X2=5.06 $Y2=1.797
r203 105 118 6.82334 $w=1.75e-07 $l=1.28328e-07 $layer=LI1_cond $X=5.435
+ $Y=1.797 $X2=5.527 $Y2=1.71
r204 105 106 15.5273 $w=1.73e-07 $l=2.45e-07 $layer=LI1_cond $X=5.435 $Y=1.797
+ $X2=5.19 $Y2=1.797
r205 101 103 39.0058 $w=2.58e-07 $l=8.8e-07 $layer=LI1_cond $X=5.06 $Y=2
+ $X2=5.06 $Y2=2.88
r206 99 117 0.0359085 $w=2.6e-07 $l=8.8e-08 $layer=LI1_cond $X=5.06 $Y=1.885
+ $X2=5.06 $Y2=1.797
r207 99 101 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=5.06 $Y=1.885
+ $X2=5.06 $Y2=2
r208 98 116 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=4.33 $Y=1.797
+ $X2=4.202 $Y2=1.797
r209 97 117 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=4.93 $Y=1.797
+ $X2=5.06 $Y2=1.797
r210 97 98 38.026 $w=1.73e-07 $l=6e-07 $layer=LI1_cond $X=4.93 $Y=1.797 $X2=4.33
+ $Y2=1.797
r211 93 95 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=4.202 $Y=2
+ $X2=4.202 $Y2=2.88
r212 91 116 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=4.202 $Y=1.885
+ $X2=4.202 $Y2=1.797
r213 91 93 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=4.202 $Y=1.885
+ $X2=4.202 $Y2=2
r214 87 115 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=4.2 $Y=0.84 $X2=4.2
+ $Y2=0.94
r215 87 89 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=4.2 $Y=0.84 $X2=4.2
+ $Y2=0.56
r216 86 113 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=3.47 $Y=1.797
+ $X2=3.342 $Y2=1.797
r217 85 116 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=4.075 $Y=1.797
+ $X2=4.202 $Y2=1.797
r218 85 86 38.3429 $w=1.73e-07 $l=6.05e-07 $layer=LI1_cond $X=4.075 $Y=1.797
+ $X2=3.47 $Y2=1.797
r219 84 112 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=3.47 $Y=0.94 $X2=3.34
+ $Y2=0.94
r220 83 115 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=4.07 $Y=0.94 $X2=4.2
+ $Y2=0.94
r221 83 84 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=4.07 $Y=0.94 $X2=3.47
+ $Y2=0.94
r222 79 81 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=3.342 $Y=2
+ $X2=3.342 $Y2=2.88
r223 77 113 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=3.342 $Y=1.885
+ $X2=3.342 $Y2=1.797
r224 77 79 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=3.342 $Y=1.885
+ $X2=3.342 $Y2=2
r225 73 112 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=3.34 $Y=0.84
+ $X2=3.34 $Y2=0.94
r226 73 75 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=3.34 $Y=0.84
+ $X2=3.34 $Y2=0.56
r227 72 111 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=2.61 $Y=1.797
+ $X2=2.482 $Y2=1.797
r228 71 113 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=3.215 $Y=1.797
+ $X2=3.342 $Y2=1.797
r229 71 72 38.3429 $w=1.73e-07 $l=6.05e-07 $layer=LI1_cond $X=3.215 $Y=1.797
+ $X2=2.61 $Y2=1.797
r230 70 110 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=2.61 $Y=0.94 $X2=2.48
+ $Y2=0.94
r231 69 112 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=3.21 $Y=0.94 $X2=3.34
+ $Y2=0.94
r232 69 70 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=3.21 $Y=0.94 $X2=2.61
+ $Y2=0.94
r233 65 67 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=2.482 $Y=2
+ $X2=2.482 $Y2=2.88
r234 63 111 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=2.482 $Y=1.885
+ $X2=2.482 $Y2=1.797
r235 63 65 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=2.482 $Y=1.885
+ $X2=2.482 $Y2=2
r236 59 110 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=2.48 $Y=0.84
+ $X2=2.48 $Y2=0.94
r237 59 61 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=2.48 $Y=0.84
+ $X2=2.48 $Y2=0.56
r238 58 109 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=1.75 $Y=1.797
+ $X2=1.622 $Y2=1.797
r239 57 111 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=2.355 $Y=1.797
+ $X2=2.482 $Y2=1.797
r240 57 58 38.3429 $w=1.73e-07 $l=6.05e-07 $layer=LI1_cond $X=2.355 $Y=1.797
+ $X2=1.75 $Y2=1.797
r241 56 108 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.75 $Y=0.94 $X2=1.62
+ $Y2=0.94
r242 55 110 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=2.35 $Y=0.94 $X2=2.48
+ $Y2=0.94
r243 55 56 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=2.35 $Y=0.94 $X2=1.75
+ $Y2=0.94
r244 51 53 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=1.622 $Y=2
+ $X2=1.622 $Y2=2.88
r245 49 109 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=1.622 $Y=1.885
+ $X2=1.622 $Y2=1.797
r246 49 51 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=1.622 $Y=1.885
+ $X2=1.622 $Y2=2
r247 45 108 0.417182 $w=2.6e-07 $l=1e-07 $layer=LI1_cond $X=1.62 $Y=0.84
+ $X2=1.62 $Y2=0.94
r248 45 47 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=1.62 $Y=0.84
+ $X2=1.62 $Y2=0.56
r249 44 107 6.97918 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=0.89 $Y=1.797
+ $X2=0.762 $Y2=1.797
r250 43 109 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=1.495 $Y=1.797
+ $X2=1.622 $Y2=1.797
r251 43 44 38.3429 $w=1.73e-07 $l=6.05e-07 $layer=LI1_cond $X=1.495 $Y=1.797
+ $X2=0.89 $Y2=1.797
r252 39 41 39.7706 $w=2.53e-07 $l=8.8e-07 $layer=LI1_cond $X=0.762 $Y=2
+ $X2=0.762 $Y2=2.88
r253 37 107 0.0291048 $w=2.55e-07 $l=8.8e-08 $layer=LI1_cond $X=0.762 $Y=1.885
+ $X2=0.762 $Y2=1.797
r254 37 39 5.19729 $w=2.53e-07 $l=1.15e-07 $layer=LI1_cond $X=0.762 $Y=1.885
+ $X2=0.762 $Y2=2
r255 35 107 6.97918 $w=1.75e-07 $l=1.27e-07 $layer=LI1_cond $X=0.635 $Y=1.797
+ $X2=0.762 $Y2=1.797
r256 35 36 18.3792 $w=1.73e-07 $l=2.9e-07 $layer=LI1_cond $X=0.635 $Y=1.797
+ $X2=0.345 $Y2=1.797
r257 33 108 6.3888 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=1.49 $Y=0.94 $X2=1.62
+ $Y2=0.94
r258 33 34 63.4955 $w=1.98e-07 $l=1.145e-06 $layer=LI1_cond $X=1.49 $Y=0.94
+ $X2=0.345 $Y2=0.94
r259 32 36 6.81835 $w=1.75e-07 $l=1.22327e-07 $layer=LI1_cond $X=0.26 $Y=1.71
+ $X2=0.345 $Y2=1.797
r260 31 34 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.26 $Y=1.04
+ $X2=0.345 $Y2=0.94
r261 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.26 $Y=1.04
+ $X2=0.26 $Y2=1.71
r262 10 103 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.835 $X2=5.06 $Y2=2.88
r263 10 101 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.835 $X2=5.06 $Y2=2
r264 9 95 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=4.06
+ $Y=1.835 $X2=4.2 $Y2=2.88
r265 9 93 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=4.06
+ $Y=1.835 $X2=4.2 $Y2=2
r266 8 81 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.835 $X2=3.34 $Y2=2.88
r267 8 79 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.835 $X2=3.34 $Y2=2
r268 7 67 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=1.835 $X2=2.48 $Y2=2.88
r269 7 65 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=1.835 $X2=2.48 $Y2=2
r270 6 53 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=2.88
r271 6 51 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=2
r272 5 41 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2.88
r273 5 39 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2
r274 4 89 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.35 $X2=4.2 $Y2=0.56
r275 3 75 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.35 $X2=3.34 $Y2=0.56
r276 2 61 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.34
+ $Y=0.35 $X2=2.48 $Y2=0.56
r277 1 47 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.35 $X2=1.62 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_8%VGND 1 2 3 4 5 18 22 26 30 32 36 39 40 42
+ 43 44 45 46 48 65 66 69 72
r61 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r62 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r63 66 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r64 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r65 63 72 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.647
+ $Y2=0
r66 63 65 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=5.52
+ $Y2=0
r67 62 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r68 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r69 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r70 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r71 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r72 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r73 53 69 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.172
+ $Y2=0
r74 53 55 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.32 $Y=0 $X2=1.68
+ $Y2=0
r75 51 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r76 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r77 48 69 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.172
+ $Y2=0
r78 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=0.72
+ $Y2=0
r79 46 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r80 46 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r81 44 61 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.6
+ $Y2=0
r82 44 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.77
+ $Y2=0
r83 42 58 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.64
+ $Y2=0
r84 42 43 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.91
+ $Y2=0
r85 41 61 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.6
+ $Y2=0
r86 41 43 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.91
+ $Y2=0
r87 39 55 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r88 39 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.92 $Y=0 $X2=2.05
+ $Y2=0
r89 38 58 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.64
+ $Y2=0
r90 38 40 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.05
+ $Y2=0
r91 34 72 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.647 $Y=0.085
+ $X2=4.647 $Y2=0
r92 34 36 16.4077 $w=2.93e-07 $l=4.2e-07 $layer=LI1_cond $X=4.647 $Y=0.085
+ $X2=4.647 $Y2=0.505
r93 33 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.9 $Y=0 $X2=3.77
+ $Y2=0
r94 32 72 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=4.647
+ $Y2=0
r95 32 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.5 $Y=0 $X2=3.9 $Y2=0
r96 28 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=0.085
+ $X2=3.77 $Y2=0
r97 28 30 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=3.77 $Y=0.085
+ $X2=3.77 $Y2=0.505
r98 24 43 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.91 $Y2=0
r99 24 26 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=2.91 $Y=0.085
+ $X2=2.91 $Y2=0.505
r100 20 40 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=0.085
+ $X2=2.05 $Y2=0
r101 20 22 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=2.05 $Y=0.085
+ $X2=2.05 $Y2=0.505
r102 16 69 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.172 $Y=0.085
+ $X2=1.172 $Y2=0
r103 16 18 16.4077 $w=2.93e-07 $l=4.2e-07 $layer=LI1_cond $X=1.172 $Y=0.085
+ $X2=1.172 $Y2=0.505
r104 5 36 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.49
+ $Y=0.35 $X2=4.63 $Y2=0.505
r105 4 30 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.35 $X2=3.77 $Y2=0.505
r106 3 26 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.77
+ $Y=0.35 $X2=2.91 $Y2=0.505
r107 2 22 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.35 $X2=2.05 $Y2=0.505
r108 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.35 $X2=1.19 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_8%VPWR 1 8 14
r68 5 14 0.00264757 $w=5.76e-06 $l=1.22e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.88 $Y2=3.208
r69 5 8 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r70 4 8 344.471 $w=1.68e-07 $l=5.28e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=5.52
+ $Y2=3.33
r71 4 5 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 1 14 2.17014e-05 $w=5.76e-06 $l=1e-09 $layer=MET1_cond $X=2.88 $Y=3.207
+ $X2=2.88 $Y2=3.208
.ends

