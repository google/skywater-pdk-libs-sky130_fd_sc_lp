* NGSPICE file created from sky130_fd_sc_lp__nand2b_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand2b_lp A_N B VGND VNB VPB VPWR Y
M1000 a_119_51# A_N a_32_51# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1001 a_277_51# B VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.176e+11p ps=1.4e+06u
M1002 Y a_32_51# a_277_51# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1003 VPWR A_N a_32_51# VPB phighvt w=1e+06u l=250000u
+  ad=6.3e+11p pd=5.26e+06u as=2.85e+11p ps=2.57e+06u
M1004 VPWR a_32_51# Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1005 VGND A_N a_119_51# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

