* NGSPICE file created from sky130_fd_sc_lp__clkbuflp_16.ext - technology: sky130A

.subckt sky130_fd_sc_lp__clkbuflp_16 A VGND VNB VPB VPWR X
M1000 X a_130_417# a_1378_47# VNB nshort w=550000u l=150000u
+  ad=7.7e+11p pd=8.3e+06u as=1.155e+11p ps=1.52e+06u
M1001 X a_130_417# a_2010_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.52e+06u
M1002 a_130_417# A a_110_47# VNB nshort w=550000u l=150000u
+  ad=3.08e+11p pd=3.32e+06u as=1.155e+11p ps=1.52e+06u
M1003 a_1852_47# a_130_417# X VNB nshort w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1004 VPWR a_130_417# X VPB phighvt w=1e+06u l=250000u
+  ad=3.33e+12p pd=3.066e+07u as=2.24e+12p ps=2.048e+07u
M1005 VPWR A a_130_417# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=8.4e+11p ps=7.68e+06u
M1006 X a_130_417# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_584_47# A a_130_417# VNB nshort w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1008 a_2010_47# a_130_417# VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.2265e+12p ps=1.326e+07u
M1009 VGND A a_584_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1378_47# a_130_417# VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_746_47# a_130_417# VGND VNB nshort w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1012 VPWR a_130_417# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_130_417# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_904_47# a_130_417# X VNB nshort w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1015 VGND a_130_417# a_1536_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.52e+06u
M1016 VPWR A a_130_417# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_130_417# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_110_47# A VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_130_417# a_904_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_130_417# a_2168_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.52e+06u
M1021 VGND A a_268_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.52e+06u
M1022 X a_130_417# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_130_417# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1062_47# a_130_417# VGND VNB nshort w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1025 a_130_417# A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_130_417# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_130_417# a_1062_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1220_47# a_130_417# X VNB nshort w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1029 VPWR A a_130_417# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1536_47# a_130_417# X VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_130_417# a_1220_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2168_47# a_130_417# X VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_268_47# A a_130_417# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1694_47# a_130_417# VGND VNB nshort w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1035 a_426_47# A VGND VNB nshort w=550000u l=150000u
+  ad=1.155e+11p pd=1.52e+06u as=0p ps=0u
M1036 X a_130_417# a_1694_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 X a_130_417# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_130_417# A a_426_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 X a_130_417# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VGND a_130_417# a_1852_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VPWR a_130_417# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR a_130_417# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VPWR a_130_417# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1044 X a_130_417# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1045 X a_130_417# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_130_417# A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_130_417# A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1048 X a_130_417# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1049 X a_130_417# a_746_47# VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

