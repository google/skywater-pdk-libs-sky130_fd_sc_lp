* File: sky130_fd_sc_lp__or4bb_lp.pex.spice
* Created: Wed Sep  2 10:33:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%A_86_21# 1 2 3 12 14 15 18 22 25 27 30 33
+ 34 35 36 37 38 39 42 44 47 48 51 53
c135 22 0 2.07706e-19 $X=0.935 $Y=2.545
c136 18 0 1.89361e-19 $X=0.865 $Y=0.445
r137 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.965
+ $Y=1.29 $X2=0.965 $Y2=1.29
r138 45 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.825 $Y=1.2
+ $X2=3.66 $Y2=1.2
r139 44 53 12.796 $w=3.48e-07 $l=4.9452e-07 $layer=LI1_cond $X=4.17 $Y=1.2
+ $X2=4.475 $Y2=0.835
r140 44 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.17 $Y=1.2
+ $X2=3.825 $Y2=1.2
r141 40 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=1.285
+ $X2=3.66 $Y2=1.2
r142 40 42 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=3.66 $Y=1.285
+ $X2=3.66 $Y2=2.145
r143 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=1.2
+ $X2=3.66 $Y2=1.2
r144 38 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.495 $Y=1.2
+ $X2=3.2 $Y2=1.2
r145 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.035 $Y=1.115
+ $X2=3.2 $Y2=1.2
r146 36 50 3.14345 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=3.035 $Y=0.945
+ $X2=3.035 $Y2=0.775
r147 36 37 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.035 $Y=0.945
+ $X2=3.035 $Y2=1.115
r148 34 50 4.62272 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.87 $Y=0.86
+ $X2=3.035 $Y2=0.775
r149 34 35 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.87 $Y=0.86
+ $X2=1.945 $Y2=0.86
r150 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.86 $Y=0.945
+ $X2=1.945 $Y2=0.86
r151 32 33 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.86 $Y=0.945
+ $X2=1.86 $Y2=1.125
r152 31 47 4.53113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.13 $Y=1.21
+ $X2=0.992 $Y2=1.21
r153 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.775 $Y=1.21
+ $X2=1.86 $Y2=1.125
r154 30 31 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.775 $Y=1.21
+ $X2=1.13 $Y2=1.21
r155 26 48 56.8556 $w=3.4e-07 $l=3.35e-07 $layer=POLY_cond $X=0.96 $Y=1.625
+ $X2=0.96 $Y2=1.29
r156 26 27 31.7294 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=0.96 $Y=1.625
+ $X2=0.96 $Y2=1.795
r157 24 48 2.54577 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=0.96 $Y=1.275
+ $X2=0.96 $Y2=1.29
r158 24 25 13.339 $w=2.45e-07 $l=7.5e-08 $layer=POLY_cond $X=0.96 $Y=1.275
+ $X2=0.96 $Y2=1.2
r159 22 27 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.935 $Y=2.545
+ $X2=0.935 $Y2=1.795
r160 16 25 13.339 $w=2.45e-07 $l=1.27083e-07 $layer=POLY_cond $X=0.865 $Y=1.125
+ $X2=0.96 $Y2=1.2
r161 16 18 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.865 $Y=1.125
+ $X2=0.865 $Y2=0.445
r162 14 25 12.4685 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.79 $Y=1.2
+ $X2=0.96 $Y2=1.2
r163 14 15 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.79 $Y=1.2
+ $X2=0.58 $Y2=1.2
r164 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.505 $Y=1.125
+ $X2=0.58 $Y2=1.2
r165 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.505 $Y=1.125
+ $X2=0.505 $Y2=0.445
r166 3 42 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.52
+ $Y=2 $X2=3.66 $Y2=2.145
r167 2 53 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.475
+ $Y=0.625 $X2=4.615 $Y2=0.835
r168 1 50 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.625 $X2=3.035 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%C_N 1 3 6 8 9 10 12 14 15 16 23
c57 16 0 1.44264e-19 $X=1.68 $Y=1.665
c58 8 0 7.13669e-20 $X=1.58 $Y=0.805
c59 6 0 1.92937e-19 $X=1.465 $Y=2.545
r60 21 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.565 $Y=1.64
+ $X2=1.655 $Y2=1.64
r61 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.64 $X2=1.565 $Y2=1.64
r62 18 21 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.465 $Y=1.64
+ $X2=1.565 $Y2=1.64
r63 16 22 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.64
+ $X2=1.565 $Y2=1.64
r64 14 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.655 $Y=1.475
+ $X2=1.655 $Y2=1.64
r65 13 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.655 $Y=0.88
+ $X2=1.655 $Y2=0.805
r66 13 14 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=1.655 $Y=0.88
+ $X2=1.655 $Y2=1.475
r67 10 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.655 $Y=0.73
+ $X2=1.655 $Y2=0.805
r68 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.655 $Y=0.73
+ $X2=1.655 $Y2=0.445
r69 8 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.58 $Y=0.805
+ $X2=1.655 $Y2=0.805
r70 8 9 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.58 $Y=0.805 $X2=1.37
+ $Y2=0.805
r71 4 18 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.805
+ $X2=1.465 $Y2=1.64
r72 4 6 183.856 $w=2.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.465 $Y=1.805
+ $X2=1.465 $Y2=2.545
r73 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.295 $Y=0.73
+ $X2=1.37 $Y2=0.805
r74 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.295 $Y=0.73 $X2=1.295
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%A_318_409# 1 2 7 8 9 11 13 16 18 19 22 25
+ 30 31 32 34 35 38 41 43 45 47 48 50 53
c140 53 0 8.04151e-20 $X=2.2 $Y=1.98
c141 50 0 6.61614e-20 $X=1.73 $Y=2.19
c142 41 0 1.58002e-19 $X=1.73 $Y=2.9
c143 38 0 1.89361e-19 $X=1.51 $Y=0.775
c144 18 0 6.50612e-20 $X=3.535 $Y=1.46
c145 7 0 1.10516e-19 $X=2.81 $Y=1.85
r146 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.2
+ $Y=1.98 $X2=2.2 $Y2=1.98
r147 50 52 10.0596 $w=5.7e-07 $l=4.7e-07 $layer=LI1_cond $X=1.73 $Y=2.15 $X2=2.2
+ $Y2=2.15
r148 47 48 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=1.05 $Y=2.065
+ $X2=1.22 $Y2=2.065
r149 43 45 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.595 $Y=0.43
+ $X2=1.87 $Y2=0.43
r150 39 50 3.93508 $w=3.3e-07 $l=3.35e-07 $layer=LI1_cond $X=1.73 $Y=2.485
+ $X2=1.73 $Y2=2.15
r151 39 41 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.73 $Y=2.485
+ $X2=1.73 $Y2=2.9
r152 37 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.51 $Y=0.595
+ $X2=1.595 $Y2=0.43
r153 37 38 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.51 $Y=0.595
+ $X2=1.51 $Y2=0.775
r154 35 50 10.1602 $w=5.7e-07 $l=2.0106e-07 $layer=LI1_cond $X=1.565 $Y=2.07
+ $X2=1.73 $Y2=2.15
r155 35 48 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.565 $Y=2.07
+ $X2=1.22 $Y2=2.07
r156 34 47 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.675 $Y=2.06
+ $X2=1.05 $Y2=2.06
r157 31 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.425 $Y=0.86
+ $X2=1.51 $Y2=0.775
r158 31 32 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.425 $Y=0.86
+ $X2=0.675 $Y2=0.86
r159 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.59 $Y=1.975
+ $X2=0.675 $Y2=2.06
r160 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.59 $Y=0.945
+ $X2=0.675 $Y2=0.86
r161 29 30 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.59 $Y=0.945
+ $X2=0.59 $Y2=1.975
r162 26 28 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=2.985 $Y=1.46
+ $X2=3.25 $Y2=1.46
r163 24 53 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.2 $Y=1.925
+ $X2=2.2 $Y2=1.98
r164 20 22 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.61 $Y=1.385
+ $X2=3.61 $Y2=0.835
r165 19 28 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.325 $Y=1.46
+ $X2=3.25 $Y2=1.46
r166 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.535 $Y=1.46
+ $X2=3.61 $Y2=1.385
r167 18 19 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.535 $Y=1.46
+ $X2=3.325 $Y2=1.46
r168 14 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.25 $Y=1.385
+ $X2=3.25 $Y2=1.46
r169 14 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.25 $Y=1.385
+ $X2=3.25 $Y2=0.835
r170 13 25 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=2.985 $Y=1.775
+ $X2=2.935 $Y2=1.85
r171 12 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.985 $Y=1.535
+ $X2=2.985 $Y2=1.46
r172 12 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.985 $Y=1.535
+ $X2=2.985 $Y2=1.775
r173 9 25 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=2.935 $Y=1.925
+ $X2=2.935 $Y2=1.85
r174 9 11 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.935 $Y=1.925
+ $X2=2.935 $Y2=2.5
r175 8 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.365 $Y=1.85
+ $X2=2.2 $Y2=1.925
r176 7 25 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.81 $Y=1.85
+ $X2=2.935 $Y2=1.85
r177 7 8 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.81 $Y=1.85
+ $X2=2.365 $Y2=1.85
r178 2 50 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=2.045 $X2=1.73 $Y2=2.19
r179 2 41 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=2.045 $X2=1.73 $Y2=2.9
r180 1 45 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.73
+ $Y=0.235 $X2=1.87 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%A_654_355# 1 2 10 11 12 13 14 15 17 19 20
+ 22 24 26 27 28 32 35 38 40 41 45 47
c115 32 0 6.64046e-20 $X=6.915 $Y=2.16
c116 28 0 6.71696e-20 $X=6.395 $Y=2.49
c117 11 0 1.23206e-19 $X=3.965 $Y=1.85
r118 47 49 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.92 $Y=0.47
+ $X2=6.92 $Y2=0.675
r119 44 45 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.56 $Y=2.24
+ $X2=6.56 $Y2=2.49
r120 41 44 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.56 $Y=2.16 $X2=6.56
+ $Y2=2.24
r121 38 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.52 $Y=2.52
+ $X2=4.52 $Y2=2.685
r122 37 40 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=2.52
+ $X2=4.685 $Y2=2.52
r123 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.52
+ $Y=2.52 $X2=4.52 $Y2=2.52
r124 35 49 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=7 $Y=2.075 $X2=7
+ $Y2=0.675
r125 33 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=2.16
+ $X2=6.56 $Y2=2.16
r126 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.915 $Y=2.16
+ $X2=7 $Y2=2.075
r127 32 33 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.915 $Y=2.16
+ $X2=6.725 $Y2=2.16
r128 28 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=2.49
+ $X2=6.56 $Y2=2.49
r129 28 40 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=6.395 $Y=2.49
+ $X2=4.685 $Y2=2.49
r130 26 52 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.43 $Y=3.075
+ $X2=4.43 $Y2=2.685
r131 22 24 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.4 $Y=1.12 $X2=4.4
+ $Y2=0.835
r132 21 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.115 $Y=1.195
+ $X2=4.04 $Y2=1.195
r133 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.325 $Y=1.195
+ $X2=4.4 $Y2=1.12
r134 20 21 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.325 $Y=1.195
+ $X2=4.115 $Y2=1.195
r135 18 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.04 $Y=1.27
+ $X2=4.04 $Y2=1.195
r136 18 19 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.04 $Y=1.27
+ $X2=4.04 $Y2=1.775
r137 15 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.04 $Y=1.12
+ $X2=4.04 $Y2=1.195
r138 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.04 $Y=1.12
+ $X2=4.04 $Y2=0.835
r139 13 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.355 $Y=3.15
+ $X2=4.43 $Y2=3.075
r140 13 14 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=4.355 $Y=3.15
+ $X2=3.52 $Y2=3.15
r141 11 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.965 $Y=1.85
+ $X2=4.04 $Y2=1.775
r142 11 12 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.965 $Y=1.85
+ $X2=3.52 $Y2=1.85
r143 8 14 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=3.395 $Y=3.075
+ $X2=3.52 $Y2=3.15
r144 8 10 142.861 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.395 $Y=3.075
+ $X2=3.395 $Y2=2.5
r145 7 12 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=3.395 $Y=1.925
+ $X2=3.52 $Y2=1.85
r146 7 10 142.861 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.395 $Y=1.925
+ $X2=3.395 $Y2=2.5
r147 2 44 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.42
+ $Y=2.095 $X2=6.56 $Y2=2.24
r148 1 47 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=6.78
+ $Y=0.235 $X2=6.92 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%B 1 3 5 6 8 9 10 12 15 17 18
c61 18 0 1.23206e-19 $X=4.56 $Y=2.035
c62 8 0 6.71696e-20 $X=5.13 $Y=1.89
c63 5 0 1.43155e-19 $X=4.83 $Y=1.815
r64 18 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.52
+ $Y=1.98 $X2=4.52 $Y2=1.98
r65 13 15 156.526 $w=2.5e-07 $l=6.3e-07 $layer=POLY_cond $X=5.255 $Y=1.965
+ $X2=5.255 $Y2=2.595
r66 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.19 $Y=1.12 $X2=5.19
+ $Y2=0.835
r67 8 13 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=5.13 $Y=1.89
+ $X2=5.255 $Y2=1.965
r68 8 9 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=5.13 $Y=1.89
+ $X2=4.905 $Y2=1.89
r69 7 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.905 $Y=1.195
+ $X2=4.83 $Y2=1.195
r70 6 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.115 $Y=1.195
+ $X2=5.19 $Y2=1.12
r71 6 7 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.115 $Y=1.195
+ $X2=4.905 $Y2=1.195
r72 5 9 22.3869 $w=2.58e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.83 $Y=1.815
+ $X2=4.905 $Y2=1.89
r73 5 21 57.9147 $w=2.58e-07 $l=3.83732e-07 $layer=POLY_cond $X=4.83 $Y=1.815
+ $X2=4.52 $Y2=1.98
r74 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.83 $Y=1.27 $X2=4.83
+ $Y2=1.195
r75 4 5 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.83 $Y=1.27 $X2=4.83
+ $Y2=1.815
r76 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.83 $Y=1.12 $X2=4.83
+ $Y2=1.195
r77 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.83 $Y=1.12 $X2=4.83
+ $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%A 3 5 6 9 14 15 18 19
c66 19 0 8.78408e-20 $X=5.755 $Y=1.71
c67 14 0 7.03397e-20 $X=5.78 $Y=1.135
r68 18 21 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.755 $Y=1.71
+ $X2=5.755 $Y2=1.875
r69 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.755 $Y=1.71
+ $X2=5.755 $Y2=1.545
r70 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.755
+ $Y=1.71 $X2=5.755 $Y2=1.71
r71 15 19 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=5.52 $Y=1.71
+ $X2=5.755 $Y2=1.71
r72 14 20 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=5.78 $Y=1.135
+ $X2=5.78 $Y2=1.545
r73 11 14 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.78 $Y=0.255
+ $X2=5.78 $Y2=1.135
r74 9 21 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=5.745 $Y=2.595
+ $X2=5.745 $Y2=1.875
r75 5 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.705 $Y=0.18
+ $X2=5.78 $Y2=0.255
r76 5 6 1440.87 $w=1.5e-07 $l=2.81e-06 $layer=POLY_cond $X=5.705 $Y=0.18
+ $X2=2.895 $Y2=0.18
r77 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.82 $Y=0.255
+ $X2=2.895 $Y2=0.18
r78 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.82 $Y=0.255 $X2=2.82
+ $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%D_N 1 3 7 11 13 14
c37 13 0 7.03397e-20 $X=6.48 $Y=1.295
c38 7 0 1.54392e-19 $X=6.345 $Y=0.445
c39 3 0 6.64046e-20 $X=6.295 $Y=2.595
c40 1 0 8.78408e-20 $X=6.295 $Y=1.905
r41 13 14 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.56 $Y=1.275
+ $X2=6.56 $Y2=1.665
r42 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.56
+ $Y=1.275 $X2=6.56 $Y2=1.275
r43 9 18 35.2629 $w=2.34e-07 $l=3.01413e-07 $layer=POLY_cond $X=6.705 $Y=1.11
+ $X2=6.475 $Y2=1.275
r44 9 11 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=6.705 $Y=1.11
+ $X2=6.705 $Y2=0.445
r45 5 18 35.2629 $w=2.34e-07 $l=2.20624e-07 $layer=POLY_cond $X=6.345 $Y=1.11
+ $X2=6.475 $Y2=1.275
r46 5 7 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=6.345 $Y=1.11
+ $X2=6.345 $Y2=0.445
r47 1 18 75.1946 $w=4.69e-07 $l=7.14353e-07 $layer=POLY_cond $X=6.295 $Y=1.905
+ $X2=6.475 $Y2=1.275
r48 1 3 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.295 $Y=1.905
+ $X2=6.295 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%X 1 2 7 8 9 10 11 12 13 40 43
c23 43 0 1.92937e-19 $X=0.24 $Y=2.405
r24 43 44 8.25644 $w=7.08e-07 $l=8e-08 $layer=LI1_cond $X=0.48 $Y=2.405 $X2=0.48
+ $Y2=2.325
r25 23 35 3.66692 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.225 $Y=0.595
+ $X2=0.225 $Y2=0.43
r26 13 47 4.80116 $w=7.08e-07 $l=2.85e-07 $layer=LI1_cond $X=0.48 $Y=2.775
+ $X2=0.48 $Y2=2.49
r27 12 47 1.39823 $w=7.08e-07 $l=8.3e-08 $layer=LI1_cond $X=0.48 $Y=2.407
+ $X2=0.48 $Y2=2.49
r28 12 43 0.0336923 $w=7.08e-07 $l=2e-09 $layer=LI1_cond $X=0.48 $Y=2.407
+ $X2=0.48 $Y2=2.405
r29 12 44 0.166364 $w=1.98e-07 $l=3e-09 $layer=LI1_cond $X=0.225 $Y=2.322
+ $X2=0.225 $Y2=2.325
r30 11 12 15.9155 $w=1.98e-07 $l=2.87e-07 $layer=LI1_cond $X=0.225 $Y=2.035
+ $X2=0.225 $Y2=2.322
r31 10 11 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=2.035
r32 9 10 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r33 8 9 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r34 7 40 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.24 $Y=0.43 $X2=0.29
+ $Y2=0.43
r35 7 35 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.24 $Y=0.43
+ $X2=0.225 $Y2=0.43
r36 7 8 17.08 $w=1.98e-07 $l=3.08e-07 $layer=LI1_cond $X=0.225 $Y=0.617
+ $X2=0.225 $Y2=0.925
r37 7 23 1.22 $w=1.98e-07 $l=2.2e-08 $layer=LI1_cond $X=0.225 $Y=0.617 $X2=0.225
+ $Y2=0.595
r38 2 47 300 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_PDIFF $count=2 $X=0.525
+ $Y=2.045 $X2=0.67 $Y2=2.49
r39 1 40 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.235 $X2=0.29 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%VPWR 1 2 9 13 15 17 22 32 33 36 39
c58 22 0 1.26713e-20 $X=5.845 $Y=3.33
c59 9 0 8.04151e-20 $X=1.2 $Y=2.5
r60 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r61 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r62 33 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33 $X2=6
+ $Y2=3.33
r63 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r64 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.01 $Y2=3.33
r65 30 32 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.96 $Y2=3.33
r66 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r67 28 29 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r68 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 25 28 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=5.52 $Y2=3.33
r70 25 26 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.2 $Y2=3.33
r72 23 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.365 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6.01 $Y2=3.33
r74 22 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r76 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.2 $Y2=3.33
r78 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 15 29 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r80 15 26 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=1.68 $Y2=3.33
r81 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=3.33
r82 11 13 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=2.935
r83 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=3.245 $X2=1.2
+ $Y2=3.33
r84 7 9 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=1.2 $Y=3.245 $X2=1.2
+ $Y2=2.5
r85 2 13 600 $w=1.7e-07 $l=9.07304e-07 $layer=licon1_PDIFF $count=1 $X=5.87
+ $Y=2.095 $X2=6.01 $Y2=2.935
r86 1 9 300 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=2.045 $X2=1.2 $Y2=2.5
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%A_505_400# 1 2 9 12
r30 12 14 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.67 $Y=2.85 $X2=2.67
+ $Y2=2.95
r31 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=2.95
+ $X2=2.67 $Y2=2.95
r32 7 9 140.594 $w=1.68e-07 $l=2.155e-06 $layer=LI1_cond $X=2.835 $Y=2.95
+ $X2=4.99 $Y2=2.95
r33 2 9 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.845
+ $Y=2.095 $X2=4.99 $Y2=2.95
r34 1 12 600 $w=1.7e-07 $l=9.19647e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=2 $X2=2.67 $Y2=2.85
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%VGND 1 2 3 4 15 19 23 25 29 32 33 34 36 45
+ 54 55 58 61 64
c86 32 0 7.13669e-20 $X=3.66 $Y=0
c87 23 0 2.97547e-19 $X=5.485 $Y=0.77
r88 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r89 62 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r90 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r91 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 55 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6
+ $Y2=0
r93 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r94 52 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.13
+ $Y2=0
r95 52 54 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.96
+ $Y2=0
r96 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r97 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r98 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r99 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r100 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r101 45 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.485
+ $Y2=0
r102 45 50 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.04
+ $Y2=0
r103 41 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.08
+ $Y2=0
r104 41 43 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=1.245 $Y=0
+ $X2=3.6 $Y2=0
r105 39 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r106 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r107 36 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.08
+ $Y2=0
r108 36 38 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=0.915 $Y=0
+ $X2=0.72 $Y2=0
r109 34 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r110 34 59 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=1.2
+ $Y2=0
r111 34 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r112 32 43 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.66 $Y=0 $X2=3.6
+ $Y2=0
r113 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.66 $Y=0 $X2=3.825
+ $Y2=0
r114 31 47 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.99 $Y=0 $X2=4.08
+ $Y2=0
r115 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=0 $X2=3.825
+ $Y2=0
r116 27 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0
r117 27 29 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.13 $Y=0.085
+ $X2=6.13 $Y2=0.445
r118 26 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.65 $Y=0 $X2=5.485
+ $Y2=0
r119 25 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.965 $Y=0 $X2=6.13
+ $Y2=0
r120 25 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.965 $Y=0
+ $X2=5.65 $Y2=0
r121 21 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.485 $Y=0.085
+ $X2=5.485 $Y2=0
r122 21 23 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=5.485 $Y=0.085
+ $X2=5.485 $Y2=0.77
r123 17 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=0.085
+ $X2=3.825 $Y2=0
r124 17 19 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=3.825 $Y=0.085
+ $X2=3.825 $Y2=0.77
r125 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=0.085
+ $X2=1.08 $Y2=0
r126 13 15 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.08 $Y=0.085
+ $X2=1.08 $Y2=0.405
r127 4 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.985
+ $Y=0.235 $X2=6.13 $Y2=0.445
r128 3 23 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=5.265
+ $Y=0.625 $X2=5.485 $Y2=0.77
r129 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.685
+ $Y=0.625 $X2=3.825 $Y2=0.77
r130 1 15 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.235 $X2=1.08 $Y2=0.405
.ends

.subckt PM_SKY130_FD_SC_LP__OR4BB_LP%A_476_125# 1 2 9 12 13 14 16 17 18 20 21 22
+ 24 26 28
c111 18 0 6.50612e-20 $X=4.175 $Y=1.55
c112 13 0 1.23187e-19 $X=4.005 $Y=2.495
r113 28 30 10.5346 $w=3.83e-07 $l=2.3e-07 $layer=LI1_cond $X=6.022 $Y=1.135
+ $X2=6.022 $Y2=1.365
r114 25 26 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.537 $Y=1.465
+ $X2=2.537 $Y2=1.635
r115 24 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.13 $Y=2.055
+ $X2=6.13 $Y2=1.365
r116 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.045 $Y=2.14
+ $X2=6.13 $Y2=2.055
r117 21 22 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=6.045 $Y=2.14
+ $X2=5.035 $Y2=2.14
r118 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.95 $Y=2.055
+ $X2=5.035 $Y2=2.14
r119 19 20 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.95 $Y=1.635
+ $X2=4.95 $Y2=2.055
r120 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.865 $Y=1.55
+ $X2=4.95 $Y2=1.635
r121 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.865 $Y=1.55
+ $X2=4.175 $Y2=1.55
r122 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.09 $Y=1.635
+ $X2=4.175 $Y2=1.55
r123 15 16 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=4.09 $Y=1.635
+ $X2=4.09 $Y2=2.41
r124 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.005 $Y=2.495
+ $X2=4.09 $Y2=2.41
r125 13 14 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.005 $Y=2.495
+ $X2=2.715 $Y2=2.495
r126 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.63 $Y=2.41
+ $X2=2.715 $Y2=2.495
r127 12 26 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.63 $Y=2.41
+ $X2=2.63 $Y2=1.635
r128 9 25 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.525 $Y=1.29
+ $X2=2.525 $Y2=1.465
r129 2 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.855
+ $Y=0.925 $X2=5.995 $Y2=1.135
r130 1 9 182 $w=1.7e-07 $l=7.33928e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.625 $X2=2.525 $Y2=1.29
.ends

