# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__nand4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.210000 0.865000 1.750000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.210000 1.285000 1.750000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.270000 1.200000 8.005000 1.515000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.210000 1.200000 9.925000 1.515000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.292800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.145000 0.955000 3.690000 1.215000 ;
        RECT 2.345000 1.775000 9.485000 1.945000 ;
        RECT 2.345000 1.945000 2.535000 3.075000 ;
        RECT 3.205000 1.945000 3.425000 3.075000 ;
        RECT 3.520000 1.215000 3.690000 1.775000 ;
        RECT 3.995000 1.945000 6.085000 2.120000 ;
        RECT 3.995000 2.120000 4.255000 3.075000 ;
        RECT 4.925000 2.120000 6.085000 2.160000 ;
        RECT 4.925000 2.160000 5.115000 3.075000 ;
        RECT 6.255000 1.685000 9.485000 1.775000 ;
        RECT 6.645000 1.945000 6.875000 3.075000 ;
        RECT 7.545000 1.945000 7.735000 3.075000 ;
        RECT 8.405000 1.945000 8.595000 3.075000 ;
        RECT 9.265000 1.945000 9.485000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.085000  0.325000  0.460000 1.040000 ;
      RECT 0.085000  1.040000  0.275000 1.930000 ;
      RECT 0.085000  1.930000  0.450000 2.340000 ;
      RECT 0.085000  2.340000  2.020000 2.510000 ;
      RECT 0.085000  2.510000  0.450000 2.940000 ;
      RECT 0.630000  0.085000  0.960000 1.040000 ;
      RECT 0.630000  2.680000  0.960000 3.245000 ;
      RECT 1.060000  1.920000  1.680000 2.170000 ;
      RECT 1.130000  0.325000  1.330000 0.615000 ;
      RECT 1.130000  0.615000  4.040000 0.785000 ;
      RECT 1.130000  0.785000  1.330000 1.040000 ;
      RECT 1.500000  0.785000  1.680000 1.920000 ;
      RECT 1.600000  0.255000  5.760000 0.425000 ;
      RECT 1.600000  0.425000  4.945000 0.445000 ;
      RECT 1.845000  2.680000  2.175000 3.245000 ;
      RECT 1.850000  1.385000  3.340000 1.605000 ;
      RECT 1.850000  1.605000  2.020000 2.340000 ;
      RECT 2.705000  2.115000  3.035000 3.245000 ;
      RECT 3.595000  2.115000  3.825000 3.245000 ;
      RECT 3.870000  0.785000  4.040000 1.415000 ;
      RECT 3.870000  1.415000  5.900000 1.605000 ;
      RECT 4.245000  0.885000  4.445000 1.055000 ;
      RECT 4.245000  1.055000  6.100000 1.245000 ;
      RECT 4.425000  2.290000  4.755000 3.245000 ;
      RECT 4.615000  0.445000  4.945000 0.885000 ;
      RECT 5.115000  0.860000  5.305000 0.960000 ;
      RECT 5.115000  0.960000  6.100000 1.055000 ;
      RECT 5.285000  2.330000  6.475000 3.245000 ;
      RECT 5.475000  0.425000  5.760000 0.790000 ;
      RECT 5.930000  0.310000  7.775000 0.520000 ;
      RECT 5.930000  0.520000  6.100000 0.960000 ;
      RECT 6.255000  2.125000  6.475000 2.330000 ;
      RECT 6.280000  0.700000  7.345000 0.860000 ;
      RECT 6.280000  0.860000  9.925000 1.030000 ;
      RECT 7.045000  2.115000  7.375000 3.245000 ;
      RECT 7.515000  0.520000  7.775000 0.690000 ;
      RECT 7.905000  2.115000  8.235000 3.245000 ;
      RECT 7.995000  0.255000  8.195000 0.860000 ;
      RECT 8.365000  0.085000  8.695000 0.690000 ;
      RECT 8.765000  2.115000  9.095000 3.245000 ;
      RECT 8.865000  0.255000  9.045000 0.860000 ;
      RECT 9.225000  0.085000  9.555000 0.690000 ;
      RECT 9.655000  1.815000  9.955000 3.245000 ;
      RECT 9.725000  0.255000  9.925000 0.860000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__nand4bb_4
END LIBRARY
