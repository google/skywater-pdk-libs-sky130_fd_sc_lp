* NGSPICE file created from sky130_fd_sc_lp__o211ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 VGND A1 a_286_65# VNB nshort w=840000u l=150000u
+  ad=6.804e+11p pd=6.66e+06u as=7.056e+11p ps=6.72e+06u
M1001 VPWR A1 a_487_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3734e+12p pd=1.226e+07u as=1.0206e+12p ps=9.18e+06u
M1002 a_286_65# B1 a_31_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=6.804e+11p ps=6.66e+06u
M1003 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.0584e+12p ps=9.24e+06u
M1004 a_487_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_286_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_31_65# B1 a_286_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_487_367# A2 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y C1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y C1 a_31_65# VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1010 a_31_65# C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_286_65# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A2 a_487_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_286_65# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

