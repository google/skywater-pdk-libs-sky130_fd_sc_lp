* File: sky130_fd_sc_lp__clkinvlp_16.pxi.spice
* Created: Wed Sep  2 09:41:05 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINVLP_16%A N_A_M1025_g N_A_M1000_g N_A_M1001_g
+ N_A_M1002_g N_A_M1005_g N_A_M1003_g N_A_M1004_g N_A_M1010_g N_A_M1007_g
+ N_A_M1006_g N_A_M1009_g N_A_M1008_g N_A_M1011_g N_A_M1031_g N_A_M1015_g
+ N_A_M1012_g N_A_M1013_g N_A_M1016_g N_A_M1014_g N_A_M1017_g N_A_M1024_g
+ N_A_M1019_g N_A_M1021_g N_A_M1018_g N_A_M1022_g N_A_M1020_g N_A_M1023_g
+ N_A_M1027_g N_A_M1026_g N_A_M1029_g N_A_M1028_g N_A_M1030_g N_A_M1032_g
+ N_A_M1034_g N_A_M1033_g N_A_c_167_n N_A_M1035_g A N_A_c_169_n N_A_c_170_n
+ N_A_c_171_n N_A_c_172_n N_A_c_173_n N_A_c_174_n N_A_c_175_n
+ PM_SKY130_FD_SC_LP__CLKINVLP_16%A
x_PM_SKY130_FD_SC_LP__CLKINVLP_16%VPWR N_VPWR_M1000_s N_VPWR_M1002_s
+ N_VPWR_M1007_s N_VPWR_M1011_s N_VPWR_M1016_s N_VPWR_M1021_s N_VPWR_M1023_s
+ N_VPWR_M1030_s N_VPWR_M1035_s N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n
+ N_VPWR_c_518_n N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n
+ N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n
+ N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n
+ N_VPWR_c_533_n VPWR N_VPWR_c_534_n N_VPWR_c_535_n N_VPWR_c_536_n
+ N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n N_VPWR_c_514_n
+ VPWR PM_SKY130_FD_SC_LP__CLKINVLP_16%VPWR
x_PM_SKY130_FD_SC_LP__CLKINVLP_16%Y N_Y_M1001_s N_Y_M1006_s N_Y_M1013_s
+ N_Y_M1018_s N_Y_M1028_s N_Y_M1000_d N_Y_M1003_d N_Y_M1009_d N_Y_M1012_d
+ N_Y_M1017_d N_Y_M1022_d N_Y_M1029_d N_Y_M1034_d N_Y_c_675_n N_Y_c_705_n
+ N_Y_c_713_n N_Y_c_720_n N_Y_c_683_n N_Y_c_730_n N_Y_c_684_n N_Y_c_676_n
+ N_Y_c_677_n N_Y_c_686_n N_Y_c_678_n N_Y_c_679_n N_Y_c_680_n N_Y_c_681_n Y
+ N_Y_c_688_n N_Y_c_689_n N_Y_c_690_n N_Y_c_691_n N_Y_c_692_n N_Y_c_693_n
+ N_Y_c_694_n N_Y_c_695_n N_Y_c_696_n N_Y_c_682_n
+ PM_SKY130_FD_SC_LP__CLKINVLP_16%Y
x_PM_SKY130_FD_SC_LP__CLKINVLP_16%VGND N_VGND_M1025_d N_VGND_M1004_d
+ N_VGND_M1031_d N_VGND_M1024_d N_VGND_M1027_d N_VGND_M1033_d N_VGND_c_919_n
+ N_VGND_c_920_n N_VGND_c_921_n N_VGND_c_922_n N_VGND_c_923_n N_VGND_c_924_n
+ N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n N_VGND_c_928_n N_VGND_c_929_n
+ VGND N_VGND_c_930_n N_VGND_c_931_n N_VGND_c_932_n N_VGND_c_933_n
+ N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n N_VGND_c_937_n VGND
+ PM_SKY130_FD_SC_LP__CLKINVLP_16%VGND
cc_1 VNB N_A_M1025_g 0.0367769f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.61
cc_2 VNB N_A_M1000_g 0.00506355f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.48
cc_3 VNB N_A_M1001_g 0.025148f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.61
cc_4 VNB N_A_M1002_g 0.00544189f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.48
cc_5 VNB N_A_M1005_g 0.0270661f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=0.61
cc_6 VNB N_A_M1003_g 0.00546844f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=2.48
cc_7 VNB N_A_M1004_g 0.0266529f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=0.61
cc_8 VNB N_A_M1010_g 0.026629f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=0.61
cc_9 VNB N_A_M1007_g 0.00546743f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=2.48
cc_10 VNB N_A_M1006_g 0.0259642f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=0.61
cc_11 VNB N_A_M1009_g 0.00509865f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.48
cc_12 VNB N_A_M1008_g 0.025945f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=0.61
cc_13 VNB N_A_M1011_g 0.00509672f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.48
cc_14 VNB N_A_M1031_g 0.0266457f $X=-0.19 $Y=-0.245 $X2=3.205 $Y2=0.61
cc_15 VNB N_A_M1015_g 0.0266475f $X=-0.19 $Y=-0.245 $X2=3.635 $Y2=0.61
cc_16 VNB N_A_M1012_g 0.00543915f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=2.48
cc_17 VNB N_A_M1013_g 0.0259447f $X=-0.19 $Y=-0.245 $X2=3.995 $Y2=0.61
cc_18 VNB N_A_M1016_g 0.00509865f $X=-0.19 $Y=-0.245 $X2=4.235 $Y2=2.48
cc_19 VNB N_A_M1014_g 0.0259642f $X=-0.19 $Y=-0.245 $X2=4.425 $Y2=0.61
cc_20 VNB N_A_M1017_g 0.00546743f $X=-0.19 $Y=-0.245 $X2=4.765 $Y2=2.48
cc_21 VNB N_A_M1024_g 0.026639f $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=0.61
cc_22 VNB N_A_M1019_g 0.026629f $X=-0.19 $Y=-0.245 $X2=5.215 $Y2=0.61
cc_23 VNB N_A_M1021_g 0.00546666f $X=-0.19 $Y=-0.245 $X2=5.295 $Y2=2.48
cc_24 VNB N_A_M1018_g 0.0259642f $X=-0.19 $Y=-0.245 $X2=5.575 $Y2=0.61
cc_25 VNB N_A_M1022_g 0.00509865f $X=-0.19 $Y=-0.245 $X2=5.825 $Y2=2.48
cc_26 VNB N_A_M1020_g 0.0259552f $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=0.61
cc_27 VNB N_A_M1023_g 0.00543887f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=2.48
cc_28 VNB N_A_M1027_g 0.0266415f $X=-0.19 $Y=-0.245 $X2=6.365 $Y2=0.61
cc_29 VNB N_A_M1026_g 0.0266488f $X=-0.19 $Y=-0.245 $X2=6.795 $Y2=0.61
cc_30 VNB N_A_M1029_g 0.00509657f $X=-0.19 $Y=-0.245 $X2=6.885 $Y2=2.48
cc_31 VNB N_A_M1028_g 0.0259552f $X=-0.19 $Y=-0.245 $X2=7.155 $Y2=0.61
cc_32 VNB N_A_M1030_g 0.00509865f $X=-0.19 $Y=-0.245 $X2=7.415 $Y2=2.48
cc_33 VNB N_A_M1032_g 0.0259539f $X=-0.19 $Y=-0.245 $X2=7.585 $Y2=0.61
cc_34 VNB N_A_M1034_g 0.00546743f $X=-0.19 $Y=-0.245 $X2=7.945 $Y2=2.48
cc_35 VNB N_A_M1033_g 0.0381984f $X=-0.19 $Y=-0.245 $X2=7.945 $Y2=0.61
cc_36 VNB N_A_c_167_n 0.435692f $X=-0.19 $Y=-0.245 $X2=8.475 $Y2=1.565
cc_37 VNB N_A_M1035_g 0.0083313f $X=-0.19 $Y=-0.245 $X2=8.475 $Y2=2.48
cc_38 VNB N_A_c_169_n 0.00214937f $X=-0.19 $Y=-0.245 $X2=3.44 $Y2=1.4
cc_39 VNB N_A_c_170_n 0.0186424f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.295
cc_40 VNB N_A_c_171_n 0.00973245f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.295
cc_41 VNB N_A_c_172_n 0.00538664f $X=-0.19 $Y=-0.245 $X2=5.04 $Y2=1.295
cc_42 VNB N_A_c_173_n 0.00322887f $X=-0.19 $Y=-0.245 $X2=6.48 $Y2=1.295
cc_43 VNB N_A_c_174_n 0.0293078f $X=-0.19 $Y=-0.245 $X2=8.4 $Y2=1.295
cc_44 VNB N_A_c_175_n 0.108638f $X=-0.19 $Y=-0.245 $X2=8.4 $Y2=1.295
cc_45 VNB N_VPWR_c_514_n 0.382608f $X=-0.19 $Y=-0.245 $X2=7.945 $Y2=0.61
cc_46 VNB N_Y_c_675_n 0.00664871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_676_n 0.00240513f $X=-0.19 $Y=-0.245 $X2=4.235 $Y2=2.48
cc_48 VNB N_Y_c_677_n 0.00215056f $X=-0.19 $Y=-0.245 $X2=4.425 $Y2=0.61
cc_49 VNB N_Y_c_678_n 8.48552e-19 $X=-0.19 $Y=-0.245 $X2=4.765 $Y2=2.48
cc_50 VNB N_Y_c_679_n 6.41415e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_Y_c_680_n 0.00155753f $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=0.61
cc_52 VNB N_Y_c_681_n 0.00143153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_Y_c_682_n 8.71722e-19 $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.407
cc_54 VNB N_VGND_c_919_n 0.0111239f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=0.61
cc_55 VNB N_VGND_c_920_n 0.0255575f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=1.565
cc_56 VNB N_VGND_c_921_n 0.00306361f $X=-0.19 $Y=-0.245 $X2=1.625 $Y2=1.235
cc_57 VNB N_VGND_c_922_n 0.00306361f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=1.235
cc_58 VNB N_VGND_c_923_n 0.00306361f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.565
cc_59 VNB N_VGND_c_924_n 0.00306361f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.235
cc_60 VNB N_VGND_c_925_n 0.0254428f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.565
cc_61 VNB N_VGND_c_926_n 0.0368108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_927_n 0.00561514f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=1.235
cc_63 VNB N_VGND_c_928_n 0.0368108f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=0.61
cc_64 VNB N_VGND_c_929_n 0.00589254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_930_n 0.0340009f $X=-0.19 $Y=-0.245 $X2=3.175 $Y2=2.48
cc_66 VNB N_VGND_c_931_n 0.0368108f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=2.48
cc_67 VNB N_VGND_c_932_n 0.0368108f $X=-0.19 $Y=-0.245 $X2=4.235 $Y2=2.48
cc_68 VNB N_VGND_c_933_n 0.0274418f $X=-0.19 $Y=-0.245 $X2=4.785 $Y2=0.61
cc_69 VNB N_VGND_c_934_n 0.546648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_935_n 0.00561514f $X=-0.19 $Y=-0.245 $X2=5.295 $Y2=2.48
cc_71 VNB N_VGND_c_936_n 0.00561514f $X=-0.19 $Y=-0.245 $X2=5.575 $Y2=1.235
cc_72 VNB N_VGND_c_937_n 0.00561514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VPB N_A_M1000_g 0.0434878f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.48
cc_74 VPB N_A_M1002_g 0.0342029f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.48
cc_75 VPB N_A_M1003_g 0.0350066f $X=-0.19 $Y=1.655 $X2=1.585 $Y2=2.48
cc_76 VPB N_A_M1007_g 0.0350057f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.48
cc_77 VPB N_A_M1009_g 0.0339077f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.48
cc_78 VPB N_A_M1011_g 0.0339001f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=2.48
cc_79 VPB N_A_M1012_g 0.0344639f $X=-0.19 $Y=1.655 $X2=3.705 $Y2=2.48
cc_80 VPB N_A_M1016_g 0.0338811f $X=-0.19 $Y=1.655 $X2=4.235 $Y2=2.48
cc_81 VPB N_A_M1017_g 0.0350057f $X=-0.19 $Y=1.655 $X2=4.765 $Y2=2.48
cc_82 VPB N_A_M1021_g 0.0350034f $X=-0.19 $Y=1.655 $X2=5.295 $Y2=2.48
cc_83 VPB N_A_M1022_g 0.033888f $X=-0.19 $Y=1.655 $X2=5.825 $Y2=2.48
cc_84 VPB N_A_M1023_g 0.034747f $X=-0.19 $Y=1.655 $X2=6.355 $Y2=2.48
cc_85 VPB N_A_M1029_g 0.0339008f $X=-0.19 $Y=1.655 $X2=6.885 $Y2=2.48
cc_86 VPB N_A_M1030_g 0.0339077f $X=-0.19 $Y=1.655 $X2=7.415 $Y2=2.48
cc_87 VPB N_A_M1034_g 0.0350057f $X=-0.19 $Y=1.655 $X2=7.945 $Y2=2.48
cc_88 VPB N_A_M1035_g 0.0472476f $X=-0.19 $Y=1.655 $X2=8.475 $Y2=2.48
cc_89 VPB N_A_c_170_n 0.00764565f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.295
cc_90 VPB N_VPWR_c_515_n 0.0112117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_516_n 0.0506365f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=0.61
cc_92 VPB N_VPWR_c_517_n 0.0199224f $X=-0.19 $Y=1.655 $X2=2.115 $Y2=2.48
cc_93 VPB N_VPWR_c_518_n 0.00535062f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=0.61
cc_94 VPB N_VPWR_c_519_n 0.00658911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_520_n 0.00535399f $X=-0.19 $Y=1.655 $X2=3.175 $Y2=2.48
cc_96 VPB N_VPWR_c_521_n 0.00698874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_522_n 0.00661398f $X=-0.19 $Y=1.655 $X2=3.705 $Y2=2.48
cc_98 VPB N_VPWR_c_523_n 0.0196786f $X=-0.19 $Y=1.655 $X2=3.995 $Y2=0.61
cc_99 VPB N_VPWR_c_524_n 0.00572628f $X=-0.19 $Y=1.655 $X2=4.235 $Y2=2.48
cc_100 VPB N_VPWR_c_525_n 0.00636813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_526_n 0.0150395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_527_n 0.0572237f $X=-0.19 $Y=1.655 $X2=4.785 $Y2=0.61
cc_103 VPB N_VPWR_c_528_n 0.0199224f $X=-0.19 $Y=1.655 $X2=5.215 $Y2=0.61
cc_104 VPB N_VPWR_c_529_n 0.00577233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_530_n 0.0199224f $X=-0.19 $Y=1.655 $X2=5.295 $Y2=2.48
cc_106 VPB N_VPWR_c_531_n 0.00577233f $X=-0.19 $Y=1.655 $X2=5.295 $Y2=2.48
cc_107 VPB N_VPWR_c_532_n 0.0199224f $X=-0.19 $Y=1.655 $X2=5.575 $Y2=1.235
cc_108 VPB N_VPWR_c_533_n 0.00577233f $X=-0.19 $Y=1.655 $X2=5.575 $Y2=0.61
cc_109 VPB N_VPWR_c_534_n 0.0199224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_535_n 0.0199224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_536_n 0.0199224f $X=-0.19 $Y=1.655 $X2=6.885 $Y2=1.565
cc_112 VPB N_VPWR_c_537_n 0.00577233f $X=-0.19 $Y=1.655 $X2=7.415 $Y2=1.565
cc_113 VPB N_VPWR_c_538_n 0.00577233f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_539_n 0.00577233f $X=-0.19 $Y=1.655 $X2=7.585 $Y2=0.61
cc_115 VPB N_VPWR_c_540_n 0.00577233f $X=-0.19 $Y=1.655 $X2=7.945 $Y2=2.48
cc_116 VPB N_VPWR_c_514_n 0.0653573f $X=-0.19 $Y=1.655 $X2=7.945 $Y2=0.61
cc_117 VPB N_Y_c_683_n 0.00232136f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_Y_c_684_n 3.86553e-19 $X=-0.19 $Y=1.655 $X2=4.235 $Y2=2.48
cc_119 VPB N_Y_c_676_n 7.58544e-19 $X=-0.19 $Y=1.655 $X2=4.235 $Y2=2.48
cc_120 VPB N_Y_c_686_n 8.36639e-19 $X=-0.19 $Y=1.655 $X2=4.765 $Y2=1.565
cc_121 VPB N_Y_c_678_n 0.00142061f $X=-0.19 $Y=1.655 $X2=4.765 $Y2=2.48
cc_122 VPB N_Y_c_688_n 0.00232136f $X=-0.19 $Y=1.655 $X2=5.575 $Y2=1.235
cc_123 VPB N_Y_c_689_n 0.00408178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_Y_c_690_n 0.00232136f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_Y_c_691_n 0.00232136f $X=-0.19 $Y=1.655 $X2=6.795 $Y2=0.61
cc_126 VPB N_Y_c_692_n 0.00408178f $X=-0.19 $Y=1.655 $X2=7.155 $Y2=0.61
cc_127 VPB N_Y_c_693_n 0.00232136f $X=-0.19 $Y=1.655 $X2=7.585 $Y2=0.61
cc_128 VPB N_Y_c_694_n 0.00408542f $X=-0.19 $Y=1.655 $X2=7.945 $Y2=1.235
cc_129 VPB N_Y_c_695_n 0.0216583f $X=-0.19 $Y=1.655 $X2=7.945 $Y2=0.61
cc_130 VPB N_Y_c_696_n 7.21307e-19 $X=-0.19 $Y=1.655 $X2=0.075 $Y2=1.18
cc_131 VPB N_Y_c_682_n 0.00212119f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.407
cc_132 N_A_M1000_g N_VPWR_c_516_n 0.0234272f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_133 N_A_M1002_g N_VPWR_c_516_n 8.05893e-19 $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_134 N_A_c_167_n N_VPWR_c_516_n 0.00122665f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_135 N_A_c_170_n N_VPWR_c_516_n 0.0278519f $X=0.24 $Y=1.295 $X2=0 $Y2=0
cc_136 N_A_c_175_n N_VPWR_c_516_n 0.00150998f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_137 N_A_M1000_g N_VPWR_c_517_n 0.00687065f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_138 N_A_M1002_g N_VPWR_c_517_n 0.00687065f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_139 N_A_M1000_g N_VPWR_c_518_n 8.69657e-19 $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_140 N_A_M1002_g N_VPWR_c_518_n 0.0212636f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_141 N_A_M1003_g N_VPWR_c_518_n 0.0212636f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_142 N_A_M1007_g N_VPWR_c_518_n 8.69657e-19 $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_143 N_A_c_167_n N_VPWR_c_518_n 5.19494e-19 $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_144 N_A_c_171_n N_VPWR_c_518_n 0.00887565f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_145 N_A_c_175_n N_VPWR_c_518_n 3.69173e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_146 N_A_M1003_g N_VPWR_c_519_n 8.69657e-19 $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_147 N_A_M1007_g N_VPWR_c_519_n 0.0212636f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_148 N_A_M1009_g N_VPWR_c_519_n 0.0212642f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_149 N_A_M1011_g N_VPWR_c_519_n 8.69657e-19 $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_150 N_A_c_167_n N_VPWR_c_519_n 0.00300581f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_151 N_A_c_171_n N_VPWR_c_519_n 0.00123069f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_152 N_A_c_175_n N_VPWR_c_519_n 0.00126121f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_153 N_A_M1009_g N_VPWR_c_520_n 8.69657e-19 $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_154 N_A_M1011_g N_VPWR_c_520_n 0.0212642f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_155 N_A_M1012_g N_VPWR_c_520_n 0.0212642f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_156 N_A_M1016_g N_VPWR_c_520_n 8.71352e-19 $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_157 N_A_c_167_n N_VPWR_c_520_n 0.00190552f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_158 N_A_c_169_n N_VPWR_c_520_n 0.00884676f $X=3.44 $Y=1.4 $X2=0 $Y2=0
cc_159 N_A_c_175_n N_VPWR_c_520_n 3.69624e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_160 N_A_M1012_g N_VPWR_c_521_n 8.71352e-19 $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_161 N_A_M1016_g N_VPWR_c_521_n 0.0212636f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_162 N_A_M1017_g N_VPWR_c_521_n 0.0214005f $X=4.765 $Y=2.48 $X2=0 $Y2=0
cc_163 N_A_M1021_g N_VPWR_c_521_n 8.69657e-19 $X=5.295 $Y=2.48 $X2=0 $Y2=0
cc_164 N_A_c_167_n N_VPWR_c_521_n 0.00300581f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_165 N_A_c_175_n N_VPWR_c_521_n 0.00171827f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_166 N_A_M1017_g N_VPWR_c_522_n 8.69657e-19 $X=4.765 $Y=2.48 $X2=0 $Y2=0
cc_167 N_A_M1021_g N_VPWR_c_522_n 0.0214689f $X=5.295 $Y=2.48 $X2=0 $Y2=0
cc_168 N_A_M1022_g N_VPWR_c_522_n 0.0200381f $X=5.825 $Y=2.48 $X2=0 $Y2=0
cc_169 N_A_M1023_g N_VPWR_c_522_n 8.23274e-19 $X=6.355 $Y=2.48 $X2=0 $Y2=0
cc_170 N_A_c_167_n N_VPWR_c_522_n 0.00300581f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_171 N_A_c_175_n N_VPWR_c_522_n 0.00153217f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_172 N_A_M1022_g N_VPWR_c_523_n 0.00651431f $X=5.825 $Y=2.48 $X2=0 $Y2=0
cc_173 N_A_M1023_g N_VPWR_c_523_n 0.00687065f $X=6.355 $Y=2.48 $X2=0 $Y2=0
cc_174 N_A_M1022_g N_VPWR_c_524_n 8.69657e-19 $X=5.825 $Y=2.48 $X2=0 $Y2=0
cc_175 N_A_M1023_g N_VPWR_c_524_n 0.0212636f $X=6.355 $Y=2.48 $X2=0 $Y2=0
cc_176 N_A_M1029_g N_VPWR_c_524_n 0.0214689f $X=6.885 $Y=2.48 $X2=0 $Y2=0
cc_177 N_A_M1030_g N_VPWR_c_524_n 8.69657e-19 $X=7.415 $Y=2.48 $X2=0 $Y2=0
cc_178 N_A_c_167_n N_VPWR_c_524_n 5.22715e-19 $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_179 N_A_c_173_n N_VPWR_c_524_n 0.00662199f $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_180 N_A_c_175_n N_VPWR_c_524_n 8.93042e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_181 N_A_M1029_g N_VPWR_c_525_n 8.69657e-19 $X=6.885 $Y=2.48 $X2=0 $Y2=0
cc_182 N_A_M1030_g N_VPWR_c_525_n 0.0213069f $X=7.415 $Y=2.48 $X2=0 $Y2=0
cc_183 N_A_M1034_g N_VPWR_c_525_n 0.0212642f $X=7.945 $Y=2.48 $X2=0 $Y2=0
cc_184 N_A_c_167_n N_VPWR_c_525_n 0.00279289f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_185 N_A_M1035_g N_VPWR_c_525_n 8.69657e-19 $X=8.475 $Y=2.48 $X2=0 $Y2=0
cc_186 N_A_c_174_n N_VPWR_c_525_n 0.00373439f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_187 N_A_c_175_n N_VPWR_c_525_n 0.00115435f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_188 N_A_M1034_g N_VPWR_c_527_n 8.05893e-19 $X=7.945 $Y=2.48 $X2=0 $Y2=0
cc_189 N_A_c_167_n N_VPWR_c_527_n 0.00232902f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_190 N_A_M1035_g N_VPWR_c_527_n 0.0236565f $X=8.475 $Y=2.48 $X2=0 $Y2=0
cc_191 N_A_c_174_n N_VPWR_c_527_n 0.00621202f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_192 N_A_M1003_g N_VPWR_c_528_n 0.00687065f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_193 N_A_M1007_g N_VPWR_c_528_n 0.00687065f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_194 N_A_M1009_g N_VPWR_c_530_n 0.00687065f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_195 N_A_M1011_g N_VPWR_c_530_n 0.00687065f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_196 N_A_M1029_g N_VPWR_c_532_n 0.00687065f $X=6.885 $Y=2.48 $X2=0 $Y2=0
cc_197 N_A_M1030_g N_VPWR_c_532_n 0.00687065f $X=7.415 $Y=2.48 $X2=0 $Y2=0
cc_198 N_A_M1012_g N_VPWR_c_534_n 0.00687065f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_199 N_A_M1016_g N_VPWR_c_534_n 0.00687065f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_200 N_A_M1017_g N_VPWR_c_535_n 0.00687065f $X=4.765 $Y=2.48 $X2=0 $Y2=0
cc_201 N_A_M1021_g N_VPWR_c_535_n 0.00687065f $X=5.295 $Y=2.48 $X2=0 $Y2=0
cc_202 N_A_M1034_g N_VPWR_c_536_n 0.00687065f $X=7.945 $Y=2.48 $X2=0 $Y2=0
cc_203 N_A_M1035_g N_VPWR_c_536_n 0.00687065f $X=8.475 $Y=2.48 $X2=0 $Y2=0
cc_204 N_A_M1000_g N_VPWR_c_514_n 0.0129282f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_205 N_A_M1002_g N_VPWR_c_514_n 0.0129282f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_206 N_A_M1003_g N_VPWR_c_514_n 0.0129282f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_207 N_A_M1007_g N_VPWR_c_514_n 0.0129282f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_208 N_A_M1009_g N_VPWR_c_514_n 0.0129282f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_209 N_A_M1011_g N_VPWR_c_514_n 0.0129282f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_210 N_A_M1012_g N_VPWR_c_514_n 0.0129282f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_211 N_A_M1016_g N_VPWR_c_514_n 0.0129282f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_212 N_A_M1017_g N_VPWR_c_514_n 0.0129282f $X=4.765 $Y=2.48 $X2=0 $Y2=0
cc_213 N_A_M1021_g N_VPWR_c_514_n 0.0129282f $X=5.295 $Y=2.48 $X2=0 $Y2=0
cc_214 N_A_M1022_g N_VPWR_c_514_n 0.0118237f $X=5.825 $Y=2.48 $X2=0 $Y2=0
cc_215 N_A_M1023_g N_VPWR_c_514_n 0.0129282f $X=6.355 $Y=2.48 $X2=0 $Y2=0
cc_216 N_A_M1029_g N_VPWR_c_514_n 0.0129282f $X=6.885 $Y=2.48 $X2=0 $Y2=0
cc_217 N_A_M1030_g N_VPWR_c_514_n 0.0129282f $X=7.415 $Y=2.48 $X2=0 $Y2=0
cc_218 N_A_M1034_g N_VPWR_c_514_n 0.0129282f $X=7.945 $Y=2.48 $X2=0 $Y2=0
cc_219 N_A_M1035_g N_VPWR_c_514_n 0.0129282f $X=8.475 $Y=2.48 $X2=0 $Y2=0
cc_220 N_A_M1025_g N_Y_c_675_n 0.0093532f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_221 N_A_M1001_g N_Y_c_675_n 0.0168059f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_222 N_A_M1005_g N_Y_c_675_n 0.0121215f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_223 N_A_M1004_g N_Y_c_675_n 0.00127327f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_224 N_A_c_167_n N_Y_c_675_n 0.00212762f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_225 N_A_c_171_n N_Y_c_675_n 0.00314436f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_226 N_A_c_175_n N_Y_c_675_n 0.00887315f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_227 N_A_M1010_g N_Y_c_705_n 0.00294952f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_228 N_A_M1006_g N_Y_c_705_n 0.0174032f $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_229 N_A_M1008_g N_Y_c_705_n 0.0174654f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_230 N_A_M1031_g N_Y_c_705_n 0.00298431f $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_231 N_A_c_167_n N_Y_c_705_n 0.00101117f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_232 N_A_c_169_n N_Y_c_705_n 2.35614e-19 $X=3.44 $Y=1.4 $X2=0 $Y2=0
cc_233 N_A_c_171_n N_Y_c_705_n 8.7935e-19 $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_234 N_A_c_175_n N_Y_c_705_n 0.0192226f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_235 N_A_M1015_g N_Y_c_713_n 0.00296326f $X=3.635 $Y=0.61 $X2=0 $Y2=0
cc_236 N_A_M1013_g N_Y_c_713_n 0.0174089f $X=3.995 $Y=0.61 $X2=0 $Y2=0
cc_237 N_A_M1014_g N_Y_c_713_n 0.017403f $X=4.425 $Y=0.61 $X2=0 $Y2=0
cc_238 N_A_M1024_g N_Y_c_713_n 0.00302176f $X=4.785 $Y=0.61 $X2=0 $Y2=0
cc_239 N_A_c_169_n N_Y_c_713_n 3.98224e-19 $X=3.44 $Y=1.4 $X2=0 $Y2=0
cc_240 N_A_c_172_n N_Y_c_713_n 0.0172617f $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_241 N_A_c_175_n N_Y_c_713_n 0.0191522f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_242 N_A_M1019_g N_Y_c_720_n 0.00295231f $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_243 N_A_M1018_g N_Y_c_720_n 0.0174146f $X=5.575 $Y=0.61 $X2=0 $Y2=0
cc_244 N_A_M1020_g N_Y_c_720_n 0.0174594f $X=6.005 $Y=0.61 $X2=0 $Y2=0
cc_245 N_A_M1027_g N_Y_c_720_n 0.00297577f $X=6.365 $Y=0.61 $X2=0 $Y2=0
cc_246 N_A_c_167_n N_Y_c_720_n 0.00101117f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_247 N_A_c_172_n N_Y_c_720_n 7.11429e-19 $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_248 N_A_c_173_n N_Y_c_720_n 3.21263e-19 $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_249 N_A_c_175_n N_Y_c_720_n 0.0192502f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_250 N_A_M1022_g N_Y_c_683_n 0.0175603f $X=5.825 $Y=2.48 $X2=0 $Y2=0
cc_251 N_A_M1023_g N_Y_c_683_n 0.0157734f $X=6.355 $Y=2.48 $X2=0 $Y2=0
cc_252 N_A_M1026_g N_Y_c_730_n 0.00298052f $X=6.795 $Y=0.61 $X2=0 $Y2=0
cc_253 N_A_M1028_g N_Y_c_730_n 0.0174817f $X=7.155 $Y=0.61 $X2=0 $Y2=0
cc_254 N_A_M1032_g N_Y_c_730_n 0.0173911f $X=7.585 $Y=0.61 $X2=0 $Y2=0
cc_255 N_A_M1033_g N_Y_c_730_n 0.00295534f $X=7.945 $Y=0.61 $X2=0 $Y2=0
cc_256 N_A_c_167_n N_Y_c_730_n 0.00101117f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_257 N_A_c_173_n N_Y_c_730_n 2.8332e-19 $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_258 N_A_c_174_n N_Y_c_730_n 9.78674e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_259 N_A_c_175_n N_Y_c_730_n 0.0192182f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_260 N_A_M1000_g N_Y_c_684_n 0.00806477f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_261 N_A_M1002_g N_Y_c_684_n 0.00584978f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_262 N_A_M1003_g N_Y_c_684_n 0.00105163f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_263 N_A_c_175_n N_Y_c_684_n 0.0014304f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_264 N_A_M1025_g N_Y_c_676_n 0.00305574f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_265 N_A_M1000_g N_Y_c_676_n 0.00395812f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_266 N_A_M1001_g N_Y_c_676_n 0.00652913f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_267 N_A_M1002_g N_Y_c_676_n 0.00470263f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_268 N_A_M1005_g N_Y_c_676_n 0.00113655f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_269 N_A_c_167_n N_Y_c_676_n 0.0192704f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_270 N_A_c_170_n N_Y_c_676_n 0.0485825f $X=0.24 $Y=1.295 $X2=0 $Y2=0
cc_271 N_A_c_171_n N_Y_c_676_n 0.0274372f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_272 N_A_c_175_n N_Y_c_676_n 0.0347027f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_273 N_A_M1006_g N_Y_c_677_n 7.28304e-19 $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_274 N_A_M1008_g N_Y_c_677_n 0.00422479f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_275 N_A_M1031_g N_Y_c_677_n 2.30958e-19 $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_276 N_A_c_167_n N_Y_c_677_n 0.035967f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_277 N_A_c_169_n N_Y_c_677_n 0.02295f $X=3.44 $Y=1.4 $X2=0 $Y2=0
cc_278 N_A_c_171_n N_Y_c_677_n 0.0232393f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_279 N_A_c_175_n N_Y_c_677_n 0.0345224f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_280 N_A_M1011_g N_Y_c_686_n 0.00109487f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_281 N_A_M1012_g N_Y_c_686_n 0.00587694f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_282 N_A_M1016_g N_Y_c_686_n 0.00534507f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_283 N_A_M1017_g N_Y_c_686_n 3.42148e-19 $X=4.765 $Y=2.48 $X2=0 $Y2=0
cc_284 N_A_c_175_n N_Y_c_686_n 0.00204152f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_285 N_A_M1012_g N_Y_c_678_n 0.0063066f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_286 N_A_M1016_g N_Y_c_678_n 0.00689888f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_287 N_A_M1017_g N_Y_c_678_n 0.00178225f $X=4.765 $Y=2.48 $X2=0 $Y2=0
cc_288 N_A_M1013_g N_Y_c_679_n 0.0040912f $X=3.995 $Y=0.61 $X2=0 $Y2=0
cc_289 N_A_M1014_g N_Y_c_679_n 7.9939e-19 $X=4.425 $Y=0.61 $X2=0 $Y2=0
cc_290 N_A_c_167_n N_Y_c_679_n 0.0341972f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_291 N_A_c_169_n N_Y_c_679_n 0.0265534f $X=3.44 $Y=1.4 $X2=0 $Y2=0
cc_292 N_A_c_175_n N_Y_c_679_n 0.0312408f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_293 N_A_M1018_g N_Y_c_680_n 7.57281e-19 $X=5.575 $Y=0.61 $X2=0 $Y2=0
cc_294 N_A_M1020_g N_Y_c_680_n 0.00418093f $X=6.005 $Y=0.61 $X2=0 $Y2=0
cc_295 N_A_c_167_n N_Y_c_680_n 0.0344394f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_296 N_A_c_172_n N_Y_c_680_n 0.0190656f $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_297 N_A_c_173_n N_Y_c_680_n 0.0249349f $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_298 N_A_c_175_n N_Y_c_680_n 0.0320752f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_299 N_A_M1026_g N_Y_c_681_n 2.34361e-19 $X=6.795 $Y=0.61 $X2=0 $Y2=0
cc_300 N_A_M1028_g N_Y_c_681_n 0.00416495f $X=7.155 $Y=0.61 $X2=0 $Y2=0
cc_301 N_A_M1032_g N_Y_c_681_n 7.09601e-19 $X=7.585 $Y=0.61 $X2=0 $Y2=0
cc_302 N_A_c_167_n N_Y_c_681_n 0.0330736f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_303 N_A_c_173_n N_Y_c_681_n 0.0160657f $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_304 N_A_c_174_n N_Y_c_681_n 0.0272125f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_305 N_A_c_175_n N_Y_c_681_n 0.0313287f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_306 N_A_M1000_g N_Y_c_688_n 0.0201351f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_307 N_A_M1002_g N_Y_c_688_n 0.0190291f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_308 N_A_M1003_g N_Y_c_688_n 3.42738e-19 $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_309 N_A_M1002_g N_Y_c_689_n 6.00676e-19 $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_310 N_A_M1003_g N_Y_c_689_n 0.0187564f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_311 N_A_M1007_g N_Y_c_689_n 0.0187564f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_312 N_A_M1009_g N_Y_c_689_n 6.00676e-19 $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_313 N_A_c_167_n N_Y_c_689_n 5.49158e-19 $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_314 N_A_c_171_n N_Y_c_689_n 0.0101708f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_315 N_A_c_175_n N_Y_c_689_n 3.81322e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_316 N_A_M1007_g N_Y_c_690_n 0.00212374f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_317 N_A_M1009_g N_Y_c_690_n 0.029853f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_318 N_A_M1011_g N_Y_c_690_n 0.029853f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_319 N_A_M1012_g N_Y_c_690_n 0.00212374f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_320 N_A_c_167_n N_Y_c_690_n 0.00352791f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_321 N_A_c_175_n N_Y_c_690_n 5.63117e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_322 N_A_M1012_g N_Y_c_691_n 0.0167627f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_323 N_A_M1016_g N_Y_c_691_n 0.0167627f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_324 N_A_M1016_g N_Y_c_692_n 6.00676e-19 $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_325 N_A_M1017_g N_Y_c_692_n 0.0187564f $X=4.765 $Y=2.48 $X2=0 $Y2=0
cc_326 N_A_M1021_g N_Y_c_692_n 0.0187564f $X=5.295 $Y=2.48 $X2=0 $Y2=0
cc_327 N_A_M1022_g N_Y_c_692_n 6.00676e-19 $X=5.825 $Y=2.48 $X2=0 $Y2=0
cc_328 N_A_c_167_n N_Y_c_692_n 5.47993e-19 $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_329 N_A_c_172_n N_Y_c_692_n 0.0101708f $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_330 N_A_c_175_n N_Y_c_692_n 3.81322e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_331 N_A_M1023_g N_Y_c_693_n 0.00212374f $X=6.355 $Y=2.48 $X2=0 $Y2=0
cc_332 N_A_M1029_g N_Y_c_693_n 0.029853f $X=6.885 $Y=2.48 $X2=0 $Y2=0
cc_333 N_A_M1030_g N_Y_c_693_n 0.029853f $X=7.415 $Y=2.48 $X2=0 $Y2=0
cc_334 N_A_M1034_g N_Y_c_693_n 0.00212374f $X=7.945 $Y=2.48 $X2=0 $Y2=0
cc_335 N_A_c_167_n N_Y_c_693_n 0.00352791f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_336 N_A_c_175_n N_Y_c_693_n 5.63117e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_337 N_A_M1030_g N_Y_c_694_n 6.00676e-19 $X=7.415 $Y=2.48 $X2=0 $Y2=0
cc_338 N_A_M1034_g N_Y_c_694_n 0.0187571f $X=7.945 $Y=2.48 $X2=0 $Y2=0
cc_339 N_A_c_167_n N_Y_c_694_n 0.00191254f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_340 N_A_M1035_g N_Y_c_694_n 0.0216295f $X=8.475 $Y=2.48 $X2=0 $Y2=0
cc_341 N_A_c_174_n N_Y_c_694_n 0.0103398f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_342 N_A_c_175_n N_Y_c_694_n 4.40983e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_343 N_A_M1000_g N_Y_c_695_n 0.00625372f $X=0.525 $Y=2.48 $X2=0 $Y2=0
cc_344 N_A_M1002_g N_Y_c_695_n 0.0120234f $X=1.055 $Y=2.48 $X2=0 $Y2=0
cc_345 N_A_M1003_g N_Y_c_695_n 0.0115941f $X=1.585 $Y=2.48 $X2=0 $Y2=0
cc_346 N_A_M1007_g N_Y_c_695_n 0.0115941f $X=2.115 $Y=2.48 $X2=0 $Y2=0
cc_347 N_A_M1009_g N_Y_c_695_n 0.0113428f $X=2.645 $Y=2.48 $X2=0 $Y2=0
cc_348 N_A_M1011_g N_Y_c_695_n 0.0124655f $X=3.175 $Y=2.48 $X2=0 $Y2=0
cc_349 N_A_M1012_g N_Y_c_695_n 0.011879f $X=3.705 $Y=2.48 $X2=0 $Y2=0
cc_350 N_A_M1016_g N_Y_c_695_n 0.0113303f $X=4.235 $Y=2.48 $X2=0 $Y2=0
cc_351 N_A_M1017_g N_Y_c_695_n 0.0116836f $X=4.765 $Y=2.48 $X2=0 $Y2=0
cc_352 N_A_M1021_g N_Y_c_695_n 0.0118235f $X=5.295 $Y=2.48 $X2=0 $Y2=0
cc_353 N_A_M1022_g N_Y_c_695_n 0.00971468f $X=5.825 $Y=2.48 $X2=0 $Y2=0
cc_354 N_A_M1023_g N_Y_c_695_n 0.0119954f $X=6.355 $Y=2.48 $X2=0 $Y2=0
cc_355 N_A_M1029_g N_Y_c_695_n 0.0126052f $X=6.885 $Y=2.48 $X2=0 $Y2=0
cc_356 N_A_M1030_g N_Y_c_695_n 0.0113707f $X=7.415 $Y=2.48 $X2=0 $Y2=0
cc_357 N_A_M1034_g N_Y_c_695_n 0.0115963f $X=7.945 $Y=2.48 $X2=0 $Y2=0
cc_358 N_A_c_167_n N_Y_c_695_n 0.00910449f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_359 N_A_c_169_n N_Y_c_695_n 0.00583575f $X=3.44 $Y=1.4 $X2=0 $Y2=0
cc_360 N_A_c_171_n N_Y_c_695_n 0.0167964f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_361 N_A_c_172_n N_Y_c_695_n 0.010794f $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_362 N_A_c_173_n N_Y_c_695_n 0.00447841f $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_363 N_A_c_174_n N_Y_c_695_n 0.00764294f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_364 N_A_c_175_n N_Y_c_695_n 0.362232f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_365 N_A_M1021_g N_Y_c_696_n 3.19008e-19 $X=5.295 $Y=2.48 $X2=0 $Y2=0
cc_366 N_A_M1022_g N_Y_c_696_n 0.00447619f $X=5.825 $Y=2.48 $X2=0 $Y2=0
cc_367 N_A_M1023_g N_Y_c_696_n 0.00474094f $X=6.355 $Y=2.48 $X2=0 $Y2=0
cc_368 N_A_M1029_g N_Y_c_696_n 7.9557e-19 $X=6.885 $Y=2.48 $X2=0 $Y2=0
cc_369 N_A_c_175_n N_Y_c_696_n 0.00162193f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_370 N_A_M1021_g N_Y_c_682_n 0.00187871f $X=5.295 $Y=2.48 $X2=0 $Y2=0
cc_371 N_A_M1022_g N_Y_c_682_n 0.00976352f $X=5.825 $Y=2.48 $X2=0 $Y2=0
cc_372 N_A_M1023_g N_Y_c_682_n 0.008518f $X=6.355 $Y=2.48 $X2=0 $Y2=0
cc_373 N_A_c_167_n N_Y_c_682_n 0.00341969f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_374 N_A_c_175_n N_Y_c_682_n 5.03028e-19 $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_375 N_A_M1025_g N_VGND_c_920_n 0.0121638f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_376 N_A_M1001_g N_VGND_c_920_n 0.00106741f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_377 N_A_c_167_n N_VGND_c_920_n 0.00118321f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_378 N_A_c_170_n N_VGND_c_920_n 0.0145155f $X=0.24 $Y=1.295 $X2=0 $Y2=0
cc_379 N_A_c_175_n N_VGND_c_920_n 0.00251493f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_380 N_A_M1005_g N_VGND_c_921_n 0.00194004f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_381 N_A_M1004_g N_VGND_c_921_n 0.0129138f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_382 N_A_M1010_g N_VGND_c_921_n 0.0131f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_383 N_A_M1006_g N_VGND_c_921_n 0.00223895f $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_384 N_A_c_167_n N_VGND_c_921_n 6.36823e-19 $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_385 N_A_c_171_n N_VGND_c_921_n 0.00780499f $X=1.2 $Y=1.295 $X2=0 $Y2=0
cc_386 N_A_c_175_n N_VGND_c_921_n 0.00259541f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_387 N_A_M1008_g N_VGND_c_922_n 0.00223895f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_388 N_A_M1031_g N_VGND_c_922_n 0.0130244f $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_389 N_A_M1015_g N_VGND_c_922_n 0.0131007f $X=3.635 $Y=0.61 $X2=0 $Y2=0
cc_390 N_A_M1013_g N_VGND_c_922_n 0.00223895f $X=3.995 $Y=0.61 $X2=0 $Y2=0
cc_391 N_A_c_167_n N_VGND_c_922_n 6.37201e-19 $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_392 N_A_c_169_n N_VGND_c_922_n 0.00731964f $X=3.44 $Y=1.4 $X2=0 $Y2=0
cc_393 N_A_c_175_n N_VGND_c_922_n 0.0082865f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_394 N_A_M1014_g N_VGND_c_923_n 0.00223895f $X=4.425 $Y=0.61 $X2=0 $Y2=0
cc_395 N_A_M1024_g N_VGND_c_923_n 0.0131f $X=4.785 $Y=0.61 $X2=0 $Y2=0
cc_396 N_A_M1019_g N_VGND_c_923_n 0.0131f $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_397 N_A_M1018_g N_VGND_c_923_n 0.00223895f $X=5.575 $Y=0.61 $X2=0 $Y2=0
cc_398 N_A_c_167_n N_VGND_c_923_n 6.35875e-19 $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_399 N_A_c_172_n N_VGND_c_923_n 0.00780499f $X=5.04 $Y=1.295 $X2=0 $Y2=0
cc_400 N_A_c_175_n N_VGND_c_923_n 0.00259541f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_401 N_A_M1020_g N_VGND_c_924_n 0.00223895f $X=6.005 $Y=0.61 $X2=0 $Y2=0
cc_402 N_A_M1027_g N_VGND_c_924_n 0.0131f $X=6.365 $Y=0.61 $X2=0 $Y2=0
cc_403 N_A_M1026_g N_VGND_c_924_n 0.0131187f $X=6.795 $Y=0.61 $X2=0 $Y2=0
cc_404 N_A_M1028_g N_VGND_c_924_n 0.00223895f $X=7.155 $Y=0.61 $X2=0 $Y2=0
cc_405 N_A_c_167_n N_VGND_c_924_n 6.354e-19 $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_406 N_A_c_173_n N_VGND_c_924_n 0.00691915f $X=6.48 $Y=1.295 $X2=0 $Y2=0
cc_407 N_A_c_175_n N_VGND_c_924_n 0.0040015f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_408 N_A_M1032_g N_VGND_c_925_n 0.00223895f $X=7.585 $Y=0.61 $X2=0 $Y2=0
cc_409 N_A_M1033_g N_VGND_c_925_n 0.0148319f $X=7.945 $Y=0.61 $X2=0 $Y2=0
cc_410 N_A_c_167_n N_VGND_c_925_n 0.00170633f $X=8.475 $Y=1.565 $X2=0 $Y2=0
cc_411 N_A_c_174_n N_VGND_c_925_n 0.00881269f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_412 N_A_c_175_n N_VGND_c_925_n 0.00811184f $X=8.4 $Y=1.295 $X2=0 $Y2=0
cc_413 N_A_M1010_g N_VGND_c_926_n 0.00407525f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_414 N_A_M1006_g N_VGND_c_926_n 0.00464284f $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_415 N_A_M1008_g N_VGND_c_926_n 0.00464284f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_416 N_A_M1031_g N_VGND_c_926_n 0.00407525f $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_417 N_A_M1026_g N_VGND_c_928_n 0.00407525f $X=6.795 $Y=0.61 $X2=0 $Y2=0
cc_418 N_A_M1028_g N_VGND_c_928_n 0.00464284f $X=7.155 $Y=0.61 $X2=0 $Y2=0
cc_419 N_A_M1032_g N_VGND_c_928_n 0.00464284f $X=7.585 $Y=0.61 $X2=0 $Y2=0
cc_420 N_A_M1033_g N_VGND_c_928_n 0.00407525f $X=7.945 $Y=0.61 $X2=0 $Y2=0
cc_421 N_A_M1025_g N_VGND_c_930_n 0.00407525f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_422 N_A_M1001_g N_VGND_c_930_n 0.00306164f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_423 N_A_M1005_g N_VGND_c_930_n 0.00460042f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_424 N_A_M1004_g N_VGND_c_930_n 0.00407525f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_425 N_A_M1015_g N_VGND_c_931_n 0.00407525f $X=3.635 $Y=0.61 $X2=0 $Y2=0
cc_426 N_A_M1013_g N_VGND_c_931_n 0.00464284f $X=3.995 $Y=0.61 $X2=0 $Y2=0
cc_427 N_A_M1014_g N_VGND_c_931_n 0.00464284f $X=4.425 $Y=0.61 $X2=0 $Y2=0
cc_428 N_A_M1024_g N_VGND_c_931_n 0.00407525f $X=4.785 $Y=0.61 $X2=0 $Y2=0
cc_429 N_A_M1019_g N_VGND_c_932_n 0.00407525f $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_430 N_A_M1018_g N_VGND_c_932_n 0.00464284f $X=5.575 $Y=0.61 $X2=0 $Y2=0
cc_431 N_A_M1020_g N_VGND_c_932_n 0.00464284f $X=6.005 $Y=0.61 $X2=0 $Y2=0
cc_432 N_A_M1027_g N_VGND_c_932_n 0.00407525f $X=6.365 $Y=0.61 $X2=0 $Y2=0
cc_433 N_A_M1025_g N_VGND_c_934_n 0.00774993f $X=0.475 $Y=0.61 $X2=0 $Y2=0
cc_434 N_A_M1001_g N_VGND_c_934_n 0.0041313f $X=0.835 $Y=0.61 $X2=0 $Y2=0
cc_435 N_A_M1005_g N_VGND_c_934_n 0.00874299f $X=1.265 $Y=0.61 $X2=0 $Y2=0
cc_436 N_A_M1004_g N_VGND_c_934_n 0.00774993f $X=1.625 $Y=0.61 $X2=0 $Y2=0
cc_437 N_A_M1010_g N_VGND_c_934_n 0.00774993f $X=2.055 $Y=0.61 $X2=0 $Y2=0
cc_438 N_A_M1006_g N_VGND_c_934_n 0.0088065f $X=2.415 $Y=0.61 $X2=0 $Y2=0
cc_439 N_A_M1008_g N_VGND_c_934_n 0.0088065f $X=2.845 $Y=0.61 $X2=0 $Y2=0
cc_440 N_A_M1031_g N_VGND_c_934_n 0.00774993f $X=3.205 $Y=0.61 $X2=0 $Y2=0
cc_441 N_A_M1015_g N_VGND_c_934_n 0.00774993f $X=3.635 $Y=0.61 $X2=0 $Y2=0
cc_442 N_A_M1013_g N_VGND_c_934_n 0.0088065f $X=3.995 $Y=0.61 $X2=0 $Y2=0
cc_443 N_A_M1014_g N_VGND_c_934_n 0.0088065f $X=4.425 $Y=0.61 $X2=0 $Y2=0
cc_444 N_A_M1024_g N_VGND_c_934_n 0.00774993f $X=4.785 $Y=0.61 $X2=0 $Y2=0
cc_445 N_A_M1019_g N_VGND_c_934_n 0.00774993f $X=5.215 $Y=0.61 $X2=0 $Y2=0
cc_446 N_A_M1018_g N_VGND_c_934_n 0.0088065f $X=5.575 $Y=0.61 $X2=0 $Y2=0
cc_447 N_A_M1020_g N_VGND_c_934_n 0.0088065f $X=6.005 $Y=0.61 $X2=0 $Y2=0
cc_448 N_A_M1027_g N_VGND_c_934_n 0.00774993f $X=6.365 $Y=0.61 $X2=0 $Y2=0
cc_449 N_A_M1026_g N_VGND_c_934_n 0.00774993f $X=6.795 $Y=0.61 $X2=0 $Y2=0
cc_450 N_A_M1028_g N_VGND_c_934_n 0.0088065f $X=7.155 $Y=0.61 $X2=0 $Y2=0
cc_451 N_A_M1032_g N_VGND_c_934_n 0.0088065f $X=7.585 $Y=0.61 $X2=0 $Y2=0
cc_452 N_A_M1033_g N_VGND_c_934_n 0.00774993f $X=7.945 $Y=0.61 $X2=0 $Y2=0
cc_453 N_VPWR_c_523_n N_Y_c_683_n 0.0171239f $X=6.455 $Y=3.33 $X2=0 $Y2=0
cc_454 N_VPWR_c_514_n N_Y_c_683_n 0.0130063f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_455 N_VPWR_c_519_n N_Y_c_677_n 0.00207514f $X=2.38 $Y=2.125 $X2=0 $Y2=0
cc_456 N_VPWR_c_520_n N_Y_c_686_n 0.0663323f $X=3.44 $Y=2.125 $X2=0 $Y2=0
cc_457 N_VPWR_c_521_n N_Y_c_686_n 0.0663323f $X=4.5 $Y=2.125 $X2=0 $Y2=0
cc_458 N_VPWR_c_521_n N_Y_c_679_n 9.95116e-19 $X=4.5 $Y=2.125 $X2=0 $Y2=0
cc_459 N_VPWR_c_522_n N_Y_c_680_n 0.00262489f $X=5.56 $Y=2.125 $X2=0 $Y2=0
cc_460 N_VPWR_c_525_n N_Y_c_681_n 4.45963e-19 $X=7.68 $Y=2.125 $X2=0 $Y2=0
cc_461 N_VPWR_c_516_n N_Y_c_688_n 0.0658767f $X=0.26 $Y=2.125 $X2=0 $Y2=0
cc_462 N_VPWR_c_517_n N_Y_c_688_n 0.0157615f $X=1.155 $Y=3.33 $X2=0 $Y2=0
cc_463 N_VPWR_c_518_n N_Y_c_688_n 0.0663595f $X=1.32 $Y=2.125 $X2=0 $Y2=0
cc_464 N_VPWR_c_514_n N_Y_c_688_n 0.0120285f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_465 N_VPWR_c_518_n N_Y_c_689_n 0.0663595f $X=1.32 $Y=2.125 $X2=0 $Y2=0
cc_466 N_VPWR_c_519_n N_Y_c_689_n 0.0663595f $X=2.38 $Y=2.125 $X2=0 $Y2=0
cc_467 N_VPWR_c_528_n N_Y_c_689_n 0.0157615f $X=2.215 $Y=3.33 $X2=0 $Y2=0
cc_468 N_VPWR_c_514_n N_Y_c_689_n 0.0120285f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_469 N_VPWR_c_519_n N_Y_c_690_n 0.0663595f $X=2.38 $Y=2.125 $X2=0 $Y2=0
cc_470 N_VPWR_c_520_n N_Y_c_690_n 0.0663595f $X=3.44 $Y=2.125 $X2=0 $Y2=0
cc_471 N_VPWR_c_530_n N_Y_c_690_n 0.0157615f $X=3.275 $Y=3.33 $X2=0 $Y2=0
cc_472 N_VPWR_c_514_n N_Y_c_690_n 0.0120285f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_473 N_VPWR_c_534_n N_Y_c_691_n 0.0157615f $X=4.335 $Y=3.33 $X2=0 $Y2=0
cc_474 N_VPWR_c_514_n N_Y_c_691_n 0.0120285f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_475 N_VPWR_c_521_n N_Y_c_692_n 0.0663595f $X=4.5 $Y=2.125 $X2=0 $Y2=0
cc_476 N_VPWR_c_522_n N_Y_c_692_n 0.0663595f $X=5.56 $Y=2.125 $X2=0 $Y2=0
cc_477 N_VPWR_c_535_n N_Y_c_692_n 0.0157615f $X=5.395 $Y=3.33 $X2=0 $Y2=0
cc_478 N_VPWR_c_514_n N_Y_c_692_n 0.0120285f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_479 N_VPWR_c_524_n N_Y_c_693_n 0.0663595f $X=6.62 $Y=2.125 $X2=0 $Y2=0
cc_480 N_VPWR_c_525_n N_Y_c_693_n 0.0663595f $X=7.68 $Y=2.125 $X2=0 $Y2=0
cc_481 N_VPWR_c_532_n N_Y_c_693_n 0.0157615f $X=7.515 $Y=3.33 $X2=0 $Y2=0
cc_482 N_VPWR_c_514_n N_Y_c_693_n 0.0120285f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_483 N_VPWR_c_525_n N_Y_c_694_n 0.0663595f $X=7.68 $Y=2.125 $X2=0 $Y2=0
cc_484 N_VPWR_c_527_n N_Y_c_694_n 0.0671438f $X=8.74 $Y=2.125 $X2=0 $Y2=0
cc_485 N_VPWR_c_536_n N_Y_c_694_n 0.0157615f $X=8.575 $Y=3.33 $X2=0 $Y2=0
cc_486 N_VPWR_c_514_n N_Y_c_694_n 0.0120285f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_487 N_VPWR_c_516_n N_Y_c_695_n 0.00575829f $X=0.26 $Y=2.125 $X2=0 $Y2=0
cc_488 N_VPWR_c_518_n N_Y_c_695_n 0.0320279f $X=1.32 $Y=2.125 $X2=0 $Y2=0
cc_489 N_VPWR_c_519_n N_Y_c_695_n 0.0344002f $X=2.38 $Y=2.125 $X2=0 $Y2=0
cc_490 N_VPWR_c_520_n N_Y_c_695_n 0.0320347f $X=3.44 $Y=2.125 $X2=0 $Y2=0
cc_491 N_VPWR_c_521_n N_Y_c_695_n 0.0352693f $X=4.5 $Y=2.125 $X2=0 $Y2=0
cc_492 N_VPWR_c_522_n N_Y_c_695_n 0.034316f $X=5.56 $Y=2.125 $X2=0 $Y2=0
cc_493 N_VPWR_c_524_n N_Y_c_695_n 0.0329035f $X=6.62 $Y=2.125 $X2=0 $Y2=0
cc_494 N_VPWR_c_525_n N_Y_c_695_n 0.0340098f $X=7.68 $Y=2.125 $X2=0 $Y2=0
cc_495 N_VPWR_c_527_n N_Y_c_695_n 0.00126886f $X=8.74 $Y=2.125 $X2=0 $Y2=0
cc_496 N_VPWR_c_522_n N_Y_c_696_n 0.0765853f $X=5.56 $Y=2.125 $X2=0 $Y2=0
cc_497 N_VPWR_c_524_n N_Y_c_696_n 0.0667114f $X=6.62 $Y=2.125 $X2=0 $Y2=0
cc_498 N_Y_c_675_n N_VGND_c_920_n 0.0331575f $X=0.765 $Y=1.01 $X2=0 $Y2=0
cc_499 N_Y_c_675_n N_VGND_c_921_n 0.0161396f $X=0.765 $Y=1.01 $X2=0 $Y2=0
cc_500 N_Y_c_705_n N_VGND_c_921_n 0.0110409f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_501 N_Y_c_705_n N_VGND_c_922_n 0.0110409f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_502 N_Y_c_713_n N_VGND_c_922_n 0.0110409f $X=4.21 $Y=0.61 $X2=0 $Y2=0
cc_503 N_Y_c_713_n N_VGND_c_923_n 0.0110409f $X=4.21 $Y=0.61 $X2=0 $Y2=0
cc_504 N_Y_c_720_n N_VGND_c_923_n 0.0110409f $X=5.79 $Y=0.61 $X2=0 $Y2=0
cc_505 N_Y_c_720_n N_VGND_c_924_n 0.0110409f $X=5.79 $Y=0.61 $X2=0 $Y2=0
cc_506 N_Y_c_730_n N_VGND_c_924_n 0.0110409f $X=7.37 $Y=0.61 $X2=0 $Y2=0
cc_507 N_Y_c_730_n N_VGND_c_925_n 0.0110409f $X=7.37 $Y=0.61 $X2=0 $Y2=0
cc_508 N_Y_c_705_n N_VGND_c_926_n 0.00846545f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_509 N_Y_c_730_n N_VGND_c_928_n 0.00846545f $X=7.37 $Y=0.61 $X2=0 $Y2=0
cc_510 N_Y_c_675_n N_VGND_c_930_n 0.0296946f $X=0.765 $Y=1.01 $X2=0 $Y2=0
cc_511 N_Y_c_713_n N_VGND_c_931_n 0.00846545f $X=4.21 $Y=0.61 $X2=0 $Y2=0
cc_512 N_Y_c_720_n N_VGND_c_932_n 0.00846545f $X=5.79 $Y=0.61 $X2=0 $Y2=0
cc_513 N_Y_c_675_n N_VGND_c_934_n 0.0212961f $X=0.765 $Y=1.01 $X2=0 $Y2=0
cc_514 N_Y_c_705_n N_VGND_c_934_n 0.0111318f $X=2.63 $Y=0.61 $X2=0 $Y2=0
cc_515 N_Y_c_713_n N_VGND_c_934_n 0.0111318f $X=4.21 $Y=0.61 $X2=0 $Y2=0
cc_516 N_Y_c_720_n N_VGND_c_934_n 0.0111318f $X=5.79 $Y=0.61 $X2=0 $Y2=0
cc_517 N_Y_c_730_n N_VGND_c_934_n 0.0111318f $X=7.37 $Y=0.61 $X2=0 $Y2=0
cc_518 N_Y_c_675_n A_268_67# 0.00528527f $X=0.765 $Y=1.01 $X2=-0.19 $Y2=-0.245
