* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2_4 A0 A1 S VGND VNB VPB VPWR X
X0 X a_359_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_287_47# A0 a_359_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 X a_359_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VPWR a_359_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 X a_359_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_359_47# A1 a_508_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_359_47# A1 a_210_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_317_367# A0 a_359_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND a_359_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 X a_359_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR a_359_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_41_367# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VGND a_41_367# a_287_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VPWR a_41_367# a_210_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_508_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_41_367# S VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VGND a_359_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_317_367# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
