* File: sky130_fd_sc_lp__o22a_m.pxi.spice
* Created: Wed Sep  2 10:20:19 2020
* 
x_PM_SKY130_FD_SC_LP__O22A_M%A_88_187# N_A_88_187#_M1008_d N_A_88_187#_M1001_d
+ N_A_88_187#_c_62_n N_A_88_187#_M1000_g N_A_88_187#_M1002_g N_A_88_187#_c_64_n
+ N_A_88_187#_c_65_n N_A_88_187#_c_66_n N_A_88_187#_c_67_n N_A_88_187#_c_108_p
+ N_A_88_187#_c_72_n N_A_88_187#_c_109_p N_A_88_187#_c_102_p N_A_88_187#_c_68_n
+ N_A_88_187#_c_69_n PM_SKY130_FD_SC_LP__O22A_M%A_88_187#
x_PM_SKY130_FD_SC_LP__O22A_M%A1 N_A1_M1007_g N_A1_M1005_g N_A1_c_148_n
+ N_A1_c_143_n N_A1_c_160_n N_A1_c_144_n A1 A1 A1 N_A1_c_146_n
+ PM_SKY130_FD_SC_LP__O22A_M%A1
x_PM_SKY130_FD_SC_LP__O22A_M%B1 N_B1_M1008_g N_B1_M1004_g N_B1_c_202_n
+ N_B1_c_203_n B1 PM_SKY130_FD_SC_LP__O22A_M%B1
x_PM_SKY130_FD_SC_LP__O22A_M%B2 N_B2_M1001_g N_B2_M1009_g N_B2_c_240_n
+ N_B2_c_241_n B2 B2 N_B2_c_243_n PM_SKY130_FD_SC_LP__O22A_M%B2
x_PM_SKY130_FD_SC_LP__O22A_M%A2 N_A2_c_271_n N_A2_M1006_g N_A2_c_273_n
+ N_A2_M1003_g A2 A2 PM_SKY130_FD_SC_LP__O22A_M%A2
x_PM_SKY130_FD_SC_LP__O22A_M%X N_X_M1002_s N_X_M1000_s N_X_c_305_n X X X X X X
+ PM_SKY130_FD_SC_LP__O22A_M%X
x_PM_SKY130_FD_SC_LP__O22A_M%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_c_321_n
+ N_VPWR_c_322_n N_VPWR_c_323_n VPWR N_VPWR_c_324_n N_VPWR_c_325_n
+ N_VPWR_c_326_n N_VPWR_c_320_n PM_SKY130_FD_SC_LP__O22A_M%VPWR
x_PM_SKY130_FD_SC_LP__O22A_M%VGND N_VGND_M1002_d N_VGND_M1003_d N_VGND_c_366_n
+ N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n VGND N_VGND_c_370_n
+ N_VGND_c_371_n N_VGND_c_372_n PM_SKY130_FD_SC_LP__O22A_M%VGND
x_PM_SKY130_FD_SC_LP__O22A_M%A_237_81# N_A_237_81#_M1007_d N_A_237_81#_M1009_d
+ N_A_237_81#_c_404_n N_A_237_81#_c_405_n N_A_237_81#_c_406_n
+ PM_SKY130_FD_SC_LP__O22A_M%A_237_81#
cc_1 VNB N_A_88_187#_c_62_n 0.0243924f $X=-0.19 $Y=-0.245 $X2=0.617 $Y2=1.428
cc_2 VNB N_A_88_187#_M1000_g 0.00271133f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.885
cc_3 VNB N_A_88_187#_c_64_n 0.0217295f $X=-0.19 $Y=-0.245 $X2=0.617 $Y2=1.605
cc_4 VNB N_A_88_187#_c_65_n 3.82471e-19 $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.1
cc_5 VNB N_A_88_187#_c_66_n 0.0194671f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.1
cc_6 VNB N_A_88_187#_c_67_n 0.0113455f $X=-0.19 $Y=-0.245 $X2=1.67 $Y2=0.9
cc_7 VNB N_A_88_187#_c_68_n 0.00416461f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.7
cc_8 VNB N_A_88_187#_c_69_n 0.0212298f $X=-0.19 $Y=-0.245 $X2=0.617 $Y2=0.935
cc_9 VNB N_A1_M1007_g 0.0243998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_143_n 0.0206075f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.935
cc_11 VNB N_A1_c_144_n 0.0427712f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.985
cc_12 VNB A1 0.0103173f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.1
cc_13 VNB N_A1_c_146_n 0.00927694f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.7
cc_14 VNB N_B1_M1008_g 0.050519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_M1009_g 0.0542335f $X=-0.19 $Y=-0.245 $X2=0.617 $Y2=1.112
cc_16 VNB N_A2_c_271_n 0.0567238f $X=-0.19 $Y=-0.245 $X2=1.695 $Y2=0.405
cc_17 VNB N_A2_M1006_g 0.0136406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_273_n 0.0179825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB A2 0.0320046f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.605
cc_20 VNB N_X_c_305_n 0.00774695f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.605
cc_21 VNB X 0.0482802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_320_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.617 $Y2=1.1
cc_23 VNB N_VGND_c_366_n 0.0119452f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.885
cc_24 VNB N_VGND_c_367_n 0.0255801f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.615
cc_25 VNB N_VGND_c_368_n 0.0419211f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.535
cc_26 VNB N_VGND_c_369_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.1
cc_27 VNB N_VGND_c_370_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.7
cc_28 VNB N_VGND_c_371_n 0.216579f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.7
cc_29 VNB N_VGND_c_372_n 0.0269996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_237_81#_c_404_n 0.00558527f $X=-0.19 $Y=-0.245 $X2=0.617 $Y2=1.112
cc_31 VNB N_A_237_81#_c_405_n 0.00276651f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.605
cc_32 VNB N_A_237_81#_c_406_n 0.00276869f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.615
cc_33 VPB N_A_88_187#_M1000_g 0.0780017f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.885
cc_34 VPB N_A_88_187#_c_65_n 0.01837f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.1
cc_35 VPB N_A_88_187#_c_72_n 0.0256231f $X=-0.19 $Y=1.655 $X2=2.09 $Y2=2.62
cc_36 VPB N_A1_M1005_g 0.0367794f $X=-0.19 $Y=1.655 $X2=0.617 $Y2=1.112
cc_37 VPB N_A1_c_148_n 0.0183924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A1_c_143_n 0.0195181f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.935
cc_39 VPB N_A1_c_144_n 0.0146535f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.985
cc_40 VPB A1 0.0339357f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.1
cc_41 VPB N_A1_c_146_n 0.0496787f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=0.7
cc_42 VPB N_B1_M1008_g 0.0220897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_B1_M1004_g 0.0370254f $X=-0.19 $Y=1.655 $X2=0.617 $Y2=1.112
cc_44 VPB N_B1_c_202_n 0.0494443f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.605
cc_45 VPB N_B1_c_203_n 0.00860416f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.885
cc_46 VPB B1 0.00368569f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.885
cc_47 VPB N_B2_M1001_g 0.0224199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_B2_M1009_g 0.00597243f $X=-0.19 $Y=1.655 $X2=0.617 $Y2=1.112
cc_49 VPB N_B2_c_240_n 0.0187158f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.885
cc_50 VPB N_B2_c_241_n 0.0147324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB B2 0.00937551f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.615
cc_52 VPB N_B2_c_243_n 0.0147337f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.535
cc_53 VPB N_A2_M1006_g 0.0622595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB X 0.0620435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_321_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.605
cc_56 VPB N_VPWR_c_322_n 0.0104933f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.885
cc_57 VPB N_VPWR_c_323_n 0.0138343f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.935
cc_58 VPB N_VPWR_c_324_n 0.0172304f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.985
cc_59 VPB N_VPWR_c_325_n 0.0565823f $X=-0.19 $Y=1.655 $X2=1.67 $Y2=0.9
cc_60 VPB N_VPWR_c_326_n 0.00510002f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=0.7
cc_61 VPB N_VPWR_c_320_n 0.0464872f $X=-0.19 $Y=1.655 $X2=0.617 $Y2=1.1
cc_62 N_A_88_187#_c_65_n N_A1_M1007_g 5.4276e-19 $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_63 N_A_88_187#_c_66_n N_A1_M1007_g 0.00842562f $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_64 N_A_88_187#_c_67_n N_A1_M1007_g 0.0124073f $X=1.67 $Y=0.9 $X2=0 $Y2=0
cc_65 N_A_88_187#_c_68_n N_A1_M1007_g 7.169e-19 $X=1.835 $Y=0.7 $X2=0 $Y2=0
cc_66 N_A_88_187#_c_69_n N_A1_M1007_g 0.0154677f $X=0.617 $Y=0.935 $X2=0 $Y2=0
cc_67 N_A_88_187#_c_67_n N_A1_c_143_n 0.0108479f $X=1.67 $Y=0.9 $X2=0 $Y2=0
cc_68 N_A_88_187#_c_68_n N_A1_c_143_n 0.0119066f $X=1.835 $Y=0.7 $X2=0 $Y2=0
cc_69 N_A_88_187#_c_62_n N_A1_c_160_n 0.0016442f $X=0.617 $Y=1.428 $X2=0 $Y2=0
cc_70 N_A_88_187#_c_65_n N_A1_c_160_n 0.0239869f $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_71 N_A_88_187#_c_67_n N_A1_c_160_n 0.0239644f $X=1.67 $Y=0.9 $X2=0 $Y2=0
cc_72 N_A_88_187#_c_62_n N_A1_c_144_n 0.0163862f $X=0.617 $Y=1.428 $X2=0 $Y2=0
cc_73 N_A_88_187#_M1000_g N_A1_c_144_n 0.00378059f $X=0.515 $Y=2.885 $X2=0 $Y2=0
cc_74 N_A_88_187#_c_65_n N_A1_c_144_n 0.0039306f $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_75 N_A_88_187#_c_66_n N_A1_c_144_n 0.0163862f $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_76 N_A_88_187#_c_67_n N_A1_c_144_n 0.00512673f $X=1.67 $Y=0.9 $X2=0 $Y2=0
cc_77 N_A_88_187#_c_67_n N_B1_M1008_g 0.0106242f $X=1.67 $Y=0.9 $X2=0 $Y2=0
cc_78 N_A_88_187#_c_68_n N_B1_M1008_g 0.00743101f $X=1.835 $Y=0.7 $X2=0 $Y2=0
cc_79 N_A_88_187#_c_72_n N_B1_M1004_g 0.0149306f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_80 N_A_88_187#_M1000_g N_B1_c_202_n 0.00797014f $X=0.515 $Y=2.885 $X2=0 $Y2=0
cc_81 N_A_88_187#_c_65_n N_B1_c_202_n 0.00292769f $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_82 N_A_88_187#_c_72_n N_B1_c_202_n 0.0134188f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_83 N_A_88_187#_M1000_g B1 5.34131e-19 $X=0.515 $Y=2.885 $X2=0 $Y2=0
cc_84 N_A_88_187#_c_65_n B1 0.014357f $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_85 N_A_88_187#_c_72_n B1 0.0109236f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_86 N_A_88_187#_c_72_n N_B2_M1001_g 0.0109749f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_87 N_A_88_187#_c_68_n N_B2_M1009_g 0.00929658f $X=1.835 $Y=0.7 $X2=0 $Y2=0
cc_88 N_A_88_187#_c_72_n N_B2_c_241_n 0.00522449f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_89 N_A_88_187#_c_72_n B2 0.0493359f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_90 N_A_88_187#_c_72_n N_A2_M1006_g 0.00502338f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_91 N_A_88_187#_c_102_p N_A2_M1006_g 0.00495675f $X=2.195 $Y=2.82 $X2=0 $Y2=0
cc_92 N_A_88_187#_c_68_n N_A2_c_273_n 8.13518e-19 $X=1.835 $Y=0.7 $X2=0 $Y2=0
cc_93 N_A_88_187#_c_68_n A2 0.00488669f $X=1.835 $Y=0.7 $X2=0 $Y2=0
cc_94 N_A_88_187#_c_69_n N_X_c_305_n 0.00174322f $X=0.617 $Y=0.935 $X2=0 $Y2=0
cc_95 N_A_88_187#_c_65_n X 0.108463f $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_96 N_A_88_187#_c_66_n X 0.0445856f $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_97 N_A_88_187#_c_108_p X 0.01322f $X=0.715 $Y=0.9 $X2=0 $Y2=0
cc_98 N_A_88_187#_c_109_p X 0.0132317f $X=0.715 $Y=2.62 $X2=0 $Y2=0
cc_99 N_A_88_187#_c_69_n X 0.00735798f $X=0.617 $Y=0.935 $X2=0 $Y2=0
cc_100 N_A_88_187#_c_72_n N_VPWR_M1000_d 0.0130176f $X=2.09 $Y=2.62 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_88_187#_c_109_p N_VPWR_M1000_d 7.38663e-19 $X=0.715 $Y=2.62 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_88_187#_M1000_g N_VPWR_c_321_n 0.0118722f $X=0.515 $Y=2.885 $X2=0
+ $Y2=0
cc_103 N_A_88_187#_c_72_n N_VPWR_c_321_n 0.0128944f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_104 N_A_88_187#_c_109_p N_VPWR_c_321_n 0.00716712f $X=0.715 $Y=2.62 $X2=0
+ $Y2=0
cc_105 N_A_88_187#_c_102_p N_VPWR_c_323_n 0.00371471f $X=2.195 $Y=2.82 $X2=0
+ $Y2=0
cc_106 N_A_88_187#_M1000_g N_VPWR_c_324_n 0.00465533f $X=0.515 $Y=2.885 $X2=0
+ $Y2=0
cc_107 N_A_88_187#_c_109_p N_VPWR_c_324_n 3.4848e-19 $X=0.715 $Y=2.62 $X2=0
+ $Y2=0
cc_108 N_A_88_187#_c_72_n N_VPWR_c_325_n 0.0193717f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_109 N_A_88_187#_c_102_p N_VPWR_c_325_n 0.00854632f $X=2.195 $Y=2.82 $X2=0
+ $Y2=0
cc_110 N_A_88_187#_M1001_d N_VPWR_c_320_n 0.00840059f $X=2.055 $Y=2.675 $X2=0
+ $Y2=0
cc_111 N_A_88_187#_M1000_g N_VPWR_c_320_n 0.0087003f $X=0.515 $Y=2.885 $X2=0
+ $Y2=0
cc_112 N_A_88_187#_c_72_n N_VPWR_c_320_n 0.0337695f $X=2.09 $Y=2.62 $X2=0 $Y2=0
cc_113 N_A_88_187#_c_109_p N_VPWR_c_320_n 0.00132454f $X=0.715 $Y=2.62 $X2=0
+ $Y2=0
cc_114 N_A_88_187#_c_102_p N_VPWR_c_320_n 0.00760156f $X=2.195 $Y=2.82 $X2=0
+ $Y2=0
cc_115 N_A_88_187#_c_72_n A_339_535# 0.00165214f $X=2.09 $Y=2.62 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A_88_187#_c_67_n N_VGND_M1002_d 0.00280695f $X=1.67 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_88_187#_c_108_p N_VGND_M1002_d 4.79672e-19 $X=0.715 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_88_187#_c_66_n N_VGND_c_366_n 8.05468e-19 $X=0.63 $Y=1.1 $X2=0 $Y2=0
cc_119 N_A_88_187#_c_67_n N_VGND_c_366_n 0.0199847f $X=1.67 $Y=0.9 $X2=0 $Y2=0
cc_120 N_A_88_187#_c_108_p N_VGND_c_366_n 0.00361359f $X=0.715 $Y=0.9 $X2=0
+ $Y2=0
cc_121 N_A_88_187#_c_69_n N_VGND_c_366_n 0.00525079f $X=0.617 $Y=0.935 $X2=0
+ $Y2=0
cc_122 N_A_88_187#_c_67_n N_VGND_c_371_n 0.00790195f $X=1.67 $Y=0.9 $X2=0 $Y2=0
cc_123 N_A_88_187#_c_108_p N_VGND_c_371_n 0.00424573f $X=0.715 $Y=0.9 $X2=0
+ $Y2=0
cc_124 N_A_88_187#_c_69_n N_VGND_c_371_n 0.00534666f $X=0.617 $Y=0.935 $X2=0
+ $Y2=0
cc_125 N_A_88_187#_c_69_n N_VGND_c_372_n 0.00548357f $X=0.617 $Y=0.935 $X2=0
+ $Y2=0
cc_126 N_A_88_187#_c_67_n N_A_237_81#_M1007_d 0.00263553f $X=1.67 $Y=0.9
+ $X2=-0.19 $Y2=-0.245
cc_127 N_A_88_187#_M1008_d N_A_237_81#_c_404_n 0.00180746f $X=1.695 $Y=0.405
+ $X2=0 $Y2=0
cc_128 N_A_88_187#_c_67_n N_A_237_81#_c_404_n 0.00383775f $X=1.67 $Y=0.9 $X2=0
+ $Y2=0
cc_129 N_A_88_187#_c_68_n N_A_237_81#_c_404_n 0.0145548f $X=1.835 $Y=0.7 $X2=0
+ $Y2=0
cc_130 N_A_88_187#_c_67_n N_A_237_81#_c_405_n 0.0192949f $X=1.67 $Y=0.9 $X2=0
+ $Y2=0
cc_131 N_A1_M1007_g N_B1_M1008_g 0.0215974f $X=1.11 $Y=0.615 $X2=0 $Y2=0
cc_132 N_A1_c_143_n N_B1_M1008_g 0.0131881f $X=2.885 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A1_c_160_n N_B1_M1008_g 0.00238428f $X=1.17 $Y=1.25 $X2=0 $Y2=0
cc_134 N_A1_c_144_n N_B1_M1008_g 0.0439966f $X=1.17 $Y=1.25 $X2=0 $Y2=0
cc_135 N_A1_c_143_n N_B1_c_202_n 0.00663531f $X=2.885 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A1_c_160_n N_B1_c_202_n 9.40141e-19 $X=1.17 $Y=1.25 $X2=0 $Y2=0
cc_137 N_A1_c_144_n N_B1_c_202_n 0.0177996f $X=1.17 $Y=1.25 $X2=0 $Y2=0
cc_138 N_A1_c_160_n B1 0.00974616f $X=1.17 $Y=1.25 $X2=0 $Y2=0
cc_139 N_A1_c_144_n B1 0.00130935f $X=1.17 $Y=1.25 $X2=0 $Y2=0
cc_140 N_A1_c_143_n N_B2_M1009_g 0.0148057f $X=2.885 $Y=1.58 $X2=0 $Y2=0
cc_141 N_A1_c_143_n B2 0.0484228f $X=2.885 $Y=1.58 $X2=0 $Y2=0
cc_142 A1 B2 0.0154556f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_143 N_A1_c_143_n N_B2_c_243_n 0.00512677f $X=2.885 $Y=1.58 $X2=0 $Y2=0
cc_144 N_A1_c_143_n N_A2_c_271_n 0.0051706f $X=2.885 $Y=1.58 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A1_c_146_n N_A2_c_271_n 2.75264e-19 $X=2.97 $Y=1.82 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A1_c_143_n N_A2_M1006_g 0.0186283f $X=2.885 $Y=1.58 $X2=0 $Y2=0
cc_147 A1 N_A2_M1006_g 0.00342252f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A1_c_146_n N_A2_M1006_g 0.0984597f $X=2.97 $Y=1.82 $X2=0 $Y2=0
cc_149 N_A1_c_143_n A2 0.0191161f $X=2.885 $Y=1.58 $X2=0 $Y2=0
cc_150 A1 A2 0.0186911f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A1_c_146_n A2 0.00160081f $X=2.97 $Y=1.82 $X2=0 $Y2=0
cc_152 N_A1_M1005_g N_VPWR_c_323_n 0.010878f $X=2.88 $Y=2.885 $X2=0 $Y2=0
cc_153 N_A1_c_148_n N_VPWR_c_323_n 7.57551e-19 $X=2.97 $Y=2.325 $X2=0 $Y2=0
cc_154 A1 N_VPWR_c_323_n 0.0111823f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A1_M1005_g N_VPWR_c_325_n 0.00486043f $X=2.88 $Y=2.885 $X2=0 $Y2=0
cc_156 N_A1_M1005_g N_VPWR_c_320_n 0.00685218f $X=2.88 $Y=2.885 $X2=0 $Y2=0
cc_157 A1 N_VPWR_c_320_n 0.00289837f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A1_M1007_g N_VGND_c_366_n 0.00258275f $X=1.11 $Y=0.615 $X2=0 $Y2=0
cc_159 N_A1_M1007_g N_VGND_c_368_n 0.00478816f $X=1.11 $Y=0.615 $X2=0 $Y2=0
cc_160 N_A1_M1007_g N_VGND_c_371_n 0.0044912f $X=1.11 $Y=0.615 $X2=0 $Y2=0
cc_161 N_A1_M1007_g N_A_237_81#_c_405_n 0.00605605f $X=1.11 $Y=0.615 $X2=0 $Y2=0
cc_162 N_B1_M1008_g N_B2_M1009_g 0.0548731f $X=1.62 $Y=0.615 $X2=0 $Y2=0
cc_163 N_B1_c_203_n N_B2_c_240_n 0.0317823f $X=1.62 $Y=2.16 $X2=0 $Y2=0
cc_164 N_B1_M1004_g N_B2_c_241_n 0.0317823f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_165 N_B1_M1008_g B2 0.00916098f $X=1.62 $Y=0.615 $X2=0 $Y2=0
cc_166 N_B1_M1004_g B2 0.00321112f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_167 N_B1_c_203_n B2 0.0127627f $X=1.62 $Y=2.16 $X2=0 $Y2=0
cc_168 B1 B2 0.0177075f $X=1.115 $Y=1.95 $X2=0 $Y2=0
cc_169 N_B1_M1008_g N_B2_c_243_n 0.0317823f $X=1.62 $Y=0.615 $X2=0 $Y2=0
cc_170 N_B1_M1004_g N_VPWR_c_321_n 0.00621833f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_171 N_B1_M1004_g N_VPWR_c_325_n 0.0042361f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_172 N_B1_M1004_g N_VPWR_c_320_n 0.00723233f $X=1.62 $Y=2.885 $X2=0 $Y2=0
cc_173 N_B1_M1008_g N_VGND_c_368_n 9.29198e-19 $X=1.62 $Y=0.615 $X2=0 $Y2=0
cc_174 N_B1_M1008_g N_A_237_81#_c_404_n 0.0102179f $X=1.62 $Y=0.615 $X2=0 $Y2=0
cc_175 N_B1_M1008_g N_A_237_81#_c_405_n 3.90742e-19 $X=1.62 $Y=0.615 $X2=0 $Y2=0
cc_176 N_B2_M1009_g N_A2_c_271_n 0.0200392f $X=2.05 $Y=0.615 $X2=-0.19
+ $Y2=-0.245
cc_177 N_B2_M1001_g N_A2_M1006_g 0.0187329f $X=1.98 $Y=2.885 $X2=0 $Y2=0
cc_178 B2 N_A2_M1006_g 0.0057391f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_179 N_B2_c_243_n N_A2_M1006_g 0.041097f $X=2.07 $Y=1.93 $X2=0 $Y2=0
cc_180 N_B2_M1009_g N_A2_c_273_n 0.0275678f $X=2.05 $Y=0.615 $X2=0 $Y2=0
cc_181 N_B2_M1009_g A2 0.00170453f $X=2.05 $Y=0.615 $X2=0 $Y2=0
cc_182 N_B2_M1001_g N_VPWR_c_325_n 0.0042361f $X=1.98 $Y=2.885 $X2=0 $Y2=0
cc_183 N_B2_M1001_g N_VPWR_c_320_n 0.00612074f $X=1.98 $Y=2.885 $X2=0 $Y2=0
cc_184 N_B2_M1009_g N_VGND_c_368_n 9.29198e-19 $X=2.05 $Y=0.615 $X2=0 $Y2=0
cc_185 N_B2_M1009_g N_A_237_81#_c_404_n 0.0131325f $X=2.05 $Y=0.615 $X2=0 $Y2=0
cc_186 N_B2_M1009_g N_A_237_81#_c_406_n 3.90742e-19 $X=2.05 $Y=0.615 $X2=0 $Y2=0
cc_187 N_A2_M1006_g N_VPWR_c_323_n 0.00209922f $X=2.52 $Y=2.885 $X2=0 $Y2=0
cc_188 N_A2_M1006_g N_VPWR_c_325_n 0.00585385f $X=2.52 $Y=2.885 $X2=0 $Y2=0
cc_189 N_A2_M1006_g N_VPWR_c_320_n 0.011101f $X=2.52 $Y=2.885 $X2=0 $Y2=0
cc_190 N_A2_c_271_n N_VGND_c_367_n 7.69862e-19 $X=2.52 $Y=1.445 $X2=0 $Y2=0
cc_191 N_A2_c_273_n N_VGND_c_367_n 0.00771883f $X=2.56 $Y=0.935 $X2=0 $Y2=0
cc_192 A2 N_VGND_c_367_n 0.0260407f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_193 N_A2_c_273_n N_VGND_c_368_n 0.00478816f $X=2.56 $Y=0.935 $X2=0 $Y2=0
cc_194 N_A2_c_273_n N_VGND_c_371_n 0.0044912f $X=2.56 $Y=0.935 $X2=0 $Y2=0
cc_195 A2 N_VGND_c_371_n 0.0143029f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_196 N_A2_c_273_n N_A_237_81#_c_406_n 0.00640878f $X=2.56 $Y=0.935 $X2=0 $Y2=0
cc_197 A2 N_A_237_81#_c_406_n 0.0016295f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_198 X N_VPWR_c_321_n 0.0066518f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_199 X N_VPWR_c_324_n 0.00990143f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_200 N_X_M1000_s N_VPWR_c_320_n 0.00503412f $X=0.155 $Y=2.675 $X2=0 $Y2=0
cc_201 X N_VPWR_c_320_n 0.00826079f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_202 N_X_c_305_n N_VGND_c_371_n 0.0112216f $X=0.305 $Y=0.55 $X2=0 $Y2=0
cc_203 N_X_c_305_n N_VGND_c_372_n 0.00929899f $X=0.305 $Y=0.55 $X2=0 $Y2=0
cc_204 N_VPWR_c_320_n A_339_535# 0.00241193f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_205 N_VPWR_c_320_n A_519_535# 0.00899413f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_206 N_VGND_c_368_n N_A_237_81#_c_404_n 0.0418379f $X=2.69 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_c_371_n N_A_237_81#_c_404_n 0.0257875f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_208 N_VGND_c_366_n N_A_237_81#_c_405_n 0.0188574f $X=0.815 $Y=0.53 $X2=0
+ $Y2=0
cc_209 N_VGND_c_368_n N_A_237_81#_c_405_n 0.0211423f $X=2.69 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_371_n N_A_237_81#_c_405_n 0.0124918f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_367_n N_A_237_81#_c_406_n 0.0195743f $X=2.855 $Y=0.55 $X2=0
+ $Y2=0
cc_212 N_VGND_c_368_n N_A_237_81#_c_406_n 0.021223f $X=2.69 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_c_371_n N_A_237_81#_c_406_n 0.0125082f $X=3.12 $Y=0 $X2=0 $Y2=0
