* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__iso0p_lp A KAPWR SLEEP VGND VNB VPB VPWR X
X0 a_342_489# A a_432_489# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND a_342_489# a_602_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_112_93# SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_27_93# SLEEP a_112_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_112_489# SLEEP KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_27_93# SLEEP a_112_489# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND a_27_93# a_340_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 KAPWR a_342_489# a_602_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_602_367# a_342_489# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_432_489# A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_340_93# A a_342_489# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 KAPWR a_27_93# a_270_489# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 a_270_489# a_27_93# a_342_489# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_602_93# a_342_489# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
