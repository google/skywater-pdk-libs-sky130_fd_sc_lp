* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fahcin_1 A B CIN VGND VNB VPB VPWR COUT SUM
X0 a_1883_395# a_1774_367# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 VGND CIN a_1774_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND a_1926_135# SUM VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND a_439_47# a_1152_389# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_1152_389# a_364_73# COUT VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 VPWR a_1926_135# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND a_29_47# a_256_87# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 a_439_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_1883_395# a_555_73# a_1926_135# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X9 a_29_47# B a_364_73# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 COUT a_555_73# a_1500_63# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_256_87# B a_555_73# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 a_1883_395# a_1774_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X13 a_364_73# a_439_47# a_256_87# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 a_1926_135# a_364_73# a_1774_367# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 a_555_73# a_439_47# a_29_47# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 a_29_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_256_87# B a_364_73# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_1500_63# CIN VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X19 a_1774_367# a_555_73# a_1926_135# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X20 COUT a_364_73# a_1500_63# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_1500_63# CIN VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_29_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_1926_135# a_364_73# a_1883_395# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 a_439_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_364_73# a_439_47# a_29_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 a_1152_389# a_555_73# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 a_29_47# B a_555_73# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 VPWR a_29_47# a_256_87# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X29 VPWR a_439_47# a_1152_389# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=150000u
X30 a_555_73# a_439_47# a_256_87# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X31 VPWR CIN a_1774_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
